module basic_1500_15000_2000_20_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_427,In_1140);
or U1 (N_1,In_167,In_526);
nand U2 (N_2,In_1463,In_1309);
and U3 (N_3,In_620,In_538);
nor U4 (N_4,In_1022,In_139);
xor U5 (N_5,In_602,In_295);
or U6 (N_6,In_240,In_97);
nor U7 (N_7,In_610,In_974);
and U8 (N_8,In_297,In_1385);
xor U9 (N_9,In_655,In_86);
or U10 (N_10,In_112,In_1497);
xor U11 (N_11,In_783,In_541);
or U12 (N_12,In_203,In_1203);
nand U13 (N_13,In_532,In_935);
or U14 (N_14,In_868,In_692);
nor U15 (N_15,In_233,In_521);
nand U16 (N_16,In_241,In_1173);
or U17 (N_17,In_817,In_424);
and U18 (N_18,In_570,In_821);
nand U19 (N_19,In_1165,In_291);
nor U20 (N_20,In_507,In_503);
nand U21 (N_21,In_1372,In_1186);
xor U22 (N_22,In_330,In_11);
xor U23 (N_23,In_1275,In_1093);
or U24 (N_24,In_172,In_451);
and U25 (N_25,In_966,In_1151);
nand U26 (N_26,In_1341,In_1109);
nand U27 (N_27,In_1192,In_211);
and U28 (N_28,In_740,In_66);
or U29 (N_29,In_1405,In_1284);
or U30 (N_30,In_511,In_769);
nor U31 (N_31,In_393,In_754);
nor U32 (N_32,In_844,In_148);
nand U33 (N_33,In_865,In_290);
nand U34 (N_34,In_1234,In_1236);
nand U35 (N_35,In_899,In_772);
nor U36 (N_36,In_1101,In_617);
or U37 (N_37,In_59,In_851);
or U38 (N_38,In_442,In_711);
xnor U39 (N_39,In_1412,In_471);
xor U40 (N_40,In_593,In_1200);
nand U41 (N_41,In_447,In_50);
or U42 (N_42,In_640,In_1273);
nand U43 (N_43,In_1055,In_27);
nor U44 (N_44,In_748,In_993);
xnor U45 (N_45,In_260,In_971);
and U46 (N_46,In_320,In_637);
and U47 (N_47,In_1382,In_536);
and U48 (N_48,In_417,In_283);
xor U49 (N_49,In_625,In_1029);
xor U50 (N_50,In_1447,In_731);
and U51 (N_51,In_520,In_159);
and U52 (N_52,In_302,In_1313);
nor U53 (N_53,In_446,In_469);
nor U54 (N_54,In_1401,In_682);
and U55 (N_55,In_182,In_799);
nand U56 (N_56,In_1123,In_587);
or U57 (N_57,In_1061,In_616);
or U58 (N_58,In_292,In_1465);
xor U59 (N_59,In_43,In_516);
or U60 (N_60,In_365,In_143);
and U61 (N_61,In_550,In_399);
nor U62 (N_62,In_515,In_905);
and U63 (N_63,In_39,In_1128);
xnor U64 (N_64,In_867,In_857);
xnor U65 (N_65,In_254,In_646);
xor U66 (N_66,In_122,In_601);
and U67 (N_67,In_269,In_923);
xnor U68 (N_68,In_586,In_873);
nand U69 (N_69,In_29,In_577);
and U70 (N_70,In_954,In_621);
and U71 (N_71,In_886,In_1133);
nand U72 (N_72,In_457,In_1145);
nand U73 (N_73,In_443,In_1352);
xor U74 (N_74,In_657,In_1479);
nand U75 (N_75,In_1419,In_709);
xor U76 (N_76,In_359,In_1271);
or U77 (N_77,In_67,In_69);
or U78 (N_78,In_1446,In_354);
nor U79 (N_79,In_893,In_287);
nand U80 (N_80,In_1077,In_1159);
or U81 (N_81,In_1373,In_1097);
or U82 (N_82,In_1066,In_733);
or U83 (N_83,In_1265,In_774);
nand U84 (N_84,In_402,In_1499);
nand U85 (N_85,In_422,In_267);
xnor U86 (N_86,In_1119,In_480);
nor U87 (N_87,In_1364,In_1094);
nand U88 (N_88,In_832,In_209);
and U89 (N_89,In_357,In_942);
nor U90 (N_90,In_430,In_53);
or U91 (N_91,In_279,In_842);
or U92 (N_92,In_998,In_611);
or U93 (N_93,In_1310,In_543);
nand U94 (N_94,In_16,In_136);
or U95 (N_95,In_331,In_225);
nand U96 (N_96,In_1169,In_1116);
xor U97 (N_97,In_834,In_1168);
or U98 (N_98,In_607,In_40);
nand U99 (N_99,In_1289,In_723);
nor U100 (N_100,In_63,In_1449);
or U101 (N_101,In_1415,In_1464);
xor U102 (N_102,In_562,In_111);
or U103 (N_103,In_419,In_551);
nand U104 (N_104,In_699,In_1069);
nand U105 (N_105,In_401,In_118);
or U106 (N_106,In_168,In_544);
xor U107 (N_107,In_374,In_667);
and U108 (N_108,In_473,In_41);
or U109 (N_109,In_1392,In_797);
or U110 (N_110,In_724,In_1141);
nor U111 (N_111,In_679,In_1046);
or U112 (N_112,In_1179,In_528);
or U113 (N_113,In_56,In_1024);
and U114 (N_114,In_1067,In_1149);
or U115 (N_115,In_864,In_1411);
xor U116 (N_116,In_623,In_109);
nor U117 (N_117,In_1207,In_1166);
nand U118 (N_118,In_612,In_147);
or U119 (N_119,In_685,In_765);
xnor U120 (N_120,In_488,In_467);
or U121 (N_121,In_631,In_653);
nor U122 (N_122,In_1150,In_713);
nand U123 (N_123,In_1158,In_256);
nand U124 (N_124,In_12,In_956);
nand U125 (N_125,In_1276,In_89);
nor U126 (N_126,In_334,In_218);
xnor U127 (N_127,In_1295,In_925);
nand U128 (N_128,In_1065,In_948);
and U129 (N_129,In_924,In_1387);
nor U130 (N_130,In_243,In_1004);
nor U131 (N_131,In_1459,In_1117);
and U132 (N_132,In_798,In_1196);
nor U133 (N_133,In_767,In_512);
nand U134 (N_134,In_936,In_1335);
or U135 (N_135,In_1118,In_1072);
nand U136 (N_136,In_1181,In_4);
xor U137 (N_137,In_449,In_1305);
and U138 (N_138,In_455,In_785);
nor U139 (N_139,In_396,In_784);
or U140 (N_140,In_164,In_1322);
or U141 (N_141,In_888,In_92);
nand U142 (N_142,In_1190,In_549);
xor U143 (N_143,In_45,In_1374);
nor U144 (N_144,In_1349,In_1278);
or U145 (N_145,In_1362,In_337);
or U146 (N_146,In_1308,In_57);
xnor U147 (N_147,In_1453,In_1475);
nor U148 (N_148,In_47,In_1157);
nor U149 (N_149,In_335,In_1365);
and U150 (N_150,In_982,In_452);
nand U151 (N_151,In_296,In_406);
or U152 (N_152,In_665,In_1484);
nand U153 (N_153,In_613,In_930);
nand U154 (N_154,In_1327,In_1017);
or U155 (N_155,In_559,In_984);
nand U156 (N_156,In_445,In_453);
or U157 (N_157,In_683,In_1469);
nor U158 (N_158,In_1445,In_1442);
and U159 (N_159,In_989,In_1059);
and U160 (N_160,In_961,In_126);
nor U161 (N_161,In_1458,In_18);
or U162 (N_162,In_792,In_588);
xnor U163 (N_163,In_470,In_928);
or U164 (N_164,In_131,In_54);
nand U165 (N_165,In_1233,In_574);
xor U166 (N_166,In_1360,In_13);
and U167 (N_167,In_818,In_650);
nor U168 (N_168,In_931,In_594);
nor U169 (N_169,In_927,In_801);
nor U170 (N_170,In_554,In_1220);
nand U171 (N_171,In_1285,In_510);
xnor U172 (N_172,In_44,In_245);
nor U173 (N_173,In_1398,In_1481);
or U174 (N_174,In_1448,In_828);
or U175 (N_175,In_173,In_1433);
or U176 (N_176,In_812,In_663);
nor U177 (N_177,In_939,In_722);
xnor U178 (N_178,In_1494,In_329);
or U179 (N_179,In_542,In_975);
nor U180 (N_180,In_1267,In_686);
xor U181 (N_181,In_229,In_973);
or U182 (N_182,In_1098,In_691);
nor U183 (N_183,In_78,In_1120);
nand U184 (N_184,In_545,In_595);
nand U185 (N_185,In_1304,In_1461);
nor U186 (N_186,In_1016,In_94);
nand U187 (N_187,In_911,In_1015);
or U188 (N_188,In_1367,In_852);
xor U189 (N_189,In_555,In_1052);
and U190 (N_190,In_238,In_589);
nand U191 (N_191,In_835,In_130);
or U192 (N_192,In_407,In_450);
and U193 (N_193,In_1426,In_1368);
and U194 (N_194,In_1070,In_894);
nor U195 (N_195,In_166,In_1081);
xnor U196 (N_196,In_24,In_1430);
and U197 (N_197,In_48,In_432);
nand U198 (N_198,In_946,In_2);
or U199 (N_199,In_194,In_462);
or U200 (N_200,In_477,In_786);
and U201 (N_201,In_478,In_82);
or U202 (N_202,In_263,In_231);
xor U203 (N_203,In_1,In_1488);
and U204 (N_204,In_749,In_394);
or U205 (N_205,In_180,In_1131);
nor U206 (N_206,In_1455,In_1084);
xnor U207 (N_207,In_0,In_853);
nor U208 (N_208,In_1450,In_933);
nand U209 (N_209,In_1359,In_71);
or U210 (N_210,In_1251,In_741);
xnor U211 (N_211,In_776,In_1164);
xor U212 (N_212,In_1031,In_116);
xor U213 (N_213,In_1228,In_929);
and U214 (N_214,In_920,In_992);
or U215 (N_215,In_433,In_866);
or U216 (N_216,In_490,In_826);
nor U217 (N_217,In_556,In_855);
xnor U218 (N_218,In_977,In_494);
or U219 (N_219,In_1254,In_1418);
nor U220 (N_220,In_115,In_1229);
and U221 (N_221,In_88,In_305);
or U222 (N_222,In_1078,In_790);
nor U223 (N_223,In_360,In_106);
nor U224 (N_224,In_1299,In_23);
and U225 (N_225,In_522,In_1427);
and U226 (N_226,In_1237,In_157);
nand U227 (N_227,In_1377,In_339);
nor U228 (N_228,In_414,In_913);
and U229 (N_229,In_747,In_689);
or U230 (N_230,In_1205,In_802);
or U231 (N_231,In_1075,In_1347);
or U232 (N_232,In_1403,In_1354);
xnor U233 (N_233,In_197,In_117);
nor U234 (N_234,In_1040,In_65);
xor U235 (N_235,In_1184,In_1311);
xnor U236 (N_236,In_727,In_482);
and U237 (N_237,In_815,In_902);
or U238 (N_238,In_598,In_608);
nand U239 (N_239,In_1369,In_379);
nand U240 (N_240,In_878,In_495);
xnor U241 (N_241,In_10,In_1030);
or U242 (N_242,In_1246,In_560);
or U243 (N_243,In_1423,In_847);
xnor U244 (N_244,In_1180,In_531);
and U245 (N_245,In_1139,In_1495);
and U246 (N_246,In_435,In_1312);
or U247 (N_247,In_1036,In_1153);
nand U248 (N_248,In_1074,In_585);
nor U249 (N_249,In_196,In_805);
and U250 (N_250,In_273,In_1307);
or U251 (N_251,In_1413,In_395);
or U252 (N_252,In_1008,In_322);
nand U253 (N_253,In_1211,In_609);
or U254 (N_254,In_30,In_428);
xnor U255 (N_255,In_883,In_1079);
or U256 (N_256,In_1404,In_259);
and U257 (N_257,In_436,In_672);
and U258 (N_258,In_654,In_988);
nor U259 (N_259,In_850,In_1187);
nand U260 (N_260,In_1417,In_141);
and U261 (N_261,In_213,In_666);
xor U262 (N_262,In_872,In_439);
xor U263 (N_263,In_804,In_1210);
and U264 (N_264,In_61,In_1318);
nor U265 (N_265,In_487,In_8);
nor U266 (N_266,In_1073,In_176);
or U267 (N_267,In_696,In_349);
nor U268 (N_268,In_125,In_794);
xnor U269 (N_269,In_508,In_1435);
nor U270 (N_270,In_958,In_871);
xnor U271 (N_271,In_768,In_1255);
and U272 (N_272,In_1122,In_1294);
xnor U273 (N_273,In_1240,In_1356);
nand U274 (N_274,In_1248,In_158);
xor U275 (N_275,In_837,In_1006);
nor U276 (N_276,In_1226,In_807);
nand U277 (N_277,In_247,In_1344);
or U278 (N_278,In_1002,In_278);
nor U279 (N_279,In_372,In_412);
xor U280 (N_280,In_1332,In_1490);
or U281 (N_281,In_309,In_932);
xor U282 (N_282,In_1298,In_519);
or U283 (N_283,In_323,In_319);
nor U284 (N_284,In_1358,In_651);
nand U285 (N_285,In_145,In_721);
or U286 (N_286,In_3,In_781);
nand U287 (N_287,In_474,In_904);
nand U288 (N_288,In_969,In_373);
nand U289 (N_289,In_880,In_527);
nor U290 (N_290,In_1477,In_1345);
and U291 (N_291,In_1043,In_1202);
xnor U292 (N_292,In_622,In_846);
or U293 (N_293,In_1178,In_953);
xor U294 (N_294,In_963,In_250);
and U295 (N_295,In_1416,In_706);
nand U296 (N_296,In_1301,In_312);
and U297 (N_297,In_1452,In_645);
and U298 (N_298,In_1256,In_207);
and U299 (N_299,In_572,In_382);
nor U300 (N_300,In_940,In_193);
nor U301 (N_301,In_415,In_947);
nand U302 (N_302,In_1083,In_1491);
or U303 (N_303,In_1085,In_600);
xor U304 (N_304,In_811,In_1217);
xnor U305 (N_305,In_228,In_903);
nand U306 (N_306,In_1383,In_1134);
xor U307 (N_307,In_921,In_6);
nor U308 (N_308,In_1363,In_26);
and U309 (N_309,In_367,In_1410);
nand U310 (N_310,In_375,In_782);
xnor U311 (N_311,In_265,In_1371);
and U312 (N_312,In_552,In_1182);
nand U313 (N_313,In_328,In_701);
nor U314 (N_314,In_1071,In_534);
nand U315 (N_315,In_313,In_590);
nor U316 (N_316,In_491,In_624);
and U317 (N_317,In_985,In_479);
xnor U318 (N_318,In_918,In_1104);
or U319 (N_319,In_299,In_1489);
and U320 (N_320,In_1395,In_677);
and U321 (N_321,In_1253,In_113);
nor U322 (N_322,In_324,In_410);
or U323 (N_323,In_1247,In_142);
and U324 (N_324,In_648,In_1167);
and U325 (N_325,In_398,In_652);
and U326 (N_326,In_85,In_140);
xor U327 (N_327,In_286,In_189);
and U328 (N_328,In_567,In_1089);
nor U329 (N_329,In_1334,In_1482);
nor U330 (N_330,In_368,In_1223);
xnor U331 (N_331,In_1121,In_957);
nand U332 (N_332,In_205,In_1257);
and U333 (N_333,In_1346,In_997);
nor U334 (N_334,In_870,In_573);
or U335 (N_335,In_734,In_1486);
xnor U336 (N_336,In_237,In_514);
xor U337 (N_337,In_775,In_458);
or U338 (N_338,In_1470,In_77);
xor U339 (N_339,In_674,In_342);
or U340 (N_340,In_192,In_919);
nor U341 (N_341,In_579,In_275);
nand U342 (N_342,In_178,In_914);
xor U343 (N_343,In_981,In_1214);
xnor U344 (N_344,In_1467,In_1431);
nor U345 (N_345,In_1056,In_738);
and U346 (N_346,In_539,In_1054);
nand U347 (N_347,In_1350,In_144);
nand U348 (N_348,In_1033,In_19);
nand U349 (N_349,In_1460,In_156);
nor U350 (N_350,In_763,In_1393);
or U351 (N_351,In_1397,In_1326);
nand U352 (N_352,In_1286,In_1197);
xnor U353 (N_353,In_163,In_1025);
xnor U354 (N_354,In_889,In_100);
and U355 (N_355,In_1476,In_162);
nor U356 (N_356,In_638,In_315);
nor U357 (N_357,In_806,In_848);
nand U358 (N_358,In_170,In_370);
nor U359 (N_359,In_174,In_860);
nand U360 (N_360,In_459,In_606);
nand U361 (N_361,In_673,In_796);
nand U362 (N_362,In_1297,In_661);
xnor U363 (N_363,In_725,In_1227);
xnor U364 (N_364,In_366,In_1045);
or U365 (N_365,In_177,In_1394);
and U366 (N_366,In_808,In_1018);
nand U367 (N_367,In_348,In_810);
nor U368 (N_368,In_108,In_153);
nor U369 (N_369,In_149,In_440);
and U370 (N_370,In_183,In_55);
nand U371 (N_371,In_475,In_1408);
xnor U372 (N_372,In_390,In_578);
or U373 (N_373,In_759,In_1296);
nor U374 (N_374,In_690,In_1142);
nor U375 (N_375,In_950,In_1336);
nand U376 (N_376,In_823,In_1343);
or U377 (N_377,In_463,In_687);
nor U378 (N_378,In_659,In_675);
xnor U379 (N_379,In_1216,In_1424);
xnor U380 (N_380,In_1287,In_425);
and U381 (N_381,In_951,In_1272);
xnor U382 (N_382,In_1132,In_1050);
or U383 (N_383,In_1241,In_962);
and U384 (N_384,In_750,In_897);
nand U385 (N_385,In_970,In_1238);
nor U386 (N_386,In_434,In_592);
and U387 (N_387,In_1155,In_755);
and U388 (N_388,In_1007,In_107);
nor U389 (N_389,In_224,In_730);
or U390 (N_390,In_1047,In_346);
nand U391 (N_391,In_1357,In_703);
nand U392 (N_392,In_210,In_84);
nor U393 (N_393,In_845,In_444);
nand U394 (N_394,In_1468,In_380);
nand U395 (N_395,In_591,In_1474);
or U396 (N_396,In_972,In_548);
nor U397 (N_397,In_403,In_517);
xnor U398 (N_398,In_1086,In_70);
and U399 (N_399,In_1269,In_1201);
or U400 (N_400,In_1351,In_1172);
or U401 (N_401,In_244,In_825);
nand U402 (N_402,In_952,In_627);
xor U403 (N_403,In_378,In_413);
or U404 (N_404,In_246,In_202);
xor U405 (N_405,In_1434,In_28);
nor U406 (N_406,In_770,In_119);
xor U407 (N_407,In_49,In_766);
and U408 (N_408,In_1090,In_1390);
nor U409 (N_409,In_1080,In_1111);
nand U410 (N_410,In_658,In_191);
xor U411 (N_411,In_1259,In_1021);
xnor U412 (N_412,In_662,In_165);
nor U413 (N_413,In_264,In_17);
nor U414 (N_414,In_1429,In_344);
nand U415 (N_415,In_1191,In_876);
and U416 (N_416,In_1028,In_926);
or U417 (N_417,In_1127,In_483);
xnor U418 (N_418,In_1399,In_881);
or U419 (N_419,In_1193,In_756);
and U420 (N_420,In_1137,In_1496);
and U421 (N_421,In_212,In_814);
or U422 (N_422,In_1044,In_1130);
xnor U423 (N_423,In_856,In_219);
or U424 (N_424,In_304,In_1420);
nor U425 (N_425,In_779,In_251);
and U426 (N_426,In_788,In_294);
xnor U427 (N_427,In_188,In_793);
or U428 (N_428,In_708,In_676);
nor U429 (N_429,In_861,In_46);
and U430 (N_430,In_137,In_1019);
xor U431 (N_431,In_1406,In_1438);
xnor U432 (N_432,In_656,In_93);
or U433 (N_433,In_227,In_288);
and U434 (N_434,In_890,In_420);
and U435 (N_435,In_1027,In_381);
xnor U436 (N_436,In_1068,In_751);
xnor U437 (N_437,In_1208,In_146);
xnor U438 (N_438,In_87,In_917);
nand U439 (N_439,In_91,In_698);
and U440 (N_440,In_341,In_276);
nor U441 (N_441,In_604,In_1219);
or U442 (N_442,In_960,In_1051);
or U443 (N_443,In_1270,In_736);
nand U444 (N_444,In_680,In_1041);
nand U445 (N_445,In_615,In_639);
nand U446 (N_446,In_79,In_1319);
nor U447 (N_447,In_582,In_105);
nor U448 (N_448,In_1260,In_300);
and U449 (N_449,In_820,In_1148);
and U450 (N_450,In_485,In_274);
nand U451 (N_451,In_1092,In_518);
nor U452 (N_452,In_190,In_764);
or U453 (N_453,In_132,In_397);
or U454 (N_454,In_1386,In_1038);
nand U455 (N_455,In_1136,In_1473);
or U456 (N_456,In_649,In_1035);
nand U457 (N_457,In_484,In_513);
nor U458 (N_458,In_314,In_1493);
and U459 (N_459,In_34,In_987);
nand U460 (N_460,In_90,In_744);
or U461 (N_461,In_1388,In_1243);
and U462 (N_462,In_581,In_1096);
nor U463 (N_463,In_910,In_1242);
nor U464 (N_464,In_1320,In_333);
and U465 (N_465,In_757,In_753);
or U466 (N_466,In_762,In_862);
nor U467 (N_467,In_760,In_558);
and U468 (N_468,In_745,In_102);
xor U469 (N_469,In_448,In_1457);
and U470 (N_470,In_1099,In_795);
nand U471 (N_471,In_1177,In_185);
nand U472 (N_472,In_277,In_1189);
nor U473 (N_473,In_1402,In_25);
xor U474 (N_474,In_206,In_1231);
or U475 (N_475,In_849,In_599);
or U476 (N_476,In_841,In_829);
or U477 (N_477,In_892,In_1209);
or U478 (N_478,In_1340,In_678);
nand U479 (N_479,In_7,In_614);
or U480 (N_480,In_391,In_38);
and U481 (N_481,In_1293,In_150);
and U482 (N_482,In_803,In_1466);
xnor U483 (N_483,In_1280,In_411);
nor U484 (N_484,In_21,In_1389);
or U485 (N_485,In_822,In_493);
nand U486 (N_486,In_874,In_752);
and U487 (N_487,In_280,In_1001);
nand U488 (N_488,In_1183,In_1268);
nor U489 (N_489,In_347,In_629);
nand U490 (N_490,In_68,In_882);
xnor U491 (N_491,In_1443,In_110);
nand U492 (N_492,In_839,In_80);
nor U493 (N_493,In_289,In_400);
or U494 (N_494,In_120,In_1300);
or U495 (N_495,In_773,In_1105);
nand U496 (N_496,In_496,In_937);
or U497 (N_497,In_199,In_771);
and U498 (N_498,In_1384,In_272);
nor U499 (N_499,In_1005,In_1391);
or U500 (N_500,In_934,In_813);
xor U501 (N_501,In_1348,In_743);
nand U502 (N_502,In_900,In_1215);
or U503 (N_503,In_502,In_1471);
xnor U504 (N_504,In_1199,In_941);
xor U505 (N_505,In_311,In_1281);
nor U506 (N_506,In_843,In_628);
or U507 (N_507,In_409,In_885);
xnor U508 (N_508,In_719,In_418);
xnor U509 (N_509,In_1436,In_20);
nand U510 (N_510,In_181,In_500);
nor U511 (N_511,In_995,In_1325);
or U512 (N_512,In_325,In_863);
nor U513 (N_513,In_9,In_1135);
or U514 (N_514,In_317,In_1212);
nand U515 (N_515,In_1370,In_376);
nand U516 (N_516,In_332,In_1113);
or U517 (N_517,In_1409,In_1026);
or U518 (N_518,In_979,In_1222);
nand U519 (N_519,In_630,In_501);
nor U520 (N_520,In_98,In_634);
nor U521 (N_521,In_670,In_831);
xor U522 (N_522,In_1487,In_99);
and U523 (N_523,In_76,In_52);
and U524 (N_524,In_566,In_859);
and U525 (N_525,In_887,In_257);
nand U526 (N_526,In_535,In_1198);
nand U527 (N_527,In_1302,In_1485);
and U528 (N_528,In_1143,In_1014);
or U529 (N_529,In_266,In_643);
and U530 (N_530,In_707,In_336);
xor U531 (N_531,In_234,In_1154);
and U532 (N_532,In_605,In_1088);
or U533 (N_533,In_704,In_1264);
nand U534 (N_534,In_389,In_64);
nor U535 (N_535,In_363,In_429);
nand U536 (N_536,In_1010,In_580);
nor U537 (N_537,In_547,In_1342);
or U538 (N_538,In_1441,In_597);
and U539 (N_539,In_705,In_356);
xnor U540 (N_540,In_103,In_1174);
nand U541 (N_541,In_476,In_208);
xnor U542 (N_542,In_1376,In_262);
and U543 (N_543,In_1058,In_565);
or U544 (N_544,In_1012,In_456);
nand U545 (N_545,In_1218,In_1023);
xnor U546 (N_546,In_1396,In_529);
nand U547 (N_547,In_42,In_1353);
and U548 (N_548,In_619,In_1125);
or U549 (N_549,In_1162,In_990);
nor U550 (N_550,In_1279,In_1091);
xnor U551 (N_551,In_1003,In_668);
xnor U552 (N_552,In_777,In_498);
nand U553 (N_553,In_1361,In_355);
and U554 (N_554,In_780,In_282);
nand U555 (N_555,In_114,In_293);
or U556 (N_556,In_854,In_1282);
xnor U557 (N_557,In_1252,In_216);
and U558 (N_558,In_664,In_60);
and U559 (N_559,In_345,In_492);
or U560 (N_560,In_352,In_466);
nor U561 (N_561,In_1274,In_468);
nor U562 (N_562,In_1103,In_1432);
xnor U563 (N_563,In_465,In_340);
nand U564 (N_564,In_1129,In_700);
and U565 (N_565,In_789,In_1032);
or U566 (N_566,In_732,In_220);
nand U567 (N_567,In_271,In_632);
xor U568 (N_568,In_1053,In_1483);
or U569 (N_569,In_201,In_169);
and U570 (N_570,In_255,In_1239);
nand U571 (N_571,In_633,In_1152);
nor U572 (N_572,In_746,In_426);
or U573 (N_573,In_200,In_726);
nor U574 (N_574,In_858,In_310);
nand U575 (N_575,In_1110,In_906);
and U576 (N_576,In_524,In_1328);
or U577 (N_577,In_1314,In_160);
xnor U578 (N_578,In_1291,In_1147);
xnor U579 (N_579,In_525,In_104);
or U580 (N_580,In_214,In_1338);
nand U581 (N_581,In_1020,In_235);
and U582 (N_582,In_833,In_499);
or U583 (N_583,In_1100,In_253);
or U584 (N_584,In_537,In_791);
and U585 (N_585,In_1263,In_1421);
or U586 (N_586,In_636,In_37);
nand U587 (N_587,In_1375,In_1306);
xnor U588 (N_588,In_239,In_307);
and U589 (N_589,In_184,In_1037);
xor U590 (N_590,In_489,In_73);
and U591 (N_591,In_1230,In_576);
or U592 (N_592,In_509,In_1454);
nor U593 (N_593,In_22,In_198);
and U594 (N_594,In_1175,In_133);
or U595 (N_595,In_15,In_405);
or U596 (N_596,In_761,In_1472);
nand U597 (N_597,In_530,In_252);
and U598 (N_598,In_879,In_955);
xnor U599 (N_599,In_408,In_964);
and U600 (N_600,In_568,In_1156);
and U601 (N_601,In_123,In_1124);
or U602 (N_602,In_75,In_1146);
or U603 (N_603,In_81,In_223);
and U604 (N_604,In_423,In_710);
nand U605 (N_605,In_1337,In_138);
and U606 (N_606,In_1425,In_1194);
or U607 (N_607,In_14,In_712);
xor U608 (N_608,In_124,In_351);
and U609 (N_609,In_626,In_230);
nand U610 (N_610,In_461,In_1266);
xor U611 (N_611,In_1204,In_1249);
nand U612 (N_612,In_702,In_1039);
nor U613 (N_613,In_717,In_569);
or U614 (N_614,In_1213,In_361);
nand U615 (N_615,In_1224,In_915);
nand U616 (N_616,In_1379,In_945);
nand U617 (N_617,In_1422,In_695);
and U618 (N_618,In_51,In_161);
xor U619 (N_619,In_460,In_171);
and U620 (N_620,In_996,In_681);
and U621 (N_621,In_1107,In_1235);
or U622 (N_622,In_809,In_306);
and U623 (N_623,In_1185,In_728);
nor U624 (N_624,In_175,In_1087);
xnor U625 (N_625,In_584,In_1317);
and U626 (N_626,In_965,In_1315);
xnor U627 (N_627,In_641,In_540);
or U628 (N_628,In_96,In_1057);
or U629 (N_629,In_35,In_303);
and U630 (N_630,In_1221,In_980);
nand U631 (N_631,In_36,In_1330);
or U632 (N_632,In_1331,In_1261);
and U633 (N_633,In_875,In_1108);
and U634 (N_634,In_481,In_404);
nand U635 (N_635,In_1414,In_800);
and U636 (N_636,In_1049,In_877);
xnor U637 (N_637,In_134,In_901);
or U638 (N_638,In_377,In_1333);
xor U639 (N_639,In_497,In_1492);
nor U640 (N_640,In_281,In_739);
nor U641 (N_641,In_431,In_222);
and U642 (N_642,In_912,In_261);
xnor U643 (N_643,In_338,In_1009);
nand U644 (N_644,In_129,In_1288);
xnor U645 (N_645,In_242,In_684);
xnor U646 (N_646,In_1176,In_1112);
or U647 (N_647,In_1063,In_991);
or U648 (N_648,In_316,In_392);
or U649 (N_649,In_1381,In_1076);
nand U650 (N_650,In_986,In_441);
or U651 (N_651,In_472,In_1262);
or U652 (N_652,In_644,In_660);
nor U653 (N_653,In_1355,In_505);
nor U654 (N_654,In_523,In_827);
nor U655 (N_655,In_838,In_1225);
or U656 (N_656,In_787,In_737);
nand U657 (N_657,In_1462,In_58);
nor U658 (N_658,In_1380,In_546);
and U659 (N_659,In_385,In_1245);
xnor U660 (N_660,In_83,In_301);
nand U661 (N_661,In_999,In_697);
xnor U662 (N_662,In_1437,In_557);
or U663 (N_663,In_186,In_95);
or U664 (N_664,In_824,In_1283);
and U665 (N_665,In_583,In_716);
nor U666 (N_666,In_1106,In_327);
xnor U667 (N_667,In_154,In_438);
xnor U668 (N_668,In_1250,In_308);
and U669 (N_669,In_386,In_285);
xor U670 (N_670,In_688,In_369);
or U671 (N_671,In_318,In_215);
nor U672 (N_672,In_350,In_729);
or U673 (N_673,In_909,In_1439);
or U674 (N_674,In_694,In_1171);
xnor U675 (N_675,In_869,In_561);
nor U676 (N_676,In_1366,In_1456);
and U677 (N_677,In_31,In_1138);
xnor U678 (N_678,In_693,In_1451);
xor U679 (N_679,In_715,In_1095);
or U680 (N_680,In_895,In_596);
nor U681 (N_681,In_101,In_635);
xnor U682 (N_682,In_916,In_1303);
nand U683 (N_683,In_1498,In_221);
nand U684 (N_684,In_384,In_284);
nor U685 (N_685,In_232,In_179);
and U686 (N_686,In_437,In_976);
nor U687 (N_687,In_504,In_236);
xnor U688 (N_688,In_758,In_1064);
nor U689 (N_689,In_938,In_454);
nand U690 (N_690,In_268,In_836);
and U691 (N_691,In_1000,In_618);
xnor U692 (N_692,In_647,In_195);
nand U693 (N_693,In_1480,In_152);
and U694 (N_694,In_249,In_563);
xor U695 (N_695,In_121,In_1060);
nand U696 (N_696,In_908,In_155);
or U697 (N_697,In_371,In_298);
or U698 (N_698,In_421,In_1034);
nand U699 (N_699,In_1048,In_416);
nor U700 (N_700,In_464,In_1163);
nand U701 (N_701,In_575,In_270);
nand U702 (N_702,In_1206,In_321);
and U703 (N_703,In_387,In_1290);
nand U704 (N_704,In_669,In_1339);
and U705 (N_705,In_1160,In_742);
xor U706 (N_706,In_1478,In_1292);
nor U707 (N_707,In_533,In_840);
and U708 (N_708,In_364,In_5);
xor U709 (N_709,In_959,In_1062);
or U710 (N_710,In_642,In_943);
xnor U711 (N_711,In_217,In_1042);
nand U712 (N_712,In_922,In_1277);
nor U713 (N_713,In_1324,In_714);
xor U714 (N_714,In_891,In_944);
or U715 (N_715,In_978,In_187);
xnor U716 (N_716,In_1011,In_720);
xnor U717 (N_717,In_898,In_1316);
nor U718 (N_718,In_33,In_258);
and U719 (N_719,In_1440,In_994);
nand U720 (N_720,In_571,In_353);
xnor U721 (N_721,In_907,In_819);
or U722 (N_722,In_74,In_1232);
and U723 (N_723,In_1114,In_1082);
nand U724 (N_724,In_1400,In_896);
nor U725 (N_725,In_1126,In_983);
nor U726 (N_726,In_778,In_603);
nor U727 (N_727,In_388,In_1444);
and U728 (N_728,In_564,In_248);
and U729 (N_729,In_486,In_718);
nor U730 (N_730,In_735,In_128);
xnor U731 (N_731,In_1115,In_1321);
xnor U732 (N_732,In_127,In_1329);
xor U733 (N_733,In_135,In_1323);
nor U734 (N_734,In_1013,In_1378);
or U735 (N_735,In_204,In_62);
or U736 (N_736,In_967,In_1258);
or U737 (N_737,In_72,In_1144);
xor U738 (N_738,In_830,In_1428);
or U739 (N_739,In_151,In_358);
xor U740 (N_740,In_968,In_383);
and U741 (N_741,In_326,In_884);
nor U742 (N_742,In_1170,In_343);
or U743 (N_743,In_1195,In_1188);
and U744 (N_744,In_1407,In_506);
nor U745 (N_745,In_32,In_362);
nand U746 (N_746,In_226,In_1161);
xnor U747 (N_747,In_1102,In_949);
nand U748 (N_748,In_671,In_816);
nor U749 (N_749,In_553,In_1244);
and U750 (N_750,N_366,N_694);
nand U751 (N_751,N_238,N_430);
xor U752 (N_752,N_535,N_434);
and U753 (N_753,N_66,N_254);
or U754 (N_754,N_656,N_168);
or U755 (N_755,N_641,N_41);
or U756 (N_756,N_745,N_147);
xor U757 (N_757,N_77,N_110);
and U758 (N_758,N_142,N_205);
xnor U759 (N_759,N_184,N_468);
nand U760 (N_760,N_637,N_732);
nor U761 (N_761,N_577,N_440);
nor U762 (N_762,N_335,N_355);
and U763 (N_763,N_331,N_385);
xnor U764 (N_764,N_558,N_10);
or U765 (N_765,N_653,N_394);
or U766 (N_766,N_396,N_740);
xnor U767 (N_767,N_138,N_616);
or U768 (N_768,N_199,N_292);
nand U769 (N_769,N_93,N_633);
xnor U770 (N_770,N_538,N_81);
nand U771 (N_771,N_129,N_201);
nand U772 (N_772,N_661,N_1);
nor U773 (N_773,N_164,N_483);
or U774 (N_774,N_617,N_230);
or U775 (N_775,N_622,N_84);
xnor U776 (N_776,N_223,N_329);
and U777 (N_777,N_166,N_314);
and U778 (N_778,N_175,N_576);
nor U779 (N_779,N_27,N_436);
xnor U780 (N_780,N_607,N_412);
or U781 (N_781,N_505,N_332);
or U782 (N_782,N_302,N_532);
or U783 (N_783,N_642,N_666);
and U784 (N_784,N_106,N_315);
or U785 (N_785,N_180,N_131);
nor U786 (N_786,N_118,N_156);
nor U787 (N_787,N_714,N_9);
nor U788 (N_788,N_197,N_425);
or U789 (N_789,N_219,N_120);
nor U790 (N_790,N_593,N_96);
and U791 (N_791,N_372,N_348);
or U792 (N_792,N_479,N_159);
nor U793 (N_793,N_549,N_744);
and U794 (N_794,N_313,N_370);
or U795 (N_795,N_361,N_588);
and U796 (N_796,N_431,N_534);
or U797 (N_797,N_171,N_403);
nor U798 (N_798,N_566,N_650);
and U799 (N_799,N_251,N_570);
nand U800 (N_800,N_443,N_13);
and U801 (N_801,N_452,N_733);
nand U802 (N_802,N_352,N_350);
or U803 (N_803,N_212,N_679);
nand U804 (N_804,N_516,N_560);
nor U805 (N_805,N_420,N_50);
or U806 (N_806,N_343,N_83);
xnor U807 (N_807,N_723,N_513);
nor U808 (N_808,N_736,N_377);
xor U809 (N_809,N_132,N_317);
or U810 (N_810,N_126,N_725);
xnor U811 (N_811,N_579,N_231);
nand U812 (N_812,N_398,N_508);
or U813 (N_813,N_260,N_305);
nand U814 (N_814,N_554,N_94);
nand U815 (N_815,N_316,N_218);
xnor U816 (N_816,N_409,N_433);
nor U817 (N_817,N_493,N_470);
nand U818 (N_818,N_486,N_457);
and U819 (N_819,N_269,N_288);
nor U820 (N_820,N_44,N_550);
nor U821 (N_821,N_676,N_621);
and U822 (N_822,N_211,N_609);
and U823 (N_823,N_318,N_151);
or U824 (N_824,N_278,N_682);
nor U825 (N_825,N_545,N_346);
and U826 (N_826,N_191,N_704);
and U827 (N_827,N_428,N_614);
nand U828 (N_828,N_24,N_178);
nand U829 (N_829,N_451,N_186);
nand U830 (N_830,N_222,N_333);
or U831 (N_831,N_562,N_606);
xnor U832 (N_832,N_46,N_737);
nor U833 (N_833,N_225,N_14);
or U834 (N_834,N_441,N_369);
and U835 (N_835,N_338,N_308);
and U836 (N_836,N_686,N_490);
xor U837 (N_837,N_456,N_651);
xor U838 (N_838,N_306,N_638);
or U839 (N_839,N_31,N_183);
nor U840 (N_840,N_255,N_37);
nand U841 (N_841,N_665,N_748);
or U842 (N_842,N_639,N_80);
nand U843 (N_843,N_735,N_192);
nand U844 (N_844,N_39,N_494);
and U845 (N_845,N_446,N_38);
and U846 (N_846,N_210,N_234);
and U847 (N_847,N_283,N_537);
nand U848 (N_848,N_585,N_613);
and U849 (N_849,N_675,N_154);
or U850 (N_850,N_224,N_7);
nor U851 (N_851,N_277,N_561);
xor U852 (N_852,N_424,N_499);
or U853 (N_853,N_271,N_23);
and U854 (N_854,N_163,N_485);
nand U855 (N_855,N_357,N_444);
xnor U856 (N_856,N_109,N_381);
nor U857 (N_857,N_722,N_134);
nand U858 (N_858,N_365,N_108);
or U859 (N_859,N_730,N_86);
or U860 (N_860,N_123,N_586);
xnor U861 (N_861,N_18,N_401);
and U862 (N_862,N_26,N_741);
nand U863 (N_863,N_276,N_360);
or U864 (N_864,N_204,N_453);
and U865 (N_865,N_474,N_598);
nand U866 (N_866,N_179,N_530);
xnor U867 (N_867,N_703,N_517);
or U868 (N_868,N_673,N_388);
nand U869 (N_869,N_267,N_423);
or U870 (N_870,N_429,N_232);
nor U871 (N_871,N_475,N_290);
nand U872 (N_872,N_248,N_282);
and U873 (N_873,N_689,N_359);
nor U874 (N_874,N_632,N_189);
and U875 (N_875,N_196,N_678);
xor U876 (N_876,N_239,N_557);
xnor U877 (N_877,N_491,N_578);
nor U878 (N_878,N_71,N_472);
nor U879 (N_879,N_62,N_384);
nor U880 (N_880,N_198,N_459);
and U881 (N_881,N_91,N_477);
or U882 (N_882,N_705,N_649);
and U883 (N_883,N_629,N_297);
or U884 (N_884,N_400,N_663);
or U885 (N_885,N_130,N_630);
and U886 (N_886,N_258,N_228);
or U887 (N_887,N_20,N_563);
nor U888 (N_888,N_515,N_362);
nor U889 (N_889,N_571,N_15);
xor U890 (N_890,N_502,N_34);
xnor U891 (N_891,N_45,N_450);
nand U892 (N_892,N_683,N_146);
nand U893 (N_893,N_449,N_700);
and U894 (N_894,N_667,N_64);
and U895 (N_895,N_458,N_647);
and U896 (N_896,N_709,N_17);
xnor U897 (N_897,N_112,N_460);
and U898 (N_898,N_695,N_90);
nor U899 (N_899,N_136,N_553);
nor U900 (N_900,N_304,N_273);
nand U901 (N_901,N_322,N_482);
nand U902 (N_902,N_411,N_393);
nand U903 (N_903,N_35,N_662);
and U904 (N_904,N_243,N_265);
nor U905 (N_905,N_437,N_710);
or U906 (N_906,N_284,N_712);
nand U907 (N_907,N_303,N_610);
and U908 (N_908,N_575,N_699);
nand U909 (N_909,N_426,N_548);
xor U910 (N_910,N_655,N_674);
nor U911 (N_911,N_49,N_392);
xnor U912 (N_912,N_729,N_286);
nand U913 (N_913,N_263,N_702);
nor U914 (N_914,N_600,N_525);
and U915 (N_915,N_659,N_56);
and U916 (N_916,N_672,N_301);
xor U917 (N_917,N_552,N_325);
or U918 (N_918,N_153,N_547);
nor U919 (N_919,N_564,N_448);
and U920 (N_920,N_85,N_170);
nand U921 (N_921,N_105,N_719);
nand U922 (N_922,N_504,N_383);
or U923 (N_923,N_711,N_680);
nor U924 (N_924,N_79,N_88);
or U925 (N_925,N_349,N_312);
xnor U926 (N_926,N_162,N_668);
xor U927 (N_927,N_418,N_309);
nor U928 (N_928,N_272,N_221);
nand U929 (N_929,N_692,N_478);
xor U930 (N_930,N_531,N_287);
and U931 (N_931,N_155,N_467);
nor U932 (N_932,N_471,N_559);
nand U933 (N_933,N_480,N_684);
or U934 (N_934,N_496,N_185);
nand U935 (N_935,N_687,N_188);
or U936 (N_936,N_6,N_209);
or U937 (N_937,N_167,N_599);
or U938 (N_938,N_533,N_462);
nand U939 (N_939,N_595,N_353);
and U940 (N_940,N_492,N_693);
and U941 (N_941,N_128,N_8);
and U942 (N_942,N_127,N_611);
xnor U943 (N_943,N_567,N_102);
and U944 (N_944,N_701,N_405);
nor U945 (N_945,N_296,N_364);
and U946 (N_946,N_82,N_635);
or U947 (N_947,N_55,N_169);
nand U948 (N_948,N_61,N_217);
nor U949 (N_949,N_351,N_310);
nand U950 (N_950,N_519,N_368);
or U951 (N_951,N_643,N_664);
xnor U952 (N_952,N_395,N_447);
and U953 (N_953,N_603,N_715);
xnor U954 (N_954,N_69,N_40);
nand U955 (N_955,N_195,N_30);
and U956 (N_956,N_582,N_21);
nand U957 (N_957,N_341,N_98);
or U958 (N_958,N_226,N_261);
or U959 (N_959,N_580,N_518);
nor U960 (N_960,N_319,N_465);
and U961 (N_961,N_640,N_503);
or U962 (N_962,N_374,N_63);
nand U963 (N_963,N_73,N_237);
xor U964 (N_964,N_140,N_371);
nor U965 (N_965,N_115,N_631);
or U966 (N_966,N_543,N_65);
nand U967 (N_967,N_207,N_696);
nand U968 (N_968,N_404,N_618);
nand U969 (N_969,N_568,N_54);
or U970 (N_970,N_125,N_143);
and U971 (N_971,N_107,N_363);
or U972 (N_972,N_121,N_501);
or U973 (N_973,N_241,N_644);
nand U974 (N_974,N_76,N_116);
nand U975 (N_975,N_193,N_605);
and U976 (N_976,N_731,N_337);
and U977 (N_977,N_47,N_187);
or U978 (N_978,N_572,N_660);
or U979 (N_979,N_620,N_122);
or U980 (N_980,N_245,N_52);
or U981 (N_981,N_11,N_262);
xnor U982 (N_982,N_367,N_594);
xnor U983 (N_983,N_53,N_509);
nand U984 (N_984,N_407,N_749);
or U985 (N_985,N_229,N_713);
nor U986 (N_986,N_546,N_438);
nand U987 (N_987,N_574,N_158);
nand U988 (N_988,N_5,N_399);
xor U989 (N_989,N_442,N_145);
and U990 (N_990,N_19,N_528);
or U991 (N_991,N_390,N_569);
or U992 (N_992,N_523,N_285);
nand U993 (N_993,N_624,N_58);
nor U994 (N_994,N_25,N_215);
nand U995 (N_995,N_133,N_173);
nor U996 (N_996,N_601,N_72);
xor U997 (N_997,N_336,N_149);
and U998 (N_998,N_615,N_101);
nand U999 (N_999,N_506,N_520);
and U1000 (N_1000,N_698,N_176);
xor U1001 (N_1001,N_32,N_628);
and U1002 (N_1002,N_657,N_74);
and U1003 (N_1003,N_268,N_59);
nor U1004 (N_1004,N_387,N_4);
xor U1005 (N_1005,N_500,N_320);
nand U1006 (N_1006,N_445,N_354);
xnor U1007 (N_1007,N_208,N_743);
xor U1008 (N_1008,N_148,N_742);
xor U1009 (N_1009,N_358,N_697);
and U1010 (N_1010,N_87,N_113);
and U1011 (N_1011,N_152,N_487);
xnor U1012 (N_1012,N_307,N_92);
nor U1013 (N_1013,N_249,N_75);
nor U1014 (N_1014,N_342,N_51);
nand U1015 (N_1015,N_619,N_78);
nand U1016 (N_1016,N_551,N_416);
xnor U1017 (N_1017,N_581,N_386);
nand U1018 (N_1018,N_608,N_669);
and U1019 (N_1019,N_300,N_590);
nand U1020 (N_1020,N_539,N_202);
and U1021 (N_1021,N_236,N_521);
nor U1022 (N_1022,N_565,N_227);
and U1023 (N_1023,N_334,N_589);
or U1024 (N_1024,N_144,N_60);
nor U1025 (N_1025,N_378,N_36);
or U1026 (N_1026,N_135,N_280);
and U1027 (N_1027,N_380,N_584);
or U1028 (N_1028,N_634,N_139);
or U1029 (N_1029,N_68,N_511);
nand U1030 (N_1030,N_321,N_541);
nand U1031 (N_1031,N_488,N_97);
and U1032 (N_1032,N_376,N_728);
xor U1033 (N_1033,N_495,N_489);
xnor U1034 (N_1034,N_252,N_356);
nand U1035 (N_1035,N_626,N_648);
xor U1036 (N_1036,N_327,N_275);
or U1037 (N_1037,N_422,N_264);
xnor U1038 (N_1038,N_244,N_279);
nor U1039 (N_1039,N_746,N_206);
nand U1040 (N_1040,N_691,N_658);
and U1041 (N_1041,N_734,N_213);
nor U1042 (N_1042,N_739,N_182);
xnor U1043 (N_1043,N_160,N_414);
or U1044 (N_1044,N_529,N_291);
xnor U1045 (N_1045,N_421,N_623);
xor U1046 (N_1046,N_645,N_95);
and U1047 (N_1047,N_281,N_165);
nand U1048 (N_1048,N_690,N_540);
and U1049 (N_1049,N_636,N_344);
and U1050 (N_1050,N_463,N_114);
or U1051 (N_1051,N_137,N_707);
nor U1052 (N_1052,N_671,N_339);
or U1053 (N_1053,N_597,N_544);
nor U1054 (N_1054,N_124,N_119);
nand U1055 (N_1055,N_382,N_726);
or U1056 (N_1056,N_612,N_413);
or U1057 (N_1057,N_330,N_514);
and U1058 (N_1058,N_573,N_161);
and U1059 (N_1059,N_246,N_242);
nor U1060 (N_1060,N_200,N_104);
xor U1061 (N_1061,N_720,N_2);
nand U1062 (N_1062,N_259,N_439);
or U1063 (N_1063,N_512,N_177);
and U1064 (N_1064,N_172,N_12);
nor U1065 (N_1065,N_727,N_294);
and U1066 (N_1066,N_587,N_627);
nor U1067 (N_1067,N_293,N_481);
xnor U1068 (N_1068,N_256,N_717);
nor U1069 (N_1069,N_625,N_716);
xnor U1070 (N_1070,N_295,N_604);
and U1071 (N_1071,N_432,N_375);
xor U1072 (N_1072,N_417,N_299);
or U1073 (N_1073,N_721,N_591);
xnor U1074 (N_1074,N_103,N_406);
or U1075 (N_1075,N_190,N_583);
nand U1076 (N_1076,N_326,N_435);
xnor U1077 (N_1077,N_270,N_454);
and U1078 (N_1078,N_289,N_253);
nand U1079 (N_1079,N_247,N_70);
nor U1080 (N_1080,N_194,N_117);
xor U1081 (N_1081,N_397,N_29);
xnor U1082 (N_1082,N_42,N_141);
and U1083 (N_1083,N_510,N_43);
and U1084 (N_1084,N_181,N_427);
and U1085 (N_1085,N_455,N_738);
and U1086 (N_1086,N_3,N_389);
or U1087 (N_1087,N_602,N_524);
or U1088 (N_1088,N_555,N_596);
nand U1089 (N_1089,N_33,N_100);
xor U1090 (N_1090,N_592,N_324);
and U1091 (N_1091,N_274,N_233);
and U1092 (N_1092,N_235,N_461);
and U1093 (N_1093,N_654,N_507);
nand U1094 (N_1094,N_340,N_379);
nand U1095 (N_1095,N_67,N_266);
nor U1096 (N_1096,N_22,N_476);
or U1097 (N_1097,N_718,N_527);
xor U1098 (N_1098,N_373,N_677);
nand U1099 (N_1099,N_174,N_298);
or U1100 (N_1100,N_542,N_150);
nand U1101 (N_1101,N_250,N_652);
xnor U1102 (N_1102,N_670,N_497);
and U1103 (N_1103,N_747,N_28);
and U1104 (N_1104,N_214,N_391);
xor U1105 (N_1105,N_203,N_688);
or U1106 (N_1106,N_16,N_706);
and U1107 (N_1107,N_257,N_419);
or U1108 (N_1108,N_473,N_0);
and U1109 (N_1109,N_402,N_311);
nor U1110 (N_1110,N_157,N_708);
xnor U1111 (N_1111,N_328,N_498);
nand U1112 (N_1112,N_240,N_556);
nand U1113 (N_1113,N_99,N_57);
and U1114 (N_1114,N_220,N_526);
nor U1115 (N_1115,N_111,N_323);
or U1116 (N_1116,N_681,N_89);
and U1117 (N_1117,N_464,N_484);
and U1118 (N_1118,N_48,N_646);
nor U1119 (N_1119,N_216,N_347);
and U1120 (N_1120,N_536,N_410);
xor U1121 (N_1121,N_415,N_469);
nand U1122 (N_1122,N_522,N_345);
nor U1123 (N_1123,N_724,N_408);
xnor U1124 (N_1124,N_466,N_685);
nand U1125 (N_1125,N_570,N_51);
nor U1126 (N_1126,N_240,N_145);
and U1127 (N_1127,N_589,N_269);
nand U1128 (N_1128,N_152,N_650);
nand U1129 (N_1129,N_158,N_252);
nor U1130 (N_1130,N_173,N_113);
or U1131 (N_1131,N_742,N_641);
nor U1132 (N_1132,N_149,N_691);
or U1133 (N_1133,N_256,N_350);
xnor U1134 (N_1134,N_506,N_486);
and U1135 (N_1135,N_5,N_567);
xor U1136 (N_1136,N_186,N_602);
and U1137 (N_1137,N_418,N_300);
xor U1138 (N_1138,N_143,N_679);
or U1139 (N_1139,N_5,N_53);
and U1140 (N_1140,N_41,N_12);
or U1141 (N_1141,N_278,N_338);
or U1142 (N_1142,N_120,N_6);
nand U1143 (N_1143,N_519,N_470);
and U1144 (N_1144,N_320,N_216);
nor U1145 (N_1145,N_425,N_654);
and U1146 (N_1146,N_417,N_567);
and U1147 (N_1147,N_570,N_452);
xor U1148 (N_1148,N_642,N_742);
xnor U1149 (N_1149,N_152,N_436);
nand U1150 (N_1150,N_586,N_342);
nand U1151 (N_1151,N_638,N_395);
or U1152 (N_1152,N_678,N_50);
or U1153 (N_1153,N_657,N_422);
xnor U1154 (N_1154,N_694,N_103);
nand U1155 (N_1155,N_91,N_544);
or U1156 (N_1156,N_377,N_713);
nor U1157 (N_1157,N_439,N_683);
nand U1158 (N_1158,N_420,N_75);
nor U1159 (N_1159,N_652,N_357);
nor U1160 (N_1160,N_471,N_172);
or U1161 (N_1161,N_616,N_137);
or U1162 (N_1162,N_508,N_396);
nor U1163 (N_1163,N_626,N_683);
and U1164 (N_1164,N_131,N_479);
and U1165 (N_1165,N_47,N_120);
xor U1166 (N_1166,N_630,N_425);
xor U1167 (N_1167,N_546,N_296);
xor U1168 (N_1168,N_475,N_297);
nand U1169 (N_1169,N_108,N_731);
nor U1170 (N_1170,N_41,N_463);
nand U1171 (N_1171,N_311,N_529);
nand U1172 (N_1172,N_344,N_640);
nand U1173 (N_1173,N_168,N_382);
or U1174 (N_1174,N_723,N_722);
and U1175 (N_1175,N_209,N_744);
nor U1176 (N_1176,N_749,N_208);
or U1177 (N_1177,N_392,N_658);
or U1178 (N_1178,N_477,N_135);
nor U1179 (N_1179,N_486,N_519);
xnor U1180 (N_1180,N_635,N_611);
nor U1181 (N_1181,N_277,N_430);
or U1182 (N_1182,N_554,N_728);
nor U1183 (N_1183,N_40,N_314);
and U1184 (N_1184,N_208,N_173);
xor U1185 (N_1185,N_225,N_373);
or U1186 (N_1186,N_583,N_447);
xnor U1187 (N_1187,N_646,N_535);
nand U1188 (N_1188,N_562,N_331);
nand U1189 (N_1189,N_209,N_494);
nor U1190 (N_1190,N_298,N_161);
nor U1191 (N_1191,N_305,N_621);
or U1192 (N_1192,N_735,N_635);
xor U1193 (N_1193,N_290,N_531);
and U1194 (N_1194,N_675,N_268);
nor U1195 (N_1195,N_483,N_549);
nor U1196 (N_1196,N_669,N_666);
xnor U1197 (N_1197,N_722,N_75);
xor U1198 (N_1198,N_59,N_561);
and U1199 (N_1199,N_448,N_543);
and U1200 (N_1200,N_340,N_190);
nor U1201 (N_1201,N_312,N_235);
nor U1202 (N_1202,N_226,N_128);
nand U1203 (N_1203,N_541,N_654);
or U1204 (N_1204,N_424,N_26);
and U1205 (N_1205,N_221,N_161);
nor U1206 (N_1206,N_290,N_472);
or U1207 (N_1207,N_596,N_561);
or U1208 (N_1208,N_530,N_542);
or U1209 (N_1209,N_554,N_130);
xnor U1210 (N_1210,N_740,N_685);
and U1211 (N_1211,N_309,N_6);
xor U1212 (N_1212,N_152,N_131);
or U1213 (N_1213,N_154,N_151);
nor U1214 (N_1214,N_114,N_190);
or U1215 (N_1215,N_230,N_220);
nor U1216 (N_1216,N_119,N_129);
xnor U1217 (N_1217,N_424,N_64);
nand U1218 (N_1218,N_534,N_356);
and U1219 (N_1219,N_632,N_266);
and U1220 (N_1220,N_85,N_220);
and U1221 (N_1221,N_603,N_243);
and U1222 (N_1222,N_612,N_402);
nor U1223 (N_1223,N_271,N_377);
xnor U1224 (N_1224,N_218,N_158);
nor U1225 (N_1225,N_122,N_264);
nor U1226 (N_1226,N_715,N_560);
nand U1227 (N_1227,N_62,N_423);
nor U1228 (N_1228,N_216,N_430);
and U1229 (N_1229,N_477,N_282);
nand U1230 (N_1230,N_200,N_316);
or U1231 (N_1231,N_732,N_569);
xor U1232 (N_1232,N_220,N_642);
xnor U1233 (N_1233,N_515,N_563);
or U1234 (N_1234,N_581,N_325);
and U1235 (N_1235,N_496,N_4);
nor U1236 (N_1236,N_424,N_184);
or U1237 (N_1237,N_380,N_319);
and U1238 (N_1238,N_258,N_639);
nand U1239 (N_1239,N_30,N_42);
and U1240 (N_1240,N_60,N_136);
xor U1241 (N_1241,N_235,N_662);
xnor U1242 (N_1242,N_381,N_368);
nand U1243 (N_1243,N_614,N_529);
xnor U1244 (N_1244,N_239,N_554);
nor U1245 (N_1245,N_68,N_36);
or U1246 (N_1246,N_407,N_705);
nor U1247 (N_1247,N_538,N_324);
nand U1248 (N_1248,N_238,N_286);
nor U1249 (N_1249,N_594,N_556);
and U1250 (N_1250,N_360,N_397);
and U1251 (N_1251,N_48,N_702);
nor U1252 (N_1252,N_521,N_136);
nand U1253 (N_1253,N_110,N_183);
nor U1254 (N_1254,N_95,N_269);
or U1255 (N_1255,N_135,N_660);
and U1256 (N_1256,N_686,N_550);
nand U1257 (N_1257,N_131,N_7);
xor U1258 (N_1258,N_11,N_309);
nand U1259 (N_1259,N_357,N_694);
or U1260 (N_1260,N_650,N_72);
nor U1261 (N_1261,N_579,N_19);
xor U1262 (N_1262,N_43,N_521);
nand U1263 (N_1263,N_76,N_484);
nor U1264 (N_1264,N_384,N_688);
nand U1265 (N_1265,N_302,N_377);
nor U1266 (N_1266,N_471,N_101);
nand U1267 (N_1267,N_522,N_485);
and U1268 (N_1268,N_202,N_57);
xor U1269 (N_1269,N_450,N_52);
and U1270 (N_1270,N_33,N_586);
nand U1271 (N_1271,N_496,N_13);
nor U1272 (N_1272,N_743,N_635);
and U1273 (N_1273,N_504,N_461);
or U1274 (N_1274,N_93,N_618);
nand U1275 (N_1275,N_172,N_740);
or U1276 (N_1276,N_710,N_524);
or U1277 (N_1277,N_588,N_241);
nor U1278 (N_1278,N_629,N_747);
nand U1279 (N_1279,N_216,N_267);
xnor U1280 (N_1280,N_243,N_521);
nor U1281 (N_1281,N_467,N_304);
nand U1282 (N_1282,N_580,N_70);
and U1283 (N_1283,N_512,N_63);
and U1284 (N_1284,N_682,N_595);
xnor U1285 (N_1285,N_487,N_539);
or U1286 (N_1286,N_149,N_321);
or U1287 (N_1287,N_349,N_461);
nor U1288 (N_1288,N_106,N_184);
nand U1289 (N_1289,N_25,N_171);
and U1290 (N_1290,N_161,N_283);
xor U1291 (N_1291,N_109,N_598);
and U1292 (N_1292,N_122,N_305);
nand U1293 (N_1293,N_311,N_596);
nand U1294 (N_1294,N_589,N_58);
or U1295 (N_1295,N_700,N_540);
or U1296 (N_1296,N_748,N_329);
and U1297 (N_1297,N_179,N_477);
nand U1298 (N_1298,N_582,N_539);
and U1299 (N_1299,N_58,N_740);
nand U1300 (N_1300,N_285,N_50);
nor U1301 (N_1301,N_725,N_184);
xnor U1302 (N_1302,N_562,N_533);
or U1303 (N_1303,N_497,N_627);
and U1304 (N_1304,N_256,N_282);
nor U1305 (N_1305,N_400,N_22);
or U1306 (N_1306,N_221,N_397);
and U1307 (N_1307,N_105,N_578);
nor U1308 (N_1308,N_482,N_406);
nor U1309 (N_1309,N_528,N_194);
nor U1310 (N_1310,N_619,N_364);
nand U1311 (N_1311,N_441,N_497);
xor U1312 (N_1312,N_360,N_498);
or U1313 (N_1313,N_21,N_531);
or U1314 (N_1314,N_735,N_592);
nor U1315 (N_1315,N_287,N_43);
nand U1316 (N_1316,N_314,N_662);
xor U1317 (N_1317,N_734,N_525);
and U1318 (N_1318,N_210,N_666);
nor U1319 (N_1319,N_716,N_188);
nor U1320 (N_1320,N_726,N_192);
xnor U1321 (N_1321,N_594,N_258);
or U1322 (N_1322,N_119,N_543);
nor U1323 (N_1323,N_407,N_212);
or U1324 (N_1324,N_171,N_357);
and U1325 (N_1325,N_556,N_351);
xor U1326 (N_1326,N_195,N_586);
nand U1327 (N_1327,N_386,N_349);
or U1328 (N_1328,N_575,N_272);
nand U1329 (N_1329,N_435,N_301);
xor U1330 (N_1330,N_676,N_488);
xnor U1331 (N_1331,N_451,N_282);
nand U1332 (N_1332,N_8,N_648);
or U1333 (N_1333,N_570,N_667);
and U1334 (N_1334,N_215,N_609);
xnor U1335 (N_1335,N_189,N_30);
nand U1336 (N_1336,N_393,N_469);
xor U1337 (N_1337,N_174,N_697);
or U1338 (N_1338,N_528,N_239);
nand U1339 (N_1339,N_244,N_92);
xor U1340 (N_1340,N_548,N_661);
nor U1341 (N_1341,N_670,N_169);
nor U1342 (N_1342,N_58,N_301);
nand U1343 (N_1343,N_175,N_651);
nand U1344 (N_1344,N_656,N_335);
or U1345 (N_1345,N_391,N_568);
or U1346 (N_1346,N_406,N_342);
nor U1347 (N_1347,N_241,N_736);
nor U1348 (N_1348,N_747,N_39);
xnor U1349 (N_1349,N_431,N_554);
or U1350 (N_1350,N_240,N_255);
nand U1351 (N_1351,N_99,N_238);
nand U1352 (N_1352,N_558,N_63);
xnor U1353 (N_1353,N_628,N_586);
nor U1354 (N_1354,N_125,N_738);
or U1355 (N_1355,N_494,N_246);
or U1356 (N_1356,N_719,N_109);
xor U1357 (N_1357,N_320,N_205);
nand U1358 (N_1358,N_466,N_621);
nor U1359 (N_1359,N_674,N_734);
or U1360 (N_1360,N_222,N_381);
nand U1361 (N_1361,N_32,N_299);
or U1362 (N_1362,N_635,N_335);
or U1363 (N_1363,N_67,N_371);
xnor U1364 (N_1364,N_373,N_338);
nand U1365 (N_1365,N_439,N_271);
and U1366 (N_1366,N_246,N_661);
and U1367 (N_1367,N_270,N_151);
or U1368 (N_1368,N_37,N_749);
nand U1369 (N_1369,N_470,N_48);
nor U1370 (N_1370,N_623,N_354);
and U1371 (N_1371,N_693,N_582);
xor U1372 (N_1372,N_11,N_197);
and U1373 (N_1373,N_135,N_526);
xnor U1374 (N_1374,N_508,N_556);
xnor U1375 (N_1375,N_2,N_565);
and U1376 (N_1376,N_427,N_145);
nor U1377 (N_1377,N_100,N_209);
and U1378 (N_1378,N_579,N_409);
nand U1379 (N_1379,N_394,N_611);
xor U1380 (N_1380,N_200,N_11);
or U1381 (N_1381,N_31,N_105);
and U1382 (N_1382,N_79,N_194);
xor U1383 (N_1383,N_281,N_465);
and U1384 (N_1384,N_505,N_589);
or U1385 (N_1385,N_132,N_561);
nor U1386 (N_1386,N_182,N_655);
and U1387 (N_1387,N_350,N_370);
xnor U1388 (N_1388,N_281,N_16);
or U1389 (N_1389,N_407,N_27);
nand U1390 (N_1390,N_351,N_292);
nor U1391 (N_1391,N_723,N_29);
nor U1392 (N_1392,N_435,N_414);
xor U1393 (N_1393,N_590,N_484);
or U1394 (N_1394,N_469,N_596);
nor U1395 (N_1395,N_399,N_427);
or U1396 (N_1396,N_435,N_515);
nand U1397 (N_1397,N_716,N_518);
and U1398 (N_1398,N_431,N_369);
or U1399 (N_1399,N_32,N_29);
and U1400 (N_1400,N_214,N_413);
xnor U1401 (N_1401,N_645,N_355);
or U1402 (N_1402,N_235,N_198);
nor U1403 (N_1403,N_186,N_292);
nand U1404 (N_1404,N_321,N_302);
and U1405 (N_1405,N_184,N_672);
and U1406 (N_1406,N_419,N_451);
or U1407 (N_1407,N_276,N_621);
nand U1408 (N_1408,N_744,N_720);
and U1409 (N_1409,N_245,N_386);
xnor U1410 (N_1410,N_159,N_42);
nor U1411 (N_1411,N_554,N_722);
nor U1412 (N_1412,N_658,N_500);
nor U1413 (N_1413,N_294,N_275);
nor U1414 (N_1414,N_338,N_574);
or U1415 (N_1415,N_261,N_551);
xnor U1416 (N_1416,N_271,N_741);
nor U1417 (N_1417,N_169,N_682);
nand U1418 (N_1418,N_322,N_403);
and U1419 (N_1419,N_136,N_233);
xor U1420 (N_1420,N_287,N_155);
nor U1421 (N_1421,N_492,N_440);
xnor U1422 (N_1422,N_699,N_40);
nor U1423 (N_1423,N_313,N_315);
and U1424 (N_1424,N_234,N_449);
xor U1425 (N_1425,N_360,N_741);
or U1426 (N_1426,N_383,N_632);
nor U1427 (N_1427,N_681,N_696);
and U1428 (N_1428,N_569,N_566);
nand U1429 (N_1429,N_648,N_316);
or U1430 (N_1430,N_705,N_293);
and U1431 (N_1431,N_698,N_351);
or U1432 (N_1432,N_455,N_207);
xor U1433 (N_1433,N_449,N_392);
and U1434 (N_1434,N_577,N_515);
xnor U1435 (N_1435,N_554,N_448);
nand U1436 (N_1436,N_660,N_30);
nand U1437 (N_1437,N_117,N_557);
or U1438 (N_1438,N_442,N_73);
and U1439 (N_1439,N_65,N_54);
nor U1440 (N_1440,N_292,N_6);
nand U1441 (N_1441,N_38,N_159);
nor U1442 (N_1442,N_749,N_11);
or U1443 (N_1443,N_436,N_68);
nand U1444 (N_1444,N_519,N_165);
or U1445 (N_1445,N_99,N_269);
and U1446 (N_1446,N_532,N_226);
xnor U1447 (N_1447,N_352,N_285);
and U1448 (N_1448,N_492,N_362);
nor U1449 (N_1449,N_409,N_637);
nor U1450 (N_1450,N_56,N_128);
or U1451 (N_1451,N_597,N_593);
and U1452 (N_1452,N_485,N_374);
nand U1453 (N_1453,N_314,N_249);
nand U1454 (N_1454,N_361,N_263);
nand U1455 (N_1455,N_139,N_422);
nor U1456 (N_1456,N_107,N_51);
and U1457 (N_1457,N_391,N_321);
or U1458 (N_1458,N_261,N_528);
nor U1459 (N_1459,N_207,N_248);
nor U1460 (N_1460,N_478,N_346);
xor U1461 (N_1461,N_587,N_589);
nand U1462 (N_1462,N_510,N_255);
and U1463 (N_1463,N_92,N_377);
or U1464 (N_1464,N_291,N_741);
nor U1465 (N_1465,N_128,N_234);
nor U1466 (N_1466,N_668,N_712);
xnor U1467 (N_1467,N_474,N_693);
nor U1468 (N_1468,N_339,N_174);
or U1469 (N_1469,N_617,N_628);
nand U1470 (N_1470,N_205,N_277);
and U1471 (N_1471,N_67,N_604);
nand U1472 (N_1472,N_561,N_543);
nor U1473 (N_1473,N_343,N_121);
or U1474 (N_1474,N_158,N_77);
and U1475 (N_1475,N_247,N_133);
or U1476 (N_1476,N_599,N_332);
xnor U1477 (N_1477,N_693,N_147);
or U1478 (N_1478,N_21,N_267);
xnor U1479 (N_1479,N_267,N_695);
and U1480 (N_1480,N_636,N_227);
nand U1481 (N_1481,N_684,N_702);
or U1482 (N_1482,N_244,N_485);
xor U1483 (N_1483,N_569,N_583);
or U1484 (N_1484,N_88,N_349);
xor U1485 (N_1485,N_396,N_102);
or U1486 (N_1486,N_670,N_711);
xor U1487 (N_1487,N_384,N_122);
or U1488 (N_1488,N_231,N_356);
xor U1489 (N_1489,N_227,N_1);
and U1490 (N_1490,N_478,N_412);
nor U1491 (N_1491,N_334,N_1);
nand U1492 (N_1492,N_683,N_438);
and U1493 (N_1493,N_208,N_627);
nand U1494 (N_1494,N_44,N_585);
or U1495 (N_1495,N_8,N_639);
nand U1496 (N_1496,N_700,N_154);
nor U1497 (N_1497,N_23,N_244);
xnor U1498 (N_1498,N_87,N_180);
nor U1499 (N_1499,N_382,N_543);
or U1500 (N_1500,N_1295,N_1352);
xor U1501 (N_1501,N_1254,N_1173);
xor U1502 (N_1502,N_1279,N_1430);
xor U1503 (N_1503,N_1443,N_1498);
nand U1504 (N_1504,N_1466,N_1458);
nand U1505 (N_1505,N_874,N_1005);
xnor U1506 (N_1506,N_984,N_829);
and U1507 (N_1507,N_764,N_893);
nand U1508 (N_1508,N_1333,N_1341);
or U1509 (N_1509,N_912,N_1322);
nor U1510 (N_1510,N_1261,N_919);
nor U1511 (N_1511,N_1469,N_1417);
nand U1512 (N_1512,N_1052,N_1349);
xnor U1513 (N_1513,N_866,N_973);
or U1514 (N_1514,N_966,N_1043);
and U1515 (N_1515,N_1362,N_1377);
and U1516 (N_1516,N_1138,N_1372);
nor U1517 (N_1517,N_989,N_1178);
xnor U1518 (N_1518,N_1350,N_1402);
nor U1519 (N_1519,N_1007,N_992);
xnor U1520 (N_1520,N_1422,N_1131);
and U1521 (N_1521,N_1166,N_882);
nor U1522 (N_1522,N_977,N_924);
or U1523 (N_1523,N_1130,N_1197);
nand U1524 (N_1524,N_800,N_1236);
or U1525 (N_1525,N_892,N_765);
nand U1526 (N_1526,N_902,N_768);
nand U1527 (N_1527,N_858,N_1171);
xnor U1528 (N_1528,N_1081,N_1202);
nand U1529 (N_1529,N_1114,N_1061);
nand U1530 (N_1530,N_1355,N_870);
nor U1531 (N_1531,N_1191,N_1012);
or U1532 (N_1532,N_759,N_873);
nor U1533 (N_1533,N_916,N_1159);
or U1534 (N_1534,N_1331,N_986);
or U1535 (N_1535,N_795,N_1426);
and U1536 (N_1536,N_1281,N_1106);
or U1537 (N_1537,N_1309,N_1205);
and U1538 (N_1538,N_1297,N_1237);
xor U1539 (N_1539,N_1014,N_1464);
or U1540 (N_1540,N_1448,N_917);
xor U1541 (N_1541,N_1453,N_1489);
nor U1542 (N_1542,N_944,N_1212);
nor U1543 (N_1543,N_1395,N_754);
nor U1544 (N_1544,N_1278,N_1463);
and U1545 (N_1545,N_1163,N_1328);
or U1546 (N_1546,N_1493,N_1234);
nand U1547 (N_1547,N_1357,N_1168);
nand U1548 (N_1548,N_1023,N_1062);
and U1549 (N_1549,N_1269,N_1070);
and U1550 (N_1550,N_950,N_817);
nand U1551 (N_1551,N_1450,N_1240);
and U1552 (N_1552,N_786,N_1113);
or U1553 (N_1553,N_1442,N_861);
nor U1554 (N_1554,N_1414,N_1326);
xnor U1555 (N_1555,N_910,N_1369);
or U1556 (N_1556,N_833,N_1193);
or U1557 (N_1557,N_813,N_1293);
nor U1558 (N_1558,N_782,N_921);
nand U1559 (N_1559,N_775,N_1003);
xor U1560 (N_1560,N_1050,N_1275);
nor U1561 (N_1561,N_1084,N_1010);
or U1562 (N_1562,N_1207,N_1145);
nor U1563 (N_1563,N_1066,N_1385);
or U1564 (N_1564,N_1413,N_1340);
nor U1565 (N_1565,N_979,N_798);
nand U1566 (N_1566,N_785,N_1313);
xnor U1567 (N_1567,N_1096,N_884);
and U1568 (N_1568,N_1072,N_1040);
and U1569 (N_1569,N_1201,N_1231);
and U1570 (N_1570,N_1058,N_1404);
nand U1571 (N_1571,N_1018,N_1223);
and U1572 (N_1572,N_1107,N_1472);
nand U1573 (N_1573,N_1488,N_951);
and U1574 (N_1574,N_1170,N_1143);
xor U1575 (N_1575,N_1270,N_1051);
nand U1576 (N_1576,N_932,N_1181);
or U1577 (N_1577,N_1255,N_1339);
nand U1578 (N_1578,N_896,N_1116);
nor U1579 (N_1579,N_1336,N_1308);
nand U1580 (N_1580,N_796,N_1054);
nor U1581 (N_1581,N_1247,N_783);
nor U1582 (N_1582,N_1048,N_1348);
and U1583 (N_1583,N_815,N_1219);
and U1584 (N_1584,N_925,N_1423);
and U1585 (N_1585,N_1174,N_975);
nor U1586 (N_1586,N_946,N_955);
nand U1587 (N_1587,N_1465,N_755);
or U1588 (N_1588,N_1155,N_805);
and U1589 (N_1589,N_1002,N_857);
xor U1590 (N_1590,N_788,N_1444);
or U1591 (N_1591,N_846,N_1361);
nor U1592 (N_1592,N_1125,N_757);
and U1593 (N_1593,N_1157,N_1120);
and U1594 (N_1594,N_1259,N_825);
nand U1595 (N_1595,N_1388,N_1343);
nand U1596 (N_1596,N_900,N_1449);
or U1597 (N_1597,N_1306,N_1277);
and U1598 (N_1598,N_806,N_790);
xnor U1599 (N_1599,N_1300,N_934);
nor U1600 (N_1600,N_1367,N_1437);
nand U1601 (N_1601,N_766,N_1042);
nor U1602 (N_1602,N_940,N_1264);
and U1603 (N_1603,N_1312,N_1016);
nor U1604 (N_1604,N_1345,N_1188);
nor U1605 (N_1605,N_830,N_1088);
nor U1606 (N_1606,N_879,N_1475);
or U1607 (N_1607,N_1126,N_1325);
xor U1608 (N_1608,N_1418,N_1029);
xor U1609 (N_1609,N_1440,N_1396);
and U1610 (N_1610,N_799,N_1015);
nor U1611 (N_1611,N_1097,N_1141);
and U1612 (N_1612,N_845,N_1401);
and U1613 (N_1613,N_850,N_1479);
xnor U1614 (N_1614,N_991,N_1447);
or U1615 (N_1615,N_1482,N_956);
nor U1616 (N_1616,N_1135,N_1260);
nor U1617 (N_1617,N_888,N_1045);
nand U1618 (N_1618,N_988,N_1287);
nand U1619 (N_1619,N_1221,N_1228);
xnor U1620 (N_1620,N_1316,N_1215);
or U1621 (N_1621,N_939,N_1085);
xor U1622 (N_1622,N_1271,N_1059);
xnor U1623 (N_1623,N_1071,N_831);
nor U1624 (N_1624,N_1195,N_981);
and U1625 (N_1625,N_1146,N_952);
or U1626 (N_1626,N_1021,N_953);
nand U1627 (N_1627,N_852,N_1124);
nor U1628 (N_1628,N_1108,N_836);
nor U1629 (N_1629,N_1365,N_1383);
or U1630 (N_1630,N_1315,N_980);
nand U1631 (N_1631,N_774,N_1429);
or U1632 (N_1632,N_942,N_1499);
or U1633 (N_1633,N_818,N_1144);
nand U1634 (N_1634,N_1397,N_1068);
xor U1635 (N_1635,N_793,N_1233);
or U1636 (N_1636,N_1153,N_1462);
nand U1637 (N_1637,N_1387,N_862);
nor U1638 (N_1638,N_1064,N_1087);
nor U1639 (N_1639,N_928,N_1338);
or U1640 (N_1640,N_1224,N_1244);
or U1641 (N_1641,N_1351,N_1276);
xnor U1642 (N_1642,N_1384,N_1209);
and U1643 (N_1643,N_773,N_983);
or U1644 (N_1644,N_963,N_1327);
or U1645 (N_1645,N_1284,N_1399);
xor U1646 (N_1646,N_840,N_1137);
nand U1647 (N_1647,N_1119,N_1394);
and U1648 (N_1648,N_753,N_1147);
nor U1649 (N_1649,N_1089,N_1329);
and U1650 (N_1650,N_876,N_1492);
nor U1651 (N_1651,N_811,N_1185);
xnor U1652 (N_1652,N_769,N_1265);
and U1653 (N_1653,N_1075,N_1100);
nand U1654 (N_1654,N_1238,N_1187);
or U1655 (N_1655,N_1156,N_1290);
xor U1656 (N_1656,N_1006,N_1026);
xnor U1657 (N_1657,N_1216,N_1353);
xor U1658 (N_1658,N_751,N_1366);
or U1659 (N_1659,N_1342,N_1410);
xnor U1660 (N_1660,N_1213,N_804);
and U1661 (N_1661,N_756,N_1301);
nand U1662 (N_1662,N_1235,N_1127);
nand U1663 (N_1663,N_1063,N_1432);
nand U1664 (N_1664,N_926,N_1198);
nand U1665 (N_1665,N_1232,N_1057);
nand U1666 (N_1666,N_909,N_851);
nand U1667 (N_1667,N_985,N_1407);
and U1668 (N_1668,N_1317,N_864);
and U1669 (N_1669,N_1041,N_885);
or U1670 (N_1670,N_1183,N_1167);
nor U1671 (N_1671,N_1477,N_1030);
nor U1672 (N_1672,N_936,N_971);
or U1673 (N_1673,N_899,N_863);
or U1674 (N_1674,N_854,N_1476);
and U1675 (N_1675,N_1379,N_1082);
nor U1676 (N_1676,N_837,N_1031);
and U1677 (N_1677,N_841,N_1434);
xnor U1678 (N_1678,N_1090,N_1467);
nor U1679 (N_1679,N_1140,N_1251);
and U1680 (N_1680,N_1027,N_1298);
nand U1681 (N_1681,N_843,N_1245);
or U1682 (N_1682,N_1334,N_1204);
xnor U1683 (N_1683,N_1321,N_886);
xor U1684 (N_1684,N_1182,N_752);
nand U1685 (N_1685,N_931,N_1494);
nor U1686 (N_1686,N_930,N_890);
nor U1687 (N_1687,N_1009,N_1373);
or U1688 (N_1688,N_1268,N_908);
nor U1689 (N_1689,N_1076,N_1389);
xnor U1690 (N_1690,N_1038,N_878);
xor U1691 (N_1691,N_1225,N_1056);
and U1692 (N_1692,N_1077,N_1128);
xnor U1693 (N_1693,N_1360,N_976);
nand U1694 (N_1694,N_1065,N_1335);
xor U1695 (N_1695,N_1046,N_933);
nor U1696 (N_1696,N_860,N_1337);
or U1697 (N_1697,N_1374,N_938);
and U1698 (N_1698,N_1400,N_810);
and U1699 (N_1699,N_762,N_1391);
nor U1700 (N_1700,N_1382,N_907);
nor U1701 (N_1701,N_1020,N_1456);
or U1702 (N_1702,N_1304,N_770);
nor U1703 (N_1703,N_871,N_835);
nor U1704 (N_1704,N_1129,N_1176);
xnor U1705 (N_1705,N_894,N_1378);
nand U1706 (N_1706,N_839,N_1017);
xnor U1707 (N_1707,N_1473,N_1266);
or U1708 (N_1708,N_889,N_990);
and U1709 (N_1709,N_993,N_945);
xor U1710 (N_1710,N_1218,N_1037);
or U1711 (N_1711,N_969,N_1206);
or U1712 (N_1712,N_1148,N_972);
nor U1713 (N_1713,N_1289,N_1452);
and U1714 (N_1714,N_809,N_923);
nor U1715 (N_1715,N_1164,N_987);
nand U1716 (N_1716,N_1019,N_1283);
nor U1717 (N_1717,N_1445,N_1495);
nor U1718 (N_1718,N_997,N_1091);
nor U1719 (N_1719,N_847,N_1274);
or U1720 (N_1720,N_819,N_1291);
and U1721 (N_1721,N_1408,N_1222);
nand U1722 (N_1722,N_1484,N_875);
or U1723 (N_1723,N_1288,N_750);
and U1724 (N_1724,N_1250,N_877);
or U1725 (N_1725,N_1226,N_1421);
nand U1726 (N_1726,N_1122,N_1123);
or U1727 (N_1727,N_767,N_1241);
nor U1728 (N_1728,N_802,N_1139);
xnor U1729 (N_1729,N_1253,N_842);
xnor U1730 (N_1730,N_1214,N_1083);
or U1731 (N_1731,N_1272,N_1133);
and U1732 (N_1732,N_1092,N_1381);
or U1733 (N_1733,N_904,N_1405);
nand U1734 (N_1734,N_1302,N_1285);
or U1735 (N_1735,N_1314,N_1386);
nand U1736 (N_1736,N_776,N_915);
xnor U1737 (N_1737,N_935,N_898);
nand U1738 (N_1738,N_1118,N_1152);
nand U1739 (N_1739,N_1239,N_1318);
or U1740 (N_1740,N_859,N_1175);
or U1741 (N_1741,N_1332,N_1249);
nand U1742 (N_1742,N_1194,N_1110);
or U1743 (N_1743,N_1371,N_832);
nor U1744 (N_1744,N_853,N_1032);
or U1745 (N_1745,N_978,N_849);
nand U1746 (N_1746,N_794,N_922);
and U1747 (N_1747,N_758,N_1210);
and U1748 (N_1748,N_1109,N_895);
xnor U1749 (N_1749,N_1177,N_1470);
nand U1750 (N_1750,N_1104,N_1098);
and U1751 (N_1751,N_855,N_838);
and U1752 (N_1752,N_1460,N_868);
nor U1753 (N_1753,N_982,N_1069);
xnor U1754 (N_1754,N_1478,N_1474);
nor U1755 (N_1755,N_848,N_1438);
or U1756 (N_1756,N_1347,N_760);
xor U1757 (N_1757,N_1103,N_1172);
xor U1758 (N_1758,N_1370,N_1451);
or U1759 (N_1759,N_1263,N_1368);
xnor U1760 (N_1760,N_1267,N_937);
and U1761 (N_1761,N_998,N_964);
and U1762 (N_1762,N_1034,N_958);
or U1763 (N_1763,N_1427,N_1162);
nor U1764 (N_1764,N_1256,N_974);
xor U1765 (N_1765,N_856,N_801);
xnor U1766 (N_1766,N_834,N_1243);
and U1767 (N_1767,N_1011,N_1189);
xor U1768 (N_1768,N_996,N_1364);
and U1769 (N_1769,N_1296,N_1203);
or U1770 (N_1770,N_781,N_1420);
nand U1771 (N_1771,N_1022,N_1099);
nor U1772 (N_1772,N_1192,N_959);
nand U1773 (N_1773,N_1008,N_995);
xor U1774 (N_1774,N_1419,N_1471);
xnor U1775 (N_1775,N_1280,N_1044);
xor U1776 (N_1776,N_1190,N_1000);
xnor U1777 (N_1777,N_901,N_999);
nand U1778 (N_1778,N_961,N_1154);
nand U1779 (N_1779,N_1258,N_891);
xor U1780 (N_1780,N_1487,N_867);
xnor U1781 (N_1781,N_1497,N_887);
and U1782 (N_1782,N_1480,N_1398);
nand U1783 (N_1783,N_1424,N_784);
nor U1784 (N_1784,N_812,N_1409);
xnor U1785 (N_1785,N_1481,N_883);
xnor U1786 (N_1786,N_1282,N_1102);
nor U1787 (N_1787,N_881,N_1319);
nor U1788 (N_1788,N_1320,N_965);
xor U1789 (N_1789,N_869,N_1229);
xor U1790 (N_1790,N_1035,N_1033);
nor U1791 (N_1791,N_947,N_913);
or U1792 (N_1792,N_761,N_1165);
nor U1793 (N_1793,N_816,N_897);
nor U1794 (N_1794,N_1230,N_1211);
nand U1795 (N_1795,N_1380,N_778);
or U1796 (N_1796,N_1094,N_1180);
or U1797 (N_1797,N_1093,N_1055);
nand U1798 (N_1798,N_1112,N_1199);
nand U1799 (N_1799,N_1428,N_1151);
xnor U1800 (N_1800,N_1134,N_1436);
nor U1801 (N_1801,N_824,N_1496);
nor U1802 (N_1802,N_1217,N_918);
xnor U1803 (N_1803,N_1025,N_780);
nand U1804 (N_1804,N_777,N_1346);
nand U1805 (N_1805,N_1344,N_791);
and U1806 (N_1806,N_880,N_1299);
and U1807 (N_1807,N_771,N_905);
xnor U1808 (N_1808,N_1095,N_1273);
and U1809 (N_1809,N_914,N_1242);
xor U1810 (N_1810,N_763,N_1179);
nand U1811 (N_1811,N_1047,N_792);
or U1812 (N_1812,N_906,N_1220);
and U1813 (N_1813,N_1406,N_1028);
xnor U1814 (N_1814,N_957,N_772);
nor U1815 (N_1815,N_1363,N_1080);
nor U1816 (N_1816,N_1142,N_787);
xnor U1817 (N_1817,N_1311,N_1485);
nand U1818 (N_1818,N_1491,N_941);
nor U1819 (N_1819,N_844,N_1415);
nor U1820 (N_1820,N_814,N_1036);
and U1821 (N_1821,N_1411,N_1049);
nor U1822 (N_1822,N_1067,N_1186);
nand U1823 (N_1823,N_1305,N_1292);
and U1824 (N_1824,N_1208,N_1433);
nand U1825 (N_1825,N_960,N_1246);
xnor U1826 (N_1826,N_967,N_1393);
xnor U1827 (N_1827,N_1486,N_1468);
nand U1828 (N_1828,N_822,N_1390);
nand U1829 (N_1829,N_1086,N_823);
and U1830 (N_1830,N_1158,N_1004);
nand U1831 (N_1831,N_1121,N_1455);
and U1832 (N_1832,N_1074,N_1150);
and U1833 (N_1833,N_911,N_1105);
nand U1834 (N_1834,N_1053,N_865);
and U1835 (N_1835,N_1457,N_1392);
xnor U1836 (N_1836,N_1149,N_1330);
nand U1837 (N_1837,N_827,N_1294);
xnor U1838 (N_1838,N_1252,N_1376);
or U1839 (N_1839,N_968,N_1184);
and U1840 (N_1840,N_1161,N_1359);
nor U1841 (N_1841,N_1459,N_1111);
nor U1842 (N_1842,N_1310,N_821);
nor U1843 (N_1843,N_1425,N_1431);
and U1844 (N_1844,N_1039,N_1132);
nand U1845 (N_1845,N_1375,N_807);
nor U1846 (N_1846,N_970,N_1060);
xor U1847 (N_1847,N_1078,N_1248);
or U1848 (N_1848,N_789,N_1435);
nand U1849 (N_1849,N_779,N_1262);
and U1850 (N_1850,N_1354,N_826);
nor U1851 (N_1851,N_1160,N_1461);
nor U1852 (N_1852,N_1257,N_1079);
or U1853 (N_1853,N_1169,N_1101);
and U1854 (N_1854,N_1412,N_1013);
nand U1855 (N_1855,N_1136,N_1073);
or U1856 (N_1856,N_1200,N_929);
and U1857 (N_1857,N_1441,N_1358);
and U1858 (N_1858,N_1115,N_1483);
nor U1859 (N_1859,N_962,N_920);
nor U1860 (N_1860,N_1286,N_927);
and U1861 (N_1861,N_1403,N_1454);
xor U1862 (N_1862,N_949,N_1490);
and U1863 (N_1863,N_1356,N_1117);
nor U1864 (N_1864,N_820,N_954);
xnor U1865 (N_1865,N_948,N_797);
nand U1866 (N_1866,N_872,N_943);
xor U1867 (N_1867,N_1227,N_1439);
xnor U1868 (N_1868,N_994,N_1307);
nor U1869 (N_1869,N_803,N_1416);
xnor U1870 (N_1870,N_1446,N_1303);
xor U1871 (N_1871,N_808,N_1196);
xnor U1872 (N_1872,N_828,N_1324);
and U1873 (N_1873,N_1024,N_1323);
nor U1874 (N_1874,N_903,N_1001);
nor U1875 (N_1875,N_816,N_1346);
or U1876 (N_1876,N_1158,N_1224);
and U1877 (N_1877,N_806,N_1463);
or U1878 (N_1878,N_790,N_1186);
nor U1879 (N_1879,N_1075,N_1058);
nand U1880 (N_1880,N_1002,N_1080);
xnor U1881 (N_1881,N_1177,N_1407);
and U1882 (N_1882,N_1226,N_1139);
or U1883 (N_1883,N_1202,N_1258);
and U1884 (N_1884,N_1448,N_809);
and U1885 (N_1885,N_821,N_873);
xnor U1886 (N_1886,N_1147,N_974);
nor U1887 (N_1887,N_1059,N_1008);
nor U1888 (N_1888,N_1455,N_864);
and U1889 (N_1889,N_1125,N_851);
or U1890 (N_1890,N_1280,N_818);
xor U1891 (N_1891,N_1134,N_1085);
and U1892 (N_1892,N_1029,N_1340);
nor U1893 (N_1893,N_881,N_977);
nor U1894 (N_1894,N_1076,N_1239);
xor U1895 (N_1895,N_851,N_874);
nand U1896 (N_1896,N_1036,N_1239);
or U1897 (N_1897,N_1287,N_1227);
or U1898 (N_1898,N_1270,N_997);
and U1899 (N_1899,N_1414,N_1457);
nand U1900 (N_1900,N_1433,N_1218);
nor U1901 (N_1901,N_1249,N_1446);
or U1902 (N_1902,N_948,N_1345);
xnor U1903 (N_1903,N_1453,N_1333);
xnor U1904 (N_1904,N_1143,N_767);
nand U1905 (N_1905,N_760,N_1436);
nand U1906 (N_1906,N_1463,N_1253);
and U1907 (N_1907,N_960,N_1239);
or U1908 (N_1908,N_1181,N_1490);
nor U1909 (N_1909,N_1201,N_1203);
nor U1910 (N_1910,N_1392,N_780);
nor U1911 (N_1911,N_943,N_1472);
and U1912 (N_1912,N_771,N_789);
nand U1913 (N_1913,N_1049,N_955);
nand U1914 (N_1914,N_908,N_934);
nor U1915 (N_1915,N_1246,N_906);
nor U1916 (N_1916,N_959,N_1006);
and U1917 (N_1917,N_1116,N_1493);
xor U1918 (N_1918,N_909,N_1379);
or U1919 (N_1919,N_1393,N_758);
and U1920 (N_1920,N_851,N_1017);
or U1921 (N_1921,N_1458,N_866);
or U1922 (N_1922,N_1128,N_894);
xor U1923 (N_1923,N_1089,N_1269);
and U1924 (N_1924,N_1440,N_833);
nand U1925 (N_1925,N_980,N_1201);
nor U1926 (N_1926,N_876,N_1375);
and U1927 (N_1927,N_1057,N_1114);
or U1928 (N_1928,N_1489,N_1091);
or U1929 (N_1929,N_1476,N_975);
nand U1930 (N_1930,N_1443,N_1421);
or U1931 (N_1931,N_1072,N_1381);
xor U1932 (N_1932,N_1317,N_1168);
nor U1933 (N_1933,N_799,N_1163);
xor U1934 (N_1934,N_1314,N_782);
nand U1935 (N_1935,N_1410,N_1222);
or U1936 (N_1936,N_997,N_1304);
nand U1937 (N_1937,N_1291,N_1338);
nor U1938 (N_1938,N_1198,N_1339);
or U1939 (N_1939,N_1060,N_906);
or U1940 (N_1940,N_1009,N_1204);
or U1941 (N_1941,N_1438,N_934);
nand U1942 (N_1942,N_792,N_938);
or U1943 (N_1943,N_1094,N_814);
or U1944 (N_1944,N_1331,N_1078);
nor U1945 (N_1945,N_1039,N_1197);
and U1946 (N_1946,N_1471,N_1116);
nand U1947 (N_1947,N_1450,N_1205);
xnor U1948 (N_1948,N_1056,N_1312);
nor U1949 (N_1949,N_1000,N_1327);
nand U1950 (N_1950,N_1279,N_1465);
or U1951 (N_1951,N_1102,N_1225);
nor U1952 (N_1952,N_1434,N_752);
and U1953 (N_1953,N_949,N_1446);
nand U1954 (N_1954,N_1326,N_1457);
nor U1955 (N_1955,N_1144,N_1424);
nand U1956 (N_1956,N_1277,N_1085);
or U1957 (N_1957,N_884,N_1445);
and U1958 (N_1958,N_1185,N_1047);
xnor U1959 (N_1959,N_872,N_993);
or U1960 (N_1960,N_952,N_1185);
nand U1961 (N_1961,N_1305,N_1266);
nand U1962 (N_1962,N_1253,N_1478);
nand U1963 (N_1963,N_1021,N_942);
nand U1964 (N_1964,N_803,N_1435);
or U1965 (N_1965,N_842,N_840);
xor U1966 (N_1966,N_922,N_1230);
xnor U1967 (N_1967,N_847,N_1099);
xor U1968 (N_1968,N_1391,N_1339);
xnor U1969 (N_1969,N_1276,N_1460);
and U1970 (N_1970,N_779,N_969);
or U1971 (N_1971,N_1070,N_1318);
nand U1972 (N_1972,N_1088,N_1132);
nand U1973 (N_1973,N_1343,N_1199);
or U1974 (N_1974,N_830,N_1403);
nor U1975 (N_1975,N_1477,N_1416);
xor U1976 (N_1976,N_1383,N_1495);
nand U1977 (N_1977,N_894,N_1482);
nor U1978 (N_1978,N_767,N_972);
xnor U1979 (N_1979,N_987,N_1169);
nor U1980 (N_1980,N_1207,N_765);
or U1981 (N_1981,N_1032,N_1140);
and U1982 (N_1982,N_1084,N_1138);
nor U1983 (N_1983,N_1009,N_1278);
xor U1984 (N_1984,N_1074,N_907);
nor U1985 (N_1985,N_954,N_1336);
xor U1986 (N_1986,N_1093,N_775);
or U1987 (N_1987,N_1203,N_1273);
or U1988 (N_1988,N_966,N_902);
xnor U1989 (N_1989,N_910,N_796);
and U1990 (N_1990,N_1438,N_840);
or U1991 (N_1991,N_1012,N_1248);
nor U1992 (N_1992,N_1173,N_1045);
or U1993 (N_1993,N_1145,N_767);
nand U1994 (N_1994,N_1113,N_1197);
or U1995 (N_1995,N_944,N_1240);
or U1996 (N_1996,N_765,N_821);
xnor U1997 (N_1997,N_1326,N_817);
nand U1998 (N_1998,N_915,N_1495);
or U1999 (N_1999,N_965,N_886);
nand U2000 (N_2000,N_1482,N_1001);
and U2001 (N_2001,N_1137,N_786);
and U2002 (N_2002,N_947,N_760);
nand U2003 (N_2003,N_911,N_778);
or U2004 (N_2004,N_1012,N_1068);
nand U2005 (N_2005,N_1129,N_779);
nand U2006 (N_2006,N_1140,N_1127);
xnor U2007 (N_2007,N_1107,N_1183);
nor U2008 (N_2008,N_1153,N_1418);
or U2009 (N_2009,N_1379,N_1003);
or U2010 (N_2010,N_1321,N_1296);
or U2011 (N_2011,N_817,N_1488);
nor U2012 (N_2012,N_1346,N_851);
or U2013 (N_2013,N_1188,N_1087);
nor U2014 (N_2014,N_1310,N_856);
nand U2015 (N_2015,N_950,N_1083);
xor U2016 (N_2016,N_886,N_1293);
or U2017 (N_2017,N_799,N_1124);
and U2018 (N_2018,N_1061,N_962);
or U2019 (N_2019,N_919,N_867);
or U2020 (N_2020,N_1152,N_1043);
nand U2021 (N_2021,N_949,N_1443);
and U2022 (N_2022,N_1171,N_1075);
and U2023 (N_2023,N_1325,N_978);
nor U2024 (N_2024,N_859,N_977);
or U2025 (N_2025,N_1325,N_848);
or U2026 (N_2026,N_1060,N_1196);
xnor U2027 (N_2027,N_808,N_1165);
nand U2028 (N_2028,N_1320,N_1420);
nor U2029 (N_2029,N_1285,N_907);
or U2030 (N_2030,N_1049,N_1127);
xnor U2031 (N_2031,N_1361,N_1023);
xor U2032 (N_2032,N_828,N_956);
nor U2033 (N_2033,N_1486,N_916);
nor U2034 (N_2034,N_1094,N_929);
nand U2035 (N_2035,N_985,N_1270);
and U2036 (N_2036,N_1228,N_873);
or U2037 (N_2037,N_1072,N_1044);
nor U2038 (N_2038,N_1465,N_1090);
nor U2039 (N_2039,N_1209,N_868);
or U2040 (N_2040,N_753,N_1386);
xnor U2041 (N_2041,N_757,N_1207);
nor U2042 (N_2042,N_1187,N_1473);
xor U2043 (N_2043,N_920,N_1115);
or U2044 (N_2044,N_1091,N_1141);
xor U2045 (N_2045,N_1189,N_829);
nand U2046 (N_2046,N_988,N_1005);
and U2047 (N_2047,N_968,N_993);
xor U2048 (N_2048,N_1117,N_829);
and U2049 (N_2049,N_1079,N_1242);
and U2050 (N_2050,N_1259,N_1234);
xnor U2051 (N_2051,N_1047,N_1020);
and U2052 (N_2052,N_1174,N_1438);
nor U2053 (N_2053,N_1365,N_769);
xnor U2054 (N_2054,N_1437,N_899);
xnor U2055 (N_2055,N_1221,N_1371);
xnor U2056 (N_2056,N_1060,N_802);
nor U2057 (N_2057,N_1219,N_899);
nand U2058 (N_2058,N_1071,N_1301);
nor U2059 (N_2059,N_1126,N_1026);
or U2060 (N_2060,N_1203,N_800);
nor U2061 (N_2061,N_1282,N_1347);
nand U2062 (N_2062,N_1143,N_1008);
xor U2063 (N_2063,N_898,N_1034);
or U2064 (N_2064,N_1011,N_881);
xor U2065 (N_2065,N_1126,N_1106);
xor U2066 (N_2066,N_869,N_919);
nand U2067 (N_2067,N_938,N_1144);
xnor U2068 (N_2068,N_982,N_1160);
nor U2069 (N_2069,N_790,N_1228);
or U2070 (N_2070,N_1124,N_1075);
or U2071 (N_2071,N_878,N_1491);
nand U2072 (N_2072,N_968,N_1343);
and U2073 (N_2073,N_1038,N_1257);
or U2074 (N_2074,N_1263,N_805);
nand U2075 (N_2075,N_907,N_876);
and U2076 (N_2076,N_1212,N_1223);
nor U2077 (N_2077,N_1138,N_1406);
nor U2078 (N_2078,N_1351,N_1148);
or U2079 (N_2079,N_1472,N_1235);
and U2080 (N_2080,N_1494,N_1133);
xor U2081 (N_2081,N_1235,N_1372);
and U2082 (N_2082,N_823,N_975);
or U2083 (N_2083,N_767,N_901);
or U2084 (N_2084,N_1222,N_760);
nor U2085 (N_2085,N_1396,N_974);
nand U2086 (N_2086,N_1200,N_955);
nor U2087 (N_2087,N_1105,N_1262);
or U2088 (N_2088,N_774,N_1219);
nor U2089 (N_2089,N_846,N_802);
and U2090 (N_2090,N_1388,N_789);
or U2091 (N_2091,N_1388,N_1042);
or U2092 (N_2092,N_1092,N_1072);
xnor U2093 (N_2093,N_866,N_1278);
and U2094 (N_2094,N_1240,N_1048);
xor U2095 (N_2095,N_975,N_853);
and U2096 (N_2096,N_873,N_1466);
nand U2097 (N_2097,N_1123,N_891);
and U2098 (N_2098,N_1009,N_844);
and U2099 (N_2099,N_1082,N_1255);
and U2100 (N_2100,N_1471,N_1239);
xor U2101 (N_2101,N_974,N_867);
and U2102 (N_2102,N_982,N_765);
or U2103 (N_2103,N_770,N_1028);
nor U2104 (N_2104,N_1045,N_828);
xor U2105 (N_2105,N_1191,N_1223);
xnor U2106 (N_2106,N_1458,N_1311);
and U2107 (N_2107,N_1193,N_1276);
or U2108 (N_2108,N_1484,N_1242);
nor U2109 (N_2109,N_1046,N_1049);
xor U2110 (N_2110,N_1485,N_1325);
and U2111 (N_2111,N_850,N_1387);
nor U2112 (N_2112,N_1013,N_1497);
xnor U2113 (N_2113,N_761,N_929);
xnor U2114 (N_2114,N_753,N_820);
nand U2115 (N_2115,N_1253,N_1496);
or U2116 (N_2116,N_1478,N_1486);
or U2117 (N_2117,N_902,N_939);
and U2118 (N_2118,N_1377,N_1056);
and U2119 (N_2119,N_1285,N_859);
and U2120 (N_2120,N_765,N_938);
xor U2121 (N_2121,N_1017,N_824);
xnor U2122 (N_2122,N_1036,N_893);
or U2123 (N_2123,N_1033,N_795);
nand U2124 (N_2124,N_1215,N_977);
nand U2125 (N_2125,N_1032,N_1147);
nand U2126 (N_2126,N_1434,N_835);
and U2127 (N_2127,N_810,N_999);
nor U2128 (N_2128,N_774,N_1168);
xor U2129 (N_2129,N_1229,N_1249);
or U2130 (N_2130,N_906,N_1014);
xor U2131 (N_2131,N_1006,N_1288);
or U2132 (N_2132,N_761,N_1436);
and U2133 (N_2133,N_821,N_1243);
nand U2134 (N_2134,N_1019,N_944);
and U2135 (N_2135,N_1023,N_934);
nand U2136 (N_2136,N_896,N_925);
nand U2137 (N_2137,N_1452,N_1049);
or U2138 (N_2138,N_1134,N_793);
nand U2139 (N_2139,N_1410,N_1198);
nor U2140 (N_2140,N_1401,N_1446);
xnor U2141 (N_2141,N_1022,N_1432);
nor U2142 (N_2142,N_1355,N_1412);
xor U2143 (N_2143,N_932,N_1290);
or U2144 (N_2144,N_1096,N_1203);
and U2145 (N_2145,N_1257,N_1229);
nor U2146 (N_2146,N_1412,N_781);
xor U2147 (N_2147,N_982,N_1272);
nand U2148 (N_2148,N_1023,N_1415);
nand U2149 (N_2149,N_1168,N_1116);
nor U2150 (N_2150,N_847,N_1214);
nand U2151 (N_2151,N_1453,N_870);
nand U2152 (N_2152,N_1048,N_1449);
and U2153 (N_2153,N_1120,N_1266);
nor U2154 (N_2154,N_842,N_1001);
nand U2155 (N_2155,N_1495,N_1490);
and U2156 (N_2156,N_906,N_1019);
nand U2157 (N_2157,N_1415,N_1120);
xnor U2158 (N_2158,N_1094,N_1455);
xnor U2159 (N_2159,N_953,N_1431);
xnor U2160 (N_2160,N_1181,N_1223);
nand U2161 (N_2161,N_858,N_795);
xnor U2162 (N_2162,N_973,N_929);
or U2163 (N_2163,N_1283,N_1112);
nor U2164 (N_2164,N_1137,N_1295);
xnor U2165 (N_2165,N_1378,N_890);
nor U2166 (N_2166,N_1022,N_1088);
nor U2167 (N_2167,N_769,N_1281);
nor U2168 (N_2168,N_1209,N_799);
nand U2169 (N_2169,N_1445,N_1346);
nand U2170 (N_2170,N_907,N_1494);
and U2171 (N_2171,N_1023,N_1098);
and U2172 (N_2172,N_1339,N_836);
or U2173 (N_2173,N_1035,N_1003);
xor U2174 (N_2174,N_770,N_760);
xnor U2175 (N_2175,N_1097,N_856);
or U2176 (N_2176,N_1026,N_1248);
or U2177 (N_2177,N_1018,N_899);
and U2178 (N_2178,N_1356,N_884);
nor U2179 (N_2179,N_1428,N_1306);
nand U2180 (N_2180,N_781,N_1175);
xor U2181 (N_2181,N_1367,N_837);
and U2182 (N_2182,N_1225,N_963);
and U2183 (N_2183,N_927,N_865);
or U2184 (N_2184,N_849,N_1213);
nand U2185 (N_2185,N_1130,N_1114);
xnor U2186 (N_2186,N_1384,N_997);
xor U2187 (N_2187,N_1066,N_932);
and U2188 (N_2188,N_801,N_1127);
nor U2189 (N_2189,N_1372,N_965);
xor U2190 (N_2190,N_935,N_885);
xor U2191 (N_2191,N_1183,N_1486);
xor U2192 (N_2192,N_886,N_1292);
and U2193 (N_2193,N_885,N_972);
nand U2194 (N_2194,N_913,N_1064);
or U2195 (N_2195,N_948,N_1148);
and U2196 (N_2196,N_752,N_833);
nor U2197 (N_2197,N_1442,N_1126);
or U2198 (N_2198,N_1229,N_866);
or U2199 (N_2199,N_1300,N_1400);
xnor U2200 (N_2200,N_906,N_1163);
nand U2201 (N_2201,N_1208,N_842);
xor U2202 (N_2202,N_1083,N_1469);
nor U2203 (N_2203,N_1337,N_793);
nand U2204 (N_2204,N_854,N_1098);
nand U2205 (N_2205,N_1192,N_1089);
nor U2206 (N_2206,N_1283,N_1460);
xnor U2207 (N_2207,N_1492,N_1218);
or U2208 (N_2208,N_1002,N_846);
xor U2209 (N_2209,N_1351,N_944);
nor U2210 (N_2210,N_798,N_763);
nand U2211 (N_2211,N_1427,N_1266);
xor U2212 (N_2212,N_1420,N_934);
nor U2213 (N_2213,N_1035,N_872);
and U2214 (N_2214,N_1253,N_1339);
xnor U2215 (N_2215,N_1049,N_1420);
nor U2216 (N_2216,N_965,N_1195);
and U2217 (N_2217,N_1442,N_891);
and U2218 (N_2218,N_1208,N_1234);
or U2219 (N_2219,N_935,N_950);
or U2220 (N_2220,N_996,N_907);
xor U2221 (N_2221,N_1229,N_1343);
nand U2222 (N_2222,N_1377,N_869);
or U2223 (N_2223,N_1343,N_1326);
xnor U2224 (N_2224,N_936,N_1273);
nand U2225 (N_2225,N_1052,N_1409);
nand U2226 (N_2226,N_1199,N_1390);
nor U2227 (N_2227,N_793,N_884);
or U2228 (N_2228,N_1379,N_1389);
or U2229 (N_2229,N_1467,N_1144);
nor U2230 (N_2230,N_987,N_1474);
xor U2231 (N_2231,N_916,N_1041);
nor U2232 (N_2232,N_1215,N_892);
or U2233 (N_2233,N_1149,N_1036);
or U2234 (N_2234,N_1290,N_1419);
or U2235 (N_2235,N_1095,N_1249);
or U2236 (N_2236,N_1421,N_1265);
or U2237 (N_2237,N_1231,N_1341);
or U2238 (N_2238,N_1328,N_1259);
or U2239 (N_2239,N_779,N_908);
and U2240 (N_2240,N_761,N_1057);
nand U2241 (N_2241,N_1113,N_1098);
or U2242 (N_2242,N_938,N_1392);
nand U2243 (N_2243,N_929,N_980);
nor U2244 (N_2244,N_1345,N_1317);
xor U2245 (N_2245,N_1255,N_1101);
and U2246 (N_2246,N_936,N_786);
or U2247 (N_2247,N_938,N_1243);
nor U2248 (N_2248,N_1183,N_1120);
xor U2249 (N_2249,N_809,N_1340);
or U2250 (N_2250,N_1860,N_1651);
and U2251 (N_2251,N_1892,N_1741);
or U2252 (N_2252,N_1996,N_1836);
nor U2253 (N_2253,N_2088,N_1762);
and U2254 (N_2254,N_1521,N_1725);
nand U2255 (N_2255,N_1753,N_1761);
and U2256 (N_2256,N_2122,N_2172);
nand U2257 (N_2257,N_2193,N_1907);
or U2258 (N_2258,N_2153,N_1712);
and U2259 (N_2259,N_1540,N_1877);
nor U2260 (N_2260,N_1891,N_2113);
and U2261 (N_2261,N_2058,N_1504);
or U2262 (N_2262,N_1642,N_2217);
xor U2263 (N_2263,N_1621,N_2069);
or U2264 (N_2264,N_1797,N_2241);
and U2265 (N_2265,N_1779,N_1803);
nor U2266 (N_2266,N_2148,N_1513);
or U2267 (N_2267,N_1850,N_1847);
and U2268 (N_2268,N_1897,N_1690);
nand U2269 (N_2269,N_2195,N_2105);
and U2270 (N_2270,N_2222,N_1695);
xnor U2271 (N_2271,N_1862,N_1856);
nand U2272 (N_2272,N_2012,N_1953);
and U2273 (N_2273,N_2084,N_1755);
nand U2274 (N_2274,N_2126,N_2001);
xor U2275 (N_2275,N_1588,N_1770);
and U2276 (N_2276,N_1631,N_1882);
and U2277 (N_2277,N_1977,N_1917);
nand U2278 (N_2278,N_1679,N_1635);
nand U2279 (N_2279,N_2213,N_1508);
or U2280 (N_2280,N_1959,N_1787);
or U2281 (N_2281,N_2067,N_1832);
or U2282 (N_2282,N_2248,N_1822);
or U2283 (N_2283,N_2235,N_2095);
xnor U2284 (N_2284,N_1763,N_1818);
and U2285 (N_2285,N_2118,N_1667);
nor U2286 (N_2286,N_2098,N_1785);
nand U2287 (N_2287,N_1782,N_1565);
nand U2288 (N_2288,N_2093,N_1937);
xnor U2289 (N_2289,N_1758,N_1826);
nand U2290 (N_2290,N_1952,N_2102);
xnor U2291 (N_2291,N_1611,N_2009);
or U2292 (N_2292,N_1967,N_1852);
xor U2293 (N_2293,N_1986,N_1825);
or U2294 (N_2294,N_2215,N_2087);
nor U2295 (N_2295,N_1881,N_1629);
nand U2296 (N_2296,N_2096,N_2013);
and U2297 (N_2297,N_1505,N_1557);
nor U2298 (N_2298,N_1678,N_1736);
or U2299 (N_2299,N_1630,N_1783);
or U2300 (N_2300,N_1872,N_1553);
nor U2301 (N_2301,N_1776,N_1926);
nor U2302 (N_2302,N_1809,N_1992);
or U2303 (N_2303,N_1805,N_1605);
xnor U2304 (N_2304,N_1824,N_1958);
and U2305 (N_2305,N_2000,N_1560);
nand U2306 (N_2306,N_1855,N_1778);
xor U2307 (N_2307,N_2233,N_1837);
and U2308 (N_2308,N_2053,N_2187);
xnor U2309 (N_2309,N_2171,N_2183);
nor U2310 (N_2310,N_1601,N_1541);
xor U2311 (N_2311,N_1893,N_1964);
or U2312 (N_2312,N_1867,N_1580);
or U2313 (N_2313,N_2236,N_1887);
xor U2314 (N_2314,N_1961,N_1931);
nor U2315 (N_2315,N_2128,N_1666);
or U2316 (N_2316,N_2040,N_1780);
nand U2317 (N_2317,N_2006,N_1752);
and U2318 (N_2318,N_2005,N_1613);
and U2319 (N_2319,N_1839,N_1890);
xnor U2320 (N_2320,N_2033,N_1791);
or U2321 (N_2321,N_1509,N_1927);
or U2322 (N_2322,N_1546,N_2054);
nor U2323 (N_2323,N_2170,N_2085);
nand U2324 (N_2324,N_1619,N_2103);
or U2325 (N_2325,N_1906,N_1547);
or U2326 (N_2326,N_1558,N_1942);
nor U2327 (N_2327,N_1863,N_1664);
and U2328 (N_2328,N_1913,N_1652);
nor U2329 (N_2329,N_1661,N_2056);
and U2330 (N_2330,N_1914,N_1561);
xnor U2331 (N_2331,N_2037,N_2201);
and U2332 (N_2332,N_1528,N_1962);
nand U2333 (N_2333,N_2240,N_1767);
nor U2334 (N_2334,N_2086,N_1811);
and U2335 (N_2335,N_1830,N_1590);
or U2336 (N_2336,N_2038,N_1639);
xor U2337 (N_2337,N_1749,N_1831);
xor U2338 (N_2338,N_1721,N_1902);
nand U2339 (N_2339,N_1555,N_2047);
nand U2340 (N_2340,N_2129,N_1771);
xnor U2341 (N_2341,N_1503,N_1754);
and U2342 (N_2342,N_2059,N_1655);
or U2343 (N_2343,N_1535,N_1674);
and U2344 (N_2344,N_1586,N_2071);
and U2345 (N_2345,N_1518,N_1781);
or U2346 (N_2346,N_1807,N_2210);
and U2347 (N_2347,N_1632,N_1742);
or U2348 (N_2348,N_1699,N_1579);
nor U2349 (N_2349,N_1599,N_1889);
and U2350 (N_2350,N_2144,N_1857);
nor U2351 (N_2351,N_2065,N_2147);
nor U2352 (N_2352,N_2208,N_2243);
xnor U2353 (N_2353,N_1979,N_1786);
and U2354 (N_2354,N_1516,N_1823);
and U2355 (N_2355,N_1724,N_1924);
nor U2356 (N_2356,N_1641,N_1600);
nor U2357 (N_2357,N_2123,N_1567);
nor U2358 (N_2358,N_1689,N_2015);
and U2359 (N_2359,N_1685,N_2036);
nand U2360 (N_2360,N_1672,N_1746);
nor U2361 (N_2361,N_1671,N_1646);
xor U2362 (N_2362,N_1829,N_1525);
or U2363 (N_2363,N_1757,N_1845);
xor U2364 (N_2364,N_1524,N_1573);
nand U2365 (N_2365,N_1769,N_2125);
and U2366 (N_2366,N_2094,N_1717);
nor U2367 (N_2367,N_1827,N_1707);
nor U2368 (N_2368,N_2074,N_1570);
and U2369 (N_2369,N_1718,N_1604);
nand U2370 (N_2370,N_1940,N_1530);
and U2371 (N_2371,N_1842,N_2112);
xor U2372 (N_2372,N_2116,N_1726);
or U2373 (N_2373,N_2200,N_1841);
nor U2374 (N_2374,N_2159,N_2081);
nor U2375 (N_2375,N_1644,N_2202);
nor U2376 (N_2376,N_1556,N_2165);
xnor U2377 (N_2377,N_2249,N_1577);
nand U2378 (N_2378,N_1676,N_1658);
xor U2379 (N_2379,N_2028,N_2162);
nor U2380 (N_2380,N_1955,N_1874);
or U2381 (N_2381,N_2152,N_1799);
nor U2382 (N_2382,N_1848,N_1909);
nand U2383 (N_2383,N_1900,N_1846);
and U2384 (N_2384,N_1812,N_1993);
and U2385 (N_2385,N_1727,N_1527);
nand U2386 (N_2386,N_1536,N_1663);
or U2387 (N_2387,N_1740,N_1988);
xor U2388 (N_2388,N_2063,N_2137);
xor U2389 (N_2389,N_2055,N_1574);
or U2390 (N_2390,N_1720,N_1697);
or U2391 (N_2391,N_1933,N_2072);
or U2392 (N_2392,N_1859,N_1999);
xnor U2393 (N_2393,N_1572,N_1735);
xnor U2394 (N_2394,N_2029,N_1972);
xor U2395 (N_2395,N_1617,N_1792);
nor U2396 (N_2396,N_1719,N_2238);
or U2397 (N_2397,N_1968,N_2083);
nor U2398 (N_2398,N_1539,N_2130);
xor U2399 (N_2399,N_2043,N_2117);
or U2400 (N_2400,N_1878,N_2226);
nor U2401 (N_2401,N_1563,N_1606);
and U2402 (N_2402,N_1510,N_1665);
nor U2403 (N_2403,N_1957,N_2207);
xor U2404 (N_2404,N_2078,N_1981);
nor U2405 (N_2405,N_1934,N_1815);
xnor U2406 (N_2406,N_1948,N_1515);
and U2407 (N_2407,N_2016,N_1844);
xnor U2408 (N_2408,N_2034,N_2120);
nand U2409 (N_2409,N_2035,N_1552);
nand U2410 (N_2410,N_1533,N_1798);
nand U2411 (N_2411,N_2014,N_1835);
or U2412 (N_2412,N_2057,N_2214);
nand U2413 (N_2413,N_1512,N_1597);
nand U2414 (N_2414,N_2149,N_1703);
xnor U2415 (N_2415,N_2090,N_1582);
nor U2416 (N_2416,N_2164,N_1609);
xor U2417 (N_2417,N_2030,N_2218);
nor U2418 (N_2418,N_2099,N_1589);
and U2419 (N_2419,N_2163,N_1559);
nor U2420 (N_2420,N_1594,N_2019);
or U2421 (N_2421,N_2133,N_1947);
nand U2422 (N_2422,N_1828,N_1616);
nor U2423 (N_2423,N_2157,N_1696);
nor U2424 (N_2424,N_2230,N_1708);
or U2425 (N_2425,N_2111,N_1866);
nor U2426 (N_2426,N_1669,N_1593);
xor U2427 (N_2427,N_2139,N_1675);
and U2428 (N_2428,N_2184,N_1873);
or U2429 (N_2429,N_1784,N_1946);
or U2430 (N_2430,N_1983,N_1875);
nand U2431 (N_2431,N_2168,N_1994);
nor U2432 (N_2432,N_2176,N_1500);
and U2433 (N_2433,N_2050,N_2108);
or U2434 (N_2434,N_1715,N_1583);
xnor U2435 (N_2435,N_1905,N_2242);
or U2436 (N_2436,N_2150,N_1728);
xnor U2437 (N_2437,N_1894,N_1932);
xnor U2438 (N_2438,N_1965,N_1941);
or U2439 (N_2439,N_1640,N_1908);
nand U2440 (N_2440,N_1864,N_1548);
and U2441 (N_2441,N_2190,N_1939);
or U2442 (N_2442,N_2064,N_2179);
xnor U2443 (N_2443,N_2232,N_1918);
xor U2444 (N_2444,N_1998,N_2075);
or U2445 (N_2445,N_2045,N_1865);
or U2446 (N_2446,N_1789,N_1562);
or U2447 (N_2447,N_1929,N_1649);
nand U2448 (N_2448,N_1969,N_2008);
and U2449 (N_2449,N_1680,N_2141);
or U2450 (N_2450,N_2219,N_2227);
xor U2451 (N_2451,N_1743,N_2181);
nand U2452 (N_2452,N_1544,N_2178);
nor U2453 (N_2453,N_1615,N_1529);
and U2454 (N_2454,N_1796,N_2132);
nor U2455 (N_2455,N_1648,N_1756);
and U2456 (N_2456,N_1634,N_2155);
nor U2457 (N_2457,N_1569,N_1705);
xor U2458 (N_2458,N_1884,N_1820);
and U2459 (N_2459,N_1816,N_1911);
nand U2460 (N_2460,N_1534,N_1773);
and U2461 (N_2461,N_1903,N_1571);
or U2462 (N_2462,N_1975,N_1899);
or U2463 (N_2463,N_1537,N_1885);
xnor U2464 (N_2464,N_2203,N_1700);
and U2465 (N_2465,N_1738,N_1576);
nor U2466 (N_2466,N_1950,N_1603);
nand U2467 (N_2467,N_2046,N_1625);
or U2468 (N_2468,N_2092,N_1764);
nand U2469 (N_2469,N_2191,N_2231);
or U2470 (N_2470,N_1624,N_1984);
nor U2471 (N_2471,N_1990,N_2107);
xnor U2472 (N_2472,N_2049,N_1714);
or U2473 (N_2473,N_1788,N_1880);
or U2474 (N_2474,N_1944,N_1922);
nand U2475 (N_2475,N_1732,N_2221);
nor U2476 (N_2476,N_1722,N_1662);
xor U2477 (N_2477,N_1550,N_1925);
nor U2478 (N_2478,N_1843,N_2166);
or U2479 (N_2479,N_1978,N_2022);
or U2480 (N_2480,N_2089,N_1748);
nor U2481 (N_2481,N_2077,N_2127);
nor U2482 (N_2482,N_1821,N_1733);
or U2483 (N_2483,N_1538,N_2110);
xnor U2484 (N_2484,N_1945,N_1686);
nor U2485 (N_2485,N_1916,N_1854);
nand U2486 (N_2486,N_1989,N_1760);
nand U2487 (N_2487,N_2194,N_1688);
and U2488 (N_2488,N_1858,N_1973);
xor U2489 (N_2489,N_2025,N_1888);
nor U2490 (N_2490,N_1731,N_1568);
nor U2491 (N_2491,N_1653,N_1677);
nand U2492 (N_2492,N_2018,N_1694);
xor U2493 (N_2493,N_2229,N_2039);
and U2494 (N_2494,N_2114,N_2091);
or U2495 (N_2495,N_1520,N_1526);
nand U2496 (N_2496,N_2121,N_1706);
nor U2497 (N_2497,N_2234,N_1711);
and U2498 (N_2498,N_1930,N_1620);
nor U2499 (N_2499,N_1692,N_2156);
nand U2500 (N_2500,N_1943,N_2115);
or U2501 (N_2501,N_1869,N_2196);
and U2502 (N_2502,N_1592,N_1584);
nor U2503 (N_2503,N_2188,N_1612);
nand U2504 (N_2504,N_1921,N_1519);
or U2505 (N_2505,N_1701,N_1982);
and U2506 (N_2506,N_1531,N_2158);
and U2507 (N_2507,N_2101,N_1564);
nand U2508 (N_2508,N_1750,N_1628);
nand U2509 (N_2509,N_2192,N_2223);
xor U2510 (N_2510,N_1581,N_1853);
nor U2511 (N_2511,N_1507,N_2204);
nor U2512 (N_2512,N_1804,N_1633);
or U2513 (N_2513,N_1623,N_1775);
and U2514 (N_2514,N_1956,N_1506);
nor U2515 (N_2515,N_1660,N_2066);
and U2516 (N_2516,N_1595,N_2174);
nand U2517 (N_2517,N_1768,N_2104);
nor U2518 (N_2518,N_1607,N_1814);
nor U2519 (N_2519,N_1650,N_1627);
or U2520 (N_2520,N_1951,N_2070);
nand U2521 (N_2521,N_1502,N_2020);
nand U2522 (N_2522,N_1614,N_1673);
and U2523 (N_2523,N_2185,N_1554);
nand U2524 (N_2524,N_2205,N_2175);
nand U2525 (N_2525,N_1643,N_1729);
or U2526 (N_2526,N_1517,N_1920);
nand U2527 (N_2527,N_2052,N_1793);
nand U2528 (N_2528,N_1549,N_2044);
xor U2529 (N_2529,N_2209,N_2142);
nand U2530 (N_2530,N_2182,N_2180);
or U2531 (N_2531,N_1511,N_1591);
nand U2532 (N_2532,N_2011,N_2220);
and U2533 (N_2533,N_2146,N_2027);
nand U2534 (N_2534,N_1849,N_1684);
nor U2535 (N_2535,N_1682,N_2051);
or U2536 (N_2536,N_1954,N_2212);
nor U2537 (N_2537,N_1834,N_1737);
nand U2538 (N_2538,N_1896,N_1985);
xnor U2539 (N_2539,N_1543,N_1710);
nand U2540 (N_2540,N_1980,N_1626);
xor U2541 (N_2541,N_1716,N_2004);
nand U2542 (N_2542,N_2177,N_2068);
nor U2543 (N_2543,N_1681,N_2237);
nand U2544 (N_2544,N_2073,N_1868);
nor U2545 (N_2545,N_1702,N_1575);
and U2546 (N_2546,N_1801,N_2145);
nand U2547 (N_2547,N_1870,N_1687);
and U2548 (N_2548,N_1545,N_1838);
or U2549 (N_2549,N_1654,N_2173);
nor U2550 (N_2550,N_1514,N_1659);
and U2551 (N_2551,N_1523,N_2106);
xnor U2552 (N_2552,N_1766,N_1883);
nor U2553 (N_2553,N_1808,N_2245);
nand U2554 (N_2554,N_1645,N_1657);
and U2555 (N_2555,N_1904,N_2062);
nor U2556 (N_2556,N_1970,N_1886);
and U2557 (N_2557,N_2143,N_1794);
nor U2558 (N_2558,N_1795,N_1532);
and U2559 (N_2559,N_1598,N_1585);
xnor U2560 (N_2560,N_1637,N_1861);
nor U2561 (N_2561,N_2109,N_2080);
xnor U2562 (N_2562,N_1963,N_1895);
xnor U2563 (N_2563,N_2206,N_1691);
or U2564 (N_2564,N_1713,N_1810);
or U2565 (N_2565,N_1851,N_1723);
and U2566 (N_2566,N_2160,N_2197);
xor U2567 (N_2567,N_1683,N_2079);
xnor U2568 (N_2568,N_1935,N_2239);
nand U2569 (N_2569,N_1739,N_1747);
nand U2570 (N_2570,N_1876,N_2031);
or U2571 (N_2571,N_1777,N_1813);
nand U2572 (N_2572,N_1938,N_2124);
xor U2573 (N_2573,N_1704,N_2097);
nor U2574 (N_2574,N_2189,N_1596);
xor U2575 (N_2575,N_1790,N_1730);
or U2576 (N_2576,N_1772,N_1608);
nor U2577 (N_2577,N_1578,N_1910);
or U2578 (N_2578,N_1636,N_2024);
xor U2579 (N_2579,N_1551,N_1936);
or U2580 (N_2580,N_1976,N_2003);
or U2581 (N_2581,N_2225,N_2198);
nand U2582 (N_2582,N_2154,N_2131);
nor U2583 (N_2583,N_1871,N_2021);
and U2584 (N_2584,N_1734,N_2246);
nor U2585 (N_2585,N_1522,N_1709);
or U2586 (N_2586,N_1602,N_2002);
nor U2587 (N_2587,N_2169,N_1802);
or U2588 (N_2588,N_1693,N_1668);
nor U2589 (N_2589,N_1923,N_2136);
nand U2590 (N_2590,N_2041,N_1618);
nor U2591 (N_2591,N_1587,N_2186);
nor U2592 (N_2592,N_1919,N_1638);
or U2593 (N_2593,N_1647,N_1759);
nor U2594 (N_2594,N_1960,N_2082);
and U2595 (N_2595,N_1774,N_2140);
nand U2596 (N_2596,N_2247,N_2211);
nor U2597 (N_2597,N_2026,N_1840);
nor U2598 (N_2598,N_1991,N_1698);
xor U2599 (N_2599,N_2151,N_2228);
and U2600 (N_2600,N_2244,N_1898);
nor U2601 (N_2601,N_1966,N_1949);
or U2602 (N_2602,N_1670,N_2010);
nand U2603 (N_2603,N_1997,N_2100);
nand U2604 (N_2604,N_1656,N_1806);
xnor U2605 (N_2605,N_2224,N_2023);
nor U2606 (N_2606,N_1622,N_1928);
nor U2607 (N_2607,N_1765,N_1915);
nor U2608 (N_2608,N_1610,N_1800);
xnor U2609 (N_2609,N_2060,N_1566);
xor U2610 (N_2610,N_1501,N_1995);
or U2611 (N_2611,N_2161,N_2042);
or U2612 (N_2612,N_2032,N_1751);
xor U2613 (N_2613,N_1817,N_2199);
nor U2614 (N_2614,N_1542,N_2061);
or U2615 (N_2615,N_1971,N_2048);
xnor U2616 (N_2616,N_1819,N_1987);
xor U2617 (N_2617,N_2134,N_2216);
or U2618 (N_2618,N_2076,N_1912);
and U2619 (N_2619,N_2017,N_1901);
nor U2620 (N_2620,N_1833,N_2135);
xor U2621 (N_2621,N_1745,N_2007);
nor U2622 (N_2622,N_2167,N_1744);
nor U2623 (N_2623,N_1974,N_1879);
nor U2624 (N_2624,N_2119,N_2138);
nor U2625 (N_2625,N_1695,N_1926);
xor U2626 (N_2626,N_1679,N_1663);
nand U2627 (N_2627,N_1558,N_1707);
and U2628 (N_2628,N_2164,N_1618);
nor U2629 (N_2629,N_2166,N_2000);
nand U2630 (N_2630,N_2126,N_1968);
xor U2631 (N_2631,N_2054,N_1942);
and U2632 (N_2632,N_2179,N_2191);
or U2633 (N_2633,N_2242,N_1859);
nor U2634 (N_2634,N_1959,N_1691);
xor U2635 (N_2635,N_1634,N_2101);
or U2636 (N_2636,N_2233,N_1501);
nor U2637 (N_2637,N_1671,N_1941);
nor U2638 (N_2638,N_2136,N_1690);
and U2639 (N_2639,N_2242,N_1773);
xnor U2640 (N_2640,N_1901,N_2056);
nand U2641 (N_2641,N_1540,N_1737);
nand U2642 (N_2642,N_2021,N_2119);
nor U2643 (N_2643,N_2094,N_1719);
and U2644 (N_2644,N_1733,N_1627);
and U2645 (N_2645,N_2050,N_1725);
xnor U2646 (N_2646,N_1578,N_1905);
xnor U2647 (N_2647,N_2007,N_2189);
or U2648 (N_2648,N_1646,N_1617);
and U2649 (N_2649,N_1874,N_2019);
and U2650 (N_2650,N_1825,N_1934);
nor U2651 (N_2651,N_1889,N_1866);
or U2652 (N_2652,N_1707,N_1578);
or U2653 (N_2653,N_1770,N_1576);
nand U2654 (N_2654,N_1755,N_2066);
or U2655 (N_2655,N_1517,N_2226);
and U2656 (N_2656,N_2124,N_2067);
nand U2657 (N_2657,N_1925,N_1992);
nand U2658 (N_2658,N_1629,N_1783);
nor U2659 (N_2659,N_1964,N_1951);
or U2660 (N_2660,N_2067,N_1660);
and U2661 (N_2661,N_1569,N_2073);
nand U2662 (N_2662,N_1763,N_1787);
and U2663 (N_2663,N_2219,N_2216);
xnor U2664 (N_2664,N_2053,N_1619);
nand U2665 (N_2665,N_1826,N_1972);
or U2666 (N_2666,N_1560,N_2024);
nand U2667 (N_2667,N_1933,N_1881);
nand U2668 (N_2668,N_1979,N_1981);
and U2669 (N_2669,N_2120,N_1883);
nor U2670 (N_2670,N_2218,N_2054);
nand U2671 (N_2671,N_1965,N_1874);
nand U2672 (N_2672,N_2006,N_1936);
or U2673 (N_2673,N_2085,N_2063);
and U2674 (N_2674,N_2243,N_1830);
xnor U2675 (N_2675,N_1924,N_1901);
xnor U2676 (N_2676,N_1701,N_2196);
and U2677 (N_2677,N_1922,N_2190);
xnor U2678 (N_2678,N_2220,N_1930);
and U2679 (N_2679,N_1507,N_1596);
and U2680 (N_2680,N_1701,N_1984);
nor U2681 (N_2681,N_2087,N_1935);
and U2682 (N_2682,N_2182,N_1774);
nand U2683 (N_2683,N_1762,N_1696);
or U2684 (N_2684,N_1835,N_2096);
and U2685 (N_2685,N_1805,N_1928);
or U2686 (N_2686,N_1836,N_1543);
nand U2687 (N_2687,N_2221,N_1877);
xnor U2688 (N_2688,N_1867,N_1956);
or U2689 (N_2689,N_2029,N_1728);
nor U2690 (N_2690,N_1667,N_2105);
xor U2691 (N_2691,N_2217,N_1686);
and U2692 (N_2692,N_2113,N_2162);
or U2693 (N_2693,N_2147,N_1736);
and U2694 (N_2694,N_1747,N_2143);
nor U2695 (N_2695,N_1805,N_1681);
xor U2696 (N_2696,N_2225,N_2011);
nand U2697 (N_2697,N_2024,N_2044);
or U2698 (N_2698,N_1562,N_1792);
nand U2699 (N_2699,N_2061,N_1979);
nand U2700 (N_2700,N_2233,N_1757);
nor U2701 (N_2701,N_1712,N_2000);
and U2702 (N_2702,N_1773,N_2020);
or U2703 (N_2703,N_1780,N_2107);
or U2704 (N_2704,N_1966,N_1504);
and U2705 (N_2705,N_1748,N_1863);
xnor U2706 (N_2706,N_1811,N_2009);
nand U2707 (N_2707,N_1509,N_2094);
xor U2708 (N_2708,N_2107,N_2193);
and U2709 (N_2709,N_1966,N_2072);
nand U2710 (N_2710,N_1566,N_1915);
nand U2711 (N_2711,N_1666,N_2086);
xnor U2712 (N_2712,N_1940,N_1678);
and U2713 (N_2713,N_1702,N_1747);
or U2714 (N_2714,N_2077,N_1705);
nor U2715 (N_2715,N_1700,N_2008);
xor U2716 (N_2716,N_1788,N_1585);
nand U2717 (N_2717,N_1774,N_1719);
and U2718 (N_2718,N_1817,N_1526);
or U2719 (N_2719,N_1990,N_1770);
nor U2720 (N_2720,N_1904,N_1879);
and U2721 (N_2721,N_2031,N_1999);
xor U2722 (N_2722,N_1523,N_1909);
xor U2723 (N_2723,N_2224,N_1532);
nand U2724 (N_2724,N_2187,N_1804);
nor U2725 (N_2725,N_1575,N_1969);
xor U2726 (N_2726,N_1929,N_2093);
and U2727 (N_2727,N_2137,N_2184);
and U2728 (N_2728,N_1722,N_1503);
or U2729 (N_2729,N_1757,N_1771);
xor U2730 (N_2730,N_2183,N_1722);
nor U2731 (N_2731,N_1963,N_1692);
xor U2732 (N_2732,N_1963,N_1794);
nor U2733 (N_2733,N_1738,N_2020);
or U2734 (N_2734,N_1906,N_2170);
and U2735 (N_2735,N_2078,N_2154);
nor U2736 (N_2736,N_1585,N_1552);
and U2737 (N_2737,N_2136,N_1904);
and U2738 (N_2738,N_1527,N_1842);
xor U2739 (N_2739,N_2163,N_1780);
and U2740 (N_2740,N_1610,N_1607);
and U2741 (N_2741,N_2014,N_2158);
and U2742 (N_2742,N_2117,N_1871);
xor U2743 (N_2743,N_1717,N_1636);
and U2744 (N_2744,N_2027,N_1973);
nand U2745 (N_2745,N_2015,N_1644);
or U2746 (N_2746,N_2058,N_1824);
nand U2747 (N_2747,N_2078,N_1616);
and U2748 (N_2748,N_2230,N_1777);
or U2749 (N_2749,N_2114,N_2008);
xor U2750 (N_2750,N_1905,N_1509);
nand U2751 (N_2751,N_1800,N_1726);
or U2752 (N_2752,N_2241,N_2105);
and U2753 (N_2753,N_1742,N_1811);
nor U2754 (N_2754,N_2059,N_2068);
xnor U2755 (N_2755,N_1950,N_1719);
or U2756 (N_2756,N_2149,N_1889);
nand U2757 (N_2757,N_1864,N_2153);
or U2758 (N_2758,N_2175,N_2182);
and U2759 (N_2759,N_2123,N_1587);
or U2760 (N_2760,N_1872,N_1730);
xor U2761 (N_2761,N_2246,N_1789);
nand U2762 (N_2762,N_1736,N_1502);
nor U2763 (N_2763,N_1721,N_1804);
nor U2764 (N_2764,N_1991,N_1663);
xor U2765 (N_2765,N_1514,N_2122);
nand U2766 (N_2766,N_1724,N_2233);
nor U2767 (N_2767,N_1628,N_1673);
or U2768 (N_2768,N_1594,N_1677);
xor U2769 (N_2769,N_1528,N_1607);
or U2770 (N_2770,N_2023,N_1644);
nor U2771 (N_2771,N_1555,N_1979);
nand U2772 (N_2772,N_2077,N_1843);
and U2773 (N_2773,N_1580,N_1998);
or U2774 (N_2774,N_2225,N_1773);
nor U2775 (N_2775,N_1995,N_1982);
nand U2776 (N_2776,N_2211,N_1812);
nor U2777 (N_2777,N_1833,N_1806);
nand U2778 (N_2778,N_1704,N_1872);
xnor U2779 (N_2779,N_2064,N_1817);
or U2780 (N_2780,N_2093,N_1646);
xor U2781 (N_2781,N_2178,N_1577);
nand U2782 (N_2782,N_1571,N_1816);
xnor U2783 (N_2783,N_1955,N_1893);
nand U2784 (N_2784,N_2163,N_1534);
nand U2785 (N_2785,N_1886,N_2199);
and U2786 (N_2786,N_2104,N_2163);
nor U2787 (N_2787,N_1618,N_1996);
nand U2788 (N_2788,N_2239,N_2228);
and U2789 (N_2789,N_2009,N_1989);
xnor U2790 (N_2790,N_1549,N_2224);
and U2791 (N_2791,N_2085,N_1697);
nor U2792 (N_2792,N_1627,N_2151);
nor U2793 (N_2793,N_2172,N_2030);
nand U2794 (N_2794,N_2197,N_1921);
nor U2795 (N_2795,N_1517,N_1942);
xor U2796 (N_2796,N_2091,N_1646);
or U2797 (N_2797,N_1641,N_1745);
nor U2798 (N_2798,N_1976,N_1565);
nand U2799 (N_2799,N_2238,N_1940);
or U2800 (N_2800,N_2103,N_1855);
nand U2801 (N_2801,N_2081,N_1721);
or U2802 (N_2802,N_1914,N_1732);
nor U2803 (N_2803,N_2123,N_1575);
xnor U2804 (N_2804,N_2037,N_1923);
nor U2805 (N_2805,N_2229,N_1745);
nand U2806 (N_2806,N_2136,N_1807);
nor U2807 (N_2807,N_1726,N_2169);
nor U2808 (N_2808,N_1739,N_1688);
xnor U2809 (N_2809,N_2215,N_2226);
and U2810 (N_2810,N_1884,N_1719);
xnor U2811 (N_2811,N_1752,N_2234);
xnor U2812 (N_2812,N_2095,N_1744);
nand U2813 (N_2813,N_1645,N_1567);
xor U2814 (N_2814,N_2248,N_1846);
nor U2815 (N_2815,N_1863,N_1956);
and U2816 (N_2816,N_1767,N_1530);
and U2817 (N_2817,N_2078,N_2018);
nand U2818 (N_2818,N_2233,N_1925);
or U2819 (N_2819,N_1723,N_1512);
nand U2820 (N_2820,N_1988,N_1656);
or U2821 (N_2821,N_2105,N_1582);
nand U2822 (N_2822,N_2097,N_1759);
xnor U2823 (N_2823,N_1619,N_2054);
xor U2824 (N_2824,N_1623,N_1638);
and U2825 (N_2825,N_1743,N_2158);
nand U2826 (N_2826,N_2005,N_1838);
xor U2827 (N_2827,N_1840,N_2242);
and U2828 (N_2828,N_1714,N_1751);
or U2829 (N_2829,N_1963,N_2069);
xor U2830 (N_2830,N_1791,N_1602);
nand U2831 (N_2831,N_1721,N_2042);
nand U2832 (N_2832,N_1992,N_1792);
nor U2833 (N_2833,N_2064,N_2033);
and U2834 (N_2834,N_1727,N_2235);
xnor U2835 (N_2835,N_1840,N_1885);
nor U2836 (N_2836,N_1920,N_1696);
xnor U2837 (N_2837,N_1730,N_2057);
and U2838 (N_2838,N_2175,N_1764);
and U2839 (N_2839,N_1773,N_1994);
or U2840 (N_2840,N_2037,N_1734);
nand U2841 (N_2841,N_1503,N_2185);
and U2842 (N_2842,N_2166,N_2167);
xor U2843 (N_2843,N_1631,N_2242);
or U2844 (N_2844,N_2043,N_1731);
or U2845 (N_2845,N_1528,N_1930);
and U2846 (N_2846,N_2156,N_2032);
nand U2847 (N_2847,N_1719,N_1558);
nand U2848 (N_2848,N_1751,N_1922);
xnor U2849 (N_2849,N_1899,N_1820);
or U2850 (N_2850,N_1577,N_1504);
nand U2851 (N_2851,N_2166,N_1824);
nor U2852 (N_2852,N_1945,N_1972);
or U2853 (N_2853,N_2060,N_2100);
nor U2854 (N_2854,N_1563,N_2208);
nor U2855 (N_2855,N_2137,N_1509);
nand U2856 (N_2856,N_1833,N_2090);
xor U2857 (N_2857,N_1503,N_1641);
nand U2858 (N_2858,N_1978,N_1550);
nor U2859 (N_2859,N_1529,N_2056);
nand U2860 (N_2860,N_1725,N_1720);
nand U2861 (N_2861,N_1550,N_1623);
nand U2862 (N_2862,N_2051,N_1515);
and U2863 (N_2863,N_1947,N_2126);
or U2864 (N_2864,N_1916,N_1900);
nand U2865 (N_2865,N_1642,N_1961);
and U2866 (N_2866,N_1570,N_2235);
or U2867 (N_2867,N_2091,N_2010);
xnor U2868 (N_2868,N_1644,N_1832);
or U2869 (N_2869,N_1708,N_1539);
and U2870 (N_2870,N_1865,N_1804);
nand U2871 (N_2871,N_2055,N_1989);
xor U2872 (N_2872,N_2005,N_2044);
nand U2873 (N_2873,N_2243,N_1951);
or U2874 (N_2874,N_1822,N_1972);
nand U2875 (N_2875,N_2220,N_2131);
or U2876 (N_2876,N_1619,N_2146);
nand U2877 (N_2877,N_1579,N_1895);
or U2878 (N_2878,N_2101,N_2067);
nor U2879 (N_2879,N_2139,N_1760);
or U2880 (N_2880,N_1622,N_1704);
nand U2881 (N_2881,N_1808,N_1948);
or U2882 (N_2882,N_1804,N_1834);
or U2883 (N_2883,N_1601,N_1531);
or U2884 (N_2884,N_1702,N_1617);
xor U2885 (N_2885,N_2014,N_1764);
xnor U2886 (N_2886,N_1806,N_1910);
nand U2887 (N_2887,N_2085,N_2062);
nor U2888 (N_2888,N_1565,N_2067);
nand U2889 (N_2889,N_1901,N_1685);
or U2890 (N_2890,N_2236,N_2221);
and U2891 (N_2891,N_1665,N_2140);
xor U2892 (N_2892,N_1554,N_1783);
and U2893 (N_2893,N_2014,N_1889);
nand U2894 (N_2894,N_1585,N_1556);
or U2895 (N_2895,N_1727,N_1617);
nand U2896 (N_2896,N_1843,N_1602);
xnor U2897 (N_2897,N_1927,N_1780);
nor U2898 (N_2898,N_2166,N_2175);
or U2899 (N_2899,N_2174,N_1775);
nand U2900 (N_2900,N_1978,N_1579);
nor U2901 (N_2901,N_1721,N_1955);
and U2902 (N_2902,N_1585,N_1703);
and U2903 (N_2903,N_1692,N_2112);
nand U2904 (N_2904,N_1794,N_1687);
and U2905 (N_2905,N_2045,N_1701);
or U2906 (N_2906,N_1688,N_1734);
and U2907 (N_2907,N_2015,N_1759);
nor U2908 (N_2908,N_1866,N_2037);
or U2909 (N_2909,N_2176,N_1550);
nand U2910 (N_2910,N_2020,N_1836);
or U2911 (N_2911,N_2171,N_2173);
or U2912 (N_2912,N_1860,N_1982);
or U2913 (N_2913,N_1984,N_2235);
xor U2914 (N_2914,N_1800,N_1784);
nor U2915 (N_2915,N_1733,N_1685);
nand U2916 (N_2916,N_1511,N_2209);
nand U2917 (N_2917,N_1931,N_1649);
or U2918 (N_2918,N_1931,N_1504);
and U2919 (N_2919,N_2117,N_2106);
nand U2920 (N_2920,N_1599,N_1575);
or U2921 (N_2921,N_1721,N_1601);
nor U2922 (N_2922,N_2000,N_1782);
or U2923 (N_2923,N_2060,N_2066);
or U2924 (N_2924,N_2204,N_2193);
nand U2925 (N_2925,N_1588,N_2156);
nand U2926 (N_2926,N_1520,N_1765);
xor U2927 (N_2927,N_1978,N_1544);
xnor U2928 (N_2928,N_2248,N_1972);
or U2929 (N_2929,N_1955,N_2221);
or U2930 (N_2930,N_1614,N_1715);
or U2931 (N_2931,N_1715,N_1934);
nor U2932 (N_2932,N_1663,N_1777);
and U2933 (N_2933,N_2152,N_1911);
or U2934 (N_2934,N_1626,N_2193);
xnor U2935 (N_2935,N_1734,N_1543);
xor U2936 (N_2936,N_1956,N_2059);
xnor U2937 (N_2937,N_1584,N_1924);
nand U2938 (N_2938,N_2075,N_2082);
nor U2939 (N_2939,N_1620,N_1710);
nor U2940 (N_2940,N_1501,N_2075);
nand U2941 (N_2941,N_1817,N_2014);
nand U2942 (N_2942,N_1875,N_2140);
nor U2943 (N_2943,N_2146,N_2009);
nor U2944 (N_2944,N_1855,N_1556);
or U2945 (N_2945,N_2093,N_1575);
nand U2946 (N_2946,N_2168,N_1695);
nand U2947 (N_2947,N_1619,N_1910);
or U2948 (N_2948,N_1896,N_1576);
and U2949 (N_2949,N_1564,N_1827);
nor U2950 (N_2950,N_2096,N_2136);
nand U2951 (N_2951,N_2170,N_1518);
or U2952 (N_2952,N_2095,N_2078);
and U2953 (N_2953,N_1994,N_2234);
or U2954 (N_2954,N_2211,N_2078);
and U2955 (N_2955,N_2082,N_1643);
and U2956 (N_2956,N_2077,N_2069);
nand U2957 (N_2957,N_1567,N_2172);
nand U2958 (N_2958,N_1903,N_1734);
and U2959 (N_2959,N_1618,N_2230);
or U2960 (N_2960,N_2240,N_2223);
nand U2961 (N_2961,N_2102,N_1760);
xor U2962 (N_2962,N_1782,N_2171);
and U2963 (N_2963,N_1758,N_1840);
nand U2964 (N_2964,N_1552,N_2016);
or U2965 (N_2965,N_2204,N_2143);
or U2966 (N_2966,N_2091,N_1914);
xor U2967 (N_2967,N_1536,N_1808);
nand U2968 (N_2968,N_1592,N_2177);
nand U2969 (N_2969,N_1685,N_2243);
nand U2970 (N_2970,N_1746,N_2003);
nor U2971 (N_2971,N_1597,N_2027);
xnor U2972 (N_2972,N_1957,N_1605);
nand U2973 (N_2973,N_1874,N_2021);
or U2974 (N_2974,N_2099,N_2009);
nand U2975 (N_2975,N_2091,N_1682);
or U2976 (N_2976,N_2165,N_2094);
nor U2977 (N_2977,N_1998,N_1548);
and U2978 (N_2978,N_1569,N_1775);
xnor U2979 (N_2979,N_1507,N_1919);
xnor U2980 (N_2980,N_1509,N_1769);
and U2981 (N_2981,N_2186,N_1958);
nand U2982 (N_2982,N_2230,N_1757);
nand U2983 (N_2983,N_2060,N_1772);
or U2984 (N_2984,N_1900,N_1711);
and U2985 (N_2985,N_1782,N_2223);
or U2986 (N_2986,N_1632,N_1990);
xnor U2987 (N_2987,N_1853,N_1868);
xor U2988 (N_2988,N_1872,N_1761);
and U2989 (N_2989,N_1763,N_1700);
xor U2990 (N_2990,N_1741,N_1666);
and U2991 (N_2991,N_2002,N_1675);
or U2992 (N_2992,N_2045,N_1908);
xnor U2993 (N_2993,N_1610,N_2208);
nand U2994 (N_2994,N_1956,N_2208);
nor U2995 (N_2995,N_1876,N_1804);
xnor U2996 (N_2996,N_1932,N_1946);
nand U2997 (N_2997,N_2015,N_1790);
nor U2998 (N_2998,N_2130,N_1790);
and U2999 (N_2999,N_1548,N_1908);
and U3000 (N_3000,N_2924,N_2748);
xnor U3001 (N_3001,N_2979,N_2600);
xor U3002 (N_3002,N_2736,N_2549);
or U3003 (N_3003,N_2268,N_2663);
nand U3004 (N_3004,N_2839,N_2881);
nor U3005 (N_3005,N_2260,N_2726);
and U3006 (N_3006,N_2838,N_2576);
nor U3007 (N_3007,N_2303,N_2717);
xnor U3008 (N_3008,N_2781,N_2400);
nand U3009 (N_3009,N_2930,N_2564);
nor U3010 (N_3010,N_2493,N_2842);
xnor U3011 (N_3011,N_2585,N_2262);
or U3012 (N_3012,N_2476,N_2652);
nand U3013 (N_3013,N_2933,N_2886);
xor U3014 (N_3014,N_2811,N_2478);
nand U3015 (N_3015,N_2257,N_2932);
xor U3016 (N_3016,N_2584,N_2951);
nand U3017 (N_3017,N_2700,N_2337);
xnor U3018 (N_3018,N_2441,N_2383);
xnor U3019 (N_3019,N_2821,N_2800);
nor U3020 (N_3020,N_2361,N_2386);
nor U3021 (N_3021,N_2854,N_2690);
xnor U3022 (N_3022,N_2485,N_2940);
nor U3023 (N_3023,N_2798,N_2752);
xor U3024 (N_3024,N_2624,N_2285);
nand U3025 (N_3025,N_2435,N_2484);
and U3026 (N_3026,N_2947,N_2394);
or U3027 (N_3027,N_2482,N_2500);
xnor U3028 (N_3028,N_2462,N_2844);
nand U3029 (N_3029,N_2437,N_2346);
nand U3030 (N_3030,N_2864,N_2675);
nor U3031 (N_3031,N_2751,N_2292);
or U3032 (N_3032,N_2625,N_2643);
and U3033 (N_3033,N_2352,N_2342);
nand U3034 (N_3034,N_2450,N_2290);
nand U3035 (N_3035,N_2962,N_2531);
xnor U3036 (N_3036,N_2742,N_2826);
nor U3037 (N_3037,N_2714,N_2323);
and U3038 (N_3038,N_2703,N_2955);
nand U3039 (N_3039,N_2495,N_2561);
and U3040 (N_3040,N_2661,N_2530);
nor U3041 (N_3041,N_2454,N_2702);
xnor U3042 (N_3042,N_2272,N_2973);
nor U3043 (N_3043,N_2764,N_2697);
xnor U3044 (N_3044,N_2626,N_2333);
nand U3045 (N_3045,N_2883,N_2521);
nand U3046 (N_3046,N_2266,N_2528);
and U3047 (N_3047,N_2720,N_2276);
or U3048 (N_3048,N_2406,N_2895);
xnor U3049 (N_3049,N_2419,N_2321);
nor U3050 (N_3050,N_2651,N_2596);
xnor U3051 (N_3051,N_2468,N_2291);
nand U3052 (N_3052,N_2264,N_2640);
and U3053 (N_3053,N_2351,N_2957);
xor U3054 (N_3054,N_2746,N_2387);
or U3055 (N_3055,N_2660,N_2674);
and U3056 (N_3056,N_2362,N_2552);
xnor U3057 (N_3057,N_2280,N_2629);
xnor U3058 (N_3058,N_2896,N_2738);
nand U3059 (N_3059,N_2536,N_2497);
nand U3060 (N_3060,N_2927,N_2318);
or U3061 (N_3061,N_2310,N_2759);
and U3062 (N_3062,N_2818,N_2725);
nand U3063 (N_3063,N_2669,N_2686);
or U3064 (N_3064,N_2486,N_2921);
and U3065 (N_3065,N_2499,N_2960);
xor U3066 (N_3066,N_2672,N_2992);
and U3067 (N_3067,N_2365,N_2556);
or U3068 (N_3068,N_2869,N_2275);
and U3069 (N_3069,N_2446,N_2622);
nand U3070 (N_3070,N_2537,N_2952);
or U3071 (N_3071,N_2460,N_2719);
or U3072 (N_3072,N_2479,N_2645);
and U3073 (N_3073,N_2656,N_2473);
nor U3074 (N_3074,N_2586,N_2964);
nand U3075 (N_3075,N_2331,N_2474);
nand U3076 (N_3076,N_2996,N_2630);
or U3077 (N_3077,N_2694,N_2442);
and U3078 (N_3078,N_2770,N_2966);
xnor U3079 (N_3079,N_2659,N_2308);
nor U3080 (N_3080,N_2529,N_2868);
nand U3081 (N_3081,N_2572,N_2670);
nand U3082 (N_3082,N_2265,N_2511);
xnor U3083 (N_3083,N_2716,N_2598);
nand U3084 (N_3084,N_2544,N_2408);
nand U3085 (N_3085,N_2783,N_2589);
xor U3086 (N_3086,N_2253,N_2425);
nand U3087 (N_3087,N_2443,N_2831);
and U3088 (N_3088,N_2754,N_2843);
or U3089 (N_3089,N_2282,N_2985);
xnor U3090 (N_3090,N_2873,N_2557);
nor U3091 (N_3091,N_2779,N_2588);
and U3092 (N_3092,N_2676,N_2477);
nand U3093 (N_3093,N_2780,N_2830);
nor U3094 (N_3094,N_2889,N_2750);
or U3095 (N_3095,N_2741,N_2677);
or U3096 (N_3096,N_2599,N_2322);
and U3097 (N_3097,N_2734,N_2617);
or U3098 (N_3098,N_2902,N_2890);
or U3099 (N_3099,N_2934,N_2887);
xnor U3100 (N_3100,N_2970,N_2872);
and U3101 (N_3101,N_2317,N_2696);
and U3102 (N_3102,N_2392,N_2802);
and U3103 (N_3103,N_2657,N_2744);
xor U3104 (N_3104,N_2963,N_2724);
nand U3105 (N_3105,N_2583,N_2638);
or U3106 (N_3106,N_2316,N_2405);
or U3107 (N_3107,N_2683,N_2749);
or U3108 (N_3108,N_2948,N_2288);
and U3109 (N_3109,N_2455,N_2628);
or U3110 (N_3110,N_2972,N_2296);
and U3111 (N_3111,N_2593,N_2635);
xor U3112 (N_3112,N_2708,N_2745);
xor U3113 (N_3113,N_2977,N_2366);
xnor U3114 (N_3114,N_2490,N_2760);
or U3115 (N_3115,N_2518,N_2367);
nand U3116 (N_3116,N_2418,N_2678);
nand U3117 (N_3117,N_2608,N_2298);
or U3118 (N_3118,N_2293,N_2397);
nor U3119 (N_3119,N_2937,N_2510);
nor U3120 (N_3120,N_2271,N_2466);
nor U3121 (N_3121,N_2691,N_2345);
nand U3122 (N_3122,N_2368,N_2816);
nand U3123 (N_3123,N_2284,N_2565);
nand U3124 (N_3124,N_2475,N_2546);
nor U3125 (N_3125,N_2515,N_2680);
or U3126 (N_3126,N_2430,N_2603);
nor U3127 (N_3127,N_2978,N_2655);
xor U3128 (N_3128,N_2620,N_2954);
and U3129 (N_3129,N_2824,N_2823);
and U3130 (N_3130,N_2314,N_2534);
xor U3131 (N_3131,N_2261,N_2481);
nor U3132 (N_3132,N_2788,N_2877);
and U3133 (N_3133,N_2447,N_2928);
or U3134 (N_3134,N_2359,N_2496);
xnor U3135 (N_3135,N_2522,N_2395);
xor U3136 (N_3136,N_2326,N_2791);
or U3137 (N_3137,N_2792,N_2273);
and U3138 (N_3138,N_2713,N_2995);
or U3139 (N_3139,N_2402,N_2743);
and U3140 (N_3140,N_2753,N_2449);
nand U3141 (N_3141,N_2832,N_2363);
and U3142 (N_3142,N_2601,N_2639);
and U3143 (N_3143,N_2820,N_2707);
xnor U3144 (N_3144,N_2968,N_2602);
xnor U3145 (N_3145,N_2355,N_2379);
xor U3146 (N_3146,N_2944,N_2946);
or U3147 (N_3147,N_2765,N_2641);
nand U3148 (N_3148,N_2941,N_2612);
and U3149 (N_3149,N_2649,N_2658);
xor U3150 (N_3150,N_2980,N_2803);
and U3151 (N_3151,N_2756,N_2906);
or U3152 (N_3152,N_2413,N_2766);
or U3153 (N_3153,N_2503,N_2856);
nand U3154 (N_3154,N_2698,N_2863);
and U3155 (N_3155,N_2464,N_2942);
or U3156 (N_3156,N_2610,N_2578);
or U3157 (N_3157,N_2739,N_2547);
or U3158 (N_3158,N_2508,N_2457);
or U3159 (N_3159,N_2782,N_2772);
or U3160 (N_3160,N_2582,N_2524);
nor U3161 (N_3161,N_2828,N_2894);
or U3162 (N_3162,N_2730,N_2827);
xnor U3163 (N_3163,N_2354,N_2277);
or U3164 (N_3164,N_2634,N_2684);
nand U3165 (N_3165,N_2568,N_2263);
and U3166 (N_3166,N_2374,N_2722);
nand U3167 (N_3167,N_2900,N_2796);
nor U3168 (N_3168,N_2778,N_2631);
nand U3169 (N_3169,N_2865,N_2252);
or U3170 (N_3170,N_2936,N_2533);
nor U3171 (N_3171,N_2988,N_2673);
or U3172 (N_3172,N_2885,N_2372);
xor U3173 (N_3173,N_2595,N_2251);
or U3174 (N_3174,N_2840,N_2502);
nor U3175 (N_3175,N_2591,N_2685);
or U3176 (N_3176,N_2404,N_2763);
and U3177 (N_3177,N_2543,N_2607);
or U3178 (N_3178,N_2539,N_2880);
and U3179 (N_3179,N_2870,N_2815);
and U3180 (N_3180,N_2859,N_2679);
nand U3181 (N_3181,N_2876,N_2846);
and U3182 (N_3182,N_2422,N_2687);
xor U3183 (N_3183,N_2695,N_2665);
and U3184 (N_3184,N_2693,N_2498);
nor U3185 (N_3185,N_2715,N_2434);
nand U3186 (N_3186,N_2401,N_2429);
nor U3187 (N_3187,N_2648,N_2965);
or U3188 (N_3188,N_2389,N_2548);
and U3189 (N_3189,N_2721,N_2259);
nor U3190 (N_3190,N_2501,N_2836);
and U3191 (N_3191,N_2909,N_2668);
nor U3192 (N_3192,N_2892,N_2535);
and U3193 (N_3193,N_2984,N_2448);
nor U3194 (N_3194,N_2705,N_2424);
and U3195 (N_3195,N_2516,N_2433);
nor U3196 (N_3196,N_2882,N_2975);
nor U3197 (N_3197,N_2338,N_2769);
or U3198 (N_3198,N_2256,N_2845);
nor U3199 (N_3199,N_2855,N_2718);
xnor U3200 (N_3200,N_2295,N_2616);
nand U3201 (N_3201,N_2336,N_2735);
nor U3202 (N_3202,N_2423,N_2623);
nor U3203 (N_3203,N_2647,N_2566);
nand U3204 (N_3204,N_2480,N_2377);
or U3205 (N_3205,N_2723,N_2286);
or U3206 (N_3206,N_2841,N_2627);
xor U3207 (N_3207,N_2594,N_2327);
xnor U3208 (N_3208,N_2709,N_2560);
and U3209 (N_3209,N_2421,N_2580);
nand U3210 (N_3210,N_2577,N_2399);
xnor U3211 (N_3211,N_2728,N_2487);
xor U3212 (N_3212,N_2306,N_2733);
or U3213 (N_3213,N_2382,N_2614);
xnor U3214 (N_3214,N_2357,N_2597);
or U3215 (N_3215,N_2908,N_2671);
nand U3216 (N_3216,N_2943,N_2618);
nand U3217 (N_3217,N_2911,N_2899);
xor U3218 (N_3218,N_2289,N_2315);
and U3219 (N_3219,N_2789,N_2350);
xnor U3220 (N_3220,N_2527,N_2507);
xor U3221 (N_3221,N_2258,N_2550);
nor U3222 (N_3222,N_2904,N_2917);
nand U3223 (N_3223,N_2545,N_2606);
xnor U3224 (N_3224,N_2312,N_2861);
and U3225 (N_3225,N_2349,N_2851);
xor U3226 (N_3226,N_2808,N_2848);
nor U3227 (N_3227,N_2274,N_2767);
or U3228 (N_3228,N_2884,N_2562);
nor U3229 (N_3229,N_2254,N_2787);
and U3230 (N_3230,N_2344,N_2692);
nand U3231 (N_3231,N_2850,N_2532);
nor U3232 (N_3232,N_2866,N_2587);
xnor U3233 (N_3233,N_2689,N_2451);
nor U3234 (N_3234,N_2991,N_2644);
nand U3235 (N_3235,N_2375,N_2431);
xor U3236 (N_3236,N_2436,N_2488);
nor U3237 (N_3237,N_2757,N_2747);
and U3238 (N_3238,N_2555,N_2740);
xor U3239 (N_3239,N_2998,N_2371);
xnor U3240 (N_3240,N_2523,N_2391);
nand U3241 (N_3241,N_2269,N_2699);
and U3242 (N_3242,N_2913,N_2795);
or U3243 (N_3243,N_2912,N_2445);
and U3244 (N_3244,N_2822,N_2444);
nand U3245 (N_3245,N_2775,N_2905);
nor U3246 (N_3246,N_2758,N_2380);
nor U3247 (N_3247,N_2340,N_2483);
nor U3248 (N_3248,N_2852,N_2939);
nor U3249 (N_3249,N_2335,N_2701);
nand U3250 (N_3250,N_2554,N_2667);
xor U3251 (N_3251,N_2898,N_2817);
xor U3252 (N_3252,N_2390,N_2903);
nor U3253 (N_3253,N_2997,N_2294);
or U3254 (N_3254,N_2819,N_2409);
or U3255 (N_3255,N_2862,N_2553);
and U3256 (N_3256,N_2491,N_2774);
nand U3257 (N_3257,N_2492,N_2926);
nand U3258 (N_3258,N_2956,N_2710);
and U3259 (N_3259,N_2918,N_2407);
xnor U3260 (N_3260,N_2297,N_2513);
nor U3261 (N_3261,N_2467,N_2410);
and U3262 (N_3262,N_2804,N_2805);
nor U3263 (N_3263,N_2329,N_2396);
xnor U3264 (N_3264,N_2320,N_2711);
or U3265 (N_3265,N_2959,N_2540);
xor U3266 (N_3266,N_2847,N_2563);
nor U3267 (N_3267,N_2915,N_2812);
and U3268 (N_3268,N_2922,N_2958);
nor U3269 (N_3269,N_2287,N_2325);
nor U3270 (N_3270,N_2737,N_2925);
nor U3271 (N_3271,N_2799,N_2637);
nor U3272 (N_3272,N_2914,N_2874);
or U3273 (N_3273,N_2786,N_2417);
or U3274 (N_3274,N_2923,N_2814);
and U3275 (N_3275,N_2609,N_2910);
and U3276 (N_3276,N_2999,N_2893);
or U3277 (N_3277,N_2319,N_2935);
and U3278 (N_3278,N_2494,N_2776);
nand U3279 (N_3279,N_2646,N_2519);
nor U3280 (N_3280,N_2837,N_2360);
or U3281 (N_3281,N_2590,N_2453);
nand U3282 (N_3282,N_2879,N_2358);
nand U3283 (N_3283,N_2981,N_2813);
xnor U3284 (N_3284,N_2688,N_2463);
xnor U3285 (N_3285,N_2777,N_2761);
nand U3286 (N_3286,N_2706,N_2255);
or U3287 (N_3287,N_2420,N_2654);
and U3288 (N_3288,N_2542,N_2681);
nand U3289 (N_3289,N_2526,N_2334);
nor U3290 (N_3290,N_2929,N_2414);
nand U3291 (N_3291,N_2611,N_2809);
and U3292 (N_3292,N_2307,N_2949);
nor U3293 (N_3293,N_2920,N_2283);
nand U3294 (N_3294,N_2330,N_2569);
nand U3295 (N_3295,N_2452,N_2994);
xnor U3296 (N_3296,N_2858,N_2916);
and U3297 (N_3297,N_2574,N_2439);
nand U3298 (N_3298,N_2621,N_2653);
nand U3299 (N_3299,N_2427,N_2299);
nor U3300 (N_3300,N_2801,N_2472);
nor U3301 (N_3301,N_2538,N_2440);
xor U3302 (N_3302,N_2993,N_2416);
or U3303 (N_3303,N_2373,N_2341);
nor U3304 (N_3304,N_2810,N_2415);
xnor U3305 (N_3305,N_2504,N_2509);
xnor U3306 (N_3306,N_2364,N_2807);
xnor U3307 (N_3307,N_2797,N_2541);
and U3308 (N_3308,N_2332,N_2381);
nand U3309 (N_3309,N_2825,N_2384);
and U3310 (N_3310,N_2302,N_2989);
nor U3311 (N_3311,N_2428,N_2470);
or U3312 (N_3312,N_2505,N_2712);
or U3313 (N_3313,N_2267,N_2833);
nand U3314 (N_3314,N_2967,N_2615);
or U3315 (N_3315,N_2512,N_2986);
nand U3316 (N_3316,N_2931,N_2938);
nor U3317 (N_3317,N_2878,N_2785);
and U3318 (N_3318,N_2969,N_2559);
and U3319 (N_3319,N_2633,N_2592);
and U3320 (N_3320,N_2990,N_2459);
and U3321 (N_3321,N_2309,N_2897);
and U3322 (N_3322,N_2328,N_2412);
or U3323 (N_3323,N_2456,N_2806);
nand U3324 (N_3324,N_2857,N_2987);
nor U3325 (N_3325,N_2773,N_2784);
xnor U3326 (N_3326,N_2982,N_2324);
nor U3327 (N_3327,N_2520,N_2729);
nor U3328 (N_3328,N_2558,N_2393);
nor U3329 (N_3329,N_2727,N_2619);
nor U3330 (N_3330,N_2571,N_2461);
or U3331 (N_3331,N_2953,N_2950);
nand U3332 (N_3332,N_2768,N_2551);
nand U3333 (N_3333,N_2343,N_2636);
nand U3334 (N_3334,N_2755,N_2731);
xor U3335 (N_3335,N_2860,N_2974);
nand U3336 (N_3336,N_2426,N_2871);
or U3337 (N_3337,N_2664,N_2570);
and U3338 (N_3338,N_2793,N_2313);
or U3339 (N_3339,N_2311,N_2613);
and U3340 (N_3340,N_2849,N_2834);
nor U3341 (N_3341,N_2579,N_2301);
and U3342 (N_3342,N_2604,N_2567);
or U3343 (N_3343,N_2983,N_2525);
xnor U3344 (N_3344,N_2506,N_2919);
nor U3345 (N_3345,N_2388,N_2348);
xnor U3346 (N_3346,N_2888,N_2250);
or U3347 (N_3347,N_2650,N_2573);
and U3348 (N_3348,N_2378,N_2835);
nor U3349 (N_3349,N_2370,N_2432);
nand U3350 (N_3350,N_2489,N_2875);
nand U3351 (N_3351,N_2971,N_2762);
nand U3352 (N_3352,N_2385,N_2339);
nor U3353 (N_3353,N_2279,N_2829);
xnor U3354 (N_3354,N_2281,N_2471);
nand U3355 (N_3355,N_2376,N_2901);
or U3356 (N_3356,N_2605,N_2771);
nand U3357 (N_3357,N_2278,N_2581);
xnor U3358 (N_3358,N_2575,N_2305);
nand U3359 (N_3359,N_2867,N_2682);
nand U3360 (N_3360,N_2853,N_2891);
nor U3361 (N_3361,N_2438,N_2465);
nand U3362 (N_3362,N_2794,N_2517);
and U3363 (N_3363,N_2411,N_2790);
and U3364 (N_3364,N_2300,N_2403);
nor U3365 (N_3365,N_2945,N_2469);
xor U3366 (N_3366,N_2398,N_2666);
and U3367 (N_3367,N_2514,N_2976);
or U3368 (N_3368,N_2662,N_2907);
and U3369 (N_3369,N_2632,N_2704);
nand U3370 (N_3370,N_2642,N_2353);
nand U3371 (N_3371,N_2304,N_2356);
and U3372 (N_3372,N_2961,N_2270);
and U3373 (N_3373,N_2458,N_2369);
xnor U3374 (N_3374,N_2732,N_2347);
or U3375 (N_3375,N_2269,N_2737);
xnor U3376 (N_3376,N_2547,N_2535);
and U3377 (N_3377,N_2331,N_2755);
nand U3378 (N_3378,N_2577,N_2954);
or U3379 (N_3379,N_2702,N_2671);
and U3380 (N_3380,N_2677,N_2939);
nand U3381 (N_3381,N_2489,N_2730);
nor U3382 (N_3382,N_2571,N_2322);
and U3383 (N_3383,N_2353,N_2738);
nor U3384 (N_3384,N_2748,N_2833);
xnor U3385 (N_3385,N_2628,N_2684);
nor U3386 (N_3386,N_2732,N_2850);
and U3387 (N_3387,N_2904,N_2657);
nand U3388 (N_3388,N_2371,N_2643);
and U3389 (N_3389,N_2912,N_2466);
nor U3390 (N_3390,N_2837,N_2872);
xor U3391 (N_3391,N_2911,N_2825);
nand U3392 (N_3392,N_2868,N_2306);
and U3393 (N_3393,N_2493,N_2934);
xor U3394 (N_3394,N_2620,N_2791);
nor U3395 (N_3395,N_2498,N_2295);
and U3396 (N_3396,N_2805,N_2852);
xnor U3397 (N_3397,N_2664,N_2766);
or U3398 (N_3398,N_2705,N_2833);
and U3399 (N_3399,N_2951,N_2305);
nor U3400 (N_3400,N_2564,N_2475);
and U3401 (N_3401,N_2646,N_2762);
xnor U3402 (N_3402,N_2255,N_2809);
xor U3403 (N_3403,N_2449,N_2519);
nor U3404 (N_3404,N_2259,N_2941);
or U3405 (N_3405,N_2624,N_2497);
and U3406 (N_3406,N_2515,N_2623);
or U3407 (N_3407,N_2466,N_2806);
or U3408 (N_3408,N_2434,N_2918);
or U3409 (N_3409,N_2404,N_2536);
nand U3410 (N_3410,N_2509,N_2929);
xnor U3411 (N_3411,N_2299,N_2560);
xor U3412 (N_3412,N_2902,N_2470);
nor U3413 (N_3413,N_2831,N_2515);
xor U3414 (N_3414,N_2445,N_2905);
xor U3415 (N_3415,N_2488,N_2949);
or U3416 (N_3416,N_2655,N_2729);
nor U3417 (N_3417,N_2313,N_2288);
xnor U3418 (N_3418,N_2385,N_2986);
nor U3419 (N_3419,N_2496,N_2809);
nor U3420 (N_3420,N_2564,N_2465);
or U3421 (N_3421,N_2546,N_2991);
or U3422 (N_3422,N_2335,N_2391);
and U3423 (N_3423,N_2978,N_2397);
or U3424 (N_3424,N_2399,N_2363);
and U3425 (N_3425,N_2274,N_2443);
nand U3426 (N_3426,N_2742,N_2374);
nor U3427 (N_3427,N_2360,N_2307);
nor U3428 (N_3428,N_2773,N_2441);
nand U3429 (N_3429,N_2933,N_2553);
or U3430 (N_3430,N_2968,N_2437);
or U3431 (N_3431,N_2719,N_2292);
and U3432 (N_3432,N_2985,N_2542);
nand U3433 (N_3433,N_2737,N_2462);
xnor U3434 (N_3434,N_2605,N_2917);
xnor U3435 (N_3435,N_2347,N_2674);
and U3436 (N_3436,N_2468,N_2363);
or U3437 (N_3437,N_2835,N_2349);
xor U3438 (N_3438,N_2579,N_2903);
nand U3439 (N_3439,N_2466,N_2765);
nor U3440 (N_3440,N_2502,N_2309);
nor U3441 (N_3441,N_2687,N_2392);
and U3442 (N_3442,N_2472,N_2716);
nor U3443 (N_3443,N_2442,N_2499);
nand U3444 (N_3444,N_2543,N_2972);
xnor U3445 (N_3445,N_2836,N_2426);
nand U3446 (N_3446,N_2813,N_2585);
xnor U3447 (N_3447,N_2596,N_2919);
nor U3448 (N_3448,N_2840,N_2609);
and U3449 (N_3449,N_2394,N_2752);
and U3450 (N_3450,N_2441,N_2814);
nor U3451 (N_3451,N_2275,N_2627);
and U3452 (N_3452,N_2837,N_2412);
nor U3453 (N_3453,N_2566,N_2774);
nor U3454 (N_3454,N_2583,N_2775);
xor U3455 (N_3455,N_2431,N_2895);
xor U3456 (N_3456,N_2839,N_2716);
or U3457 (N_3457,N_2862,N_2977);
nor U3458 (N_3458,N_2636,N_2973);
or U3459 (N_3459,N_2747,N_2556);
and U3460 (N_3460,N_2678,N_2413);
and U3461 (N_3461,N_2620,N_2413);
xnor U3462 (N_3462,N_2684,N_2811);
or U3463 (N_3463,N_2950,N_2281);
xnor U3464 (N_3464,N_2481,N_2614);
or U3465 (N_3465,N_2561,N_2384);
nand U3466 (N_3466,N_2597,N_2997);
xnor U3467 (N_3467,N_2996,N_2815);
and U3468 (N_3468,N_2792,N_2556);
or U3469 (N_3469,N_2782,N_2460);
nand U3470 (N_3470,N_2579,N_2707);
or U3471 (N_3471,N_2828,N_2588);
and U3472 (N_3472,N_2999,N_2697);
xor U3473 (N_3473,N_2520,N_2413);
and U3474 (N_3474,N_2387,N_2979);
or U3475 (N_3475,N_2911,N_2840);
or U3476 (N_3476,N_2642,N_2985);
xnor U3477 (N_3477,N_2471,N_2351);
nand U3478 (N_3478,N_2475,N_2850);
or U3479 (N_3479,N_2623,N_2782);
nor U3480 (N_3480,N_2748,N_2322);
or U3481 (N_3481,N_2369,N_2702);
or U3482 (N_3482,N_2638,N_2844);
or U3483 (N_3483,N_2699,N_2538);
or U3484 (N_3484,N_2843,N_2305);
xnor U3485 (N_3485,N_2363,N_2853);
or U3486 (N_3486,N_2472,N_2523);
nor U3487 (N_3487,N_2300,N_2738);
xor U3488 (N_3488,N_2683,N_2458);
nand U3489 (N_3489,N_2489,N_2285);
xor U3490 (N_3490,N_2345,N_2533);
and U3491 (N_3491,N_2611,N_2640);
nor U3492 (N_3492,N_2471,N_2298);
or U3493 (N_3493,N_2543,N_2513);
and U3494 (N_3494,N_2782,N_2887);
xor U3495 (N_3495,N_2892,N_2473);
and U3496 (N_3496,N_2482,N_2732);
nor U3497 (N_3497,N_2393,N_2600);
xnor U3498 (N_3498,N_2871,N_2525);
nand U3499 (N_3499,N_2662,N_2575);
nor U3500 (N_3500,N_2799,N_2646);
and U3501 (N_3501,N_2713,N_2864);
nand U3502 (N_3502,N_2501,N_2628);
nor U3503 (N_3503,N_2627,N_2780);
nand U3504 (N_3504,N_2507,N_2846);
or U3505 (N_3505,N_2938,N_2295);
or U3506 (N_3506,N_2408,N_2598);
xnor U3507 (N_3507,N_2456,N_2720);
and U3508 (N_3508,N_2526,N_2400);
or U3509 (N_3509,N_2704,N_2336);
nand U3510 (N_3510,N_2792,N_2839);
xor U3511 (N_3511,N_2707,N_2581);
nand U3512 (N_3512,N_2376,N_2935);
and U3513 (N_3513,N_2272,N_2803);
nand U3514 (N_3514,N_2870,N_2570);
nand U3515 (N_3515,N_2566,N_2630);
or U3516 (N_3516,N_2608,N_2414);
and U3517 (N_3517,N_2491,N_2330);
or U3518 (N_3518,N_2867,N_2317);
nor U3519 (N_3519,N_2594,N_2344);
nor U3520 (N_3520,N_2541,N_2852);
and U3521 (N_3521,N_2798,N_2618);
xnor U3522 (N_3522,N_2735,N_2531);
nand U3523 (N_3523,N_2274,N_2485);
and U3524 (N_3524,N_2293,N_2963);
and U3525 (N_3525,N_2817,N_2657);
nand U3526 (N_3526,N_2687,N_2558);
nand U3527 (N_3527,N_2932,N_2612);
xnor U3528 (N_3528,N_2816,N_2920);
nand U3529 (N_3529,N_2947,N_2508);
nor U3530 (N_3530,N_2972,N_2354);
xnor U3531 (N_3531,N_2615,N_2532);
or U3532 (N_3532,N_2987,N_2585);
and U3533 (N_3533,N_2544,N_2987);
nor U3534 (N_3534,N_2662,N_2648);
nor U3535 (N_3535,N_2337,N_2264);
nand U3536 (N_3536,N_2823,N_2945);
xor U3537 (N_3537,N_2989,N_2379);
nor U3538 (N_3538,N_2546,N_2470);
nor U3539 (N_3539,N_2737,N_2896);
xnor U3540 (N_3540,N_2534,N_2341);
nor U3541 (N_3541,N_2986,N_2586);
nor U3542 (N_3542,N_2501,N_2358);
and U3543 (N_3543,N_2899,N_2693);
nand U3544 (N_3544,N_2590,N_2535);
and U3545 (N_3545,N_2550,N_2397);
and U3546 (N_3546,N_2402,N_2722);
nand U3547 (N_3547,N_2630,N_2987);
nand U3548 (N_3548,N_2867,N_2966);
xnor U3549 (N_3549,N_2436,N_2803);
or U3550 (N_3550,N_2564,N_2677);
nor U3551 (N_3551,N_2612,N_2467);
nor U3552 (N_3552,N_2400,N_2255);
xor U3553 (N_3553,N_2572,N_2869);
or U3554 (N_3554,N_2658,N_2889);
and U3555 (N_3555,N_2924,N_2752);
or U3556 (N_3556,N_2950,N_2289);
xnor U3557 (N_3557,N_2595,N_2493);
nand U3558 (N_3558,N_2815,N_2313);
or U3559 (N_3559,N_2731,N_2644);
and U3560 (N_3560,N_2308,N_2828);
nand U3561 (N_3561,N_2335,N_2742);
nand U3562 (N_3562,N_2714,N_2910);
and U3563 (N_3563,N_2544,N_2565);
xnor U3564 (N_3564,N_2709,N_2727);
nand U3565 (N_3565,N_2693,N_2629);
nand U3566 (N_3566,N_2450,N_2990);
nor U3567 (N_3567,N_2636,N_2392);
xor U3568 (N_3568,N_2684,N_2878);
xnor U3569 (N_3569,N_2687,N_2813);
and U3570 (N_3570,N_2565,N_2609);
nor U3571 (N_3571,N_2425,N_2418);
nor U3572 (N_3572,N_2443,N_2318);
nand U3573 (N_3573,N_2353,N_2469);
nor U3574 (N_3574,N_2499,N_2290);
and U3575 (N_3575,N_2945,N_2583);
xnor U3576 (N_3576,N_2963,N_2898);
nor U3577 (N_3577,N_2616,N_2282);
nand U3578 (N_3578,N_2969,N_2600);
nor U3579 (N_3579,N_2672,N_2836);
or U3580 (N_3580,N_2331,N_2563);
nor U3581 (N_3581,N_2537,N_2795);
nor U3582 (N_3582,N_2341,N_2651);
and U3583 (N_3583,N_2426,N_2648);
xor U3584 (N_3584,N_2975,N_2956);
nor U3585 (N_3585,N_2269,N_2643);
nand U3586 (N_3586,N_2612,N_2444);
nor U3587 (N_3587,N_2402,N_2470);
nor U3588 (N_3588,N_2909,N_2889);
xor U3589 (N_3589,N_2807,N_2887);
nor U3590 (N_3590,N_2304,N_2960);
xnor U3591 (N_3591,N_2526,N_2365);
nand U3592 (N_3592,N_2583,N_2458);
or U3593 (N_3593,N_2256,N_2703);
or U3594 (N_3594,N_2834,N_2437);
nand U3595 (N_3595,N_2428,N_2520);
nand U3596 (N_3596,N_2374,N_2637);
nor U3597 (N_3597,N_2503,N_2665);
or U3598 (N_3598,N_2356,N_2952);
xnor U3599 (N_3599,N_2708,N_2515);
nor U3600 (N_3600,N_2463,N_2438);
nor U3601 (N_3601,N_2491,N_2921);
xnor U3602 (N_3602,N_2777,N_2901);
nor U3603 (N_3603,N_2551,N_2275);
nand U3604 (N_3604,N_2348,N_2682);
and U3605 (N_3605,N_2265,N_2409);
nand U3606 (N_3606,N_2453,N_2991);
xor U3607 (N_3607,N_2385,N_2407);
nand U3608 (N_3608,N_2369,N_2555);
nand U3609 (N_3609,N_2386,N_2275);
nand U3610 (N_3610,N_2955,N_2795);
nor U3611 (N_3611,N_2792,N_2777);
or U3612 (N_3612,N_2896,N_2622);
and U3613 (N_3613,N_2413,N_2460);
and U3614 (N_3614,N_2578,N_2639);
or U3615 (N_3615,N_2424,N_2301);
nor U3616 (N_3616,N_2430,N_2421);
or U3617 (N_3617,N_2343,N_2396);
nor U3618 (N_3618,N_2810,N_2664);
or U3619 (N_3619,N_2337,N_2754);
xnor U3620 (N_3620,N_2503,N_2852);
xnor U3621 (N_3621,N_2712,N_2535);
nor U3622 (N_3622,N_2569,N_2636);
nor U3623 (N_3623,N_2806,N_2779);
xnor U3624 (N_3624,N_2348,N_2804);
and U3625 (N_3625,N_2338,N_2365);
xor U3626 (N_3626,N_2880,N_2578);
xor U3627 (N_3627,N_2353,N_2833);
nor U3628 (N_3628,N_2507,N_2277);
xnor U3629 (N_3629,N_2576,N_2367);
xor U3630 (N_3630,N_2444,N_2436);
nand U3631 (N_3631,N_2445,N_2683);
or U3632 (N_3632,N_2811,N_2979);
or U3633 (N_3633,N_2786,N_2814);
or U3634 (N_3634,N_2320,N_2307);
nor U3635 (N_3635,N_2932,N_2920);
xor U3636 (N_3636,N_2323,N_2828);
xnor U3637 (N_3637,N_2272,N_2282);
xnor U3638 (N_3638,N_2348,N_2874);
xor U3639 (N_3639,N_2347,N_2471);
and U3640 (N_3640,N_2915,N_2859);
and U3641 (N_3641,N_2700,N_2484);
and U3642 (N_3642,N_2499,N_2319);
nor U3643 (N_3643,N_2889,N_2695);
nand U3644 (N_3644,N_2784,N_2663);
or U3645 (N_3645,N_2251,N_2870);
or U3646 (N_3646,N_2624,N_2933);
and U3647 (N_3647,N_2705,N_2744);
nand U3648 (N_3648,N_2704,N_2857);
and U3649 (N_3649,N_2263,N_2781);
nor U3650 (N_3650,N_2953,N_2271);
xor U3651 (N_3651,N_2738,N_2576);
and U3652 (N_3652,N_2709,N_2297);
xnor U3653 (N_3653,N_2397,N_2953);
nand U3654 (N_3654,N_2601,N_2511);
nor U3655 (N_3655,N_2855,N_2781);
or U3656 (N_3656,N_2649,N_2771);
xor U3657 (N_3657,N_2991,N_2601);
and U3658 (N_3658,N_2850,N_2440);
and U3659 (N_3659,N_2365,N_2676);
nand U3660 (N_3660,N_2565,N_2814);
nand U3661 (N_3661,N_2781,N_2499);
or U3662 (N_3662,N_2908,N_2498);
nor U3663 (N_3663,N_2512,N_2582);
nor U3664 (N_3664,N_2648,N_2330);
and U3665 (N_3665,N_2924,N_2730);
xor U3666 (N_3666,N_2740,N_2857);
or U3667 (N_3667,N_2452,N_2792);
nand U3668 (N_3668,N_2775,N_2893);
and U3669 (N_3669,N_2342,N_2289);
or U3670 (N_3670,N_2558,N_2816);
xnor U3671 (N_3671,N_2465,N_2983);
nor U3672 (N_3672,N_2510,N_2922);
and U3673 (N_3673,N_2409,N_2542);
xnor U3674 (N_3674,N_2873,N_2263);
and U3675 (N_3675,N_2307,N_2789);
nor U3676 (N_3676,N_2694,N_2989);
and U3677 (N_3677,N_2408,N_2759);
nand U3678 (N_3678,N_2924,N_2317);
or U3679 (N_3679,N_2955,N_2538);
xnor U3680 (N_3680,N_2822,N_2585);
nor U3681 (N_3681,N_2388,N_2765);
and U3682 (N_3682,N_2784,N_2957);
and U3683 (N_3683,N_2654,N_2744);
nand U3684 (N_3684,N_2835,N_2312);
nand U3685 (N_3685,N_2774,N_2731);
and U3686 (N_3686,N_2775,N_2412);
and U3687 (N_3687,N_2375,N_2589);
nor U3688 (N_3688,N_2355,N_2596);
nor U3689 (N_3689,N_2546,N_2751);
and U3690 (N_3690,N_2268,N_2592);
xnor U3691 (N_3691,N_2682,N_2319);
and U3692 (N_3692,N_2734,N_2842);
nor U3693 (N_3693,N_2385,N_2439);
xor U3694 (N_3694,N_2577,N_2753);
or U3695 (N_3695,N_2362,N_2882);
xnor U3696 (N_3696,N_2390,N_2877);
xor U3697 (N_3697,N_2704,N_2334);
nor U3698 (N_3698,N_2967,N_2748);
nand U3699 (N_3699,N_2999,N_2684);
and U3700 (N_3700,N_2743,N_2540);
xnor U3701 (N_3701,N_2822,N_2929);
nor U3702 (N_3702,N_2870,N_2428);
nand U3703 (N_3703,N_2993,N_2648);
or U3704 (N_3704,N_2984,N_2307);
xnor U3705 (N_3705,N_2898,N_2836);
nand U3706 (N_3706,N_2709,N_2670);
xnor U3707 (N_3707,N_2462,N_2760);
xnor U3708 (N_3708,N_2849,N_2422);
nand U3709 (N_3709,N_2529,N_2335);
xor U3710 (N_3710,N_2581,N_2928);
nand U3711 (N_3711,N_2972,N_2976);
nand U3712 (N_3712,N_2978,N_2795);
xor U3713 (N_3713,N_2448,N_2599);
nand U3714 (N_3714,N_2420,N_2263);
or U3715 (N_3715,N_2621,N_2340);
nor U3716 (N_3716,N_2661,N_2946);
and U3717 (N_3717,N_2762,N_2341);
nor U3718 (N_3718,N_2635,N_2293);
xor U3719 (N_3719,N_2286,N_2796);
xor U3720 (N_3720,N_2771,N_2782);
xor U3721 (N_3721,N_2715,N_2930);
xnor U3722 (N_3722,N_2956,N_2875);
nand U3723 (N_3723,N_2322,N_2450);
nor U3724 (N_3724,N_2761,N_2437);
or U3725 (N_3725,N_2874,N_2588);
nand U3726 (N_3726,N_2278,N_2271);
nor U3727 (N_3727,N_2539,N_2501);
and U3728 (N_3728,N_2966,N_2324);
xnor U3729 (N_3729,N_2650,N_2360);
and U3730 (N_3730,N_2566,N_2805);
xnor U3731 (N_3731,N_2454,N_2850);
and U3732 (N_3732,N_2468,N_2710);
and U3733 (N_3733,N_2800,N_2578);
xor U3734 (N_3734,N_2983,N_2317);
nor U3735 (N_3735,N_2442,N_2916);
nand U3736 (N_3736,N_2328,N_2640);
nor U3737 (N_3737,N_2520,N_2830);
nand U3738 (N_3738,N_2804,N_2571);
nor U3739 (N_3739,N_2783,N_2711);
and U3740 (N_3740,N_2377,N_2552);
and U3741 (N_3741,N_2665,N_2825);
and U3742 (N_3742,N_2745,N_2604);
nor U3743 (N_3743,N_2655,N_2499);
nand U3744 (N_3744,N_2654,N_2762);
nor U3745 (N_3745,N_2921,N_2929);
nor U3746 (N_3746,N_2352,N_2664);
or U3747 (N_3747,N_2443,N_2750);
xor U3748 (N_3748,N_2899,N_2654);
or U3749 (N_3749,N_2938,N_2933);
xor U3750 (N_3750,N_3180,N_3076);
nand U3751 (N_3751,N_3380,N_3018);
or U3752 (N_3752,N_3310,N_3266);
or U3753 (N_3753,N_3295,N_3680);
xor U3754 (N_3754,N_3745,N_3517);
nor U3755 (N_3755,N_3388,N_3248);
nand U3756 (N_3756,N_3640,N_3424);
xor U3757 (N_3757,N_3730,N_3327);
nand U3758 (N_3758,N_3017,N_3510);
nand U3759 (N_3759,N_3151,N_3397);
or U3760 (N_3760,N_3457,N_3613);
and U3761 (N_3761,N_3121,N_3437);
nor U3762 (N_3762,N_3594,N_3707);
nor U3763 (N_3763,N_3672,N_3498);
xor U3764 (N_3764,N_3738,N_3678);
xor U3765 (N_3765,N_3058,N_3372);
nand U3766 (N_3766,N_3186,N_3591);
xnor U3767 (N_3767,N_3556,N_3500);
nand U3768 (N_3768,N_3114,N_3302);
nand U3769 (N_3769,N_3547,N_3393);
or U3770 (N_3770,N_3697,N_3411);
nand U3771 (N_3771,N_3638,N_3196);
xor U3772 (N_3772,N_3321,N_3528);
and U3773 (N_3773,N_3088,N_3491);
nor U3774 (N_3774,N_3013,N_3334);
or U3775 (N_3775,N_3568,N_3176);
or U3776 (N_3776,N_3709,N_3601);
nor U3777 (N_3777,N_3669,N_3376);
or U3778 (N_3778,N_3642,N_3548);
nand U3779 (N_3779,N_3091,N_3209);
and U3780 (N_3780,N_3219,N_3314);
xnor U3781 (N_3781,N_3071,N_3615);
or U3782 (N_3782,N_3499,N_3065);
and U3783 (N_3783,N_3489,N_3352);
and U3784 (N_3784,N_3541,N_3732);
nor U3785 (N_3785,N_3276,N_3513);
nand U3786 (N_3786,N_3394,N_3118);
xnor U3787 (N_3787,N_3259,N_3455);
and U3788 (N_3788,N_3687,N_3663);
xor U3789 (N_3789,N_3264,N_3622);
nor U3790 (N_3790,N_3268,N_3449);
and U3791 (N_3791,N_3152,N_3445);
xnor U3792 (N_3792,N_3520,N_3512);
and U3793 (N_3793,N_3336,N_3433);
nor U3794 (N_3794,N_3718,N_3285);
and U3795 (N_3795,N_3325,N_3049);
nor U3796 (N_3796,N_3181,N_3293);
xor U3797 (N_3797,N_3197,N_3704);
nand U3798 (N_3798,N_3363,N_3626);
xor U3799 (N_3799,N_3679,N_3708);
xor U3800 (N_3800,N_3421,N_3515);
nand U3801 (N_3801,N_3215,N_3565);
and U3802 (N_3802,N_3340,N_3202);
and U3803 (N_3803,N_3208,N_3419);
nor U3804 (N_3804,N_3272,N_3237);
or U3805 (N_3805,N_3214,N_3521);
and U3806 (N_3806,N_3037,N_3170);
nand U3807 (N_3807,N_3353,N_3232);
and U3808 (N_3808,N_3281,N_3641);
or U3809 (N_3809,N_3221,N_3073);
or U3810 (N_3810,N_3684,N_3172);
xor U3811 (N_3811,N_3169,N_3584);
nand U3812 (N_3812,N_3700,N_3081);
nor U3813 (N_3813,N_3090,N_3370);
nor U3814 (N_3814,N_3650,N_3223);
or U3815 (N_3815,N_3705,N_3654);
nand U3816 (N_3816,N_3724,N_3525);
and U3817 (N_3817,N_3486,N_3261);
nor U3818 (N_3818,N_3183,N_3153);
nor U3819 (N_3819,N_3531,N_3624);
and U3820 (N_3820,N_3101,N_3593);
xor U3821 (N_3821,N_3407,N_3140);
xor U3822 (N_3822,N_3304,N_3729);
xnor U3823 (N_3823,N_3092,N_3216);
nor U3824 (N_3824,N_3212,N_3689);
or U3825 (N_3825,N_3280,N_3112);
xor U3826 (N_3826,N_3061,N_3116);
xnor U3827 (N_3827,N_3612,N_3126);
xnor U3828 (N_3828,N_3365,N_3441);
or U3829 (N_3829,N_3720,N_3734);
or U3830 (N_3830,N_3168,N_3006);
nand U3831 (N_3831,N_3296,N_3432);
and U3832 (N_3832,N_3435,N_3623);
xor U3833 (N_3833,N_3303,N_3416);
nand U3834 (N_3834,N_3288,N_3369);
and U3835 (N_3835,N_3198,N_3564);
nand U3836 (N_3836,N_3649,N_3731);
nand U3837 (N_3837,N_3406,N_3374);
nand U3838 (N_3838,N_3082,N_3291);
nor U3839 (N_3839,N_3159,N_3614);
xor U3840 (N_3840,N_3287,N_3021);
nand U3841 (N_3841,N_3269,N_3001);
nand U3842 (N_3842,N_3175,N_3298);
and U3843 (N_3843,N_3238,N_3185);
and U3844 (N_3844,N_3342,N_3326);
and U3845 (N_3845,N_3561,N_3546);
and U3846 (N_3846,N_3355,N_3733);
xor U3847 (N_3847,N_3620,N_3532);
xnor U3848 (N_3848,N_3586,N_3273);
nor U3849 (N_3849,N_3600,N_3358);
or U3850 (N_3850,N_3097,N_3165);
or U3851 (N_3851,N_3211,N_3572);
nor U3852 (N_3852,N_3089,N_3711);
nand U3853 (N_3853,N_3670,N_3201);
or U3854 (N_3854,N_3274,N_3147);
xnor U3855 (N_3855,N_3414,N_3359);
xnor U3856 (N_3856,N_3228,N_3322);
nand U3857 (N_3857,N_3047,N_3244);
xor U3858 (N_3858,N_3659,N_3579);
and U3859 (N_3859,N_3190,N_3119);
or U3860 (N_3860,N_3390,N_3361);
or U3861 (N_3861,N_3467,N_3179);
nand U3862 (N_3862,N_3505,N_3519);
and U3863 (N_3863,N_3706,N_3002);
nor U3864 (N_3864,N_3554,N_3571);
xnor U3865 (N_3865,N_3408,N_3702);
xor U3866 (N_3866,N_3044,N_3712);
nand U3867 (N_3867,N_3124,N_3339);
and U3868 (N_3868,N_3616,N_3052);
nor U3869 (N_3869,N_3748,N_3569);
or U3870 (N_3870,N_3386,N_3282);
and U3871 (N_3871,N_3643,N_3074);
or U3872 (N_3872,N_3206,N_3580);
or U3873 (N_3873,N_3671,N_3028);
nand U3874 (N_3874,N_3027,N_3418);
and U3875 (N_3875,N_3559,N_3462);
or U3876 (N_3876,N_3648,N_3381);
nor U3877 (N_3877,N_3155,N_3451);
xor U3878 (N_3878,N_3736,N_3725);
and U3879 (N_3879,N_3133,N_3200);
nand U3880 (N_3880,N_3127,N_3246);
xor U3881 (N_3881,N_3496,N_3098);
and U3882 (N_3882,N_3283,N_3038);
xor U3883 (N_3883,N_3444,N_3628);
or U3884 (N_3884,N_3573,N_3617);
or U3885 (N_3885,N_3583,N_3239);
and U3886 (N_3886,N_3247,N_3317);
nand U3887 (N_3887,N_3661,N_3301);
xnor U3888 (N_3888,N_3167,N_3135);
and U3889 (N_3889,N_3578,N_3427);
nand U3890 (N_3890,N_3425,N_3651);
nand U3891 (N_3891,N_3292,N_3509);
and U3892 (N_3892,N_3235,N_3335);
or U3893 (N_3893,N_3178,N_3014);
and U3894 (N_3894,N_3514,N_3251);
or U3895 (N_3895,N_3463,N_3193);
and U3896 (N_3896,N_3194,N_3117);
or U3897 (N_3897,N_3694,N_3540);
nand U3898 (N_3898,N_3069,N_3619);
xnor U3899 (N_3899,N_3067,N_3043);
and U3900 (N_3900,N_3157,N_3275);
and U3901 (N_3901,N_3503,N_3122);
nand U3902 (N_3902,N_3577,N_3439);
xor U3903 (N_3903,N_3045,N_3338);
or U3904 (N_3904,N_3551,N_3562);
or U3905 (N_3905,N_3132,N_3453);
nand U3906 (N_3906,N_3046,N_3536);
nor U3907 (N_3907,N_3710,N_3681);
or U3908 (N_3908,N_3364,N_3440);
nand U3909 (N_3909,N_3396,N_3316);
nor U3910 (N_3910,N_3100,N_3438);
and U3911 (N_3911,N_3610,N_3652);
xor U3912 (N_3912,N_3351,N_3692);
xor U3913 (N_3913,N_3078,N_3599);
nand U3914 (N_3914,N_3740,N_3262);
or U3915 (N_3915,N_3534,N_3068);
nand U3916 (N_3916,N_3004,N_3606);
and U3917 (N_3917,N_3000,N_3625);
and U3918 (N_3918,N_3313,N_3328);
nand U3919 (N_3919,N_3420,N_3025);
nand U3920 (N_3920,N_3504,N_3523);
nor U3921 (N_3921,N_3587,N_3156);
nor U3922 (N_3922,N_3057,N_3324);
and U3923 (N_3923,N_3062,N_3323);
nand U3924 (N_3924,N_3252,N_3137);
xnor U3925 (N_3925,N_3744,N_3737);
xnor U3926 (N_3926,N_3241,N_3631);
or U3927 (N_3927,N_3443,N_3297);
nor U3928 (N_3928,N_3431,N_3348);
or U3929 (N_3929,N_3476,N_3596);
nor U3930 (N_3930,N_3686,N_3655);
xor U3931 (N_3931,N_3145,N_3405);
nor U3932 (N_3932,N_3031,N_3229);
nor U3933 (N_3933,N_3401,N_3494);
or U3934 (N_3934,N_3409,N_3426);
nor U3935 (N_3935,N_3570,N_3138);
and U3936 (N_3936,N_3227,N_3522);
and U3937 (N_3937,N_3222,N_3154);
nand U3938 (N_3938,N_3713,N_3721);
and U3939 (N_3939,N_3653,N_3130);
nor U3940 (N_3940,N_3477,N_3039);
nor U3941 (N_3941,N_3646,N_3403);
and U3942 (N_3942,N_3174,N_3389);
xor U3943 (N_3943,N_3309,N_3460);
or U3944 (N_3944,N_3189,N_3267);
or U3945 (N_3945,N_3430,N_3470);
xnor U3946 (N_3946,N_3107,N_3367);
and U3947 (N_3947,N_3487,N_3633);
or U3948 (N_3948,N_3055,N_3345);
nor U3949 (N_3949,N_3258,N_3527);
nor U3950 (N_3950,N_3341,N_3675);
and U3951 (N_3951,N_3123,N_3716);
nand U3952 (N_3952,N_3290,N_3609);
xnor U3953 (N_3953,N_3243,N_3539);
nand U3954 (N_3954,N_3300,N_3464);
xnor U3955 (N_3955,N_3256,N_3093);
and U3956 (N_3956,N_3743,N_3051);
xnor U3957 (N_3957,N_3682,N_3422);
or U3958 (N_3958,N_3299,N_3080);
and U3959 (N_3959,N_3226,N_3289);
xor U3960 (N_3960,N_3668,N_3413);
or U3961 (N_3961,N_3096,N_3493);
and U3962 (N_3962,N_3020,N_3161);
or U3963 (N_3963,N_3630,N_3105);
or U3964 (N_3964,N_3203,N_3371);
xnor U3965 (N_3965,N_3735,N_3749);
nor U3966 (N_3966,N_3319,N_3146);
and U3967 (N_3967,N_3488,N_3010);
xnor U3968 (N_3968,N_3234,N_3306);
nand U3969 (N_3969,N_3662,N_3109);
or U3970 (N_3970,N_3608,N_3332);
and U3971 (N_3971,N_3484,N_3549);
xor U3972 (N_3972,N_3245,N_3184);
and U3973 (N_3973,N_3207,N_3019);
and U3974 (N_3974,N_3485,N_3472);
nor U3975 (N_3975,N_3660,N_3113);
nor U3976 (N_3976,N_3158,N_3452);
xor U3977 (N_3977,N_3727,N_3588);
or U3978 (N_3978,N_3217,N_3473);
xnor U3979 (N_3979,N_3307,N_3347);
and U3980 (N_3980,N_3033,N_3656);
and U3981 (N_3981,N_3085,N_3382);
nor U3982 (N_3982,N_3070,N_3331);
nor U3983 (N_3983,N_3379,N_3602);
xnor U3984 (N_3984,N_3538,N_3150);
and U3985 (N_3985,N_3412,N_3349);
xor U3986 (N_3986,N_3059,N_3305);
or U3987 (N_3987,N_3318,N_3357);
nor U3988 (N_3988,N_3557,N_3746);
or U3989 (N_3989,N_3026,N_3337);
nand U3990 (N_3990,N_3605,N_3698);
nand U3991 (N_3991,N_3213,N_3507);
nand U3992 (N_3992,N_3575,N_3501);
or U3993 (N_3993,N_3526,N_3007);
and U3994 (N_3994,N_3607,N_3343);
or U3995 (N_3995,N_3644,N_3005);
nor U3996 (N_3996,N_3717,N_3048);
nand U3997 (N_3997,N_3257,N_3474);
and U3998 (N_3998,N_3029,N_3436);
nand U3999 (N_3999,N_3447,N_3634);
or U4000 (N_4000,N_3225,N_3254);
and U4001 (N_4001,N_3611,N_3270);
and U4002 (N_4002,N_3576,N_3286);
nor U4003 (N_4003,N_3446,N_3134);
nor U4004 (N_4004,N_3592,N_3567);
or U4005 (N_4005,N_3676,N_3191);
nor U4006 (N_4006,N_3008,N_3518);
nand U4007 (N_4007,N_3516,N_3263);
nor U4008 (N_4008,N_3434,N_3482);
xnor U4009 (N_4009,N_3148,N_3106);
or U4010 (N_4010,N_3461,N_3469);
and U4011 (N_4011,N_3639,N_3036);
and U4012 (N_4012,N_3162,N_3354);
or U4013 (N_4013,N_3308,N_3350);
nand U4014 (N_4014,N_3391,N_3344);
nand U4015 (N_4015,N_3034,N_3277);
or U4016 (N_4016,N_3693,N_3084);
and U4017 (N_4017,N_3204,N_3621);
xnor U4018 (N_4018,N_3603,N_3552);
nor U4019 (N_4019,N_3072,N_3373);
nor U4020 (N_4020,N_3050,N_3714);
or U4021 (N_4021,N_3255,N_3495);
or U4022 (N_4022,N_3465,N_3701);
nor U4023 (N_4023,N_3728,N_3040);
xnor U4024 (N_4024,N_3657,N_3368);
or U4025 (N_4025,N_3558,N_3177);
nand U4026 (N_4026,N_3312,N_3079);
xor U4027 (N_4027,N_3492,N_3233);
and U4028 (N_4028,N_3722,N_3077);
nand U4029 (N_4029,N_3220,N_3094);
or U4030 (N_4030,N_3023,N_3399);
xor U4031 (N_4031,N_3099,N_3129);
xor U4032 (N_4032,N_3497,N_3636);
nand U4033 (N_4033,N_3378,N_3739);
nand U4034 (N_4034,N_3395,N_3468);
xor U4035 (N_4035,N_3141,N_3015);
nand U4036 (N_4036,N_3423,N_3479);
or U4037 (N_4037,N_3673,N_3160);
nor U4038 (N_4038,N_3404,N_3715);
nor U4039 (N_4039,N_3210,N_3511);
or U4040 (N_4040,N_3398,N_3553);
and U4041 (N_4041,N_3171,N_3481);
nor U4042 (N_4042,N_3115,N_3502);
nor U4043 (N_4043,N_3480,N_3083);
nor U4044 (N_4044,N_3530,N_3011);
nand U4045 (N_4045,N_3240,N_3086);
nor U4046 (N_4046,N_3647,N_3265);
nor U4047 (N_4047,N_3585,N_3719);
nand U4048 (N_4048,N_3205,N_3103);
nor U4049 (N_4049,N_3278,N_3544);
and U4050 (N_4050,N_3066,N_3362);
nor U4051 (N_4051,N_3533,N_3450);
and U4052 (N_4052,N_3417,N_3104);
nand U4053 (N_4053,N_3560,N_3110);
nand U4054 (N_4054,N_3555,N_3645);
and U4055 (N_4055,N_3635,N_3236);
and U4056 (N_4056,N_3582,N_3144);
or U4057 (N_4057,N_3022,N_3674);
or U4058 (N_4058,N_3415,N_3375);
xor U4059 (N_4059,N_3111,N_3095);
or U4060 (N_4060,N_3087,N_3448);
or U4061 (N_4061,N_3333,N_3723);
and U4062 (N_4062,N_3429,N_3030);
and U4063 (N_4063,N_3163,N_3629);
nor U4064 (N_4064,N_3218,N_3060);
nand U4065 (N_4065,N_3315,N_3590);
and U4066 (N_4066,N_3566,N_3695);
xor U4067 (N_4067,N_3294,N_3075);
or U4068 (N_4068,N_3542,N_3064);
and U4069 (N_4069,N_3128,N_3677);
or U4070 (N_4070,N_3009,N_3666);
or U4071 (N_4071,N_3042,N_3392);
and U4072 (N_4072,N_3598,N_3199);
or U4073 (N_4073,N_3454,N_3537);
nor U4074 (N_4074,N_3136,N_3524);
and U4075 (N_4075,N_3475,N_3187);
nand U4076 (N_4076,N_3320,N_3279);
nor U4077 (N_4077,N_3550,N_3195);
xor U4078 (N_4078,N_3330,N_3260);
nand U4079 (N_4079,N_3627,N_3231);
nor U4080 (N_4080,N_3574,N_3054);
xor U4081 (N_4081,N_3188,N_3166);
xor U4082 (N_4082,N_3329,N_3597);
xor U4083 (N_4083,N_3637,N_3618);
or U4084 (N_4084,N_3589,N_3685);
xor U4085 (N_4085,N_3683,N_3053);
and U4086 (N_4086,N_3667,N_3466);
and U4087 (N_4087,N_3024,N_3665);
or U4088 (N_4088,N_3699,N_3125);
nand U4089 (N_4089,N_3490,N_3703);
nor U4090 (N_4090,N_3529,N_3164);
xor U4091 (N_4091,N_3563,N_3271);
and U4092 (N_4092,N_3149,N_3506);
nand U4093 (N_4093,N_3032,N_3366);
and U4094 (N_4094,N_3108,N_3632);
xor U4095 (N_4095,N_3224,N_3696);
and U4096 (N_4096,N_3483,N_3192);
or U4097 (N_4097,N_3131,N_3410);
or U4098 (N_4098,N_3041,N_3384);
and U4099 (N_4099,N_3387,N_3690);
and U4100 (N_4100,N_3535,N_3253);
nor U4101 (N_4101,N_3383,N_3726);
nor U4102 (N_4102,N_3471,N_3456);
nand U4103 (N_4103,N_3143,N_3581);
xor U4104 (N_4104,N_3346,N_3139);
xor U4105 (N_4105,N_3142,N_3063);
nor U4106 (N_4106,N_3459,N_3056);
and U4107 (N_4107,N_3400,N_3664);
xor U4108 (N_4108,N_3747,N_3658);
nor U4109 (N_4109,N_3120,N_3356);
nand U4110 (N_4110,N_3102,N_3508);
and U4111 (N_4111,N_3012,N_3545);
nand U4112 (N_4112,N_3230,N_3242);
and U4113 (N_4113,N_3284,N_3003);
nor U4114 (N_4114,N_3688,N_3402);
xnor U4115 (N_4115,N_3385,N_3428);
nand U4116 (N_4116,N_3741,N_3377);
nor U4117 (N_4117,N_3311,N_3360);
or U4118 (N_4118,N_3595,N_3543);
or U4119 (N_4119,N_3458,N_3604);
or U4120 (N_4120,N_3016,N_3182);
nand U4121 (N_4121,N_3742,N_3035);
xor U4122 (N_4122,N_3250,N_3249);
xor U4123 (N_4123,N_3478,N_3442);
nor U4124 (N_4124,N_3691,N_3173);
and U4125 (N_4125,N_3181,N_3034);
and U4126 (N_4126,N_3252,N_3420);
xnor U4127 (N_4127,N_3451,N_3370);
xor U4128 (N_4128,N_3104,N_3467);
xnor U4129 (N_4129,N_3606,N_3286);
xor U4130 (N_4130,N_3468,N_3135);
nand U4131 (N_4131,N_3262,N_3173);
xnor U4132 (N_4132,N_3079,N_3291);
and U4133 (N_4133,N_3079,N_3733);
or U4134 (N_4134,N_3657,N_3004);
and U4135 (N_4135,N_3269,N_3484);
or U4136 (N_4136,N_3372,N_3240);
xor U4137 (N_4137,N_3602,N_3669);
xnor U4138 (N_4138,N_3051,N_3600);
and U4139 (N_4139,N_3547,N_3730);
nand U4140 (N_4140,N_3318,N_3026);
nor U4141 (N_4141,N_3165,N_3561);
xnor U4142 (N_4142,N_3621,N_3033);
nand U4143 (N_4143,N_3395,N_3020);
or U4144 (N_4144,N_3161,N_3600);
xnor U4145 (N_4145,N_3664,N_3396);
xor U4146 (N_4146,N_3148,N_3288);
or U4147 (N_4147,N_3570,N_3582);
or U4148 (N_4148,N_3335,N_3230);
nand U4149 (N_4149,N_3250,N_3639);
or U4150 (N_4150,N_3013,N_3534);
nand U4151 (N_4151,N_3334,N_3017);
or U4152 (N_4152,N_3138,N_3488);
nor U4153 (N_4153,N_3140,N_3059);
nand U4154 (N_4154,N_3556,N_3255);
nand U4155 (N_4155,N_3504,N_3705);
and U4156 (N_4156,N_3045,N_3150);
and U4157 (N_4157,N_3465,N_3124);
xnor U4158 (N_4158,N_3664,N_3445);
and U4159 (N_4159,N_3529,N_3659);
and U4160 (N_4160,N_3608,N_3177);
or U4161 (N_4161,N_3101,N_3199);
nor U4162 (N_4162,N_3493,N_3163);
and U4163 (N_4163,N_3748,N_3580);
or U4164 (N_4164,N_3371,N_3113);
nor U4165 (N_4165,N_3419,N_3282);
or U4166 (N_4166,N_3705,N_3677);
or U4167 (N_4167,N_3049,N_3367);
xor U4168 (N_4168,N_3614,N_3474);
and U4169 (N_4169,N_3200,N_3644);
xnor U4170 (N_4170,N_3671,N_3280);
nand U4171 (N_4171,N_3306,N_3398);
nand U4172 (N_4172,N_3059,N_3330);
and U4173 (N_4173,N_3414,N_3464);
or U4174 (N_4174,N_3438,N_3287);
and U4175 (N_4175,N_3231,N_3157);
or U4176 (N_4176,N_3071,N_3269);
nand U4177 (N_4177,N_3011,N_3325);
and U4178 (N_4178,N_3625,N_3226);
and U4179 (N_4179,N_3215,N_3360);
or U4180 (N_4180,N_3355,N_3559);
or U4181 (N_4181,N_3477,N_3233);
and U4182 (N_4182,N_3708,N_3607);
or U4183 (N_4183,N_3241,N_3466);
nand U4184 (N_4184,N_3280,N_3550);
nor U4185 (N_4185,N_3649,N_3205);
nor U4186 (N_4186,N_3233,N_3730);
nor U4187 (N_4187,N_3540,N_3244);
and U4188 (N_4188,N_3137,N_3535);
or U4189 (N_4189,N_3346,N_3340);
nand U4190 (N_4190,N_3171,N_3299);
nor U4191 (N_4191,N_3353,N_3008);
and U4192 (N_4192,N_3286,N_3505);
xnor U4193 (N_4193,N_3089,N_3325);
and U4194 (N_4194,N_3389,N_3082);
or U4195 (N_4195,N_3256,N_3357);
nand U4196 (N_4196,N_3213,N_3745);
xnor U4197 (N_4197,N_3721,N_3711);
nor U4198 (N_4198,N_3451,N_3716);
nand U4199 (N_4199,N_3705,N_3710);
nand U4200 (N_4200,N_3128,N_3730);
nand U4201 (N_4201,N_3297,N_3435);
or U4202 (N_4202,N_3532,N_3550);
xnor U4203 (N_4203,N_3071,N_3466);
nand U4204 (N_4204,N_3272,N_3243);
nor U4205 (N_4205,N_3126,N_3689);
or U4206 (N_4206,N_3224,N_3346);
nand U4207 (N_4207,N_3544,N_3016);
or U4208 (N_4208,N_3706,N_3207);
nor U4209 (N_4209,N_3398,N_3510);
nor U4210 (N_4210,N_3327,N_3393);
nor U4211 (N_4211,N_3697,N_3189);
or U4212 (N_4212,N_3718,N_3136);
or U4213 (N_4213,N_3445,N_3398);
or U4214 (N_4214,N_3456,N_3002);
xor U4215 (N_4215,N_3538,N_3383);
nor U4216 (N_4216,N_3727,N_3396);
nand U4217 (N_4217,N_3420,N_3284);
nand U4218 (N_4218,N_3183,N_3062);
nor U4219 (N_4219,N_3291,N_3266);
xnor U4220 (N_4220,N_3537,N_3253);
nand U4221 (N_4221,N_3627,N_3008);
xnor U4222 (N_4222,N_3097,N_3275);
nand U4223 (N_4223,N_3315,N_3014);
and U4224 (N_4224,N_3662,N_3631);
nor U4225 (N_4225,N_3468,N_3543);
nor U4226 (N_4226,N_3605,N_3129);
nor U4227 (N_4227,N_3600,N_3240);
nand U4228 (N_4228,N_3047,N_3097);
nor U4229 (N_4229,N_3290,N_3520);
and U4230 (N_4230,N_3613,N_3292);
or U4231 (N_4231,N_3387,N_3369);
or U4232 (N_4232,N_3257,N_3309);
nand U4233 (N_4233,N_3078,N_3668);
or U4234 (N_4234,N_3527,N_3512);
nand U4235 (N_4235,N_3481,N_3705);
xnor U4236 (N_4236,N_3671,N_3305);
nand U4237 (N_4237,N_3470,N_3231);
and U4238 (N_4238,N_3415,N_3102);
or U4239 (N_4239,N_3100,N_3008);
or U4240 (N_4240,N_3560,N_3197);
xor U4241 (N_4241,N_3313,N_3164);
nor U4242 (N_4242,N_3299,N_3501);
or U4243 (N_4243,N_3175,N_3480);
xor U4244 (N_4244,N_3205,N_3468);
xnor U4245 (N_4245,N_3448,N_3327);
or U4246 (N_4246,N_3343,N_3206);
nor U4247 (N_4247,N_3578,N_3603);
xor U4248 (N_4248,N_3237,N_3723);
and U4249 (N_4249,N_3624,N_3146);
or U4250 (N_4250,N_3556,N_3582);
xor U4251 (N_4251,N_3299,N_3069);
xor U4252 (N_4252,N_3056,N_3274);
nor U4253 (N_4253,N_3651,N_3606);
and U4254 (N_4254,N_3416,N_3719);
or U4255 (N_4255,N_3658,N_3651);
nor U4256 (N_4256,N_3295,N_3736);
nand U4257 (N_4257,N_3051,N_3094);
nor U4258 (N_4258,N_3029,N_3618);
and U4259 (N_4259,N_3671,N_3450);
nor U4260 (N_4260,N_3484,N_3276);
and U4261 (N_4261,N_3220,N_3217);
or U4262 (N_4262,N_3282,N_3108);
xor U4263 (N_4263,N_3350,N_3078);
or U4264 (N_4264,N_3549,N_3244);
or U4265 (N_4265,N_3349,N_3592);
and U4266 (N_4266,N_3694,N_3355);
nor U4267 (N_4267,N_3177,N_3683);
nand U4268 (N_4268,N_3163,N_3203);
nor U4269 (N_4269,N_3262,N_3213);
xor U4270 (N_4270,N_3503,N_3590);
or U4271 (N_4271,N_3496,N_3628);
nor U4272 (N_4272,N_3631,N_3669);
nor U4273 (N_4273,N_3478,N_3232);
nand U4274 (N_4274,N_3009,N_3709);
xor U4275 (N_4275,N_3552,N_3547);
and U4276 (N_4276,N_3354,N_3336);
or U4277 (N_4277,N_3181,N_3712);
or U4278 (N_4278,N_3083,N_3516);
xor U4279 (N_4279,N_3203,N_3647);
or U4280 (N_4280,N_3116,N_3076);
or U4281 (N_4281,N_3417,N_3482);
nand U4282 (N_4282,N_3606,N_3326);
nand U4283 (N_4283,N_3276,N_3212);
nand U4284 (N_4284,N_3307,N_3435);
or U4285 (N_4285,N_3187,N_3018);
and U4286 (N_4286,N_3206,N_3498);
xnor U4287 (N_4287,N_3246,N_3710);
nor U4288 (N_4288,N_3112,N_3216);
nor U4289 (N_4289,N_3464,N_3289);
nor U4290 (N_4290,N_3024,N_3646);
and U4291 (N_4291,N_3240,N_3050);
nand U4292 (N_4292,N_3200,N_3265);
xor U4293 (N_4293,N_3033,N_3425);
and U4294 (N_4294,N_3713,N_3362);
nand U4295 (N_4295,N_3687,N_3606);
nor U4296 (N_4296,N_3067,N_3203);
xor U4297 (N_4297,N_3049,N_3096);
or U4298 (N_4298,N_3574,N_3137);
nor U4299 (N_4299,N_3636,N_3491);
nand U4300 (N_4300,N_3665,N_3517);
xnor U4301 (N_4301,N_3198,N_3296);
nor U4302 (N_4302,N_3201,N_3558);
nor U4303 (N_4303,N_3472,N_3745);
nor U4304 (N_4304,N_3471,N_3321);
and U4305 (N_4305,N_3009,N_3169);
nor U4306 (N_4306,N_3245,N_3297);
nand U4307 (N_4307,N_3682,N_3295);
nor U4308 (N_4308,N_3053,N_3337);
and U4309 (N_4309,N_3297,N_3325);
and U4310 (N_4310,N_3558,N_3520);
xor U4311 (N_4311,N_3453,N_3546);
nand U4312 (N_4312,N_3012,N_3214);
nand U4313 (N_4313,N_3204,N_3671);
and U4314 (N_4314,N_3735,N_3746);
nand U4315 (N_4315,N_3580,N_3111);
nor U4316 (N_4316,N_3036,N_3198);
nor U4317 (N_4317,N_3685,N_3304);
and U4318 (N_4318,N_3242,N_3404);
nand U4319 (N_4319,N_3487,N_3677);
and U4320 (N_4320,N_3614,N_3104);
or U4321 (N_4321,N_3679,N_3400);
or U4322 (N_4322,N_3479,N_3281);
nand U4323 (N_4323,N_3230,N_3133);
xnor U4324 (N_4324,N_3175,N_3128);
xor U4325 (N_4325,N_3413,N_3200);
nor U4326 (N_4326,N_3197,N_3523);
xor U4327 (N_4327,N_3084,N_3199);
nor U4328 (N_4328,N_3581,N_3696);
nor U4329 (N_4329,N_3679,N_3472);
nor U4330 (N_4330,N_3599,N_3425);
xnor U4331 (N_4331,N_3493,N_3669);
nor U4332 (N_4332,N_3620,N_3318);
or U4333 (N_4333,N_3505,N_3631);
nor U4334 (N_4334,N_3569,N_3218);
or U4335 (N_4335,N_3623,N_3713);
or U4336 (N_4336,N_3731,N_3008);
xnor U4337 (N_4337,N_3109,N_3539);
xnor U4338 (N_4338,N_3376,N_3005);
xnor U4339 (N_4339,N_3245,N_3270);
nor U4340 (N_4340,N_3689,N_3145);
nor U4341 (N_4341,N_3571,N_3433);
and U4342 (N_4342,N_3091,N_3502);
and U4343 (N_4343,N_3179,N_3495);
nor U4344 (N_4344,N_3745,N_3648);
nand U4345 (N_4345,N_3425,N_3641);
nand U4346 (N_4346,N_3735,N_3048);
or U4347 (N_4347,N_3504,N_3588);
nand U4348 (N_4348,N_3278,N_3468);
xnor U4349 (N_4349,N_3111,N_3259);
nor U4350 (N_4350,N_3519,N_3498);
nor U4351 (N_4351,N_3704,N_3083);
nand U4352 (N_4352,N_3430,N_3438);
or U4353 (N_4353,N_3447,N_3284);
nand U4354 (N_4354,N_3369,N_3144);
xnor U4355 (N_4355,N_3397,N_3465);
nand U4356 (N_4356,N_3469,N_3409);
xnor U4357 (N_4357,N_3526,N_3698);
nor U4358 (N_4358,N_3595,N_3012);
xor U4359 (N_4359,N_3550,N_3498);
nor U4360 (N_4360,N_3309,N_3039);
nor U4361 (N_4361,N_3051,N_3610);
or U4362 (N_4362,N_3715,N_3020);
nand U4363 (N_4363,N_3460,N_3050);
and U4364 (N_4364,N_3733,N_3457);
nor U4365 (N_4365,N_3544,N_3583);
nor U4366 (N_4366,N_3551,N_3628);
or U4367 (N_4367,N_3644,N_3571);
nor U4368 (N_4368,N_3620,N_3116);
xnor U4369 (N_4369,N_3063,N_3195);
nor U4370 (N_4370,N_3244,N_3555);
or U4371 (N_4371,N_3656,N_3024);
nor U4372 (N_4372,N_3354,N_3714);
nor U4373 (N_4373,N_3690,N_3591);
nand U4374 (N_4374,N_3438,N_3588);
and U4375 (N_4375,N_3324,N_3368);
nand U4376 (N_4376,N_3694,N_3596);
xor U4377 (N_4377,N_3181,N_3484);
nor U4378 (N_4378,N_3704,N_3620);
and U4379 (N_4379,N_3560,N_3031);
nor U4380 (N_4380,N_3449,N_3061);
and U4381 (N_4381,N_3211,N_3051);
xor U4382 (N_4382,N_3727,N_3269);
nor U4383 (N_4383,N_3005,N_3229);
or U4384 (N_4384,N_3230,N_3040);
and U4385 (N_4385,N_3706,N_3219);
nand U4386 (N_4386,N_3446,N_3520);
nor U4387 (N_4387,N_3658,N_3660);
or U4388 (N_4388,N_3135,N_3614);
xnor U4389 (N_4389,N_3604,N_3220);
and U4390 (N_4390,N_3264,N_3287);
and U4391 (N_4391,N_3211,N_3651);
and U4392 (N_4392,N_3396,N_3490);
xnor U4393 (N_4393,N_3625,N_3749);
xor U4394 (N_4394,N_3017,N_3165);
nor U4395 (N_4395,N_3072,N_3643);
or U4396 (N_4396,N_3396,N_3214);
xor U4397 (N_4397,N_3483,N_3334);
and U4398 (N_4398,N_3081,N_3207);
nor U4399 (N_4399,N_3682,N_3620);
nand U4400 (N_4400,N_3320,N_3354);
xnor U4401 (N_4401,N_3698,N_3470);
or U4402 (N_4402,N_3196,N_3586);
xnor U4403 (N_4403,N_3296,N_3127);
and U4404 (N_4404,N_3349,N_3037);
and U4405 (N_4405,N_3510,N_3678);
xnor U4406 (N_4406,N_3686,N_3505);
or U4407 (N_4407,N_3747,N_3640);
and U4408 (N_4408,N_3688,N_3324);
or U4409 (N_4409,N_3415,N_3027);
xnor U4410 (N_4410,N_3548,N_3256);
or U4411 (N_4411,N_3606,N_3171);
and U4412 (N_4412,N_3648,N_3308);
or U4413 (N_4413,N_3665,N_3615);
nand U4414 (N_4414,N_3243,N_3121);
xnor U4415 (N_4415,N_3329,N_3675);
xnor U4416 (N_4416,N_3393,N_3740);
or U4417 (N_4417,N_3340,N_3629);
and U4418 (N_4418,N_3350,N_3208);
and U4419 (N_4419,N_3092,N_3018);
and U4420 (N_4420,N_3726,N_3321);
nor U4421 (N_4421,N_3514,N_3551);
nand U4422 (N_4422,N_3072,N_3468);
and U4423 (N_4423,N_3310,N_3219);
nand U4424 (N_4424,N_3119,N_3433);
nor U4425 (N_4425,N_3337,N_3351);
xor U4426 (N_4426,N_3635,N_3207);
nand U4427 (N_4427,N_3590,N_3091);
or U4428 (N_4428,N_3340,N_3694);
or U4429 (N_4429,N_3275,N_3579);
or U4430 (N_4430,N_3697,N_3184);
or U4431 (N_4431,N_3030,N_3489);
or U4432 (N_4432,N_3649,N_3736);
or U4433 (N_4433,N_3403,N_3548);
nand U4434 (N_4434,N_3478,N_3063);
or U4435 (N_4435,N_3404,N_3123);
nand U4436 (N_4436,N_3636,N_3321);
nand U4437 (N_4437,N_3015,N_3338);
or U4438 (N_4438,N_3162,N_3269);
and U4439 (N_4439,N_3522,N_3375);
xor U4440 (N_4440,N_3182,N_3265);
nand U4441 (N_4441,N_3276,N_3057);
or U4442 (N_4442,N_3301,N_3440);
nand U4443 (N_4443,N_3349,N_3552);
and U4444 (N_4444,N_3026,N_3463);
or U4445 (N_4445,N_3018,N_3131);
nor U4446 (N_4446,N_3682,N_3444);
nand U4447 (N_4447,N_3142,N_3161);
xor U4448 (N_4448,N_3177,N_3277);
nand U4449 (N_4449,N_3023,N_3703);
and U4450 (N_4450,N_3698,N_3617);
nor U4451 (N_4451,N_3195,N_3643);
and U4452 (N_4452,N_3328,N_3284);
nand U4453 (N_4453,N_3712,N_3175);
and U4454 (N_4454,N_3320,N_3593);
nor U4455 (N_4455,N_3264,N_3306);
and U4456 (N_4456,N_3719,N_3498);
or U4457 (N_4457,N_3181,N_3522);
xnor U4458 (N_4458,N_3036,N_3356);
or U4459 (N_4459,N_3604,N_3486);
and U4460 (N_4460,N_3705,N_3137);
xnor U4461 (N_4461,N_3363,N_3550);
or U4462 (N_4462,N_3604,N_3039);
nor U4463 (N_4463,N_3219,N_3202);
or U4464 (N_4464,N_3029,N_3399);
or U4465 (N_4465,N_3135,N_3153);
nor U4466 (N_4466,N_3046,N_3053);
xnor U4467 (N_4467,N_3127,N_3420);
xnor U4468 (N_4468,N_3275,N_3241);
or U4469 (N_4469,N_3525,N_3469);
xnor U4470 (N_4470,N_3703,N_3589);
or U4471 (N_4471,N_3501,N_3664);
or U4472 (N_4472,N_3044,N_3735);
xor U4473 (N_4473,N_3650,N_3091);
xnor U4474 (N_4474,N_3581,N_3669);
or U4475 (N_4475,N_3672,N_3151);
or U4476 (N_4476,N_3710,N_3286);
nor U4477 (N_4477,N_3382,N_3548);
nor U4478 (N_4478,N_3216,N_3491);
and U4479 (N_4479,N_3226,N_3420);
nand U4480 (N_4480,N_3410,N_3146);
or U4481 (N_4481,N_3585,N_3703);
xnor U4482 (N_4482,N_3054,N_3247);
nor U4483 (N_4483,N_3651,N_3361);
and U4484 (N_4484,N_3363,N_3607);
xnor U4485 (N_4485,N_3247,N_3160);
and U4486 (N_4486,N_3398,N_3161);
xor U4487 (N_4487,N_3304,N_3202);
and U4488 (N_4488,N_3520,N_3398);
or U4489 (N_4489,N_3176,N_3739);
or U4490 (N_4490,N_3675,N_3547);
nand U4491 (N_4491,N_3336,N_3234);
and U4492 (N_4492,N_3669,N_3658);
or U4493 (N_4493,N_3038,N_3126);
xnor U4494 (N_4494,N_3298,N_3519);
xor U4495 (N_4495,N_3613,N_3141);
xnor U4496 (N_4496,N_3218,N_3669);
nand U4497 (N_4497,N_3353,N_3420);
nand U4498 (N_4498,N_3284,N_3694);
nor U4499 (N_4499,N_3395,N_3359);
nor U4500 (N_4500,N_3933,N_4422);
or U4501 (N_4501,N_4130,N_4420);
or U4502 (N_4502,N_4315,N_4248);
nor U4503 (N_4503,N_3858,N_4151);
or U4504 (N_4504,N_4265,N_4343);
nand U4505 (N_4505,N_3902,N_4192);
nand U4506 (N_4506,N_3810,N_4199);
or U4507 (N_4507,N_4235,N_3940);
nor U4508 (N_4508,N_4414,N_4037);
and U4509 (N_4509,N_4081,N_3977);
or U4510 (N_4510,N_4345,N_4243);
xor U4511 (N_4511,N_4089,N_4026);
xor U4512 (N_4512,N_4217,N_3793);
nand U4513 (N_4513,N_4004,N_4373);
and U4514 (N_4514,N_4189,N_4178);
and U4515 (N_4515,N_4425,N_3838);
and U4516 (N_4516,N_4197,N_4277);
nand U4517 (N_4517,N_3777,N_4423);
xor U4518 (N_4518,N_4119,N_4249);
nor U4519 (N_4519,N_3848,N_3784);
nand U4520 (N_4520,N_4206,N_4124);
and U4521 (N_4521,N_3853,N_4355);
or U4522 (N_4522,N_4335,N_4103);
and U4523 (N_4523,N_3964,N_3898);
nor U4524 (N_4524,N_3942,N_3766);
and U4525 (N_4525,N_4366,N_4498);
nand U4526 (N_4526,N_3854,N_3887);
nor U4527 (N_4527,N_3789,N_4097);
and U4528 (N_4528,N_3871,N_4030);
or U4529 (N_4529,N_3973,N_3862);
and U4530 (N_4530,N_3995,N_4012);
xor U4531 (N_4531,N_3948,N_4136);
xnor U4532 (N_4532,N_4442,N_3791);
or U4533 (N_4533,N_4281,N_4144);
or U4534 (N_4534,N_3957,N_3774);
xor U4535 (N_4535,N_4094,N_3983);
nand U4536 (N_4536,N_4402,N_3767);
or U4537 (N_4537,N_3958,N_4150);
or U4538 (N_4538,N_4287,N_4256);
xor U4539 (N_4539,N_4318,N_4351);
and U4540 (N_4540,N_4399,N_4176);
and U4541 (N_4541,N_3931,N_3753);
nand U4542 (N_4542,N_3929,N_3844);
xnor U4543 (N_4543,N_3779,N_4194);
or U4544 (N_4544,N_4198,N_4040);
and U4545 (N_4545,N_4481,N_4226);
and U4546 (N_4546,N_4053,N_4464);
nand U4547 (N_4547,N_4163,N_3930);
and U4548 (N_4548,N_4262,N_3895);
nand U4549 (N_4549,N_4042,N_4110);
nor U4550 (N_4550,N_4382,N_4025);
xor U4551 (N_4551,N_4024,N_4453);
xor U4552 (N_4552,N_3785,N_4175);
nand U4553 (N_4553,N_4485,N_4329);
or U4554 (N_4554,N_4247,N_3927);
or U4555 (N_4555,N_4046,N_3924);
or U4556 (N_4556,N_4048,N_3832);
xor U4557 (N_4557,N_4061,N_4098);
nand U4558 (N_4558,N_4107,N_4146);
nor U4559 (N_4559,N_4190,N_4203);
or U4560 (N_4560,N_4072,N_3870);
or U4561 (N_4561,N_4236,N_4033);
or U4562 (N_4562,N_3765,N_4191);
xnor U4563 (N_4563,N_4322,N_4029);
nor U4564 (N_4564,N_4079,N_4108);
and U4565 (N_4565,N_3894,N_4237);
and U4566 (N_4566,N_3962,N_4337);
and U4567 (N_4567,N_3943,N_4353);
or U4568 (N_4568,N_3825,N_4044);
or U4569 (N_4569,N_4045,N_4240);
nand U4570 (N_4570,N_4187,N_3761);
and U4571 (N_4571,N_3999,N_4261);
and U4572 (N_4572,N_4439,N_3897);
nor U4573 (N_4573,N_4090,N_4251);
nor U4574 (N_4574,N_3802,N_4415);
nand U4575 (N_4575,N_4100,N_4312);
nand U4576 (N_4576,N_4210,N_3780);
nor U4577 (N_4577,N_4444,N_4465);
nor U4578 (N_4578,N_4070,N_3826);
and U4579 (N_4579,N_3880,N_4474);
nor U4580 (N_4580,N_4458,N_4413);
and U4581 (N_4581,N_4358,N_4067);
nand U4582 (N_4582,N_3807,N_4400);
or U4583 (N_4583,N_4138,N_4409);
and U4584 (N_4584,N_4260,N_4367);
xor U4585 (N_4585,N_4091,N_3952);
and U4586 (N_4586,N_4371,N_3944);
and U4587 (N_4587,N_4306,N_3863);
xor U4588 (N_4588,N_3829,N_4112);
nand U4589 (N_4589,N_3831,N_4158);
or U4590 (N_4590,N_3969,N_4106);
nand U4591 (N_4591,N_4344,N_3959);
nand U4592 (N_4592,N_3903,N_3889);
or U4593 (N_4593,N_4228,N_4011);
and U4594 (N_4594,N_4102,N_4115);
xnor U4595 (N_4595,N_3769,N_4374);
or U4596 (N_4596,N_4380,N_4405);
and U4597 (N_4597,N_3755,N_3875);
nor U4598 (N_4598,N_3915,N_4055);
or U4599 (N_4599,N_3884,N_3941);
xor U4600 (N_4600,N_3905,N_3859);
nand U4601 (N_4601,N_4491,N_3792);
xor U4602 (N_4602,N_3847,N_3781);
nand U4603 (N_4603,N_4200,N_4370);
or U4604 (N_4604,N_4290,N_4139);
nand U4605 (N_4605,N_4336,N_4171);
or U4606 (N_4606,N_4276,N_4041);
nand U4607 (N_4607,N_4239,N_4404);
nand U4608 (N_4608,N_4227,N_4284);
or U4609 (N_4609,N_4417,N_4252);
nand U4610 (N_4610,N_4185,N_4034);
and U4611 (N_4611,N_4216,N_3932);
and U4612 (N_4612,N_4142,N_3773);
xor U4613 (N_4613,N_4093,N_4186);
or U4614 (N_4614,N_4452,N_4148);
xor U4615 (N_4615,N_4495,N_4323);
nor U4616 (N_4616,N_4454,N_4433);
or U4617 (N_4617,N_4401,N_4319);
or U4618 (N_4618,N_4478,N_4294);
nand U4619 (N_4619,N_4273,N_4487);
xor U4620 (N_4620,N_4377,N_4407);
or U4621 (N_4621,N_3770,N_4208);
nor U4622 (N_4622,N_4177,N_4238);
nor U4623 (N_4623,N_4493,N_4320);
xor U4624 (N_4624,N_3809,N_4468);
or U4625 (N_4625,N_4475,N_4170);
and U4626 (N_4626,N_4035,N_4381);
nor U4627 (N_4627,N_4007,N_3975);
nor U4628 (N_4628,N_4376,N_4307);
and U4629 (N_4629,N_3833,N_3771);
nor U4630 (N_4630,N_4255,N_4101);
or U4631 (N_4631,N_3830,N_4328);
and U4632 (N_4632,N_4223,N_3778);
and U4633 (N_4633,N_3996,N_3811);
xnor U4634 (N_4634,N_4435,N_3790);
xnor U4635 (N_4635,N_4310,N_4398);
nand U4636 (N_4636,N_4372,N_4445);
nand U4637 (N_4637,N_4285,N_3994);
or U4638 (N_4638,N_3827,N_4340);
nor U4639 (N_4639,N_3814,N_4071);
and U4640 (N_4640,N_3951,N_4088);
and U4641 (N_4641,N_3945,N_3872);
or U4642 (N_4642,N_3913,N_3794);
xor U4643 (N_4643,N_3968,N_3805);
and U4644 (N_4644,N_4009,N_4326);
and U4645 (N_4645,N_3860,N_4293);
xor U4646 (N_4646,N_4050,N_3804);
nand U4647 (N_4647,N_3786,N_4448);
or U4648 (N_4648,N_4105,N_4135);
xor U4649 (N_4649,N_4424,N_3992);
xnor U4650 (N_4650,N_3934,N_3974);
nand U4651 (N_4651,N_3890,N_4184);
nor U4652 (N_4652,N_3764,N_4164);
nand U4653 (N_4653,N_4008,N_4469);
nand U4654 (N_4654,N_3938,N_4378);
or U4655 (N_4655,N_4379,N_4488);
xnor U4656 (N_4656,N_4418,N_3856);
nand U4657 (N_4657,N_3752,N_4117);
or U4658 (N_4658,N_4292,N_4232);
nor U4659 (N_4659,N_3857,N_4368);
or U4660 (N_4660,N_4393,N_4268);
or U4661 (N_4661,N_4043,N_4038);
nor U4662 (N_4662,N_4122,N_4324);
xnor U4663 (N_4663,N_4313,N_4015);
xor U4664 (N_4664,N_4204,N_3783);
and U4665 (N_4665,N_4411,N_4113);
and U4666 (N_4666,N_3998,N_4394);
nand U4667 (N_4667,N_3882,N_4086);
nand U4668 (N_4668,N_3993,N_3806);
or U4669 (N_4669,N_4395,N_4054);
xnor U4670 (N_4670,N_3828,N_4314);
and U4671 (N_4671,N_4215,N_4327);
xnor U4672 (N_4672,N_4047,N_4220);
nor U4673 (N_4673,N_3982,N_3812);
or U4674 (N_4674,N_3762,N_4157);
nor U4675 (N_4675,N_4257,N_4279);
and U4676 (N_4676,N_3839,N_4169);
xnor U4677 (N_4677,N_4354,N_4118);
or U4678 (N_4678,N_4317,N_4229);
nor U4679 (N_4679,N_4309,N_4278);
nor U4680 (N_4680,N_3985,N_4429);
xor U4681 (N_4681,N_3947,N_3950);
nor U4682 (N_4682,N_3849,N_4111);
and U4683 (N_4683,N_4494,N_4341);
and U4684 (N_4684,N_4068,N_4263);
nand U4685 (N_4685,N_4168,N_4010);
and U4686 (N_4686,N_4365,N_3820);
or U4687 (N_4687,N_4001,N_4470);
xnor U4688 (N_4688,N_4385,N_3817);
or U4689 (N_4689,N_4457,N_3978);
and U4690 (N_4690,N_4451,N_4346);
xor U4691 (N_4691,N_4426,N_4259);
xnor U4692 (N_4692,N_4264,N_4304);
and U4693 (N_4693,N_3936,N_4212);
xor U4694 (N_4694,N_3920,N_4497);
xnor U4695 (N_4695,N_4356,N_4021);
or U4696 (N_4696,N_4123,N_3799);
xnor U4697 (N_4697,N_3991,N_4121);
nor U4698 (N_4698,N_3757,N_4300);
nand U4699 (N_4699,N_3750,N_4408);
nor U4700 (N_4700,N_3795,N_4338);
or U4701 (N_4701,N_4253,N_4137);
nor U4702 (N_4702,N_4149,N_3855);
nor U4703 (N_4703,N_4173,N_3987);
nor U4704 (N_4704,N_3888,N_4431);
and U4705 (N_4705,N_4182,N_4074);
and U4706 (N_4706,N_4258,N_4441);
nand U4707 (N_4707,N_4286,N_3923);
xor U4708 (N_4708,N_4369,N_4443);
and U4709 (N_4709,N_4109,N_3912);
or U4710 (N_4710,N_3949,N_3960);
and U4711 (N_4711,N_3843,N_3989);
xor U4712 (N_4712,N_4126,N_3821);
and U4713 (N_4713,N_4062,N_4480);
and U4714 (N_4714,N_4036,N_4233);
xor U4715 (N_4715,N_3919,N_4181);
or U4716 (N_4716,N_4219,N_3967);
or U4717 (N_4717,N_3892,N_4143);
nor U4718 (N_4718,N_4153,N_3842);
nand U4719 (N_4719,N_3867,N_4213);
nor U4720 (N_4720,N_3914,N_4428);
or U4721 (N_4721,N_3834,N_4436);
nand U4722 (N_4722,N_4162,N_4364);
xor U4723 (N_4723,N_4360,N_4455);
and U4724 (N_4724,N_4282,N_4174);
or U4725 (N_4725,N_4202,N_4056);
nand U4726 (N_4726,N_3921,N_3824);
nor U4727 (N_4727,N_3782,N_4069);
or U4728 (N_4728,N_3758,N_4179);
or U4729 (N_4729,N_4270,N_4195);
nor U4730 (N_4730,N_4450,N_3864);
and U4731 (N_4731,N_3896,N_4078);
xor U4732 (N_4732,N_4254,N_4283);
nor U4733 (N_4733,N_4499,N_4114);
nor U4734 (N_4734,N_3865,N_4154);
xor U4735 (N_4735,N_4473,N_3988);
nand U4736 (N_4736,N_4084,N_4492);
and U4737 (N_4737,N_4039,N_4155);
or U4738 (N_4738,N_4230,N_4180);
xnor U4739 (N_4739,N_3954,N_4348);
nor U4740 (N_4740,N_4161,N_3970);
xor U4741 (N_4741,N_4476,N_3852);
nand U4742 (N_4742,N_4363,N_4057);
nor U4743 (N_4743,N_3851,N_3916);
nor U4744 (N_4744,N_4172,N_4095);
nor U4745 (N_4745,N_3840,N_3917);
nand U4746 (N_4746,N_3891,N_4006);
and U4747 (N_4747,N_4438,N_4332);
and U4748 (N_4748,N_4269,N_3972);
and U4749 (N_4749,N_3937,N_4303);
or U4750 (N_4750,N_4201,N_4390);
xor U4751 (N_4751,N_3986,N_4460);
xnor U4752 (N_4752,N_3953,N_4224);
nor U4753 (N_4753,N_3874,N_4383);
or U4754 (N_4754,N_3751,N_4244);
and U4755 (N_4755,N_3886,N_4387);
or U4756 (N_4756,N_3926,N_4389);
xnor U4757 (N_4757,N_4352,N_3918);
nand U4758 (N_4758,N_4075,N_4274);
and U4759 (N_4759,N_3869,N_4388);
and U4760 (N_4760,N_4267,N_4246);
nand U4761 (N_4761,N_4092,N_4132);
and U4762 (N_4762,N_4116,N_4466);
nand U4763 (N_4763,N_4359,N_4131);
and U4764 (N_4764,N_4082,N_3906);
and U4765 (N_4765,N_4362,N_3881);
nor U4766 (N_4766,N_4479,N_4334);
or U4767 (N_4767,N_3823,N_4017);
nand U4768 (N_4768,N_4005,N_4333);
xor U4769 (N_4769,N_4083,N_3835);
nor U4770 (N_4770,N_4016,N_4166);
nor U4771 (N_4771,N_3979,N_4463);
or U4772 (N_4772,N_4211,N_4221);
nand U4773 (N_4773,N_4266,N_3801);
xor U4774 (N_4774,N_4060,N_4077);
or U4775 (N_4775,N_3797,N_4250);
nand U4776 (N_4776,N_4271,N_4496);
xor U4777 (N_4777,N_3868,N_4298);
nor U4778 (N_4778,N_3883,N_4027);
nand U4779 (N_4779,N_4280,N_3796);
or U4780 (N_4780,N_4301,N_3808);
and U4781 (N_4781,N_4434,N_3873);
nand U4782 (N_4782,N_3798,N_4490);
nand U4783 (N_4783,N_4134,N_3910);
nand U4784 (N_4784,N_4218,N_3966);
xor U4785 (N_4785,N_4140,N_4342);
nor U4786 (N_4786,N_3813,N_4296);
nand U4787 (N_4787,N_4145,N_3815);
and U4788 (N_4788,N_4449,N_3900);
nor U4789 (N_4789,N_4477,N_4416);
or U4790 (N_4790,N_4205,N_4288);
nand U4791 (N_4791,N_3878,N_4063);
xnor U4792 (N_4792,N_4437,N_4347);
or U4793 (N_4793,N_3955,N_3772);
nand U4794 (N_4794,N_4125,N_4207);
xnor U4795 (N_4795,N_4272,N_4225);
nand U4796 (N_4796,N_3935,N_4156);
nand U4797 (N_4797,N_3984,N_3850);
or U4798 (N_4798,N_3946,N_4305);
nand U4799 (N_4799,N_4193,N_4308);
xnor U4800 (N_4800,N_4299,N_3965);
nor U4801 (N_4801,N_4023,N_4003);
and U4802 (N_4802,N_3956,N_4331);
xnor U4803 (N_4803,N_4461,N_4427);
nor U4804 (N_4804,N_4412,N_4440);
or U4805 (N_4805,N_4482,N_4222);
nor U4806 (N_4806,N_4080,N_4421);
xnor U4807 (N_4807,N_4245,N_4013);
nand U4808 (N_4808,N_4316,N_4052);
or U4809 (N_4809,N_4165,N_3841);
and U4810 (N_4810,N_4014,N_4188);
xnor U4811 (N_4811,N_4000,N_4297);
nand U4812 (N_4812,N_3961,N_3763);
or U4813 (N_4813,N_4214,N_4032);
or U4814 (N_4814,N_3909,N_3756);
and U4815 (N_4815,N_3899,N_4391);
or U4816 (N_4816,N_4311,N_4141);
xor U4817 (N_4817,N_3925,N_4325);
or U4818 (N_4818,N_3822,N_4486);
nor U4819 (N_4819,N_3836,N_3788);
xnor U4820 (N_4820,N_4002,N_4241);
nand U4821 (N_4821,N_4489,N_4484);
nor U4822 (N_4822,N_3928,N_3922);
xor U4823 (N_4823,N_4049,N_4096);
nand U4824 (N_4824,N_4321,N_3800);
nor U4825 (N_4825,N_3754,N_4403);
or U4826 (N_4826,N_4058,N_3866);
and U4827 (N_4827,N_3803,N_4330);
xor U4828 (N_4828,N_4059,N_4350);
xor U4829 (N_4829,N_3846,N_4467);
xnor U4830 (N_4830,N_4128,N_4031);
xor U4831 (N_4831,N_4018,N_4483);
or U4832 (N_4832,N_4349,N_4152);
xor U4833 (N_4833,N_3819,N_3976);
or U4834 (N_4834,N_3845,N_4386);
and U4835 (N_4835,N_3861,N_4064);
nand U4836 (N_4836,N_4375,N_4462);
and U4837 (N_4837,N_3990,N_4242);
nor U4838 (N_4838,N_4446,N_4459);
and U4839 (N_4839,N_4087,N_4159);
nand U4840 (N_4840,N_4085,N_3776);
xnor U4841 (N_4841,N_4447,N_4384);
and U4842 (N_4842,N_3904,N_4076);
xnor U4843 (N_4843,N_3885,N_4120);
or U4844 (N_4844,N_4432,N_4302);
and U4845 (N_4845,N_4051,N_4147);
nand U4846 (N_4846,N_4361,N_4456);
and U4847 (N_4847,N_3980,N_4209);
xnor U4848 (N_4848,N_4406,N_3876);
nand U4849 (N_4849,N_3877,N_4339);
nand U4850 (N_4850,N_4073,N_4020);
nand U4851 (N_4851,N_4231,N_4410);
and U4852 (N_4852,N_3907,N_3879);
nand U4853 (N_4853,N_4295,N_4028);
nand U4854 (N_4854,N_4196,N_4167);
and U4855 (N_4855,N_4275,N_3818);
xnor U4856 (N_4856,N_4472,N_4289);
or U4857 (N_4857,N_3963,N_4430);
and U4858 (N_4858,N_3981,N_3939);
nor U4859 (N_4859,N_3997,N_4104);
xor U4860 (N_4860,N_4397,N_3908);
xor U4861 (N_4861,N_4127,N_4065);
nand U4862 (N_4862,N_3775,N_4392);
and U4863 (N_4863,N_4066,N_3837);
or U4864 (N_4864,N_3893,N_4133);
or U4865 (N_4865,N_4129,N_4019);
nand U4866 (N_4866,N_3816,N_4291);
nor U4867 (N_4867,N_4357,N_3787);
or U4868 (N_4868,N_3760,N_4234);
xnor U4869 (N_4869,N_3901,N_4022);
or U4870 (N_4870,N_4396,N_4419);
nand U4871 (N_4871,N_3759,N_4099);
and U4872 (N_4872,N_4471,N_3971);
or U4873 (N_4873,N_3911,N_4183);
xor U4874 (N_4874,N_4160,N_3768);
or U4875 (N_4875,N_4227,N_3912);
nor U4876 (N_4876,N_4340,N_4118);
nand U4877 (N_4877,N_4473,N_4019);
xor U4878 (N_4878,N_3772,N_4357);
nor U4879 (N_4879,N_4449,N_4496);
nand U4880 (N_4880,N_4034,N_3959);
or U4881 (N_4881,N_4229,N_3896);
and U4882 (N_4882,N_4271,N_4165);
nand U4883 (N_4883,N_4365,N_4325);
or U4884 (N_4884,N_3922,N_4021);
or U4885 (N_4885,N_4034,N_4029);
nand U4886 (N_4886,N_4136,N_4417);
xnor U4887 (N_4887,N_3783,N_4030);
nand U4888 (N_4888,N_4336,N_4352);
nand U4889 (N_4889,N_3921,N_4216);
xor U4890 (N_4890,N_4437,N_4088);
or U4891 (N_4891,N_4074,N_4206);
nor U4892 (N_4892,N_3928,N_4488);
or U4893 (N_4893,N_4277,N_4422);
and U4894 (N_4894,N_4484,N_4185);
xor U4895 (N_4895,N_4213,N_3813);
nor U4896 (N_4896,N_3954,N_4363);
and U4897 (N_4897,N_4360,N_4321);
xnor U4898 (N_4898,N_4065,N_3991);
xor U4899 (N_4899,N_4104,N_4456);
xnor U4900 (N_4900,N_4424,N_4479);
or U4901 (N_4901,N_3828,N_4066);
xnor U4902 (N_4902,N_4408,N_4292);
xnor U4903 (N_4903,N_3768,N_4428);
or U4904 (N_4904,N_4273,N_3906);
nor U4905 (N_4905,N_4041,N_3904);
xor U4906 (N_4906,N_3931,N_4356);
and U4907 (N_4907,N_4046,N_3753);
xnor U4908 (N_4908,N_4455,N_4159);
and U4909 (N_4909,N_3996,N_4155);
nand U4910 (N_4910,N_3830,N_4089);
xor U4911 (N_4911,N_4258,N_4197);
or U4912 (N_4912,N_3979,N_3760);
or U4913 (N_4913,N_3819,N_4069);
xor U4914 (N_4914,N_3937,N_3869);
nand U4915 (N_4915,N_4142,N_4446);
nor U4916 (N_4916,N_3759,N_4229);
nor U4917 (N_4917,N_4252,N_4223);
or U4918 (N_4918,N_4272,N_4327);
xnor U4919 (N_4919,N_4062,N_4001);
nor U4920 (N_4920,N_4017,N_4209);
nor U4921 (N_4921,N_4085,N_4459);
or U4922 (N_4922,N_3866,N_4478);
xor U4923 (N_4923,N_4194,N_4391);
and U4924 (N_4924,N_4140,N_4423);
nor U4925 (N_4925,N_3832,N_4220);
nor U4926 (N_4926,N_4366,N_4119);
nor U4927 (N_4927,N_4111,N_3779);
and U4928 (N_4928,N_3751,N_4474);
nand U4929 (N_4929,N_3927,N_4000);
or U4930 (N_4930,N_4107,N_3781);
and U4931 (N_4931,N_3807,N_4087);
nor U4932 (N_4932,N_4048,N_4452);
and U4933 (N_4933,N_4452,N_3945);
or U4934 (N_4934,N_3768,N_3880);
nand U4935 (N_4935,N_4489,N_4260);
or U4936 (N_4936,N_4056,N_4329);
and U4937 (N_4937,N_3850,N_3909);
and U4938 (N_4938,N_4321,N_3984);
nand U4939 (N_4939,N_4267,N_4496);
nand U4940 (N_4940,N_4354,N_3768);
xor U4941 (N_4941,N_3800,N_3997);
or U4942 (N_4942,N_4344,N_3916);
and U4943 (N_4943,N_4035,N_4195);
nor U4944 (N_4944,N_3859,N_4073);
or U4945 (N_4945,N_4103,N_3980);
nor U4946 (N_4946,N_4037,N_3853);
nand U4947 (N_4947,N_4387,N_4051);
nand U4948 (N_4948,N_4478,N_4475);
and U4949 (N_4949,N_4337,N_3848);
nor U4950 (N_4950,N_4088,N_4008);
nand U4951 (N_4951,N_4020,N_4244);
nor U4952 (N_4952,N_3796,N_3773);
xor U4953 (N_4953,N_4098,N_3821);
xnor U4954 (N_4954,N_4103,N_4276);
nor U4955 (N_4955,N_3764,N_3944);
nand U4956 (N_4956,N_3839,N_4322);
nand U4957 (N_4957,N_3761,N_3983);
xnor U4958 (N_4958,N_4134,N_3796);
xor U4959 (N_4959,N_3958,N_4247);
xor U4960 (N_4960,N_3894,N_4041);
and U4961 (N_4961,N_4169,N_4248);
and U4962 (N_4962,N_4197,N_4323);
and U4963 (N_4963,N_4270,N_3871);
nand U4964 (N_4964,N_4054,N_3931);
nand U4965 (N_4965,N_4137,N_4485);
xnor U4966 (N_4966,N_4333,N_4022);
nor U4967 (N_4967,N_3890,N_3985);
or U4968 (N_4968,N_3856,N_4246);
and U4969 (N_4969,N_3821,N_4042);
nor U4970 (N_4970,N_4061,N_4360);
nand U4971 (N_4971,N_4082,N_3775);
nor U4972 (N_4972,N_4482,N_4157);
xnor U4973 (N_4973,N_4206,N_4165);
nor U4974 (N_4974,N_3774,N_3987);
or U4975 (N_4975,N_3966,N_4350);
nand U4976 (N_4976,N_4020,N_4136);
xor U4977 (N_4977,N_4121,N_4134);
and U4978 (N_4978,N_4116,N_4103);
and U4979 (N_4979,N_3758,N_3908);
xnor U4980 (N_4980,N_4198,N_4358);
nand U4981 (N_4981,N_4118,N_4405);
or U4982 (N_4982,N_4174,N_3908);
nand U4983 (N_4983,N_4198,N_4328);
or U4984 (N_4984,N_4162,N_4268);
nand U4985 (N_4985,N_4119,N_4086);
xnor U4986 (N_4986,N_4291,N_3942);
or U4987 (N_4987,N_4062,N_4267);
and U4988 (N_4988,N_4232,N_4137);
and U4989 (N_4989,N_3835,N_3974);
or U4990 (N_4990,N_4322,N_4394);
nand U4991 (N_4991,N_4097,N_4088);
and U4992 (N_4992,N_4036,N_4430);
and U4993 (N_4993,N_4069,N_4135);
nor U4994 (N_4994,N_3796,N_3988);
nand U4995 (N_4995,N_4151,N_4428);
xnor U4996 (N_4996,N_3911,N_3801);
xnor U4997 (N_4997,N_4211,N_4061);
or U4998 (N_4998,N_4055,N_3806);
or U4999 (N_4999,N_3848,N_3889);
xor U5000 (N_5000,N_4487,N_4270);
nand U5001 (N_5001,N_4197,N_4477);
nor U5002 (N_5002,N_4389,N_4394);
xnor U5003 (N_5003,N_4343,N_4407);
nand U5004 (N_5004,N_4357,N_3975);
or U5005 (N_5005,N_4424,N_4209);
and U5006 (N_5006,N_4313,N_3906);
nor U5007 (N_5007,N_4040,N_4046);
nor U5008 (N_5008,N_3783,N_4419);
or U5009 (N_5009,N_4030,N_4458);
nor U5010 (N_5010,N_3779,N_3899);
xnor U5011 (N_5011,N_3811,N_4447);
or U5012 (N_5012,N_3881,N_4273);
nor U5013 (N_5013,N_3864,N_4085);
xnor U5014 (N_5014,N_3773,N_4130);
or U5015 (N_5015,N_3756,N_3760);
xor U5016 (N_5016,N_4376,N_4063);
xor U5017 (N_5017,N_3778,N_4297);
and U5018 (N_5018,N_4138,N_3932);
or U5019 (N_5019,N_4471,N_3988);
and U5020 (N_5020,N_3954,N_4430);
or U5021 (N_5021,N_4446,N_3825);
xnor U5022 (N_5022,N_4068,N_4339);
nor U5023 (N_5023,N_4288,N_4404);
or U5024 (N_5024,N_4245,N_4121);
and U5025 (N_5025,N_4384,N_3853);
xor U5026 (N_5026,N_4110,N_4148);
nor U5027 (N_5027,N_3763,N_4169);
and U5028 (N_5028,N_4327,N_4160);
xnor U5029 (N_5029,N_4357,N_3944);
or U5030 (N_5030,N_3804,N_4176);
nand U5031 (N_5031,N_4245,N_4276);
xor U5032 (N_5032,N_4342,N_3948);
nor U5033 (N_5033,N_4309,N_4259);
nand U5034 (N_5034,N_4032,N_4324);
xnor U5035 (N_5035,N_4110,N_3931);
nand U5036 (N_5036,N_3809,N_4243);
nor U5037 (N_5037,N_4153,N_4358);
xor U5038 (N_5038,N_4168,N_3778);
nand U5039 (N_5039,N_3968,N_4454);
or U5040 (N_5040,N_4116,N_4376);
or U5041 (N_5041,N_4028,N_3900);
xor U5042 (N_5042,N_4191,N_4143);
nand U5043 (N_5043,N_3751,N_3925);
or U5044 (N_5044,N_4000,N_4014);
xor U5045 (N_5045,N_4232,N_4216);
and U5046 (N_5046,N_4243,N_4395);
nor U5047 (N_5047,N_4048,N_3981);
nor U5048 (N_5048,N_3769,N_4237);
xor U5049 (N_5049,N_4199,N_4394);
xnor U5050 (N_5050,N_4096,N_4367);
xnor U5051 (N_5051,N_4338,N_4443);
xnor U5052 (N_5052,N_4242,N_4389);
and U5053 (N_5053,N_3958,N_4489);
nor U5054 (N_5054,N_3848,N_3772);
nand U5055 (N_5055,N_3793,N_4327);
or U5056 (N_5056,N_4217,N_4295);
nor U5057 (N_5057,N_4386,N_3842);
xnor U5058 (N_5058,N_3810,N_4360);
nand U5059 (N_5059,N_4245,N_4168);
xnor U5060 (N_5060,N_3924,N_4207);
and U5061 (N_5061,N_4392,N_4285);
or U5062 (N_5062,N_4071,N_4167);
nor U5063 (N_5063,N_4252,N_4088);
and U5064 (N_5064,N_3974,N_3922);
nor U5065 (N_5065,N_3791,N_3787);
nand U5066 (N_5066,N_3910,N_4284);
and U5067 (N_5067,N_4348,N_4321);
and U5068 (N_5068,N_4419,N_3843);
nor U5069 (N_5069,N_4261,N_4478);
nand U5070 (N_5070,N_4175,N_4360);
nand U5071 (N_5071,N_4180,N_4405);
or U5072 (N_5072,N_4405,N_4309);
xor U5073 (N_5073,N_3880,N_4117);
and U5074 (N_5074,N_3795,N_4188);
and U5075 (N_5075,N_4439,N_4290);
nor U5076 (N_5076,N_3903,N_4281);
or U5077 (N_5077,N_4010,N_4317);
nor U5078 (N_5078,N_3775,N_3902);
and U5079 (N_5079,N_4135,N_4094);
xnor U5080 (N_5080,N_4017,N_3781);
nand U5081 (N_5081,N_4297,N_3925);
and U5082 (N_5082,N_3976,N_4496);
or U5083 (N_5083,N_4180,N_3766);
or U5084 (N_5084,N_3760,N_3975);
nor U5085 (N_5085,N_3892,N_4464);
xnor U5086 (N_5086,N_3914,N_4225);
nand U5087 (N_5087,N_4296,N_4259);
nor U5088 (N_5088,N_4439,N_3765);
xor U5089 (N_5089,N_3824,N_3985);
nand U5090 (N_5090,N_3815,N_3960);
or U5091 (N_5091,N_4442,N_4365);
nand U5092 (N_5092,N_4365,N_3998);
nand U5093 (N_5093,N_3986,N_4184);
nor U5094 (N_5094,N_3772,N_4099);
and U5095 (N_5095,N_3981,N_4299);
nand U5096 (N_5096,N_4096,N_4253);
nand U5097 (N_5097,N_4342,N_4289);
nand U5098 (N_5098,N_3917,N_4245);
xnor U5099 (N_5099,N_3864,N_3968);
nand U5100 (N_5100,N_4416,N_4402);
and U5101 (N_5101,N_3918,N_4232);
and U5102 (N_5102,N_4339,N_3767);
or U5103 (N_5103,N_4329,N_3761);
xnor U5104 (N_5104,N_3949,N_3810);
nor U5105 (N_5105,N_3910,N_4479);
xnor U5106 (N_5106,N_4230,N_4171);
and U5107 (N_5107,N_4311,N_3779);
or U5108 (N_5108,N_4293,N_4436);
or U5109 (N_5109,N_3988,N_3783);
and U5110 (N_5110,N_4009,N_3764);
xor U5111 (N_5111,N_4384,N_4440);
or U5112 (N_5112,N_4236,N_4169);
or U5113 (N_5113,N_4109,N_4004);
nand U5114 (N_5114,N_3862,N_3753);
or U5115 (N_5115,N_3988,N_3835);
nor U5116 (N_5116,N_3922,N_4397);
nor U5117 (N_5117,N_4441,N_4481);
xor U5118 (N_5118,N_4358,N_3970);
or U5119 (N_5119,N_4216,N_3936);
xor U5120 (N_5120,N_3965,N_4293);
or U5121 (N_5121,N_4099,N_4470);
or U5122 (N_5122,N_4212,N_3901);
and U5123 (N_5123,N_4143,N_4036);
and U5124 (N_5124,N_3823,N_4143);
xor U5125 (N_5125,N_3899,N_3940);
xnor U5126 (N_5126,N_4325,N_3936);
nand U5127 (N_5127,N_4101,N_4141);
nand U5128 (N_5128,N_4290,N_4313);
xnor U5129 (N_5129,N_4137,N_4376);
and U5130 (N_5130,N_4094,N_4251);
or U5131 (N_5131,N_4346,N_4397);
or U5132 (N_5132,N_4046,N_4377);
xor U5133 (N_5133,N_3851,N_4025);
nand U5134 (N_5134,N_3776,N_4227);
xnor U5135 (N_5135,N_4328,N_3750);
or U5136 (N_5136,N_4408,N_4307);
xnor U5137 (N_5137,N_3999,N_3875);
and U5138 (N_5138,N_4250,N_4352);
or U5139 (N_5139,N_3772,N_4421);
or U5140 (N_5140,N_4248,N_3994);
and U5141 (N_5141,N_4364,N_4423);
nor U5142 (N_5142,N_4174,N_4488);
nor U5143 (N_5143,N_3949,N_4463);
xor U5144 (N_5144,N_4192,N_4300);
nor U5145 (N_5145,N_4368,N_4215);
and U5146 (N_5146,N_4399,N_4460);
nor U5147 (N_5147,N_4289,N_3839);
or U5148 (N_5148,N_3873,N_3869);
xor U5149 (N_5149,N_4260,N_4145);
and U5150 (N_5150,N_4368,N_4331);
xnor U5151 (N_5151,N_3818,N_3970);
nand U5152 (N_5152,N_3920,N_3800);
nor U5153 (N_5153,N_4292,N_4313);
xor U5154 (N_5154,N_3936,N_4120);
nor U5155 (N_5155,N_4028,N_4096);
nand U5156 (N_5156,N_4401,N_4250);
nor U5157 (N_5157,N_3836,N_4428);
xnor U5158 (N_5158,N_3783,N_4012);
and U5159 (N_5159,N_4113,N_3814);
xnor U5160 (N_5160,N_3865,N_3965);
nand U5161 (N_5161,N_4323,N_4383);
or U5162 (N_5162,N_3976,N_4431);
nand U5163 (N_5163,N_4481,N_3950);
and U5164 (N_5164,N_4327,N_4189);
and U5165 (N_5165,N_3847,N_4327);
nand U5166 (N_5166,N_3886,N_3830);
nor U5167 (N_5167,N_4253,N_4213);
nand U5168 (N_5168,N_4294,N_4137);
or U5169 (N_5169,N_3791,N_3909);
nand U5170 (N_5170,N_4137,N_4194);
xor U5171 (N_5171,N_3918,N_3775);
xnor U5172 (N_5172,N_4438,N_4409);
or U5173 (N_5173,N_3885,N_4069);
or U5174 (N_5174,N_3937,N_4422);
nor U5175 (N_5175,N_4222,N_3917);
nand U5176 (N_5176,N_4160,N_4057);
xor U5177 (N_5177,N_4324,N_4232);
or U5178 (N_5178,N_4152,N_3987);
and U5179 (N_5179,N_4260,N_4302);
and U5180 (N_5180,N_4338,N_4481);
or U5181 (N_5181,N_4305,N_4269);
and U5182 (N_5182,N_4071,N_4304);
nor U5183 (N_5183,N_4420,N_4323);
and U5184 (N_5184,N_4143,N_4328);
nor U5185 (N_5185,N_4315,N_3883);
xor U5186 (N_5186,N_4079,N_3924);
nor U5187 (N_5187,N_3862,N_3996);
or U5188 (N_5188,N_4192,N_4428);
and U5189 (N_5189,N_4430,N_4120);
and U5190 (N_5190,N_4222,N_4309);
or U5191 (N_5191,N_4008,N_4232);
or U5192 (N_5192,N_4490,N_4201);
or U5193 (N_5193,N_4493,N_3762);
xnor U5194 (N_5194,N_3931,N_3976);
and U5195 (N_5195,N_4167,N_3924);
xnor U5196 (N_5196,N_3887,N_4333);
and U5197 (N_5197,N_4356,N_3945);
xor U5198 (N_5198,N_3922,N_4173);
and U5199 (N_5199,N_3817,N_4256);
xor U5200 (N_5200,N_4072,N_4142);
nor U5201 (N_5201,N_4053,N_4143);
nand U5202 (N_5202,N_3868,N_4287);
nor U5203 (N_5203,N_4474,N_4055);
xnor U5204 (N_5204,N_3791,N_3984);
nand U5205 (N_5205,N_4255,N_4108);
nand U5206 (N_5206,N_4156,N_4066);
nor U5207 (N_5207,N_3857,N_4055);
xnor U5208 (N_5208,N_4323,N_4132);
nand U5209 (N_5209,N_4148,N_4095);
and U5210 (N_5210,N_4039,N_4470);
or U5211 (N_5211,N_4058,N_4095);
and U5212 (N_5212,N_3860,N_4365);
nor U5213 (N_5213,N_4499,N_4278);
or U5214 (N_5214,N_3980,N_4176);
or U5215 (N_5215,N_4346,N_3764);
nor U5216 (N_5216,N_4285,N_4192);
and U5217 (N_5217,N_4182,N_3975);
or U5218 (N_5218,N_4499,N_3850);
or U5219 (N_5219,N_3993,N_4285);
nor U5220 (N_5220,N_4207,N_4005);
nor U5221 (N_5221,N_3816,N_3785);
xnor U5222 (N_5222,N_4355,N_3751);
and U5223 (N_5223,N_4269,N_4457);
and U5224 (N_5224,N_4350,N_3775);
and U5225 (N_5225,N_3988,N_4477);
nor U5226 (N_5226,N_4493,N_4112);
nand U5227 (N_5227,N_4246,N_3786);
or U5228 (N_5228,N_4331,N_4056);
and U5229 (N_5229,N_4213,N_4463);
or U5230 (N_5230,N_3759,N_4327);
nand U5231 (N_5231,N_4468,N_4022);
or U5232 (N_5232,N_4399,N_3855);
xnor U5233 (N_5233,N_4392,N_4357);
nand U5234 (N_5234,N_4269,N_4424);
or U5235 (N_5235,N_4054,N_3843);
nand U5236 (N_5236,N_4414,N_3960);
nor U5237 (N_5237,N_4010,N_3880);
and U5238 (N_5238,N_4348,N_4467);
nor U5239 (N_5239,N_3896,N_3865);
nor U5240 (N_5240,N_3795,N_4329);
xnor U5241 (N_5241,N_4101,N_4398);
nand U5242 (N_5242,N_4363,N_3833);
or U5243 (N_5243,N_3917,N_3869);
nor U5244 (N_5244,N_4360,N_3770);
nand U5245 (N_5245,N_4060,N_3752);
and U5246 (N_5246,N_3777,N_4441);
xnor U5247 (N_5247,N_4334,N_3845);
and U5248 (N_5248,N_4231,N_3942);
and U5249 (N_5249,N_4163,N_4031);
or U5250 (N_5250,N_5103,N_4952);
and U5251 (N_5251,N_4985,N_4947);
or U5252 (N_5252,N_4524,N_4971);
nor U5253 (N_5253,N_5055,N_4720);
or U5254 (N_5254,N_4745,N_5040);
or U5255 (N_5255,N_5099,N_5197);
nand U5256 (N_5256,N_4906,N_4702);
nand U5257 (N_5257,N_5125,N_4931);
nand U5258 (N_5258,N_4588,N_4851);
nor U5259 (N_5259,N_5143,N_4757);
and U5260 (N_5260,N_4534,N_4553);
and U5261 (N_5261,N_4867,N_4555);
or U5262 (N_5262,N_4568,N_4894);
nand U5263 (N_5263,N_5079,N_4628);
xnor U5264 (N_5264,N_4937,N_5088);
nand U5265 (N_5265,N_4900,N_4919);
and U5266 (N_5266,N_4823,N_4573);
or U5267 (N_5267,N_4871,N_4543);
or U5268 (N_5268,N_5224,N_5012);
or U5269 (N_5269,N_5043,N_4872);
and U5270 (N_5270,N_4523,N_5131);
nand U5271 (N_5271,N_4596,N_5170);
nor U5272 (N_5272,N_4511,N_5073);
and U5273 (N_5273,N_4846,N_5048);
nor U5274 (N_5274,N_5248,N_4860);
xnor U5275 (N_5275,N_4814,N_4820);
and U5276 (N_5276,N_4782,N_4911);
xor U5277 (N_5277,N_5185,N_4870);
nand U5278 (N_5278,N_4558,N_4815);
and U5279 (N_5279,N_4941,N_4625);
nor U5280 (N_5280,N_5009,N_5148);
nand U5281 (N_5281,N_5041,N_4658);
xor U5282 (N_5282,N_5172,N_4569);
nor U5283 (N_5283,N_5100,N_4994);
xnor U5284 (N_5284,N_4875,N_4806);
nand U5285 (N_5285,N_4661,N_4984);
or U5286 (N_5286,N_4873,N_4791);
nand U5287 (N_5287,N_5188,N_5246);
or U5288 (N_5288,N_5124,N_4956);
and U5289 (N_5289,N_4618,N_4863);
nor U5290 (N_5290,N_4684,N_4903);
nand U5291 (N_5291,N_4611,N_4563);
or U5292 (N_5292,N_5039,N_4804);
and U5293 (N_5293,N_4608,N_4507);
nor U5294 (N_5294,N_4575,N_5011);
and U5295 (N_5295,N_5085,N_4795);
and U5296 (N_5296,N_4794,N_5204);
nand U5297 (N_5297,N_4570,N_4832);
or U5298 (N_5298,N_4803,N_5208);
and U5299 (N_5299,N_4564,N_4807);
or U5300 (N_5300,N_4584,N_5061);
or U5301 (N_5301,N_4622,N_5215);
nand U5302 (N_5302,N_5193,N_5194);
nor U5303 (N_5303,N_4812,N_4682);
nor U5304 (N_5304,N_5093,N_4601);
nand U5305 (N_5305,N_4697,N_4982);
or U5306 (N_5306,N_4891,N_4770);
or U5307 (N_5307,N_4805,N_4515);
nor U5308 (N_5308,N_5161,N_4551);
nand U5309 (N_5309,N_5044,N_5116);
xor U5310 (N_5310,N_4946,N_4710);
nand U5311 (N_5311,N_4735,N_5151);
and U5312 (N_5312,N_4880,N_4530);
or U5313 (N_5313,N_5008,N_5056);
or U5314 (N_5314,N_4707,N_5214);
or U5315 (N_5315,N_4525,N_4856);
and U5316 (N_5316,N_5126,N_5200);
nor U5317 (N_5317,N_4818,N_5095);
xnor U5318 (N_5318,N_5166,N_4904);
xnor U5319 (N_5319,N_4948,N_5175);
and U5320 (N_5320,N_5066,N_4849);
nor U5321 (N_5321,N_4708,N_4582);
and U5322 (N_5322,N_5024,N_4790);
and U5323 (N_5323,N_5062,N_4781);
or U5324 (N_5324,N_4830,N_5105);
xor U5325 (N_5325,N_5106,N_5077);
nor U5326 (N_5326,N_4560,N_5155);
or U5327 (N_5327,N_4606,N_5178);
nor U5328 (N_5328,N_4991,N_4884);
or U5329 (N_5329,N_4506,N_4912);
or U5330 (N_5330,N_4885,N_5081);
xor U5331 (N_5331,N_4689,N_4562);
and U5332 (N_5332,N_5157,N_5144);
nand U5333 (N_5333,N_4843,N_4918);
xnor U5334 (N_5334,N_5243,N_5137);
nor U5335 (N_5335,N_4852,N_4504);
and U5336 (N_5336,N_4855,N_5226);
and U5337 (N_5337,N_4580,N_4597);
and U5338 (N_5338,N_4537,N_4974);
and U5339 (N_5339,N_5003,N_4896);
and U5340 (N_5340,N_4652,N_4769);
xor U5341 (N_5341,N_4718,N_5084);
or U5342 (N_5342,N_5018,N_4716);
xnor U5343 (N_5343,N_4839,N_4943);
xor U5344 (N_5344,N_4999,N_5059);
or U5345 (N_5345,N_4890,N_4737);
xnor U5346 (N_5346,N_4747,N_4698);
nand U5347 (N_5347,N_5113,N_4888);
nand U5348 (N_5348,N_4759,N_4993);
and U5349 (N_5349,N_4917,N_4785);
xor U5350 (N_5350,N_4895,N_4767);
xnor U5351 (N_5351,N_4811,N_4674);
xnor U5352 (N_5352,N_4522,N_5069);
nand U5353 (N_5353,N_4734,N_4930);
and U5354 (N_5354,N_5191,N_4922);
or U5355 (N_5355,N_4679,N_4741);
xnor U5356 (N_5356,N_4983,N_4585);
xnor U5357 (N_5357,N_4714,N_4605);
or U5358 (N_5358,N_5181,N_5201);
nor U5359 (N_5359,N_4541,N_4826);
nor U5360 (N_5360,N_5187,N_4756);
or U5361 (N_5361,N_4742,N_5104);
xnor U5362 (N_5362,N_5049,N_4838);
or U5363 (N_5363,N_4627,N_5046);
or U5364 (N_5364,N_4824,N_4579);
nor U5365 (N_5365,N_4772,N_4744);
nand U5366 (N_5366,N_4669,N_5127);
xor U5367 (N_5367,N_4594,N_5112);
nor U5368 (N_5368,N_4547,N_4681);
nand U5369 (N_5369,N_5004,N_4548);
or U5370 (N_5370,N_5064,N_4591);
and U5371 (N_5371,N_4763,N_4552);
nand U5372 (N_5372,N_4603,N_5117);
xnor U5373 (N_5373,N_5230,N_5177);
nor U5374 (N_5374,N_5021,N_4528);
xnor U5375 (N_5375,N_5228,N_4510);
or U5376 (N_5376,N_4639,N_4914);
nand U5377 (N_5377,N_5219,N_4925);
nand U5378 (N_5378,N_5130,N_4612);
nor U5379 (N_5379,N_5220,N_5247);
or U5380 (N_5380,N_4527,N_4899);
nor U5381 (N_5381,N_4644,N_4960);
nand U5382 (N_5382,N_4724,N_5183);
or U5383 (N_5383,N_4561,N_5235);
and U5384 (N_5384,N_4683,N_5216);
xnor U5385 (N_5385,N_4544,N_5240);
nor U5386 (N_5386,N_4926,N_5168);
or U5387 (N_5387,N_4972,N_4513);
nor U5388 (N_5388,N_4953,N_4670);
and U5389 (N_5389,N_4802,N_4559);
and U5390 (N_5390,N_4779,N_5067);
nand U5391 (N_5391,N_4538,N_4809);
nand U5392 (N_5392,N_5122,N_4910);
or U5393 (N_5393,N_5160,N_4761);
nand U5394 (N_5394,N_4746,N_4633);
nor U5395 (N_5395,N_5023,N_5233);
and U5396 (N_5396,N_5006,N_5107);
and U5397 (N_5397,N_5232,N_4648);
nor U5398 (N_5398,N_4987,N_4672);
xor U5399 (N_5399,N_4593,N_5225);
and U5400 (N_5400,N_4813,N_5020);
and U5401 (N_5401,N_4576,N_5182);
nor U5402 (N_5402,N_5002,N_4651);
xor U5403 (N_5403,N_4663,N_5237);
nor U5404 (N_5404,N_4728,N_5190);
nand U5405 (N_5405,N_4637,N_4620);
and U5406 (N_5406,N_4965,N_4955);
xnor U5407 (N_5407,N_4920,N_4869);
and U5408 (N_5408,N_4566,N_5153);
nand U5409 (N_5409,N_4825,N_5118);
nand U5410 (N_5410,N_5196,N_4934);
xnor U5411 (N_5411,N_5054,N_4655);
xor U5412 (N_5412,N_5179,N_4610);
and U5413 (N_5413,N_4600,N_5090);
nand U5414 (N_5414,N_5038,N_4961);
nor U5415 (N_5415,N_4771,N_4615);
nor U5416 (N_5416,N_5205,N_5025);
nor U5417 (N_5417,N_4862,N_4653);
and U5418 (N_5418,N_5019,N_4951);
or U5419 (N_5419,N_5078,N_4879);
nor U5420 (N_5420,N_5029,N_4660);
and U5421 (N_5421,N_4709,N_4789);
nor U5422 (N_5422,N_4516,N_4508);
xor U5423 (N_5423,N_5030,N_4755);
and U5424 (N_5424,N_4532,N_4845);
xnor U5425 (N_5425,N_4536,N_4963);
and U5426 (N_5426,N_5022,N_5229);
xnor U5427 (N_5427,N_5097,N_4859);
nor U5428 (N_5428,N_5089,N_4602);
xnor U5429 (N_5429,N_4662,N_5010);
and U5430 (N_5430,N_4822,N_4666);
and U5431 (N_5431,N_5086,N_4954);
nand U5432 (N_5432,N_4529,N_4964);
nand U5433 (N_5433,N_5026,N_4887);
or U5434 (N_5434,N_5005,N_4969);
and U5435 (N_5435,N_4857,N_4801);
nor U5436 (N_5436,N_4793,N_5108);
xnor U5437 (N_5437,N_5050,N_4743);
nand U5438 (N_5438,N_5211,N_4768);
nand U5439 (N_5439,N_4630,N_4977);
and U5440 (N_5440,N_5028,N_5109);
nor U5441 (N_5441,N_5147,N_4694);
nand U5442 (N_5442,N_4695,N_4753);
and U5443 (N_5443,N_5245,N_4642);
xnor U5444 (N_5444,N_5110,N_4667);
or U5445 (N_5445,N_4866,N_4719);
nand U5446 (N_5446,N_4700,N_4533);
xor U5447 (N_5447,N_4916,N_4928);
and U5448 (N_5448,N_5244,N_5132);
nand U5449 (N_5449,N_5167,N_4998);
xnor U5450 (N_5450,N_5159,N_4908);
nand U5451 (N_5451,N_4675,N_5027);
nand U5452 (N_5452,N_4861,N_5034);
xor U5453 (N_5453,N_5149,N_4936);
nor U5454 (N_5454,N_5176,N_4898);
nor U5455 (N_5455,N_5037,N_4545);
nor U5456 (N_5456,N_5072,N_5134);
nand U5457 (N_5457,N_5063,N_4780);
or U5458 (N_5458,N_4577,N_4995);
nor U5459 (N_5459,N_4976,N_4848);
xor U5460 (N_5460,N_4877,N_4712);
xnor U5461 (N_5461,N_4819,N_5000);
xnor U5462 (N_5462,N_4574,N_5053);
xor U5463 (N_5463,N_5007,N_4876);
xnor U5464 (N_5464,N_4927,N_5140);
xor U5465 (N_5465,N_4766,N_4565);
nand U5466 (N_5466,N_4854,N_4640);
nor U5467 (N_5467,N_4874,N_4722);
and U5468 (N_5468,N_4760,N_5206);
and U5469 (N_5469,N_5111,N_5202);
and U5470 (N_5470,N_4514,N_4500);
nand U5471 (N_5471,N_5171,N_4711);
nand U5472 (N_5472,N_5123,N_5222);
or U5473 (N_5473,N_4783,N_4986);
nor U5474 (N_5474,N_4990,N_4645);
nor U5475 (N_5475,N_4542,N_4988);
and U5476 (N_5476,N_5133,N_4557);
and U5477 (N_5477,N_4502,N_4554);
nand U5478 (N_5478,N_4732,N_4629);
and U5479 (N_5479,N_4787,N_5032);
or U5480 (N_5480,N_4656,N_4773);
or U5481 (N_5481,N_5249,N_5114);
and U5482 (N_5482,N_4721,N_5075);
nand U5483 (N_5483,N_5065,N_5051);
and U5484 (N_5484,N_4828,N_5236);
or U5485 (N_5485,N_5074,N_4730);
and U5486 (N_5486,N_5164,N_4808);
nand U5487 (N_5487,N_4583,N_5238);
or U5488 (N_5488,N_5223,N_4680);
xor U5489 (N_5489,N_4868,N_4967);
nor U5490 (N_5490,N_4671,N_5057);
xor U5491 (N_5491,N_4798,N_4751);
or U5492 (N_5492,N_4665,N_5087);
nor U5493 (N_5493,N_5145,N_5115);
and U5494 (N_5494,N_4571,N_4973);
xor U5495 (N_5495,N_5121,N_4733);
or U5496 (N_5496,N_5068,N_4792);
nor U5497 (N_5497,N_5083,N_5239);
and U5498 (N_5498,N_4691,N_5080);
and U5499 (N_5499,N_5082,N_5154);
xnor U5500 (N_5500,N_5227,N_5203);
or U5501 (N_5501,N_5158,N_4831);
xor U5502 (N_5502,N_4587,N_5128);
nand U5503 (N_5503,N_4617,N_4784);
nor U5504 (N_5504,N_5234,N_4817);
or U5505 (N_5505,N_4750,N_4979);
nand U5506 (N_5506,N_4677,N_5016);
and U5507 (N_5507,N_5071,N_4858);
and U5508 (N_5508,N_4723,N_4847);
nand U5509 (N_5509,N_4567,N_4821);
or U5510 (N_5510,N_4643,N_4520);
nor U5511 (N_5511,N_4609,N_4889);
and U5512 (N_5512,N_5060,N_5180);
or U5513 (N_5513,N_4749,N_4764);
nand U5514 (N_5514,N_5186,N_4727);
xor U5515 (N_5515,N_5045,N_4886);
and U5516 (N_5516,N_5094,N_4589);
or U5517 (N_5517,N_5241,N_4631);
and U5518 (N_5518,N_4853,N_4923);
and U5519 (N_5519,N_4657,N_4717);
xnor U5520 (N_5520,N_4646,N_5218);
nand U5521 (N_5521,N_4512,N_4850);
or U5522 (N_5522,N_4586,N_4765);
or U5523 (N_5523,N_5119,N_5096);
nand U5524 (N_5524,N_5173,N_4678);
nor U5525 (N_5525,N_4844,N_5169);
and U5526 (N_5526,N_4797,N_4882);
or U5527 (N_5527,N_4736,N_5212);
nand U5528 (N_5528,N_5142,N_4800);
and U5529 (N_5529,N_4624,N_4932);
or U5530 (N_5530,N_4676,N_5138);
nor U5531 (N_5531,N_4842,N_4739);
and U5532 (N_5532,N_5102,N_4539);
or U5533 (N_5533,N_5209,N_4726);
and U5534 (N_5534,N_5184,N_4957);
nor U5535 (N_5535,N_4688,N_4929);
or U5536 (N_5536,N_4833,N_5129);
and U5537 (N_5537,N_4690,N_5101);
nor U5538 (N_5538,N_4942,N_4595);
nand U5539 (N_5539,N_4664,N_5242);
xnor U5540 (N_5540,N_4958,N_5031);
nor U5541 (N_5541,N_4635,N_5058);
or U5542 (N_5542,N_4944,N_5052);
nand U5543 (N_5543,N_4864,N_5013);
nor U5544 (N_5544,N_4686,N_4962);
xor U5545 (N_5545,N_4775,N_4693);
nand U5546 (N_5546,N_4827,N_4614);
nor U5547 (N_5547,N_4550,N_5070);
or U5548 (N_5548,N_4715,N_5047);
nand U5549 (N_5549,N_4668,N_4786);
xor U5550 (N_5550,N_4924,N_4578);
or U5551 (N_5551,N_5152,N_4796);
or U5552 (N_5552,N_4997,N_5198);
nand U5553 (N_5553,N_4503,N_4501);
or U5554 (N_5554,N_4754,N_4572);
or U5555 (N_5555,N_4518,N_4685);
nand U5556 (N_5556,N_4829,N_4913);
and U5557 (N_5557,N_4978,N_5139);
nand U5558 (N_5558,N_5042,N_4613);
nor U5559 (N_5559,N_4907,N_4654);
and U5560 (N_5560,N_5221,N_4725);
nand U5561 (N_5561,N_4788,N_4604);
or U5562 (N_5562,N_5035,N_5120);
or U5563 (N_5563,N_5150,N_5091);
xnor U5564 (N_5564,N_5146,N_4531);
nor U5565 (N_5565,N_4881,N_4989);
nor U5566 (N_5566,N_4902,N_4526);
xor U5567 (N_5567,N_4626,N_4598);
nor U5568 (N_5568,N_4883,N_5192);
or U5569 (N_5569,N_4647,N_4621);
nand U5570 (N_5570,N_5189,N_4938);
or U5571 (N_5571,N_4703,N_4901);
or U5572 (N_5572,N_5199,N_4673);
nor U5573 (N_5573,N_4619,N_4540);
nand U5574 (N_5574,N_4992,N_4752);
nand U5575 (N_5575,N_4940,N_4696);
and U5576 (N_5576,N_4649,N_4581);
nor U5577 (N_5577,N_4701,N_4777);
and U5578 (N_5578,N_4748,N_4840);
nor U5579 (N_5579,N_4950,N_5136);
or U5580 (N_5580,N_4740,N_4549);
or U5581 (N_5581,N_4841,N_4933);
or U5582 (N_5582,N_4634,N_4758);
nor U5583 (N_5583,N_4632,N_4865);
and U5584 (N_5584,N_4909,N_5165);
nand U5585 (N_5585,N_5036,N_4935);
and U5586 (N_5586,N_4546,N_4836);
and U5587 (N_5587,N_5098,N_4692);
xnor U5588 (N_5588,N_4893,N_5033);
and U5589 (N_5589,N_5076,N_4650);
xnor U5590 (N_5590,N_4731,N_4945);
nand U5591 (N_5591,N_4704,N_4713);
xnor U5592 (N_5592,N_4970,N_4980);
nand U5593 (N_5593,N_5001,N_5014);
and U5594 (N_5594,N_4519,N_4975);
and U5595 (N_5595,N_4517,N_5174);
and U5596 (N_5596,N_4949,N_4959);
nand U5597 (N_5597,N_5141,N_4592);
xnor U5598 (N_5598,N_4778,N_4623);
nor U5599 (N_5599,N_4687,N_4607);
nor U5600 (N_5600,N_5162,N_4599);
or U5601 (N_5601,N_4521,N_4799);
xnor U5602 (N_5602,N_4638,N_4636);
xnor U5603 (N_5603,N_5195,N_4966);
or U5604 (N_5604,N_4939,N_4705);
and U5605 (N_5605,N_4837,N_4996);
xor U5606 (N_5606,N_5017,N_5207);
nand U5607 (N_5607,N_5217,N_4762);
nand U5608 (N_5608,N_4905,N_4738);
or U5609 (N_5609,N_4706,N_4897);
or U5610 (N_5610,N_4659,N_4968);
nand U5611 (N_5611,N_4878,N_4816);
nand U5612 (N_5612,N_4981,N_5210);
nand U5613 (N_5613,N_4505,N_4915);
xor U5614 (N_5614,N_4509,N_4535);
or U5615 (N_5615,N_4810,N_5231);
or U5616 (N_5616,N_4834,N_4921);
nor U5617 (N_5617,N_5015,N_5092);
nand U5618 (N_5618,N_4729,N_4616);
or U5619 (N_5619,N_4556,N_4835);
xnor U5620 (N_5620,N_4641,N_5213);
and U5621 (N_5621,N_4776,N_4892);
or U5622 (N_5622,N_5135,N_4774);
xnor U5623 (N_5623,N_4699,N_5163);
and U5624 (N_5624,N_5156,N_4590);
nor U5625 (N_5625,N_5181,N_4736);
xor U5626 (N_5626,N_4933,N_4778);
nor U5627 (N_5627,N_4755,N_5160);
nor U5628 (N_5628,N_4648,N_5199);
nand U5629 (N_5629,N_5218,N_4936);
or U5630 (N_5630,N_4937,N_4650);
nor U5631 (N_5631,N_5056,N_5188);
nand U5632 (N_5632,N_5150,N_5015);
nand U5633 (N_5633,N_4528,N_5049);
xnor U5634 (N_5634,N_5081,N_5130);
nand U5635 (N_5635,N_5030,N_4808);
nor U5636 (N_5636,N_5179,N_4976);
nor U5637 (N_5637,N_4605,N_4652);
or U5638 (N_5638,N_4772,N_4528);
or U5639 (N_5639,N_5170,N_4934);
and U5640 (N_5640,N_4754,N_5170);
and U5641 (N_5641,N_4536,N_4933);
and U5642 (N_5642,N_4862,N_4666);
nand U5643 (N_5643,N_5041,N_4652);
nor U5644 (N_5644,N_5168,N_4677);
or U5645 (N_5645,N_5127,N_4557);
or U5646 (N_5646,N_4590,N_5242);
xor U5647 (N_5647,N_4600,N_4888);
xnor U5648 (N_5648,N_4502,N_4683);
or U5649 (N_5649,N_5025,N_4590);
or U5650 (N_5650,N_5228,N_4836);
or U5651 (N_5651,N_4649,N_4948);
and U5652 (N_5652,N_4742,N_5014);
nor U5653 (N_5653,N_5054,N_4544);
xor U5654 (N_5654,N_4644,N_5245);
xnor U5655 (N_5655,N_5246,N_4742);
nand U5656 (N_5656,N_5221,N_5021);
or U5657 (N_5657,N_4865,N_4507);
nand U5658 (N_5658,N_4667,N_5009);
nor U5659 (N_5659,N_4735,N_4763);
and U5660 (N_5660,N_4842,N_4592);
xnor U5661 (N_5661,N_4873,N_5146);
and U5662 (N_5662,N_4933,N_4904);
nor U5663 (N_5663,N_4642,N_5028);
nor U5664 (N_5664,N_5196,N_4875);
and U5665 (N_5665,N_4993,N_4642);
or U5666 (N_5666,N_4935,N_4511);
or U5667 (N_5667,N_4814,N_5015);
nand U5668 (N_5668,N_4965,N_5244);
or U5669 (N_5669,N_4868,N_4605);
and U5670 (N_5670,N_5216,N_5156);
and U5671 (N_5671,N_4997,N_5040);
and U5672 (N_5672,N_4971,N_4790);
or U5673 (N_5673,N_4740,N_4625);
or U5674 (N_5674,N_4778,N_4869);
xor U5675 (N_5675,N_4972,N_5020);
nand U5676 (N_5676,N_4759,N_4653);
nand U5677 (N_5677,N_4851,N_4522);
and U5678 (N_5678,N_5188,N_4934);
or U5679 (N_5679,N_5023,N_5165);
nor U5680 (N_5680,N_5056,N_4551);
nor U5681 (N_5681,N_4868,N_4768);
nor U5682 (N_5682,N_4675,N_5203);
nand U5683 (N_5683,N_5206,N_4578);
xor U5684 (N_5684,N_5102,N_4788);
or U5685 (N_5685,N_4926,N_5176);
nor U5686 (N_5686,N_5206,N_5002);
xor U5687 (N_5687,N_4964,N_4738);
nand U5688 (N_5688,N_5173,N_4701);
or U5689 (N_5689,N_5012,N_4877);
nand U5690 (N_5690,N_4842,N_4907);
or U5691 (N_5691,N_5041,N_5164);
or U5692 (N_5692,N_4575,N_4814);
nor U5693 (N_5693,N_5116,N_4895);
xnor U5694 (N_5694,N_4632,N_5214);
or U5695 (N_5695,N_4776,N_5226);
nand U5696 (N_5696,N_4596,N_5247);
nand U5697 (N_5697,N_5093,N_5215);
and U5698 (N_5698,N_5184,N_4720);
and U5699 (N_5699,N_5243,N_4828);
nor U5700 (N_5700,N_4929,N_5006);
nand U5701 (N_5701,N_4743,N_4735);
or U5702 (N_5702,N_4701,N_4602);
or U5703 (N_5703,N_5069,N_5108);
nor U5704 (N_5704,N_4806,N_5175);
nor U5705 (N_5705,N_4632,N_5048);
or U5706 (N_5706,N_4964,N_4527);
or U5707 (N_5707,N_4563,N_4692);
or U5708 (N_5708,N_4922,N_5115);
or U5709 (N_5709,N_4895,N_4879);
or U5710 (N_5710,N_4843,N_4872);
and U5711 (N_5711,N_4779,N_4682);
or U5712 (N_5712,N_4798,N_4775);
xor U5713 (N_5713,N_5148,N_4956);
and U5714 (N_5714,N_4875,N_4864);
or U5715 (N_5715,N_4556,N_4903);
nor U5716 (N_5716,N_5102,N_4821);
nor U5717 (N_5717,N_4784,N_4746);
or U5718 (N_5718,N_4908,N_4550);
xnor U5719 (N_5719,N_4639,N_4599);
nand U5720 (N_5720,N_5074,N_5109);
xor U5721 (N_5721,N_4896,N_4971);
nand U5722 (N_5722,N_4878,N_5091);
nand U5723 (N_5723,N_5245,N_4831);
nor U5724 (N_5724,N_4613,N_4971);
xor U5725 (N_5725,N_4704,N_5140);
xnor U5726 (N_5726,N_4561,N_5248);
or U5727 (N_5727,N_4776,N_4983);
and U5728 (N_5728,N_4836,N_4693);
nand U5729 (N_5729,N_4637,N_4855);
nor U5730 (N_5730,N_4838,N_4743);
and U5731 (N_5731,N_5105,N_5060);
xnor U5732 (N_5732,N_4983,N_5171);
xor U5733 (N_5733,N_5222,N_5099);
or U5734 (N_5734,N_5126,N_5168);
and U5735 (N_5735,N_4787,N_4780);
nand U5736 (N_5736,N_4714,N_4857);
xnor U5737 (N_5737,N_4539,N_4576);
nand U5738 (N_5738,N_5109,N_5004);
nand U5739 (N_5739,N_5104,N_5013);
and U5740 (N_5740,N_4983,N_5092);
nand U5741 (N_5741,N_5200,N_5226);
nand U5742 (N_5742,N_5159,N_5120);
nor U5743 (N_5743,N_5049,N_5215);
xor U5744 (N_5744,N_4875,N_4787);
nor U5745 (N_5745,N_4886,N_5222);
xor U5746 (N_5746,N_4806,N_4626);
or U5747 (N_5747,N_4741,N_4858);
nand U5748 (N_5748,N_4884,N_4773);
xnor U5749 (N_5749,N_4696,N_4513);
nor U5750 (N_5750,N_4784,N_4984);
nor U5751 (N_5751,N_5004,N_4555);
and U5752 (N_5752,N_4516,N_4500);
nand U5753 (N_5753,N_5130,N_4613);
or U5754 (N_5754,N_4740,N_4787);
xor U5755 (N_5755,N_5103,N_4796);
and U5756 (N_5756,N_4628,N_4572);
nand U5757 (N_5757,N_4554,N_4584);
nor U5758 (N_5758,N_4650,N_4819);
xor U5759 (N_5759,N_4848,N_4526);
nand U5760 (N_5760,N_4671,N_4859);
nor U5761 (N_5761,N_4731,N_4623);
nor U5762 (N_5762,N_4710,N_4584);
or U5763 (N_5763,N_4716,N_5194);
nand U5764 (N_5764,N_4882,N_4524);
nand U5765 (N_5765,N_5143,N_4709);
nand U5766 (N_5766,N_5228,N_4552);
and U5767 (N_5767,N_4787,N_4558);
nand U5768 (N_5768,N_4999,N_4514);
nor U5769 (N_5769,N_4690,N_4878);
and U5770 (N_5770,N_4938,N_5206);
nor U5771 (N_5771,N_5041,N_4865);
nand U5772 (N_5772,N_4611,N_5160);
nor U5773 (N_5773,N_4947,N_4631);
nor U5774 (N_5774,N_4812,N_4721);
nand U5775 (N_5775,N_5055,N_4601);
nand U5776 (N_5776,N_4906,N_4852);
and U5777 (N_5777,N_4758,N_4598);
nand U5778 (N_5778,N_4696,N_4735);
or U5779 (N_5779,N_4907,N_4871);
xnor U5780 (N_5780,N_4925,N_4711);
or U5781 (N_5781,N_5162,N_4848);
xor U5782 (N_5782,N_5207,N_4913);
nand U5783 (N_5783,N_5128,N_5190);
and U5784 (N_5784,N_5194,N_4809);
nand U5785 (N_5785,N_4940,N_5169);
nor U5786 (N_5786,N_4748,N_4802);
xor U5787 (N_5787,N_4955,N_4681);
nor U5788 (N_5788,N_4695,N_4613);
nand U5789 (N_5789,N_5190,N_5072);
nand U5790 (N_5790,N_4971,N_5045);
nand U5791 (N_5791,N_5145,N_4574);
and U5792 (N_5792,N_5020,N_4655);
and U5793 (N_5793,N_5151,N_4806);
and U5794 (N_5794,N_4511,N_4851);
xor U5795 (N_5795,N_5085,N_5227);
or U5796 (N_5796,N_4553,N_5073);
xor U5797 (N_5797,N_5210,N_5197);
xor U5798 (N_5798,N_4930,N_5047);
xnor U5799 (N_5799,N_4928,N_4510);
or U5800 (N_5800,N_4518,N_4612);
and U5801 (N_5801,N_4781,N_4872);
and U5802 (N_5802,N_4733,N_5022);
xor U5803 (N_5803,N_4582,N_5046);
nand U5804 (N_5804,N_4634,N_4973);
and U5805 (N_5805,N_4970,N_5093);
and U5806 (N_5806,N_4954,N_5221);
nand U5807 (N_5807,N_5022,N_4999);
and U5808 (N_5808,N_4971,N_5157);
xor U5809 (N_5809,N_4731,N_4627);
and U5810 (N_5810,N_4525,N_5083);
and U5811 (N_5811,N_4871,N_5031);
nor U5812 (N_5812,N_4515,N_5131);
or U5813 (N_5813,N_4955,N_4727);
and U5814 (N_5814,N_4780,N_4961);
or U5815 (N_5815,N_4761,N_4681);
nor U5816 (N_5816,N_4663,N_4580);
nand U5817 (N_5817,N_5074,N_4932);
or U5818 (N_5818,N_4940,N_5149);
nor U5819 (N_5819,N_4655,N_4573);
or U5820 (N_5820,N_5027,N_5066);
and U5821 (N_5821,N_4701,N_4680);
and U5822 (N_5822,N_5035,N_4595);
nand U5823 (N_5823,N_4918,N_4571);
nor U5824 (N_5824,N_4606,N_4527);
nor U5825 (N_5825,N_5219,N_5005);
nand U5826 (N_5826,N_4521,N_4674);
and U5827 (N_5827,N_5043,N_4702);
nand U5828 (N_5828,N_5108,N_5247);
or U5829 (N_5829,N_5139,N_4804);
nand U5830 (N_5830,N_5125,N_4580);
nor U5831 (N_5831,N_4876,N_4786);
nor U5832 (N_5832,N_4638,N_4915);
xnor U5833 (N_5833,N_4886,N_5038);
nand U5834 (N_5834,N_5177,N_4682);
and U5835 (N_5835,N_5126,N_4596);
nand U5836 (N_5836,N_5070,N_4756);
nor U5837 (N_5837,N_4500,N_5150);
nand U5838 (N_5838,N_4562,N_5085);
and U5839 (N_5839,N_5060,N_5119);
or U5840 (N_5840,N_4614,N_4894);
nor U5841 (N_5841,N_4770,N_5072);
nand U5842 (N_5842,N_4557,N_4864);
nand U5843 (N_5843,N_5147,N_4587);
and U5844 (N_5844,N_5009,N_5220);
or U5845 (N_5845,N_4892,N_5186);
nor U5846 (N_5846,N_4967,N_4568);
or U5847 (N_5847,N_4624,N_4655);
or U5848 (N_5848,N_5232,N_4825);
and U5849 (N_5849,N_5046,N_5155);
xnor U5850 (N_5850,N_4738,N_5127);
or U5851 (N_5851,N_5183,N_5165);
and U5852 (N_5852,N_5006,N_5216);
nor U5853 (N_5853,N_4604,N_4682);
and U5854 (N_5854,N_5045,N_4619);
or U5855 (N_5855,N_5153,N_4682);
nand U5856 (N_5856,N_5173,N_4821);
and U5857 (N_5857,N_4519,N_4739);
nand U5858 (N_5858,N_4504,N_4641);
and U5859 (N_5859,N_5047,N_4888);
xor U5860 (N_5860,N_4717,N_4832);
or U5861 (N_5861,N_4944,N_4524);
xnor U5862 (N_5862,N_4568,N_4934);
and U5863 (N_5863,N_5185,N_4721);
nor U5864 (N_5864,N_5120,N_5205);
nand U5865 (N_5865,N_4999,N_5032);
or U5866 (N_5866,N_5204,N_4592);
or U5867 (N_5867,N_4538,N_5208);
xor U5868 (N_5868,N_5051,N_4506);
and U5869 (N_5869,N_5022,N_5226);
nand U5870 (N_5870,N_4741,N_4656);
nand U5871 (N_5871,N_4582,N_4734);
or U5872 (N_5872,N_4998,N_5147);
xnor U5873 (N_5873,N_4544,N_5216);
xnor U5874 (N_5874,N_5150,N_4556);
nand U5875 (N_5875,N_4568,N_4744);
xnor U5876 (N_5876,N_4621,N_4738);
xor U5877 (N_5877,N_5171,N_4755);
or U5878 (N_5878,N_4987,N_4599);
xor U5879 (N_5879,N_4534,N_5212);
nand U5880 (N_5880,N_5123,N_4790);
and U5881 (N_5881,N_4511,N_4607);
and U5882 (N_5882,N_4858,N_5171);
nor U5883 (N_5883,N_4807,N_4624);
nand U5884 (N_5884,N_4894,N_4534);
nor U5885 (N_5885,N_4999,N_4862);
nor U5886 (N_5886,N_4791,N_5142);
nand U5887 (N_5887,N_4913,N_4682);
nor U5888 (N_5888,N_5216,N_4594);
or U5889 (N_5889,N_4602,N_4827);
nor U5890 (N_5890,N_4923,N_5202);
nor U5891 (N_5891,N_5049,N_4782);
or U5892 (N_5892,N_5009,N_4614);
or U5893 (N_5893,N_5225,N_5196);
nand U5894 (N_5894,N_4534,N_4764);
and U5895 (N_5895,N_5152,N_5229);
and U5896 (N_5896,N_4854,N_5015);
and U5897 (N_5897,N_5170,N_4722);
nor U5898 (N_5898,N_4575,N_4830);
xnor U5899 (N_5899,N_5212,N_4772);
nor U5900 (N_5900,N_4535,N_5163);
or U5901 (N_5901,N_5010,N_4550);
or U5902 (N_5902,N_4782,N_4542);
or U5903 (N_5903,N_4579,N_4721);
and U5904 (N_5904,N_4865,N_4868);
nand U5905 (N_5905,N_4621,N_4544);
xnor U5906 (N_5906,N_4942,N_4785);
nand U5907 (N_5907,N_4739,N_4738);
and U5908 (N_5908,N_5105,N_5017);
xor U5909 (N_5909,N_4689,N_4773);
and U5910 (N_5910,N_4591,N_5096);
nand U5911 (N_5911,N_4511,N_4587);
or U5912 (N_5912,N_4680,N_4957);
and U5913 (N_5913,N_4959,N_4673);
nor U5914 (N_5914,N_4567,N_5201);
or U5915 (N_5915,N_5143,N_5049);
xnor U5916 (N_5916,N_4525,N_5115);
nand U5917 (N_5917,N_4927,N_5089);
nor U5918 (N_5918,N_5161,N_4547);
nand U5919 (N_5919,N_5170,N_5061);
nand U5920 (N_5920,N_4705,N_5231);
or U5921 (N_5921,N_4630,N_5045);
and U5922 (N_5922,N_5113,N_5083);
and U5923 (N_5923,N_5170,N_5202);
nand U5924 (N_5924,N_4945,N_5053);
or U5925 (N_5925,N_5217,N_4680);
nand U5926 (N_5926,N_4683,N_5111);
nor U5927 (N_5927,N_5061,N_4546);
nor U5928 (N_5928,N_5215,N_4516);
and U5929 (N_5929,N_4913,N_4678);
nor U5930 (N_5930,N_5115,N_5111);
nand U5931 (N_5931,N_4911,N_4972);
nor U5932 (N_5932,N_4703,N_5167);
xor U5933 (N_5933,N_4816,N_4873);
xor U5934 (N_5934,N_4771,N_5003);
or U5935 (N_5935,N_5116,N_4533);
or U5936 (N_5936,N_4979,N_4782);
nand U5937 (N_5937,N_4625,N_4939);
xnor U5938 (N_5938,N_4666,N_5044);
and U5939 (N_5939,N_5014,N_4980);
nand U5940 (N_5940,N_4758,N_4681);
nor U5941 (N_5941,N_5011,N_4659);
nand U5942 (N_5942,N_4907,N_4784);
nor U5943 (N_5943,N_5113,N_4992);
nor U5944 (N_5944,N_4999,N_5099);
xor U5945 (N_5945,N_4658,N_4775);
nor U5946 (N_5946,N_4870,N_4962);
and U5947 (N_5947,N_4632,N_5231);
nor U5948 (N_5948,N_4965,N_4521);
nor U5949 (N_5949,N_5229,N_4848);
and U5950 (N_5950,N_5227,N_4731);
and U5951 (N_5951,N_4541,N_4953);
nor U5952 (N_5952,N_4850,N_4603);
and U5953 (N_5953,N_5001,N_4715);
xor U5954 (N_5954,N_5136,N_4579);
or U5955 (N_5955,N_4736,N_4879);
nor U5956 (N_5956,N_4871,N_5171);
nand U5957 (N_5957,N_4788,N_4894);
or U5958 (N_5958,N_4582,N_4658);
nor U5959 (N_5959,N_4581,N_4622);
or U5960 (N_5960,N_4686,N_4594);
or U5961 (N_5961,N_4903,N_5136);
or U5962 (N_5962,N_4660,N_4529);
nor U5963 (N_5963,N_4571,N_5134);
nand U5964 (N_5964,N_4837,N_5058);
and U5965 (N_5965,N_4738,N_5019);
nand U5966 (N_5966,N_5049,N_4527);
nand U5967 (N_5967,N_4628,N_5249);
nor U5968 (N_5968,N_5000,N_5222);
nand U5969 (N_5969,N_5174,N_4765);
nand U5970 (N_5970,N_4828,N_4726);
xnor U5971 (N_5971,N_4993,N_4878);
xor U5972 (N_5972,N_4673,N_5022);
or U5973 (N_5973,N_4543,N_5011);
xnor U5974 (N_5974,N_4580,N_4645);
xor U5975 (N_5975,N_4608,N_5128);
xnor U5976 (N_5976,N_4755,N_4679);
nor U5977 (N_5977,N_5010,N_4982);
xor U5978 (N_5978,N_5202,N_4908);
nor U5979 (N_5979,N_4760,N_5190);
nand U5980 (N_5980,N_5153,N_5248);
and U5981 (N_5981,N_5198,N_4734);
and U5982 (N_5982,N_5186,N_4779);
or U5983 (N_5983,N_4564,N_4682);
nand U5984 (N_5984,N_5180,N_4523);
xnor U5985 (N_5985,N_5068,N_4514);
nor U5986 (N_5986,N_4725,N_5088);
nor U5987 (N_5987,N_4764,N_4628);
nor U5988 (N_5988,N_5095,N_4999);
and U5989 (N_5989,N_4904,N_4746);
xnor U5990 (N_5990,N_4893,N_4840);
and U5991 (N_5991,N_4835,N_4739);
nor U5992 (N_5992,N_5062,N_4642);
and U5993 (N_5993,N_4772,N_5186);
xnor U5994 (N_5994,N_4847,N_5131);
or U5995 (N_5995,N_4753,N_4588);
and U5996 (N_5996,N_5198,N_4532);
xor U5997 (N_5997,N_5041,N_4530);
and U5998 (N_5998,N_4664,N_4981);
and U5999 (N_5999,N_5113,N_5047);
and U6000 (N_6000,N_5505,N_5358);
nand U6001 (N_6001,N_5584,N_5481);
xnor U6002 (N_6002,N_5471,N_5656);
nor U6003 (N_6003,N_5486,N_5359);
nor U6004 (N_6004,N_5620,N_5690);
nand U6005 (N_6005,N_5939,N_5305);
and U6006 (N_6006,N_5614,N_5654);
or U6007 (N_6007,N_5983,N_5876);
or U6008 (N_6008,N_5364,N_5804);
or U6009 (N_6009,N_5677,N_5896);
and U6010 (N_6010,N_5310,N_5856);
or U6011 (N_6011,N_5565,N_5631);
nand U6012 (N_6012,N_5749,N_5919);
nor U6013 (N_6013,N_5659,N_5688);
and U6014 (N_6014,N_5523,N_5957);
xor U6015 (N_6015,N_5385,N_5517);
and U6016 (N_6016,N_5904,N_5586);
nor U6017 (N_6017,N_5765,N_5768);
xor U6018 (N_6018,N_5321,N_5449);
nor U6019 (N_6019,N_5526,N_5662);
nand U6020 (N_6020,N_5929,N_5763);
and U6021 (N_6021,N_5412,N_5282);
and U6022 (N_6022,N_5545,N_5989);
nand U6023 (N_6023,N_5493,N_5743);
and U6024 (N_6024,N_5529,N_5918);
xor U6025 (N_6025,N_5316,N_5426);
xor U6026 (N_6026,N_5834,N_5599);
nor U6027 (N_6027,N_5346,N_5858);
and U6028 (N_6028,N_5648,N_5562);
nor U6029 (N_6029,N_5891,N_5559);
and U6030 (N_6030,N_5377,N_5499);
or U6031 (N_6031,N_5561,N_5937);
nor U6032 (N_6032,N_5522,N_5827);
xnor U6033 (N_6033,N_5831,N_5387);
nand U6034 (N_6034,N_5616,N_5572);
nor U6035 (N_6035,N_5794,N_5269);
and U6036 (N_6036,N_5521,N_5798);
nor U6037 (N_6037,N_5888,N_5301);
nor U6038 (N_6038,N_5382,N_5409);
or U6039 (N_6039,N_5868,N_5520);
and U6040 (N_6040,N_5940,N_5622);
and U6041 (N_6041,N_5698,N_5514);
and U6042 (N_6042,N_5259,N_5276);
xnor U6043 (N_6043,N_5598,N_5476);
and U6044 (N_6044,N_5440,N_5920);
and U6045 (N_6045,N_5328,N_5578);
xnor U6046 (N_6046,N_5960,N_5826);
and U6047 (N_6047,N_5341,N_5390);
nor U6048 (N_6048,N_5907,N_5905);
or U6049 (N_6049,N_5571,N_5557);
and U6050 (N_6050,N_5825,N_5287);
nor U6051 (N_6051,N_5815,N_5878);
nor U6052 (N_6052,N_5666,N_5435);
nor U6053 (N_6053,N_5954,N_5619);
nand U6054 (N_6054,N_5258,N_5291);
nand U6055 (N_6055,N_5946,N_5386);
nand U6056 (N_6056,N_5976,N_5901);
nand U6057 (N_6057,N_5711,N_5309);
and U6058 (N_6058,N_5267,N_5932);
or U6059 (N_6059,N_5780,N_5326);
nor U6060 (N_6060,N_5478,N_5632);
and U6061 (N_6061,N_5781,N_5956);
or U6062 (N_6062,N_5357,N_5883);
xnor U6063 (N_6063,N_5761,N_5495);
and U6064 (N_6064,N_5997,N_5706);
and U6065 (N_6065,N_5560,N_5685);
and U6066 (N_6066,N_5348,N_5992);
and U6067 (N_6067,N_5371,N_5772);
nor U6068 (N_6068,N_5759,N_5353);
xnor U6069 (N_6069,N_5338,N_5516);
and U6070 (N_6070,N_5424,N_5935);
and U6071 (N_6071,N_5702,N_5882);
nand U6072 (N_6072,N_5871,N_5959);
and U6073 (N_6073,N_5621,N_5398);
and U6074 (N_6074,N_5392,N_5552);
nand U6075 (N_6075,N_5419,N_5263);
or U6076 (N_6076,N_5617,N_5474);
xnor U6077 (N_6077,N_5953,N_5579);
nor U6078 (N_6078,N_5397,N_5757);
nand U6079 (N_6079,N_5463,N_5543);
or U6080 (N_6080,N_5410,N_5497);
or U6081 (N_6081,N_5381,N_5861);
or U6082 (N_6082,N_5694,N_5865);
xor U6083 (N_6083,N_5756,N_5597);
and U6084 (N_6084,N_5777,N_5480);
or U6085 (N_6085,N_5404,N_5796);
xor U6086 (N_6086,N_5418,N_5963);
xnor U6087 (N_6087,N_5949,N_5285);
or U6088 (N_6088,N_5642,N_5665);
and U6089 (N_6089,N_5279,N_5573);
or U6090 (N_6090,N_5300,N_5890);
xnor U6091 (N_6091,N_5867,N_5695);
nand U6092 (N_6092,N_5933,N_5802);
and U6093 (N_6093,N_5697,N_5958);
and U6094 (N_6094,N_5549,N_5721);
nor U6095 (N_6095,N_5807,N_5917);
or U6096 (N_6096,N_5680,N_5313);
xor U6097 (N_6097,N_5658,N_5910);
nand U6098 (N_6098,N_5824,N_5509);
xor U6099 (N_6099,N_5335,N_5699);
nor U6100 (N_6100,N_5678,N_5964);
nand U6101 (N_6101,N_5587,N_5539);
and U6102 (N_6102,N_5769,N_5663);
xor U6103 (N_6103,N_5512,N_5754);
and U6104 (N_6104,N_5361,N_5446);
xnor U6105 (N_6105,N_5811,N_5906);
and U6106 (N_6106,N_5808,N_5594);
nor U6107 (N_6107,N_5576,N_5912);
xor U6108 (N_6108,N_5582,N_5724);
xnor U6109 (N_6109,N_5644,N_5840);
nor U6110 (N_6110,N_5613,N_5433);
or U6111 (N_6111,N_5455,N_5875);
nor U6112 (N_6112,N_5299,N_5558);
nor U6113 (N_6113,N_5720,N_5286);
xor U6114 (N_6114,N_5710,N_5337);
nor U6115 (N_6115,N_5612,N_5730);
nor U6116 (N_6116,N_5672,N_5589);
and U6117 (N_6117,N_5814,N_5687);
or U6118 (N_6118,N_5555,N_5519);
xnor U6119 (N_6119,N_5745,N_5592);
and U6120 (N_6120,N_5792,N_5783);
nand U6121 (N_6121,N_5444,N_5773);
nor U6122 (N_6122,N_5511,N_5360);
xnor U6123 (N_6123,N_5674,N_5640);
xnor U6124 (N_6124,N_5641,N_5835);
nand U6125 (N_6125,N_5948,N_5403);
or U6126 (N_6126,N_5566,N_5268);
nor U6127 (N_6127,N_5971,N_5965);
xnor U6128 (N_6128,N_5507,N_5515);
xnor U6129 (N_6129,N_5547,N_5319);
xor U6130 (N_6130,N_5334,N_5770);
nor U6131 (N_6131,N_5823,N_5731);
and U6132 (N_6132,N_5980,N_5950);
nor U6133 (N_6133,N_5430,N_5943);
xnor U6134 (N_6134,N_5760,N_5624);
nor U6135 (N_6135,N_5652,N_5885);
xor U6136 (N_6136,N_5266,N_5421);
xor U6137 (N_6137,N_5329,N_5298);
xor U6138 (N_6138,N_5289,N_5567);
nand U6139 (N_6139,N_5942,N_5366);
or U6140 (N_6140,N_5590,N_5563);
nor U6141 (N_6141,N_5717,N_5785);
and U6142 (N_6142,N_5502,N_5854);
and U6143 (N_6143,N_5633,N_5669);
nand U6144 (N_6144,N_5927,N_5836);
nand U6145 (N_6145,N_5741,N_5609);
nand U6146 (N_6146,N_5962,N_5275);
or U6147 (N_6147,N_5848,N_5909);
xor U6148 (N_6148,N_5355,N_5250);
nor U6149 (N_6149,N_5857,N_5703);
and U6150 (N_6150,N_5908,N_5924);
nor U6151 (N_6151,N_5413,N_5391);
nor U6152 (N_6152,N_5574,N_5998);
nand U6153 (N_6153,N_5603,N_5568);
and U6154 (N_6154,N_5961,N_5860);
or U6155 (N_6155,N_5414,N_5607);
xor U6156 (N_6156,N_5251,N_5693);
nor U6157 (N_6157,N_5981,N_5786);
xnor U6158 (N_6158,N_5884,N_5593);
and U6159 (N_6159,N_5849,N_5626);
and U6160 (N_6160,N_5683,N_5634);
xnor U6161 (N_6161,N_5722,N_5846);
nand U6162 (N_6162,N_5540,N_5454);
and U6163 (N_6163,N_5452,N_5365);
nor U6164 (N_6164,N_5525,N_5911);
xor U6165 (N_6165,N_5368,N_5635);
nor U6166 (N_6166,N_5342,N_5302);
xnor U6167 (N_6167,N_5931,N_5708);
nor U6168 (N_6168,N_5821,N_5344);
nor U6169 (N_6169,N_5257,N_5615);
nand U6170 (N_6170,N_5689,N_5376);
or U6171 (N_6171,N_5967,N_5822);
and U6172 (N_6172,N_5886,N_5556);
nand U6173 (N_6173,N_5401,N_5716);
and U6174 (N_6174,N_5748,N_5870);
xnor U6175 (N_6175,N_5349,N_5915);
or U6176 (N_6176,N_5438,N_5692);
or U6177 (N_6177,N_5639,N_5793);
nor U6178 (N_6178,N_5696,N_5787);
nand U6179 (N_6179,N_5707,N_5432);
nand U6180 (N_6180,N_5548,N_5325);
nand U6181 (N_6181,N_5406,N_5384);
xnor U6182 (N_6182,N_5637,N_5420);
nand U6183 (N_6183,N_5926,N_5468);
nor U6184 (N_6184,N_5475,N_5736);
or U6185 (N_6185,N_5375,N_5766);
and U6186 (N_6186,N_5874,N_5427);
or U6187 (N_6187,N_5537,N_5664);
and U6188 (N_6188,N_5892,N_5531);
nor U6189 (N_6189,N_5354,N_5280);
xnor U6190 (N_6190,N_5800,N_5378);
nor U6191 (N_6191,N_5852,N_5496);
xor U6192 (N_6192,N_5513,N_5504);
nor U6193 (N_6193,N_5510,N_5979);
and U6194 (N_6194,N_5746,N_5484);
xnor U6195 (N_6195,N_5944,N_5439);
or U6196 (N_6196,N_5791,N_5994);
or U6197 (N_6197,N_5459,N_5799);
nand U6198 (N_6198,N_5618,N_5491);
or U6199 (N_6199,N_5370,N_5832);
xnor U6200 (N_6200,N_5623,N_5859);
and U6201 (N_6201,N_5894,N_5755);
and U6202 (N_6202,N_5996,N_5869);
nand U6203 (N_6203,N_5945,N_5638);
xnor U6204 (N_6204,N_5788,N_5372);
and U6205 (N_6205,N_5564,N_5281);
or U6206 (N_6206,N_5645,N_5803);
or U6207 (N_6207,N_5383,N_5987);
xnor U6208 (N_6208,N_5627,N_5294);
nand U6209 (N_6209,N_5367,N_5661);
or U6210 (N_6210,N_5501,N_5500);
and U6211 (N_6211,N_5657,N_5828);
xnor U6212 (N_6212,N_5396,N_5443);
or U6213 (N_6213,N_5629,N_5879);
and U6214 (N_6214,N_5389,N_5817);
or U6215 (N_6215,N_5318,N_5925);
or U6216 (N_6216,N_5352,N_5679);
nand U6217 (N_6217,N_5388,N_5457);
xor U6218 (N_6218,N_5668,N_5415);
nor U6219 (N_6219,N_5608,N_5993);
and U6220 (N_6220,N_5734,N_5819);
or U6221 (N_6221,N_5751,N_5725);
or U6222 (N_6222,N_5843,N_5542);
nor U6223 (N_6223,N_5982,N_5782);
nand U6224 (N_6224,N_5728,N_5533);
nand U6225 (N_6225,N_5900,N_5393);
or U6226 (N_6226,N_5467,N_5465);
xnor U6227 (N_6227,N_5585,N_5270);
nand U6228 (N_6228,N_5830,N_5534);
xor U6229 (N_6229,N_5308,N_5527);
nor U6230 (N_6230,N_5739,N_5262);
or U6231 (N_6231,N_5758,N_5253);
nor U6232 (N_6232,N_5649,N_5673);
nand U6233 (N_6233,N_5841,N_5974);
xnor U6234 (N_6234,N_5343,N_5999);
xnor U6235 (N_6235,N_5317,N_5577);
and U6236 (N_6236,N_5735,N_5880);
xor U6237 (N_6237,N_5411,N_5417);
or U6238 (N_6238,N_5686,N_5536);
nand U6239 (N_6239,N_5273,N_5283);
xnor U6240 (N_6240,N_5336,N_5727);
and U6241 (N_6241,N_5704,N_5379);
nor U6242 (N_6242,N_5719,N_5889);
nand U6243 (N_6243,N_5818,N_5469);
nand U6244 (N_6244,N_5535,N_5899);
and U6245 (N_6245,N_5580,N_5277);
or U6246 (N_6246,N_5296,N_5995);
nor U6247 (N_6247,N_5356,N_5646);
or U6248 (N_6248,N_5255,N_5492);
nor U6249 (N_6249,N_5778,N_5851);
nand U6250 (N_6250,N_5464,N_5332);
xnor U6251 (N_6251,N_5812,N_5729);
and U6252 (N_6252,N_5847,N_5307);
xor U6253 (N_6253,N_5458,N_5330);
or U6254 (N_6254,N_5625,N_5952);
xnor U6255 (N_6255,N_5333,N_5647);
and U6256 (N_6256,N_5487,N_5605);
or U6257 (N_6257,N_5866,N_5312);
or U6258 (N_6258,N_5604,N_5714);
nand U6259 (N_6259,N_5553,N_5709);
xnor U6260 (N_6260,N_5477,N_5339);
nor U6261 (N_6261,N_5350,N_5887);
xor U6262 (N_6262,N_5284,N_5450);
and U6263 (N_6263,N_5256,N_5570);
and U6264 (N_6264,N_5839,N_5790);
xor U6265 (N_6265,N_5797,N_5295);
nor U6266 (N_6266,N_5304,N_5643);
nor U6267 (N_6267,N_5423,N_5479);
nand U6268 (N_6268,N_5569,N_5506);
and U6269 (N_6269,N_5340,N_5715);
and U6270 (N_6270,N_5528,N_5445);
nor U6271 (N_6271,N_5872,N_5855);
xor U6272 (N_6272,N_5877,N_5290);
xor U6273 (N_6273,N_5809,N_5737);
and U6274 (N_6274,N_5744,N_5740);
or U6275 (N_6275,N_5903,N_5820);
or U6276 (N_6276,N_5705,N_5611);
nor U6277 (N_6277,N_5742,N_5498);
or U6278 (N_6278,N_5676,N_5544);
or U6279 (N_6279,N_5524,N_5532);
xor U6280 (N_6280,N_5873,N_5916);
and U6281 (N_6281,N_5436,N_5779);
xor U6282 (N_6282,N_5466,N_5898);
or U6283 (N_6283,N_5970,N_5303);
and U6284 (N_6284,N_5315,N_5682);
or U6285 (N_6285,N_5893,N_5601);
and U6286 (N_6286,N_5591,N_5451);
and U6287 (N_6287,N_5395,N_5650);
or U6288 (N_6288,N_5951,N_5684);
xor U6289 (N_6289,N_5272,N_5374);
xnor U6290 (N_6290,N_5844,N_5806);
and U6291 (N_6291,N_5628,N_5984);
xnor U6292 (N_6292,N_5726,N_5816);
and U6293 (N_6293,N_5408,N_5394);
or U6294 (N_6294,N_5482,N_5947);
and U6295 (N_6295,N_5362,N_5462);
xor U6296 (N_6296,N_5853,N_5972);
xor U6297 (N_6297,N_5837,N_5265);
xnor U6298 (N_6298,N_5402,N_5829);
or U6299 (N_6299,N_5595,N_5986);
or U6300 (N_6300,N_5764,N_5936);
xor U6301 (N_6301,N_5311,N_5771);
xnor U6302 (N_6302,N_5271,N_5448);
or U6303 (N_6303,N_5314,N_5700);
and U6304 (N_6304,N_5470,N_5456);
xnor U6305 (N_6305,N_5508,N_5551);
xor U6306 (N_6306,N_5288,N_5518);
xnor U6307 (N_6307,N_5322,N_5363);
xor U6308 (N_6308,N_5345,N_5431);
and U6309 (N_6309,N_5541,N_5554);
nor U6310 (N_6310,N_5713,N_5845);
xor U6311 (N_6311,N_5733,N_5838);
nand U6312 (N_6312,N_5968,N_5297);
nor U6313 (N_6313,N_5400,N_5938);
xnor U6314 (N_6314,N_5373,N_5775);
or U6315 (N_6315,N_5813,N_5442);
and U6316 (N_6316,N_5895,N_5913);
or U6317 (N_6317,N_5453,N_5437);
xor U6318 (N_6318,N_5575,N_5934);
or U6319 (N_6319,N_5583,N_5399);
or U6320 (N_6320,N_5795,N_5973);
or U6321 (N_6321,N_5600,N_5490);
or U6322 (N_6322,N_5407,N_5784);
and U6323 (N_6323,N_5293,N_5331);
and U6324 (N_6324,N_5347,N_5588);
or U6325 (N_6325,N_5955,N_5850);
xnor U6326 (N_6326,N_5606,N_5789);
xor U6327 (N_6327,N_5546,N_5767);
nand U6328 (N_6328,N_5667,N_5750);
and U6329 (N_6329,N_5655,N_5923);
xor U6330 (N_6330,N_5380,N_5675);
nand U6331 (N_6331,N_5966,N_5636);
nand U6332 (N_6332,N_5862,N_5902);
nor U6333 (N_6333,N_5712,N_5774);
nand U6334 (N_6334,N_5292,N_5753);
and U6335 (N_6335,N_5985,N_5425);
xnor U6336 (N_6336,N_5941,N_5723);
nor U6337 (N_6337,N_5278,N_5416);
and U6338 (N_6338,N_5428,N_5473);
or U6339 (N_6339,N_5261,N_5581);
and U6340 (N_6340,N_5842,N_5660);
or U6341 (N_6341,N_5969,N_5732);
or U6342 (N_6342,N_5460,N_5488);
nor U6343 (N_6343,N_5977,N_5441);
xnor U6344 (N_6344,N_5671,N_5429);
nand U6345 (N_6345,N_5434,N_5461);
nand U6346 (N_6346,N_5805,N_5405);
xnor U6347 (N_6347,N_5762,N_5485);
nand U6348 (N_6348,N_5738,N_5254);
and U6349 (N_6349,N_5550,N_5610);
or U6350 (N_6350,N_5991,N_5320);
nor U6351 (N_6351,N_5921,N_5327);
or U6352 (N_6352,N_5833,N_5494);
or U6353 (N_6353,N_5530,N_5447);
xor U6354 (N_6354,N_5747,N_5701);
xor U6355 (N_6355,N_5914,N_5990);
nand U6356 (N_6356,N_5988,N_5670);
nor U6357 (N_6357,N_5928,N_5252);
or U6358 (N_6358,N_5691,N_5653);
and U6359 (N_6359,N_5881,N_5260);
xnor U6360 (N_6360,N_5503,N_5538);
nor U6361 (N_6361,N_5472,N_5274);
or U6362 (N_6362,N_5489,N_5264);
nor U6363 (N_6363,N_5369,N_5324);
nand U6364 (N_6364,N_5975,N_5801);
nor U6365 (N_6365,N_5718,N_5351);
xnor U6366 (N_6366,N_5306,N_5422);
xnor U6367 (N_6367,N_5863,N_5930);
or U6368 (N_6368,N_5864,N_5651);
or U6369 (N_6369,N_5752,N_5978);
xor U6370 (N_6370,N_5483,N_5602);
or U6371 (N_6371,N_5596,N_5810);
or U6372 (N_6372,N_5776,N_5323);
xor U6373 (N_6373,N_5681,N_5922);
xor U6374 (N_6374,N_5630,N_5897);
and U6375 (N_6375,N_5386,N_5835);
and U6376 (N_6376,N_5945,N_5514);
or U6377 (N_6377,N_5440,N_5404);
xor U6378 (N_6378,N_5769,N_5950);
xor U6379 (N_6379,N_5349,N_5638);
nand U6380 (N_6380,N_5706,N_5349);
nor U6381 (N_6381,N_5795,N_5408);
or U6382 (N_6382,N_5880,N_5626);
xor U6383 (N_6383,N_5980,N_5494);
xor U6384 (N_6384,N_5632,N_5633);
or U6385 (N_6385,N_5912,N_5293);
xnor U6386 (N_6386,N_5666,N_5530);
or U6387 (N_6387,N_5845,N_5506);
and U6388 (N_6388,N_5391,N_5478);
or U6389 (N_6389,N_5273,N_5945);
xnor U6390 (N_6390,N_5370,N_5920);
nor U6391 (N_6391,N_5320,N_5630);
nand U6392 (N_6392,N_5779,N_5529);
and U6393 (N_6393,N_5453,N_5264);
nor U6394 (N_6394,N_5802,N_5803);
or U6395 (N_6395,N_5364,N_5274);
or U6396 (N_6396,N_5998,N_5946);
nor U6397 (N_6397,N_5309,N_5654);
nor U6398 (N_6398,N_5610,N_5942);
and U6399 (N_6399,N_5837,N_5841);
nor U6400 (N_6400,N_5397,N_5490);
nand U6401 (N_6401,N_5409,N_5559);
xor U6402 (N_6402,N_5395,N_5997);
and U6403 (N_6403,N_5303,N_5840);
xnor U6404 (N_6404,N_5692,N_5994);
or U6405 (N_6405,N_5644,N_5802);
and U6406 (N_6406,N_5578,N_5777);
or U6407 (N_6407,N_5389,N_5319);
or U6408 (N_6408,N_5994,N_5680);
nor U6409 (N_6409,N_5310,N_5335);
xnor U6410 (N_6410,N_5929,N_5874);
xor U6411 (N_6411,N_5948,N_5283);
or U6412 (N_6412,N_5495,N_5778);
or U6413 (N_6413,N_5318,N_5265);
nand U6414 (N_6414,N_5645,N_5333);
xor U6415 (N_6415,N_5653,N_5309);
or U6416 (N_6416,N_5410,N_5703);
xor U6417 (N_6417,N_5366,N_5525);
xor U6418 (N_6418,N_5384,N_5627);
or U6419 (N_6419,N_5338,N_5373);
nor U6420 (N_6420,N_5701,N_5735);
xnor U6421 (N_6421,N_5447,N_5861);
xnor U6422 (N_6422,N_5572,N_5456);
or U6423 (N_6423,N_5464,N_5269);
nor U6424 (N_6424,N_5549,N_5783);
or U6425 (N_6425,N_5673,N_5485);
or U6426 (N_6426,N_5479,N_5612);
or U6427 (N_6427,N_5429,N_5299);
nor U6428 (N_6428,N_5255,N_5577);
or U6429 (N_6429,N_5771,N_5990);
nand U6430 (N_6430,N_5829,N_5306);
xnor U6431 (N_6431,N_5987,N_5712);
nand U6432 (N_6432,N_5556,N_5982);
or U6433 (N_6433,N_5524,N_5981);
and U6434 (N_6434,N_5295,N_5328);
nor U6435 (N_6435,N_5515,N_5644);
nor U6436 (N_6436,N_5934,N_5255);
and U6437 (N_6437,N_5299,N_5391);
and U6438 (N_6438,N_5988,N_5919);
and U6439 (N_6439,N_5476,N_5516);
xnor U6440 (N_6440,N_5952,N_5778);
or U6441 (N_6441,N_5276,N_5666);
and U6442 (N_6442,N_5322,N_5994);
or U6443 (N_6443,N_5811,N_5750);
nand U6444 (N_6444,N_5808,N_5838);
nand U6445 (N_6445,N_5535,N_5280);
and U6446 (N_6446,N_5656,N_5995);
nand U6447 (N_6447,N_5821,N_5947);
or U6448 (N_6448,N_5931,N_5319);
and U6449 (N_6449,N_5923,N_5699);
or U6450 (N_6450,N_5675,N_5814);
or U6451 (N_6451,N_5915,N_5264);
nand U6452 (N_6452,N_5283,N_5263);
nor U6453 (N_6453,N_5542,N_5431);
or U6454 (N_6454,N_5976,N_5817);
nor U6455 (N_6455,N_5274,N_5314);
or U6456 (N_6456,N_5426,N_5917);
xnor U6457 (N_6457,N_5929,N_5435);
and U6458 (N_6458,N_5561,N_5452);
nor U6459 (N_6459,N_5875,N_5585);
xnor U6460 (N_6460,N_5384,N_5584);
or U6461 (N_6461,N_5632,N_5952);
nand U6462 (N_6462,N_5337,N_5799);
and U6463 (N_6463,N_5818,N_5392);
nor U6464 (N_6464,N_5672,N_5254);
nand U6465 (N_6465,N_5598,N_5551);
nand U6466 (N_6466,N_5257,N_5958);
or U6467 (N_6467,N_5570,N_5658);
and U6468 (N_6468,N_5331,N_5296);
and U6469 (N_6469,N_5285,N_5970);
xor U6470 (N_6470,N_5409,N_5842);
and U6471 (N_6471,N_5635,N_5611);
and U6472 (N_6472,N_5692,N_5803);
nor U6473 (N_6473,N_5766,N_5597);
xnor U6474 (N_6474,N_5646,N_5759);
xor U6475 (N_6475,N_5524,N_5947);
or U6476 (N_6476,N_5752,N_5376);
nor U6477 (N_6477,N_5913,N_5934);
nand U6478 (N_6478,N_5621,N_5917);
and U6479 (N_6479,N_5796,N_5399);
or U6480 (N_6480,N_5330,N_5913);
nor U6481 (N_6481,N_5596,N_5291);
nand U6482 (N_6482,N_5500,N_5686);
or U6483 (N_6483,N_5750,N_5743);
nor U6484 (N_6484,N_5744,N_5333);
nor U6485 (N_6485,N_5866,N_5683);
nand U6486 (N_6486,N_5297,N_5318);
or U6487 (N_6487,N_5724,N_5450);
and U6488 (N_6488,N_5582,N_5830);
and U6489 (N_6489,N_5572,N_5875);
nand U6490 (N_6490,N_5343,N_5700);
nor U6491 (N_6491,N_5860,N_5769);
and U6492 (N_6492,N_5465,N_5923);
or U6493 (N_6493,N_5334,N_5477);
nand U6494 (N_6494,N_5719,N_5621);
nand U6495 (N_6495,N_5483,N_5392);
nand U6496 (N_6496,N_5731,N_5699);
xor U6497 (N_6497,N_5263,N_5252);
xnor U6498 (N_6498,N_5329,N_5864);
nand U6499 (N_6499,N_5636,N_5765);
or U6500 (N_6500,N_5659,N_5897);
or U6501 (N_6501,N_5991,N_5382);
and U6502 (N_6502,N_5263,N_5722);
and U6503 (N_6503,N_5996,N_5368);
or U6504 (N_6504,N_5581,N_5526);
nand U6505 (N_6505,N_5664,N_5508);
and U6506 (N_6506,N_5493,N_5545);
xor U6507 (N_6507,N_5800,N_5563);
xor U6508 (N_6508,N_5550,N_5378);
xor U6509 (N_6509,N_5461,N_5561);
xor U6510 (N_6510,N_5675,N_5385);
or U6511 (N_6511,N_5379,N_5735);
and U6512 (N_6512,N_5862,N_5637);
or U6513 (N_6513,N_5908,N_5976);
nand U6514 (N_6514,N_5673,N_5543);
xor U6515 (N_6515,N_5885,N_5716);
nor U6516 (N_6516,N_5897,N_5403);
or U6517 (N_6517,N_5843,N_5700);
and U6518 (N_6518,N_5526,N_5468);
or U6519 (N_6519,N_5835,N_5398);
xor U6520 (N_6520,N_5282,N_5376);
and U6521 (N_6521,N_5394,N_5384);
and U6522 (N_6522,N_5801,N_5341);
nand U6523 (N_6523,N_5933,N_5639);
nand U6524 (N_6524,N_5402,N_5362);
or U6525 (N_6525,N_5809,N_5791);
nor U6526 (N_6526,N_5451,N_5533);
or U6527 (N_6527,N_5315,N_5283);
xnor U6528 (N_6528,N_5854,N_5439);
nand U6529 (N_6529,N_5541,N_5851);
nor U6530 (N_6530,N_5770,N_5669);
nand U6531 (N_6531,N_5305,N_5440);
nor U6532 (N_6532,N_5609,N_5536);
xnor U6533 (N_6533,N_5983,N_5360);
xor U6534 (N_6534,N_5476,N_5752);
nor U6535 (N_6535,N_5664,N_5436);
xor U6536 (N_6536,N_5764,N_5814);
nor U6537 (N_6537,N_5777,N_5824);
nor U6538 (N_6538,N_5304,N_5540);
nor U6539 (N_6539,N_5981,N_5844);
and U6540 (N_6540,N_5572,N_5452);
nor U6541 (N_6541,N_5282,N_5452);
nand U6542 (N_6542,N_5530,N_5807);
nand U6543 (N_6543,N_5562,N_5550);
or U6544 (N_6544,N_5589,N_5939);
nand U6545 (N_6545,N_5982,N_5675);
nand U6546 (N_6546,N_5542,N_5520);
and U6547 (N_6547,N_5368,N_5925);
nor U6548 (N_6548,N_5597,N_5467);
xor U6549 (N_6549,N_5477,N_5399);
or U6550 (N_6550,N_5724,N_5921);
nor U6551 (N_6551,N_5762,N_5351);
nor U6552 (N_6552,N_5559,N_5650);
and U6553 (N_6553,N_5922,N_5535);
xor U6554 (N_6554,N_5410,N_5851);
xnor U6555 (N_6555,N_5688,N_5958);
and U6556 (N_6556,N_5855,N_5363);
nor U6557 (N_6557,N_5520,N_5443);
nand U6558 (N_6558,N_5438,N_5422);
xor U6559 (N_6559,N_5280,N_5274);
or U6560 (N_6560,N_5746,N_5893);
nor U6561 (N_6561,N_5538,N_5778);
or U6562 (N_6562,N_5321,N_5731);
nor U6563 (N_6563,N_5482,N_5980);
and U6564 (N_6564,N_5772,N_5399);
and U6565 (N_6565,N_5411,N_5636);
nand U6566 (N_6566,N_5917,N_5859);
and U6567 (N_6567,N_5696,N_5265);
and U6568 (N_6568,N_5527,N_5327);
nor U6569 (N_6569,N_5962,N_5762);
xnor U6570 (N_6570,N_5775,N_5259);
nor U6571 (N_6571,N_5667,N_5524);
nor U6572 (N_6572,N_5390,N_5663);
xnor U6573 (N_6573,N_5253,N_5276);
xnor U6574 (N_6574,N_5467,N_5359);
nand U6575 (N_6575,N_5838,N_5856);
xnor U6576 (N_6576,N_5688,N_5562);
and U6577 (N_6577,N_5324,N_5602);
nor U6578 (N_6578,N_5488,N_5968);
or U6579 (N_6579,N_5425,N_5428);
or U6580 (N_6580,N_5513,N_5703);
xor U6581 (N_6581,N_5569,N_5933);
nor U6582 (N_6582,N_5324,N_5253);
or U6583 (N_6583,N_5378,N_5718);
nand U6584 (N_6584,N_5445,N_5708);
xnor U6585 (N_6585,N_5344,N_5293);
and U6586 (N_6586,N_5575,N_5598);
and U6587 (N_6587,N_5619,N_5408);
nand U6588 (N_6588,N_5344,N_5542);
nor U6589 (N_6589,N_5469,N_5962);
nand U6590 (N_6590,N_5810,N_5419);
and U6591 (N_6591,N_5506,N_5668);
xnor U6592 (N_6592,N_5509,N_5297);
and U6593 (N_6593,N_5535,N_5796);
xnor U6594 (N_6594,N_5331,N_5900);
nand U6595 (N_6595,N_5612,N_5264);
or U6596 (N_6596,N_5291,N_5883);
nor U6597 (N_6597,N_5870,N_5895);
or U6598 (N_6598,N_5323,N_5330);
xnor U6599 (N_6599,N_5724,N_5462);
and U6600 (N_6600,N_5561,N_5503);
nor U6601 (N_6601,N_5555,N_5883);
nand U6602 (N_6602,N_5909,N_5640);
or U6603 (N_6603,N_5952,N_5800);
and U6604 (N_6604,N_5406,N_5299);
nand U6605 (N_6605,N_5517,N_5542);
nand U6606 (N_6606,N_5527,N_5298);
nand U6607 (N_6607,N_5687,N_5581);
or U6608 (N_6608,N_5893,N_5261);
xor U6609 (N_6609,N_5459,N_5449);
xnor U6610 (N_6610,N_5925,N_5659);
xnor U6611 (N_6611,N_5386,N_5724);
or U6612 (N_6612,N_5421,N_5808);
or U6613 (N_6613,N_5421,N_5602);
and U6614 (N_6614,N_5522,N_5935);
nor U6615 (N_6615,N_5327,N_5539);
or U6616 (N_6616,N_5290,N_5288);
and U6617 (N_6617,N_5813,N_5373);
xor U6618 (N_6618,N_5638,N_5711);
and U6619 (N_6619,N_5329,N_5406);
xor U6620 (N_6620,N_5525,N_5741);
and U6621 (N_6621,N_5488,N_5601);
and U6622 (N_6622,N_5460,N_5873);
and U6623 (N_6623,N_5410,N_5380);
or U6624 (N_6624,N_5513,N_5573);
or U6625 (N_6625,N_5551,N_5665);
and U6626 (N_6626,N_5932,N_5826);
nand U6627 (N_6627,N_5860,N_5277);
xnor U6628 (N_6628,N_5621,N_5859);
or U6629 (N_6629,N_5482,N_5395);
or U6630 (N_6630,N_5828,N_5784);
or U6631 (N_6631,N_5883,N_5633);
or U6632 (N_6632,N_5605,N_5265);
or U6633 (N_6633,N_5252,N_5735);
and U6634 (N_6634,N_5583,N_5594);
xor U6635 (N_6635,N_5373,N_5281);
nand U6636 (N_6636,N_5334,N_5627);
nor U6637 (N_6637,N_5767,N_5376);
and U6638 (N_6638,N_5705,N_5526);
nor U6639 (N_6639,N_5699,N_5724);
xor U6640 (N_6640,N_5869,N_5331);
and U6641 (N_6641,N_5279,N_5749);
nor U6642 (N_6642,N_5895,N_5899);
xor U6643 (N_6643,N_5774,N_5498);
nand U6644 (N_6644,N_5714,N_5389);
xor U6645 (N_6645,N_5251,N_5920);
and U6646 (N_6646,N_5309,N_5421);
or U6647 (N_6647,N_5817,N_5878);
xor U6648 (N_6648,N_5775,N_5684);
nand U6649 (N_6649,N_5729,N_5568);
nor U6650 (N_6650,N_5554,N_5391);
and U6651 (N_6651,N_5638,N_5572);
nand U6652 (N_6652,N_5261,N_5784);
nor U6653 (N_6653,N_5285,N_5664);
nand U6654 (N_6654,N_5572,N_5295);
and U6655 (N_6655,N_5724,N_5888);
nor U6656 (N_6656,N_5494,N_5929);
or U6657 (N_6657,N_5569,N_5701);
xor U6658 (N_6658,N_5987,N_5572);
xnor U6659 (N_6659,N_5517,N_5479);
xor U6660 (N_6660,N_5713,N_5545);
nand U6661 (N_6661,N_5431,N_5962);
xor U6662 (N_6662,N_5615,N_5384);
and U6663 (N_6663,N_5278,N_5324);
nand U6664 (N_6664,N_5829,N_5358);
or U6665 (N_6665,N_5394,N_5963);
nand U6666 (N_6666,N_5373,N_5672);
nor U6667 (N_6667,N_5435,N_5355);
xnor U6668 (N_6668,N_5300,N_5602);
xor U6669 (N_6669,N_5705,N_5694);
or U6670 (N_6670,N_5312,N_5394);
xor U6671 (N_6671,N_5273,N_5752);
nand U6672 (N_6672,N_5905,N_5744);
or U6673 (N_6673,N_5559,N_5537);
nand U6674 (N_6674,N_5251,N_5429);
xnor U6675 (N_6675,N_5566,N_5989);
xor U6676 (N_6676,N_5855,N_5588);
nor U6677 (N_6677,N_5390,N_5551);
nand U6678 (N_6678,N_5739,N_5769);
nand U6679 (N_6679,N_5704,N_5463);
or U6680 (N_6680,N_5763,N_5546);
or U6681 (N_6681,N_5540,N_5826);
nor U6682 (N_6682,N_5629,N_5796);
nand U6683 (N_6683,N_5680,N_5959);
nand U6684 (N_6684,N_5888,N_5676);
or U6685 (N_6685,N_5964,N_5888);
nor U6686 (N_6686,N_5461,N_5404);
xor U6687 (N_6687,N_5306,N_5258);
xor U6688 (N_6688,N_5572,N_5947);
nand U6689 (N_6689,N_5605,N_5442);
xor U6690 (N_6690,N_5679,N_5323);
xnor U6691 (N_6691,N_5639,N_5975);
or U6692 (N_6692,N_5301,N_5459);
or U6693 (N_6693,N_5897,N_5496);
xor U6694 (N_6694,N_5607,N_5844);
xor U6695 (N_6695,N_5927,N_5393);
or U6696 (N_6696,N_5497,N_5615);
nor U6697 (N_6697,N_5286,N_5700);
xnor U6698 (N_6698,N_5981,N_5678);
xnor U6699 (N_6699,N_5552,N_5510);
nor U6700 (N_6700,N_5564,N_5437);
xnor U6701 (N_6701,N_5307,N_5725);
xnor U6702 (N_6702,N_5738,N_5355);
nand U6703 (N_6703,N_5332,N_5290);
or U6704 (N_6704,N_5374,N_5317);
and U6705 (N_6705,N_5746,N_5268);
nor U6706 (N_6706,N_5796,N_5997);
and U6707 (N_6707,N_5507,N_5705);
and U6708 (N_6708,N_5520,N_5722);
and U6709 (N_6709,N_5561,N_5932);
xor U6710 (N_6710,N_5761,N_5794);
nor U6711 (N_6711,N_5713,N_5528);
xor U6712 (N_6712,N_5278,N_5381);
and U6713 (N_6713,N_5770,N_5437);
nor U6714 (N_6714,N_5710,N_5527);
or U6715 (N_6715,N_5677,N_5918);
nand U6716 (N_6716,N_5556,N_5815);
nand U6717 (N_6717,N_5538,N_5621);
or U6718 (N_6718,N_5375,N_5725);
xor U6719 (N_6719,N_5719,N_5985);
nand U6720 (N_6720,N_5503,N_5504);
and U6721 (N_6721,N_5971,N_5747);
nand U6722 (N_6722,N_5454,N_5988);
xor U6723 (N_6723,N_5590,N_5333);
nor U6724 (N_6724,N_5325,N_5999);
and U6725 (N_6725,N_5285,N_5253);
xor U6726 (N_6726,N_5560,N_5426);
or U6727 (N_6727,N_5656,N_5463);
nand U6728 (N_6728,N_5750,N_5359);
and U6729 (N_6729,N_5552,N_5814);
nand U6730 (N_6730,N_5485,N_5277);
xor U6731 (N_6731,N_5615,N_5391);
nor U6732 (N_6732,N_5439,N_5772);
xnor U6733 (N_6733,N_5878,N_5407);
and U6734 (N_6734,N_5642,N_5668);
nand U6735 (N_6735,N_5745,N_5765);
and U6736 (N_6736,N_5563,N_5793);
and U6737 (N_6737,N_5577,N_5393);
nand U6738 (N_6738,N_5543,N_5650);
xor U6739 (N_6739,N_5561,N_5796);
xor U6740 (N_6740,N_5614,N_5586);
nand U6741 (N_6741,N_5446,N_5263);
xor U6742 (N_6742,N_5651,N_5471);
nor U6743 (N_6743,N_5737,N_5948);
or U6744 (N_6744,N_5739,N_5831);
xnor U6745 (N_6745,N_5291,N_5919);
or U6746 (N_6746,N_5679,N_5850);
and U6747 (N_6747,N_5605,N_5481);
or U6748 (N_6748,N_5305,N_5308);
nand U6749 (N_6749,N_5258,N_5738);
xnor U6750 (N_6750,N_6449,N_6090);
nor U6751 (N_6751,N_6218,N_6233);
xor U6752 (N_6752,N_6248,N_6683);
or U6753 (N_6753,N_6058,N_6190);
nor U6754 (N_6754,N_6268,N_6083);
xnor U6755 (N_6755,N_6521,N_6575);
nand U6756 (N_6756,N_6510,N_6681);
nor U6757 (N_6757,N_6003,N_6250);
or U6758 (N_6758,N_6089,N_6165);
and U6759 (N_6759,N_6118,N_6104);
nand U6760 (N_6760,N_6106,N_6001);
nor U6761 (N_6761,N_6359,N_6548);
and U6762 (N_6762,N_6467,N_6578);
xnor U6763 (N_6763,N_6205,N_6701);
nand U6764 (N_6764,N_6581,N_6245);
xnor U6765 (N_6765,N_6124,N_6039);
nor U6766 (N_6766,N_6673,N_6518);
xnor U6767 (N_6767,N_6476,N_6226);
nor U6768 (N_6768,N_6473,N_6225);
nor U6769 (N_6769,N_6685,N_6399);
nand U6770 (N_6770,N_6224,N_6554);
nor U6771 (N_6771,N_6046,N_6731);
nor U6772 (N_6772,N_6597,N_6735);
and U6773 (N_6773,N_6532,N_6588);
nand U6774 (N_6774,N_6453,N_6197);
and U6775 (N_6775,N_6024,N_6527);
or U6776 (N_6776,N_6624,N_6331);
and U6777 (N_6777,N_6401,N_6499);
or U6778 (N_6778,N_6481,N_6659);
xnor U6779 (N_6779,N_6494,N_6227);
nor U6780 (N_6780,N_6706,N_6274);
nand U6781 (N_6781,N_6035,N_6145);
nand U6782 (N_6782,N_6488,N_6458);
xnor U6783 (N_6783,N_6194,N_6468);
xor U6784 (N_6784,N_6579,N_6219);
and U6785 (N_6785,N_6451,N_6123);
xnor U6786 (N_6786,N_6541,N_6516);
nand U6787 (N_6787,N_6114,N_6170);
or U6788 (N_6788,N_6444,N_6350);
xnor U6789 (N_6789,N_6718,N_6018);
nor U6790 (N_6790,N_6013,N_6695);
nor U6791 (N_6791,N_6049,N_6103);
or U6792 (N_6792,N_6610,N_6356);
or U6793 (N_6793,N_6639,N_6668);
nand U6794 (N_6794,N_6726,N_6280);
nor U6795 (N_6795,N_6709,N_6590);
and U6796 (N_6796,N_6383,N_6071);
xnor U6797 (N_6797,N_6396,N_6121);
and U6798 (N_6798,N_6625,N_6747);
and U6799 (N_6799,N_6189,N_6550);
nand U6800 (N_6800,N_6415,N_6580);
nor U6801 (N_6801,N_6295,N_6495);
and U6802 (N_6802,N_6077,N_6178);
nor U6803 (N_6803,N_6098,N_6043);
nand U6804 (N_6804,N_6207,N_6397);
and U6805 (N_6805,N_6725,N_6109);
and U6806 (N_6806,N_6287,N_6710);
and U6807 (N_6807,N_6559,N_6188);
or U6808 (N_6808,N_6220,N_6424);
xnor U6809 (N_6809,N_6199,N_6093);
or U6810 (N_6810,N_6445,N_6158);
or U6811 (N_6811,N_6347,N_6513);
and U6812 (N_6812,N_6727,N_6688);
nand U6813 (N_6813,N_6493,N_6169);
and U6814 (N_6814,N_6557,N_6479);
nor U6815 (N_6815,N_6708,N_6616);
xor U6816 (N_6816,N_6334,N_6368);
and U6817 (N_6817,N_6247,N_6583);
or U6818 (N_6818,N_6357,N_6386);
or U6819 (N_6819,N_6021,N_6714);
xor U6820 (N_6820,N_6587,N_6120);
or U6821 (N_6821,N_6582,N_6733);
nor U6822 (N_6822,N_6029,N_6129);
nand U6823 (N_6823,N_6429,N_6661);
or U6824 (N_6824,N_6407,N_6348);
or U6825 (N_6825,N_6705,N_6414);
or U6826 (N_6826,N_6064,N_6540);
and U6827 (N_6827,N_6384,N_6455);
xor U6828 (N_6828,N_6471,N_6151);
xor U6829 (N_6829,N_6674,N_6627);
or U6830 (N_6830,N_6477,N_6128);
xnor U6831 (N_6831,N_6440,N_6028);
nor U6832 (N_6832,N_6671,N_6275);
nand U6833 (N_6833,N_6149,N_6339);
xor U6834 (N_6834,N_6343,N_6044);
xor U6835 (N_6835,N_6056,N_6305);
xor U6836 (N_6836,N_6208,N_6301);
and U6837 (N_6837,N_6351,N_6643);
xnor U6838 (N_6838,N_6652,N_6378);
nor U6839 (N_6839,N_6241,N_6641);
or U6840 (N_6840,N_6312,N_6594);
nor U6841 (N_6841,N_6341,N_6690);
xor U6842 (N_6842,N_6100,N_6411);
and U6843 (N_6843,N_6257,N_6080);
nor U6844 (N_6844,N_6537,N_6655);
or U6845 (N_6845,N_6460,N_6298);
and U6846 (N_6846,N_6577,N_6484);
xnor U6847 (N_6847,N_6657,N_6108);
or U6848 (N_6848,N_6586,N_6558);
or U6849 (N_6849,N_6605,N_6536);
nor U6850 (N_6850,N_6125,N_6620);
nand U6851 (N_6851,N_6722,N_6006);
and U6852 (N_6852,N_6418,N_6526);
and U6853 (N_6853,N_6677,N_6382);
nand U6854 (N_6854,N_6117,N_6525);
or U6855 (N_6855,N_6078,N_6094);
xor U6856 (N_6856,N_6087,N_6408);
xor U6857 (N_6857,N_6571,N_6387);
nor U6858 (N_6858,N_6309,N_6565);
or U6859 (N_6859,N_6353,N_6167);
or U6860 (N_6860,N_6395,N_6676);
nand U6861 (N_6861,N_6215,N_6463);
and U6862 (N_6862,N_6004,N_6279);
nand U6863 (N_6863,N_6036,N_6329);
nor U6864 (N_6864,N_6156,N_6574);
and U6865 (N_6865,N_6293,N_6107);
xor U6866 (N_6866,N_6232,N_6263);
or U6867 (N_6867,N_6719,N_6288);
xnor U6868 (N_6868,N_6475,N_6569);
nand U6869 (N_6869,N_6622,N_6011);
xor U6870 (N_6870,N_6512,N_6133);
nor U6871 (N_6871,N_6642,N_6336);
xnor U6872 (N_6872,N_6529,N_6713);
nand U6873 (N_6873,N_6323,N_6490);
xor U6874 (N_6874,N_6134,N_6530);
or U6875 (N_6875,N_6195,N_6127);
or U6876 (N_6876,N_6730,N_6648);
or U6877 (N_6877,N_6313,N_6697);
or U6878 (N_6878,N_6181,N_6744);
xor U6879 (N_6879,N_6228,N_6647);
nand U6880 (N_6880,N_6054,N_6084);
xnor U6881 (N_6881,N_6073,N_6509);
and U6882 (N_6882,N_6180,N_6609);
and U6883 (N_6883,N_6556,N_6693);
or U6884 (N_6884,N_6212,N_6566);
or U6885 (N_6885,N_6691,N_6503);
nor U6886 (N_6886,N_6079,N_6159);
nor U6887 (N_6887,N_6342,N_6322);
xor U6888 (N_6888,N_6522,N_6636);
and U6889 (N_6889,N_6489,N_6626);
and U6890 (N_6890,N_6294,N_6326);
and U6891 (N_6891,N_6187,N_6173);
xor U6892 (N_6892,N_6560,N_6286);
nand U6893 (N_6893,N_6254,N_6454);
or U6894 (N_6894,N_6113,N_6604);
nand U6895 (N_6895,N_6650,N_6016);
nand U6896 (N_6896,N_6026,N_6613);
or U6897 (N_6897,N_6595,N_6086);
or U6898 (N_6898,N_6060,N_6632);
or U6899 (N_6899,N_6355,N_6171);
and U6900 (N_6900,N_6014,N_6373);
xor U6901 (N_6901,N_6439,N_6174);
and U6902 (N_6902,N_6282,N_6672);
xor U6903 (N_6903,N_6211,N_6221);
nor U6904 (N_6904,N_6122,N_6005);
and U6905 (N_6905,N_6161,N_6349);
and U6906 (N_6906,N_6296,N_6692);
nand U6907 (N_6907,N_6419,N_6277);
nand U6908 (N_6908,N_6664,N_6095);
or U6909 (N_6909,N_6130,N_6551);
nor U6910 (N_6910,N_6185,N_6409);
nor U6911 (N_6911,N_6404,N_6164);
or U6912 (N_6912,N_6059,N_6539);
nor U6913 (N_6913,N_6748,N_6135);
nor U6914 (N_6914,N_6362,N_6564);
nand U6915 (N_6915,N_6266,N_6278);
and U6916 (N_6916,N_6191,N_6593);
nor U6917 (N_6917,N_6370,N_6491);
xnor U6918 (N_6918,N_6741,N_6700);
or U6919 (N_6919,N_6160,N_6289);
and U6920 (N_6920,N_6737,N_6315);
nand U6921 (N_6921,N_6447,N_6327);
and U6922 (N_6922,N_6022,N_6423);
xor U6923 (N_6923,N_6469,N_6470);
nand U6924 (N_6924,N_6738,N_6547);
nand U6925 (N_6925,N_6517,N_6267);
or U6926 (N_6926,N_6328,N_6291);
and U6927 (N_6927,N_6679,N_6506);
nor U6928 (N_6928,N_6111,N_6363);
and U6929 (N_6929,N_6507,N_6192);
and U6930 (N_6930,N_6137,N_6466);
xor U6931 (N_6931,N_6237,N_6658);
xor U6932 (N_6932,N_6482,N_6146);
and U6933 (N_6933,N_6153,N_6422);
or U6934 (N_6934,N_6544,N_6391);
nand U6935 (N_6935,N_6175,N_6502);
nor U6936 (N_6936,N_6033,N_6410);
nand U6937 (N_6937,N_6459,N_6320);
nor U6938 (N_6938,N_6591,N_6306);
nor U6939 (N_6939,N_6038,N_6635);
and U6940 (N_6940,N_6150,N_6702);
or U6941 (N_6941,N_6061,N_6088);
nor U6942 (N_6942,N_6157,N_6523);
nor U6943 (N_6943,N_6740,N_6400);
or U6944 (N_6944,N_6416,N_6015);
nor U6945 (N_6945,N_6143,N_6155);
nand U6946 (N_6946,N_6040,N_6736);
and U6947 (N_6947,N_6222,N_6682);
and U6948 (N_6948,N_6621,N_6303);
xor U6949 (N_6949,N_6649,N_6075);
or U6950 (N_6950,N_6520,N_6390);
xor U6951 (N_6951,N_6567,N_6456);
nor U6952 (N_6952,N_6229,N_6589);
nand U6953 (N_6953,N_6256,N_6009);
or U6954 (N_6954,N_6426,N_6235);
or U6955 (N_6955,N_6265,N_6317);
xor U6956 (N_6956,N_6182,N_6533);
nor U6957 (N_6957,N_6485,N_6728);
or U6958 (N_6958,N_6048,N_6515);
xnor U6959 (N_6959,N_6501,N_6433);
or U6960 (N_6960,N_6606,N_6213);
and U6961 (N_6961,N_6644,N_6542);
xor U6962 (N_6962,N_6394,N_6438);
nand U6963 (N_6963,N_6253,N_6596);
xor U6964 (N_6964,N_6615,N_6259);
nor U6965 (N_6965,N_6119,N_6608);
xnor U6966 (N_6966,N_6217,N_6202);
xor U6967 (N_6967,N_6549,N_6629);
or U6968 (N_6968,N_6371,N_6645);
xnor U6969 (N_6969,N_6201,N_6214);
xor U6970 (N_6970,N_6176,N_6264);
nand U6971 (N_6971,N_6154,N_6545);
nor U6972 (N_6972,N_6553,N_6742);
nor U6973 (N_6973,N_6561,N_6050);
nor U6974 (N_6974,N_6552,N_6534);
nor U6975 (N_6975,N_6101,N_6019);
and U6976 (N_6976,N_6734,N_6462);
and U6977 (N_6977,N_6074,N_6319);
or U6978 (N_6978,N_6576,N_6746);
nand U6979 (N_6979,N_6234,N_6498);
nand U6980 (N_6980,N_6538,N_6297);
xor U6981 (N_6981,N_6066,N_6242);
and U6982 (N_6982,N_6115,N_6251);
nor U6983 (N_6983,N_6500,N_6562);
xnor U6984 (N_6984,N_6206,N_6599);
and U6985 (N_6985,N_6346,N_6179);
xnor U6986 (N_6986,N_6375,N_6030);
and U6987 (N_6987,N_6099,N_6653);
nor U6988 (N_6988,N_6745,N_6421);
nor U6989 (N_6989,N_6186,N_6318);
nand U6990 (N_6990,N_6435,N_6132);
nand U6991 (N_6991,N_6619,N_6209);
nand U6992 (N_6992,N_6689,N_6367);
nand U6993 (N_6993,N_6360,N_6743);
or U6994 (N_6994,N_6299,N_6252);
xnor U6995 (N_6995,N_6258,N_6112);
nor U6996 (N_6996,N_6662,N_6721);
nor U6997 (N_6997,N_6568,N_6666);
or U6998 (N_6998,N_6448,N_6302);
nand U6999 (N_6999,N_6210,N_6330);
xnor U7000 (N_7000,N_6017,N_6430);
and U7001 (N_7001,N_6425,N_6678);
and U7002 (N_7002,N_6139,N_6405);
or U7003 (N_7003,N_6651,N_6497);
nand U7004 (N_7004,N_6193,N_6260);
xnor U7005 (N_7005,N_6531,N_6524);
nand U7006 (N_7006,N_6634,N_6603);
xnor U7007 (N_7007,N_6045,N_6204);
xor U7008 (N_7008,N_6380,N_6474);
or U7009 (N_7009,N_6105,N_6618);
xor U7010 (N_7010,N_6203,N_6116);
or U7011 (N_7011,N_6344,N_6273);
xnor U7012 (N_7012,N_6431,N_6374);
or U7013 (N_7013,N_6249,N_6398);
and U7014 (N_7014,N_6031,N_6729);
xnor U7015 (N_7015,N_6446,N_6010);
or U7016 (N_7016,N_6667,N_6163);
and U7017 (N_7017,N_6707,N_6262);
and U7018 (N_7018,N_6441,N_6670);
nand U7019 (N_7019,N_6640,N_6126);
xor U7020 (N_7020,N_6572,N_6168);
nand U7021 (N_7021,N_6376,N_6081);
and U7022 (N_7022,N_6023,N_6366);
and U7023 (N_7023,N_6177,N_6053);
xor U7024 (N_7024,N_6669,N_6085);
nand U7025 (N_7025,N_6570,N_6261);
nand U7026 (N_7026,N_6680,N_6592);
and U7027 (N_7027,N_6442,N_6243);
nor U7028 (N_7028,N_6340,N_6246);
xnor U7029 (N_7029,N_6236,N_6352);
nand U7030 (N_7030,N_6230,N_6543);
nand U7031 (N_7031,N_6285,N_6717);
nand U7032 (N_7032,N_6281,N_6183);
nor U7033 (N_7033,N_6147,N_6598);
and U7034 (N_7034,N_6712,N_6388);
or U7035 (N_7035,N_6141,N_6427);
nor U7036 (N_7036,N_6076,N_6244);
nor U7037 (N_7037,N_6223,N_6068);
or U7038 (N_7038,N_6654,N_6412);
nor U7039 (N_7039,N_6720,N_6434);
nand U7040 (N_7040,N_6051,N_6631);
and U7041 (N_7041,N_6699,N_6162);
xor U7042 (N_7042,N_6486,N_6063);
or U7043 (N_7043,N_6369,N_6239);
and U7044 (N_7044,N_6216,N_6337);
and U7045 (N_7045,N_6437,N_6292);
nand U7046 (N_7046,N_6514,N_6097);
or U7047 (N_7047,N_6240,N_6623);
nor U7048 (N_7048,N_6276,N_6614);
or U7049 (N_7049,N_6505,N_6008);
nand U7050 (N_7050,N_6546,N_6308);
and U7051 (N_7051,N_6283,N_6316);
nand U7052 (N_7052,N_6660,N_6696);
and U7053 (N_7053,N_6361,N_6102);
and U7054 (N_7054,N_6496,N_6110);
and U7055 (N_7055,N_6612,N_6304);
nand U7056 (N_7056,N_6508,N_6034);
nor U7057 (N_7057,N_6739,N_6480);
or U7058 (N_7058,N_6602,N_6062);
xnor U7059 (N_7059,N_6172,N_6617);
nor U7060 (N_7060,N_6002,N_6335);
or U7061 (N_7061,N_6403,N_6472);
xor U7062 (N_7062,N_6140,N_6300);
and U7063 (N_7063,N_6646,N_6633);
or U7064 (N_7064,N_6535,N_6715);
nand U7065 (N_7065,N_6067,N_6184);
xnor U7066 (N_7066,N_6096,N_6724);
or U7067 (N_7067,N_6354,N_6377);
nand U7068 (N_7068,N_6684,N_6381);
xor U7069 (N_7069,N_6457,N_6432);
xnor U7070 (N_7070,N_6487,N_6321);
xor U7071 (N_7071,N_6255,N_6231);
or U7072 (N_7072,N_6511,N_6042);
xnor U7073 (N_7073,N_6152,N_6379);
and U7074 (N_7074,N_6032,N_6392);
and U7075 (N_7075,N_6136,N_6436);
or U7076 (N_7076,N_6492,N_6464);
or U7077 (N_7077,N_6365,N_6338);
xor U7078 (N_7078,N_6314,N_6333);
nand U7079 (N_7079,N_6325,N_6465);
and U7080 (N_7080,N_6057,N_6082);
nor U7081 (N_7081,N_6238,N_6389);
nor U7082 (N_7082,N_6041,N_6012);
xnor U7083 (N_7083,N_6025,N_6638);
or U7084 (N_7084,N_6372,N_6732);
nand U7085 (N_7085,N_6271,N_6047);
and U7086 (N_7086,N_6364,N_6284);
xor U7087 (N_7087,N_6450,N_6611);
xnor U7088 (N_7088,N_6663,N_6332);
and U7089 (N_7089,N_6142,N_6417);
and U7090 (N_7090,N_6483,N_6452);
and U7091 (N_7091,N_6072,N_6665);
nor U7092 (N_7092,N_6393,N_6148);
or U7093 (N_7093,N_6420,N_6461);
or U7094 (N_7094,N_6065,N_6091);
nand U7095 (N_7095,N_6675,N_6601);
or U7096 (N_7096,N_6052,N_6694);
nand U7097 (N_7097,N_6385,N_6528);
xor U7098 (N_7098,N_6749,N_6584);
or U7099 (N_7099,N_6563,N_6131);
or U7100 (N_7100,N_6272,N_6585);
and U7101 (N_7101,N_6716,N_6310);
and U7102 (N_7102,N_6628,N_6200);
and U7103 (N_7103,N_6711,N_6607);
and U7104 (N_7104,N_6270,N_6704);
xnor U7105 (N_7105,N_6345,N_6723);
and U7106 (N_7106,N_6703,N_6196);
nand U7107 (N_7107,N_6027,N_6656);
and U7108 (N_7108,N_6070,N_6600);
xnor U7109 (N_7109,N_6144,N_6358);
nand U7110 (N_7110,N_6324,N_6698);
and U7111 (N_7111,N_6007,N_6687);
or U7112 (N_7112,N_6519,N_6269);
or U7113 (N_7113,N_6307,N_6637);
nand U7114 (N_7114,N_6555,N_6478);
nand U7115 (N_7115,N_6020,N_6428);
nor U7116 (N_7116,N_6630,N_6092);
xor U7117 (N_7117,N_6166,N_6406);
or U7118 (N_7118,N_6686,N_6413);
and U7119 (N_7119,N_6443,N_6198);
nor U7120 (N_7120,N_6069,N_6573);
nand U7121 (N_7121,N_6138,N_6402);
or U7122 (N_7122,N_6290,N_6037);
and U7123 (N_7123,N_6504,N_6311);
or U7124 (N_7124,N_6000,N_6055);
nand U7125 (N_7125,N_6372,N_6518);
nor U7126 (N_7126,N_6516,N_6089);
and U7127 (N_7127,N_6150,N_6322);
or U7128 (N_7128,N_6009,N_6021);
or U7129 (N_7129,N_6059,N_6250);
nor U7130 (N_7130,N_6118,N_6232);
or U7131 (N_7131,N_6086,N_6587);
nor U7132 (N_7132,N_6283,N_6254);
nand U7133 (N_7133,N_6065,N_6602);
or U7134 (N_7134,N_6352,N_6295);
nand U7135 (N_7135,N_6161,N_6521);
xor U7136 (N_7136,N_6524,N_6397);
and U7137 (N_7137,N_6418,N_6259);
or U7138 (N_7138,N_6620,N_6401);
nor U7139 (N_7139,N_6086,N_6057);
nor U7140 (N_7140,N_6355,N_6341);
nand U7141 (N_7141,N_6726,N_6417);
xnor U7142 (N_7142,N_6468,N_6230);
nor U7143 (N_7143,N_6254,N_6679);
or U7144 (N_7144,N_6414,N_6279);
nor U7145 (N_7145,N_6221,N_6490);
and U7146 (N_7146,N_6650,N_6210);
or U7147 (N_7147,N_6167,N_6122);
nor U7148 (N_7148,N_6184,N_6375);
nor U7149 (N_7149,N_6087,N_6509);
and U7150 (N_7150,N_6197,N_6341);
xor U7151 (N_7151,N_6399,N_6628);
and U7152 (N_7152,N_6358,N_6452);
xor U7153 (N_7153,N_6341,N_6538);
or U7154 (N_7154,N_6372,N_6678);
and U7155 (N_7155,N_6407,N_6103);
xnor U7156 (N_7156,N_6500,N_6481);
or U7157 (N_7157,N_6037,N_6166);
or U7158 (N_7158,N_6466,N_6651);
nand U7159 (N_7159,N_6275,N_6481);
or U7160 (N_7160,N_6175,N_6090);
or U7161 (N_7161,N_6315,N_6045);
and U7162 (N_7162,N_6492,N_6735);
and U7163 (N_7163,N_6571,N_6711);
nand U7164 (N_7164,N_6436,N_6279);
nor U7165 (N_7165,N_6591,N_6294);
nand U7166 (N_7166,N_6220,N_6135);
nor U7167 (N_7167,N_6383,N_6284);
nand U7168 (N_7168,N_6068,N_6003);
or U7169 (N_7169,N_6660,N_6608);
nor U7170 (N_7170,N_6015,N_6013);
or U7171 (N_7171,N_6385,N_6218);
and U7172 (N_7172,N_6247,N_6347);
nand U7173 (N_7173,N_6743,N_6711);
xnor U7174 (N_7174,N_6384,N_6374);
and U7175 (N_7175,N_6304,N_6268);
xor U7176 (N_7176,N_6632,N_6254);
nor U7177 (N_7177,N_6578,N_6133);
and U7178 (N_7178,N_6161,N_6360);
nor U7179 (N_7179,N_6296,N_6465);
xnor U7180 (N_7180,N_6601,N_6747);
nand U7181 (N_7181,N_6227,N_6045);
nand U7182 (N_7182,N_6032,N_6552);
or U7183 (N_7183,N_6016,N_6389);
nor U7184 (N_7184,N_6529,N_6376);
and U7185 (N_7185,N_6022,N_6675);
and U7186 (N_7186,N_6723,N_6176);
and U7187 (N_7187,N_6036,N_6037);
and U7188 (N_7188,N_6362,N_6226);
or U7189 (N_7189,N_6183,N_6659);
and U7190 (N_7190,N_6675,N_6511);
xor U7191 (N_7191,N_6703,N_6168);
and U7192 (N_7192,N_6702,N_6499);
nor U7193 (N_7193,N_6618,N_6184);
nand U7194 (N_7194,N_6206,N_6294);
nand U7195 (N_7195,N_6577,N_6613);
or U7196 (N_7196,N_6510,N_6132);
or U7197 (N_7197,N_6140,N_6039);
or U7198 (N_7198,N_6049,N_6260);
xnor U7199 (N_7199,N_6270,N_6245);
or U7200 (N_7200,N_6059,N_6709);
nor U7201 (N_7201,N_6152,N_6409);
nand U7202 (N_7202,N_6069,N_6603);
or U7203 (N_7203,N_6239,N_6541);
or U7204 (N_7204,N_6469,N_6081);
nand U7205 (N_7205,N_6098,N_6702);
xor U7206 (N_7206,N_6003,N_6019);
xnor U7207 (N_7207,N_6517,N_6075);
nand U7208 (N_7208,N_6155,N_6598);
nor U7209 (N_7209,N_6056,N_6627);
xnor U7210 (N_7210,N_6083,N_6384);
nor U7211 (N_7211,N_6492,N_6336);
and U7212 (N_7212,N_6457,N_6675);
nor U7213 (N_7213,N_6444,N_6573);
nor U7214 (N_7214,N_6134,N_6497);
xor U7215 (N_7215,N_6685,N_6447);
or U7216 (N_7216,N_6263,N_6282);
xor U7217 (N_7217,N_6437,N_6679);
nand U7218 (N_7218,N_6173,N_6079);
nor U7219 (N_7219,N_6060,N_6363);
nor U7220 (N_7220,N_6596,N_6437);
and U7221 (N_7221,N_6674,N_6626);
nor U7222 (N_7222,N_6148,N_6088);
nor U7223 (N_7223,N_6049,N_6550);
nor U7224 (N_7224,N_6115,N_6663);
xnor U7225 (N_7225,N_6403,N_6658);
and U7226 (N_7226,N_6444,N_6428);
nor U7227 (N_7227,N_6407,N_6437);
and U7228 (N_7228,N_6427,N_6228);
xnor U7229 (N_7229,N_6033,N_6459);
and U7230 (N_7230,N_6530,N_6235);
and U7231 (N_7231,N_6126,N_6283);
or U7232 (N_7232,N_6536,N_6294);
nor U7233 (N_7233,N_6591,N_6244);
and U7234 (N_7234,N_6385,N_6008);
nor U7235 (N_7235,N_6186,N_6732);
or U7236 (N_7236,N_6247,N_6373);
nand U7237 (N_7237,N_6506,N_6507);
or U7238 (N_7238,N_6683,N_6579);
or U7239 (N_7239,N_6186,N_6523);
or U7240 (N_7240,N_6665,N_6702);
or U7241 (N_7241,N_6434,N_6308);
or U7242 (N_7242,N_6642,N_6288);
nand U7243 (N_7243,N_6524,N_6313);
and U7244 (N_7244,N_6153,N_6264);
nand U7245 (N_7245,N_6387,N_6421);
nand U7246 (N_7246,N_6219,N_6636);
nor U7247 (N_7247,N_6222,N_6476);
and U7248 (N_7248,N_6422,N_6543);
nor U7249 (N_7249,N_6439,N_6243);
xor U7250 (N_7250,N_6228,N_6015);
xor U7251 (N_7251,N_6218,N_6424);
and U7252 (N_7252,N_6448,N_6211);
xor U7253 (N_7253,N_6295,N_6729);
nand U7254 (N_7254,N_6032,N_6257);
nand U7255 (N_7255,N_6136,N_6611);
nor U7256 (N_7256,N_6105,N_6737);
xnor U7257 (N_7257,N_6517,N_6068);
xnor U7258 (N_7258,N_6744,N_6021);
nand U7259 (N_7259,N_6457,N_6290);
xnor U7260 (N_7260,N_6152,N_6727);
nand U7261 (N_7261,N_6703,N_6513);
nand U7262 (N_7262,N_6263,N_6630);
xor U7263 (N_7263,N_6104,N_6727);
and U7264 (N_7264,N_6690,N_6479);
nor U7265 (N_7265,N_6455,N_6626);
nor U7266 (N_7266,N_6051,N_6047);
nand U7267 (N_7267,N_6294,N_6619);
nand U7268 (N_7268,N_6319,N_6046);
nor U7269 (N_7269,N_6187,N_6201);
nor U7270 (N_7270,N_6716,N_6030);
and U7271 (N_7271,N_6252,N_6672);
xor U7272 (N_7272,N_6196,N_6722);
or U7273 (N_7273,N_6545,N_6230);
nor U7274 (N_7274,N_6053,N_6615);
nand U7275 (N_7275,N_6665,N_6736);
nor U7276 (N_7276,N_6386,N_6413);
nand U7277 (N_7277,N_6186,N_6224);
nand U7278 (N_7278,N_6062,N_6490);
nor U7279 (N_7279,N_6580,N_6257);
or U7280 (N_7280,N_6089,N_6159);
and U7281 (N_7281,N_6201,N_6603);
and U7282 (N_7282,N_6393,N_6000);
xor U7283 (N_7283,N_6617,N_6283);
nor U7284 (N_7284,N_6722,N_6375);
xor U7285 (N_7285,N_6710,N_6715);
nand U7286 (N_7286,N_6010,N_6558);
nor U7287 (N_7287,N_6650,N_6451);
nor U7288 (N_7288,N_6032,N_6551);
or U7289 (N_7289,N_6316,N_6473);
nand U7290 (N_7290,N_6139,N_6343);
nor U7291 (N_7291,N_6647,N_6112);
nor U7292 (N_7292,N_6546,N_6021);
and U7293 (N_7293,N_6352,N_6658);
xnor U7294 (N_7294,N_6302,N_6693);
or U7295 (N_7295,N_6637,N_6448);
xor U7296 (N_7296,N_6276,N_6392);
or U7297 (N_7297,N_6118,N_6510);
or U7298 (N_7298,N_6237,N_6082);
nand U7299 (N_7299,N_6635,N_6400);
nor U7300 (N_7300,N_6338,N_6631);
or U7301 (N_7301,N_6667,N_6644);
nand U7302 (N_7302,N_6458,N_6437);
nand U7303 (N_7303,N_6423,N_6067);
or U7304 (N_7304,N_6138,N_6407);
or U7305 (N_7305,N_6186,N_6389);
and U7306 (N_7306,N_6739,N_6208);
or U7307 (N_7307,N_6363,N_6397);
or U7308 (N_7308,N_6177,N_6117);
nand U7309 (N_7309,N_6168,N_6096);
nand U7310 (N_7310,N_6559,N_6088);
or U7311 (N_7311,N_6638,N_6697);
xnor U7312 (N_7312,N_6070,N_6569);
nand U7313 (N_7313,N_6057,N_6378);
nor U7314 (N_7314,N_6365,N_6103);
and U7315 (N_7315,N_6544,N_6705);
nand U7316 (N_7316,N_6703,N_6069);
and U7317 (N_7317,N_6586,N_6683);
xnor U7318 (N_7318,N_6606,N_6180);
nand U7319 (N_7319,N_6055,N_6664);
nor U7320 (N_7320,N_6643,N_6035);
xor U7321 (N_7321,N_6351,N_6141);
and U7322 (N_7322,N_6143,N_6058);
nor U7323 (N_7323,N_6395,N_6495);
nand U7324 (N_7324,N_6471,N_6239);
and U7325 (N_7325,N_6577,N_6184);
xnor U7326 (N_7326,N_6030,N_6491);
nand U7327 (N_7327,N_6568,N_6251);
nor U7328 (N_7328,N_6692,N_6339);
and U7329 (N_7329,N_6435,N_6243);
and U7330 (N_7330,N_6734,N_6618);
xor U7331 (N_7331,N_6024,N_6126);
nand U7332 (N_7332,N_6146,N_6651);
and U7333 (N_7333,N_6450,N_6358);
xnor U7334 (N_7334,N_6608,N_6360);
nand U7335 (N_7335,N_6739,N_6721);
nor U7336 (N_7336,N_6183,N_6094);
nand U7337 (N_7337,N_6199,N_6243);
or U7338 (N_7338,N_6587,N_6545);
xnor U7339 (N_7339,N_6188,N_6083);
nand U7340 (N_7340,N_6470,N_6000);
xor U7341 (N_7341,N_6153,N_6120);
nand U7342 (N_7342,N_6407,N_6629);
xnor U7343 (N_7343,N_6083,N_6607);
or U7344 (N_7344,N_6748,N_6531);
nand U7345 (N_7345,N_6642,N_6542);
xor U7346 (N_7346,N_6498,N_6157);
nor U7347 (N_7347,N_6729,N_6434);
or U7348 (N_7348,N_6466,N_6547);
xor U7349 (N_7349,N_6243,N_6598);
nand U7350 (N_7350,N_6543,N_6130);
xor U7351 (N_7351,N_6705,N_6312);
or U7352 (N_7352,N_6662,N_6466);
xnor U7353 (N_7353,N_6643,N_6592);
nand U7354 (N_7354,N_6215,N_6656);
or U7355 (N_7355,N_6647,N_6543);
nor U7356 (N_7356,N_6290,N_6623);
nor U7357 (N_7357,N_6496,N_6436);
and U7358 (N_7358,N_6687,N_6348);
nand U7359 (N_7359,N_6297,N_6674);
nor U7360 (N_7360,N_6535,N_6139);
nor U7361 (N_7361,N_6217,N_6712);
nand U7362 (N_7362,N_6474,N_6340);
or U7363 (N_7363,N_6488,N_6725);
xor U7364 (N_7364,N_6304,N_6683);
or U7365 (N_7365,N_6054,N_6722);
or U7366 (N_7366,N_6051,N_6129);
nand U7367 (N_7367,N_6642,N_6340);
and U7368 (N_7368,N_6677,N_6701);
nand U7369 (N_7369,N_6058,N_6250);
nand U7370 (N_7370,N_6681,N_6580);
xnor U7371 (N_7371,N_6589,N_6056);
xnor U7372 (N_7372,N_6500,N_6166);
or U7373 (N_7373,N_6355,N_6672);
nor U7374 (N_7374,N_6722,N_6167);
nor U7375 (N_7375,N_6252,N_6274);
nand U7376 (N_7376,N_6203,N_6332);
nand U7377 (N_7377,N_6497,N_6184);
and U7378 (N_7378,N_6504,N_6107);
and U7379 (N_7379,N_6101,N_6295);
xor U7380 (N_7380,N_6651,N_6653);
nand U7381 (N_7381,N_6048,N_6554);
xnor U7382 (N_7382,N_6714,N_6669);
xnor U7383 (N_7383,N_6296,N_6178);
or U7384 (N_7384,N_6533,N_6459);
xor U7385 (N_7385,N_6090,N_6083);
nand U7386 (N_7386,N_6180,N_6434);
nor U7387 (N_7387,N_6111,N_6096);
nor U7388 (N_7388,N_6030,N_6455);
and U7389 (N_7389,N_6458,N_6312);
or U7390 (N_7390,N_6344,N_6010);
nor U7391 (N_7391,N_6350,N_6178);
or U7392 (N_7392,N_6504,N_6486);
xnor U7393 (N_7393,N_6455,N_6289);
and U7394 (N_7394,N_6029,N_6182);
or U7395 (N_7395,N_6176,N_6307);
nor U7396 (N_7396,N_6594,N_6458);
nor U7397 (N_7397,N_6330,N_6451);
and U7398 (N_7398,N_6684,N_6594);
and U7399 (N_7399,N_6404,N_6648);
xnor U7400 (N_7400,N_6286,N_6596);
nor U7401 (N_7401,N_6396,N_6137);
xnor U7402 (N_7402,N_6014,N_6601);
nand U7403 (N_7403,N_6457,N_6047);
or U7404 (N_7404,N_6353,N_6269);
and U7405 (N_7405,N_6233,N_6121);
xnor U7406 (N_7406,N_6226,N_6725);
nor U7407 (N_7407,N_6576,N_6060);
nor U7408 (N_7408,N_6723,N_6560);
xnor U7409 (N_7409,N_6517,N_6580);
nand U7410 (N_7410,N_6362,N_6092);
nand U7411 (N_7411,N_6420,N_6210);
and U7412 (N_7412,N_6260,N_6353);
nor U7413 (N_7413,N_6007,N_6270);
and U7414 (N_7414,N_6269,N_6239);
xnor U7415 (N_7415,N_6051,N_6353);
nand U7416 (N_7416,N_6368,N_6543);
or U7417 (N_7417,N_6079,N_6528);
xnor U7418 (N_7418,N_6003,N_6385);
and U7419 (N_7419,N_6648,N_6693);
or U7420 (N_7420,N_6621,N_6339);
nor U7421 (N_7421,N_6633,N_6448);
nor U7422 (N_7422,N_6457,N_6487);
nand U7423 (N_7423,N_6297,N_6399);
nand U7424 (N_7424,N_6390,N_6700);
nand U7425 (N_7425,N_6141,N_6650);
and U7426 (N_7426,N_6440,N_6233);
nor U7427 (N_7427,N_6018,N_6574);
and U7428 (N_7428,N_6428,N_6731);
and U7429 (N_7429,N_6656,N_6629);
and U7430 (N_7430,N_6708,N_6291);
and U7431 (N_7431,N_6042,N_6551);
xnor U7432 (N_7432,N_6559,N_6268);
and U7433 (N_7433,N_6025,N_6651);
or U7434 (N_7434,N_6585,N_6075);
nand U7435 (N_7435,N_6183,N_6112);
or U7436 (N_7436,N_6524,N_6462);
xnor U7437 (N_7437,N_6063,N_6120);
and U7438 (N_7438,N_6458,N_6166);
nor U7439 (N_7439,N_6586,N_6287);
xnor U7440 (N_7440,N_6392,N_6474);
and U7441 (N_7441,N_6337,N_6033);
nand U7442 (N_7442,N_6120,N_6699);
xor U7443 (N_7443,N_6193,N_6042);
xor U7444 (N_7444,N_6169,N_6162);
or U7445 (N_7445,N_6675,N_6179);
xor U7446 (N_7446,N_6281,N_6720);
and U7447 (N_7447,N_6593,N_6573);
nand U7448 (N_7448,N_6207,N_6244);
or U7449 (N_7449,N_6067,N_6655);
xnor U7450 (N_7450,N_6352,N_6587);
xor U7451 (N_7451,N_6251,N_6058);
or U7452 (N_7452,N_6345,N_6144);
nand U7453 (N_7453,N_6053,N_6376);
nand U7454 (N_7454,N_6118,N_6381);
and U7455 (N_7455,N_6435,N_6280);
and U7456 (N_7456,N_6074,N_6470);
or U7457 (N_7457,N_6547,N_6032);
or U7458 (N_7458,N_6198,N_6317);
nand U7459 (N_7459,N_6156,N_6666);
and U7460 (N_7460,N_6384,N_6166);
and U7461 (N_7461,N_6245,N_6062);
nand U7462 (N_7462,N_6381,N_6457);
or U7463 (N_7463,N_6626,N_6483);
nand U7464 (N_7464,N_6321,N_6219);
xnor U7465 (N_7465,N_6220,N_6262);
nor U7466 (N_7466,N_6531,N_6259);
or U7467 (N_7467,N_6724,N_6017);
nand U7468 (N_7468,N_6234,N_6572);
nand U7469 (N_7469,N_6518,N_6180);
and U7470 (N_7470,N_6360,N_6419);
nand U7471 (N_7471,N_6311,N_6730);
or U7472 (N_7472,N_6201,N_6152);
nor U7473 (N_7473,N_6292,N_6398);
or U7474 (N_7474,N_6315,N_6674);
and U7475 (N_7475,N_6190,N_6542);
xor U7476 (N_7476,N_6414,N_6399);
nor U7477 (N_7477,N_6520,N_6304);
xor U7478 (N_7478,N_6427,N_6269);
and U7479 (N_7479,N_6564,N_6336);
or U7480 (N_7480,N_6209,N_6361);
or U7481 (N_7481,N_6383,N_6539);
or U7482 (N_7482,N_6452,N_6229);
or U7483 (N_7483,N_6413,N_6677);
xnor U7484 (N_7484,N_6283,N_6729);
xor U7485 (N_7485,N_6446,N_6502);
xor U7486 (N_7486,N_6077,N_6008);
xor U7487 (N_7487,N_6289,N_6138);
or U7488 (N_7488,N_6334,N_6070);
and U7489 (N_7489,N_6709,N_6422);
or U7490 (N_7490,N_6683,N_6619);
nand U7491 (N_7491,N_6729,N_6136);
nand U7492 (N_7492,N_6539,N_6516);
nor U7493 (N_7493,N_6711,N_6491);
xor U7494 (N_7494,N_6218,N_6055);
or U7495 (N_7495,N_6632,N_6406);
or U7496 (N_7496,N_6530,N_6430);
xnor U7497 (N_7497,N_6299,N_6151);
xnor U7498 (N_7498,N_6639,N_6228);
xnor U7499 (N_7499,N_6395,N_6274);
xor U7500 (N_7500,N_7234,N_6783);
or U7501 (N_7501,N_7349,N_6831);
xor U7502 (N_7502,N_6968,N_6973);
nand U7503 (N_7503,N_7355,N_6914);
and U7504 (N_7504,N_6789,N_7160);
nand U7505 (N_7505,N_7258,N_7126);
nand U7506 (N_7506,N_6998,N_6787);
nor U7507 (N_7507,N_7291,N_7076);
or U7508 (N_7508,N_7282,N_7351);
and U7509 (N_7509,N_7147,N_6900);
nor U7510 (N_7510,N_6989,N_6902);
xor U7511 (N_7511,N_7273,N_7064);
or U7512 (N_7512,N_6921,N_7209);
nor U7513 (N_7513,N_7012,N_6993);
nor U7514 (N_7514,N_7132,N_7178);
nand U7515 (N_7515,N_6962,N_6959);
nor U7516 (N_7516,N_6799,N_7109);
nor U7517 (N_7517,N_7242,N_7368);
xor U7518 (N_7518,N_6843,N_6837);
or U7519 (N_7519,N_7146,N_6961);
and U7520 (N_7520,N_6956,N_7302);
or U7521 (N_7521,N_7155,N_7461);
nor U7522 (N_7522,N_7432,N_6826);
xnor U7523 (N_7523,N_7344,N_7374);
nand U7524 (N_7524,N_7231,N_7100);
or U7525 (N_7525,N_7085,N_7218);
xor U7526 (N_7526,N_6770,N_6964);
and U7527 (N_7527,N_7340,N_7304);
nand U7528 (N_7528,N_6990,N_7263);
nor U7529 (N_7529,N_6876,N_6920);
xor U7530 (N_7530,N_7407,N_7277);
and U7531 (N_7531,N_6965,N_6909);
nand U7532 (N_7532,N_7393,N_6946);
or U7533 (N_7533,N_7294,N_6923);
nand U7534 (N_7534,N_7203,N_7055);
xor U7535 (N_7535,N_7071,N_7322);
nor U7536 (N_7536,N_6814,N_7091);
nor U7537 (N_7537,N_6986,N_7397);
nor U7538 (N_7538,N_6769,N_6980);
nor U7539 (N_7539,N_6791,N_7281);
nor U7540 (N_7540,N_7078,N_7326);
and U7541 (N_7541,N_6917,N_7303);
xnor U7542 (N_7542,N_7066,N_7089);
or U7543 (N_7543,N_6856,N_7013);
nor U7544 (N_7544,N_7020,N_7140);
nand U7545 (N_7545,N_7454,N_7062);
xor U7546 (N_7546,N_6882,N_7241);
nand U7547 (N_7547,N_6774,N_7093);
xor U7548 (N_7548,N_7321,N_7341);
and U7549 (N_7549,N_7310,N_7348);
and U7550 (N_7550,N_7269,N_7034);
or U7551 (N_7551,N_7206,N_7058);
xor U7552 (N_7552,N_6889,N_7193);
nor U7553 (N_7553,N_7312,N_7365);
nor U7554 (N_7554,N_7042,N_6981);
and U7555 (N_7555,N_7196,N_7026);
or U7556 (N_7556,N_7445,N_6807);
xnor U7557 (N_7557,N_7223,N_6940);
nand U7558 (N_7558,N_7039,N_7446);
xor U7559 (N_7559,N_6937,N_7080);
and U7560 (N_7560,N_7198,N_6978);
and U7561 (N_7561,N_7429,N_7334);
xor U7562 (N_7562,N_7005,N_6879);
nand U7563 (N_7563,N_7128,N_7017);
and U7564 (N_7564,N_7179,N_7157);
and U7565 (N_7565,N_6844,N_6898);
nor U7566 (N_7566,N_7450,N_7376);
nand U7567 (N_7567,N_7127,N_7171);
nand U7568 (N_7568,N_7214,N_7098);
nor U7569 (N_7569,N_7219,N_7243);
and U7570 (N_7570,N_6951,N_7447);
and U7571 (N_7571,N_7136,N_6872);
and U7572 (N_7572,N_7029,N_7475);
or U7573 (N_7573,N_6975,N_6773);
nor U7574 (N_7574,N_7370,N_7133);
nor U7575 (N_7575,N_6772,N_7107);
xor U7576 (N_7576,N_6829,N_7489);
nand U7577 (N_7577,N_6835,N_7087);
and U7578 (N_7578,N_7083,N_7197);
and U7579 (N_7579,N_6750,N_6913);
and U7580 (N_7580,N_7435,N_6796);
xnor U7581 (N_7581,N_7460,N_7194);
and U7582 (N_7582,N_7498,N_7410);
or U7583 (N_7583,N_7164,N_7471);
nand U7584 (N_7584,N_6929,N_6958);
or U7585 (N_7585,N_6931,N_7396);
or U7586 (N_7586,N_7323,N_7182);
and U7587 (N_7587,N_6957,N_6926);
and U7588 (N_7588,N_7215,N_6764);
nor U7589 (N_7589,N_7297,N_7459);
nor U7590 (N_7590,N_7324,N_7168);
nor U7591 (N_7591,N_7217,N_7059);
or U7592 (N_7592,N_7079,N_7189);
nand U7593 (N_7593,N_7047,N_6869);
nor U7594 (N_7594,N_6955,N_6935);
or U7595 (N_7595,N_7329,N_6974);
and U7596 (N_7596,N_7077,N_7254);
nor U7597 (N_7597,N_7262,N_7307);
nor U7598 (N_7598,N_7375,N_7249);
or U7599 (N_7599,N_6776,N_6997);
and U7600 (N_7600,N_7113,N_6820);
or U7601 (N_7601,N_6943,N_6852);
and U7602 (N_7602,N_6782,N_7339);
and U7603 (N_7603,N_6758,N_7050);
xor U7604 (N_7604,N_6918,N_7406);
nor U7605 (N_7605,N_7296,N_7444);
and U7606 (N_7606,N_6803,N_7224);
xor U7607 (N_7607,N_7068,N_6751);
or U7608 (N_7608,N_7252,N_7208);
nor U7609 (N_7609,N_7442,N_7280);
nand U7610 (N_7610,N_7037,N_7118);
nand U7611 (N_7611,N_6806,N_7373);
and U7612 (N_7612,N_7007,N_7283);
nor U7613 (N_7613,N_6985,N_7449);
and U7614 (N_7614,N_7404,N_7465);
xor U7615 (N_7615,N_6868,N_7130);
or U7616 (N_7616,N_6878,N_6757);
or U7617 (N_7617,N_7401,N_7385);
nand U7618 (N_7618,N_7038,N_7416);
nor U7619 (N_7619,N_7371,N_6819);
nor U7620 (N_7620,N_7388,N_7092);
nor U7621 (N_7621,N_7046,N_7412);
nand U7622 (N_7622,N_7463,N_6939);
xnor U7623 (N_7623,N_6983,N_7239);
nor U7624 (N_7624,N_7285,N_7353);
or U7625 (N_7625,N_6862,N_7073);
or U7626 (N_7626,N_7377,N_7305);
nor U7627 (N_7627,N_6895,N_6960);
nor U7628 (N_7628,N_7448,N_7279);
nor U7629 (N_7629,N_6833,N_7210);
and U7630 (N_7630,N_7174,N_7230);
nand U7631 (N_7631,N_7086,N_7065);
or U7632 (N_7632,N_7161,N_7261);
nand U7633 (N_7633,N_7021,N_6984);
nand U7634 (N_7634,N_7473,N_6930);
nor U7635 (N_7635,N_7030,N_6786);
nand U7636 (N_7636,N_6875,N_7169);
nor U7637 (N_7637,N_7335,N_6848);
or U7638 (N_7638,N_7120,N_7163);
and U7639 (N_7639,N_7331,N_7006);
xnor U7640 (N_7640,N_7337,N_6827);
xor U7641 (N_7641,N_7137,N_7286);
or U7642 (N_7642,N_6849,N_7345);
nor U7643 (N_7643,N_7325,N_7199);
and U7644 (N_7644,N_7248,N_6987);
or U7645 (N_7645,N_7056,N_7306);
xnor U7646 (N_7646,N_7316,N_6775);
nand U7647 (N_7647,N_6952,N_6867);
xnor U7648 (N_7648,N_7457,N_7019);
and U7649 (N_7649,N_6892,N_7229);
nand U7650 (N_7650,N_7255,N_7278);
nor U7651 (N_7651,N_6780,N_7496);
nor U7652 (N_7652,N_7419,N_7499);
and U7653 (N_7653,N_6784,N_7008);
nor U7654 (N_7654,N_7400,N_6756);
nand U7655 (N_7655,N_6795,N_6907);
and U7656 (N_7656,N_6860,N_6881);
xnor U7657 (N_7657,N_7170,N_7270);
xnor U7658 (N_7658,N_6953,N_7200);
or U7659 (N_7659,N_6847,N_6912);
xor U7660 (N_7660,N_7380,N_6821);
nor U7661 (N_7661,N_7367,N_7315);
and U7662 (N_7662,N_7403,N_6877);
and U7663 (N_7663,N_7011,N_6880);
and U7664 (N_7664,N_7390,N_7320);
nand U7665 (N_7665,N_7096,N_7060);
or U7666 (N_7666,N_6781,N_6950);
nand U7667 (N_7667,N_6967,N_7010);
nand U7668 (N_7668,N_6841,N_7453);
xnor U7669 (N_7669,N_7481,N_7031);
nand U7670 (N_7670,N_7265,N_7186);
nand U7671 (N_7671,N_7480,N_7221);
and U7672 (N_7672,N_7434,N_6753);
nand U7673 (N_7673,N_7359,N_7028);
and U7674 (N_7674,N_6846,N_6948);
or U7675 (N_7675,N_7384,N_7094);
xnor U7676 (N_7676,N_6808,N_7417);
nand U7677 (N_7677,N_7382,N_7222);
nor U7678 (N_7678,N_7486,N_7308);
xnor U7679 (N_7679,N_7418,N_6905);
nor U7680 (N_7680,N_7441,N_7158);
nand U7681 (N_7681,N_7119,N_7167);
xor U7682 (N_7682,N_7328,N_7350);
nor U7683 (N_7683,N_6768,N_7057);
or U7684 (N_7684,N_7378,N_7421);
xor U7685 (N_7685,N_7386,N_6911);
and U7686 (N_7686,N_7183,N_7069);
or U7687 (N_7687,N_7491,N_7338);
nand U7688 (N_7688,N_6766,N_7451);
nand U7689 (N_7689,N_6798,N_6863);
and U7690 (N_7690,N_7260,N_6949);
nand U7691 (N_7691,N_7228,N_6971);
nor U7692 (N_7692,N_7372,N_6793);
nand U7693 (N_7693,N_7000,N_7099);
xor U7694 (N_7694,N_6828,N_7275);
nor U7695 (N_7695,N_6797,N_6976);
or U7696 (N_7696,N_6865,N_6840);
nand U7697 (N_7697,N_6922,N_7129);
nor U7698 (N_7698,N_7131,N_7470);
or U7699 (N_7699,N_7485,N_7356);
xor U7700 (N_7700,N_6830,N_6979);
and U7701 (N_7701,N_7138,N_7268);
nand U7702 (N_7702,N_7436,N_7456);
nor U7703 (N_7703,N_7154,N_7300);
or U7704 (N_7704,N_7488,N_6904);
xnor U7705 (N_7705,N_6812,N_7327);
or U7706 (N_7706,N_7121,N_7469);
nand U7707 (N_7707,N_7088,N_7188);
nor U7708 (N_7708,N_6761,N_7181);
or U7709 (N_7709,N_7479,N_7317);
nor U7710 (N_7710,N_7298,N_7438);
or U7711 (N_7711,N_6896,N_7225);
or U7712 (N_7712,N_6901,N_6916);
nand U7713 (N_7713,N_6836,N_6947);
or U7714 (N_7714,N_7431,N_7244);
xnor U7715 (N_7715,N_6899,N_6825);
xnor U7716 (N_7716,N_7187,N_6972);
xor U7717 (N_7717,N_7259,N_6815);
nand U7718 (N_7718,N_7141,N_7311);
and U7719 (N_7719,N_6924,N_7398);
nand U7720 (N_7720,N_7052,N_7105);
xnor U7721 (N_7721,N_6897,N_7016);
and U7722 (N_7722,N_7004,N_7430);
xnor U7723 (N_7723,N_7180,N_6982);
xnor U7724 (N_7724,N_7114,N_7101);
nor U7725 (N_7725,N_7212,N_6887);
or U7726 (N_7726,N_6938,N_7392);
or U7727 (N_7727,N_6858,N_7240);
nor U7728 (N_7728,N_7264,N_7112);
xnor U7729 (N_7729,N_7455,N_6928);
nor U7730 (N_7730,N_7097,N_7414);
or U7731 (N_7731,N_6888,N_6919);
nor U7732 (N_7732,N_7207,N_7483);
nor U7733 (N_7733,N_7405,N_7074);
nor U7734 (N_7734,N_6861,N_6908);
xnor U7735 (N_7735,N_6942,N_7015);
nand U7736 (N_7736,N_7271,N_7415);
and U7737 (N_7737,N_7108,N_7428);
nand U7738 (N_7738,N_6870,N_7025);
nand U7739 (N_7739,N_6866,N_7205);
or U7740 (N_7740,N_7072,N_7408);
xnor U7741 (N_7741,N_6785,N_7149);
nor U7742 (N_7742,N_7246,N_7361);
xnor U7743 (N_7743,N_6755,N_7202);
and U7744 (N_7744,N_6915,N_7123);
xnor U7745 (N_7745,N_7266,N_6765);
nor U7746 (N_7746,N_7357,N_6963);
and U7747 (N_7747,N_7102,N_6816);
and U7748 (N_7748,N_6894,N_7022);
or U7749 (N_7749,N_6969,N_6954);
and U7750 (N_7750,N_7095,N_7233);
and U7751 (N_7751,N_7173,N_7220);
nand U7752 (N_7752,N_7413,N_7067);
nor U7753 (N_7753,N_7314,N_7043);
nand U7754 (N_7754,N_7145,N_6855);
xor U7755 (N_7755,N_6767,N_6805);
or U7756 (N_7756,N_7175,N_6991);
xnor U7757 (N_7757,N_7362,N_7125);
and U7758 (N_7758,N_6792,N_7290);
or U7759 (N_7759,N_6934,N_7216);
xor U7760 (N_7760,N_7443,N_6891);
nand U7761 (N_7761,N_7497,N_6811);
nor U7762 (N_7762,N_7150,N_7153);
and U7763 (N_7763,N_7192,N_7110);
xor U7764 (N_7764,N_6910,N_6996);
and U7765 (N_7765,N_6801,N_7389);
xnor U7766 (N_7766,N_6977,N_7292);
and U7767 (N_7767,N_7477,N_6800);
or U7768 (N_7768,N_7383,N_6871);
and U7769 (N_7769,N_7176,N_7253);
and U7770 (N_7770,N_7476,N_7295);
or U7771 (N_7771,N_7256,N_7204);
nor U7772 (N_7772,N_7053,N_7054);
and U7773 (N_7773,N_7166,N_6762);
and U7774 (N_7774,N_7287,N_7422);
or U7775 (N_7775,N_7284,N_6763);
nand U7776 (N_7776,N_7104,N_7232);
or U7777 (N_7777,N_7184,N_7274);
or U7778 (N_7778,N_7162,N_7117);
or U7779 (N_7779,N_6817,N_7075);
nand U7780 (N_7780,N_6992,N_7381);
or U7781 (N_7781,N_7009,N_7342);
nand U7782 (N_7782,N_7464,N_7023);
or U7783 (N_7783,N_7152,N_7044);
nand U7784 (N_7784,N_7041,N_7245);
nor U7785 (N_7785,N_7051,N_6851);
or U7786 (N_7786,N_7111,N_7411);
xnor U7787 (N_7787,N_7213,N_7135);
nand U7788 (N_7788,N_7366,N_7048);
xor U7789 (N_7789,N_7492,N_7084);
nor U7790 (N_7790,N_7346,N_7301);
xnor U7791 (N_7791,N_6794,N_7336);
and U7792 (N_7792,N_7201,N_7035);
xor U7793 (N_7793,N_7433,N_7251);
xor U7794 (N_7794,N_7276,N_7495);
xnor U7795 (N_7795,N_7364,N_6834);
or U7796 (N_7796,N_7474,N_7144);
or U7797 (N_7797,N_7352,N_7379);
or U7798 (N_7798,N_6839,N_6813);
or U7799 (N_7799,N_7437,N_7330);
nand U7800 (N_7800,N_7402,N_6809);
xor U7801 (N_7801,N_7103,N_7309);
xnor U7802 (N_7802,N_6760,N_7190);
nand U7803 (N_7803,N_6788,N_6838);
nor U7804 (N_7804,N_6864,N_6771);
nand U7805 (N_7805,N_7002,N_6927);
or U7806 (N_7806,N_7358,N_7090);
nand U7807 (N_7807,N_6857,N_7116);
nand U7808 (N_7808,N_7409,N_6854);
or U7809 (N_7809,N_7003,N_7354);
or U7810 (N_7810,N_7293,N_7333);
nor U7811 (N_7811,N_6884,N_7177);
or U7812 (N_7812,N_7458,N_6886);
nor U7813 (N_7813,N_7484,N_6883);
nand U7814 (N_7814,N_6941,N_7142);
or U7815 (N_7815,N_6999,N_6754);
xor U7816 (N_7816,N_6778,N_7440);
nand U7817 (N_7817,N_6804,N_7018);
nand U7818 (N_7818,N_7387,N_7238);
xor U7819 (N_7819,N_7399,N_7363);
xnor U7820 (N_7820,N_7045,N_7143);
xnor U7821 (N_7821,N_6845,N_7395);
nor U7822 (N_7822,N_6874,N_7425);
and U7823 (N_7823,N_7001,N_7360);
and U7824 (N_7824,N_6818,N_6906);
and U7825 (N_7825,N_7493,N_7250);
nor U7826 (N_7826,N_7332,N_6823);
and U7827 (N_7827,N_7426,N_7288);
nor U7828 (N_7828,N_7191,N_6759);
or U7829 (N_7829,N_7227,N_7134);
nand U7830 (N_7830,N_7462,N_7427);
and U7831 (N_7831,N_6873,N_7313);
or U7832 (N_7832,N_7257,N_7472);
nor U7833 (N_7833,N_7369,N_6994);
xor U7834 (N_7834,N_7343,N_6925);
nor U7835 (N_7835,N_7151,N_6850);
nor U7836 (N_7836,N_7319,N_6859);
nand U7837 (N_7837,N_7478,N_7049);
xnor U7838 (N_7838,N_7272,N_7036);
xnor U7839 (N_7839,N_6936,N_7211);
nor U7840 (N_7840,N_7027,N_6970);
nand U7841 (N_7841,N_6822,N_6988);
nor U7842 (N_7842,N_7156,N_7139);
nor U7843 (N_7843,N_6790,N_7237);
xnor U7844 (N_7844,N_7247,N_7494);
xnor U7845 (N_7845,N_7172,N_7423);
nand U7846 (N_7846,N_7148,N_7040);
or U7847 (N_7847,N_7490,N_6777);
xor U7848 (N_7848,N_6824,N_7487);
nor U7849 (N_7849,N_7394,N_6966);
nor U7850 (N_7850,N_6945,N_6903);
and U7851 (N_7851,N_7014,N_7482);
or U7852 (N_7852,N_7424,N_7115);
nand U7853 (N_7853,N_6752,N_6779);
xnor U7854 (N_7854,N_6810,N_7391);
nand U7855 (N_7855,N_6832,N_7032);
or U7856 (N_7856,N_7081,N_7024);
xnor U7857 (N_7857,N_6933,N_7124);
xnor U7858 (N_7858,N_7420,N_7318);
or U7859 (N_7859,N_7122,N_7347);
nor U7860 (N_7860,N_7061,N_7165);
nand U7861 (N_7861,N_7466,N_7033);
or U7862 (N_7862,N_6893,N_7185);
or U7863 (N_7863,N_6995,N_6944);
nor U7864 (N_7864,N_6802,N_7468);
xnor U7865 (N_7865,N_6885,N_7267);
nor U7866 (N_7866,N_7289,N_7467);
and U7867 (N_7867,N_7063,N_6853);
or U7868 (N_7868,N_7452,N_7236);
nor U7869 (N_7869,N_7235,N_7106);
and U7870 (N_7870,N_7082,N_6932);
and U7871 (N_7871,N_7299,N_7195);
nor U7872 (N_7872,N_7226,N_7439);
nor U7873 (N_7873,N_7159,N_6842);
nand U7874 (N_7874,N_7070,N_6890);
or U7875 (N_7875,N_6921,N_7231);
nor U7876 (N_7876,N_6919,N_7196);
xor U7877 (N_7877,N_6930,N_7344);
nor U7878 (N_7878,N_7112,N_7487);
nand U7879 (N_7879,N_7286,N_7425);
and U7880 (N_7880,N_7436,N_7216);
or U7881 (N_7881,N_6784,N_6980);
or U7882 (N_7882,N_6940,N_6783);
nor U7883 (N_7883,N_7048,N_7176);
nand U7884 (N_7884,N_7002,N_7155);
xor U7885 (N_7885,N_6976,N_7061);
nor U7886 (N_7886,N_7489,N_7353);
nand U7887 (N_7887,N_7353,N_7022);
or U7888 (N_7888,N_7173,N_6948);
nand U7889 (N_7889,N_7188,N_6788);
nor U7890 (N_7890,N_7434,N_7378);
nand U7891 (N_7891,N_6771,N_7085);
or U7892 (N_7892,N_6771,N_7220);
or U7893 (N_7893,N_7395,N_6788);
or U7894 (N_7894,N_6796,N_6871);
nand U7895 (N_7895,N_7420,N_6852);
or U7896 (N_7896,N_7344,N_7019);
xnor U7897 (N_7897,N_6840,N_7371);
nor U7898 (N_7898,N_7044,N_7164);
nand U7899 (N_7899,N_7028,N_6776);
xnor U7900 (N_7900,N_7145,N_7442);
nand U7901 (N_7901,N_7160,N_7295);
nor U7902 (N_7902,N_6888,N_7178);
xor U7903 (N_7903,N_7103,N_7272);
and U7904 (N_7904,N_6779,N_7155);
nand U7905 (N_7905,N_7193,N_7225);
xor U7906 (N_7906,N_7253,N_7138);
or U7907 (N_7907,N_7175,N_7315);
nor U7908 (N_7908,N_6917,N_6754);
or U7909 (N_7909,N_7421,N_6971);
xor U7910 (N_7910,N_7378,N_7352);
xnor U7911 (N_7911,N_7107,N_7239);
and U7912 (N_7912,N_6910,N_7034);
nor U7913 (N_7913,N_6820,N_7265);
or U7914 (N_7914,N_6783,N_6935);
and U7915 (N_7915,N_7463,N_7272);
xor U7916 (N_7916,N_6815,N_6792);
nand U7917 (N_7917,N_7181,N_7089);
nor U7918 (N_7918,N_6873,N_7444);
nor U7919 (N_7919,N_7422,N_7275);
xor U7920 (N_7920,N_7286,N_7014);
and U7921 (N_7921,N_7010,N_6959);
xor U7922 (N_7922,N_7232,N_7475);
nand U7923 (N_7923,N_7021,N_6943);
xnor U7924 (N_7924,N_7433,N_6903);
nand U7925 (N_7925,N_7472,N_6983);
or U7926 (N_7926,N_7116,N_7002);
and U7927 (N_7927,N_7123,N_7180);
xor U7928 (N_7928,N_7160,N_6856);
xnor U7929 (N_7929,N_7132,N_6867);
nand U7930 (N_7930,N_7122,N_6753);
or U7931 (N_7931,N_6903,N_7260);
nor U7932 (N_7932,N_7120,N_7151);
or U7933 (N_7933,N_7209,N_7170);
nor U7934 (N_7934,N_7256,N_6823);
xor U7935 (N_7935,N_7463,N_7392);
nor U7936 (N_7936,N_7169,N_6964);
nand U7937 (N_7937,N_6863,N_6817);
xor U7938 (N_7938,N_7090,N_7351);
xnor U7939 (N_7939,N_7193,N_7276);
nand U7940 (N_7940,N_6997,N_6768);
xor U7941 (N_7941,N_6803,N_7154);
nand U7942 (N_7942,N_7336,N_6925);
xor U7943 (N_7943,N_7431,N_6855);
and U7944 (N_7944,N_7098,N_7436);
nand U7945 (N_7945,N_7408,N_6938);
nor U7946 (N_7946,N_6798,N_7240);
and U7947 (N_7947,N_7282,N_7349);
xnor U7948 (N_7948,N_7268,N_7179);
xor U7949 (N_7949,N_6976,N_7280);
and U7950 (N_7950,N_7315,N_6823);
nand U7951 (N_7951,N_6896,N_7426);
and U7952 (N_7952,N_6766,N_6810);
xor U7953 (N_7953,N_7286,N_7485);
xnor U7954 (N_7954,N_6960,N_7498);
and U7955 (N_7955,N_7099,N_6876);
nor U7956 (N_7956,N_7392,N_6907);
xor U7957 (N_7957,N_6772,N_7132);
nand U7958 (N_7958,N_7360,N_7111);
nor U7959 (N_7959,N_7292,N_6758);
xnor U7960 (N_7960,N_7490,N_7067);
nand U7961 (N_7961,N_6935,N_7483);
xor U7962 (N_7962,N_6903,N_7249);
or U7963 (N_7963,N_7439,N_6879);
nand U7964 (N_7964,N_7391,N_7046);
nand U7965 (N_7965,N_6777,N_7054);
and U7966 (N_7966,N_7197,N_7105);
xor U7967 (N_7967,N_7296,N_7004);
nor U7968 (N_7968,N_7403,N_7272);
xnor U7969 (N_7969,N_7305,N_6837);
nand U7970 (N_7970,N_7080,N_7434);
nor U7971 (N_7971,N_7371,N_6936);
nand U7972 (N_7972,N_7254,N_6857);
or U7973 (N_7973,N_6890,N_6966);
nand U7974 (N_7974,N_6851,N_6991);
nor U7975 (N_7975,N_7325,N_6822);
xor U7976 (N_7976,N_7176,N_6934);
nor U7977 (N_7977,N_7341,N_7297);
xor U7978 (N_7978,N_7231,N_7134);
xnor U7979 (N_7979,N_7335,N_6909);
or U7980 (N_7980,N_7495,N_6813);
xnor U7981 (N_7981,N_6839,N_6946);
nor U7982 (N_7982,N_7079,N_7016);
or U7983 (N_7983,N_7479,N_7496);
nand U7984 (N_7984,N_7328,N_7063);
nand U7985 (N_7985,N_6959,N_7137);
nand U7986 (N_7986,N_6809,N_6980);
nand U7987 (N_7987,N_6924,N_6930);
and U7988 (N_7988,N_7457,N_7231);
nand U7989 (N_7989,N_7239,N_7317);
nor U7990 (N_7990,N_6948,N_7258);
nor U7991 (N_7991,N_7063,N_7175);
nor U7992 (N_7992,N_7449,N_6762);
and U7993 (N_7993,N_7031,N_7389);
or U7994 (N_7994,N_7399,N_6854);
nor U7995 (N_7995,N_7147,N_7208);
or U7996 (N_7996,N_7135,N_7229);
nand U7997 (N_7997,N_7165,N_6930);
xor U7998 (N_7998,N_6850,N_6795);
nor U7999 (N_7999,N_6757,N_6824);
nor U8000 (N_8000,N_7127,N_6875);
nand U8001 (N_8001,N_6955,N_6864);
xnor U8002 (N_8002,N_6790,N_6920);
and U8003 (N_8003,N_6797,N_6805);
nand U8004 (N_8004,N_7249,N_7150);
and U8005 (N_8005,N_6852,N_7235);
or U8006 (N_8006,N_7023,N_7321);
or U8007 (N_8007,N_7298,N_7129);
and U8008 (N_8008,N_7493,N_7390);
nor U8009 (N_8009,N_7328,N_6765);
or U8010 (N_8010,N_6785,N_7120);
and U8011 (N_8011,N_6869,N_7315);
or U8012 (N_8012,N_7431,N_7062);
xnor U8013 (N_8013,N_7056,N_6823);
or U8014 (N_8014,N_7080,N_7453);
nor U8015 (N_8015,N_7055,N_7069);
or U8016 (N_8016,N_7005,N_7225);
nor U8017 (N_8017,N_7467,N_6778);
or U8018 (N_8018,N_7209,N_7314);
or U8019 (N_8019,N_7352,N_6823);
xor U8020 (N_8020,N_7271,N_6984);
nor U8021 (N_8021,N_7031,N_6803);
or U8022 (N_8022,N_6872,N_6895);
xor U8023 (N_8023,N_7387,N_6916);
and U8024 (N_8024,N_7190,N_7253);
nor U8025 (N_8025,N_7015,N_6778);
nand U8026 (N_8026,N_7394,N_7328);
nand U8027 (N_8027,N_7333,N_7453);
nand U8028 (N_8028,N_7119,N_6774);
nand U8029 (N_8029,N_7408,N_7360);
xor U8030 (N_8030,N_7210,N_6980);
nor U8031 (N_8031,N_6940,N_7483);
or U8032 (N_8032,N_7303,N_7310);
or U8033 (N_8033,N_7434,N_6852);
xor U8034 (N_8034,N_7265,N_7015);
and U8035 (N_8035,N_7304,N_7057);
and U8036 (N_8036,N_7399,N_6753);
nor U8037 (N_8037,N_7306,N_7051);
and U8038 (N_8038,N_6905,N_7183);
xnor U8039 (N_8039,N_7187,N_7186);
xor U8040 (N_8040,N_6924,N_7435);
nand U8041 (N_8041,N_6775,N_7084);
xor U8042 (N_8042,N_7298,N_7110);
or U8043 (N_8043,N_6984,N_7034);
nand U8044 (N_8044,N_7330,N_7395);
nor U8045 (N_8045,N_6994,N_7180);
or U8046 (N_8046,N_6786,N_7117);
and U8047 (N_8047,N_7144,N_7058);
xnor U8048 (N_8048,N_7345,N_7472);
and U8049 (N_8049,N_6813,N_7123);
xnor U8050 (N_8050,N_7193,N_7443);
or U8051 (N_8051,N_6914,N_7320);
xnor U8052 (N_8052,N_6920,N_7158);
and U8053 (N_8053,N_7405,N_7048);
nor U8054 (N_8054,N_7365,N_7448);
nand U8055 (N_8055,N_6922,N_6964);
and U8056 (N_8056,N_7031,N_7081);
or U8057 (N_8057,N_7234,N_7209);
or U8058 (N_8058,N_6821,N_7426);
nand U8059 (N_8059,N_7072,N_7446);
nand U8060 (N_8060,N_6834,N_6773);
or U8061 (N_8061,N_7113,N_6765);
or U8062 (N_8062,N_7344,N_6759);
nor U8063 (N_8063,N_7414,N_7188);
nor U8064 (N_8064,N_6781,N_6817);
nor U8065 (N_8065,N_7225,N_6946);
and U8066 (N_8066,N_7027,N_7094);
xnor U8067 (N_8067,N_7165,N_7125);
or U8068 (N_8068,N_6799,N_7036);
and U8069 (N_8069,N_7000,N_7179);
nor U8070 (N_8070,N_7107,N_7461);
and U8071 (N_8071,N_7381,N_7457);
nor U8072 (N_8072,N_6871,N_7476);
xnor U8073 (N_8073,N_7177,N_7358);
nor U8074 (N_8074,N_6933,N_7455);
or U8075 (N_8075,N_7395,N_6870);
or U8076 (N_8076,N_6861,N_7228);
xor U8077 (N_8077,N_7094,N_7018);
or U8078 (N_8078,N_6808,N_7441);
and U8079 (N_8079,N_7376,N_7343);
nand U8080 (N_8080,N_7249,N_6825);
xnor U8081 (N_8081,N_6825,N_7260);
or U8082 (N_8082,N_6958,N_6774);
or U8083 (N_8083,N_7106,N_6864);
or U8084 (N_8084,N_7459,N_7455);
and U8085 (N_8085,N_7048,N_7498);
nand U8086 (N_8086,N_7416,N_7254);
and U8087 (N_8087,N_7396,N_7159);
and U8088 (N_8088,N_7244,N_6927);
or U8089 (N_8089,N_6825,N_7225);
xor U8090 (N_8090,N_7081,N_7339);
nor U8091 (N_8091,N_6876,N_7034);
xor U8092 (N_8092,N_7097,N_7056);
nor U8093 (N_8093,N_7218,N_7469);
or U8094 (N_8094,N_7494,N_7036);
nor U8095 (N_8095,N_7280,N_7218);
and U8096 (N_8096,N_7103,N_7006);
xor U8097 (N_8097,N_6839,N_7044);
nand U8098 (N_8098,N_7209,N_7380);
or U8099 (N_8099,N_6761,N_7300);
nand U8100 (N_8100,N_6939,N_7447);
and U8101 (N_8101,N_6834,N_7350);
nor U8102 (N_8102,N_7174,N_6833);
or U8103 (N_8103,N_6809,N_6882);
or U8104 (N_8104,N_6827,N_7250);
or U8105 (N_8105,N_7220,N_7101);
nor U8106 (N_8106,N_7156,N_7273);
nor U8107 (N_8107,N_7218,N_7242);
and U8108 (N_8108,N_6785,N_7112);
nand U8109 (N_8109,N_7026,N_7250);
nor U8110 (N_8110,N_7187,N_7164);
and U8111 (N_8111,N_7117,N_7150);
or U8112 (N_8112,N_6909,N_7221);
nor U8113 (N_8113,N_7399,N_7222);
or U8114 (N_8114,N_6788,N_6976);
nor U8115 (N_8115,N_7345,N_6902);
nand U8116 (N_8116,N_7341,N_7391);
or U8117 (N_8117,N_7459,N_7326);
and U8118 (N_8118,N_6957,N_6856);
and U8119 (N_8119,N_6939,N_7203);
and U8120 (N_8120,N_7175,N_7466);
xnor U8121 (N_8121,N_6767,N_7465);
and U8122 (N_8122,N_6820,N_7399);
and U8123 (N_8123,N_7370,N_7058);
nand U8124 (N_8124,N_7272,N_6888);
nor U8125 (N_8125,N_6946,N_7088);
or U8126 (N_8126,N_6971,N_7146);
and U8127 (N_8127,N_7467,N_7288);
or U8128 (N_8128,N_7434,N_7146);
nor U8129 (N_8129,N_6884,N_7486);
xor U8130 (N_8130,N_7080,N_7373);
nor U8131 (N_8131,N_7258,N_6780);
and U8132 (N_8132,N_7068,N_7114);
and U8133 (N_8133,N_6949,N_6843);
or U8134 (N_8134,N_7319,N_7335);
and U8135 (N_8135,N_7130,N_7293);
xnor U8136 (N_8136,N_7077,N_7288);
or U8137 (N_8137,N_7414,N_6967);
or U8138 (N_8138,N_7165,N_6956);
nor U8139 (N_8139,N_6779,N_6766);
nand U8140 (N_8140,N_7032,N_7245);
nor U8141 (N_8141,N_6825,N_6834);
xor U8142 (N_8142,N_7440,N_7419);
and U8143 (N_8143,N_6849,N_6944);
nor U8144 (N_8144,N_6966,N_7372);
nand U8145 (N_8145,N_7478,N_7470);
or U8146 (N_8146,N_6928,N_6790);
and U8147 (N_8147,N_6838,N_7178);
and U8148 (N_8148,N_6950,N_7298);
nand U8149 (N_8149,N_7052,N_7020);
nor U8150 (N_8150,N_7419,N_6956);
nand U8151 (N_8151,N_7274,N_7381);
xnor U8152 (N_8152,N_6961,N_7393);
xnor U8153 (N_8153,N_6758,N_6932);
or U8154 (N_8154,N_6777,N_7273);
and U8155 (N_8155,N_6883,N_6926);
nand U8156 (N_8156,N_6981,N_7140);
or U8157 (N_8157,N_6886,N_7366);
xnor U8158 (N_8158,N_6805,N_6794);
nand U8159 (N_8159,N_7491,N_6975);
nor U8160 (N_8160,N_7370,N_6898);
and U8161 (N_8161,N_7179,N_7397);
or U8162 (N_8162,N_6902,N_6855);
nor U8163 (N_8163,N_6820,N_7011);
or U8164 (N_8164,N_7354,N_7281);
nand U8165 (N_8165,N_7069,N_7388);
nor U8166 (N_8166,N_6935,N_7127);
nor U8167 (N_8167,N_6869,N_7155);
nor U8168 (N_8168,N_7368,N_7424);
nand U8169 (N_8169,N_7488,N_7380);
and U8170 (N_8170,N_7203,N_6769);
and U8171 (N_8171,N_7123,N_6805);
nand U8172 (N_8172,N_7123,N_6761);
nor U8173 (N_8173,N_7469,N_7227);
and U8174 (N_8174,N_6906,N_7180);
nor U8175 (N_8175,N_7295,N_6946);
nor U8176 (N_8176,N_7389,N_6937);
and U8177 (N_8177,N_6940,N_6886);
nand U8178 (N_8178,N_7335,N_7457);
nand U8179 (N_8179,N_7338,N_7070);
xor U8180 (N_8180,N_6786,N_7175);
xor U8181 (N_8181,N_6962,N_6994);
or U8182 (N_8182,N_7132,N_7100);
nand U8183 (N_8183,N_7364,N_6928);
and U8184 (N_8184,N_7398,N_7385);
xnor U8185 (N_8185,N_6918,N_7055);
nand U8186 (N_8186,N_7071,N_7029);
and U8187 (N_8187,N_6898,N_6753);
nor U8188 (N_8188,N_7280,N_7350);
nor U8189 (N_8189,N_7410,N_7305);
or U8190 (N_8190,N_6877,N_7371);
nand U8191 (N_8191,N_7160,N_7039);
or U8192 (N_8192,N_6971,N_7089);
and U8193 (N_8193,N_6753,N_7435);
nand U8194 (N_8194,N_7302,N_7308);
nand U8195 (N_8195,N_7013,N_7422);
xor U8196 (N_8196,N_6989,N_7080);
or U8197 (N_8197,N_7212,N_6804);
nor U8198 (N_8198,N_6990,N_7343);
nand U8199 (N_8199,N_6893,N_7342);
xnor U8200 (N_8200,N_7383,N_7360);
nor U8201 (N_8201,N_7402,N_7281);
or U8202 (N_8202,N_6808,N_7051);
nand U8203 (N_8203,N_7407,N_6768);
xor U8204 (N_8204,N_6987,N_7343);
xor U8205 (N_8205,N_7215,N_7020);
nand U8206 (N_8206,N_6758,N_7497);
xnor U8207 (N_8207,N_7101,N_7449);
nor U8208 (N_8208,N_7331,N_7254);
and U8209 (N_8209,N_7440,N_7347);
and U8210 (N_8210,N_7461,N_7088);
and U8211 (N_8211,N_7034,N_6847);
nor U8212 (N_8212,N_6898,N_6981);
nor U8213 (N_8213,N_6953,N_7246);
xor U8214 (N_8214,N_7066,N_7216);
or U8215 (N_8215,N_6998,N_7065);
or U8216 (N_8216,N_7268,N_7107);
nand U8217 (N_8217,N_7088,N_7481);
and U8218 (N_8218,N_6821,N_6897);
nor U8219 (N_8219,N_7215,N_6758);
or U8220 (N_8220,N_7037,N_7411);
nand U8221 (N_8221,N_7339,N_7364);
and U8222 (N_8222,N_7300,N_7066);
and U8223 (N_8223,N_7481,N_6998);
and U8224 (N_8224,N_7166,N_6813);
xnor U8225 (N_8225,N_7437,N_7235);
and U8226 (N_8226,N_7195,N_7028);
or U8227 (N_8227,N_7187,N_6880);
xor U8228 (N_8228,N_7310,N_7355);
xor U8229 (N_8229,N_6753,N_7112);
or U8230 (N_8230,N_7464,N_7395);
and U8231 (N_8231,N_7156,N_7053);
xnor U8232 (N_8232,N_7247,N_7012);
or U8233 (N_8233,N_6990,N_7259);
xor U8234 (N_8234,N_7330,N_7388);
or U8235 (N_8235,N_7297,N_7212);
and U8236 (N_8236,N_6811,N_6910);
nor U8237 (N_8237,N_7295,N_6884);
xnor U8238 (N_8238,N_7360,N_7180);
xor U8239 (N_8239,N_7262,N_7158);
and U8240 (N_8240,N_6957,N_7252);
nand U8241 (N_8241,N_6769,N_7209);
nand U8242 (N_8242,N_6875,N_7265);
xor U8243 (N_8243,N_7034,N_6803);
nor U8244 (N_8244,N_7101,N_7136);
nand U8245 (N_8245,N_7161,N_6962);
nor U8246 (N_8246,N_7316,N_6913);
nand U8247 (N_8247,N_7168,N_7090);
nor U8248 (N_8248,N_6769,N_6796);
xnor U8249 (N_8249,N_6790,N_7206);
nor U8250 (N_8250,N_8108,N_8226);
or U8251 (N_8251,N_8014,N_7739);
nand U8252 (N_8252,N_8143,N_7531);
or U8253 (N_8253,N_7829,N_8135);
and U8254 (N_8254,N_7873,N_8104);
or U8255 (N_8255,N_7765,N_7535);
and U8256 (N_8256,N_7591,N_8086);
or U8257 (N_8257,N_8157,N_8244);
nand U8258 (N_8258,N_7619,N_7760);
xor U8259 (N_8259,N_7952,N_7746);
or U8260 (N_8260,N_7823,N_8103);
or U8261 (N_8261,N_8061,N_7945);
nand U8262 (N_8262,N_8243,N_7964);
xor U8263 (N_8263,N_7686,N_7502);
or U8264 (N_8264,N_7525,N_7902);
nand U8265 (N_8265,N_7658,N_8122);
nor U8266 (N_8266,N_7824,N_8238);
nor U8267 (N_8267,N_8242,N_7917);
xnor U8268 (N_8268,N_7642,N_7710);
xor U8269 (N_8269,N_7646,N_7708);
xnor U8270 (N_8270,N_8126,N_8218);
and U8271 (N_8271,N_7817,N_7992);
or U8272 (N_8272,N_7779,N_7684);
and U8273 (N_8273,N_8015,N_7866);
and U8274 (N_8274,N_8141,N_7890);
or U8275 (N_8275,N_7532,N_8233);
nor U8276 (N_8276,N_8113,N_7828);
xnor U8277 (N_8277,N_7534,N_7566);
nor U8278 (N_8278,N_7986,N_8118);
nor U8279 (N_8279,N_7682,N_7975);
or U8280 (N_8280,N_7640,N_8094);
nor U8281 (N_8281,N_7764,N_7941);
or U8282 (N_8282,N_8160,N_7622);
or U8283 (N_8283,N_7604,N_7745);
and U8284 (N_8284,N_8105,N_7568);
xor U8285 (N_8285,N_7643,N_7996);
nor U8286 (N_8286,N_7972,N_8140);
and U8287 (N_8287,N_7961,N_7834);
or U8288 (N_8288,N_8182,N_8077);
xor U8289 (N_8289,N_7599,N_8235);
or U8290 (N_8290,N_8054,N_7989);
nor U8291 (N_8291,N_8180,N_8032);
and U8292 (N_8292,N_7762,N_8188);
xor U8293 (N_8293,N_7889,N_8205);
and U8294 (N_8294,N_7785,N_7722);
or U8295 (N_8295,N_7512,N_7700);
nand U8296 (N_8296,N_7656,N_7691);
and U8297 (N_8297,N_7618,N_7954);
xor U8298 (N_8298,N_7935,N_7901);
xnor U8299 (N_8299,N_8234,N_7672);
and U8300 (N_8300,N_8149,N_8021);
nand U8301 (N_8301,N_7578,N_7925);
and U8302 (N_8302,N_8178,N_7826);
xnor U8303 (N_8303,N_7895,N_7805);
or U8304 (N_8304,N_7825,N_7988);
nor U8305 (N_8305,N_7795,N_7606);
nor U8306 (N_8306,N_7997,N_7868);
xor U8307 (N_8307,N_8246,N_7729);
nand U8308 (N_8308,N_7685,N_7908);
and U8309 (N_8309,N_7832,N_7918);
nand U8310 (N_8310,N_8227,N_8042);
and U8311 (N_8311,N_7709,N_7649);
or U8312 (N_8312,N_8045,N_7536);
or U8313 (N_8313,N_8080,N_8120);
nor U8314 (N_8314,N_7724,N_7523);
nand U8315 (N_8315,N_7524,N_7590);
nand U8316 (N_8316,N_7963,N_8138);
or U8317 (N_8317,N_7584,N_7737);
or U8318 (N_8318,N_7600,N_8079);
xnor U8319 (N_8319,N_8147,N_7513);
nor U8320 (N_8320,N_7893,N_8100);
xor U8321 (N_8321,N_7620,N_8039);
or U8322 (N_8322,N_7645,N_7693);
xnor U8323 (N_8323,N_8137,N_7511);
nand U8324 (N_8324,N_7863,N_7850);
xnor U8325 (N_8325,N_7597,N_7831);
or U8326 (N_8326,N_8187,N_7688);
and U8327 (N_8327,N_7929,N_7652);
or U8328 (N_8328,N_8085,N_7968);
nor U8329 (N_8329,N_7521,N_8223);
xnor U8330 (N_8330,N_7923,N_7812);
xor U8331 (N_8331,N_7806,N_7987);
nand U8332 (N_8332,N_8175,N_8241);
nand U8333 (N_8333,N_8169,N_7696);
and U8334 (N_8334,N_7697,N_7938);
nor U8335 (N_8335,N_7603,N_8065);
nand U8336 (N_8336,N_7638,N_7569);
xor U8337 (N_8337,N_7689,N_7849);
nand U8338 (N_8338,N_7843,N_7811);
nor U8339 (N_8339,N_8196,N_8035);
or U8340 (N_8340,N_7706,N_7628);
and U8341 (N_8341,N_7506,N_8151);
nand U8342 (N_8342,N_7616,N_7860);
and U8343 (N_8343,N_8165,N_7567);
nor U8344 (N_8344,N_7687,N_7756);
or U8345 (N_8345,N_7520,N_7884);
or U8346 (N_8346,N_7916,N_8066);
nor U8347 (N_8347,N_7799,N_7920);
nand U8348 (N_8348,N_7728,N_8220);
xor U8349 (N_8349,N_7958,N_7538);
nand U8350 (N_8350,N_7668,N_7576);
xor U8351 (N_8351,N_8133,N_7654);
or U8352 (N_8352,N_7936,N_7796);
nand U8353 (N_8353,N_8199,N_7882);
and U8354 (N_8354,N_7951,N_7841);
or U8355 (N_8355,N_7803,N_8029);
nor U8356 (N_8356,N_7983,N_7851);
xor U8357 (N_8357,N_7790,N_8225);
nand U8358 (N_8358,N_8146,N_8091);
nor U8359 (N_8359,N_7778,N_7580);
or U8360 (N_8360,N_8174,N_8047);
and U8361 (N_8361,N_7814,N_8222);
and U8362 (N_8362,N_7744,N_7942);
nor U8363 (N_8363,N_7894,N_8150);
nand U8364 (N_8364,N_7801,N_7653);
nand U8365 (N_8365,N_7934,N_7683);
nand U8366 (N_8366,N_7897,N_7807);
nor U8367 (N_8367,N_8060,N_7820);
xnor U8368 (N_8368,N_8072,N_8069);
nor U8369 (N_8369,N_7982,N_7639);
xnor U8370 (N_8370,N_7822,N_7571);
or U8371 (N_8371,N_7671,N_7690);
or U8372 (N_8372,N_7699,N_7607);
xnor U8373 (N_8373,N_7940,N_7927);
and U8374 (N_8374,N_7818,N_7510);
or U8375 (N_8375,N_7809,N_7769);
and U8376 (N_8376,N_7853,N_7577);
or U8377 (N_8377,N_8158,N_8007);
or U8378 (N_8378,N_7953,N_8041);
and U8379 (N_8379,N_8051,N_8012);
nor U8380 (N_8380,N_7838,N_7768);
nor U8381 (N_8381,N_7859,N_7957);
nand U8382 (N_8382,N_8183,N_7657);
nand U8383 (N_8383,N_8232,N_7854);
nor U8384 (N_8384,N_7904,N_7899);
or U8385 (N_8385,N_7614,N_8101);
nor U8386 (N_8386,N_7847,N_7558);
nor U8387 (N_8387,N_7501,N_8185);
and U8388 (N_8388,N_8209,N_8081);
nor U8389 (N_8389,N_7922,N_7973);
xor U8390 (N_8390,N_7780,N_8073);
xnor U8391 (N_8391,N_7991,N_8154);
or U8392 (N_8392,N_8228,N_7594);
and U8393 (N_8393,N_7694,N_7881);
xor U8394 (N_8394,N_7971,N_7837);
xor U8395 (N_8395,N_7673,N_7727);
xnor U8396 (N_8396,N_8026,N_7743);
nor U8397 (N_8397,N_7912,N_7979);
xnor U8398 (N_8398,N_7886,N_8134);
nor U8399 (N_8399,N_8170,N_8167);
xor U8400 (N_8400,N_8111,N_7835);
nand U8401 (N_8401,N_7741,N_7667);
or U8402 (N_8402,N_7869,N_7602);
or U8403 (N_8403,N_8123,N_7574);
nand U8404 (N_8404,N_8239,N_8215);
or U8405 (N_8405,N_7755,N_8190);
nand U8406 (N_8406,N_7840,N_7615);
xnor U8407 (N_8407,N_7621,N_7816);
nand U8408 (N_8408,N_7583,N_8128);
xnor U8409 (N_8409,N_7518,N_7937);
and U8410 (N_8410,N_8097,N_7582);
nand U8411 (N_8411,N_7990,N_8152);
nor U8412 (N_8412,N_7862,N_7549);
nor U8413 (N_8413,N_7770,N_8189);
xor U8414 (N_8414,N_7877,N_7794);
nor U8415 (N_8415,N_7924,N_8142);
nor U8416 (N_8416,N_7575,N_8159);
or U8417 (N_8417,N_8231,N_7802);
nor U8418 (N_8418,N_8092,N_8020);
or U8419 (N_8419,N_7675,N_7980);
xnor U8420 (N_8420,N_8095,N_7844);
or U8421 (N_8421,N_7871,N_7752);
nor U8422 (N_8422,N_7857,N_7633);
nor U8423 (N_8423,N_8206,N_7872);
or U8424 (N_8424,N_7514,N_8040);
nand U8425 (N_8425,N_8207,N_7641);
xor U8426 (N_8426,N_8213,N_8139);
nand U8427 (N_8427,N_7733,N_7933);
nand U8428 (N_8428,N_7730,N_8071);
xnor U8429 (N_8429,N_8116,N_8049);
and U8430 (N_8430,N_8063,N_7855);
and U8431 (N_8431,N_7928,N_7867);
nor U8432 (N_8432,N_7742,N_7692);
and U8433 (N_8433,N_8121,N_8181);
and U8434 (N_8434,N_8186,N_8155);
nand U8435 (N_8435,N_8229,N_7681);
and U8436 (N_8436,N_8098,N_7879);
nor U8437 (N_8437,N_7508,N_7763);
or U8438 (N_8438,N_8062,N_8176);
or U8439 (N_8439,N_7856,N_7542);
nand U8440 (N_8440,N_8070,N_7720);
nand U8441 (N_8441,N_8038,N_8217);
nand U8442 (N_8442,N_7962,N_8096);
and U8443 (N_8443,N_7662,N_7792);
or U8444 (N_8444,N_7800,N_7553);
nand U8445 (N_8445,N_7605,N_8053);
and U8446 (N_8446,N_7703,N_7715);
and U8447 (N_8447,N_7978,N_8212);
xor U8448 (N_8448,N_7726,N_7959);
nand U8449 (N_8449,N_8002,N_7913);
xor U8450 (N_8450,N_8153,N_7588);
nand U8451 (N_8451,N_8127,N_7533);
and U8452 (N_8452,N_7637,N_8088);
xnor U8453 (N_8453,N_7595,N_7999);
nor U8454 (N_8454,N_7680,N_7707);
and U8455 (N_8455,N_8168,N_8249);
or U8456 (N_8456,N_7892,N_7677);
or U8457 (N_8457,N_7556,N_7581);
nand U8458 (N_8458,N_7970,N_7914);
and U8459 (N_8459,N_8030,N_7659);
or U8460 (N_8460,N_7788,N_7655);
and U8461 (N_8461,N_7716,N_7617);
nand U8462 (N_8462,N_8197,N_8119);
or U8463 (N_8463,N_7725,N_7804);
nor U8464 (N_8464,N_8093,N_7723);
nor U8465 (N_8465,N_7557,N_8194);
or U8466 (N_8466,N_7827,N_7839);
or U8467 (N_8467,N_7539,N_8166);
and U8468 (N_8468,N_7547,N_7887);
xor U8469 (N_8469,N_7550,N_7573);
or U8470 (N_8470,N_7977,N_7561);
and U8471 (N_8471,N_7836,N_7878);
xor U8472 (N_8472,N_7787,N_8203);
xnor U8473 (N_8473,N_7864,N_8240);
xnor U8474 (N_8474,N_8107,N_7736);
xnor U8475 (N_8475,N_7630,N_7585);
and U8476 (N_8476,N_7503,N_8237);
nand U8477 (N_8477,N_8136,N_8075);
nor U8478 (N_8478,N_7905,N_8099);
and U8479 (N_8479,N_8184,N_8214);
nor U8480 (N_8480,N_8004,N_7526);
nand U8481 (N_8481,N_8008,N_8083);
or U8482 (N_8482,N_7903,N_8089);
and U8483 (N_8483,N_7842,N_7593);
nand U8484 (N_8484,N_7915,N_7559);
or U8485 (N_8485,N_8018,N_7735);
nand U8486 (N_8486,N_7519,N_8028);
nor U8487 (N_8487,N_7896,N_7898);
nand U8488 (N_8488,N_7679,N_7664);
and U8489 (N_8489,N_7663,N_8017);
or U8490 (N_8490,N_7965,N_8248);
and U8491 (N_8491,N_7625,N_7740);
and U8492 (N_8492,N_8058,N_7563);
nand U8493 (N_8493,N_7782,N_8023);
nand U8494 (N_8494,N_7966,N_7738);
or U8495 (N_8495,N_8144,N_8109);
or U8496 (N_8496,N_8076,N_7516);
xor U8497 (N_8497,N_7974,N_7946);
nor U8498 (N_8498,N_7791,N_8090);
and U8499 (N_8499,N_7609,N_8162);
or U8500 (N_8500,N_7624,N_7852);
or U8501 (N_8501,N_8210,N_7956);
nand U8502 (N_8502,N_7711,N_7732);
xnor U8503 (N_8503,N_7527,N_8013);
nand U8504 (N_8504,N_7775,N_7589);
nor U8505 (N_8505,N_7717,N_7921);
or U8506 (N_8506,N_8031,N_8036);
nand U8507 (N_8507,N_7552,N_7949);
or U8508 (N_8508,N_7670,N_8172);
nor U8509 (N_8509,N_7880,N_8124);
and U8510 (N_8510,N_7598,N_7955);
or U8511 (N_8511,N_7650,N_7810);
nand U8512 (N_8512,N_7613,N_8164);
nand U8513 (N_8513,N_7704,N_7660);
or U8514 (N_8514,N_7555,N_7906);
and U8515 (N_8515,N_7540,N_7734);
and U8516 (N_8516,N_7932,N_7751);
nor U8517 (N_8517,N_7783,N_7909);
xor U8518 (N_8518,N_8048,N_8208);
xor U8519 (N_8519,N_7784,N_8025);
or U8520 (N_8520,N_7786,N_7611);
xnor U8521 (N_8521,N_7910,N_8037);
and U8522 (N_8522,N_8236,N_7610);
and U8523 (N_8523,N_8115,N_8106);
xnor U8524 (N_8524,N_8056,N_7874);
nand U8525 (N_8525,N_7623,N_7712);
nor U8526 (N_8526,N_7774,N_7939);
nor U8527 (N_8527,N_7608,N_8132);
and U8528 (N_8528,N_8192,N_7793);
and U8529 (N_8529,N_8084,N_7947);
or U8530 (N_8530,N_8010,N_7661);
nor U8531 (N_8531,N_7517,N_7579);
nand U8532 (N_8532,N_7900,N_7926);
xnor U8533 (N_8533,N_8082,N_7813);
and U8534 (N_8534,N_7572,N_7976);
and U8535 (N_8535,N_7530,N_7592);
or U8536 (N_8536,N_8078,N_7626);
and U8537 (N_8537,N_8173,N_8163);
nor U8538 (N_8538,N_7870,N_7754);
xor U8539 (N_8539,N_7848,N_7701);
nand U8540 (N_8540,N_8202,N_7644);
or U8541 (N_8541,N_8171,N_8057);
nand U8542 (N_8542,N_7985,N_8130);
xor U8543 (N_8543,N_7674,N_8156);
nor U8544 (N_8544,N_7981,N_7930);
nor U8545 (N_8545,N_7647,N_7773);
nor U8546 (N_8546,N_7718,N_7676);
nand U8547 (N_8547,N_8044,N_7543);
xor U8548 (N_8548,N_7969,N_8204);
or U8549 (N_8549,N_7865,N_8005);
nor U8550 (N_8550,N_8043,N_8230);
nand U8551 (N_8551,N_8191,N_7815);
nand U8552 (N_8552,N_7819,N_7705);
xor U8553 (N_8553,N_7601,N_7500);
and U8554 (N_8554,N_7570,N_7846);
and U8555 (N_8555,N_8019,N_7509);
nor U8556 (N_8556,N_7781,N_8195);
and U8557 (N_8557,N_8221,N_7797);
nand U8558 (N_8558,N_8193,N_7875);
or U8559 (N_8559,N_7504,N_7919);
xnor U8560 (N_8560,N_7544,N_7960);
or U8561 (N_8561,N_8000,N_7507);
nand U8562 (N_8562,N_7776,N_7721);
nand U8563 (N_8563,N_8145,N_8027);
nand U8564 (N_8564,N_7631,N_8050);
or U8565 (N_8565,N_7548,N_7562);
and U8566 (N_8566,N_7761,N_7749);
or U8567 (N_8567,N_7876,N_8129);
or U8568 (N_8568,N_7789,N_7944);
nand U8569 (N_8569,N_7714,N_8003);
or U8570 (N_8570,N_7702,N_7546);
or U8571 (N_8571,N_7515,N_7528);
nor U8572 (N_8572,N_7907,N_7665);
nand U8573 (N_8573,N_7713,N_7545);
and U8574 (N_8574,N_7750,N_8052);
xnor U8575 (N_8575,N_7747,N_8211);
nor U8576 (N_8576,N_7636,N_7541);
xnor U8577 (N_8577,N_7596,N_7967);
nand U8578 (N_8578,N_8064,N_7943);
or U8579 (N_8579,N_7767,N_8046);
xnor U8580 (N_8580,N_8022,N_7948);
and U8581 (N_8581,N_7529,N_7883);
and U8582 (N_8582,N_8068,N_7522);
and U8583 (N_8583,N_8016,N_7748);
xor U8584 (N_8584,N_7833,N_8001);
nand U8585 (N_8585,N_7911,N_7719);
nor U8586 (N_8586,N_7931,N_7505);
or U8587 (N_8587,N_8067,N_8247);
and U8588 (N_8588,N_7629,N_8200);
and U8589 (N_8589,N_7731,N_7560);
and U8590 (N_8590,N_8087,N_7888);
nor U8591 (N_8591,N_7757,N_8112);
nand U8592 (N_8592,N_7891,N_7669);
xor U8593 (N_8593,N_7861,N_7993);
xnor U8594 (N_8594,N_7758,N_7753);
xnor U8595 (N_8595,N_8177,N_8245);
nor U8596 (N_8596,N_7551,N_7771);
xor U8597 (N_8597,N_7759,N_7695);
or U8598 (N_8598,N_8219,N_8009);
and U8599 (N_8599,N_7777,N_8055);
nor U8600 (N_8600,N_7565,N_7648);
nand U8601 (N_8601,N_7698,N_7798);
or U8602 (N_8602,N_7666,N_7537);
or U8603 (N_8603,N_7564,N_7766);
and U8604 (N_8604,N_7885,N_7994);
xnor U8605 (N_8605,N_7830,N_7821);
xnor U8606 (N_8606,N_8117,N_7858);
nor U8607 (N_8607,N_8074,N_8006);
and U8608 (N_8608,N_8114,N_8110);
nor U8609 (N_8609,N_8125,N_7587);
and U8610 (N_8610,N_7984,N_7612);
or U8611 (N_8611,N_7950,N_8011);
or U8612 (N_8612,N_7845,N_7635);
or U8613 (N_8613,N_8198,N_7634);
xnor U8614 (N_8614,N_7627,N_8148);
or U8615 (N_8615,N_8131,N_7998);
and U8616 (N_8616,N_8024,N_8161);
or U8617 (N_8617,N_8224,N_8216);
or U8618 (N_8618,N_7554,N_7995);
nand U8619 (N_8619,N_7678,N_8034);
nor U8620 (N_8620,N_8201,N_7632);
nand U8621 (N_8621,N_8179,N_7772);
nor U8622 (N_8622,N_8033,N_7808);
or U8623 (N_8623,N_7586,N_8059);
or U8624 (N_8624,N_8102,N_7651);
nor U8625 (N_8625,N_7738,N_8005);
or U8626 (N_8626,N_7885,N_7975);
or U8627 (N_8627,N_7529,N_7738);
or U8628 (N_8628,N_7956,N_8099);
and U8629 (N_8629,N_8204,N_7626);
xnor U8630 (N_8630,N_7587,N_7765);
and U8631 (N_8631,N_7772,N_7893);
nor U8632 (N_8632,N_8057,N_7925);
and U8633 (N_8633,N_7833,N_8034);
nor U8634 (N_8634,N_8030,N_8029);
xnor U8635 (N_8635,N_7622,N_7538);
xnor U8636 (N_8636,N_7878,N_7503);
nand U8637 (N_8637,N_7709,N_8050);
or U8638 (N_8638,N_8086,N_8115);
or U8639 (N_8639,N_7835,N_7506);
and U8640 (N_8640,N_7626,N_8249);
nor U8641 (N_8641,N_7841,N_7670);
and U8642 (N_8642,N_7546,N_8202);
nand U8643 (N_8643,N_7773,N_7786);
or U8644 (N_8644,N_7756,N_8069);
nand U8645 (N_8645,N_8057,N_7771);
xor U8646 (N_8646,N_7797,N_7550);
nand U8647 (N_8647,N_8245,N_7961);
nand U8648 (N_8648,N_8146,N_7559);
nor U8649 (N_8649,N_7720,N_7661);
nor U8650 (N_8650,N_7644,N_7970);
or U8651 (N_8651,N_7721,N_7668);
or U8652 (N_8652,N_7532,N_7828);
nand U8653 (N_8653,N_7504,N_8234);
nor U8654 (N_8654,N_8133,N_7895);
nor U8655 (N_8655,N_7884,N_8023);
xor U8656 (N_8656,N_8054,N_7749);
nand U8657 (N_8657,N_7574,N_7745);
nand U8658 (N_8658,N_7878,N_8031);
nor U8659 (N_8659,N_7762,N_7928);
nand U8660 (N_8660,N_7585,N_8161);
nor U8661 (N_8661,N_8161,N_7671);
and U8662 (N_8662,N_8109,N_7722);
nand U8663 (N_8663,N_7594,N_7924);
nor U8664 (N_8664,N_8206,N_7821);
and U8665 (N_8665,N_8034,N_8134);
and U8666 (N_8666,N_7542,N_7826);
nor U8667 (N_8667,N_8005,N_7647);
xor U8668 (N_8668,N_7791,N_8219);
and U8669 (N_8669,N_7929,N_7978);
xnor U8670 (N_8670,N_8159,N_7862);
or U8671 (N_8671,N_7818,N_7649);
nor U8672 (N_8672,N_8165,N_7769);
and U8673 (N_8673,N_7878,N_8242);
or U8674 (N_8674,N_8103,N_7951);
nand U8675 (N_8675,N_8192,N_8237);
or U8676 (N_8676,N_7925,N_7915);
xnor U8677 (N_8677,N_7794,N_8202);
or U8678 (N_8678,N_7506,N_7943);
nor U8679 (N_8679,N_7788,N_7577);
or U8680 (N_8680,N_7932,N_8140);
nand U8681 (N_8681,N_7771,N_7950);
or U8682 (N_8682,N_7889,N_8081);
or U8683 (N_8683,N_8207,N_8085);
and U8684 (N_8684,N_7978,N_7752);
or U8685 (N_8685,N_8091,N_7791);
nor U8686 (N_8686,N_8005,N_7588);
nor U8687 (N_8687,N_8166,N_7752);
or U8688 (N_8688,N_8197,N_7679);
xor U8689 (N_8689,N_7973,N_7905);
and U8690 (N_8690,N_8030,N_7634);
nor U8691 (N_8691,N_7827,N_8038);
nand U8692 (N_8692,N_7771,N_7981);
and U8693 (N_8693,N_7882,N_8217);
xor U8694 (N_8694,N_7563,N_7898);
nand U8695 (N_8695,N_7654,N_7914);
and U8696 (N_8696,N_7758,N_7840);
or U8697 (N_8697,N_7641,N_7793);
nor U8698 (N_8698,N_7833,N_7543);
and U8699 (N_8699,N_8153,N_7552);
nand U8700 (N_8700,N_8182,N_7505);
xnor U8701 (N_8701,N_7754,N_7966);
or U8702 (N_8702,N_7906,N_8207);
nand U8703 (N_8703,N_8170,N_7748);
or U8704 (N_8704,N_8205,N_7911);
nand U8705 (N_8705,N_7785,N_8197);
and U8706 (N_8706,N_7900,N_7568);
xnor U8707 (N_8707,N_7775,N_7846);
and U8708 (N_8708,N_8075,N_7519);
nand U8709 (N_8709,N_8225,N_8073);
or U8710 (N_8710,N_8132,N_8187);
xnor U8711 (N_8711,N_7771,N_7742);
nor U8712 (N_8712,N_7736,N_7564);
nand U8713 (N_8713,N_7686,N_7825);
nor U8714 (N_8714,N_7716,N_7774);
nand U8715 (N_8715,N_8106,N_8134);
nor U8716 (N_8716,N_7754,N_7695);
nand U8717 (N_8717,N_7500,N_7567);
or U8718 (N_8718,N_7869,N_7942);
or U8719 (N_8719,N_7675,N_7609);
or U8720 (N_8720,N_8026,N_8116);
nor U8721 (N_8721,N_7901,N_7881);
and U8722 (N_8722,N_7667,N_8056);
xor U8723 (N_8723,N_7758,N_7806);
or U8724 (N_8724,N_8060,N_7766);
or U8725 (N_8725,N_8100,N_8000);
nor U8726 (N_8726,N_7642,N_8177);
and U8727 (N_8727,N_8023,N_7689);
and U8728 (N_8728,N_7763,N_7866);
and U8729 (N_8729,N_7650,N_7724);
or U8730 (N_8730,N_7559,N_8194);
or U8731 (N_8731,N_7648,N_7961);
and U8732 (N_8732,N_8030,N_7520);
or U8733 (N_8733,N_7851,N_7748);
or U8734 (N_8734,N_7510,N_7713);
or U8735 (N_8735,N_7914,N_7559);
or U8736 (N_8736,N_8052,N_7801);
and U8737 (N_8737,N_7623,N_8052);
and U8738 (N_8738,N_8207,N_7918);
xor U8739 (N_8739,N_7556,N_7708);
nand U8740 (N_8740,N_7546,N_7891);
nor U8741 (N_8741,N_8180,N_8107);
or U8742 (N_8742,N_8180,N_7506);
and U8743 (N_8743,N_7789,N_7936);
or U8744 (N_8744,N_8143,N_8240);
nand U8745 (N_8745,N_7830,N_7628);
nor U8746 (N_8746,N_8224,N_7726);
or U8747 (N_8747,N_8192,N_7858);
or U8748 (N_8748,N_8242,N_7714);
or U8749 (N_8749,N_8079,N_7988);
nand U8750 (N_8750,N_8101,N_7518);
xnor U8751 (N_8751,N_7615,N_8029);
xor U8752 (N_8752,N_8217,N_7608);
xor U8753 (N_8753,N_8176,N_8163);
xnor U8754 (N_8754,N_7898,N_7597);
nand U8755 (N_8755,N_8174,N_8235);
or U8756 (N_8756,N_7647,N_7632);
nand U8757 (N_8757,N_7658,N_7840);
or U8758 (N_8758,N_8079,N_7665);
xor U8759 (N_8759,N_8187,N_7687);
or U8760 (N_8760,N_8095,N_7867);
or U8761 (N_8761,N_7553,N_7856);
and U8762 (N_8762,N_8184,N_7644);
nand U8763 (N_8763,N_7722,N_7943);
xor U8764 (N_8764,N_7661,N_7913);
nand U8765 (N_8765,N_8224,N_8018);
or U8766 (N_8766,N_7605,N_7785);
and U8767 (N_8767,N_8077,N_7624);
nor U8768 (N_8768,N_8127,N_7650);
xor U8769 (N_8769,N_7569,N_7613);
or U8770 (N_8770,N_7751,N_7676);
or U8771 (N_8771,N_7763,N_7673);
or U8772 (N_8772,N_8033,N_7781);
xnor U8773 (N_8773,N_7786,N_7748);
xnor U8774 (N_8774,N_7534,N_8024);
and U8775 (N_8775,N_7820,N_7780);
nor U8776 (N_8776,N_8183,N_7727);
or U8777 (N_8777,N_7926,N_7948);
nand U8778 (N_8778,N_7584,N_8100);
or U8779 (N_8779,N_7660,N_7917);
or U8780 (N_8780,N_7527,N_7767);
nand U8781 (N_8781,N_7821,N_7946);
or U8782 (N_8782,N_7725,N_7667);
nor U8783 (N_8783,N_8055,N_8072);
and U8784 (N_8784,N_8197,N_7869);
or U8785 (N_8785,N_7855,N_8121);
or U8786 (N_8786,N_7605,N_7742);
and U8787 (N_8787,N_7963,N_7579);
nor U8788 (N_8788,N_8238,N_7959);
nand U8789 (N_8789,N_7761,N_7864);
xor U8790 (N_8790,N_8217,N_7710);
nand U8791 (N_8791,N_7553,N_8110);
nor U8792 (N_8792,N_8064,N_7614);
or U8793 (N_8793,N_7844,N_7860);
nor U8794 (N_8794,N_8068,N_7880);
nor U8795 (N_8795,N_7918,N_7927);
xnor U8796 (N_8796,N_8222,N_8084);
or U8797 (N_8797,N_7688,N_8177);
nor U8798 (N_8798,N_7508,N_8063);
nor U8799 (N_8799,N_7673,N_7610);
or U8800 (N_8800,N_8233,N_7786);
nand U8801 (N_8801,N_7567,N_7594);
or U8802 (N_8802,N_7898,N_8021);
nand U8803 (N_8803,N_7592,N_8026);
xor U8804 (N_8804,N_8182,N_7555);
nand U8805 (N_8805,N_7789,N_7756);
nand U8806 (N_8806,N_7888,N_8112);
xor U8807 (N_8807,N_8192,N_8216);
nand U8808 (N_8808,N_7844,N_8139);
or U8809 (N_8809,N_8101,N_7539);
and U8810 (N_8810,N_7604,N_7764);
or U8811 (N_8811,N_7839,N_7519);
and U8812 (N_8812,N_7887,N_8093);
and U8813 (N_8813,N_7557,N_7597);
nand U8814 (N_8814,N_7542,N_7740);
and U8815 (N_8815,N_8190,N_7908);
or U8816 (N_8816,N_7733,N_8026);
or U8817 (N_8817,N_7876,N_8142);
nand U8818 (N_8818,N_8194,N_7592);
xor U8819 (N_8819,N_7558,N_7903);
xor U8820 (N_8820,N_7525,N_8204);
xor U8821 (N_8821,N_8124,N_7884);
and U8822 (N_8822,N_8081,N_8104);
nand U8823 (N_8823,N_7629,N_7758);
or U8824 (N_8824,N_7688,N_8248);
or U8825 (N_8825,N_8222,N_8090);
nand U8826 (N_8826,N_7721,N_7720);
nand U8827 (N_8827,N_7721,N_7834);
and U8828 (N_8828,N_7780,N_8248);
and U8829 (N_8829,N_8160,N_7844);
nor U8830 (N_8830,N_7564,N_8190);
and U8831 (N_8831,N_7602,N_7648);
xnor U8832 (N_8832,N_8244,N_7810);
and U8833 (N_8833,N_7881,N_8190);
and U8834 (N_8834,N_8188,N_8047);
xnor U8835 (N_8835,N_8147,N_7652);
or U8836 (N_8836,N_8244,N_7784);
nor U8837 (N_8837,N_8007,N_7603);
or U8838 (N_8838,N_8034,N_8236);
and U8839 (N_8839,N_7932,N_8091);
xnor U8840 (N_8840,N_7705,N_7571);
nor U8841 (N_8841,N_7667,N_8052);
and U8842 (N_8842,N_7892,N_8033);
nand U8843 (N_8843,N_8180,N_7863);
xor U8844 (N_8844,N_8103,N_7588);
or U8845 (N_8845,N_7715,N_7943);
or U8846 (N_8846,N_8171,N_8021);
and U8847 (N_8847,N_8149,N_7966);
xnor U8848 (N_8848,N_8000,N_7570);
nand U8849 (N_8849,N_8182,N_8234);
xnor U8850 (N_8850,N_8129,N_7961);
or U8851 (N_8851,N_8245,N_7544);
and U8852 (N_8852,N_7929,N_7607);
or U8853 (N_8853,N_7654,N_7656);
xor U8854 (N_8854,N_8073,N_8095);
xor U8855 (N_8855,N_7959,N_7891);
or U8856 (N_8856,N_8117,N_7763);
xor U8857 (N_8857,N_7581,N_7707);
or U8858 (N_8858,N_8127,N_7903);
nand U8859 (N_8859,N_7739,N_8048);
and U8860 (N_8860,N_7656,N_7773);
xor U8861 (N_8861,N_7787,N_8188);
xnor U8862 (N_8862,N_8232,N_8078);
or U8863 (N_8863,N_8192,N_8166);
or U8864 (N_8864,N_7820,N_7748);
xnor U8865 (N_8865,N_7871,N_8197);
xor U8866 (N_8866,N_7833,N_7958);
nor U8867 (N_8867,N_7536,N_8102);
xor U8868 (N_8868,N_7926,N_7928);
and U8869 (N_8869,N_7990,N_7603);
nor U8870 (N_8870,N_8066,N_8172);
and U8871 (N_8871,N_7670,N_7745);
nand U8872 (N_8872,N_7995,N_7786);
nand U8873 (N_8873,N_7663,N_7669);
and U8874 (N_8874,N_7690,N_8084);
nand U8875 (N_8875,N_7564,N_7872);
nor U8876 (N_8876,N_7954,N_7579);
nand U8877 (N_8877,N_7631,N_8089);
and U8878 (N_8878,N_7944,N_7957);
xor U8879 (N_8879,N_7674,N_7821);
xor U8880 (N_8880,N_8169,N_7731);
xnor U8881 (N_8881,N_7528,N_7805);
nor U8882 (N_8882,N_8082,N_7861);
and U8883 (N_8883,N_8035,N_7895);
nor U8884 (N_8884,N_8086,N_7745);
xor U8885 (N_8885,N_8150,N_7875);
or U8886 (N_8886,N_7529,N_8110);
xor U8887 (N_8887,N_7653,N_7880);
and U8888 (N_8888,N_7725,N_8084);
xnor U8889 (N_8889,N_7568,N_8237);
nor U8890 (N_8890,N_7869,N_8022);
and U8891 (N_8891,N_7527,N_7854);
nand U8892 (N_8892,N_7719,N_7627);
xor U8893 (N_8893,N_8027,N_7874);
nand U8894 (N_8894,N_7704,N_7948);
nor U8895 (N_8895,N_7995,N_7964);
nand U8896 (N_8896,N_7929,N_7778);
and U8897 (N_8897,N_7559,N_7995);
nand U8898 (N_8898,N_7882,N_7723);
xor U8899 (N_8899,N_8090,N_8210);
or U8900 (N_8900,N_7813,N_7559);
or U8901 (N_8901,N_7738,N_7765);
nand U8902 (N_8902,N_7636,N_8247);
nand U8903 (N_8903,N_8025,N_7742);
xor U8904 (N_8904,N_7732,N_7786);
nor U8905 (N_8905,N_7840,N_7889);
nor U8906 (N_8906,N_8027,N_7769);
or U8907 (N_8907,N_8201,N_7795);
and U8908 (N_8908,N_7723,N_7560);
xor U8909 (N_8909,N_7761,N_7653);
or U8910 (N_8910,N_8248,N_7587);
and U8911 (N_8911,N_8163,N_7635);
nand U8912 (N_8912,N_8115,N_7561);
and U8913 (N_8913,N_7508,N_7765);
or U8914 (N_8914,N_7751,N_7643);
nor U8915 (N_8915,N_7734,N_7815);
nor U8916 (N_8916,N_7706,N_8206);
and U8917 (N_8917,N_7618,N_8063);
or U8918 (N_8918,N_7597,N_7731);
nand U8919 (N_8919,N_8043,N_7776);
xor U8920 (N_8920,N_7836,N_7704);
nand U8921 (N_8921,N_8227,N_7944);
and U8922 (N_8922,N_7542,N_7572);
and U8923 (N_8923,N_8209,N_8084);
and U8924 (N_8924,N_7513,N_7899);
xnor U8925 (N_8925,N_7539,N_7651);
nor U8926 (N_8926,N_7504,N_7802);
or U8927 (N_8927,N_8083,N_7599);
xor U8928 (N_8928,N_7502,N_7530);
xor U8929 (N_8929,N_7682,N_7617);
or U8930 (N_8930,N_7609,N_7834);
and U8931 (N_8931,N_8120,N_7955);
xnor U8932 (N_8932,N_7628,N_7653);
nor U8933 (N_8933,N_7563,N_7663);
nand U8934 (N_8934,N_7768,N_8127);
or U8935 (N_8935,N_8140,N_8205);
or U8936 (N_8936,N_8211,N_7695);
and U8937 (N_8937,N_7903,N_8063);
or U8938 (N_8938,N_7734,N_7607);
nand U8939 (N_8939,N_7777,N_8039);
nor U8940 (N_8940,N_8183,N_7950);
nor U8941 (N_8941,N_7518,N_8023);
or U8942 (N_8942,N_7712,N_8055);
or U8943 (N_8943,N_7730,N_7625);
nor U8944 (N_8944,N_8053,N_7844);
nor U8945 (N_8945,N_7616,N_8011);
and U8946 (N_8946,N_7617,N_8023);
or U8947 (N_8947,N_7953,N_7534);
xor U8948 (N_8948,N_7714,N_8191);
and U8949 (N_8949,N_7615,N_8012);
xnor U8950 (N_8950,N_8183,N_7620);
nand U8951 (N_8951,N_7598,N_7838);
and U8952 (N_8952,N_7878,N_8021);
xor U8953 (N_8953,N_8211,N_7673);
nor U8954 (N_8954,N_7924,N_7993);
xor U8955 (N_8955,N_7594,N_8195);
xor U8956 (N_8956,N_7789,N_7895);
or U8957 (N_8957,N_8030,N_7528);
xor U8958 (N_8958,N_7600,N_8137);
or U8959 (N_8959,N_7589,N_7684);
and U8960 (N_8960,N_7610,N_7930);
nand U8961 (N_8961,N_8068,N_8004);
nand U8962 (N_8962,N_7668,N_8172);
and U8963 (N_8963,N_7825,N_7501);
nand U8964 (N_8964,N_7610,N_7919);
and U8965 (N_8965,N_8050,N_7839);
nand U8966 (N_8966,N_7916,N_7587);
nand U8967 (N_8967,N_7664,N_7829);
and U8968 (N_8968,N_8100,N_8119);
xor U8969 (N_8969,N_8234,N_7622);
and U8970 (N_8970,N_7716,N_7940);
nand U8971 (N_8971,N_7899,N_8017);
nand U8972 (N_8972,N_7715,N_7645);
or U8973 (N_8973,N_7757,N_7789);
nor U8974 (N_8974,N_7665,N_7837);
and U8975 (N_8975,N_7641,N_8104);
nand U8976 (N_8976,N_8045,N_7762);
and U8977 (N_8977,N_7756,N_7763);
nand U8978 (N_8978,N_8041,N_7907);
or U8979 (N_8979,N_7592,N_7517);
and U8980 (N_8980,N_7896,N_7686);
xnor U8981 (N_8981,N_7533,N_7500);
nor U8982 (N_8982,N_7548,N_7587);
and U8983 (N_8983,N_7737,N_7745);
or U8984 (N_8984,N_8001,N_8200);
and U8985 (N_8985,N_7747,N_8114);
nor U8986 (N_8986,N_7619,N_7919);
or U8987 (N_8987,N_8214,N_8245);
nor U8988 (N_8988,N_7593,N_7936);
xnor U8989 (N_8989,N_7634,N_8233);
nor U8990 (N_8990,N_7797,N_8020);
or U8991 (N_8991,N_8209,N_8055);
xor U8992 (N_8992,N_7981,N_7760);
and U8993 (N_8993,N_7903,N_7666);
xnor U8994 (N_8994,N_8065,N_7581);
and U8995 (N_8995,N_7555,N_7828);
xor U8996 (N_8996,N_8035,N_7800);
xnor U8997 (N_8997,N_7779,N_7578);
and U8998 (N_8998,N_7939,N_8233);
or U8999 (N_8999,N_8089,N_8178);
and U9000 (N_9000,N_8263,N_8730);
xor U9001 (N_9001,N_8967,N_8689);
xor U9002 (N_9002,N_8917,N_8254);
nand U9003 (N_9003,N_8934,N_8463);
xnor U9004 (N_9004,N_8586,N_8672);
and U9005 (N_9005,N_8850,N_8705);
nand U9006 (N_9006,N_8511,N_8845);
and U9007 (N_9007,N_8686,N_8522);
nor U9008 (N_9008,N_8506,N_8420);
or U9009 (N_9009,N_8537,N_8837);
nor U9010 (N_9010,N_8616,N_8653);
xnor U9011 (N_9011,N_8380,N_8859);
or U9012 (N_9012,N_8631,N_8717);
xnor U9013 (N_9013,N_8444,N_8430);
and U9014 (N_9014,N_8601,N_8514);
and U9015 (N_9015,N_8334,N_8714);
or U9016 (N_9016,N_8827,N_8995);
xnor U9017 (N_9017,N_8292,N_8610);
nor U9018 (N_9018,N_8919,N_8501);
nand U9019 (N_9019,N_8895,N_8635);
nor U9020 (N_9020,N_8922,N_8440);
xnor U9021 (N_9021,N_8516,N_8748);
nor U9022 (N_9022,N_8694,N_8603);
and U9023 (N_9023,N_8290,N_8452);
nor U9024 (N_9024,N_8571,N_8346);
xnor U9025 (N_9025,N_8553,N_8413);
and U9026 (N_9026,N_8756,N_8617);
xnor U9027 (N_9027,N_8579,N_8417);
and U9028 (N_9028,N_8453,N_8728);
nor U9029 (N_9029,N_8785,N_8867);
nand U9030 (N_9030,N_8797,N_8989);
nand U9031 (N_9031,N_8426,N_8803);
nand U9032 (N_9032,N_8261,N_8834);
xor U9033 (N_9033,N_8580,N_8367);
nand U9034 (N_9034,N_8805,N_8721);
and U9035 (N_9035,N_8732,N_8351);
nand U9036 (N_9036,N_8814,N_8884);
or U9037 (N_9037,N_8646,N_8977);
nand U9038 (N_9038,N_8527,N_8606);
nor U9039 (N_9039,N_8352,N_8636);
or U9040 (N_9040,N_8353,N_8270);
and U9041 (N_9041,N_8670,N_8633);
or U9042 (N_9042,N_8543,N_8323);
xnor U9043 (N_9043,N_8675,N_8948);
and U9044 (N_9044,N_8360,N_8354);
nand U9045 (N_9045,N_8704,N_8472);
or U9046 (N_9046,N_8999,N_8986);
nor U9047 (N_9047,N_8916,N_8820);
xnor U9048 (N_9048,N_8990,N_8259);
xor U9049 (N_9049,N_8959,N_8398);
nor U9050 (N_9050,N_8528,N_8577);
nand U9051 (N_9051,N_8678,N_8298);
nand U9052 (N_9052,N_8824,N_8602);
nand U9053 (N_9053,N_8681,N_8376);
xor U9054 (N_9054,N_8775,N_8296);
or U9055 (N_9055,N_8768,N_8829);
xnor U9056 (N_9056,N_8666,N_8790);
or U9057 (N_9057,N_8862,N_8906);
and U9058 (N_9058,N_8943,N_8929);
xor U9059 (N_9059,N_8379,N_8719);
and U9060 (N_9060,N_8718,N_8655);
nand U9061 (N_9061,N_8903,N_8411);
and U9062 (N_9062,N_8918,N_8826);
nand U9063 (N_9063,N_8572,N_8536);
nor U9064 (N_9064,N_8341,N_8585);
nand U9065 (N_9065,N_8474,N_8268);
or U9066 (N_9066,N_8578,N_8358);
nand U9067 (N_9067,N_8615,N_8569);
nand U9068 (N_9068,N_8725,N_8915);
nand U9069 (N_9069,N_8520,N_8400);
nor U9070 (N_9070,N_8713,N_8455);
or U9071 (N_9071,N_8484,N_8285);
or U9072 (N_9072,N_8703,N_8423);
nor U9073 (N_9073,N_8876,N_8921);
xor U9074 (N_9074,N_8691,N_8424);
or U9075 (N_9075,N_8562,N_8871);
or U9076 (N_9076,N_8560,N_8992);
xnor U9077 (N_9077,N_8326,N_8330);
or U9078 (N_9078,N_8628,N_8370);
or U9079 (N_9079,N_8264,N_8547);
nor U9080 (N_9080,N_8923,N_8589);
or U9081 (N_9081,N_8657,N_8644);
xor U9082 (N_9082,N_8548,N_8737);
and U9083 (N_9083,N_8676,N_8954);
and U9084 (N_9084,N_8960,N_8744);
or U9085 (N_9085,N_8322,N_8723);
xor U9086 (N_9086,N_8462,N_8498);
nor U9087 (N_9087,N_8561,N_8928);
and U9088 (N_9088,N_8769,N_8503);
or U9089 (N_9089,N_8621,N_8434);
xnor U9090 (N_9090,N_8564,N_8623);
nand U9091 (N_9091,N_8940,N_8611);
nor U9092 (N_9092,N_8594,N_8902);
nand U9093 (N_9093,N_8702,N_8410);
or U9094 (N_9094,N_8979,N_8500);
and U9095 (N_9095,N_8483,N_8557);
or U9096 (N_9096,N_8407,N_8946);
xnor U9097 (N_9097,N_8529,N_8302);
xor U9098 (N_9098,N_8480,N_8901);
xor U9099 (N_9099,N_8396,N_8493);
and U9100 (N_9100,N_8652,N_8552);
or U9101 (N_9101,N_8349,N_8894);
or U9102 (N_9102,N_8466,N_8993);
nand U9103 (N_9103,N_8831,N_8763);
xor U9104 (N_9104,N_8853,N_8679);
nor U9105 (N_9105,N_8605,N_8599);
nand U9106 (N_9106,N_8315,N_8852);
nand U9107 (N_9107,N_8565,N_8937);
xor U9108 (N_9108,N_8377,N_8740);
xnor U9109 (N_9109,N_8549,N_8668);
nand U9110 (N_9110,N_8425,N_8688);
and U9111 (N_9111,N_8684,N_8486);
or U9112 (N_9112,N_8978,N_8471);
xnor U9113 (N_9113,N_8278,N_8447);
xnor U9114 (N_9114,N_8275,N_8970);
nand U9115 (N_9115,N_8707,N_8613);
nor U9116 (N_9116,N_8545,N_8739);
and U9117 (N_9117,N_8595,N_8421);
nand U9118 (N_9118,N_8745,N_8406);
nand U9119 (N_9119,N_8294,N_8587);
nor U9120 (N_9120,N_8658,N_8950);
and U9121 (N_9121,N_8271,N_8764);
nand U9122 (N_9122,N_8865,N_8771);
nand U9123 (N_9123,N_8706,N_8303);
and U9124 (N_9124,N_8632,N_8808);
nor U9125 (N_9125,N_8932,N_8575);
nor U9126 (N_9126,N_8695,N_8625);
or U9127 (N_9127,N_8325,N_8418);
nor U9128 (N_9128,N_8619,N_8807);
nand U9129 (N_9129,N_8281,N_8328);
nand U9130 (N_9130,N_8724,N_8314);
or U9131 (N_9131,N_8373,N_8470);
nor U9132 (N_9132,N_8436,N_8766);
and U9133 (N_9133,N_8609,N_8816);
nor U9134 (N_9134,N_8499,N_8883);
nand U9135 (N_9135,N_8386,N_8487);
nor U9136 (N_9136,N_8854,N_8291);
and U9137 (N_9137,N_8843,N_8512);
nand U9138 (N_9138,N_8382,N_8318);
nand U9139 (N_9139,N_8947,N_8262);
or U9140 (N_9140,N_8600,N_8277);
nand U9141 (N_9141,N_8709,N_8980);
xnor U9142 (N_9142,N_8755,N_8389);
nor U9143 (N_9143,N_8792,N_8985);
and U9144 (N_9144,N_8583,N_8945);
and U9145 (N_9145,N_8332,N_8910);
nor U9146 (N_9146,N_8907,N_8914);
and U9147 (N_9147,N_8267,N_8598);
nor U9148 (N_9148,N_8629,N_8645);
or U9149 (N_9149,N_8478,N_8662);
or U9150 (N_9150,N_8319,N_8445);
nand U9151 (N_9151,N_8881,N_8806);
or U9152 (N_9152,N_8698,N_8639);
xor U9153 (N_9153,N_8309,N_8521);
or U9154 (N_9154,N_8339,N_8607);
or U9155 (N_9155,N_8833,N_8951);
nor U9156 (N_9156,N_8981,N_8530);
nand U9157 (N_9157,N_8348,N_8855);
or U9158 (N_9158,N_8873,N_8663);
or U9159 (N_9159,N_8699,N_8782);
or U9160 (N_9160,N_8804,N_8716);
and U9161 (N_9161,N_8773,N_8643);
nand U9162 (N_9162,N_8523,N_8847);
xor U9163 (N_9163,N_8933,N_8519);
nor U9164 (N_9164,N_8693,N_8612);
xor U9165 (N_9165,N_8671,N_8415);
xnor U9166 (N_9166,N_8255,N_8375);
xnor U9167 (N_9167,N_8435,N_8443);
xor U9168 (N_9168,N_8627,N_8293);
or U9169 (N_9169,N_8822,N_8473);
or U9170 (N_9170,N_8485,N_8531);
xnor U9171 (N_9171,N_8419,N_8535);
and U9172 (N_9172,N_8251,N_8856);
xor U9173 (N_9173,N_8956,N_8458);
or U9174 (N_9174,N_8273,N_8680);
and U9175 (N_9175,N_8930,N_8384);
nor U9176 (N_9176,N_8971,N_8696);
and U9177 (N_9177,N_8720,N_8767);
nor U9178 (N_9178,N_8863,N_8568);
nand U9179 (N_9179,N_8432,N_8563);
and U9180 (N_9180,N_8659,N_8975);
nand U9181 (N_9181,N_8872,N_8591);
or U9182 (N_9182,N_8582,N_8321);
nand U9183 (N_9183,N_8540,N_8801);
and U9184 (N_9184,N_8825,N_8690);
and U9185 (N_9185,N_8338,N_8712);
nand U9186 (N_9186,N_8620,N_8656);
nor U9187 (N_9187,N_8626,N_8835);
xnor U9188 (N_9188,N_8288,N_8687);
xor U9189 (N_9189,N_8700,N_8556);
and U9190 (N_9190,N_8994,N_8282);
or U9191 (N_9191,N_8253,N_8900);
and U9192 (N_9192,N_8592,N_8538);
and U9193 (N_9193,N_8965,N_8555);
and U9194 (N_9194,N_8284,N_8887);
nand U9195 (N_9195,N_8403,N_8622);
or U9196 (N_9196,N_8495,N_8988);
nand U9197 (N_9197,N_8342,N_8673);
and U9198 (N_9198,N_8554,N_8828);
nor U9199 (N_9199,N_8817,N_8750);
nor U9200 (N_9200,N_8559,N_8905);
nand U9201 (N_9201,N_8972,N_8727);
nand U9202 (N_9202,N_8812,N_8889);
nand U9203 (N_9203,N_8795,N_8541);
or U9204 (N_9204,N_8310,N_8283);
and U9205 (N_9205,N_8550,N_8793);
and U9206 (N_9206,N_8810,N_8844);
nor U9207 (N_9207,N_8879,N_8904);
and U9208 (N_9208,N_8931,N_8692);
or U9209 (N_9209,N_8614,N_8335);
and U9210 (N_9210,N_8874,N_8449);
nand U9211 (N_9211,N_8502,N_8343);
nor U9212 (N_9212,N_8701,N_8774);
or U9213 (N_9213,N_8953,N_8401);
nand U9214 (N_9214,N_8414,N_8295);
and U9215 (N_9215,N_8276,N_8504);
or U9216 (N_9216,N_8710,N_8597);
nand U9217 (N_9217,N_8256,N_8925);
and U9218 (N_9218,N_8839,N_8497);
or U9219 (N_9219,N_8908,N_8742);
xnor U9220 (N_9220,N_8383,N_8593);
xor U9221 (N_9221,N_8467,N_8404);
xnor U9222 (N_9222,N_8637,N_8454);
or U9223 (N_9223,N_8913,N_8860);
nand U9224 (N_9224,N_8316,N_8340);
nand U9225 (N_9225,N_8751,N_8753);
and U9226 (N_9226,N_8890,N_8469);
nand U9227 (N_9227,N_8488,N_8783);
xor U9228 (N_9228,N_8539,N_8422);
and U9229 (N_9229,N_8258,N_8306);
nand U9230 (N_9230,N_8747,N_8715);
or U9231 (N_9231,N_8868,N_8708);
or U9232 (N_9232,N_8787,N_8451);
and U9233 (N_9233,N_8558,N_8650);
and U9234 (N_9234,N_8957,N_8460);
nor U9235 (N_9235,N_8477,N_8331);
nand U9236 (N_9236,N_8963,N_8534);
xor U9237 (N_9237,N_8363,N_8909);
nor U9238 (N_9238,N_8926,N_8280);
nand U9239 (N_9239,N_8492,N_8777);
or U9240 (N_9240,N_8266,N_8395);
nand U9241 (N_9241,N_8784,N_8911);
xnor U9242 (N_9242,N_8387,N_8697);
nand U9243 (N_9243,N_8546,N_8481);
and U9244 (N_9244,N_8362,N_8788);
nor U9245 (N_9245,N_8974,N_8991);
nor U9246 (N_9246,N_8821,N_8998);
or U9247 (N_9247,N_8935,N_8412);
xnor U9248 (N_9248,N_8786,N_8364);
nand U9249 (N_9249,N_8405,N_8757);
nand U9250 (N_9250,N_8897,N_8566);
xor U9251 (N_9251,N_8476,N_8870);
nor U9252 (N_9252,N_8733,N_8823);
nor U9253 (N_9253,N_8944,N_8838);
nand U9254 (N_9254,N_8429,N_8955);
nand U9255 (N_9255,N_8260,N_8427);
or U9256 (N_9256,N_8301,N_8796);
and U9257 (N_9257,N_8596,N_8711);
nand U9258 (N_9258,N_8347,N_8857);
nand U9259 (N_9259,N_8736,N_8490);
nor U9260 (N_9260,N_8968,N_8861);
xor U9261 (N_9261,N_8374,N_8297);
nand U9262 (N_9262,N_8896,N_8641);
xnor U9263 (N_9263,N_8976,N_8830);
and U9264 (N_9264,N_8941,N_8532);
or U9265 (N_9265,N_8997,N_8327);
or U9266 (N_9266,N_8344,N_8329);
or U9267 (N_9267,N_8842,N_8982);
nand U9268 (N_9268,N_8576,N_8669);
and U9269 (N_9269,N_8402,N_8508);
or U9270 (N_9270,N_8448,N_8608);
nand U9271 (N_9271,N_8858,N_8388);
and U9272 (N_9272,N_8815,N_8464);
nand U9273 (N_9273,N_8397,N_8677);
and U9274 (N_9274,N_8682,N_8505);
nor U9275 (N_9275,N_8762,N_8252);
xor U9276 (N_9276,N_8938,N_8781);
and U9277 (N_9277,N_8927,N_8969);
xor U9278 (N_9278,N_8851,N_8468);
and U9279 (N_9279,N_8289,N_8973);
nand U9280 (N_9280,N_8356,N_8507);
xor U9281 (N_9281,N_8765,N_8489);
nand U9282 (N_9282,N_8864,N_8813);
or U9283 (N_9283,N_8409,N_8912);
nor U9284 (N_9284,N_8408,N_8726);
nand U9285 (N_9285,N_8588,N_8450);
or U9286 (N_9286,N_8551,N_8664);
nand U9287 (N_9287,N_8840,N_8966);
and U9288 (N_9288,N_8518,N_8604);
or U9289 (N_9289,N_8634,N_8924);
xnor U9290 (N_9290,N_8875,N_8456);
xnor U9291 (N_9291,N_8308,N_8433);
and U9292 (N_9292,N_8819,N_8274);
xnor U9293 (N_9293,N_8882,N_8761);
nand U9294 (N_9294,N_8743,N_8355);
nand U9295 (N_9295,N_8399,N_8891);
and U9296 (N_9296,N_8533,N_8651);
and U9297 (N_9297,N_8479,N_8654);
xor U9298 (N_9298,N_8371,N_8286);
and U9299 (N_9299,N_8381,N_8836);
xnor U9300 (N_9300,N_8811,N_8385);
nor U9301 (N_9301,N_8939,N_8320);
or U9302 (N_9302,N_8789,N_8250);
xnor U9303 (N_9303,N_8517,N_8892);
xor U9304 (N_9304,N_8758,N_8642);
or U9305 (N_9305,N_8630,N_8752);
xor U9306 (N_9306,N_8393,N_8898);
or U9307 (N_9307,N_8265,N_8494);
nand U9308 (N_9308,N_8359,N_8446);
and U9309 (N_9309,N_8665,N_8513);
or U9310 (N_9310,N_8461,N_8899);
or U9311 (N_9311,N_8350,N_8849);
xnor U9312 (N_9312,N_8759,N_8667);
nor U9313 (N_9313,N_8311,N_8734);
xor U9314 (N_9314,N_8780,N_8640);
and U9315 (N_9315,N_8958,N_8324);
and U9316 (N_9316,N_8770,N_8526);
xnor U9317 (N_9317,N_8269,N_8869);
nand U9318 (N_9318,N_8618,N_8567);
or U9319 (N_9319,N_8394,N_8313);
and U9320 (N_9320,N_8584,N_8841);
or U9321 (N_9321,N_8305,N_8416);
and U9322 (N_9322,N_8441,N_8439);
nor U9323 (N_9323,N_8648,N_8800);
nand U9324 (N_9324,N_8333,N_8952);
and U9325 (N_9325,N_8866,N_8888);
nor U9326 (N_9326,N_8573,N_8660);
xnor U9327 (N_9327,N_8590,N_8345);
or U9328 (N_9328,N_8936,N_8457);
and U9329 (N_9329,N_8496,N_8459);
and U9330 (N_9330,N_8515,N_8964);
nand U9331 (N_9331,N_8776,N_8674);
or U9332 (N_9332,N_8299,N_8337);
nor U9333 (N_9333,N_8920,N_8818);
nand U9334 (N_9334,N_8731,N_8846);
and U9335 (N_9335,N_8525,N_8391);
xnor U9336 (N_9336,N_8361,N_8638);
nand U9337 (N_9337,N_8544,N_8312);
or U9338 (N_9338,N_8392,N_8794);
or U9339 (N_9339,N_8257,N_8791);
nor U9340 (N_9340,N_8649,N_8437);
nand U9341 (N_9341,N_8877,N_8749);
nor U9342 (N_9342,N_8428,N_8746);
or U9343 (N_9343,N_8741,N_8366);
and U9344 (N_9344,N_8685,N_8799);
nand U9345 (N_9345,N_8482,N_8369);
or U9346 (N_9346,N_8510,N_8279);
or U9347 (N_9347,N_8996,N_8683);
nand U9348 (N_9348,N_8809,N_8307);
nand U9349 (N_9349,N_8722,N_8893);
nor U9350 (N_9350,N_8475,N_8832);
xor U9351 (N_9351,N_8438,N_8987);
nand U9352 (N_9352,N_8570,N_8984);
nand U9353 (N_9353,N_8779,N_8983);
xor U9354 (N_9354,N_8754,N_8880);
nand U9355 (N_9355,N_8878,N_8772);
and U9356 (N_9356,N_8509,N_8942);
and U9357 (N_9357,N_8336,N_8729);
and U9358 (N_9358,N_8661,N_8574);
and U9359 (N_9359,N_8581,N_8304);
and U9360 (N_9360,N_8961,N_8524);
nand U9361 (N_9361,N_8778,N_8798);
and U9362 (N_9362,N_8465,N_8287);
or U9363 (N_9363,N_8542,N_8848);
nor U9364 (N_9364,N_8624,N_8760);
and U9365 (N_9365,N_8735,N_8802);
xor U9366 (N_9366,N_8962,N_8431);
xnor U9367 (N_9367,N_8885,N_8886);
nor U9368 (N_9368,N_8738,N_8949);
nor U9369 (N_9369,N_8390,N_8647);
and U9370 (N_9370,N_8491,N_8378);
nand U9371 (N_9371,N_8372,N_8368);
or U9372 (N_9372,N_8317,N_8272);
nor U9373 (N_9373,N_8442,N_8365);
and U9374 (N_9374,N_8300,N_8357);
nand U9375 (N_9375,N_8904,N_8430);
nand U9376 (N_9376,N_8336,N_8696);
or U9377 (N_9377,N_8587,N_8741);
nand U9378 (N_9378,N_8861,N_8394);
or U9379 (N_9379,N_8730,N_8548);
xor U9380 (N_9380,N_8645,N_8671);
nand U9381 (N_9381,N_8743,N_8633);
and U9382 (N_9382,N_8752,N_8623);
nor U9383 (N_9383,N_8802,N_8663);
or U9384 (N_9384,N_8996,N_8311);
and U9385 (N_9385,N_8301,N_8285);
or U9386 (N_9386,N_8288,N_8267);
and U9387 (N_9387,N_8936,N_8806);
nand U9388 (N_9388,N_8485,N_8490);
xor U9389 (N_9389,N_8384,N_8772);
or U9390 (N_9390,N_8725,N_8392);
nor U9391 (N_9391,N_8544,N_8609);
nor U9392 (N_9392,N_8641,N_8649);
nor U9393 (N_9393,N_8737,N_8517);
nor U9394 (N_9394,N_8250,N_8669);
and U9395 (N_9395,N_8284,N_8748);
or U9396 (N_9396,N_8499,N_8503);
nor U9397 (N_9397,N_8568,N_8316);
and U9398 (N_9398,N_8495,N_8434);
xnor U9399 (N_9399,N_8549,N_8845);
nand U9400 (N_9400,N_8645,N_8737);
or U9401 (N_9401,N_8428,N_8453);
nand U9402 (N_9402,N_8716,N_8256);
or U9403 (N_9403,N_8336,N_8952);
xnor U9404 (N_9404,N_8667,N_8373);
nor U9405 (N_9405,N_8947,N_8787);
and U9406 (N_9406,N_8958,N_8821);
xor U9407 (N_9407,N_8618,N_8258);
xor U9408 (N_9408,N_8453,N_8581);
or U9409 (N_9409,N_8290,N_8484);
or U9410 (N_9410,N_8526,N_8714);
nor U9411 (N_9411,N_8759,N_8684);
nand U9412 (N_9412,N_8431,N_8489);
or U9413 (N_9413,N_8618,N_8612);
and U9414 (N_9414,N_8966,N_8415);
nand U9415 (N_9415,N_8884,N_8761);
or U9416 (N_9416,N_8699,N_8798);
nor U9417 (N_9417,N_8670,N_8688);
xnor U9418 (N_9418,N_8859,N_8613);
nand U9419 (N_9419,N_8830,N_8736);
or U9420 (N_9420,N_8422,N_8961);
xor U9421 (N_9421,N_8753,N_8876);
nor U9422 (N_9422,N_8338,N_8581);
and U9423 (N_9423,N_8866,N_8511);
and U9424 (N_9424,N_8987,N_8571);
nand U9425 (N_9425,N_8748,N_8554);
and U9426 (N_9426,N_8707,N_8382);
and U9427 (N_9427,N_8631,N_8914);
and U9428 (N_9428,N_8511,N_8749);
and U9429 (N_9429,N_8423,N_8580);
nand U9430 (N_9430,N_8845,N_8455);
or U9431 (N_9431,N_8986,N_8557);
and U9432 (N_9432,N_8507,N_8317);
and U9433 (N_9433,N_8964,N_8304);
and U9434 (N_9434,N_8817,N_8753);
nor U9435 (N_9435,N_8660,N_8773);
nand U9436 (N_9436,N_8815,N_8570);
or U9437 (N_9437,N_8619,N_8903);
nand U9438 (N_9438,N_8561,N_8456);
and U9439 (N_9439,N_8690,N_8894);
or U9440 (N_9440,N_8350,N_8791);
and U9441 (N_9441,N_8321,N_8429);
xnor U9442 (N_9442,N_8890,N_8885);
xnor U9443 (N_9443,N_8995,N_8911);
and U9444 (N_9444,N_8879,N_8399);
nor U9445 (N_9445,N_8960,N_8637);
xor U9446 (N_9446,N_8893,N_8697);
xor U9447 (N_9447,N_8782,N_8789);
or U9448 (N_9448,N_8331,N_8674);
or U9449 (N_9449,N_8965,N_8424);
xor U9450 (N_9450,N_8942,N_8536);
and U9451 (N_9451,N_8732,N_8714);
nor U9452 (N_9452,N_8831,N_8915);
xor U9453 (N_9453,N_8338,N_8259);
or U9454 (N_9454,N_8639,N_8681);
xnor U9455 (N_9455,N_8694,N_8546);
nand U9456 (N_9456,N_8531,N_8701);
or U9457 (N_9457,N_8410,N_8384);
or U9458 (N_9458,N_8736,N_8859);
nor U9459 (N_9459,N_8323,N_8724);
nand U9460 (N_9460,N_8704,N_8675);
xor U9461 (N_9461,N_8264,N_8563);
nand U9462 (N_9462,N_8499,N_8767);
and U9463 (N_9463,N_8741,N_8351);
nor U9464 (N_9464,N_8379,N_8827);
or U9465 (N_9465,N_8331,N_8679);
nor U9466 (N_9466,N_8935,N_8739);
xor U9467 (N_9467,N_8940,N_8596);
nand U9468 (N_9468,N_8453,N_8838);
and U9469 (N_9469,N_8721,N_8963);
and U9470 (N_9470,N_8279,N_8801);
nor U9471 (N_9471,N_8820,N_8337);
nor U9472 (N_9472,N_8349,N_8854);
xnor U9473 (N_9473,N_8827,N_8470);
and U9474 (N_9474,N_8492,N_8345);
nand U9475 (N_9475,N_8522,N_8349);
or U9476 (N_9476,N_8601,N_8909);
or U9477 (N_9477,N_8284,N_8690);
xnor U9478 (N_9478,N_8609,N_8797);
and U9479 (N_9479,N_8881,N_8618);
nor U9480 (N_9480,N_8971,N_8925);
nor U9481 (N_9481,N_8857,N_8367);
or U9482 (N_9482,N_8855,N_8773);
nor U9483 (N_9483,N_8788,N_8385);
xnor U9484 (N_9484,N_8727,N_8790);
nor U9485 (N_9485,N_8303,N_8771);
nor U9486 (N_9486,N_8304,N_8441);
and U9487 (N_9487,N_8268,N_8935);
nor U9488 (N_9488,N_8804,N_8749);
or U9489 (N_9489,N_8430,N_8393);
and U9490 (N_9490,N_8416,N_8939);
nor U9491 (N_9491,N_8527,N_8853);
nand U9492 (N_9492,N_8338,N_8525);
nor U9493 (N_9493,N_8853,N_8327);
nor U9494 (N_9494,N_8810,N_8412);
xor U9495 (N_9495,N_8293,N_8756);
nand U9496 (N_9496,N_8322,N_8738);
or U9497 (N_9497,N_8680,N_8765);
xor U9498 (N_9498,N_8920,N_8707);
nand U9499 (N_9499,N_8723,N_8885);
nand U9500 (N_9500,N_8829,N_8993);
nand U9501 (N_9501,N_8302,N_8715);
or U9502 (N_9502,N_8808,N_8443);
nor U9503 (N_9503,N_8353,N_8761);
xnor U9504 (N_9504,N_8752,N_8767);
nor U9505 (N_9505,N_8965,N_8996);
nand U9506 (N_9506,N_8789,N_8279);
and U9507 (N_9507,N_8276,N_8957);
or U9508 (N_9508,N_8597,N_8583);
and U9509 (N_9509,N_8858,N_8586);
and U9510 (N_9510,N_8945,N_8470);
xor U9511 (N_9511,N_8609,N_8499);
and U9512 (N_9512,N_8976,N_8871);
xor U9513 (N_9513,N_8664,N_8679);
nor U9514 (N_9514,N_8881,N_8947);
xor U9515 (N_9515,N_8417,N_8534);
nand U9516 (N_9516,N_8663,N_8311);
nand U9517 (N_9517,N_8848,N_8740);
nor U9518 (N_9518,N_8501,N_8490);
and U9519 (N_9519,N_8965,N_8841);
or U9520 (N_9520,N_8622,N_8955);
or U9521 (N_9521,N_8705,N_8974);
xor U9522 (N_9522,N_8615,N_8533);
xnor U9523 (N_9523,N_8783,N_8319);
nor U9524 (N_9524,N_8452,N_8312);
nand U9525 (N_9525,N_8520,N_8875);
nand U9526 (N_9526,N_8282,N_8987);
nand U9527 (N_9527,N_8380,N_8546);
nor U9528 (N_9528,N_8324,N_8582);
xnor U9529 (N_9529,N_8494,N_8766);
and U9530 (N_9530,N_8468,N_8709);
or U9531 (N_9531,N_8487,N_8408);
nor U9532 (N_9532,N_8709,N_8448);
xor U9533 (N_9533,N_8905,N_8705);
or U9534 (N_9534,N_8718,N_8575);
or U9535 (N_9535,N_8968,N_8781);
nand U9536 (N_9536,N_8392,N_8503);
xor U9537 (N_9537,N_8295,N_8437);
xnor U9538 (N_9538,N_8761,N_8507);
nor U9539 (N_9539,N_8270,N_8879);
nor U9540 (N_9540,N_8346,N_8704);
and U9541 (N_9541,N_8737,N_8510);
xor U9542 (N_9542,N_8414,N_8694);
nor U9543 (N_9543,N_8885,N_8854);
and U9544 (N_9544,N_8955,N_8418);
or U9545 (N_9545,N_8978,N_8855);
nor U9546 (N_9546,N_8361,N_8655);
and U9547 (N_9547,N_8839,N_8319);
nor U9548 (N_9548,N_8943,N_8434);
or U9549 (N_9549,N_8991,N_8305);
or U9550 (N_9550,N_8251,N_8836);
and U9551 (N_9551,N_8797,N_8489);
nor U9552 (N_9552,N_8922,N_8593);
xor U9553 (N_9553,N_8974,N_8925);
or U9554 (N_9554,N_8328,N_8392);
xor U9555 (N_9555,N_8613,N_8417);
or U9556 (N_9556,N_8531,N_8816);
nor U9557 (N_9557,N_8629,N_8809);
nor U9558 (N_9558,N_8447,N_8311);
nor U9559 (N_9559,N_8380,N_8592);
xor U9560 (N_9560,N_8473,N_8448);
or U9561 (N_9561,N_8307,N_8895);
nor U9562 (N_9562,N_8611,N_8605);
xnor U9563 (N_9563,N_8882,N_8312);
nand U9564 (N_9564,N_8908,N_8898);
or U9565 (N_9565,N_8957,N_8906);
nand U9566 (N_9566,N_8883,N_8406);
nand U9567 (N_9567,N_8894,N_8605);
or U9568 (N_9568,N_8871,N_8891);
nor U9569 (N_9569,N_8392,N_8522);
nand U9570 (N_9570,N_8257,N_8696);
nor U9571 (N_9571,N_8278,N_8320);
and U9572 (N_9572,N_8462,N_8555);
and U9573 (N_9573,N_8933,N_8605);
and U9574 (N_9574,N_8874,N_8536);
nor U9575 (N_9575,N_8731,N_8940);
xor U9576 (N_9576,N_8825,N_8359);
and U9577 (N_9577,N_8516,N_8923);
nand U9578 (N_9578,N_8532,N_8352);
and U9579 (N_9579,N_8796,N_8652);
and U9580 (N_9580,N_8420,N_8441);
nand U9581 (N_9581,N_8597,N_8456);
or U9582 (N_9582,N_8432,N_8998);
or U9583 (N_9583,N_8625,N_8325);
or U9584 (N_9584,N_8302,N_8911);
or U9585 (N_9585,N_8636,N_8810);
nor U9586 (N_9586,N_8623,N_8288);
xor U9587 (N_9587,N_8876,N_8866);
xor U9588 (N_9588,N_8482,N_8528);
nand U9589 (N_9589,N_8301,N_8839);
nor U9590 (N_9590,N_8290,N_8829);
xor U9591 (N_9591,N_8850,N_8251);
nor U9592 (N_9592,N_8754,N_8987);
and U9593 (N_9593,N_8534,N_8463);
and U9594 (N_9594,N_8470,N_8768);
nor U9595 (N_9595,N_8813,N_8916);
and U9596 (N_9596,N_8341,N_8609);
nor U9597 (N_9597,N_8402,N_8313);
and U9598 (N_9598,N_8347,N_8400);
nand U9599 (N_9599,N_8434,N_8833);
xor U9600 (N_9600,N_8257,N_8523);
and U9601 (N_9601,N_8956,N_8793);
nor U9602 (N_9602,N_8626,N_8318);
nor U9603 (N_9603,N_8360,N_8362);
nand U9604 (N_9604,N_8721,N_8462);
nand U9605 (N_9605,N_8308,N_8829);
and U9606 (N_9606,N_8822,N_8819);
nand U9607 (N_9607,N_8469,N_8628);
nor U9608 (N_9608,N_8381,N_8566);
xnor U9609 (N_9609,N_8280,N_8356);
xor U9610 (N_9610,N_8742,N_8885);
nand U9611 (N_9611,N_8931,N_8749);
nand U9612 (N_9612,N_8873,N_8938);
nor U9613 (N_9613,N_8334,N_8796);
nand U9614 (N_9614,N_8519,N_8250);
nand U9615 (N_9615,N_8456,N_8507);
nand U9616 (N_9616,N_8632,N_8750);
or U9617 (N_9617,N_8262,N_8917);
xnor U9618 (N_9618,N_8325,N_8382);
and U9619 (N_9619,N_8649,N_8309);
nor U9620 (N_9620,N_8553,N_8698);
xnor U9621 (N_9621,N_8649,N_8388);
and U9622 (N_9622,N_8381,N_8360);
nand U9623 (N_9623,N_8975,N_8689);
xnor U9624 (N_9624,N_8801,N_8818);
nor U9625 (N_9625,N_8668,N_8915);
xnor U9626 (N_9626,N_8926,N_8904);
xor U9627 (N_9627,N_8735,N_8798);
nor U9628 (N_9628,N_8957,N_8959);
nand U9629 (N_9629,N_8561,N_8725);
and U9630 (N_9630,N_8877,N_8449);
or U9631 (N_9631,N_8670,N_8635);
and U9632 (N_9632,N_8290,N_8293);
or U9633 (N_9633,N_8579,N_8606);
xor U9634 (N_9634,N_8602,N_8449);
nand U9635 (N_9635,N_8485,N_8583);
nand U9636 (N_9636,N_8873,N_8448);
or U9637 (N_9637,N_8618,N_8890);
and U9638 (N_9638,N_8872,N_8696);
and U9639 (N_9639,N_8874,N_8529);
and U9640 (N_9640,N_8829,N_8715);
or U9641 (N_9641,N_8643,N_8698);
or U9642 (N_9642,N_8741,N_8385);
and U9643 (N_9643,N_8722,N_8548);
nor U9644 (N_9644,N_8377,N_8558);
xor U9645 (N_9645,N_8879,N_8431);
or U9646 (N_9646,N_8789,N_8640);
or U9647 (N_9647,N_8298,N_8761);
nand U9648 (N_9648,N_8640,N_8683);
nand U9649 (N_9649,N_8395,N_8348);
nor U9650 (N_9650,N_8370,N_8442);
xnor U9651 (N_9651,N_8895,N_8792);
nor U9652 (N_9652,N_8577,N_8388);
xor U9653 (N_9653,N_8500,N_8517);
or U9654 (N_9654,N_8637,N_8360);
xnor U9655 (N_9655,N_8963,N_8434);
or U9656 (N_9656,N_8357,N_8980);
xnor U9657 (N_9657,N_8457,N_8836);
or U9658 (N_9658,N_8530,N_8916);
or U9659 (N_9659,N_8598,N_8884);
nand U9660 (N_9660,N_8320,N_8734);
and U9661 (N_9661,N_8838,N_8970);
and U9662 (N_9662,N_8455,N_8497);
or U9663 (N_9663,N_8402,N_8936);
and U9664 (N_9664,N_8337,N_8871);
xor U9665 (N_9665,N_8536,N_8588);
nand U9666 (N_9666,N_8988,N_8843);
nor U9667 (N_9667,N_8839,N_8660);
nand U9668 (N_9668,N_8451,N_8796);
or U9669 (N_9669,N_8569,N_8273);
xnor U9670 (N_9670,N_8330,N_8741);
nand U9671 (N_9671,N_8802,N_8603);
or U9672 (N_9672,N_8852,N_8430);
and U9673 (N_9673,N_8521,N_8893);
and U9674 (N_9674,N_8490,N_8423);
xnor U9675 (N_9675,N_8561,N_8472);
nor U9676 (N_9676,N_8301,N_8438);
or U9677 (N_9677,N_8655,N_8678);
or U9678 (N_9678,N_8429,N_8371);
nor U9679 (N_9679,N_8947,N_8461);
nand U9680 (N_9680,N_8916,N_8381);
and U9681 (N_9681,N_8587,N_8719);
and U9682 (N_9682,N_8251,N_8587);
and U9683 (N_9683,N_8809,N_8532);
nand U9684 (N_9684,N_8553,N_8496);
or U9685 (N_9685,N_8720,N_8528);
nor U9686 (N_9686,N_8968,N_8288);
nand U9687 (N_9687,N_8513,N_8580);
nor U9688 (N_9688,N_8320,N_8728);
xnor U9689 (N_9689,N_8383,N_8676);
and U9690 (N_9690,N_8986,N_8617);
and U9691 (N_9691,N_8636,N_8274);
nand U9692 (N_9692,N_8695,N_8785);
or U9693 (N_9693,N_8554,N_8448);
and U9694 (N_9694,N_8722,N_8991);
or U9695 (N_9695,N_8735,N_8433);
xor U9696 (N_9696,N_8569,N_8717);
and U9697 (N_9697,N_8379,N_8759);
xor U9698 (N_9698,N_8994,N_8338);
xor U9699 (N_9699,N_8917,N_8829);
and U9700 (N_9700,N_8608,N_8489);
and U9701 (N_9701,N_8677,N_8990);
nand U9702 (N_9702,N_8327,N_8371);
nand U9703 (N_9703,N_8907,N_8638);
nor U9704 (N_9704,N_8483,N_8702);
xor U9705 (N_9705,N_8940,N_8935);
or U9706 (N_9706,N_8674,N_8926);
and U9707 (N_9707,N_8302,N_8638);
or U9708 (N_9708,N_8871,N_8306);
and U9709 (N_9709,N_8442,N_8970);
and U9710 (N_9710,N_8849,N_8594);
nand U9711 (N_9711,N_8486,N_8444);
or U9712 (N_9712,N_8410,N_8476);
nor U9713 (N_9713,N_8290,N_8562);
nor U9714 (N_9714,N_8514,N_8397);
nor U9715 (N_9715,N_8251,N_8497);
nand U9716 (N_9716,N_8479,N_8502);
xnor U9717 (N_9717,N_8868,N_8949);
xnor U9718 (N_9718,N_8417,N_8358);
nor U9719 (N_9719,N_8436,N_8270);
nor U9720 (N_9720,N_8861,N_8675);
and U9721 (N_9721,N_8743,N_8295);
and U9722 (N_9722,N_8929,N_8939);
nor U9723 (N_9723,N_8317,N_8708);
xnor U9724 (N_9724,N_8364,N_8698);
nand U9725 (N_9725,N_8755,N_8885);
nand U9726 (N_9726,N_8843,N_8719);
xnor U9727 (N_9727,N_8368,N_8833);
xor U9728 (N_9728,N_8332,N_8522);
and U9729 (N_9729,N_8724,N_8889);
xnor U9730 (N_9730,N_8531,N_8953);
nand U9731 (N_9731,N_8517,N_8337);
or U9732 (N_9732,N_8617,N_8551);
xnor U9733 (N_9733,N_8719,N_8823);
and U9734 (N_9734,N_8769,N_8617);
nand U9735 (N_9735,N_8625,N_8816);
nor U9736 (N_9736,N_8892,N_8938);
xnor U9737 (N_9737,N_8360,N_8686);
xnor U9738 (N_9738,N_8356,N_8352);
nor U9739 (N_9739,N_8512,N_8778);
or U9740 (N_9740,N_8365,N_8706);
and U9741 (N_9741,N_8269,N_8846);
or U9742 (N_9742,N_8262,N_8487);
or U9743 (N_9743,N_8637,N_8969);
xnor U9744 (N_9744,N_8360,N_8350);
or U9745 (N_9745,N_8397,N_8292);
or U9746 (N_9746,N_8592,N_8734);
nor U9747 (N_9747,N_8296,N_8801);
xor U9748 (N_9748,N_8966,N_8438);
and U9749 (N_9749,N_8265,N_8401);
nand U9750 (N_9750,N_9629,N_9715);
or U9751 (N_9751,N_9139,N_9743);
nand U9752 (N_9752,N_9465,N_9452);
xnor U9753 (N_9753,N_9354,N_9342);
nor U9754 (N_9754,N_9279,N_9632);
and U9755 (N_9755,N_9109,N_9086);
and U9756 (N_9756,N_9462,N_9219);
or U9757 (N_9757,N_9188,N_9107);
xnor U9758 (N_9758,N_9013,N_9010);
xor U9759 (N_9759,N_9403,N_9582);
or U9760 (N_9760,N_9589,N_9607);
nor U9761 (N_9761,N_9301,N_9432);
or U9762 (N_9762,N_9409,N_9055);
and U9763 (N_9763,N_9084,N_9627);
or U9764 (N_9764,N_9089,N_9346);
xor U9765 (N_9765,N_9154,N_9674);
nand U9766 (N_9766,N_9093,N_9562);
nor U9767 (N_9767,N_9115,N_9208);
or U9768 (N_9768,N_9518,N_9027);
nand U9769 (N_9769,N_9413,N_9591);
xor U9770 (N_9770,N_9337,N_9274);
or U9771 (N_9771,N_9426,N_9399);
nor U9772 (N_9772,N_9046,N_9473);
and U9773 (N_9773,N_9125,N_9456);
and U9774 (N_9774,N_9670,N_9169);
xor U9775 (N_9775,N_9039,N_9643);
nor U9776 (N_9776,N_9335,N_9710);
or U9777 (N_9777,N_9034,N_9166);
and U9778 (N_9778,N_9733,N_9564);
xnor U9779 (N_9779,N_9317,N_9334);
nor U9780 (N_9780,N_9680,N_9183);
nor U9781 (N_9781,N_9129,N_9022);
or U9782 (N_9782,N_9150,N_9729);
and U9783 (N_9783,N_9076,N_9061);
nand U9784 (N_9784,N_9740,N_9230);
nand U9785 (N_9785,N_9234,N_9706);
and U9786 (N_9786,N_9072,N_9289);
and U9787 (N_9787,N_9100,N_9396);
and U9788 (N_9788,N_9491,N_9365);
and U9789 (N_9789,N_9269,N_9622);
nor U9790 (N_9790,N_9492,N_9592);
nand U9791 (N_9791,N_9532,N_9387);
nor U9792 (N_9792,N_9425,N_9420);
nand U9793 (N_9793,N_9558,N_9471);
nand U9794 (N_9794,N_9737,N_9173);
or U9795 (N_9795,N_9616,N_9723);
or U9796 (N_9796,N_9391,N_9232);
nor U9797 (N_9797,N_9451,N_9094);
nand U9798 (N_9798,N_9065,N_9583);
nand U9799 (N_9799,N_9698,N_9570);
and U9800 (N_9800,N_9085,N_9685);
xor U9801 (N_9801,N_9559,N_9073);
xor U9802 (N_9802,N_9579,N_9136);
xor U9803 (N_9803,N_9291,N_9598);
nor U9804 (N_9804,N_9043,N_9023);
or U9805 (N_9805,N_9679,N_9481);
nand U9806 (N_9806,N_9653,N_9675);
xor U9807 (N_9807,N_9542,N_9028);
or U9808 (N_9808,N_9207,N_9480);
and U9809 (N_9809,N_9175,N_9709);
nor U9810 (N_9810,N_9398,N_9529);
nor U9811 (N_9811,N_9550,N_9624);
and U9812 (N_9812,N_9021,N_9286);
xnor U9813 (N_9813,N_9442,N_9747);
xor U9814 (N_9814,N_9329,N_9678);
and U9815 (N_9815,N_9356,N_9513);
nand U9816 (N_9816,N_9372,N_9225);
and U9817 (N_9817,N_9204,N_9051);
nor U9818 (N_9818,N_9066,N_9476);
or U9819 (N_9819,N_9263,N_9435);
nand U9820 (N_9820,N_9172,N_9145);
or U9821 (N_9821,N_9433,N_9516);
and U9822 (N_9822,N_9191,N_9295);
or U9823 (N_9823,N_9368,N_9437);
xnor U9824 (N_9824,N_9748,N_9749);
or U9825 (N_9825,N_9272,N_9251);
nand U9826 (N_9826,N_9378,N_9484);
or U9827 (N_9827,N_9738,N_9180);
and U9828 (N_9828,N_9255,N_9408);
nand U9829 (N_9829,N_9415,N_9626);
and U9830 (N_9830,N_9528,N_9104);
and U9831 (N_9831,N_9651,N_9290);
nand U9832 (N_9832,N_9602,N_9495);
xnor U9833 (N_9833,N_9474,N_9047);
or U9834 (N_9834,N_9363,N_9319);
nand U9835 (N_9835,N_9575,N_9736);
nor U9836 (N_9836,N_9177,N_9099);
nor U9837 (N_9837,N_9386,N_9667);
nand U9838 (N_9838,N_9135,N_9041);
and U9839 (N_9839,N_9599,N_9217);
or U9840 (N_9840,N_9276,N_9253);
or U9841 (N_9841,N_9257,N_9282);
nand U9842 (N_9842,N_9436,N_9467);
xor U9843 (N_9843,N_9083,N_9355);
nor U9844 (N_9844,N_9193,N_9470);
or U9845 (N_9845,N_9333,N_9123);
xnor U9846 (N_9846,N_9503,N_9233);
xnor U9847 (N_9847,N_9687,N_9647);
xnor U9848 (N_9848,N_9254,N_9485);
xnor U9849 (N_9849,N_9042,N_9049);
xnor U9850 (N_9850,N_9308,N_9725);
nand U9851 (N_9851,N_9714,N_9210);
and U9852 (N_9852,N_9587,N_9130);
or U9853 (N_9853,N_9520,N_9053);
nand U9854 (N_9854,N_9739,N_9159);
nor U9855 (N_9855,N_9434,N_9641);
nor U9856 (N_9856,N_9557,N_9661);
xnor U9857 (N_9857,N_9197,N_9478);
nand U9858 (N_9858,N_9300,N_9345);
nand U9859 (N_9859,N_9138,N_9414);
xor U9860 (N_9860,N_9638,N_9475);
or U9861 (N_9861,N_9157,N_9140);
nand U9862 (N_9862,N_9548,N_9744);
nor U9863 (N_9863,N_9278,N_9584);
nand U9864 (N_9864,N_9459,N_9577);
nand U9865 (N_9865,N_9350,N_9037);
xor U9866 (N_9866,N_9538,N_9162);
xor U9867 (N_9867,N_9691,N_9701);
or U9868 (N_9868,N_9155,N_9310);
nor U9869 (N_9869,N_9383,N_9273);
nor U9870 (N_9870,N_9699,N_9018);
xnor U9871 (N_9871,N_9305,N_9181);
xor U9872 (N_9872,N_9460,N_9686);
nand U9873 (N_9873,N_9655,N_9215);
and U9874 (N_9874,N_9585,N_9328);
nand U9875 (N_9875,N_9344,N_9332);
and U9876 (N_9876,N_9447,N_9095);
and U9877 (N_9877,N_9298,N_9488);
and U9878 (N_9878,N_9341,N_9149);
xor U9879 (N_9879,N_9718,N_9430);
nor U9880 (N_9880,N_9271,N_9652);
or U9881 (N_9881,N_9620,N_9506);
xnor U9882 (N_9882,N_9270,N_9657);
xor U9883 (N_9883,N_9262,N_9444);
nor U9884 (N_9884,N_9666,N_9654);
xor U9885 (N_9885,N_9292,N_9318);
or U9886 (N_9886,N_9200,N_9347);
nor U9887 (N_9887,N_9745,N_9229);
nand U9888 (N_9888,N_9016,N_9057);
or U9889 (N_9889,N_9025,N_9572);
nor U9890 (N_9890,N_9507,N_9428);
nand U9891 (N_9891,N_9288,N_9091);
nor U9892 (N_9892,N_9320,N_9369);
nand U9893 (N_9893,N_9418,N_9256);
nor U9894 (N_9894,N_9631,N_9165);
nor U9895 (N_9895,N_9127,N_9331);
nor U9896 (N_9896,N_9174,N_9316);
nand U9897 (N_9897,N_9192,N_9058);
or U9898 (N_9898,N_9067,N_9133);
nand U9899 (N_9899,N_9194,N_9722);
and U9900 (N_9900,N_9509,N_9006);
nand U9901 (N_9901,N_9458,N_9704);
and U9902 (N_9902,N_9000,N_9517);
nand U9903 (N_9903,N_9164,N_9479);
and U9904 (N_9904,N_9726,N_9106);
xor U9905 (N_9905,N_9358,N_9730);
xnor U9906 (N_9906,N_9222,N_9658);
xnor U9907 (N_9907,N_9688,N_9179);
nor U9908 (N_9908,N_9032,N_9070);
nor U9909 (N_9909,N_9359,N_9096);
and U9910 (N_9910,N_9201,N_9392);
xnor U9911 (N_9911,N_9078,N_9656);
nand U9912 (N_9912,N_9161,N_9040);
and U9913 (N_9913,N_9168,N_9496);
and U9914 (N_9914,N_9245,N_9593);
or U9915 (N_9915,N_9497,N_9281);
nand U9916 (N_9916,N_9499,N_9595);
xor U9917 (N_9917,N_9732,N_9510);
or U9918 (N_9918,N_9186,N_9526);
xnor U9919 (N_9919,N_9393,N_9122);
or U9920 (N_9920,N_9716,N_9148);
nand U9921 (N_9921,N_9411,N_9068);
and U9922 (N_9922,N_9494,N_9446);
and U9923 (N_9923,N_9594,N_9394);
and U9924 (N_9924,N_9634,N_9611);
or U9925 (N_9925,N_9567,N_9178);
or U9926 (N_9926,N_9486,N_9689);
nor U9927 (N_9927,N_9206,N_9375);
nor U9928 (N_9928,N_9108,N_9609);
or U9929 (N_9929,N_9468,N_9457);
nor U9930 (N_9930,N_9676,N_9530);
nor U9931 (N_9931,N_9578,N_9250);
nand U9932 (N_9932,N_9236,N_9199);
and U9933 (N_9933,N_9639,N_9400);
xnor U9934 (N_9934,N_9581,N_9142);
nand U9935 (N_9935,N_9170,N_9297);
nor U9936 (N_9936,N_9268,N_9552);
nor U9937 (N_9937,N_9090,N_9302);
and U9938 (N_9938,N_9241,N_9543);
and U9939 (N_9939,N_9321,N_9098);
xor U9940 (N_9940,N_9216,N_9322);
nor U9941 (N_9941,N_9146,N_9644);
nand U9942 (N_9942,N_9304,N_9012);
nand U9943 (N_9943,N_9031,N_9610);
or U9944 (N_9944,N_9226,N_9693);
xnor U9945 (N_9945,N_9692,N_9235);
nand U9946 (N_9946,N_9381,N_9612);
and U9947 (N_9947,N_9118,N_9614);
and U9948 (N_9948,N_9101,N_9671);
nand U9949 (N_9949,N_9605,N_9126);
and U9950 (N_9950,N_9364,N_9527);
or U9951 (N_9951,N_9303,N_9002);
xnor U9952 (N_9952,N_9015,N_9209);
and U9953 (N_9953,N_9522,N_9063);
nand U9954 (N_9954,N_9327,N_9697);
nand U9955 (N_9955,N_9665,N_9114);
or U9956 (N_9956,N_9681,N_9533);
nand U9957 (N_9957,N_9071,N_9546);
nand U9958 (N_9958,N_9519,N_9026);
nor U9959 (N_9959,N_9640,N_9137);
nand U9960 (N_9960,N_9454,N_9504);
or U9961 (N_9961,N_9306,N_9370);
nand U9962 (N_9962,N_9044,N_9703);
and U9963 (N_9963,N_9664,N_9330);
xor U9964 (N_9964,N_9410,N_9429);
or U9965 (N_9965,N_9160,N_9036);
nor U9966 (N_9966,N_9555,N_9621);
nand U9967 (N_9967,N_9134,N_9284);
nor U9968 (N_9968,N_9143,N_9185);
nand U9969 (N_9969,N_9153,N_9079);
and U9970 (N_9970,N_9511,N_9625);
nand U9971 (N_9971,N_9218,N_9469);
nand U9972 (N_9972,N_9352,N_9353);
nand U9973 (N_9973,N_9196,N_9111);
nand U9974 (N_9974,N_9544,N_9315);
or U9975 (N_9975,N_9561,N_9240);
and U9976 (N_9976,N_9694,N_9417);
and U9977 (N_9977,N_9682,N_9376);
nor U9978 (N_9978,N_9379,N_9672);
and U9979 (N_9979,N_9662,N_9151);
and U9980 (N_9980,N_9014,N_9385);
xor U9981 (N_9981,N_9244,N_9087);
and U9982 (N_9982,N_9380,N_9650);
nand U9983 (N_9983,N_9711,N_9113);
nand U9984 (N_9984,N_9586,N_9549);
nor U9985 (N_9985,N_9060,N_9734);
nor U9986 (N_9986,N_9539,N_9167);
and U9987 (N_9987,N_9349,N_9074);
nor U9988 (N_9988,N_9228,N_9412);
and U9989 (N_9989,N_9569,N_9189);
and U9990 (N_9990,N_9545,N_9357);
xnor U9991 (N_9991,N_9407,N_9141);
nor U9992 (N_9992,N_9487,N_9563);
nor U9993 (N_9993,N_9742,N_9246);
nand U9994 (N_9994,N_9466,N_9008);
and U9995 (N_9995,N_9597,N_9131);
nand U9996 (N_9996,N_9190,N_9309);
and U9997 (N_9997,N_9649,N_9541);
or U9998 (N_9998,N_9102,N_9119);
nor U9999 (N_9999,N_9038,N_9117);
xor U10000 (N_10000,N_9052,N_9382);
and U10001 (N_10001,N_9677,N_9293);
or U10002 (N_10002,N_9600,N_9259);
and U10003 (N_10003,N_9231,N_9395);
nand U10004 (N_10004,N_9673,N_9648);
or U10005 (N_10005,N_9202,N_9311);
nor U10006 (N_10006,N_9237,N_9384);
xor U10007 (N_10007,N_9182,N_9397);
nand U10008 (N_10008,N_9048,N_9588);
xor U10009 (N_10009,N_9265,N_9735);
and U10010 (N_10010,N_9668,N_9266);
nor U10011 (N_10011,N_9700,N_9500);
nand U10012 (N_10012,N_9323,N_9020);
or U10013 (N_10013,N_9371,N_9324);
nor U10014 (N_10014,N_9580,N_9717);
nor U10015 (N_10015,N_9275,N_9184);
nor U10016 (N_10016,N_9659,N_9314);
nand U10017 (N_10017,N_9419,N_9390);
or U10018 (N_10018,N_9472,N_9283);
nand U10019 (N_10019,N_9551,N_9252);
or U10020 (N_10020,N_9374,N_9388);
nor U10021 (N_10021,N_9069,N_9628);
xor U10022 (N_10022,N_9059,N_9029);
nor U10023 (N_10023,N_9260,N_9512);
nor U10024 (N_10024,N_9493,N_9402);
or U10025 (N_10025,N_9404,N_9004);
nor U10026 (N_10026,N_9105,N_9171);
xor U10027 (N_10027,N_9630,N_9731);
nor U10028 (N_10028,N_9615,N_9361);
nor U10029 (N_10029,N_9075,N_9007);
nor U10030 (N_10030,N_9445,N_9097);
and U10031 (N_10031,N_9195,N_9427);
nor U10032 (N_10032,N_9019,N_9566);
or U10033 (N_10033,N_9116,N_9277);
nor U10034 (N_10034,N_9741,N_9464);
and U10035 (N_10035,N_9326,N_9565);
nand U10036 (N_10036,N_9642,N_9176);
nand U10037 (N_10037,N_9448,N_9213);
and U10038 (N_10038,N_9124,N_9351);
nand U10039 (N_10039,N_9502,N_9081);
nand U10040 (N_10040,N_9571,N_9221);
nand U10041 (N_10041,N_9348,N_9637);
nor U10042 (N_10042,N_9024,N_9377);
nor U10043 (N_10043,N_9483,N_9045);
or U10044 (N_10044,N_9212,N_9477);
nor U10045 (N_10045,N_9088,N_9056);
or U10046 (N_10046,N_9011,N_9623);
nor U10047 (N_10047,N_9121,N_9050);
nand U10048 (N_10048,N_9439,N_9205);
nor U10049 (N_10049,N_9713,N_9147);
or U10050 (N_10050,N_9163,N_9198);
xnor U10051 (N_10051,N_9247,N_9707);
nand U10052 (N_10052,N_9373,N_9505);
nand U10053 (N_10053,N_9401,N_9336);
and U10054 (N_10054,N_9525,N_9267);
xor U10055 (N_10055,N_9660,N_9720);
nor U10056 (N_10056,N_9453,N_9280);
xor U10057 (N_10057,N_9423,N_9537);
xor U10058 (N_10058,N_9482,N_9461);
or U10059 (N_10059,N_9515,N_9243);
or U10060 (N_10060,N_9003,N_9531);
and U10061 (N_10061,N_9223,N_9001);
nor U10062 (N_10062,N_9064,N_9128);
nand U10063 (N_10063,N_9455,N_9695);
nand U10064 (N_10064,N_9239,N_9663);
xnor U10065 (N_10065,N_9633,N_9556);
nor U10066 (N_10066,N_9005,N_9405);
and U10067 (N_10067,N_9683,N_9144);
nand U10068 (N_10068,N_9719,N_9554);
and U10069 (N_10069,N_9211,N_9261);
nor U10070 (N_10070,N_9406,N_9062);
and U10071 (N_10071,N_9514,N_9635);
nand U10072 (N_10072,N_9340,N_9618);
nand U10073 (N_10073,N_9523,N_9367);
or U10074 (N_10074,N_9416,N_9590);
and U10075 (N_10075,N_9501,N_9112);
xor U10076 (N_10076,N_9534,N_9238);
nand U10077 (N_10077,N_9035,N_9712);
nand U10078 (N_10078,N_9613,N_9536);
nor U10079 (N_10079,N_9366,N_9287);
nor U10080 (N_10080,N_9617,N_9343);
nor U10081 (N_10081,N_9489,N_9708);
xnor U10082 (N_10082,N_9441,N_9009);
nor U10083 (N_10083,N_9574,N_9440);
or U10084 (N_10084,N_9152,N_9490);
nand U10085 (N_10085,N_9431,N_9450);
xnor U10086 (N_10086,N_9339,N_9463);
and U10087 (N_10087,N_9521,N_9438);
and U10088 (N_10088,N_9264,N_9285);
nand U10089 (N_10089,N_9158,N_9156);
nand U10090 (N_10090,N_9362,N_9608);
nand U10091 (N_10091,N_9547,N_9313);
and U10092 (N_10092,N_9424,N_9082);
and U10093 (N_10093,N_9422,N_9077);
nand U10094 (N_10094,N_9030,N_9645);
xnor U10095 (N_10095,N_9338,N_9258);
and U10096 (N_10096,N_9203,N_9248);
and U10097 (N_10097,N_9576,N_9603);
nand U10098 (N_10098,N_9296,N_9242);
or U10099 (N_10099,N_9421,N_9033);
or U10100 (N_10100,N_9702,N_9110);
and U10101 (N_10101,N_9601,N_9535);
or U10102 (N_10102,N_9669,N_9724);
nor U10103 (N_10103,N_9604,N_9017);
and U10104 (N_10104,N_9294,N_9214);
xor U10105 (N_10105,N_9498,N_9249);
nand U10106 (N_10106,N_9560,N_9636);
nor U10107 (N_10107,N_9596,N_9092);
nor U10108 (N_10108,N_9187,N_9299);
nand U10109 (N_10109,N_9690,N_9553);
nand U10110 (N_10110,N_9360,N_9705);
nor U10111 (N_10111,N_9443,N_9540);
nand U10112 (N_10112,N_9227,N_9746);
xnor U10113 (N_10113,N_9619,N_9684);
or U10114 (N_10114,N_9646,N_9220);
nor U10115 (N_10115,N_9389,N_9449);
xor U10116 (N_10116,N_9696,N_9080);
nor U10117 (N_10117,N_9508,N_9728);
or U10118 (N_10118,N_9132,N_9224);
xnor U10119 (N_10119,N_9325,N_9727);
nand U10120 (N_10120,N_9054,N_9721);
nand U10121 (N_10121,N_9606,N_9120);
nand U10122 (N_10122,N_9568,N_9312);
or U10123 (N_10123,N_9524,N_9103);
nor U10124 (N_10124,N_9307,N_9573);
nand U10125 (N_10125,N_9676,N_9455);
nor U10126 (N_10126,N_9543,N_9047);
nor U10127 (N_10127,N_9724,N_9039);
or U10128 (N_10128,N_9726,N_9203);
or U10129 (N_10129,N_9253,N_9705);
and U10130 (N_10130,N_9564,N_9659);
nand U10131 (N_10131,N_9279,N_9453);
xor U10132 (N_10132,N_9733,N_9497);
nand U10133 (N_10133,N_9266,N_9430);
nand U10134 (N_10134,N_9119,N_9521);
or U10135 (N_10135,N_9126,N_9604);
nor U10136 (N_10136,N_9624,N_9189);
xnor U10137 (N_10137,N_9437,N_9607);
nand U10138 (N_10138,N_9687,N_9318);
nand U10139 (N_10139,N_9112,N_9124);
or U10140 (N_10140,N_9177,N_9392);
or U10141 (N_10141,N_9655,N_9127);
nor U10142 (N_10142,N_9118,N_9713);
nor U10143 (N_10143,N_9063,N_9286);
xnor U10144 (N_10144,N_9637,N_9504);
and U10145 (N_10145,N_9181,N_9254);
or U10146 (N_10146,N_9098,N_9334);
and U10147 (N_10147,N_9139,N_9480);
nand U10148 (N_10148,N_9271,N_9664);
nor U10149 (N_10149,N_9705,N_9063);
and U10150 (N_10150,N_9076,N_9260);
or U10151 (N_10151,N_9704,N_9228);
xor U10152 (N_10152,N_9677,N_9161);
xor U10153 (N_10153,N_9414,N_9621);
xnor U10154 (N_10154,N_9536,N_9200);
or U10155 (N_10155,N_9168,N_9182);
or U10156 (N_10156,N_9517,N_9217);
or U10157 (N_10157,N_9546,N_9744);
nor U10158 (N_10158,N_9008,N_9475);
nand U10159 (N_10159,N_9059,N_9706);
nand U10160 (N_10160,N_9075,N_9729);
nor U10161 (N_10161,N_9259,N_9241);
nand U10162 (N_10162,N_9040,N_9061);
and U10163 (N_10163,N_9553,N_9716);
nand U10164 (N_10164,N_9545,N_9056);
xnor U10165 (N_10165,N_9264,N_9372);
or U10166 (N_10166,N_9238,N_9472);
nor U10167 (N_10167,N_9527,N_9105);
and U10168 (N_10168,N_9401,N_9009);
or U10169 (N_10169,N_9518,N_9026);
nor U10170 (N_10170,N_9005,N_9308);
nor U10171 (N_10171,N_9232,N_9361);
and U10172 (N_10172,N_9162,N_9484);
nor U10173 (N_10173,N_9526,N_9468);
xor U10174 (N_10174,N_9042,N_9489);
xor U10175 (N_10175,N_9221,N_9692);
or U10176 (N_10176,N_9588,N_9272);
nor U10177 (N_10177,N_9471,N_9357);
nand U10178 (N_10178,N_9133,N_9613);
and U10179 (N_10179,N_9727,N_9708);
or U10180 (N_10180,N_9233,N_9203);
nand U10181 (N_10181,N_9500,N_9670);
and U10182 (N_10182,N_9665,N_9566);
and U10183 (N_10183,N_9013,N_9181);
xnor U10184 (N_10184,N_9186,N_9122);
xor U10185 (N_10185,N_9555,N_9730);
nand U10186 (N_10186,N_9553,N_9552);
xor U10187 (N_10187,N_9310,N_9593);
nand U10188 (N_10188,N_9557,N_9445);
xnor U10189 (N_10189,N_9445,N_9255);
nand U10190 (N_10190,N_9025,N_9509);
nand U10191 (N_10191,N_9201,N_9222);
xnor U10192 (N_10192,N_9424,N_9406);
xnor U10193 (N_10193,N_9486,N_9573);
nor U10194 (N_10194,N_9128,N_9576);
and U10195 (N_10195,N_9718,N_9286);
or U10196 (N_10196,N_9635,N_9023);
nand U10197 (N_10197,N_9588,N_9463);
and U10198 (N_10198,N_9138,N_9713);
and U10199 (N_10199,N_9457,N_9097);
or U10200 (N_10200,N_9445,N_9670);
nor U10201 (N_10201,N_9428,N_9457);
and U10202 (N_10202,N_9422,N_9158);
or U10203 (N_10203,N_9014,N_9287);
xor U10204 (N_10204,N_9577,N_9699);
nand U10205 (N_10205,N_9569,N_9710);
and U10206 (N_10206,N_9011,N_9580);
nand U10207 (N_10207,N_9607,N_9384);
nor U10208 (N_10208,N_9278,N_9235);
xor U10209 (N_10209,N_9179,N_9646);
or U10210 (N_10210,N_9395,N_9293);
xnor U10211 (N_10211,N_9331,N_9507);
nor U10212 (N_10212,N_9382,N_9518);
and U10213 (N_10213,N_9084,N_9209);
xnor U10214 (N_10214,N_9595,N_9487);
or U10215 (N_10215,N_9007,N_9748);
nor U10216 (N_10216,N_9121,N_9485);
nor U10217 (N_10217,N_9740,N_9633);
nor U10218 (N_10218,N_9312,N_9413);
nand U10219 (N_10219,N_9351,N_9558);
and U10220 (N_10220,N_9522,N_9576);
xor U10221 (N_10221,N_9214,N_9219);
xnor U10222 (N_10222,N_9546,N_9405);
and U10223 (N_10223,N_9359,N_9258);
and U10224 (N_10224,N_9112,N_9494);
nand U10225 (N_10225,N_9645,N_9421);
xor U10226 (N_10226,N_9474,N_9417);
nand U10227 (N_10227,N_9658,N_9746);
nor U10228 (N_10228,N_9004,N_9603);
xor U10229 (N_10229,N_9403,N_9227);
xor U10230 (N_10230,N_9723,N_9368);
or U10231 (N_10231,N_9645,N_9261);
nand U10232 (N_10232,N_9107,N_9060);
nor U10233 (N_10233,N_9074,N_9576);
or U10234 (N_10234,N_9679,N_9029);
nor U10235 (N_10235,N_9050,N_9103);
nor U10236 (N_10236,N_9175,N_9734);
nand U10237 (N_10237,N_9198,N_9500);
or U10238 (N_10238,N_9118,N_9512);
nor U10239 (N_10239,N_9478,N_9287);
nor U10240 (N_10240,N_9681,N_9146);
or U10241 (N_10241,N_9705,N_9321);
and U10242 (N_10242,N_9023,N_9356);
nor U10243 (N_10243,N_9090,N_9126);
or U10244 (N_10244,N_9679,N_9498);
and U10245 (N_10245,N_9414,N_9372);
xnor U10246 (N_10246,N_9212,N_9679);
nand U10247 (N_10247,N_9209,N_9555);
and U10248 (N_10248,N_9232,N_9116);
xnor U10249 (N_10249,N_9015,N_9448);
nor U10250 (N_10250,N_9704,N_9529);
and U10251 (N_10251,N_9539,N_9316);
and U10252 (N_10252,N_9174,N_9511);
xnor U10253 (N_10253,N_9135,N_9084);
nand U10254 (N_10254,N_9342,N_9301);
and U10255 (N_10255,N_9304,N_9371);
or U10256 (N_10256,N_9014,N_9610);
nand U10257 (N_10257,N_9121,N_9454);
or U10258 (N_10258,N_9123,N_9199);
and U10259 (N_10259,N_9071,N_9313);
nor U10260 (N_10260,N_9047,N_9597);
nand U10261 (N_10261,N_9199,N_9547);
xnor U10262 (N_10262,N_9741,N_9125);
nand U10263 (N_10263,N_9006,N_9208);
and U10264 (N_10264,N_9040,N_9539);
nor U10265 (N_10265,N_9093,N_9490);
and U10266 (N_10266,N_9412,N_9078);
xor U10267 (N_10267,N_9194,N_9431);
xor U10268 (N_10268,N_9490,N_9480);
nor U10269 (N_10269,N_9545,N_9094);
or U10270 (N_10270,N_9435,N_9013);
nand U10271 (N_10271,N_9598,N_9533);
or U10272 (N_10272,N_9185,N_9304);
nand U10273 (N_10273,N_9430,N_9597);
and U10274 (N_10274,N_9285,N_9038);
nand U10275 (N_10275,N_9061,N_9501);
and U10276 (N_10276,N_9189,N_9006);
or U10277 (N_10277,N_9107,N_9013);
xor U10278 (N_10278,N_9121,N_9243);
and U10279 (N_10279,N_9688,N_9736);
nand U10280 (N_10280,N_9272,N_9437);
nand U10281 (N_10281,N_9127,N_9399);
nor U10282 (N_10282,N_9339,N_9567);
nand U10283 (N_10283,N_9671,N_9476);
or U10284 (N_10284,N_9562,N_9188);
or U10285 (N_10285,N_9714,N_9081);
xor U10286 (N_10286,N_9578,N_9338);
or U10287 (N_10287,N_9060,N_9313);
xnor U10288 (N_10288,N_9190,N_9654);
nor U10289 (N_10289,N_9226,N_9558);
nand U10290 (N_10290,N_9733,N_9670);
nor U10291 (N_10291,N_9093,N_9577);
xnor U10292 (N_10292,N_9189,N_9179);
nand U10293 (N_10293,N_9424,N_9377);
and U10294 (N_10294,N_9607,N_9141);
nor U10295 (N_10295,N_9641,N_9482);
xor U10296 (N_10296,N_9730,N_9420);
nor U10297 (N_10297,N_9121,N_9357);
nor U10298 (N_10298,N_9148,N_9256);
or U10299 (N_10299,N_9174,N_9686);
and U10300 (N_10300,N_9654,N_9680);
and U10301 (N_10301,N_9486,N_9177);
nand U10302 (N_10302,N_9108,N_9105);
nand U10303 (N_10303,N_9006,N_9473);
xnor U10304 (N_10304,N_9213,N_9472);
or U10305 (N_10305,N_9516,N_9380);
or U10306 (N_10306,N_9107,N_9046);
and U10307 (N_10307,N_9181,N_9190);
nor U10308 (N_10308,N_9349,N_9499);
xor U10309 (N_10309,N_9077,N_9696);
xor U10310 (N_10310,N_9124,N_9434);
nor U10311 (N_10311,N_9284,N_9008);
or U10312 (N_10312,N_9293,N_9107);
nand U10313 (N_10313,N_9713,N_9171);
xor U10314 (N_10314,N_9516,N_9039);
nor U10315 (N_10315,N_9736,N_9038);
xor U10316 (N_10316,N_9248,N_9714);
and U10317 (N_10317,N_9353,N_9044);
xnor U10318 (N_10318,N_9555,N_9115);
nand U10319 (N_10319,N_9480,N_9201);
and U10320 (N_10320,N_9402,N_9743);
or U10321 (N_10321,N_9067,N_9098);
or U10322 (N_10322,N_9480,N_9524);
and U10323 (N_10323,N_9449,N_9660);
and U10324 (N_10324,N_9208,N_9457);
nor U10325 (N_10325,N_9266,N_9575);
xnor U10326 (N_10326,N_9710,N_9734);
nand U10327 (N_10327,N_9605,N_9165);
and U10328 (N_10328,N_9692,N_9639);
nor U10329 (N_10329,N_9618,N_9282);
nor U10330 (N_10330,N_9303,N_9610);
xor U10331 (N_10331,N_9193,N_9443);
or U10332 (N_10332,N_9330,N_9223);
xor U10333 (N_10333,N_9131,N_9637);
or U10334 (N_10334,N_9514,N_9405);
or U10335 (N_10335,N_9189,N_9400);
or U10336 (N_10336,N_9298,N_9106);
or U10337 (N_10337,N_9233,N_9101);
nand U10338 (N_10338,N_9102,N_9166);
nor U10339 (N_10339,N_9057,N_9467);
xnor U10340 (N_10340,N_9726,N_9606);
and U10341 (N_10341,N_9357,N_9556);
nand U10342 (N_10342,N_9359,N_9560);
nor U10343 (N_10343,N_9701,N_9485);
xor U10344 (N_10344,N_9142,N_9418);
nor U10345 (N_10345,N_9455,N_9439);
xor U10346 (N_10346,N_9036,N_9663);
and U10347 (N_10347,N_9130,N_9360);
or U10348 (N_10348,N_9568,N_9344);
and U10349 (N_10349,N_9284,N_9644);
or U10350 (N_10350,N_9300,N_9168);
and U10351 (N_10351,N_9230,N_9427);
and U10352 (N_10352,N_9207,N_9506);
or U10353 (N_10353,N_9530,N_9250);
xor U10354 (N_10354,N_9109,N_9328);
and U10355 (N_10355,N_9395,N_9343);
nand U10356 (N_10356,N_9165,N_9749);
xnor U10357 (N_10357,N_9140,N_9516);
nor U10358 (N_10358,N_9384,N_9226);
or U10359 (N_10359,N_9530,N_9295);
nor U10360 (N_10360,N_9479,N_9427);
xor U10361 (N_10361,N_9065,N_9499);
and U10362 (N_10362,N_9127,N_9285);
and U10363 (N_10363,N_9456,N_9341);
and U10364 (N_10364,N_9039,N_9155);
and U10365 (N_10365,N_9480,N_9026);
and U10366 (N_10366,N_9596,N_9259);
xnor U10367 (N_10367,N_9701,N_9544);
or U10368 (N_10368,N_9167,N_9610);
xor U10369 (N_10369,N_9398,N_9302);
or U10370 (N_10370,N_9391,N_9561);
or U10371 (N_10371,N_9224,N_9273);
nand U10372 (N_10372,N_9621,N_9601);
and U10373 (N_10373,N_9701,N_9009);
nor U10374 (N_10374,N_9188,N_9065);
and U10375 (N_10375,N_9115,N_9511);
nand U10376 (N_10376,N_9468,N_9237);
and U10377 (N_10377,N_9630,N_9258);
and U10378 (N_10378,N_9378,N_9647);
and U10379 (N_10379,N_9468,N_9584);
nand U10380 (N_10380,N_9236,N_9655);
xor U10381 (N_10381,N_9122,N_9376);
nor U10382 (N_10382,N_9042,N_9333);
and U10383 (N_10383,N_9399,N_9437);
nor U10384 (N_10384,N_9170,N_9703);
or U10385 (N_10385,N_9525,N_9706);
xor U10386 (N_10386,N_9543,N_9153);
nand U10387 (N_10387,N_9676,N_9188);
xnor U10388 (N_10388,N_9315,N_9000);
nand U10389 (N_10389,N_9639,N_9749);
xor U10390 (N_10390,N_9337,N_9520);
and U10391 (N_10391,N_9738,N_9670);
or U10392 (N_10392,N_9316,N_9080);
and U10393 (N_10393,N_9591,N_9530);
nor U10394 (N_10394,N_9017,N_9731);
nand U10395 (N_10395,N_9036,N_9689);
nor U10396 (N_10396,N_9691,N_9091);
xor U10397 (N_10397,N_9683,N_9495);
and U10398 (N_10398,N_9665,N_9050);
or U10399 (N_10399,N_9641,N_9540);
nor U10400 (N_10400,N_9502,N_9064);
nand U10401 (N_10401,N_9470,N_9156);
nand U10402 (N_10402,N_9407,N_9123);
nand U10403 (N_10403,N_9618,N_9612);
xnor U10404 (N_10404,N_9030,N_9332);
xnor U10405 (N_10405,N_9547,N_9259);
xor U10406 (N_10406,N_9621,N_9254);
and U10407 (N_10407,N_9428,N_9266);
and U10408 (N_10408,N_9353,N_9557);
or U10409 (N_10409,N_9142,N_9744);
nor U10410 (N_10410,N_9067,N_9481);
xor U10411 (N_10411,N_9416,N_9201);
and U10412 (N_10412,N_9523,N_9694);
nor U10413 (N_10413,N_9159,N_9177);
or U10414 (N_10414,N_9068,N_9640);
xnor U10415 (N_10415,N_9513,N_9334);
or U10416 (N_10416,N_9434,N_9654);
xnor U10417 (N_10417,N_9034,N_9540);
or U10418 (N_10418,N_9636,N_9506);
nand U10419 (N_10419,N_9104,N_9256);
and U10420 (N_10420,N_9604,N_9206);
nor U10421 (N_10421,N_9129,N_9505);
and U10422 (N_10422,N_9353,N_9680);
and U10423 (N_10423,N_9046,N_9124);
xnor U10424 (N_10424,N_9162,N_9625);
xor U10425 (N_10425,N_9354,N_9004);
or U10426 (N_10426,N_9699,N_9476);
or U10427 (N_10427,N_9083,N_9171);
nor U10428 (N_10428,N_9485,N_9208);
nand U10429 (N_10429,N_9456,N_9328);
or U10430 (N_10430,N_9672,N_9040);
xnor U10431 (N_10431,N_9556,N_9044);
xor U10432 (N_10432,N_9627,N_9121);
nor U10433 (N_10433,N_9710,N_9641);
nand U10434 (N_10434,N_9533,N_9706);
nand U10435 (N_10435,N_9188,N_9677);
or U10436 (N_10436,N_9432,N_9569);
nor U10437 (N_10437,N_9331,N_9105);
nand U10438 (N_10438,N_9468,N_9380);
nand U10439 (N_10439,N_9498,N_9664);
xor U10440 (N_10440,N_9594,N_9632);
nand U10441 (N_10441,N_9176,N_9738);
xnor U10442 (N_10442,N_9700,N_9724);
nand U10443 (N_10443,N_9608,N_9181);
or U10444 (N_10444,N_9111,N_9379);
or U10445 (N_10445,N_9084,N_9227);
nand U10446 (N_10446,N_9410,N_9275);
nor U10447 (N_10447,N_9110,N_9583);
nor U10448 (N_10448,N_9064,N_9609);
nand U10449 (N_10449,N_9525,N_9286);
and U10450 (N_10450,N_9525,N_9463);
or U10451 (N_10451,N_9583,N_9025);
nor U10452 (N_10452,N_9297,N_9157);
xor U10453 (N_10453,N_9271,N_9236);
nor U10454 (N_10454,N_9135,N_9614);
or U10455 (N_10455,N_9660,N_9736);
or U10456 (N_10456,N_9725,N_9319);
and U10457 (N_10457,N_9120,N_9297);
and U10458 (N_10458,N_9709,N_9112);
nor U10459 (N_10459,N_9379,N_9742);
xnor U10460 (N_10460,N_9648,N_9433);
and U10461 (N_10461,N_9397,N_9571);
nand U10462 (N_10462,N_9172,N_9126);
xnor U10463 (N_10463,N_9165,N_9503);
or U10464 (N_10464,N_9604,N_9176);
and U10465 (N_10465,N_9589,N_9598);
and U10466 (N_10466,N_9733,N_9059);
xnor U10467 (N_10467,N_9322,N_9031);
and U10468 (N_10468,N_9336,N_9325);
or U10469 (N_10469,N_9684,N_9436);
nor U10470 (N_10470,N_9522,N_9189);
or U10471 (N_10471,N_9325,N_9317);
and U10472 (N_10472,N_9467,N_9038);
or U10473 (N_10473,N_9462,N_9600);
xnor U10474 (N_10474,N_9414,N_9370);
or U10475 (N_10475,N_9004,N_9697);
xor U10476 (N_10476,N_9428,N_9178);
xor U10477 (N_10477,N_9018,N_9640);
nor U10478 (N_10478,N_9643,N_9148);
nand U10479 (N_10479,N_9054,N_9240);
xor U10480 (N_10480,N_9603,N_9410);
xor U10481 (N_10481,N_9498,N_9553);
or U10482 (N_10482,N_9597,N_9356);
nor U10483 (N_10483,N_9152,N_9298);
nor U10484 (N_10484,N_9058,N_9017);
nand U10485 (N_10485,N_9619,N_9615);
xor U10486 (N_10486,N_9017,N_9052);
xor U10487 (N_10487,N_9009,N_9455);
or U10488 (N_10488,N_9628,N_9418);
or U10489 (N_10489,N_9266,N_9074);
and U10490 (N_10490,N_9711,N_9453);
nor U10491 (N_10491,N_9413,N_9597);
and U10492 (N_10492,N_9630,N_9367);
and U10493 (N_10493,N_9538,N_9123);
or U10494 (N_10494,N_9424,N_9113);
or U10495 (N_10495,N_9344,N_9709);
xor U10496 (N_10496,N_9363,N_9195);
and U10497 (N_10497,N_9430,N_9521);
or U10498 (N_10498,N_9169,N_9001);
nor U10499 (N_10499,N_9122,N_9298);
or U10500 (N_10500,N_9812,N_10498);
and U10501 (N_10501,N_9934,N_9840);
nor U10502 (N_10502,N_10449,N_10202);
nor U10503 (N_10503,N_9987,N_10243);
and U10504 (N_10504,N_9835,N_9807);
nor U10505 (N_10505,N_10357,N_9904);
or U10506 (N_10506,N_9828,N_10444);
and U10507 (N_10507,N_10104,N_10028);
nor U10508 (N_10508,N_10231,N_10300);
nand U10509 (N_10509,N_10225,N_10322);
nand U10510 (N_10510,N_10380,N_10160);
or U10511 (N_10511,N_10046,N_10060);
and U10512 (N_10512,N_10239,N_9774);
nand U10513 (N_10513,N_10329,N_10353);
or U10514 (N_10514,N_10155,N_10032);
or U10515 (N_10515,N_10027,N_10149);
nor U10516 (N_10516,N_9929,N_10014);
and U10517 (N_10517,N_10327,N_10354);
or U10518 (N_10518,N_10118,N_10065);
nor U10519 (N_10519,N_10184,N_10342);
nand U10520 (N_10520,N_10236,N_10404);
nor U10521 (N_10521,N_9930,N_9790);
xor U10522 (N_10522,N_10424,N_10000);
xnor U10523 (N_10523,N_10262,N_10072);
nor U10524 (N_10524,N_10246,N_10473);
and U10525 (N_10525,N_10080,N_9811);
nand U10526 (N_10526,N_10494,N_10281);
nand U10527 (N_10527,N_10333,N_9967);
xor U10528 (N_10528,N_10311,N_10011);
or U10529 (N_10529,N_10098,N_9938);
or U10530 (N_10530,N_9975,N_10176);
and U10531 (N_10531,N_10377,N_10356);
nor U10532 (N_10532,N_9997,N_10147);
xor U10533 (N_10533,N_10298,N_9942);
and U10534 (N_10534,N_10285,N_9796);
nand U10535 (N_10535,N_9896,N_10439);
nor U10536 (N_10536,N_9946,N_10163);
or U10537 (N_10537,N_9958,N_10470);
nor U10538 (N_10538,N_10240,N_10260);
nand U10539 (N_10539,N_9925,N_10426);
or U10540 (N_10540,N_10370,N_9950);
and U10541 (N_10541,N_10049,N_10233);
or U10542 (N_10542,N_10219,N_10195);
or U10543 (N_10543,N_10463,N_9851);
and U10544 (N_10544,N_10208,N_10096);
and U10545 (N_10545,N_9799,N_9860);
or U10546 (N_10546,N_9924,N_10466);
nand U10547 (N_10547,N_9966,N_9960);
nor U10548 (N_10548,N_10362,N_10255);
xnor U10549 (N_10549,N_10499,N_10484);
and U10550 (N_10550,N_10335,N_10472);
and U10551 (N_10551,N_9819,N_10400);
nand U10552 (N_10552,N_10074,N_9874);
nand U10553 (N_10553,N_10128,N_10086);
xor U10554 (N_10554,N_10339,N_9843);
or U10555 (N_10555,N_10073,N_10417);
nand U10556 (N_10556,N_9775,N_9913);
nand U10557 (N_10557,N_10307,N_10309);
nor U10558 (N_10558,N_9973,N_10363);
nand U10559 (N_10559,N_10067,N_10460);
and U10560 (N_10560,N_10313,N_9881);
or U10561 (N_10561,N_10197,N_10321);
nand U10562 (N_10562,N_9902,N_10413);
nor U10563 (N_10563,N_9970,N_9992);
nand U10564 (N_10564,N_10178,N_10268);
nor U10565 (N_10565,N_10475,N_10314);
and U10566 (N_10566,N_9991,N_10157);
nand U10567 (N_10567,N_10066,N_9772);
nor U10568 (N_10568,N_10398,N_9816);
nand U10569 (N_10569,N_9903,N_9858);
xor U10570 (N_10570,N_10192,N_10402);
nor U10571 (N_10571,N_9824,N_9755);
nor U10572 (N_10572,N_9797,N_9849);
nand U10573 (N_10573,N_9953,N_10312);
nor U10574 (N_10574,N_10301,N_10454);
nand U10575 (N_10575,N_10257,N_9832);
or U10576 (N_10576,N_10493,N_10133);
or U10577 (N_10577,N_10438,N_10292);
and U10578 (N_10578,N_9815,N_10266);
and U10579 (N_10579,N_9866,N_9752);
or U10580 (N_10580,N_9834,N_10267);
nor U10581 (N_10581,N_10087,N_10082);
and U10582 (N_10582,N_9994,N_10403);
xnor U10583 (N_10583,N_10289,N_9969);
nand U10584 (N_10584,N_9952,N_10319);
or U10585 (N_10585,N_9825,N_9844);
nor U10586 (N_10586,N_10084,N_9871);
and U10587 (N_10587,N_10071,N_9859);
and U10588 (N_10588,N_9919,N_9916);
and U10589 (N_10589,N_10304,N_9936);
xor U10590 (N_10590,N_10456,N_10089);
nand U10591 (N_10591,N_10044,N_10200);
or U10592 (N_10592,N_9764,N_9931);
or U10593 (N_10593,N_9898,N_10121);
and U10594 (N_10594,N_10323,N_10389);
nor U10595 (N_10595,N_10083,N_10381);
xnor U10596 (N_10596,N_10405,N_9935);
xnor U10597 (N_10597,N_9804,N_9750);
and U10598 (N_10598,N_10461,N_10177);
and U10599 (N_10599,N_10009,N_10110);
or U10600 (N_10600,N_10124,N_9761);
nand U10601 (N_10601,N_10294,N_10056);
or U10602 (N_10602,N_10416,N_10112);
nor U10603 (N_10603,N_10491,N_10085);
xor U10604 (N_10604,N_10410,N_10159);
xor U10605 (N_10605,N_9780,N_10373);
and U10606 (N_10606,N_10041,N_9959);
nor U10607 (N_10607,N_10282,N_10434);
xnor U10608 (N_10608,N_9854,N_9912);
nor U10609 (N_10609,N_10278,N_10440);
or U10610 (N_10610,N_10020,N_10395);
and U10611 (N_10611,N_10306,N_10366);
or U10612 (N_10612,N_9964,N_10308);
nand U10613 (N_10613,N_10015,N_10185);
nor U10614 (N_10614,N_10336,N_9805);
or U10615 (N_10615,N_9763,N_10069);
and U10616 (N_10616,N_9940,N_10375);
or U10617 (N_10617,N_10148,N_10430);
and U10618 (N_10618,N_10025,N_10303);
nand U10619 (N_10619,N_9830,N_10062);
xor U10620 (N_10620,N_9795,N_10419);
or U10621 (N_10621,N_10481,N_10194);
nand U10622 (N_10622,N_9949,N_9981);
nor U10623 (N_10623,N_10130,N_9888);
nor U10624 (N_10624,N_10222,N_9922);
nand U10625 (N_10625,N_10038,N_9899);
and U10626 (N_10626,N_10120,N_10145);
xor U10627 (N_10627,N_10190,N_9754);
and U10628 (N_10628,N_10253,N_10106);
nand U10629 (N_10629,N_10443,N_10490);
and U10630 (N_10630,N_10227,N_10181);
or U10631 (N_10631,N_9789,N_10427);
and U10632 (N_10632,N_9901,N_9999);
nor U10633 (N_10633,N_9769,N_10302);
nand U10634 (N_10634,N_10168,N_10094);
nor U10635 (N_10635,N_10226,N_9788);
nor U10636 (N_10636,N_9822,N_9996);
xor U10637 (N_10637,N_10088,N_10012);
nand U10638 (N_10638,N_10483,N_9883);
nor U10639 (N_10639,N_10437,N_10391);
nand U10640 (N_10640,N_9890,N_10035);
or U10641 (N_10641,N_9873,N_9777);
xnor U10642 (N_10642,N_9986,N_10407);
nand U10643 (N_10643,N_10414,N_10379);
and U10644 (N_10644,N_10230,N_10093);
and U10645 (N_10645,N_10330,N_10068);
or U10646 (N_10646,N_10175,N_10408);
nor U10647 (N_10647,N_10270,N_10114);
and U10648 (N_10648,N_9794,N_9932);
nand U10649 (N_10649,N_10052,N_9906);
or U10650 (N_10650,N_9918,N_10248);
nor U10651 (N_10651,N_10325,N_10468);
nor U10652 (N_10652,N_10397,N_10209);
xnor U10653 (N_10653,N_9846,N_10001);
nand U10654 (N_10654,N_10228,N_9965);
nor U10655 (N_10655,N_10210,N_10450);
nor U10656 (N_10656,N_10164,N_10345);
nand U10657 (N_10657,N_9884,N_9878);
or U10658 (N_10658,N_10191,N_10256);
nor U10659 (N_10659,N_9869,N_10057);
or U10660 (N_10660,N_10316,N_10154);
and U10661 (N_10661,N_9827,N_9993);
xor U10662 (N_10662,N_10299,N_10105);
or U10663 (N_10663,N_9765,N_10347);
nand U10664 (N_10664,N_9882,N_10421);
and U10665 (N_10665,N_10205,N_10351);
xor U10666 (N_10666,N_10077,N_9855);
or U10667 (N_10667,N_9886,N_10007);
nand U10668 (N_10668,N_10271,N_10261);
nor U10669 (N_10669,N_10406,N_9998);
nand U10670 (N_10670,N_9809,N_10127);
nand U10671 (N_10671,N_9892,N_10445);
xor U10672 (N_10672,N_9864,N_9785);
nor U10673 (N_10673,N_9900,N_9910);
or U10674 (N_10674,N_10331,N_10305);
nor U10675 (N_10675,N_10295,N_10064);
and U10676 (N_10676,N_9753,N_10103);
nand U10677 (N_10677,N_10097,N_10396);
nor U10678 (N_10678,N_9792,N_9826);
or U10679 (N_10679,N_10040,N_9856);
nor U10680 (N_10680,N_10346,N_9823);
and U10681 (N_10681,N_9927,N_9894);
and U10682 (N_10682,N_10425,N_9852);
nand U10683 (N_10683,N_10182,N_10029);
nor U10684 (N_10684,N_10109,N_10360);
and U10685 (N_10685,N_10388,N_9984);
xnor U10686 (N_10686,N_10435,N_9814);
nor U10687 (N_10687,N_9982,N_10171);
xor U10688 (N_10688,N_10247,N_9872);
nor U10689 (N_10689,N_9939,N_10348);
xnor U10690 (N_10690,N_10265,N_9870);
and U10691 (N_10691,N_9955,N_10287);
xor U10692 (N_10692,N_10174,N_10497);
and U10693 (N_10693,N_10075,N_10030);
nor U10694 (N_10694,N_10022,N_10196);
nand U10695 (N_10695,N_10367,N_10100);
nor U10696 (N_10696,N_9914,N_10179);
nor U10697 (N_10697,N_9808,N_10245);
nand U10698 (N_10698,N_10252,N_10169);
nand U10699 (N_10699,N_10477,N_10051);
and U10700 (N_10700,N_10018,N_10368);
and U10701 (N_10701,N_10047,N_9787);
or U10702 (N_10702,N_10144,N_10392);
xnor U10703 (N_10703,N_10412,N_9968);
nand U10704 (N_10704,N_9836,N_10172);
xor U10705 (N_10705,N_10332,N_10183);
or U10706 (N_10706,N_9778,N_10250);
nor U10707 (N_10707,N_10315,N_9956);
nand U10708 (N_10708,N_10320,N_10409);
and U10709 (N_10709,N_10272,N_10277);
and U10710 (N_10710,N_10070,N_9756);
or U10711 (N_10711,N_9776,N_10214);
xnor U10712 (N_10712,N_10037,N_10188);
or U10713 (N_10713,N_10199,N_10283);
xnor U10714 (N_10714,N_9865,N_10079);
or U10715 (N_10715,N_10126,N_10386);
and U10716 (N_10716,N_10170,N_10476);
nand U10717 (N_10717,N_10341,N_10310);
and U10718 (N_10718,N_10153,N_10152);
or U10719 (N_10719,N_10165,N_10193);
and U10720 (N_10720,N_10486,N_10137);
and U10721 (N_10721,N_10166,N_10223);
nor U10722 (N_10722,N_9782,N_10053);
nand U10723 (N_10723,N_10213,N_9909);
nor U10724 (N_10724,N_9798,N_10150);
and U10725 (N_10725,N_9897,N_10431);
and U10726 (N_10726,N_10420,N_10384);
nand U10727 (N_10727,N_10487,N_9926);
xor U10728 (N_10728,N_10048,N_10198);
or U10729 (N_10729,N_10436,N_10429);
or U10730 (N_10730,N_10369,N_9760);
or U10731 (N_10731,N_9905,N_9977);
nand U10732 (N_10732,N_9880,N_10116);
xnor U10733 (N_10733,N_10374,N_9850);
and U10734 (N_10734,N_9766,N_10350);
nand U10735 (N_10735,N_9885,N_9895);
and U10736 (N_10736,N_10016,N_9944);
nor U10737 (N_10737,N_10274,N_9838);
nand U10738 (N_10738,N_9862,N_10344);
nand U10739 (N_10739,N_10258,N_10474);
or U10740 (N_10740,N_10146,N_9820);
nor U10741 (N_10741,N_9893,N_9813);
nand U10742 (N_10742,N_10269,N_9793);
nor U10743 (N_10743,N_10099,N_10390);
nor U10744 (N_10744,N_10338,N_9784);
or U10745 (N_10745,N_9971,N_9781);
or U10746 (N_10746,N_9947,N_10156);
or U10747 (N_10747,N_10232,N_10365);
nand U10748 (N_10748,N_10275,N_10288);
xor U10749 (N_10749,N_9861,N_10091);
xnor U10750 (N_10750,N_10102,N_10031);
nand U10751 (N_10751,N_10054,N_9875);
nand U10752 (N_10752,N_9801,N_9907);
xnor U10753 (N_10753,N_10061,N_10151);
xnor U10754 (N_10754,N_9941,N_10076);
xor U10755 (N_10755,N_10143,N_10024);
and U10756 (N_10756,N_10382,N_9933);
or U10757 (N_10757,N_9779,N_9948);
and U10758 (N_10758,N_9770,N_10212);
xnor U10759 (N_10759,N_10286,N_10393);
nor U10760 (N_10760,N_10058,N_10224);
xor U10761 (N_10761,N_9983,N_10115);
nor U10762 (N_10762,N_10081,N_10415);
nor U10763 (N_10763,N_10385,N_10036);
or U10764 (N_10764,N_9945,N_10092);
xor U10765 (N_10765,N_10432,N_9767);
nor U10766 (N_10766,N_9980,N_9877);
and U10767 (N_10767,N_10485,N_9847);
xor U10768 (N_10768,N_9803,N_10394);
and U10769 (N_10769,N_9802,N_9995);
and U10770 (N_10770,N_10447,N_9937);
or U10771 (N_10771,N_10111,N_10372);
nand U10772 (N_10772,N_10162,N_9887);
nor U10773 (N_10773,N_10167,N_10488);
or U10774 (N_10774,N_10008,N_10465);
and U10775 (N_10775,N_10448,N_9868);
nand U10776 (N_10776,N_10234,N_9821);
xnor U10777 (N_10777,N_10003,N_10441);
nand U10778 (N_10778,N_9943,N_10376);
xnor U10779 (N_10779,N_10482,N_10129);
and U10780 (N_10780,N_10423,N_10019);
and U10781 (N_10781,N_10383,N_10279);
nand U10782 (N_10782,N_9915,N_9920);
xor U10783 (N_10783,N_10358,N_10471);
nand U10784 (N_10784,N_10023,N_10211);
or U10785 (N_10785,N_10055,N_9976);
and U10786 (N_10786,N_10340,N_10050);
xor U10787 (N_10787,N_10229,N_9957);
nand U10788 (N_10788,N_9891,N_9974);
xor U10789 (N_10789,N_10293,N_10043);
nand U10790 (N_10790,N_10095,N_10203);
or U10791 (N_10791,N_10280,N_10122);
and U10792 (N_10792,N_10002,N_10489);
or U10793 (N_10793,N_9985,N_10242);
nand U10794 (N_10794,N_9833,N_10459);
and U10795 (N_10795,N_10378,N_9989);
nand U10796 (N_10796,N_10238,N_9800);
nor U10797 (N_10797,N_10207,N_10158);
or U10798 (N_10798,N_10453,N_10276);
nand U10799 (N_10799,N_9876,N_9786);
nand U10800 (N_10800,N_9759,N_10254);
or U10801 (N_10801,N_10428,N_9921);
nor U10802 (N_10802,N_9839,N_10467);
nand U10803 (N_10803,N_10249,N_10399);
or U10804 (N_10804,N_10411,N_9963);
or U10805 (N_10805,N_10297,N_10101);
and U10806 (N_10806,N_10123,N_10464);
xnor U10807 (N_10807,N_9951,N_9863);
or U10808 (N_10808,N_10218,N_10187);
xor U10809 (N_10809,N_10140,N_10478);
xor U10810 (N_10810,N_10433,N_10161);
nor U10811 (N_10811,N_9908,N_10215);
and U10812 (N_10812,N_9879,N_10131);
and U10813 (N_10813,N_9757,N_9988);
and U10814 (N_10814,N_10479,N_9829);
nor U10815 (N_10815,N_10042,N_9867);
nor U10816 (N_10816,N_10469,N_10141);
nor U10817 (N_10817,N_9768,N_9954);
nor U10818 (N_10818,N_9990,N_9773);
or U10819 (N_10819,N_10349,N_10021);
nor U10820 (N_10820,N_10216,N_10446);
nor U10821 (N_10821,N_9857,N_10401);
nor U10822 (N_10822,N_10217,N_10013);
and U10823 (N_10823,N_10180,N_10005);
nor U10824 (N_10824,N_10136,N_10026);
nor U10825 (N_10825,N_10142,N_10273);
and U10826 (N_10826,N_10045,N_10359);
or U10827 (N_10827,N_10455,N_10119);
and U10828 (N_10828,N_10034,N_10039);
or U10829 (N_10829,N_9928,N_9783);
xnor U10830 (N_10830,N_9791,N_10004);
or U10831 (N_10831,N_10496,N_10259);
nor U10832 (N_10832,N_10387,N_10006);
nand U10833 (N_10833,N_10204,N_10296);
xnor U10834 (N_10834,N_10201,N_10113);
nand U10835 (N_10835,N_9853,N_9758);
or U10836 (N_10836,N_10244,N_10059);
or U10837 (N_10837,N_10371,N_10017);
nand U10838 (N_10838,N_10189,N_10139);
nor U10839 (N_10839,N_9978,N_10221);
nand U10840 (N_10840,N_10352,N_10290);
nor U10841 (N_10841,N_10492,N_10173);
nand U10842 (N_10842,N_10033,N_9842);
nand U10843 (N_10843,N_10452,N_10284);
and U10844 (N_10844,N_9831,N_9845);
nor U10845 (N_10845,N_10324,N_10355);
nand U10846 (N_10846,N_9771,N_9841);
nand U10847 (N_10847,N_10462,N_10343);
and U10848 (N_10848,N_9979,N_9889);
xnor U10849 (N_10849,N_9917,N_10326);
and U10850 (N_10850,N_10251,N_10328);
and U10851 (N_10851,N_10108,N_9848);
xnor U10852 (N_10852,N_9751,N_10125);
nor U10853 (N_10853,N_10291,N_10334);
nor U10854 (N_10854,N_10317,N_10138);
and U10855 (N_10855,N_10422,N_9762);
xor U10856 (N_10856,N_10135,N_10318);
nand U10857 (N_10857,N_9962,N_9961);
or U10858 (N_10858,N_10480,N_10263);
xor U10859 (N_10859,N_9923,N_9810);
nand U10860 (N_10860,N_10442,N_10264);
nand U10861 (N_10861,N_10364,N_10458);
nor U10862 (N_10862,N_10361,N_10418);
or U10863 (N_10863,N_9806,N_10457);
or U10864 (N_10864,N_10220,N_10107);
or U10865 (N_10865,N_10134,N_10495);
or U10866 (N_10866,N_10241,N_10010);
nand U10867 (N_10867,N_10117,N_10132);
nand U10868 (N_10868,N_10186,N_9817);
nor U10869 (N_10869,N_10206,N_9972);
or U10870 (N_10870,N_10237,N_10090);
and U10871 (N_10871,N_10063,N_10337);
nor U10872 (N_10872,N_10451,N_9818);
xor U10873 (N_10873,N_10235,N_10078);
xnor U10874 (N_10874,N_9837,N_9911);
xnor U10875 (N_10875,N_10132,N_10454);
nor U10876 (N_10876,N_9916,N_9751);
xor U10877 (N_10877,N_10158,N_10475);
and U10878 (N_10878,N_10480,N_10441);
nand U10879 (N_10879,N_10012,N_9851);
nor U10880 (N_10880,N_9983,N_10048);
or U10881 (N_10881,N_9976,N_9802);
nand U10882 (N_10882,N_9986,N_10119);
and U10883 (N_10883,N_10274,N_10099);
or U10884 (N_10884,N_10106,N_10206);
and U10885 (N_10885,N_9826,N_10377);
or U10886 (N_10886,N_10229,N_9823);
xnor U10887 (N_10887,N_9868,N_10174);
or U10888 (N_10888,N_9930,N_9942);
or U10889 (N_10889,N_10399,N_9898);
and U10890 (N_10890,N_10244,N_9800);
xor U10891 (N_10891,N_10339,N_10312);
and U10892 (N_10892,N_9958,N_10339);
xor U10893 (N_10893,N_10365,N_10076);
and U10894 (N_10894,N_10100,N_9820);
or U10895 (N_10895,N_10051,N_10332);
and U10896 (N_10896,N_10398,N_10493);
nor U10897 (N_10897,N_9968,N_10152);
nor U10898 (N_10898,N_10245,N_10392);
xnor U10899 (N_10899,N_10292,N_10167);
nand U10900 (N_10900,N_10136,N_10355);
nor U10901 (N_10901,N_10407,N_9751);
nand U10902 (N_10902,N_10146,N_10151);
nand U10903 (N_10903,N_10445,N_10077);
nor U10904 (N_10904,N_9838,N_9925);
or U10905 (N_10905,N_10017,N_9755);
or U10906 (N_10906,N_10453,N_10430);
or U10907 (N_10907,N_9844,N_10248);
nor U10908 (N_10908,N_10372,N_10046);
nor U10909 (N_10909,N_10318,N_10413);
nand U10910 (N_10910,N_10181,N_10046);
nand U10911 (N_10911,N_10181,N_9960);
and U10912 (N_10912,N_9787,N_10182);
nand U10913 (N_10913,N_10149,N_9764);
nand U10914 (N_10914,N_10288,N_10341);
or U10915 (N_10915,N_10455,N_10037);
nand U10916 (N_10916,N_10025,N_10461);
nand U10917 (N_10917,N_10134,N_10459);
and U10918 (N_10918,N_10108,N_10112);
and U10919 (N_10919,N_9930,N_10013);
or U10920 (N_10920,N_10200,N_10239);
xnor U10921 (N_10921,N_10209,N_10164);
nor U10922 (N_10922,N_9869,N_10073);
or U10923 (N_10923,N_10350,N_10316);
or U10924 (N_10924,N_10248,N_10031);
nor U10925 (N_10925,N_10010,N_10329);
or U10926 (N_10926,N_9879,N_10210);
and U10927 (N_10927,N_10245,N_10469);
and U10928 (N_10928,N_10022,N_10452);
and U10929 (N_10929,N_9876,N_10316);
nand U10930 (N_10930,N_10071,N_10323);
xnor U10931 (N_10931,N_10459,N_10004);
xnor U10932 (N_10932,N_9917,N_9998);
nor U10933 (N_10933,N_10319,N_10317);
nand U10934 (N_10934,N_10428,N_10160);
nor U10935 (N_10935,N_10076,N_10402);
nand U10936 (N_10936,N_10339,N_10427);
nor U10937 (N_10937,N_10234,N_10157);
or U10938 (N_10938,N_10250,N_10046);
nor U10939 (N_10939,N_10219,N_9973);
and U10940 (N_10940,N_9816,N_9780);
nand U10941 (N_10941,N_10486,N_10253);
and U10942 (N_10942,N_10342,N_9995);
nand U10943 (N_10943,N_10197,N_10176);
and U10944 (N_10944,N_9887,N_10224);
or U10945 (N_10945,N_10431,N_9952);
xor U10946 (N_10946,N_9756,N_9871);
or U10947 (N_10947,N_10275,N_9826);
xor U10948 (N_10948,N_10188,N_10280);
nor U10949 (N_10949,N_10003,N_10135);
and U10950 (N_10950,N_10123,N_9882);
xnor U10951 (N_10951,N_10147,N_10171);
or U10952 (N_10952,N_10183,N_10320);
and U10953 (N_10953,N_10079,N_9901);
and U10954 (N_10954,N_9927,N_10448);
and U10955 (N_10955,N_10319,N_10042);
nand U10956 (N_10956,N_10392,N_10460);
nand U10957 (N_10957,N_10336,N_10206);
xor U10958 (N_10958,N_9955,N_10046);
xor U10959 (N_10959,N_10469,N_10169);
nand U10960 (N_10960,N_10269,N_9841);
or U10961 (N_10961,N_9994,N_9968);
nor U10962 (N_10962,N_10110,N_10361);
nand U10963 (N_10963,N_9942,N_9815);
xnor U10964 (N_10964,N_9840,N_9933);
and U10965 (N_10965,N_10039,N_9930);
and U10966 (N_10966,N_9905,N_10440);
xor U10967 (N_10967,N_10476,N_9944);
xnor U10968 (N_10968,N_9934,N_10156);
or U10969 (N_10969,N_10371,N_9828);
nand U10970 (N_10970,N_10463,N_9787);
xnor U10971 (N_10971,N_10343,N_10442);
and U10972 (N_10972,N_10498,N_10461);
nor U10973 (N_10973,N_9837,N_10177);
nor U10974 (N_10974,N_10278,N_10150);
nand U10975 (N_10975,N_9936,N_10227);
or U10976 (N_10976,N_10367,N_10000);
nand U10977 (N_10977,N_10486,N_10316);
or U10978 (N_10978,N_9955,N_10424);
and U10979 (N_10979,N_10230,N_10136);
and U10980 (N_10980,N_10493,N_10323);
nor U10981 (N_10981,N_9907,N_10294);
nand U10982 (N_10982,N_10422,N_9879);
nand U10983 (N_10983,N_9817,N_10091);
nand U10984 (N_10984,N_10149,N_10068);
xor U10985 (N_10985,N_9820,N_10159);
or U10986 (N_10986,N_10088,N_10363);
nor U10987 (N_10987,N_10494,N_10311);
xnor U10988 (N_10988,N_10193,N_10172);
nand U10989 (N_10989,N_9929,N_9783);
nand U10990 (N_10990,N_10278,N_9791);
xor U10991 (N_10991,N_10313,N_9784);
nor U10992 (N_10992,N_10014,N_9848);
or U10993 (N_10993,N_9956,N_10303);
xnor U10994 (N_10994,N_9922,N_10088);
xnor U10995 (N_10995,N_10225,N_10431);
or U10996 (N_10996,N_10144,N_10418);
nand U10997 (N_10997,N_9948,N_10484);
xor U10998 (N_10998,N_9754,N_9815);
or U10999 (N_10999,N_10342,N_9990);
nor U11000 (N_11000,N_10266,N_9838);
nand U11001 (N_11001,N_10380,N_10434);
nor U11002 (N_11002,N_10241,N_10165);
nand U11003 (N_11003,N_10366,N_10192);
and U11004 (N_11004,N_9917,N_10341);
and U11005 (N_11005,N_10038,N_9853);
and U11006 (N_11006,N_9949,N_9954);
and U11007 (N_11007,N_10397,N_10384);
and U11008 (N_11008,N_9827,N_9846);
and U11009 (N_11009,N_10293,N_9816);
or U11010 (N_11010,N_9873,N_9791);
nand U11011 (N_11011,N_10163,N_9908);
nand U11012 (N_11012,N_10218,N_10109);
and U11013 (N_11013,N_9857,N_10101);
and U11014 (N_11014,N_10292,N_10082);
nand U11015 (N_11015,N_10393,N_9949);
xnor U11016 (N_11016,N_10404,N_10290);
xor U11017 (N_11017,N_10263,N_9978);
nand U11018 (N_11018,N_9867,N_10459);
xor U11019 (N_11019,N_10266,N_10310);
and U11020 (N_11020,N_10464,N_10074);
nand U11021 (N_11021,N_10014,N_10192);
nand U11022 (N_11022,N_10437,N_9954);
and U11023 (N_11023,N_10029,N_10020);
nor U11024 (N_11024,N_10410,N_9866);
xnor U11025 (N_11025,N_10027,N_9818);
nand U11026 (N_11026,N_10077,N_10251);
or U11027 (N_11027,N_9877,N_10463);
and U11028 (N_11028,N_9768,N_9763);
nor U11029 (N_11029,N_9804,N_10168);
or U11030 (N_11030,N_10125,N_10101);
nor U11031 (N_11031,N_9940,N_10145);
xor U11032 (N_11032,N_9866,N_9996);
and U11033 (N_11033,N_10462,N_9817);
nor U11034 (N_11034,N_9825,N_9837);
and U11035 (N_11035,N_10219,N_10057);
nand U11036 (N_11036,N_10242,N_10382);
nor U11037 (N_11037,N_10007,N_10258);
nor U11038 (N_11038,N_10134,N_9978);
nand U11039 (N_11039,N_9817,N_9895);
nand U11040 (N_11040,N_9998,N_9939);
nand U11041 (N_11041,N_9935,N_10156);
or U11042 (N_11042,N_9958,N_9819);
and U11043 (N_11043,N_10491,N_10271);
nor U11044 (N_11044,N_10270,N_10381);
and U11045 (N_11045,N_10151,N_10197);
and U11046 (N_11046,N_10210,N_10370);
nand U11047 (N_11047,N_9760,N_10143);
or U11048 (N_11048,N_9768,N_10481);
nand U11049 (N_11049,N_10236,N_10093);
nor U11050 (N_11050,N_10000,N_9815);
nor U11051 (N_11051,N_9956,N_10086);
nand U11052 (N_11052,N_9772,N_10255);
and U11053 (N_11053,N_10266,N_9908);
and U11054 (N_11054,N_10084,N_10203);
nor U11055 (N_11055,N_9923,N_10432);
or U11056 (N_11056,N_10096,N_9980);
or U11057 (N_11057,N_10465,N_10078);
or U11058 (N_11058,N_9802,N_9935);
and U11059 (N_11059,N_10344,N_9864);
xor U11060 (N_11060,N_10263,N_9997);
nor U11061 (N_11061,N_9815,N_9854);
nand U11062 (N_11062,N_10049,N_10294);
nor U11063 (N_11063,N_10068,N_10475);
xor U11064 (N_11064,N_9983,N_10164);
xor U11065 (N_11065,N_10434,N_10128);
and U11066 (N_11066,N_10130,N_10267);
and U11067 (N_11067,N_9807,N_10444);
nand U11068 (N_11068,N_10497,N_10335);
or U11069 (N_11069,N_10167,N_10350);
nor U11070 (N_11070,N_10315,N_10337);
and U11071 (N_11071,N_9896,N_9966);
or U11072 (N_11072,N_10356,N_10274);
xor U11073 (N_11073,N_10236,N_9837);
and U11074 (N_11074,N_10476,N_10276);
xnor U11075 (N_11075,N_10155,N_9979);
or U11076 (N_11076,N_9798,N_10418);
xor U11077 (N_11077,N_9859,N_9831);
nor U11078 (N_11078,N_9894,N_9852);
nand U11079 (N_11079,N_10114,N_9940);
nor U11080 (N_11080,N_10365,N_9930);
and U11081 (N_11081,N_10211,N_10294);
nand U11082 (N_11082,N_9864,N_10303);
nor U11083 (N_11083,N_10283,N_10295);
and U11084 (N_11084,N_9796,N_10122);
xnor U11085 (N_11085,N_10459,N_10119);
and U11086 (N_11086,N_10119,N_10431);
and U11087 (N_11087,N_10122,N_9988);
xor U11088 (N_11088,N_10071,N_10208);
and U11089 (N_11089,N_9926,N_10090);
nand U11090 (N_11090,N_10313,N_10443);
and U11091 (N_11091,N_10363,N_10158);
xor U11092 (N_11092,N_10032,N_9873);
xor U11093 (N_11093,N_10120,N_9981);
or U11094 (N_11094,N_9928,N_10205);
nand U11095 (N_11095,N_10048,N_10143);
or U11096 (N_11096,N_9757,N_10114);
xor U11097 (N_11097,N_10345,N_10114);
xnor U11098 (N_11098,N_10371,N_10427);
or U11099 (N_11099,N_10142,N_10356);
and U11100 (N_11100,N_10159,N_10102);
nand U11101 (N_11101,N_10354,N_10439);
nand U11102 (N_11102,N_10083,N_10298);
nand U11103 (N_11103,N_9906,N_9943);
nand U11104 (N_11104,N_10055,N_10130);
and U11105 (N_11105,N_10487,N_10474);
and U11106 (N_11106,N_9806,N_9871);
or U11107 (N_11107,N_9803,N_10279);
or U11108 (N_11108,N_10052,N_10491);
nor U11109 (N_11109,N_10488,N_10293);
or U11110 (N_11110,N_10029,N_9827);
and U11111 (N_11111,N_10208,N_10154);
or U11112 (N_11112,N_10084,N_9860);
xor U11113 (N_11113,N_10174,N_10377);
and U11114 (N_11114,N_9866,N_9870);
nand U11115 (N_11115,N_9750,N_10007);
xor U11116 (N_11116,N_10288,N_10228);
nor U11117 (N_11117,N_9788,N_9996);
xor U11118 (N_11118,N_10102,N_10426);
and U11119 (N_11119,N_10222,N_9882);
or U11120 (N_11120,N_10175,N_9854);
nor U11121 (N_11121,N_9756,N_10379);
and U11122 (N_11122,N_10249,N_10201);
nor U11123 (N_11123,N_9879,N_10086);
xor U11124 (N_11124,N_10219,N_9787);
xnor U11125 (N_11125,N_10497,N_10470);
nand U11126 (N_11126,N_10221,N_9852);
nand U11127 (N_11127,N_10446,N_10401);
nand U11128 (N_11128,N_10157,N_10097);
nor U11129 (N_11129,N_10200,N_9941);
or U11130 (N_11130,N_10142,N_9939);
nand U11131 (N_11131,N_9860,N_9753);
nand U11132 (N_11132,N_10387,N_9949);
and U11133 (N_11133,N_9969,N_10092);
or U11134 (N_11134,N_10040,N_10260);
xnor U11135 (N_11135,N_10031,N_10357);
nor U11136 (N_11136,N_9843,N_10446);
nor U11137 (N_11137,N_9840,N_10209);
or U11138 (N_11138,N_9868,N_10207);
nand U11139 (N_11139,N_10265,N_10475);
and U11140 (N_11140,N_9839,N_10278);
xnor U11141 (N_11141,N_9805,N_10164);
or U11142 (N_11142,N_9879,N_9873);
and U11143 (N_11143,N_9991,N_10016);
and U11144 (N_11144,N_10485,N_10492);
or U11145 (N_11145,N_9772,N_9910);
nor U11146 (N_11146,N_9861,N_10295);
or U11147 (N_11147,N_10163,N_10174);
or U11148 (N_11148,N_9904,N_9818);
and U11149 (N_11149,N_9777,N_10350);
nor U11150 (N_11150,N_10478,N_9796);
or U11151 (N_11151,N_10329,N_10004);
and U11152 (N_11152,N_9762,N_9892);
and U11153 (N_11153,N_10303,N_10068);
or U11154 (N_11154,N_10333,N_10219);
xnor U11155 (N_11155,N_10216,N_9861);
xor U11156 (N_11156,N_10013,N_10117);
nand U11157 (N_11157,N_10191,N_10469);
or U11158 (N_11158,N_10238,N_9956);
or U11159 (N_11159,N_10489,N_10343);
nor U11160 (N_11160,N_9840,N_10297);
nand U11161 (N_11161,N_10113,N_9817);
xnor U11162 (N_11162,N_10023,N_9846);
xnor U11163 (N_11163,N_9801,N_9999);
or U11164 (N_11164,N_10159,N_10493);
nor U11165 (N_11165,N_10277,N_9877);
nor U11166 (N_11166,N_9917,N_9898);
nor U11167 (N_11167,N_9759,N_10382);
nand U11168 (N_11168,N_9795,N_10175);
nor U11169 (N_11169,N_9999,N_9979);
xnor U11170 (N_11170,N_10357,N_10113);
or U11171 (N_11171,N_9836,N_10372);
nor U11172 (N_11172,N_10064,N_10246);
xor U11173 (N_11173,N_10373,N_10383);
or U11174 (N_11174,N_10047,N_10409);
and U11175 (N_11175,N_9865,N_10483);
nand U11176 (N_11176,N_9852,N_10093);
nand U11177 (N_11177,N_10024,N_9832);
nor U11178 (N_11178,N_10308,N_10247);
xnor U11179 (N_11179,N_10217,N_9819);
nor U11180 (N_11180,N_10478,N_9829);
xnor U11181 (N_11181,N_10170,N_10111);
xnor U11182 (N_11182,N_10364,N_9939);
xnor U11183 (N_11183,N_10478,N_10303);
and U11184 (N_11184,N_9750,N_9902);
nand U11185 (N_11185,N_9781,N_9964);
nand U11186 (N_11186,N_10308,N_9979);
and U11187 (N_11187,N_10004,N_10048);
xor U11188 (N_11188,N_10059,N_10344);
xor U11189 (N_11189,N_10242,N_10490);
xnor U11190 (N_11190,N_10043,N_9939);
xnor U11191 (N_11191,N_10193,N_9890);
or U11192 (N_11192,N_10029,N_9904);
and U11193 (N_11193,N_10166,N_10274);
or U11194 (N_11194,N_10409,N_9983);
nand U11195 (N_11195,N_10455,N_10189);
nand U11196 (N_11196,N_10190,N_10473);
and U11197 (N_11197,N_9867,N_10021);
xor U11198 (N_11198,N_10101,N_9958);
xnor U11199 (N_11199,N_9889,N_10194);
xnor U11200 (N_11200,N_9764,N_10389);
or U11201 (N_11201,N_10012,N_9916);
nor U11202 (N_11202,N_10254,N_10497);
xor U11203 (N_11203,N_10161,N_9913);
and U11204 (N_11204,N_10368,N_10056);
nand U11205 (N_11205,N_10455,N_9874);
nand U11206 (N_11206,N_10052,N_9813);
xor U11207 (N_11207,N_9949,N_9940);
nand U11208 (N_11208,N_10410,N_10379);
or U11209 (N_11209,N_10420,N_10189);
xnor U11210 (N_11210,N_10251,N_10049);
and U11211 (N_11211,N_10043,N_10036);
and U11212 (N_11212,N_10387,N_10448);
and U11213 (N_11213,N_9958,N_10485);
and U11214 (N_11214,N_10165,N_9894);
nor U11215 (N_11215,N_9825,N_10164);
nand U11216 (N_11216,N_10168,N_9862);
and U11217 (N_11217,N_9799,N_10043);
xnor U11218 (N_11218,N_9753,N_9950);
nor U11219 (N_11219,N_10126,N_10051);
xnor U11220 (N_11220,N_10182,N_9823);
or U11221 (N_11221,N_10411,N_10299);
or U11222 (N_11222,N_9798,N_10011);
nor U11223 (N_11223,N_9997,N_9972);
xor U11224 (N_11224,N_10162,N_10323);
and U11225 (N_11225,N_9787,N_9783);
and U11226 (N_11226,N_10116,N_10402);
and U11227 (N_11227,N_10207,N_10338);
xor U11228 (N_11228,N_9753,N_10299);
and U11229 (N_11229,N_10431,N_10149);
or U11230 (N_11230,N_9774,N_9945);
xor U11231 (N_11231,N_9857,N_10037);
nand U11232 (N_11232,N_10330,N_9826);
nand U11233 (N_11233,N_10171,N_9825);
xor U11234 (N_11234,N_9755,N_10380);
and U11235 (N_11235,N_10263,N_10301);
or U11236 (N_11236,N_10469,N_10453);
xor U11237 (N_11237,N_9927,N_10477);
nor U11238 (N_11238,N_9955,N_10435);
xnor U11239 (N_11239,N_10388,N_10210);
nand U11240 (N_11240,N_9750,N_10449);
nand U11241 (N_11241,N_9862,N_10297);
xor U11242 (N_11242,N_10258,N_10154);
nand U11243 (N_11243,N_10196,N_10429);
or U11244 (N_11244,N_9892,N_10082);
nor U11245 (N_11245,N_10197,N_9835);
or U11246 (N_11246,N_10240,N_9897);
xor U11247 (N_11247,N_10052,N_10153);
nor U11248 (N_11248,N_10314,N_10147);
nand U11249 (N_11249,N_9786,N_10400);
or U11250 (N_11250,N_10785,N_11238);
nor U11251 (N_11251,N_10717,N_10938);
or U11252 (N_11252,N_10862,N_10823);
xor U11253 (N_11253,N_11051,N_10536);
xnor U11254 (N_11254,N_10657,N_11185);
nor U11255 (N_11255,N_10602,N_10550);
or U11256 (N_11256,N_10836,N_11093);
or U11257 (N_11257,N_11079,N_10746);
xnor U11258 (N_11258,N_10666,N_10560);
nor U11259 (N_11259,N_10669,N_10813);
xnor U11260 (N_11260,N_10769,N_10854);
xnor U11261 (N_11261,N_10936,N_11186);
xnor U11262 (N_11262,N_11031,N_10719);
xnor U11263 (N_11263,N_10696,N_10502);
xnor U11264 (N_11264,N_10538,N_10601);
nand U11265 (N_11265,N_11157,N_10868);
xnor U11266 (N_11266,N_11010,N_10688);
nand U11267 (N_11267,N_10874,N_11043);
xor U11268 (N_11268,N_10807,N_11170);
nor U11269 (N_11269,N_11022,N_10737);
nand U11270 (N_11270,N_10681,N_11064);
xor U11271 (N_11271,N_10768,N_11182);
and U11272 (N_11272,N_11129,N_10610);
or U11273 (N_11273,N_11040,N_10570);
nand U11274 (N_11274,N_10912,N_11008);
xor U11275 (N_11275,N_10950,N_10526);
nor U11276 (N_11276,N_11023,N_11132);
nand U11277 (N_11277,N_10900,N_10662);
and U11278 (N_11278,N_11071,N_10604);
nand U11279 (N_11279,N_10791,N_10953);
and U11280 (N_11280,N_11004,N_10845);
nor U11281 (N_11281,N_10521,N_10996);
or U11282 (N_11282,N_10647,N_10650);
nand U11283 (N_11283,N_10642,N_10545);
nand U11284 (N_11284,N_10920,N_10815);
nor U11285 (N_11285,N_11111,N_10588);
and U11286 (N_11286,N_10529,N_10629);
xor U11287 (N_11287,N_10742,N_10562);
nand U11288 (N_11288,N_11224,N_11136);
xor U11289 (N_11289,N_10584,N_10625);
nor U11290 (N_11290,N_10730,N_11065);
xor U11291 (N_11291,N_11125,N_10693);
or U11292 (N_11292,N_11037,N_10672);
nand U11293 (N_11293,N_10922,N_11137);
nand U11294 (N_11294,N_11141,N_10827);
nand U11295 (N_11295,N_10598,N_10821);
or U11296 (N_11296,N_10853,N_10665);
nand U11297 (N_11297,N_10701,N_10964);
nand U11298 (N_11298,N_10939,N_11124);
nand U11299 (N_11299,N_11200,N_11147);
and U11300 (N_11300,N_10962,N_11122);
nor U11301 (N_11301,N_10524,N_10776);
nor U11302 (N_11302,N_10808,N_11116);
and U11303 (N_11303,N_11095,N_11001);
xor U11304 (N_11304,N_10937,N_10978);
and U11305 (N_11305,N_10990,N_10794);
and U11306 (N_11306,N_10704,N_11107);
and U11307 (N_11307,N_10613,N_11167);
nand U11308 (N_11308,N_11187,N_10885);
nor U11309 (N_11309,N_10555,N_11068);
and U11310 (N_11310,N_11056,N_10979);
xor U11311 (N_11311,N_10606,N_11081);
nand U11312 (N_11312,N_11102,N_10508);
or U11313 (N_11313,N_10914,N_11180);
or U11314 (N_11314,N_10582,N_11015);
and U11315 (N_11315,N_10822,N_10585);
and U11316 (N_11316,N_11208,N_10563);
or U11317 (N_11317,N_10987,N_11154);
and U11318 (N_11318,N_10576,N_11127);
xnor U11319 (N_11319,N_10965,N_10879);
nand U11320 (N_11320,N_10590,N_11084);
xor U11321 (N_11321,N_11087,N_10773);
nand U11322 (N_11322,N_10787,N_10556);
xnor U11323 (N_11323,N_10675,N_10631);
or U11324 (N_11324,N_10649,N_10852);
xnor U11325 (N_11325,N_11097,N_10680);
or U11326 (N_11326,N_10851,N_10795);
or U11327 (N_11327,N_10518,N_10640);
or U11328 (N_11328,N_10998,N_10933);
xnor U11329 (N_11329,N_10744,N_11126);
or U11330 (N_11330,N_11235,N_11233);
and U11331 (N_11331,N_10715,N_10617);
or U11332 (N_11332,N_10857,N_10739);
xnor U11333 (N_11333,N_10837,N_11074);
nand U11334 (N_11334,N_10750,N_10980);
xnor U11335 (N_11335,N_10552,N_10881);
or U11336 (N_11336,N_10786,N_10756);
and U11337 (N_11337,N_10952,N_11131);
nand U11338 (N_11338,N_11177,N_10759);
or U11339 (N_11339,N_11165,N_11205);
xnor U11340 (N_11340,N_10943,N_10743);
nand U11341 (N_11341,N_11006,N_11130);
xnor U11342 (N_11342,N_10973,N_10895);
or U11343 (N_11343,N_10517,N_10932);
nor U11344 (N_11344,N_10622,N_10697);
or U11345 (N_11345,N_10793,N_10513);
xnor U11346 (N_11346,N_10948,N_10784);
nor U11347 (N_11347,N_11120,N_10525);
and U11348 (N_11348,N_10692,N_10831);
and U11349 (N_11349,N_11145,N_11025);
xnor U11350 (N_11350,N_10543,N_10615);
nand U11351 (N_11351,N_11139,N_10982);
or U11352 (N_11352,N_10753,N_10581);
nand U11353 (N_11353,N_10911,N_11032);
xor U11354 (N_11354,N_11232,N_10894);
nand U11355 (N_11355,N_10796,N_10703);
or U11356 (N_11356,N_11227,N_11039);
nand U11357 (N_11357,N_10720,N_11195);
nor U11358 (N_11358,N_11105,N_11078);
nand U11359 (N_11359,N_10907,N_10658);
nor U11360 (N_11360,N_11153,N_11099);
nor U11361 (N_11361,N_10684,N_10924);
and U11362 (N_11362,N_11229,N_10967);
nor U11363 (N_11363,N_11035,N_11096);
or U11364 (N_11364,N_10981,N_11183);
or U11365 (N_11365,N_10740,N_10515);
nor U11366 (N_11366,N_11036,N_10781);
and U11367 (N_11367,N_10700,N_10890);
or U11368 (N_11368,N_10505,N_11248);
xor U11369 (N_11369,N_10702,N_10520);
xnor U11370 (N_11370,N_11149,N_10527);
nor U11371 (N_11371,N_10523,N_10541);
xor U11372 (N_11372,N_11173,N_10705);
xor U11373 (N_11373,N_10583,N_10600);
and U11374 (N_11374,N_10869,N_10906);
nor U11375 (N_11375,N_10970,N_11181);
xor U11376 (N_11376,N_10902,N_10501);
nor U11377 (N_11377,N_10861,N_11226);
nand U11378 (N_11378,N_11223,N_10865);
nor U11379 (N_11379,N_10754,N_11191);
xnor U11380 (N_11380,N_10644,N_10516);
xor U11381 (N_11381,N_10572,N_10997);
nand U11382 (N_11382,N_11076,N_11013);
or U11383 (N_11383,N_10548,N_10530);
and U11384 (N_11384,N_10579,N_10713);
or U11385 (N_11385,N_11077,N_11174);
and U11386 (N_11386,N_10736,N_10767);
or U11387 (N_11387,N_10820,N_10689);
and U11388 (N_11388,N_10867,N_11134);
or U11389 (N_11389,N_11020,N_11242);
or U11390 (N_11390,N_10599,N_11166);
nor U11391 (N_11391,N_10637,N_10695);
nor U11392 (N_11392,N_10630,N_10766);
xor U11393 (N_11393,N_10838,N_10848);
or U11394 (N_11394,N_10918,N_10778);
or U11395 (N_11395,N_11176,N_10956);
or U11396 (N_11396,N_10984,N_10844);
nor U11397 (N_11397,N_11220,N_10547);
nand U11398 (N_11398,N_10834,N_11201);
xnor U11399 (N_11399,N_10648,N_11090);
xnor U11400 (N_11400,N_10714,N_10955);
xor U11401 (N_11401,N_10624,N_10816);
and U11402 (N_11402,N_10655,N_10988);
or U11403 (N_11403,N_11206,N_11222);
nand U11404 (N_11404,N_11236,N_10765);
nand U11405 (N_11405,N_10986,N_11058);
nand U11406 (N_11406,N_10575,N_10534);
xnor U11407 (N_11407,N_10620,N_10958);
and U11408 (N_11408,N_11002,N_10549);
nor U11409 (N_11409,N_10917,N_10770);
nor U11410 (N_11410,N_10814,N_10663);
xnor U11411 (N_11411,N_10634,N_11048);
nor U11412 (N_11412,N_11009,N_10780);
and U11413 (N_11413,N_10916,N_10927);
or U11414 (N_11414,N_10614,N_10905);
nand U11415 (N_11415,N_10835,N_10903);
nand U11416 (N_11416,N_11160,N_11158);
nor U11417 (N_11417,N_10993,N_11184);
or U11418 (N_11418,N_11024,N_11060);
nor U11419 (N_11419,N_10828,N_11249);
nand U11420 (N_11420,N_11190,N_11104);
and U11421 (N_11421,N_10687,N_10930);
and U11422 (N_11422,N_11045,N_11210);
or U11423 (N_11423,N_11192,N_11218);
xnor U11424 (N_11424,N_10764,N_10519);
xnor U11425 (N_11425,N_11217,N_11196);
or U11426 (N_11426,N_11207,N_10945);
xnor U11427 (N_11427,N_10654,N_11148);
and U11428 (N_11428,N_10858,N_11019);
xnor U11429 (N_11429,N_11152,N_11155);
or U11430 (N_11430,N_10578,N_10567);
nor U11431 (N_11431,N_10755,N_10694);
xor U11432 (N_11432,N_10532,N_10731);
nand U11433 (N_11433,N_11188,N_10896);
xor U11434 (N_11434,N_10718,N_10925);
and U11435 (N_11435,N_11189,N_11012);
or U11436 (N_11436,N_11000,N_10760);
nor U11437 (N_11437,N_11247,N_10609);
xor U11438 (N_11438,N_10656,N_11098);
nor U11439 (N_11439,N_11085,N_10799);
nor U11440 (N_11440,N_10651,N_11029);
or U11441 (N_11441,N_10514,N_11164);
or U11442 (N_11442,N_11027,N_10589);
nand U11443 (N_11443,N_11135,N_10817);
or U11444 (N_11444,N_10554,N_11143);
nand U11445 (N_11445,N_10832,N_10723);
nand U11446 (N_11446,N_10597,N_10863);
nand U11447 (N_11447,N_11138,N_10818);
and U11448 (N_11448,N_11061,N_10957);
nand U11449 (N_11449,N_11030,N_10876);
or U11450 (N_11450,N_10611,N_10686);
xnor U11451 (N_11451,N_11112,N_10711);
nand U11452 (N_11452,N_10893,N_10829);
nand U11453 (N_11453,N_11144,N_11199);
nand U11454 (N_11454,N_10733,N_10745);
and U11455 (N_11455,N_10994,N_10540);
xor U11456 (N_11456,N_11016,N_10882);
xnor U11457 (N_11457,N_11162,N_10741);
nor U11458 (N_11458,N_11005,N_10974);
or U11459 (N_11459,N_10564,N_11197);
nand U11460 (N_11460,N_10819,N_11119);
and U11461 (N_11461,N_10878,N_11066);
xor U11462 (N_11462,N_10735,N_11054);
or U11463 (N_11463,N_11042,N_10645);
xnor U11464 (N_11464,N_10747,N_10929);
xnor U11465 (N_11465,N_11204,N_11055);
and U11466 (N_11466,N_10716,N_10727);
nor U11467 (N_11467,N_11161,N_10643);
or U11468 (N_11468,N_10603,N_10830);
nor U11469 (N_11469,N_11169,N_10800);
and U11470 (N_11470,N_10752,N_11225);
and U11471 (N_11471,N_11194,N_10999);
and U11472 (N_11472,N_10533,N_10709);
and U11473 (N_11473,N_10571,N_10618);
nor U11474 (N_11474,N_10725,N_10995);
and U11475 (N_11475,N_10909,N_11246);
xor U11476 (N_11476,N_10636,N_10626);
and U11477 (N_11477,N_10921,N_10803);
nor U11478 (N_11478,N_11014,N_11245);
xor U11479 (N_11479,N_11011,N_10691);
xor U11480 (N_11480,N_10859,N_10612);
or U11481 (N_11481,N_10596,N_11133);
xor U11482 (N_11482,N_10698,N_10839);
or U11483 (N_11483,N_11057,N_10772);
and U11484 (N_11484,N_11021,N_10985);
and U11485 (N_11485,N_10935,N_10748);
and U11486 (N_11486,N_10674,N_11228);
nand U11487 (N_11487,N_10855,N_11086);
nand U11488 (N_11488,N_10586,N_10664);
or U11489 (N_11489,N_11067,N_10919);
or U11490 (N_11490,N_11109,N_10559);
nand U11491 (N_11491,N_11175,N_10783);
nand U11492 (N_11492,N_11215,N_11114);
xor U11493 (N_11493,N_10595,N_10591);
nand U11494 (N_11494,N_10531,N_10528);
xor U11495 (N_11495,N_10889,N_10946);
and U11496 (N_11496,N_10677,N_10627);
nand U11497 (N_11497,N_11083,N_10811);
xnor U11498 (N_11498,N_11115,N_11072);
and U11499 (N_11499,N_10635,N_10989);
or U11500 (N_11500,N_10565,N_10971);
or U11501 (N_11501,N_10668,N_11212);
or U11502 (N_11502,N_10749,N_11214);
xor U11503 (N_11503,N_10667,N_10726);
nand U11504 (N_11504,N_11047,N_10771);
xor U11505 (N_11505,N_11213,N_11151);
nand U11506 (N_11506,N_10774,N_10789);
and U11507 (N_11507,N_10509,N_10673);
nor U11508 (N_11508,N_10500,N_11202);
and U11509 (N_11509,N_10699,N_11219);
xnor U11510 (N_11510,N_10763,N_11007);
xor U11511 (N_11511,N_10577,N_10537);
and U11512 (N_11512,N_10864,N_10875);
nor U11513 (N_11513,N_10758,N_11243);
nor U11514 (N_11514,N_10729,N_11075);
or U11515 (N_11515,N_11106,N_10963);
xnor U11516 (N_11516,N_11080,N_10908);
xor U11517 (N_11517,N_10913,N_10804);
nand U11518 (N_11518,N_10573,N_10991);
nand U11519 (N_11519,N_11092,N_11123);
or U11520 (N_11520,N_10976,N_10825);
xnor U11521 (N_11521,N_11150,N_11203);
nand U11522 (N_11522,N_10632,N_10891);
or U11523 (N_11523,N_10915,N_11159);
nor U11524 (N_11524,N_11231,N_10638);
nor U11525 (N_11525,N_10826,N_11052);
or U11526 (N_11526,N_10898,N_11073);
and U11527 (N_11527,N_10506,N_10551);
nor U11528 (N_11528,N_10507,N_10969);
nand U11529 (N_11529,N_10685,N_10738);
or U11530 (N_11530,N_10659,N_10558);
nand U11531 (N_11531,N_10646,N_11103);
nor U11532 (N_11532,N_10872,N_10608);
nor U11533 (N_11533,N_10671,N_10623);
or U11534 (N_11534,N_10503,N_10840);
nand U11535 (N_11535,N_10975,N_10569);
or U11536 (N_11536,N_10775,N_11146);
nor U11537 (N_11537,N_10676,N_10757);
nand U11538 (N_11538,N_10683,N_11003);
and U11539 (N_11539,N_10542,N_10546);
or U11540 (N_11540,N_10941,N_10751);
nand U11541 (N_11541,N_10724,N_10802);
or U11542 (N_11542,N_10873,N_10904);
nand U11543 (N_11543,N_10926,N_11168);
or U11544 (N_11544,N_10710,N_11049);
xnor U11545 (N_11545,N_10883,N_10587);
nor U11546 (N_11546,N_11034,N_10899);
and U11547 (N_11547,N_10923,N_10806);
nand U11548 (N_11548,N_10721,N_10708);
and U11549 (N_11549,N_10949,N_10512);
nor U11550 (N_11550,N_11053,N_10707);
xnor U11551 (N_11551,N_10847,N_11237);
or U11552 (N_11552,N_10824,N_10849);
or U11553 (N_11553,N_11100,N_10934);
and U11554 (N_11554,N_10884,N_10959);
nor U11555 (N_11555,N_10901,N_10605);
nor U11556 (N_11556,N_11239,N_10619);
and U11557 (N_11557,N_11178,N_11017);
and U11558 (N_11558,N_10722,N_10607);
xor U11559 (N_11559,N_10566,N_10641);
nand U11560 (N_11560,N_10593,N_10968);
nand U11561 (N_11561,N_10616,N_11026);
and U11562 (N_11562,N_11221,N_11118);
xor U11563 (N_11563,N_11241,N_10972);
and U11564 (N_11564,N_10511,N_11121);
nor U11565 (N_11565,N_10553,N_10782);
nand U11566 (N_11566,N_10797,N_10877);
nor U11567 (N_11567,N_10679,N_10670);
and U11568 (N_11568,N_10628,N_10846);
and U11569 (N_11569,N_11193,N_10897);
and U11570 (N_11570,N_10522,N_11028);
xnor U11571 (N_11571,N_10888,N_11211);
nor U11572 (N_11572,N_11038,N_10940);
nand U11573 (N_11573,N_10561,N_10510);
nor U11574 (N_11574,N_11117,N_10880);
nor U11575 (N_11575,N_10960,N_10942);
xnor U11576 (N_11576,N_11088,N_10841);
and U11577 (N_11577,N_10728,N_11059);
or U11578 (N_11578,N_10690,N_11091);
xor U11579 (N_11579,N_10805,N_10792);
nor U11580 (N_11580,N_11198,N_11156);
nand U11581 (N_11581,N_10810,N_11082);
xor U11582 (N_11582,N_11089,N_11172);
and U11583 (N_11583,N_10944,N_10860);
nor U11584 (N_11584,N_11179,N_10621);
or U11585 (N_11585,N_11240,N_11033);
nand U11586 (N_11586,N_10931,N_10761);
and U11587 (N_11587,N_11050,N_10801);
nor U11588 (N_11588,N_11142,N_11044);
or U11589 (N_11589,N_10557,N_10504);
nor U11590 (N_11590,N_10734,N_10954);
or U11591 (N_11591,N_10887,N_10535);
xnor U11592 (N_11592,N_10809,N_10633);
nand U11593 (N_11593,N_11171,N_10788);
and U11594 (N_11594,N_10812,N_11128);
nand U11595 (N_11595,N_10660,N_10779);
xnor U11596 (N_11596,N_10706,N_10592);
nor U11597 (N_11597,N_10661,N_11230);
and U11598 (N_11598,N_10951,N_11209);
nor U11599 (N_11599,N_11113,N_10870);
xnor U11600 (N_11600,N_11094,N_10712);
nor U11601 (N_11601,N_10886,N_10544);
xor U11602 (N_11602,N_10539,N_10594);
or U11603 (N_11603,N_10871,N_11108);
or U11604 (N_11604,N_10892,N_10790);
and U11605 (N_11605,N_11063,N_10910);
and U11606 (N_11606,N_10639,N_10574);
nand U11607 (N_11607,N_10652,N_10947);
or U11608 (N_11608,N_10732,N_10966);
nor U11609 (N_11609,N_10580,N_10856);
and U11610 (N_11610,N_10843,N_11216);
xnor U11611 (N_11611,N_11062,N_10762);
and U11612 (N_11612,N_11101,N_11041);
or U11613 (N_11613,N_11140,N_10833);
nand U11614 (N_11614,N_11234,N_10983);
and U11615 (N_11615,N_11070,N_10866);
or U11616 (N_11616,N_10568,N_11110);
nor U11617 (N_11617,N_10850,N_10977);
xor U11618 (N_11618,N_11244,N_11018);
nor U11619 (N_11619,N_10842,N_10992);
nand U11620 (N_11620,N_10798,N_11163);
and U11621 (N_11621,N_10928,N_10961);
and U11622 (N_11622,N_10678,N_10653);
xnor U11623 (N_11623,N_10777,N_11046);
nor U11624 (N_11624,N_11069,N_10682);
or U11625 (N_11625,N_11242,N_10946);
and U11626 (N_11626,N_10635,N_10932);
and U11627 (N_11627,N_10809,N_10916);
or U11628 (N_11628,N_10956,N_10943);
xnor U11629 (N_11629,N_10519,N_11035);
nor U11630 (N_11630,N_11134,N_10857);
or U11631 (N_11631,N_10833,N_10655);
or U11632 (N_11632,N_11090,N_10875);
xor U11633 (N_11633,N_10740,N_10877);
or U11634 (N_11634,N_11062,N_10996);
nand U11635 (N_11635,N_11203,N_10804);
or U11636 (N_11636,N_11091,N_10535);
nand U11637 (N_11637,N_10731,N_11113);
xor U11638 (N_11638,N_10963,N_11044);
and U11639 (N_11639,N_10587,N_10924);
nor U11640 (N_11640,N_10880,N_10934);
and U11641 (N_11641,N_10512,N_10594);
nand U11642 (N_11642,N_10929,N_11092);
and U11643 (N_11643,N_11077,N_11005);
and U11644 (N_11644,N_10760,N_10507);
and U11645 (N_11645,N_11192,N_10660);
nor U11646 (N_11646,N_11150,N_10782);
or U11647 (N_11647,N_10980,N_10983);
nand U11648 (N_11648,N_10906,N_11215);
xor U11649 (N_11649,N_11207,N_10757);
nor U11650 (N_11650,N_10650,N_11225);
nand U11651 (N_11651,N_10794,N_10872);
and U11652 (N_11652,N_11222,N_10962);
and U11653 (N_11653,N_11016,N_10899);
nor U11654 (N_11654,N_10790,N_10800);
xnor U11655 (N_11655,N_10811,N_11016);
and U11656 (N_11656,N_10541,N_11121);
xor U11657 (N_11657,N_10907,N_10826);
nor U11658 (N_11658,N_10974,N_10655);
and U11659 (N_11659,N_10754,N_10820);
nand U11660 (N_11660,N_11086,N_10904);
and U11661 (N_11661,N_10739,N_10562);
or U11662 (N_11662,N_10841,N_10506);
nor U11663 (N_11663,N_11073,N_11173);
xor U11664 (N_11664,N_11116,N_10718);
and U11665 (N_11665,N_10833,N_10979);
nor U11666 (N_11666,N_11038,N_10977);
nand U11667 (N_11667,N_10758,N_11161);
xnor U11668 (N_11668,N_10703,N_10766);
nor U11669 (N_11669,N_11164,N_10712);
or U11670 (N_11670,N_11083,N_10928);
xnor U11671 (N_11671,N_10836,N_10979);
nand U11672 (N_11672,N_10531,N_11100);
xor U11673 (N_11673,N_10834,N_10639);
and U11674 (N_11674,N_10773,N_10689);
nor U11675 (N_11675,N_11137,N_10644);
and U11676 (N_11676,N_10753,N_10931);
nand U11677 (N_11677,N_10508,N_10807);
xnor U11678 (N_11678,N_10865,N_11022);
nand U11679 (N_11679,N_11227,N_10721);
xnor U11680 (N_11680,N_10933,N_10981);
xnor U11681 (N_11681,N_10619,N_11148);
or U11682 (N_11682,N_10864,N_11104);
and U11683 (N_11683,N_11011,N_10759);
nand U11684 (N_11684,N_10606,N_10837);
or U11685 (N_11685,N_11194,N_11193);
xnor U11686 (N_11686,N_10782,N_10752);
nor U11687 (N_11687,N_10868,N_10527);
xor U11688 (N_11688,N_10577,N_11172);
nand U11689 (N_11689,N_11094,N_10689);
nor U11690 (N_11690,N_11152,N_11061);
or U11691 (N_11691,N_10689,N_10792);
nor U11692 (N_11692,N_11054,N_10983);
xor U11693 (N_11693,N_10547,N_11204);
nand U11694 (N_11694,N_10799,N_11067);
nor U11695 (N_11695,N_11080,N_10513);
xnor U11696 (N_11696,N_10759,N_11090);
or U11697 (N_11697,N_10612,N_10990);
xnor U11698 (N_11698,N_10618,N_11212);
or U11699 (N_11699,N_10974,N_11148);
nor U11700 (N_11700,N_10978,N_10605);
nor U11701 (N_11701,N_11005,N_10538);
and U11702 (N_11702,N_11173,N_10828);
xnor U11703 (N_11703,N_10769,N_11093);
and U11704 (N_11704,N_10714,N_10622);
and U11705 (N_11705,N_10725,N_10501);
and U11706 (N_11706,N_10803,N_11232);
nor U11707 (N_11707,N_10906,N_10865);
nor U11708 (N_11708,N_11189,N_10712);
and U11709 (N_11709,N_10937,N_11044);
nand U11710 (N_11710,N_10555,N_10516);
nand U11711 (N_11711,N_10973,N_10576);
nor U11712 (N_11712,N_10508,N_11065);
xor U11713 (N_11713,N_11118,N_10862);
nand U11714 (N_11714,N_10596,N_11043);
nand U11715 (N_11715,N_10903,N_11081);
or U11716 (N_11716,N_11129,N_11109);
and U11717 (N_11717,N_11030,N_11115);
or U11718 (N_11718,N_10594,N_10624);
xor U11719 (N_11719,N_10709,N_10512);
xnor U11720 (N_11720,N_11204,N_10678);
and U11721 (N_11721,N_10713,N_11209);
nand U11722 (N_11722,N_11139,N_10903);
nor U11723 (N_11723,N_11201,N_10848);
nand U11724 (N_11724,N_11077,N_10866);
nand U11725 (N_11725,N_10613,N_10585);
xor U11726 (N_11726,N_11075,N_10851);
and U11727 (N_11727,N_10588,N_10604);
xor U11728 (N_11728,N_10799,N_10696);
or U11729 (N_11729,N_10631,N_10587);
and U11730 (N_11730,N_10719,N_10894);
or U11731 (N_11731,N_11210,N_11032);
nand U11732 (N_11732,N_10696,N_10542);
or U11733 (N_11733,N_11040,N_10825);
xnor U11734 (N_11734,N_11077,N_11119);
nand U11735 (N_11735,N_10526,N_10577);
and U11736 (N_11736,N_10916,N_10939);
xor U11737 (N_11737,N_11242,N_11176);
xnor U11738 (N_11738,N_10792,N_10514);
xnor U11739 (N_11739,N_10604,N_11055);
xor U11740 (N_11740,N_10955,N_10731);
or U11741 (N_11741,N_11010,N_11015);
nor U11742 (N_11742,N_10575,N_11057);
nor U11743 (N_11743,N_10691,N_10674);
xor U11744 (N_11744,N_10839,N_10919);
xor U11745 (N_11745,N_11127,N_10579);
nor U11746 (N_11746,N_10894,N_10508);
nand U11747 (N_11747,N_11212,N_11033);
nand U11748 (N_11748,N_10784,N_11067);
and U11749 (N_11749,N_11211,N_10563);
nor U11750 (N_11750,N_10535,N_10949);
xor U11751 (N_11751,N_10529,N_10927);
nor U11752 (N_11752,N_11201,N_11024);
xor U11753 (N_11753,N_10500,N_10780);
nor U11754 (N_11754,N_10765,N_10683);
nand U11755 (N_11755,N_10528,N_10799);
or U11756 (N_11756,N_11215,N_10615);
xor U11757 (N_11757,N_11054,N_10703);
nor U11758 (N_11758,N_11239,N_10968);
and U11759 (N_11759,N_11020,N_11171);
nand U11760 (N_11760,N_11249,N_10886);
nor U11761 (N_11761,N_10786,N_10535);
or U11762 (N_11762,N_10661,N_11191);
xnor U11763 (N_11763,N_10764,N_10646);
xor U11764 (N_11764,N_11186,N_10808);
nor U11765 (N_11765,N_10917,N_10721);
xnor U11766 (N_11766,N_11198,N_10709);
xor U11767 (N_11767,N_11183,N_10819);
nand U11768 (N_11768,N_10883,N_10510);
and U11769 (N_11769,N_10862,N_10634);
nand U11770 (N_11770,N_11159,N_10862);
xor U11771 (N_11771,N_11213,N_10727);
and U11772 (N_11772,N_11186,N_10820);
and U11773 (N_11773,N_10967,N_10786);
nand U11774 (N_11774,N_10862,N_10507);
and U11775 (N_11775,N_11073,N_10948);
nand U11776 (N_11776,N_10702,N_11197);
xnor U11777 (N_11777,N_11049,N_10611);
or U11778 (N_11778,N_10546,N_10578);
xor U11779 (N_11779,N_11135,N_11087);
nand U11780 (N_11780,N_10670,N_10824);
or U11781 (N_11781,N_11217,N_10946);
and U11782 (N_11782,N_10878,N_10693);
nand U11783 (N_11783,N_10701,N_11053);
xnor U11784 (N_11784,N_10975,N_11184);
xor U11785 (N_11785,N_10851,N_11246);
or U11786 (N_11786,N_11012,N_10653);
or U11787 (N_11787,N_10951,N_10869);
and U11788 (N_11788,N_11043,N_10608);
and U11789 (N_11789,N_10676,N_11223);
or U11790 (N_11790,N_10585,N_10659);
xor U11791 (N_11791,N_10929,N_10996);
nand U11792 (N_11792,N_10992,N_11228);
nor U11793 (N_11793,N_10671,N_10651);
nor U11794 (N_11794,N_11101,N_10717);
or U11795 (N_11795,N_10986,N_10778);
xor U11796 (N_11796,N_11051,N_10802);
nor U11797 (N_11797,N_10511,N_11140);
nand U11798 (N_11798,N_10786,N_11040);
and U11799 (N_11799,N_10575,N_10742);
nand U11800 (N_11800,N_11020,N_10542);
or U11801 (N_11801,N_10834,N_10913);
nand U11802 (N_11802,N_11123,N_11019);
and U11803 (N_11803,N_10812,N_10570);
or U11804 (N_11804,N_10939,N_10505);
xor U11805 (N_11805,N_10784,N_10597);
or U11806 (N_11806,N_11015,N_10737);
or U11807 (N_11807,N_11085,N_10958);
nand U11808 (N_11808,N_11120,N_10535);
nand U11809 (N_11809,N_11193,N_10978);
and U11810 (N_11810,N_10758,N_10977);
xnor U11811 (N_11811,N_10584,N_11053);
xnor U11812 (N_11812,N_10511,N_11031);
or U11813 (N_11813,N_10906,N_10955);
and U11814 (N_11814,N_10587,N_10845);
xnor U11815 (N_11815,N_10624,N_10681);
nand U11816 (N_11816,N_10719,N_11048);
nand U11817 (N_11817,N_11082,N_10550);
nand U11818 (N_11818,N_11195,N_10885);
and U11819 (N_11819,N_10899,N_11109);
xnor U11820 (N_11820,N_10631,N_10983);
nand U11821 (N_11821,N_10984,N_11021);
xnor U11822 (N_11822,N_10621,N_10965);
nor U11823 (N_11823,N_10746,N_10949);
nand U11824 (N_11824,N_11135,N_10563);
or U11825 (N_11825,N_11019,N_11188);
and U11826 (N_11826,N_10608,N_10830);
or U11827 (N_11827,N_11031,N_10548);
and U11828 (N_11828,N_10941,N_10891);
and U11829 (N_11829,N_11195,N_11170);
and U11830 (N_11830,N_11181,N_10956);
xnor U11831 (N_11831,N_10591,N_10677);
or U11832 (N_11832,N_11054,N_10839);
or U11833 (N_11833,N_10884,N_11166);
xor U11834 (N_11834,N_10521,N_11167);
or U11835 (N_11835,N_10998,N_11169);
xor U11836 (N_11836,N_11236,N_11185);
and U11837 (N_11837,N_10563,N_10624);
nor U11838 (N_11838,N_10979,N_10678);
nor U11839 (N_11839,N_10850,N_10830);
xnor U11840 (N_11840,N_10539,N_10783);
or U11841 (N_11841,N_10533,N_10975);
nor U11842 (N_11842,N_10986,N_10873);
or U11843 (N_11843,N_10544,N_10865);
and U11844 (N_11844,N_10946,N_10508);
xnor U11845 (N_11845,N_11048,N_10973);
or U11846 (N_11846,N_10643,N_10687);
xnor U11847 (N_11847,N_10641,N_10960);
xnor U11848 (N_11848,N_10564,N_11214);
nand U11849 (N_11849,N_10854,N_11065);
nand U11850 (N_11850,N_11057,N_10789);
xor U11851 (N_11851,N_11084,N_10839);
xnor U11852 (N_11852,N_10893,N_11063);
nor U11853 (N_11853,N_10783,N_11083);
nand U11854 (N_11854,N_10764,N_11159);
and U11855 (N_11855,N_11170,N_10603);
or U11856 (N_11856,N_10876,N_10725);
nor U11857 (N_11857,N_10939,N_10950);
nor U11858 (N_11858,N_10856,N_10735);
nand U11859 (N_11859,N_10988,N_10888);
or U11860 (N_11860,N_10868,N_10889);
and U11861 (N_11861,N_10923,N_10896);
xnor U11862 (N_11862,N_11229,N_10619);
and U11863 (N_11863,N_10852,N_11228);
nor U11864 (N_11864,N_11201,N_10688);
and U11865 (N_11865,N_11035,N_10861);
or U11866 (N_11866,N_11160,N_11242);
nand U11867 (N_11867,N_10583,N_10912);
nand U11868 (N_11868,N_10813,N_11233);
nor U11869 (N_11869,N_10981,N_10602);
nor U11870 (N_11870,N_11118,N_11138);
xnor U11871 (N_11871,N_11194,N_11032);
xnor U11872 (N_11872,N_10569,N_10502);
or U11873 (N_11873,N_10583,N_10798);
nand U11874 (N_11874,N_11152,N_11125);
or U11875 (N_11875,N_10934,N_10799);
nor U11876 (N_11876,N_10748,N_10937);
or U11877 (N_11877,N_10569,N_11192);
or U11878 (N_11878,N_10594,N_11027);
or U11879 (N_11879,N_10662,N_10671);
and U11880 (N_11880,N_10736,N_10713);
nor U11881 (N_11881,N_10642,N_10964);
xor U11882 (N_11882,N_10992,N_10824);
nand U11883 (N_11883,N_10505,N_10705);
nor U11884 (N_11884,N_10909,N_10578);
xnor U11885 (N_11885,N_10995,N_10570);
and U11886 (N_11886,N_10540,N_10662);
nand U11887 (N_11887,N_10641,N_10747);
or U11888 (N_11888,N_10904,N_11081);
or U11889 (N_11889,N_10703,N_10516);
nor U11890 (N_11890,N_11237,N_10740);
nor U11891 (N_11891,N_10783,N_10695);
nand U11892 (N_11892,N_10814,N_11010);
or U11893 (N_11893,N_11145,N_10777);
and U11894 (N_11894,N_10886,N_10924);
nand U11895 (N_11895,N_10625,N_10815);
nand U11896 (N_11896,N_10605,N_11112);
xnor U11897 (N_11897,N_11144,N_10591);
and U11898 (N_11898,N_10534,N_11083);
nand U11899 (N_11899,N_11085,N_10886);
xnor U11900 (N_11900,N_11139,N_11200);
xnor U11901 (N_11901,N_10940,N_10526);
nand U11902 (N_11902,N_10544,N_11185);
and U11903 (N_11903,N_11063,N_10716);
nand U11904 (N_11904,N_11113,N_10858);
or U11905 (N_11905,N_10681,N_10603);
and U11906 (N_11906,N_10990,N_10541);
or U11907 (N_11907,N_10610,N_10629);
xor U11908 (N_11908,N_10531,N_10899);
nand U11909 (N_11909,N_10512,N_10954);
xor U11910 (N_11910,N_10527,N_10514);
or U11911 (N_11911,N_10845,N_10739);
nand U11912 (N_11912,N_11149,N_10934);
and U11913 (N_11913,N_11171,N_11139);
nand U11914 (N_11914,N_10664,N_10545);
nor U11915 (N_11915,N_11234,N_10550);
and U11916 (N_11916,N_10953,N_11223);
nor U11917 (N_11917,N_11065,N_11111);
or U11918 (N_11918,N_10975,N_10759);
and U11919 (N_11919,N_11009,N_10725);
nand U11920 (N_11920,N_10982,N_11081);
nand U11921 (N_11921,N_10796,N_10941);
nand U11922 (N_11922,N_10788,N_10560);
nor U11923 (N_11923,N_11109,N_10887);
nor U11924 (N_11924,N_10974,N_10619);
or U11925 (N_11925,N_10668,N_11086);
nand U11926 (N_11926,N_10878,N_10629);
xor U11927 (N_11927,N_11132,N_11106);
nor U11928 (N_11928,N_10825,N_11170);
nand U11929 (N_11929,N_10753,N_10958);
and U11930 (N_11930,N_11004,N_11228);
or U11931 (N_11931,N_10506,N_10938);
xnor U11932 (N_11932,N_10527,N_10611);
and U11933 (N_11933,N_10829,N_11027);
xnor U11934 (N_11934,N_11178,N_10980);
xor U11935 (N_11935,N_11025,N_10723);
nand U11936 (N_11936,N_10961,N_10981);
nand U11937 (N_11937,N_11020,N_10605);
and U11938 (N_11938,N_10555,N_11158);
nand U11939 (N_11939,N_11101,N_10852);
or U11940 (N_11940,N_10937,N_10835);
and U11941 (N_11941,N_11168,N_10944);
xor U11942 (N_11942,N_10603,N_10919);
xnor U11943 (N_11943,N_11085,N_10859);
and U11944 (N_11944,N_10787,N_10544);
and U11945 (N_11945,N_10957,N_10754);
or U11946 (N_11946,N_11080,N_10655);
nor U11947 (N_11947,N_10813,N_10635);
and U11948 (N_11948,N_11206,N_11066);
xor U11949 (N_11949,N_10742,N_11248);
and U11950 (N_11950,N_11108,N_11159);
xnor U11951 (N_11951,N_10788,N_10961);
and U11952 (N_11952,N_11072,N_10525);
nand U11953 (N_11953,N_10802,N_11092);
and U11954 (N_11954,N_10631,N_10721);
nor U11955 (N_11955,N_10645,N_11001);
nor U11956 (N_11956,N_10584,N_11148);
and U11957 (N_11957,N_10844,N_11245);
or U11958 (N_11958,N_10915,N_10977);
nor U11959 (N_11959,N_11244,N_11045);
nand U11960 (N_11960,N_10811,N_11128);
or U11961 (N_11961,N_10929,N_10595);
nand U11962 (N_11962,N_11177,N_10522);
nand U11963 (N_11963,N_10675,N_10701);
and U11964 (N_11964,N_11229,N_10522);
or U11965 (N_11965,N_11176,N_11038);
nand U11966 (N_11966,N_10777,N_11234);
or U11967 (N_11967,N_10940,N_10942);
nor U11968 (N_11968,N_10607,N_10557);
and U11969 (N_11969,N_10797,N_11107);
and U11970 (N_11970,N_10567,N_11140);
nand U11971 (N_11971,N_10656,N_10862);
xor U11972 (N_11972,N_11173,N_11198);
and U11973 (N_11973,N_11147,N_10596);
nor U11974 (N_11974,N_10795,N_10631);
nor U11975 (N_11975,N_10656,N_11100);
xnor U11976 (N_11976,N_11210,N_10566);
and U11977 (N_11977,N_10936,N_10887);
nand U11978 (N_11978,N_11139,N_10590);
and U11979 (N_11979,N_10807,N_10882);
and U11980 (N_11980,N_10594,N_10686);
or U11981 (N_11981,N_11182,N_11096);
or U11982 (N_11982,N_10969,N_10505);
nand U11983 (N_11983,N_10535,N_10987);
nor U11984 (N_11984,N_11199,N_10847);
nor U11985 (N_11985,N_10683,N_10843);
nor U11986 (N_11986,N_11007,N_11234);
nand U11987 (N_11987,N_11132,N_11140);
nand U11988 (N_11988,N_10899,N_10609);
or U11989 (N_11989,N_10726,N_10666);
nand U11990 (N_11990,N_10882,N_11137);
nand U11991 (N_11991,N_11138,N_10530);
xnor U11992 (N_11992,N_10749,N_10652);
nand U11993 (N_11993,N_10780,N_11031);
xnor U11994 (N_11994,N_10712,N_11106);
and U11995 (N_11995,N_10939,N_10809);
or U11996 (N_11996,N_10797,N_11143);
nand U11997 (N_11997,N_11145,N_10631);
nor U11998 (N_11998,N_10784,N_10606);
xnor U11999 (N_11999,N_10677,N_10869);
or U12000 (N_12000,N_11646,N_11893);
or U12001 (N_12001,N_11948,N_11934);
nor U12002 (N_12002,N_11476,N_11597);
and U12003 (N_12003,N_11531,N_11935);
nor U12004 (N_12004,N_11255,N_11324);
nand U12005 (N_12005,N_11551,N_11391);
nand U12006 (N_12006,N_11485,N_11899);
nand U12007 (N_12007,N_11705,N_11608);
and U12008 (N_12008,N_11858,N_11456);
or U12009 (N_12009,N_11349,N_11575);
xor U12010 (N_12010,N_11572,N_11801);
xor U12011 (N_12011,N_11779,N_11778);
or U12012 (N_12012,N_11536,N_11716);
and U12013 (N_12013,N_11861,N_11663);
or U12014 (N_12014,N_11432,N_11777);
nand U12015 (N_12015,N_11402,N_11812);
xor U12016 (N_12016,N_11684,N_11322);
and U12017 (N_12017,N_11878,N_11541);
nor U12018 (N_12018,N_11366,N_11973);
or U12019 (N_12019,N_11958,N_11920);
nor U12020 (N_12020,N_11339,N_11767);
xor U12021 (N_12021,N_11637,N_11983);
nor U12022 (N_12022,N_11997,N_11954);
or U12023 (N_12023,N_11522,N_11872);
or U12024 (N_12024,N_11383,N_11832);
or U12025 (N_12025,N_11772,N_11454);
and U12026 (N_12026,N_11963,N_11765);
nor U12027 (N_12027,N_11901,N_11844);
xnor U12028 (N_12028,N_11481,N_11826);
or U12029 (N_12029,N_11250,N_11873);
or U12030 (N_12030,N_11857,N_11927);
xor U12031 (N_12031,N_11361,N_11883);
nand U12032 (N_12032,N_11253,N_11664);
or U12033 (N_12033,N_11569,N_11396);
xnor U12034 (N_12034,N_11760,N_11841);
or U12035 (N_12035,N_11519,N_11823);
or U12036 (N_12036,N_11513,N_11981);
or U12037 (N_12037,N_11980,N_11377);
xnor U12038 (N_12038,N_11840,N_11769);
or U12039 (N_12039,N_11284,N_11923);
or U12040 (N_12040,N_11375,N_11782);
and U12041 (N_12041,N_11443,N_11412);
nand U12042 (N_12042,N_11437,N_11265);
and U12043 (N_12043,N_11296,N_11492);
nand U12044 (N_12044,N_11933,N_11763);
xor U12045 (N_12045,N_11517,N_11313);
or U12046 (N_12046,N_11896,N_11268);
xor U12047 (N_12047,N_11276,N_11468);
nor U12048 (N_12048,N_11364,N_11709);
nor U12049 (N_12049,N_11286,N_11588);
or U12050 (N_12050,N_11537,N_11732);
or U12051 (N_12051,N_11843,N_11549);
nand U12052 (N_12052,N_11404,N_11411);
nor U12053 (N_12053,N_11926,N_11881);
and U12054 (N_12054,N_11967,N_11849);
and U12055 (N_12055,N_11304,N_11379);
and U12056 (N_12056,N_11479,N_11816);
nand U12057 (N_12057,N_11644,N_11871);
and U12058 (N_12058,N_11472,N_11343);
nand U12059 (N_12059,N_11256,N_11312);
xor U12060 (N_12060,N_11853,N_11660);
nor U12061 (N_12061,N_11665,N_11384);
or U12062 (N_12062,N_11814,N_11419);
xor U12063 (N_12063,N_11356,N_11682);
nor U12064 (N_12064,N_11574,N_11949);
and U12065 (N_12065,N_11819,N_11876);
xnor U12066 (N_12066,N_11627,N_11774);
or U12067 (N_12067,N_11734,N_11631);
or U12068 (N_12068,N_11736,N_11251);
nor U12069 (N_12069,N_11333,N_11484);
nand U12070 (N_12070,N_11348,N_11420);
and U12071 (N_12071,N_11994,N_11982);
xor U12072 (N_12072,N_11510,N_11578);
nand U12073 (N_12073,N_11680,N_11565);
and U12074 (N_12074,N_11698,N_11652);
nor U12075 (N_12075,N_11672,N_11602);
and U12076 (N_12076,N_11700,N_11723);
and U12077 (N_12077,N_11547,N_11919);
and U12078 (N_12078,N_11441,N_11839);
and U12079 (N_12079,N_11619,N_11585);
xor U12080 (N_12080,N_11358,N_11270);
and U12081 (N_12081,N_11532,N_11793);
or U12082 (N_12082,N_11753,N_11498);
xor U12083 (N_12083,N_11946,N_11300);
nor U12084 (N_12084,N_11810,N_11376);
nand U12085 (N_12085,N_11499,N_11340);
xnor U12086 (N_12086,N_11696,N_11786);
or U12087 (N_12087,N_11798,N_11647);
and U12088 (N_12088,N_11850,N_11712);
xnor U12089 (N_12089,N_11368,N_11489);
or U12090 (N_12090,N_11668,N_11606);
and U12091 (N_12091,N_11689,N_11889);
xnor U12092 (N_12092,N_11905,N_11972);
nor U12093 (N_12093,N_11568,N_11721);
nor U12094 (N_12094,N_11950,N_11483);
and U12095 (N_12095,N_11325,N_11285);
or U12096 (N_12096,N_11415,N_11875);
xor U12097 (N_12097,N_11938,N_11761);
and U12098 (N_12098,N_11309,N_11351);
or U12099 (N_12099,N_11342,N_11471);
nand U12100 (N_12100,N_11720,N_11638);
nor U12101 (N_12101,N_11708,N_11687);
xor U12102 (N_12102,N_11310,N_11903);
nor U12103 (N_12103,N_11970,N_11922);
nor U12104 (N_12104,N_11542,N_11442);
or U12105 (N_12105,N_11388,N_11620);
nand U12106 (N_12106,N_11341,N_11681);
nor U12107 (N_12107,N_11653,N_11847);
xnor U12108 (N_12108,N_11392,N_11314);
xor U12109 (N_12109,N_11504,N_11534);
and U12110 (N_12110,N_11776,N_11624);
nor U12111 (N_12111,N_11451,N_11543);
and U12112 (N_12112,N_11280,N_11688);
nand U12113 (N_12113,N_11262,N_11929);
xnor U12114 (N_12114,N_11530,N_11453);
nand U12115 (N_12115,N_11957,N_11822);
and U12116 (N_12116,N_11544,N_11915);
and U12117 (N_12117,N_11830,N_11868);
and U12118 (N_12118,N_11320,N_11704);
nor U12119 (N_12119,N_11986,N_11390);
and U12120 (N_12120,N_11666,N_11387);
xor U12121 (N_12121,N_11748,N_11621);
xor U12122 (N_12122,N_11365,N_11703);
nand U12123 (N_12123,N_11610,N_11693);
or U12124 (N_12124,N_11879,N_11740);
nand U12125 (N_12125,N_11673,N_11766);
or U12126 (N_12126,N_11560,N_11591);
or U12127 (N_12127,N_11880,N_11589);
and U12128 (N_12128,N_11975,N_11452);
nand U12129 (N_12129,N_11338,N_11992);
and U12130 (N_12130,N_11439,N_11525);
or U12131 (N_12131,N_11527,N_11482);
nor U12132 (N_12132,N_11465,N_11506);
xnor U12133 (N_12133,N_11677,N_11892);
and U12134 (N_12134,N_11713,N_11811);
xnor U12135 (N_12135,N_11838,N_11557);
and U12136 (N_12136,N_11942,N_11900);
xor U12137 (N_12137,N_11350,N_11413);
or U12138 (N_12138,N_11287,N_11932);
xor U12139 (N_12139,N_11891,N_11882);
nand U12140 (N_12140,N_11429,N_11722);
nor U12141 (N_12141,N_11446,N_11979);
nor U12142 (N_12142,N_11533,N_11458);
or U12143 (N_12143,N_11553,N_11865);
or U12144 (N_12144,N_11433,N_11371);
nor U12145 (N_12145,N_11308,N_11555);
or U12146 (N_12146,N_11486,N_11791);
or U12147 (N_12147,N_11617,N_11321);
or U12148 (N_12148,N_11480,N_11971);
nand U12149 (N_12149,N_11599,N_11794);
or U12150 (N_12150,N_11742,N_11735);
or U12151 (N_12151,N_11961,N_11408);
xnor U12152 (N_12152,N_11616,N_11715);
xor U12153 (N_12153,N_11659,N_11870);
nand U12154 (N_12154,N_11434,N_11579);
nand U12155 (N_12155,N_11906,N_11497);
xnor U12156 (N_12156,N_11758,N_11477);
and U12157 (N_12157,N_11491,N_11969);
or U12158 (N_12158,N_11302,N_11630);
xnor U12159 (N_12159,N_11977,N_11488);
xnor U12160 (N_12160,N_11473,N_11425);
or U12161 (N_12161,N_11692,N_11757);
nand U12162 (N_12162,N_11360,N_11277);
nand U12163 (N_12163,N_11877,N_11526);
nor U12164 (N_12164,N_11584,N_11912);
and U12165 (N_12165,N_11357,N_11271);
and U12166 (N_12166,N_11267,N_11540);
nand U12167 (N_12167,N_11363,N_11707);
and U12168 (N_12168,N_11595,N_11347);
nand U12169 (N_12169,N_11475,N_11943);
nand U12170 (N_12170,N_11931,N_11636);
nor U12171 (N_12171,N_11406,N_11947);
xnor U12172 (N_12172,N_11305,N_11604);
nand U12173 (N_12173,N_11648,N_11625);
nor U12174 (N_12174,N_11487,N_11515);
nand U12175 (N_12175,N_11694,N_11651);
nor U12176 (N_12176,N_11645,N_11329);
and U12177 (N_12177,N_11805,N_11252);
or U12178 (N_12178,N_11331,N_11261);
or U12179 (N_12179,N_11508,N_11334);
nor U12180 (N_12180,N_11953,N_11385);
nand U12181 (N_12181,N_11924,N_11447);
and U12182 (N_12182,N_11895,N_11768);
nor U12183 (N_12183,N_11936,N_11728);
nor U12184 (N_12184,N_11785,N_11435);
xnor U12185 (N_12185,N_11800,N_11496);
nor U12186 (N_12186,N_11378,N_11829);
nand U12187 (N_12187,N_11685,N_11890);
nand U12188 (N_12188,N_11918,N_11848);
xor U12189 (N_12189,N_11764,N_11581);
or U12190 (N_12190,N_11611,N_11306);
or U12191 (N_12191,N_11614,N_11797);
or U12192 (N_12192,N_11490,N_11478);
nand U12193 (N_12193,N_11298,N_11632);
and U12194 (N_12194,N_11593,N_11559);
and U12195 (N_12195,N_11457,N_11423);
or U12196 (N_12196,N_11416,N_11438);
xnor U12197 (N_12197,N_11440,N_11539);
xor U12198 (N_12198,N_11724,N_11643);
nand U12199 (N_12199,N_11731,N_11374);
or U12200 (N_12200,N_11675,N_11886);
nand U12201 (N_12201,N_11548,N_11501);
or U12202 (N_12202,N_11678,N_11701);
or U12203 (N_12203,N_11956,N_11573);
nand U12204 (N_12204,N_11470,N_11729);
and U12205 (N_12205,N_11974,N_11834);
and U12206 (N_12206,N_11474,N_11299);
or U12207 (N_12207,N_11421,N_11609);
and U12208 (N_12208,N_11381,N_11626);
nand U12209 (N_12209,N_11528,N_11907);
xor U12210 (N_12210,N_11295,N_11293);
xor U12211 (N_12211,N_11607,N_11633);
and U12212 (N_12212,N_11372,N_11422);
xor U12213 (N_12213,N_11916,N_11711);
nand U12214 (N_12214,N_11804,N_11662);
or U12215 (N_12215,N_11649,N_11564);
nor U12216 (N_12216,N_11303,N_11409);
nor U12217 (N_12217,N_11874,N_11898);
and U12218 (N_12218,N_11796,N_11326);
nand U12219 (N_12219,N_11674,N_11462);
nand U12220 (N_12220,N_11683,N_11275);
nand U12221 (N_12221,N_11833,N_11799);
and U12222 (N_12222,N_11866,N_11828);
or U12223 (N_12223,N_11460,N_11571);
nand U12224 (N_12224,N_11596,N_11818);
nor U12225 (N_12225,N_11398,N_11512);
xnor U12226 (N_12226,N_11669,N_11657);
and U12227 (N_12227,N_11788,N_11820);
and U12228 (N_12228,N_11427,N_11913);
or U12229 (N_12229,N_11273,N_11998);
nor U12230 (N_12230,N_11639,N_11952);
or U12231 (N_12231,N_11968,N_11355);
and U12232 (N_12232,N_11759,N_11466);
nand U12233 (N_12233,N_11562,N_11815);
or U12234 (N_12234,N_11335,N_11332);
nand U12235 (N_12235,N_11990,N_11399);
or U12236 (N_12236,N_11289,N_11941);
or U12237 (N_12237,N_11353,N_11556);
xor U12238 (N_12238,N_11789,N_11613);
nand U12239 (N_12239,N_11410,N_11706);
or U12240 (N_12240,N_11783,N_11369);
and U12241 (N_12241,N_11751,N_11746);
nand U12242 (N_12242,N_11635,N_11655);
nor U12243 (N_12243,N_11566,N_11449);
or U12244 (N_12244,N_11962,N_11395);
nor U12245 (N_12245,N_11576,N_11825);
xor U12246 (N_12246,N_11911,N_11642);
nor U12247 (N_12247,N_11373,N_11301);
nand U12248 (N_12248,N_11787,N_11773);
and U12249 (N_12249,N_11586,N_11554);
or U12250 (N_12250,N_11336,N_11455);
or U12251 (N_12251,N_11494,N_11521);
or U12252 (N_12252,N_11529,N_11538);
nand U12253 (N_12253,N_11545,N_11756);
or U12254 (N_12254,N_11362,N_11945);
and U12255 (N_12255,N_11516,N_11955);
and U12256 (N_12256,N_11603,N_11897);
nand U12257 (N_12257,N_11254,N_11999);
xor U12258 (N_12258,N_11450,N_11869);
nor U12259 (N_12259,N_11623,N_11726);
nand U12260 (N_12260,N_11330,N_11702);
nand U12261 (N_12261,N_11634,N_11993);
xnor U12262 (N_12262,N_11459,N_11401);
and U12263 (N_12263,N_11743,N_11288);
xor U12264 (N_12264,N_11754,N_11930);
and U12265 (N_12265,N_11405,N_11505);
nor U12266 (N_12266,N_11940,N_11750);
or U12267 (N_12267,N_11699,N_11518);
and U12268 (N_12268,N_11282,N_11563);
and U12269 (N_12269,N_11592,N_11266);
xor U12270 (N_12270,N_11752,N_11960);
xor U12271 (N_12271,N_11928,N_11502);
nor U12272 (N_12272,N_11985,N_11714);
or U12273 (N_12273,N_11661,N_11802);
or U12274 (N_12274,N_11976,N_11775);
or U12275 (N_12275,N_11780,N_11686);
nor U12276 (N_12276,N_11283,N_11717);
or U12277 (N_12277,N_11264,N_11813);
and U12278 (N_12278,N_11784,N_11817);
nor U12279 (N_12279,N_11725,N_11317);
xor U12280 (N_12280,N_11978,N_11503);
or U12281 (N_12281,N_11656,N_11436);
and U12282 (N_12282,N_11337,N_11670);
nor U12283 (N_12283,N_11951,N_11426);
nand U12284 (N_12284,N_11444,N_11908);
or U12285 (N_12285,N_11749,N_11386);
nor U12286 (N_12286,N_11939,N_11618);
or U12287 (N_12287,N_11964,N_11430);
nand U12288 (N_12288,N_11561,N_11272);
nor U12289 (N_12289,N_11658,N_11598);
nand U12290 (N_12290,N_11382,N_11417);
nand U12291 (N_12291,N_11380,N_11552);
nor U12292 (N_12292,N_11583,N_11281);
and U12293 (N_12293,N_11654,N_11570);
nand U12294 (N_12294,N_11862,N_11846);
xnor U12295 (N_12295,N_11352,N_11744);
and U12296 (N_12296,N_11524,N_11629);
or U12297 (N_12297,N_11991,N_11467);
or U12298 (N_12298,N_11842,N_11307);
xnor U12299 (N_12299,N_11274,N_11921);
or U12300 (N_12300,N_11263,N_11984);
and U12301 (N_12301,N_11690,N_11959);
or U12302 (N_12302,N_11558,N_11792);
nor U12303 (N_12303,N_11867,N_11745);
xor U12304 (N_12304,N_11888,N_11316);
or U12305 (N_12305,N_11925,N_11431);
or U12306 (N_12306,N_11546,N_11612);
xor U12307 (N_12307,N_11394,N_11507);
or U12308 (N_12308,N_11495,N_11730);
or U12309 (N_12309,N_11737,N_11493);
or U12310 (N_12310,N_11428,N_11509);
nor U12311 (N_12311,N_11836,N_11323);
nand U12312 (N_12312,N_11600,N_11909);
and U12313 (N_12313,N_11260,N_11400);
nand U12314 (N_12314,N_11258,N_11781);
nor U12315 (N_12315,N_11710,N_11397);
nor U12316 (N_12316,N_11719,N_11821);
or U12317 (N_12317,N_11628,N_11667);
xnor U12318 (N_12318,N_11424,N_11835);
or U12319 (N_12319,N_11463,N_11418);
nor U12320 (N_12320,N_11580,N_11594);
nor U12321 (N_12321,N_11727,N_11741);
or U12322 (N_12322,N_11859,N_11290);
nor U12323 (N_12323,N_11311,N_11762);
and U12324 (N_12324,N_11641,N_11448);
and U12325 (N_12325,N_11550,N_11902);
nor U12326 (N_12326,N_11315,N_11577);
nor U12327 (N_12327,N_11297,N_11739);
xor U12328 (N_12328,N_11691,N_11988);
and U12329 (N_12329,N_11601,N_11318);
nand U12330 (N_12330,N_11770,N_11346);
nand U12331 (N_12331,N_11500,N_11855);
xor U12332 (N_12332,N_11278,N_11851);
nor U12333 (N_12333,N_11514,N_11987);
and U12334 (N_12334,N_11747,N_11294);
and U12335 (N_12335,N_11856,N_11523);
and U12336 (N_12336,N_11885,N_11937);
xor U12337 (N_12337,N_11864,N_11671);
nor U12338 (N_12338,N_11806,N_11738);
and U12339 (N_12339,N_11718,N_11319);
nor U12340 (N_12340,N_11966,N_11852);
nor U12341 (N_12341,N_11605,N_11445);
xor U12342 (N_12342,N_11697,N_11863);
nor U12343 (N_12343,N_11679,N_11354);
and U12344 (N_12344,N_11567,N_11854);
xnor U12345 (N_12345,N_11389,N_11894);
nor U12346 (N_12346,N_11257,N_11464);
nand U12347 (N_12347,N_11884,N_11291);
or U12348 (N_12348,N_11590,N_11461);
nor U12349 (N_12349,N_11269,N_11837);
and U12350 (N_12350,N_11587,N_11535);
or U12351 (N_12351,N_11904,N_11279);
and U12352 (N_12352,N_11914,N_11520);
nand U12353 (N_12353,N_11845,N_11359);
or U12354 (N_12354,N_11917,N_11989);
xnor U12355 (N_12355,N_11860,N_11790);
or U12356 (N_12356,N_11414,N_11824);
nor U12357 (N_12357,N_11831,N_11345);
nand U12358 (N_12358,N_11393,N_11695);
xor U12359 (N_12359,N_11809,N_11582);
or U12360 (N_12360,N_11327,N_11755);
xnor U12361 (N_12361,N_11771,N_11640);
nand U12362 (N_12362,N_11733,N_11622);
nand U12363 (N_12363,N_11996,N_11676);
xnor U12364 (N_12364,N_11292,N_11944);
nor U12365 (N_12365,N_11808,N_11259);
and U12366 (N_12366,N_11344,N_11803);
xor U12367 (N_12367,N_11795,N_11403);
nand U12368 (N_12368,N_11511,N_11995);
xnor U12369 (N_12369,N_11407,N_11650);
nor U12370 (N_12370,N_11887,N_11328);
or U12371 (N_12371,N_11827,N_11370);
or U12372 (N_12372,N_11469,N_11807);
nand U12373 (N_12373,N_11615,N_11367);
nor U12374 (N_12374,N_11910,N_11965);
xnor U12375 (N_12375,N_11332,N_11391);
or U12376 (N_12376,N_11396,N_11687);
nor U12377 (N_12377,N_11776,N_11684);
nor U12378 (N_12378,N_11960,N_11403);
nor U12379 (N_12379,N_11680,N_11511);
or U12380 (N_12380,N_11844,N_11675);
nand U12381 (N_12381,N_11805,N_11726);
nand U12382 (N_12382,N_11831,N_11464);
nor U12383 (N_12383,N_11764,N_11361);
or U12384 (N_12384,N_11323,N_11845);
or U12385 (N_12385,N_11927,N_11611);
or U12386 (N_12386,N_11841,N_11423);
or U12387 (N_12387,N_11490,N_11585);
nand U12388 (N_12388,N_11796,N_11288);
and U12389 (N_12389,N_11898,N_11552);
and U12390 (N_12390,N_11828,N_11615);
nand U12391 (N_12391,N_11607,N_11850);
or U12392 (N_12392,N_11627,N_11325);
nand U12393 (N_12393,N_11354,N_11376);
and U12394 (N_12394,N_11828,N_11661);
xor U12395 (N_12395,N_11863,N_11688);
or U12396 (N_12396,N_11859,N_11971);
and U12397 (N_12397,N_11655,N_11895);
and U12398 (N_12398,N_11744,N_11829);
nand U12399 (N_12399,N_11916,N_11384);
xnor U12400 (N_12400,N_11740,N_11565);
and U12401 (N_12401,N_11581,N_11622);
nand U12402 (N_12402,N_11798,N_11826);
xor U12403 (N_12403,N_11818,N_11349);
xor U12404 (N_12404,N_11537,N_11828);
and U12405 (N_12405,N_11600,N_11434);
nor U12406 (N_12406,N_11807,N_11498);
xor U12407 (N_12407,N_11370,N_11803);
xor U12408 (N_12408,N_11585,N_11826);
nor U12409 (N_12409,N_11629,N_11667);
nand U12410 (N_12410,N_11941,N_11321);
xor U12411 (N_12411,N_11956,N_11895);
or U12412 (N_12412,N_11670,N_11784);
and U12413 (N_12413,N_11335,N_11957);
nor U12414 (N_12414,N_11852,N_11761);
xor U12415 (N_12415,N_11590,N_11534);
xor U12416 (N_12416,N_11922,N_11262);
nand U12417 (N_12417,N_11805,N_11510);
or U12418 (N_12418,N_11447,N_11285);
or U12419 (N_12419,N_11629,N_11583);
xnor U12420 (N_12420,N_11297,N_11631);
xor U12421 (N_12421,N_11655,N_11857);
nand U12422 (N_12422,N_11773,N_11590);
or U12423 (N_12423,N_11282,N_11648);
xor U12424 (N_12424,N_11805,N_11766);
nand U12425 (N_12425,N_11507,N_11658);
nand U12426 (N_12426,N_11736,N_11638);
xor U12427 (N_12427,N_11325,N_11472);
and U12428 (N_12428,N_11389,N_11879);
or U12429 (N_12429,N_11642,N_11406);
nand U12430 (N_12430,N_11859,N_11719);
xnor U12431 (N_12431,N_11513,N_11687);
xor U12432 (N_12432,N_11401,N_11727);
or U12433 (N_12433,N_11799,N_11291);
nor U12434 (N_12434,N_11680,N_11908);
xnor U12435 (N_12435,N_11693,N_11548);
and U12436 (N_12436,N_11813,N_11622);
nor U12437 (N_12437,N_11451,N_11650);
or U12438 (N_12438,N_11564,N_11865);
nand U12439 (N_12439,N_11955,N_11830);
nor U12440 (N_12440,N_11881,N_11569);
nor U12441 (N_12441,N_11386,N_11488);
nand U12442 (N_12442,N_11468,N_11952);
or U12443 (N_12443,N_11920,N_11780);
or U12444 (N_12444,N_11637,N_11813);
nor U12445 (N_12445,N_11402,N_11418);
xor U12446 (N_12446,N_11543,N_11362);
or U12447 (N_12447,N_11343,N_11727);
or U12448 (N_12448,N_11306,N_11910);
or U12449 (N_12449,N_11852,N_11699);
or U12450 (N_12450,N_11416,N_11711);
or U12451 (N_12451,N_11428,N_11308);
xnor U12452 (N_12452,N_11761,N_11907);
and U12453 (N_12453,N_11345,N_11745);
xnor U12454 (N_12454,N_11828,N_11853);
nand U12455 (N_12455,N_11738,N_11938);
nor U12456 (N_12456,N_11257,N_11890);
nor U12457 (N_12457,N_11719,N_11788);
nor U12458 (N_12458,N_11550,N_11674);
nand U12459 (N_12459,N_11542,N_11763);
nor U12460 (N_12460,N_11596,N_11834);
and U12461 (N_12461,N_11773,N_11974);
or U12462 (N_12462,N_11767,N_11361);
nor U12463 (N_12463,N_11990,N_11398);
nand U12464 (N_12464,N_11386,N_11325);
nor U12465 (N_12465,N_11726,N_11708);
xor U12466 (N_12466,N_11335,N_11580);
nor U12467 (N_12467,N_11363,N_11717);
nand U12468 (N_12468,N_11286,N_11545);
or U12469 (N_12469,N_11650,N_11767);
or U12470 (N_12470,N_11834,N_11416);
nor U12471 (N_12471,N_11458,N_11769);
nor U12472 (N_12472,N_11916,N_11639);
or U12473 (N_12473,N_11683,N_11543);
xnor U12474 (N_12474,N_11650,N_11750);
or U12475 (N_12475,N_11799,N_11941);
nand U12476 (N_12476,N_11568,N_11765);
nand U12477 (N_12477,N_11489,N_11483);
xor U12478 (N_12478,N_11770,N_11680);
nor U12479 (N_12479,N_11650,N_11600);
nand U12480 (N_12480,N_11712,N_11472);
nor U12481 (N_12481,N_11924,N_11734);
xnor U12482 (N_12482,N_11953,N_11295);
nor U12483 (N_12483,N_11974,N_11317);
or U12484 (N_12484,N_11832,N_11379);
or U12485 (N_12485,N_11440,N_11878);
or U12486 (N_12486,N_11459,N_11627);
nand U12487 (N_12487,N_11632,N_11935);
xnor U12488 (N_12488,N_11549,N_11627);
and U12489 (N_12489,N_11978,N_11576);
nor U12490 (N_12490,N_11921,N_11430);
or U12491 (N_12491,N_11854,N_11664);
nand U12492 (N_12492,N_11580,N_11947);
nand U12493 (N_12493,N_11329,N_11706);
or U12494 (N_12494,N_11953,N_11806);
nand U12495 (N_12495,N_11849,N_11755);
or U12496 (N_12496,N_11272,N_11444);
or U12497 (N_12497,N_11832,N_11426);
xor U12498 (N_12498,N_11607,N_11359);
nor U12499 (N_12499,N_11380,N_11935);
or U12500 (N_12500,N_11587,N_11330);
nor U12501 (N_12501,N_11423,N_11726);
and U12502 (N_12502,N_11303,N_11279);
and U12503 (N_12503,N_11743,N_11711);
and U12504 (N_12504,N_11996,N_11981);
or U12505 (N_12505,N_11713,N_11884);
or U12506 (N_12506,N_11764,N_11491);
nand U12507 (N_12507,N_11862,N_11829);
xnor U12508 (N_12508,N_11913,N_11918);
xnor U12509 (N_12509,N_11652,N_11321);
xnor U12510 (N_12510,N_11929,N_11654);
and U12511 (N_12511,N_11519,N_11866);
nor U12512 (N_12512,N_11685,N_11317);
and U12513 (N_12513,N_11519,N_11426);
or U12514 (N_12514,N_11889,N_11291);
nand U12515 (N_12515,N_11377,N_11686);
and U12516 (N_12516,N_11555,N_11587);
nand U12517 (N_12517,N_11761,N_11758);
xnor U12518 (N_12518,N_11944,N_11412);
and U12519 (N_12519,N_11629,N_11809);
or U12520 (N_12520,N_11794,N_11347);
or U12521 (N_12521,N_11621,N_11423);
nand U12522 (N_12522,N_11692,N_11530);
and U12523 (N_12523,N_11666,N_11704);
nand U12524 (N_12524,N_11724,N_11777);
xor U12525 (N_12525,N_11754,N_11662);
or U12526 (N_12526,N_11950,N_11861);
and U12527 (N_12527,N_11328,N_11915);
nand U12528 (N_12528,N_11907,N_11614);
and U12529 (N_12529,N_11798,N_11277);
nand U12530 (N_12530,N_11919,N_11818);
nor U12531 (N_12531,N_11367,N_11687);
or U12532 (N_12532,N_11862,N_11920);
xnor U12533 (N_12533,N_11759,N_11955);
or U12534 (N_12534,N_11655,N_11583);
nand U12535 (N_12535,N_11375,N_11274);
xnor U12536 (N_12536,N_11447,N_11855);
xnor U12537 (N_12537,N_11365,N_11270);
nor U12538 (N_12538,N_11350,N_11965);
xnor U12539 (N_12539,N_11549,N_11929);
nor U12540 (N_12540,N_11313,N_11919);
nand U12541 (N_12541,N_11464,N_11427);
or U12542 (N_12542,N_11418,N_11946);
or U12543 (N_12543,N_11528,N_11542);
nor U12544 (N_12544,N_11552,N_11749);
nand U12545 (N_12545,N_11511,N_11730);
xnor U12546 (N_12546,N_11880,N_11416);
and U12547 (N_12547,N_11504,N_11718);
nor U12548 (N_12548,N_11632,N_11873);
and U12549 (N_12549,N_11865,N_11870);
nor U12550 (N_12550,N_11998,N_11823);
nor U12551 (N_12551,N_11684,N_11957);
or U12552 (N_12552,N_11280,N_11595);
xnor U12553 (N_12553,N_11736,N_11605);
nor U12554 (N_12554,N_11376,N_11803);
nor U12555 (N_12555,N_11860,N_11421);
or U12556 (N_12556,N_11444,N_11659);
xnor U12557 (N_12557,N_11534,N_11651);
nand U12558 (N_12558,N_11294,N_11859);
nand U12559 (N_12559,N_11444,N_11632);
nor U12560 (N_12560,N_11981,N_11483);
or U12561 (N_12561,N_11723,N_11802);
xor U12562 (N_12562,N_11546,N_11485);
and U12563 (N_12563,N_11405,N_11886);
xnor U12564 (N_12564,N_11636,N_11615);
and U12565 (N_12565,N_11723,N_11984);
or U12566 (N_12566,N_11843,N_11995);
xor U12567 (N_12567,N_11468,N_11694);
or U12568 (N_12568,N_11269,N_11842);
xnor U12569 (N_12569,N_11522,N_11312);
xnor U12570 (N_12570,N_11453,N_11884);
nor U12571 (N_12571,N_11905,N_11339);
nand U12572 (N_12572,N_11690,N_11547);
and U12573 (N_12573,N_11887,N_11850);
nand U12574 (N_12574,N_11796,N_11811);
xor U12575 (N_12575,N_11612,N_11524);
xor U12576 (N_12576,N_11924,N_11976);
and U12577 (N_12577,N_11604,N_11891);
xor U12578 (N_12578,N_11367,N_11564);
nor U12579 (N_12579,N_11716,N_11720);
nand U12580 (N_12580,N_11668,N_11260);
and U12581 (N_12581,N_11732,N_11497);
nor U12582 (N_12582,N_11298,N_11824);
or U12583 (N_12583,N_11835,N_11934);
nor U12584 (N_12584,N_11920,N_11356);
nand U12585 (N_12585,N_11583,N_11439);
nor U12586 (N_12586,N_11281,N_11820);
or U12587 (N_12587,N_11516,N_11409);
and U12588 (N_12588,N_11926,N_11615);
or U12589 (N_12589,N_11663,N_11794);
or U12590 (N_12590,N_11876,N_11430);
xor U12591 (N_12591,N_11602,N_11313);
and U12592 (N_12592,N_11416,N_11657);
nor U12593 (N_12593,N_11828,N_11978);
and U12594 (N_12594,N_11431,N_11263);
or U12595 (N_12595,N_11697,N_11583);
nand U12596 (N_12596,N_11571,N_11978);
and U12597 (N_12597,N_11319,N_11567);
and U12598 (N_12598,N_11450,N_11768);
xor U12599 (N_12599,N_11946,N_11279);
nor U12600 (N_12600,N_11755,N_11912);
nand U12601 (N_12601,N_11790,N_11964);
nor U12602 (N_12602,N_11472,N_11522);
nor U12603 (N_12603,N_11982,N_11927);
and U12604 (N_12604,N_11965,N_11489);
xnor U12605 (N_12605,N_11975,N_11276);
nand U12606 (N_12606,N_11342,N_11822);
and U12607 (N_12607,N_11575,N_11917);
nand U12608 (N_12608,N_11796,N_11685);
and U12609 (N_12609,N_11866,N_11951);
nor U12610 (N_12610,N_11355,N_11485);
nor U12611 (N_12611,N_11393,N_11510);
nand U12612 (N_12612,N_11454,N_11406);
nand U12613 (N_12613,N_11709,N_11716);
and U12614 (N_12614,N_11545,N_11436);
or U12615 (N_12615,N_11342,N_11977);
xor U12616 (N_12616,N_11456,N_11988);
and U12617 (N_12617,N_11846,N_11443);
nand U12618 (N_12618,N_11291,N_11308);
or U12619 (N_12619,N_11862,N_11315);
nand U12620 (N_12620,N_11927,N_11532);
nor U12621 (N_12621,N_11310,N_11590);
nor U12622 (N_12622,N_11421,N_11641);
xor U12623 (N_12623,N_11977,N_11412);
or U12624 (N_12624,N_11439,N_11723);
and U12625 (N_12625,N_11631,N_11450);
or U12626 (N_12626,N_11816,N_11674);
nand U12627 (N_12627,N_11351,N_11707);
or U12628 (N_12628,N_11468,N_11949);
or U12629 (N_12629,N_11695,N_11995);
xor U12630 (N_12630,N_11448,N_11650);
and U12631 (N_12631,N_11451,N_11506);
nor U12632 (N_12632,N_11453,N_11797);
nor U12633 (N_12633,N_11673,N_11496);
xnor U12634 (N_12634,N_11691,N_11734);
or U12635 (N_12635,N_11782,N_11444);
xnor U12636 (N_12636,N_11910,N_11429);
nand U12637 (N_12637,N_11743,N_11937);
nand U12638 (N_12638,N_11357,N_11553);
nor U12639 (N_12639,N_11316,N_11594);
nand U12640 (N_12640,N_11969,N_11597);
or U12641 (N_12641,N_11963,N_11772);
nand U12642 (N_12642,N_11290,N_11653);
xor U12643 (N_12643,N_11817,N_11854);
xnor U12644 (N_12644,N_11351,N_11279);
xnor U12645 (N_12645,N_11584,N_11264);
nand U12646 (N_12646,N_11838,N_11517);
and U12647 (N_12647,N_11369,N_11263);
and U12648 (N_12648,N_11891,N_11818);
or U12649 (N_12649,N_11352,N_11930);
and U12650 (N_12650,N_11925,N_11794);
and U12651 (N_12651,N_11514,N_11624);
nand U12652 (N_12652,N_11982,N_11703);
nor U12653 (N_12653,N_11936,N_11884);
nor U12654 (N_12654,N_11511,N_11858);
xor U12655 (N_12655,N_11452,N_11391);
or U12656 (N_12656,N_11402,N_11860);
xor U12657 (N_12657,N_11533,N_11282);
nor U12658 (N_12658,N_11716,N_11270);
nor U12659 (N_12659,N_11953,N_11601);
and U12660 (N_12660,N_11830,N_11677);
xor U12661 (N_12661,N_11427,N_11689);
nor U12662 (N_12662,N_11761,N_11574);
and U12663 (N_12663,N_11612,N_11505);
xor U12664 (N_12664,N_11259,N_11705);
xnor U12665 (N_12665,N_11573,N_11473);
xnor U12666 (N_12666,N_11603,N_11261);
and U12667 (N_12667,N_11339,N_11359);
nor U12668 (N_12668,N_11567,N_11658);
or U12669 (N_12669,N_11374,N_11895);
nand U12670 (N_12670,N_11495,N_11571);
and U12671 (N_12671,N_11788,N_11284);
or U12672 (N_12672,N_11339,N_11816);
xnor U12673 (N_12673,N_11924,N_11956);
nand U12674 (N_12674,N_11979,N_11854);
nand U12675 (N_12675,N_11755,N_11831);
and U12676 (N_12676,N_11703,N_11821);
nand U12677 (N_12677,N_11473,N_11721);
nand U12678 (N_12678,N_11971,N_11311);
xnor U12679 (N_12679,N_11316,N_11320);
nand U12680 (N_12680,N_11765,N_11773);
nand U12681 (N_12681,N_11754,N_11820);
or U12682 (N_12682,N_11861,N_11386);
nor U12683 (N_12683,N_11397,N_11365);
or U12684 (N_12684,N_11549,N_11780);
and U12685 (N_12685,N_11492,N_11470);
and U12686 (N_12686,N_11310,N_11309);
nand U12687 (N_12687,N_11755,N_11564);
and U12688 (N_12688,N_11552,N_11850);
xor U12689 (N_12689,N_11888,N_11597);
xnor U12690 (N_12690,N_11944,N_11700);
nand U12691 (N_12691,N_11451,N_11493);
and U12692 (N_12692,N_11360,N_11354);
nor U12693 (N_12693,N_11703,N_11440);
nor U12694 (N_12694,N_11681,N_11468);
and U12695 (N_12695,N_11412,N_11994);
or U12696 (N_12696,N_11290,N_11660);
xor U12697 (N_12697,N_11766,N_11294);
or U12698 (N_12698,N_11707,N_11600);
xnor U12699 (N_12699,N_11550,N_11792);
or U12700 (N_12700,N_11488,N_11625);
and U12701 (N_12701,N_11741,N_11773);
xnor U12702 (N_12702,N_11717,N_11920);
nor U12703 (N_12703,N_11440,N_11798);
nor U12704 (N_12704,N_11436,N_11899);
and U12705 (N_12705,N_11955,N_11966);
or U12706 (N_12706,N_11638,N_11416);
or U12707 (N_12707,N_11605,N_11985);
or U12708 (N_12708,N_11335,N_11854);
nor U12709 (N_12709,N_11855,N_11423);
and U12710 (N_12710,N_11355,N_11931);
nor U12711 (N_12711,N_11829,N_11745);
nor U12712 (N_12712,N_11902,N_11529);
nor U12713 (N_12713,N_11392,N_11439);
xnor U12714 (N_12714,N_11421,N_11254);
xor U12715 (N_12715,N_11615,N_11470);
or U12716 (N_12716,N_11267,N_11777);
nand U12717 (N_12717,N_11338,N_11251);
or U12718 (N_12718,N_11378,N_11275);
or U12719 (N_12719,N_11372,N_11729);
nor U12720 (N_12720,N_11925,N_11468);
nand U12721 (N_12721,N_11920,N_11600);
nor U12722 (N_12722,N_11715,N_11590);
xnor U12723 (N_12723,N_11256,N_11859);
and U12724 (N_12724,N_11474,N_11642);
nor U12725 (N_12725,N_11983,N_11851);
nand U12726 (N_12726,N_11677,N_11747);
and U12727 (N_12727,N_11708,N_11816);
and U12728 (N_12728,N_11649,N_11271);
nor U12729 (N_12729,N_11419,N_11937);
and U12730 (N_12730,N_11281,N_11847);
xor U12731 (N_12731,N_11911,N_11555);
or U12732 (N_12732,N_11878,N_11307);
or U12733 (N_12733,N_11804,N_11908);
nand U12734 (N_12734,N_11909,N_11507);
or U12735 (N_12735,N_11550,N_11369);
nor U12736 (N_12736,N_11824,N_11291);
nor U12737 (N_12737,N_11553,N_11373);
nor U12738 (N_12738,N_11823,N_11588);
nor U12739 (N_12739,N_11666,N_11424);
or U12740 (N_12740,N_11567,N_11562);
nand U12741 (N_12741,N_11571,N_11306);
xor U12742 (N_12742,N_11299,N_11520);
nand U12743 (N_12743,N_11329,N_11630);
and U12744 (N_12744,N_11741,N_11575);
nand U12745 (N_12745,N_11692,N_11332);
nor U12746 (N_12746,N_11765,N_11769);
nor U12747 (N_12747,N_11846,N_11969);
xnor U12748 (N_12748,N_11512,N_11731);
or U12749 (N_12749,N_11662,N_11736);
nand U12750 (N_12750,N_12608,N_12376);
and U12751 (N_12751,N_12749,N_12296);
nand U12752 (N_12752,N_12463,N_12494);
xnor U12753 (N_12753,N_12212,N_12012);
nor U12754 (N_12754,N_12254,N_12439);
and U12755 (N_12755,N_12113,N_12028);
xor U12756 (N_12756,N_12442,N_12483);
and U12757 (N_12757,N_12189,N_12098);
nand U12758 (N_12758,N_12378,N_12214);
nor U12759 (N_12759,N_12509,N_12050);
xor U12760 (N_12760,N_12153,N_12635);
xor U12761 (N_12761,N_12404,N_12495);
xor U12762 (N_12762,N_12419,N_12699);
and U12763 (N_12763,N_12106,N_12628);
xnor U12764 (N_12764,N_12530,N_12643);
and U12765 (N_12765,N_12338,N_12625);
nor U12766 (N_12766,N_12668,N_12232);
nand U12767 (N_12767,N_12058,N_12267);
nor U12768 (N_12768,N_12728,N_12662);
and U12769 (N_12769,N_12371,N_12229);
or U12770 (N_12770,N_12335,N_12682);
or U12771 (N_12771,N_12710,N_12572);
and U12772 (N_12772,N_12131,N_12285);
and U12773 (N_12773,N_12745,N_12155);
nand U12774 (N_12774,N_12319,N_12422);
nor U12775 (N_12775,N_12451,N_12248);
nand U12776 (N_12776,N_12041,N_12708);
nor U12777 (N_12777,N_12362,N_12427);
nand U12778 (N_12778,N_12613,N_12271);
or U12779 (N_12779,N_12262,N_12421);
nor U12780 (N_12780,N_12533,N_12581);
and U12781 (N_12781,N_12353,N_12663);
xnor U12782 (N_12782,N_12377,N_12257);
or U12783 (N_12783,N_12301,N_12316);
nor U12784 (N_12784,N_12469,N_12460);
nand U12785 (N_12785,N_12722,N_12644);
xor U12786 (N_12786,N_12182,N_12083);
xnor U12787 (N_12787,N_12206,N_12243);
nand U12788 (N_12788,N_12748,N_12132);
nand U12789 (N_12789,N_12430,N_12357);
nor U12790 (N_12790,N_12691,N_12160);
nand U12791 (N_12791,N_12033,N_12194);
or U12792 (N_12792,N_12384,N_12448);
or U12793 (N_12793,N_12230,N_12096);
and U12794 (N_12794,N_12547,N_12679);
or U12795 (N_12795,N_12388,N_12688);
nor U12796 (N_12796,N_12031,N_12087);
nand U12797 (N_12797,N_12200,N_12245);
and U12798 (N_12798,N_12361,N_12555);
and U12799 (N_12799,N_12350,N_12081);
nor U12800 (N_12800,N_12345,N_12615);
and U12801 (N_12801,N_12524,N_12619);
nand U12802 (N_12802,N_12225,N_12544);
nand U12803 (N_12803,N_12649,N_12346);
xor U12804 (N_12804,N_12702,N_12193);
xnor U12805 (N_12805,N_12043,N_12008);
or U12806 (N_12806,N_12094,N_12284);
or U12807 (N_12807,N_12228,N_12409);
nor U12808 (N_12808,N_12030,N_12576);
and U12809 (N_12809,N_12372,N_12580);
nor U12810 (N_12810,N_12671,N_12542);
nand U12811 (N_12811,N_12501,N_12486);
and U12812 (N_12812,N_12076,N_12648);
nor U12813 (N_12813,N_12569,N_12412);
nand U12814 (N_12814,N_12235,N_12307);
xnor U12815 (N_12815,N_12575,N_12612);
nor U12816 (N_12816,N_12700,N_12201);
and U12817 (N_12817,N_12017,N_12253);
nand U12818 (N_12818,N_12694,N_12207);
and U12819 (N_12819,N_12603,N_12443);
or U12820 (N_12820,N_12147,N_12027);
xnor U12821 (N_12821,N_12173,N_12592);
nor U12822 (N_12822,N_12393,N_12016);
nor U12823 (N_12823,N_12598,N_12221);
and U12824 (N_12824,N_12269,N_12610);
or U12825 (N_12825,N_12310,N_12117);
xor U12826 (N_12826,N_12666,N_12367);
nor U12827 (N_12827,N_12046,N_12684);
nor U12828 (N_12828,N_12109,N_12716);
or U12829 (N_12829,N_12312,N_12244);
or U12830 (N_12830,N_12045,N_12311);
xnor U12831 (N_12831,N_12313,N_12291);
nand U12832 (N_12832,N_12480,N_12647);
and U12833 (N_12833,N_12713,N_12392);
nand U12834 (N_12834,N_12134,N_12192);
nand U12835 (N_12835,N_12366,N_12237);
nor U12836 (N_12836,N_12018,N_12162);
and U12837 (N_12837,N_12185,N_12519);
or U12838 (N_12838,N_12434,N_12557);
or U12839 (N_12839,N_12239,N_12064);
or U12840 (N_12840,N_12508,N_12633);
and U12841 (N_12841,N_12139,N_12156);
xor U12842 (N_12842,N_12154,N_12698);
xor U12843 (N_12843,N_12099,N_12420);
and U12844 (N_12844,N_12681,N_12596);
or U12845 (N_12845,N_12616,N_12079);
xnor U12846 (N_12846,N_12329,N_12072);
and U12847 (N_12847,N_12704,N_12145);
and U12848 (N_12848,N_12102,N_12341);
nor U12849 (N_12849,N_12082,N_12303);
nor U12850 (N_12850,N_12656,N_12258);
and U12851 (N_12851,N_12013,N_12578);
nor U12852 (N_12852,N_12732,N_12223);
nor U12853 (N_12853,N_12380,N_12274);
xor U12854 (N_12854,N_12373,N_12571);
nor U12855 (N_12855,N_12288,N_12693);
nor U12856 (N_12856,N_12276,N_12188);
xor U12857 (N_12857,N_12078,N_12405);
nor U12858 (N_12858,N_12548,N_12023);
nor U12859 (N_12859,N_12044,N_12523);
nor U12860 (N_12860,N_12461,N_12573);
nand U12861 (N_12861,N_12715,N_12141);
and U12862 (N_12862,N_12462,N_12455);
or U12863 (N_12863,N_12263,N_12747);
nor U12864 (N_12864,N_12306,N_12642);
and U12865 (N_12865,N_12652,N_12720);
and U12866 (N_12866,N_12231,N_12560);
or U12867 (N_12867,N_12414,N_12309);
xnor U12868 (N_12868,N_12181,N_12056);
nor U12869 (N_12869,N_12165,N_12163);
and U12870 (N_12870,N_12665,N_12426);
nand U12871 (N_12871,N_12279,N_12100);
or U12872 (N_12872,N_12124,N_12600);
or U12873 (N_12873,N_12559,N_12204);
and U12874 (N_12874,N_12042,N_12746);
and U12875 (N_12875,N_12342,N_12111);
or U12876 (N_12876,N_12191,N_12048);
xnor U12877 (N_12877,N_12084,N_12609);
nor U12878 (N_12878,N_12391,N_12522);
nand U12879 (N_12879,N_12438,N_12019);
and U12880 (N_12880,N_12593,N_12352);
nor U12881 (N_12881,N_12157,N_12236);
nor U12882 (N_12882,N_12721,N_12112);
nand U12883 (N_12883,N_12707,N_12278);
nand U12884 (N_12884,N_12604,N_12539);
nand U12885 (N_12885,N_12205,N_12458);
or U12886 (N_12886,N_12742,N_12450);
and U12887 (N_12887,N_12097,N_12328);
nor U12888 (N_12888,N_12270,N_12088);
nor U12889 (N_12889,N_12020,N_12176);
and U12890 (N_12890,N_12537,N_12424);
and U12891 (N_12891,N_12007,N_12282);
and U12892 (N_12892,N_12227,N_12026);
or U12893 (N_12893,N_12242,N_12725);
nand U12894 (N_12894,N_12595,N_12300);
or U12895 (N_12895,N_12037,N_12472);
nor U12896 (N_12896,N_12068,N_12213);
nor U12897 (N_12897,N_12121,N_12401);
or U12898 (N_12898,N_12740,N_12314);
or U12899 (N_12899,N_12009,N_12375);
xnor U12900 (N_12900,N_12597,N_12622);
nor U12901 (N_12901,N_12203,N_12520);
xor U12902 (N_12902,N_12272,N_12340);
and U12903 (N_12903,N_12660,N_12219);
and U12904 (N_12904,N_12251,N_12063);
xor U12905 (N_12905,N_12585,N_12632);
nor U12906 (N_12906,N_12090,N_12621);
xor U12907 (N_12907,N_12122,N_12114);
xnor U12908 (N_12908,N_12677,N_12051);
nor U12909 (N_12909,N_12526,N_12158);
or U12910 (N_12910,N_12498,N_12432);
nand U12911 (N_12911,N_12680,N_12011);
xnor U12912 (N_12912,N_12718,N_12637);
or U12913 (N_12913,N_12172,N_12566);
nand U12914 (N_12914,N_12170,N_12387);
and U12915 (N_12915,N_12297,N_12260);
nor U12916 (N_12916,N_12567,N_12014);
and U12917 (N_12917,N_12607,N_12712);
and U12918 (N_12918,N_12075,N_12558);
xnor U12919 (N_12919,N_12330,N_12413);
nand U12920 (N_12920,N_12734,N_12292);
xor U12921 (N_12921,N_12453,N_12178);
or U12922 (N_12922,N_12151,N_12315);
xor U12923 (N_12923,N_12705,N_12743);
or U12924 (N_12924,N_12664,N_12323);
and U12925 (N_12925,N_12174,N_12324);
nor U12926 (N_12926,N_12266,N_12080);
xnor U12927 (N_12927,N_12479,N_12208);
nand U12928 (N_12928,N_12322,N_12727);
nor U12929 (N_12929,N_12126,N_12529);
or U12930 (N_12930,N_12510,N_12118);
xnor U12931 (N_12931,N_12629,N_12196);
xor U12932 (N_12932,N_12360,N_12059);
nor U12933 (N_12933,N_12645,N_12583);
and U12934 (N_12934,N_12137,N_12218);
nor U12935 (N_12935,N_12431,N_12354);
or U12936 (N_12936,N_12234,N_12085);
and U12937 (N_12937,N_12444,N_12128);
nor U12938 (N_12938,N_12395,N_12491);
nand U12939 (N_12939,N_12408,N_12478);
nor U12940 (N_12940,N_12369,N_12298);
and U12941 (N_12941,N_12249,N_12066);
nand U12942 (N_12942,N_12211,N_12689);
xnor U12943 (N_12943,N_12299,N_12657);
and U12944 (N_12944,N_12105,N_12611);
nor U12945 (N_12945,N_12073,N_12166);
nand U12946 (N_12946,N_12104,N_12737);
nand U12947 (N_12947,N_12029,N_12197);
and U12948 (N_12948,N_12654,N_12586);
nor U12949 (N_12949,N_12255,N_12714);
and U12950 (N_12950,N_12474,N_12636);
and U12951 (N_12951,N_12195,N_12568);
xor U12952 (N_12952,N_12717,N_12129);
and U12953 (N_12953,N_12209,N_12119);
or U12954 (N_12954,N_12302,N_12496);
nor U12955 (N_12955,N_12459,N_12565);
nor U12956 (N_12956,N_12464,N_12161);
or U12957 (N_12957,N_12475,N_12022);
or U12958 (N_12958,N_12120,N_12490);
nand U12959 (N_12959,N_12334,N_12488);
or U12960 (N_12960,N_12256,N_12482);
nand U12961 (N_12961,N_12418,N_12579);
xnor U12962 (N_12962,N_12074,N_12061);
or U12963 (N_12963,N_12445,N_12729);
nor U12964 (N_12964,N_12135,N_12744);
nand U12965 (N_12965,N_12040,N_12514);
and U12966 (N_12966,N_12452,N_12039);
xor U12967 (N_12967,N_12261,N_12731);
and U12968 (N_12968,N_12551,N_12626);
and U12969 (N_12969,N_12321,N_12674);
or U12970 (N_12970,N_12561,N_12473);
nand U12971 (N_12971,N_12423,N_12703);
or U12972 (N_12972,N_12187,N_12304);
nor U12973 (N_12973,N_12673,N_12407);
and U12974 (N_12974,N_12497,N_12400);
nor U12975 (N_12975,N_12183,N_12148);
or U12976 (N_12976,N_12325,N_12159);
or U12977 (N_12977,N_12133,N_12634);
or U12978 (N_12978,N_12351,N_12308);
xnor U12979 (N_12979,N_12277,N_12049);
nor U12980 (N_12980,N_12268,N_12365);
nor U12981 (N_12981,N_12339,N_12287);
nand U12982 (N_12982,N_12294,N_12525);
nor U12983 (N_12983,N_12184,N_12527);
xor U12984 (N_12984,N_12620,N_12021);
or U12985 (N_12985,N_12363,N_12317);
xor U12986 (N_12986,N_12487,N_12534);
xnor U12987 (N_12987,N_12541,N_12577);
nor U12988 (N_12988,N_12631,N_12247);
nor U12989 (N_12989,N_12676,N_12669);
xor U12990 (N_12990,N_12538,N_12252);
nor U12991 (N_12991,N_12347,N_12549);
nand U12992 (N_12992,N_12697,N_12108);
xor U12993 (N_12993,N_12146,N_12150);
nand U12994 (N_12994,N_12441,N_12553);
or U12995 (N_12995,N_12217,N_12695);
or U12996 (N_12996,N_12701,N_12499);
or U12997 (N_12997,N_12706,N_12617);
nor U12998 (N_12998,N_12331,N_12337);
nand U12999 (N_12999,N_12675,N_12429);
xnor U13000 (N_13000,N_12658,N_12374);
nor U13001 (N_13001,N_12167,N_12425);
nor U13002 (N_13002,N_12428,N_12103);
xnor U13003 (N_13003,N_12683,N_12326);
xor U13004 (N_13004,N_12741,N_12417);
and U13005 (N_13005,N_12723,N_12179);
nand U13006 (N_13006,N_12370,N_12069);
xor U13007 (N_13007,N_12506,N_12513);
nand U13008 (N_13008,N_12493,N_12053);
or U13009 (N_13009,N_12433,N_12259);
or U13010 (N_13010,N_12110,N_12368);
nand U13011 (N_13011,N_12588,N_12002);
nand U13012 (N_13012,N_12724,N_12359);
nor U13013 (N_13013,N_12152,N_12180);
nand U13014 (N_13014,N_12336,N_12032);
xnor U13015 (N_13015,N_12627,N_12071);
nand U13016 (N_13016,N_12327,N_12563);
and U13017 (N_13017,N_12504,N_12047);
nor U13018 (N_13018,N_12065,N_12564);
xnor U13019 (N_13019,N_12398,N_12403);
xnor U13020 (N_13020,N_12517,N_12457);
nand U13021 (N_13021,N_12599,N_12305);
or U13022 (N_13022,N_12385,N_12485);
or U13023 (N_13023,N_12436,N_12630);
xnor U13024 (N_13024,N_12562,N_12587);
nor U13025 (N_13025,N_12062,N_12171);
nor U13026 (N_13026,N_12005,N_12512);
or U13027 (N_13027,N_12397,N_12000);
nand U13028 (N_13028,N_12383,N_12659);
nand U13029 (N_13029,N_12574,N_12224);
xor U13030 (N_13030,N_12144,N_12736);
and U13031 (N_13031,N_12435,N_12690);
xor U13032 (N_13032,N_12216,N_12468);
nand U13033 (N_13033,N_12024,N_12006);
and U13034 (N_13034,N_12500,N_12550);
nor U13035 (N_13035,N_12003,N_12091);
xnor U13036 (N_13036,N_12531,N_12618);
nand U13037 (N_13037,N_12582,N_12624);
and U13038 (N_13038,N_12052,N_12015);
nor U13039 (N_13039,N_12246,N_12602);
nor U13040 (N_13040,N_12605,N_12670);
and U13041 (N_13041,N_12735,N_12601);
and U13042 (N_13042,N_12655,N_12025);
nand U13043 (N_13043,N_12343,N_12210);
or U13044 (N_13044,N_12169,N_12402);
nor U13045 (N_13045,N_12719,N_12467);
nand U13046 (N_13046,N_12730,N_12382);
nand U13047 (N_13047,N_12265,N_12589);
xor U13048 (N_13048,N_12381,N_12440);
or U13049 (N_13049,N_12502,N_12454);
xor U13050 (N_13050,N_12010,N_12416);
xor U13051 (N_13051,N_12686,N_12295);
and U13052 (N_13052,N_12465,N_12389);
or U13053 (N_13053,N_12358,N_12034);
nand U13054 (N_13054,N_12226,N_12484);
and U13055 (N_13055,N_12503,N_12142);
xnor U13056 (N_13056,N_12344,N_12738);
or U13057 (N_13057,N_12116,N_12198);
xnor U13058 (N_13058,N_12584,N_12515);
nor U13059 (N_13059,N_12687,N_12177);
nor U13060 (N_13060,N_12481,N_12623);
or U13061 (N_13061,N_12661,N_12552);
or U13062 (N_13062,N_12241,N_12250);
nand U13063 (N_13063,N_12471,N_12411);
nor U13064 (N_13064,N_12168,N_12115);
xor U13065 (N_13065,N_12275,N_12001);
xor U13066 (N_13066,N_12556,N_12641);
or U13067 (N_13067,N_12545,N_12726);
xnor U13068 (N_13068,N_12590,N_12492);
nand U13069 (N_13069,N_12280,N_12739);
or U13070 (N_13070,N_12386,N_12646);
or U13071 (N_13071,N_12415,N_12390);
or U13072 (N_13072,N_12543,N_12202);
or U13073 (N_13073,N_12220,N_12190);
nor U13074 (N_13074,N_12709,N_12692);
nand U13075 (N_13075,N_12678,N_12070);
xor U13076 (N_13076,N_12143,N_12399);
and U13077 (N_13077,N_12449,N_12651);
nand U13078 (N_13078,N_12470,N_12355);
xnor U13079 (N_13079,N_12238,N_12333);
nor U13080 (N_13080,N_12286,N_12518);
xnor U13081 (N_13081,N_12136,N_12004);
nor U13082 (N_13082,N_12149,N_12591);
and U13083 (N_13083,N_12614,N_12289);
xnor U13084 (N_13084,N_12290,N_12406);
nand U13085 (N_13085,N_12293,N_12396);
and U13086 (N_13086,N_12379,N_12233);
or U13087 (N_13087,N_12067,N_12650);
xnor U13088 (N_13088,N_12055,N_12077);
or U13089 (N_13089,N_12535,N_12038);
and U13090 (N_13090,N_12199,N_12095);
xnor U13091 (N_13091,N_12638,N_12511);
and U13092 (N_13092,N_12540,N_12318);
and U13093 (N_13093,N_12332,N_12036);
nand U13094 (N_13094,N_12507,N_12653);
nor U13095 (N_13095,N_12594,N_12639);
nand U13096 (N_13096,N_12127,N_12528);
nand U13097 (N_13097,N_12356,N_12093);
and U13098 (N_13098,N_12057,N_12505);
and U13099 (N_13099,N_12516,N_12283);
xnor U13100 (N_13100,N_12060,N_12546);
nand U13101 (N_13101,N_12521,N_12476);
and U13102 (N_13102,N_12281,N_12035);
nor U13103 (N_13103,N_12264,N_12733);
nand U13104 (N_13104,N_12054,N_12089);
xor U13105 (N_13105,N_12685,N_12536);
and U13106 (N_13106,N_12532,N_12466);
nor U13107 (N_13107,N_12711,N_12570);
nand U13108 (N_13108,N_12667,N_12125);
nor U13109 (N_13109,N_12186,N_12456);
or U13110 (N_13110,N_12086,N_12273);
and U13111 (N_13111,N_12696,N_12489);
nor U13112 (N_13112,N_12092,N_12240);
nor U13113 (N_13113,N_12477,N_12410);
xor U13114 (N_13114,N_12123,N_12222);
nor U13115 (N_13115,N_12672,N_12320);
or U13116 (N_13116,N_12394,N_12640);
or U13117 (N_13117,N_12447,N_12140);
or U13118 (N_13118,N_12107,N_12364);
xor U13119 (N_13119,N_12175,N_12164);
nand U13120 (N_13120,N_12215,N_12348);
nand U13121 (N_13121,N_12130,N_12101);
nor U13122 (N_13122,N_12138,N_12349);
or U13123 (N_13123,N_12446,N_12606);
or U13124 (N_13124,N_12554,N_12437);
nand U13125 (N_13125,N_12540,N_12748);
and U13126 (N_13126,N_12176,N_12043);
nor U13127 (N_13127,N_12685,N_12584);
xor U13128 (N_13128,N_12354,N_12445);
nor U13129 (N_13129,N_12448,N_12029);
xor U13130 (N_13130,N_12265,N_12519);
and U13131 (N_13131,N_12179,N_12196);
xor U13132 (N_13132,N_12533,N_12097);
nand U13133 (N_13133,N_12480,N_12205);
nor U13134 (N_13134,N_12084,N_12174);
or U13135 (N_13135,N_12178,N_12437);
xnor U13136 (N_13136,N_12601,N_12391);
nand U13137 (N_13137,N_12178,N_12363);
nor U13138 (N_13138,N_12106,N_12167);
nand U13139 (N_13139,N_12689,N_12165);
nand U13140 (N_13140,N_12453,N_12544);
nand U13141 (N_13141,N_12511,N_12123);
nor U13142 (N_13142,N_12120,N_12030);
nand U13143 (N_13143,N_12627,N_12366);
nor U13144 (N_13144,N_12277,N_12612);
nor U13145 (N_13145,N_12209,N_12386);
nand U13146 (N_13146,N_12636,N_12323);
and U13147 (N_13147,N_12371,N_12513);
or U13148 (N_13148,N_12251,N_12439);
or U13149 (N_13149,N_12338,N_12475);
or U13150 (N_13150,N_12014,N_12378);
xnor U13151 (N_13151,N_12215,N_12120);
nor U13152 (N_13152,N_12436,N_12487);
or U13153 (N_13153,N_12037,N_12249);
nand U13154 (N_13154,N_12033,N_12058);
xnor U13155 (N_13155,N_12203,N_12116);
nand U13156 (N_13156,N_12048,N_12279);
nand U13157 (N_13157,N_12313,N_12324);
nor U13158 (N_13158,N_12684,N_12543);
nand U13159 (N_13159,N_12745,N_12370);
nor U13160 (N_13160,N_12566,N_12514);
nor U13161 (N_13161,N_12121,N_12011);
nor U13162 (N_13162,N_12299,N_12646);
or U13163 (N_13163,N_12346,N_12188);
nand U13164 (N_13164,N_12705,N_12408);
nor U13165 (N_13165,N_12648,N_12275);
xnor U13166 (N_13166,N_12194,N_12437);
xor U13167 (N_13167,N_12047,N_12169);
nand U13168 (N_13168,N_12662,N_12317);
xor U13169 (N_13169,N_12728,N_12339);
nor U13170 (N_13170,N_12747,N_12332);
nand U13171 (N_13171,N_12222,N_12596);
or U13172 (N_13172,N_12516,N_12089);
nor U13173 (N_13173,N_12703,N_12509);
and U13174 (N_13174,N_12049,N_12596);
and U13175 (N_13175,N_12105,N_12652);
nor U13176 (N_13176,N_12304,N_12660);
or U13177 (N_13177,N_12027,N_12221);
nand U13178 (N_13178,N_12308,N_12438);
xor U13179 (N_13179,N_12442,N_12109);
and U13180 (N_13180,N_12171,N_12339);
and U13181 (N_13181,N_12650,N_12292);
nor U13182 (N_13182,N_12116,N_12445);
nor U13183 (N_13183,N_12193,N_12232);
nor U13184 (N_13184,N_12016,N_12411);
nand U13185 (N_13185,N_12244,N_12501);
or U13186 (N_13186,N_12378,N_12202);
xnor U13187 (N_13187,N_12140,N_12644);
xnor U13188 (N_13188,N_12105,N_12005);
and U13189 (N_13189,N_12469,N_12620);
nand U13190 (N_13190,N_12088,N_12173);
nand U13191 (N_13191,N_12008,N_12482);
xor U13192 (N_13192,N_12730,N_12083);
or U13193 (N_13193,N_12005,N_12694);
nor U13194 (N_13194,N_12438,N_12439);
nand U13195 (N_13195,N_12229,N_12710);
or U13196 (N_13196,N_12625,N_12559);
nor U13197 (N_13197,N_12381,N_12718);
xor U13198 (N_13198,N_12460,N_12711);
and U13199 (N_13199,N_12386,N_12032);
and U13200 (N_13200,N_12027,N_12115);
xor U13201 (N_13201,N_12596,N_12331);
and U13202 (N_13202,N_12715,N_12738);
nand U13203 (N_13203,N_12295,N_12420);
and U13204 (N_13204,N_12342,N_12457);
nand U13205 (N_13205,N_12728,N_12025);
or U13206 (N_13206,N_12273,N_12052);
and U13207 (N_13207,N_12458,N_12443);
nor U13208 (N_13208,N_12557,N_12607);
and U13209 (N_13209,N_12247,N_12441);
nand U13210 (N_13210,N_12552,N_12024);
or U13211 (N_13211,N_12120,N_12123);
xnor U13212 (N_13212,N_12586,N_12213);
nand U13213 (N_13213,N_12407,N_12685);
nor U13214 (N_13214,N_12136,N_12586);
and U13215 (N_13215,N_12387,N_12184);
nor U13216 (N_13216,N_12226,N_12682);
and U13217 (N_13217,N_12337,N_12404);
nand U13218 (N_13218,N_12669,N_12526);
nand U13219 (N_13219,N_12063,N_12709);
or U13220 (N_13220,N_12593,N_12283);
or U13221 (N_13221,N_12152,N_12658);
and U13222 (N_13222,N_12424,N_12715);
nand U13223 (N_13223,N_12473,N_12466);
xor U13224 (N_13224,N_12410,N_12392);
nor U13225 (N_13225,N_12122,N_12193);
xnor U13226 (N_13226,N_12708,N_12536);
and U13227 (N_13227,N_12680,N_12630);
or U13228 (N_13228,N_12689,N_12357);
nand U13229 (N_13229,N_12030,N_12041);
nand U13230 (N_13230,N_12195,N_12737);
and U13231 (N_13231,N_12293,N_12356);
nand U13232 (N_13232,N_12594,N_12302);
or U13233 (N_13233,N_12667,N_12671);
and U13234 (N_13234,N_12568,N_12541);
or U13235 (N_13235,N_12019,N_12390);
and U13236 (N_13236,N_12172,N_12526);
nor U13237 (N_13237,N_12041,N_12435);
nor U13238 (N_13238,N_12341,N_12184);
or U13239 (N_13239,N_12214,N_12041);
or U13240 (N_13240,N_12479,N_12042);
nor U13241 (N_13241,N_12047,N_12103);
nand U13242 (N_13242,N_12509,N_12268);
or U13243 (N_13243,N_12663,N_12674);
xor U13244 (N_13244,N_12455,N_12344);
and U13245 (N_13245,N_12626,N_12706);
nor U13246 (N_13246,N_12254,N_12337);
nand U13247 (N_13247,N_12703,N_12604);
and U13248 (N_13248,N_12481,N_12582);
nor U13249 (N_13249,N_12289,N_12662);
nor U13250 (N_13250,N_12584,N_12249);
xor U13251 (N_13251,N_12121,N_12654);
and U13252 (N_13252,N_12000,N_12620);
nor U13253 (N_13253,N_12510,N_12651);
nor U13254 (N_13254,N_12749,N_12434);
xor U13255 (N_13255,N_12176,N_12078);
nor U13256 (N_13256,N_12260,N_12411);
nand U13257 (N_13257,N_12649,N_12701);
xnor U13258 (N_13258,N_12574,N_12705);
nand U13259 (N_13259,N_12737,N_12420);
or U13260 (N_13260,N_12449,N_12246);
xnor U13261 (N_13261,N_12377,N_12077);
or U13262 (N_13262,N_12209,N_12251);
or U13263 (N_13263,N_12051,N_12497);
or U13264 (N_13264,N_12523,N_12138);
nand U13265 (N_13265,N_12103,N_12658);
or U13266 (N_13266,N_12215,N_12150);
and U13267 (N_13267,N_12736,N_12197);
or U13268 (N_13268,N_12042,N_12357);
xor U13269 (N_13269,N_12321,N_12244);
nand U13270 (N_13270,N_12080,N_12558);
or U13271 (N_13271,N_12536,N_12085);
and U13272 (N_13272,N_12244,N_12146);
nand U13273 (N_13273,N_12385,N_12017);
or U13274 (N_13274,N_12324,N_12604);
and U13275 (N_13275,N_12190,N_12110);
or U13276 (N_13276,N_12142,N_12314);
or U13277 (N_13277,N_12583,N_12575);
nor U13278 (N_13278,N_12223,N_12069);
or U13279 (N_13279,N_12251,N_12012);
xnor U13280 (N_13280,N_12485,N_12170);
nor U13281 (N_13281,N_12470,N_12690);
xor U13282 (N_13282,N_12504,N_12183);
or U13283 (N_13283,N_12387,N_12178);
nand U13284 (N_13284,N_12678,N_12247);
and U13285 (N_13285,N_12375,N_12352);
or U13286 (N_13286,N_12737,N_12051);
nand U13287 (N_13287,N_12269,N_12039);
or U13288 (N_13288,N_12745,N_12196);
or U13289 (N_13289,N_12372,N_12017);
nor U13290 (N_13290,N_12364,N_12098);
nor U13291 (N_13291,N_12271,N_12458);
nand U13292 (N_13292,N_12743,N_12511);
or U13293 (N_13293,N_12253,N_12038);
xor U13294 (N_13294,N_12664,N_12451);
and U13295 (N_13295,N_12323,N_12468);
nor U13296 (N_13296,N_12462,N_12598);
nor U13297 (N_13297,N_12621,N_12326);
nor U13298 (N_13298,N_12466,N_12286);
xnor U13299 (N_13299,N_12278,N_12483);
or U13300 (N_13300,N_12644,N_12345);
nor U13301 (N_13301,N_12076,N_12115);
nor U13302 (N_13302,N_12062,N_12213);
nor U13303 (N_13303,N_12549,N_12276);
xor U13304 (N_13304,N_12589,N_12635);
nor U13305 (N_13305,N_12699,N_12362);
nand U13306 (N_13306,N_12339,N_12173);
nor U13307 (N_13307,N_12266,N_12551);
xor U13308 (N_13308,N_12492,N_12137);
xnor U13309 (N_13309,N_12691,N_12388);
nor U13310 (N_13310,N_12494,N_12519);
nor U13311 (N_13311,N_12473,N_12583);
nor U13312 (N_13312,N_12031,N_12574);
nor U13313 (N_13313,N_12311,N_12634);
or U13314 (N_13314,N_12367,N_12725);
xnor U13315 (N_13315,N_12250,N_12448);
nor U13316 (N_13316,N_12030,N_12559);
and U13317 (N_13317,N_12622,N_12514);
nand U13318 (N_13318,N_12043,N_12689);
and U13319 (N_13319,N_12699,N_12118);
and U13320 (N_13320,N_12702,N_12131);
and U13321 (N_13321,N_12096,N_12313);
nand U13322 (N_13322,N_12207,N_12472);
and U13323 (N_13323,N_12152,N_12743);
nor U13324 (N_13324,N_12499,N_12733);
and U13325 (N_13325,N_12305,N_12654);
nand U13326 (N_13326,N_12369,N_12618);
and U13327 (N_13327,N_12336,N_12483);
nand U13328 (N_13328,N_12134,N_12504);
and U13329 (N_13329,N_12402,N_12504);
and U13330 (N_13330,N_12415,N_12061);
xnor U13331 (N_13331,N_12326,N_12092);
nand U13332 (N_13332,N_12617,N_12623);
or U13333 (N_13333,N_12342,N_12000);
or U13334 (N_13334,N_12318,N_12305);
nor U13335 (N_13335,N_12594,N_12495);
nand U13336 (N_13336,N_12002,N_12235);
nand U13337 (N_13337,N_12734,N_12005);
xnor U13338 (N_13338,N_12193,N_12585);
nand U13339 (N_13339,N_12054,N_12153);
or U13340 (N_13340,N_12012,N_12491);
nor U13341 (N_13341,N_12342,N_12583);
and U13342 (N_13342,N_12309,N_12481);
or U13343 (N_13343,N_12434,N_12737);
nand U13344 (N_13344,N_12476,N_12376);
xor U13345 (N_13345,N_12247,N_12260);
and U13346 (N_13346,N_12060,N_12669);
and U13347 (N_13347,N_12721,N_12249);
and U13348 (N_13348,N_12628,N_12021);
nor U13349 (N_13349,N_12298,N_12735);
nor U13350 (N_13350,N_12213,N_12084);
and U13351 (N_13351,N_12016,N_12158);
and U13352 (N_13352,N_12731,N_12725);
or U13353 (N_13353,N_12693,N_12571);
nor U13354 (N_13354,N_12250,N_12662);
or U13355 (N_13355,N_12443,N_12676);
xnor U13356 (N_13356,N_12596,N_12515);
nand U13357 (N_13357,N_12598,N_12681);
or U13358 (N_13358,N_12013,N_12002);
or U13359 (N_13359,N_12536,N_12592);
and U13360 (N_13360,N_12335,N_12727);
nor U13361 (N_13361,N_12673,N_12153);
or U13362 (N_13362,N_12092,N_12073);
xor U13363 (N_13363,N_12350,N_12205);
nand U13364 (N_13364,N_12614,N_12029);
xor U13365 (N_13365,N_12489,N_12124);
xor U13366 (N_13366,N_12579,N_12513);
nand U13367 (N_13367,N_12741,N_12606);
nor U13368 (N_13368,N_12305,N_12179);
and U13369 (N_13369,N_12511,N_12518);
nor U13370 (N_13370,N_12311,N_12329);
xnor U13371 (N_13371,N_12448,N_12249);
nand U13372 (N_13372,N_12067,N_12135);
or U13373 (N_13373,N_12279,N_12096);
nor U13374 (N_13374,N_12204,N_12446);
or U13375 (N_13375,N_12428,N_12524);
nor U13376 (N_13376,N_12604,N_12354);
nand U13377 (N_13377,N_12625,N_12743);
or U13378 (N_13378,N_12009,N_12028);
nand U13379 (N_13379,N_12713,N_12520);
nor U13380 (N_13380,N_12366,N_12394);
nor U13381 (N_13381,N_12198,N_12558);
or U13382 (N_13382,N_12598,N_12112);
nand U13383 (N_13383,N_12292,N_12223);
xnor U13384 (N_13384,N_12485,N_12465);
nor U13385 (N_13385,N_12155,N_12506);
and U13386 (N_13386,N_12519,N_12603);
nand U13387 (N_13387,N_12414,N_12481);
xor U13388 (N_13388,N_12222,N_12073);
or U13389 (N_13389,N_12729,N_12524);
or U13390 (N_13390,N_12470,N_12580);
or U13391 (N_13391,N_12536,N_12390);
and U13392 (N_13392,N_12213,N_12024);
nand U13393 (N_13393,N_12501,N_12225);
or U13394 (N_13394,N_12449,N_12123);
nand U13395 (N_13395,N_12108,N_12561);
or U13396 (N_13396,N_12174,N_12152);
nand U13397 (N_13397,N_12067,N_12463);
or U13398 (N_13398,N_12061,N_12631);
or U13399 (N_13399,N_12430,N_12493);
nor U13400 (N_13400,N_12389,N_12680);
nand U13401 (N_13401,N_12363,N_12017);
nor U13402 (N_13402,N_12317,N_12227);
nand U13403 (N_13403,N_12061,N_12207);
and U13404 (N_13404,N_12551,N_12425);
or U13405 (N_13405,N_12556,N_12496);
or U13406 (N_13406,N_12148,N_12195);
xor U13407 (N_13407,N_12001,N_12398);
or U13408 (N_13408,N_12632,N_12212);
nand U13409 (N_13409,N_12715,N_12732);
nand U13410 (N_13410,N_12312,N_12521);
and U13411 (N_13411,N_12348,N_12544);
xnor U13412 (N_13412,N_12577,N_12669);
nor U13413 (N_13413,N_12287,N_12589);
or U13414 (N_13414,N_12079,N_12008);
xnor U13415 (N_13415,N_12696,N_12452);
nor U13416 (N_13416,N_12253,N_12443);
nor U13417 (N_13417,N_12619,N_12059);
nor U13418 (N_13418,N_12506,N_12440);
and U13419 (N_13419,N_12051,N_12685);
or U13420 (N_13420,N_12389,N_12227);
or U13421 (N_13421,N_12221,N_12642);
and U13422 (N_13422,N_12173,N_12385);
and U13423 (N_13423,N_12611,N_12243);
nor U13424 (N_13424,N_12002,N_12158);
nor U13425 (N_13425,N_12541,N_12259);
nor U13426 (N_13426,N_12297,N_12643);
and U13427 (N_13427,N_12373,N_12217);
xor U13428 (N_13428,N_12612,N_12703);
nor U13429 (N_13429,N_12078,N_12269);
or U13430 (N_13430,N_12358,N_12628);
and U13431 (N_13431,N_12662,N_12140);
nand U13432 (N_13432,N_12726,N_12040);
xor U13433 (N_13433,N_12336,N_12118);
xnor U13434 (N_13434,N_12350,N_12256);
and U13435 (N_13435,N_12608,N_12437);
or U13436 (N_13436,N_12404,N_12016);
nor U13437 (N_13437,N_12297,N_12230);
and U13438 (N_13438,N_12229,N_12022);
nand U13439 (N_13439,N_12245,N_12181);
nand U13440 (N_13440,N_12235,N_12074);
or U13441 (N_13441,N_12448,N_12435);
nor U13442 (N_13442,N_12230,N_12578);
nand U13443 (N_13443,N_12012,N_12061);
xnor U13444 (N_13444,N_12348,N_12369);
and U13445 (N_13445,N_12623,N_12043);
nand U13446 (N_13446,N_12589,N_12560);
nand U13447 (N_13447,N_12174,N_12676);
nor U13448 (N_13448,N_12574,N_12665);
nor U13449 (N_13449,N_12423,N_12399);
or U13450 (N_13450,N_12044,N_12695);
or U13451 (N_13451,N_12292,N_12468);
nor U13452 (N_13452,N_12119,N_12374);
and U13453 (N_13453,N_12663,N_12090);
or U13454 (N_13454,N_12195,N_12183);
nand U13455 (N_13455,N_12724,N_12394);
and U13456 (N_13456,N_12745,N_12088);
nor U13457 (N_13457,N_12086,N_12405);
or U13458 (N_13458,N_12062,N_12211);
and U13459 (N_13459,N_12218,N_12048);
xnor U13460 (N_13460,N_12370,N_12526);
and U13461 (N_13461,N_12135,N_12084);
and U13462 (N_13462,N_12538,N_12626);
and U13463 (N_13463,N_12557,N_12109);
nand U13464 (N_13464,N_12731,N_12574);
nand U13465 (N_13465,N_12074,N_12342);
nand U13466 (N_13466,N_12070,N_12193);
nand U13467 (N_13467,N_12586,N_12643);
nand U13468 (N_13468,N_12333,N_12019);
xnor U13469 (N_13469,N_12224,N_12441);
xnor U13470 (N_13470,N_12573,N_12658);
or U13471 (N_13471,N_12413,N_12434);
or U13472 (N_13472,N_12520,N_12690);
xnor U13473 (N_13473,N_12569,N_12238);
xor U13474 (N_13474,N_12014,N_12473);
nand U13475 (N_13475,N_12131,N_12672);
or U13476 (N_13476,N_12718,N_12469);
nor U13477 (N_13477,N_12127,N_12346);
or U13478 (N_13478,N_12215,N_12019);
nand U13479 (N_13479,N_12091,N_12474);
nor U13480 (N_13480,N_12207,N_12182);
nor U13481 (N_13481,N_12186,N_12354);
nand U13482 (N_13482,N_12728,N_12240);
or U13483 (N_13483,N_12366,N_12434);
and U13484 (N_13484,N_12728,N_12099);
or U13485 (N_13485,N_12228,N_12492);
nor U13486 (N_13486,N_12405,N_12572);
or U13487 (N_13487,N_12310,N_12029);
or U13488 (N_13488,N_12483,N_12475);
nor U13489 (N_13489,N_12516,N_12258);
xnor U13490 (N_13490,N_12607,N_12483);
nand U13491 (N_13491,N_12130,N_12227);
nor U13492 (N_13492,N_12160,N_12737);
xor U13493 (N_13493,N_12331,N_12579);
or U13494 (N_13494,N_12375,N_12662);
and U13495 (N_13495,N_12623,N_12292);
nor U13496 (N_13496,N_12336,N_12360);
nor U13497 (N_13497,N_12053,N_12427);
or U13498 (N_13498,N_12287,N_12117);
xnor U13499 (N_13499,N_12150,N_12482);
nor U13500 (N_13500,N_12917,N_13490);
or U13501 (N_13501,N_12805,N_13189);
nor U13502 (N_13502,N_12883,N_13188);
nor U13503 (N_13503,N_13328,N_13002);
nand U13504 (N_13504,N_13420,N_13007);
or U13505 (N_13505,N_12819,N_13322);
and U13506 (N_13506,N_13321,N_13346);
nor U13507 (N_13507,N_13125,N_13158);
and U13508 (N_13508,N_13449,N_12762);
and U13509 (N_13509,N_13411,N_13419);
and U13510 (N_13510,N_13394,N_13171);
nand U13511 (N_13511,N_12918,N_12873);
nand U13512 (N_13512,N_13210,N_12812);
and U13513 (N_13513,N_13454,N_12890);
or U13514 (N_13514,N_12941,N_13202);
and U13515 (N_13515,N_13478,N_13013);
nand U13516 (N_13516,N_12752,N_13426);
nor U13517 (N_13517,N_13495,N_13384);
xnor U13518 (N_13518,N_13003,N_13349);
or U13519 (N_13519,N_13156,N_12754);
nor U13520 (N_13520,N_12802,N_13076);
nor U13521 (N_13521,N_13198,N_12895);
xor U13522 (N_13522,N_12949,N_13011);
xor U13523 (N_13523,N_12875,N_13369);
or U13524 (N_13524,N_12986,N_13285);
or U13525 (N_13525,N_12830,N_13139);
or U13526 (N_13526,N_12982,N_12954);
and U13527 (N_13527,N_13123,N_13250);
nand U13528 (N_13528,N_13414,N_13018);
and U13529 (N_13529,N_12851,N_12758);
nor U13530 (N_13530,N_13450,N_13067);
xnor U13531 (N_13531,N_13364,N_13054);
or U13532 (N_13532,N_13209,N_13493);
nor U13533 (N_13533,N_12791,N_13084);
xor U13534 (N_13534,N_13023,N_13387);
nand U13535 (N_13535,N_12811,N_13088);
nor U13536 (N_13536,N_13017,N_12960);
nor U13537 (N_13537,N_12947,N_13208);
and U13538 (N_13538,N_13117,N_13243);
xnor U13539 (N_13539,N_13448,N_13264);
and U13540 (N_13540,N_12871,N_13473);
xnor U13541 (N_13541,N_12850,N_13082);
nand U13542 (N_13542,N_12985,N_13444);
or U13543 (N_13543,N_12767,N_13096);
nor U13544 (N_13544,N_13235,N_13383);
xnor U13545 (N_13545,N_12860,N_13291);
xor U13546 (N_13546,N_13300,N_12885);
nor U13547 (N_13547,N_13019,N_13487);
and U13548 (N_13548,N_13040,N_13029);
xor U13549 (N_13549,N_13386,N_12872);
xor U13550 (N_13550,N_13148,N_13233);
nor U13551 (N_13551,N_13406,N_12928);
xor U13552 (N_13552,N_12927,N_13429);
and U13553 (N_13553,N_13111,N_13275);
xnor U13554 (N_13554,N_13035,N_12820);
xnor U13555 (N_13555,N_12966,N_13348);
nor U13556 (N_13556,N_12901,N_13178);
xnor U13557 (N_13557,N_13432,N_12987);
nor U13558 (N_13558,N_12995,N_13359);
nand U13559 (N_13559,N_12929,N_13227);
nand U13560 (N_13560,N_13279,N_12996);
xnor U13561 (N_13561,N_12834,N_13200);
nor U13562 (N_13562,N_13492,N_13457);
nor U13563 (N_13563,N_13446,N_13480);
nor U13564 (N_13564,N_12897,N_13032);
xor U13565 (N_13565,N_12953,N_13497);
nor U13566 (N_13566,N_13132,N_13355);
and U13567 (N_13567,N_13004,N_12755);
nor U13568 (N_13568,N_13255,N_13037);
nor U13569 (N_13569,N_13216,N_13219);
nand U13570 (N_13570,N_12876,N_13046);
and U13571 (N_13571,N_12836,N_13162);
nand U13572 (N_13572,N_12951,N_13159);
and U13573 (N_13573,N_13458,N_13164);
nor U13574 (N_13574,N_13177,N_13295);
or U13575 (N_13575,N_13447,N_13230);
and U13576 (N_13576,N_13065,N_13267);
nand U13577 (N_13577,N_13324,N_13168);
xor U13578 (N_13578,N_13270,N_13001);
and U13579 (N_13579,N_13073,N_13083);
and U13580 (N_13580,N_12807,N_13127);
nor U13581 (N_13581,N_12790,N_13408);
nor U13582 (N_13582,N_12920,N_12843);
or U13583 (N_13583,N_13424,N_13000);
and U13584 (N_13584,N_13190,N_13247);
nor U13585 (N_13585,N_13144,N_13263);
nand U13586 (N_13586,N_13167,N_13421);
xor U13587 (N_13587,N_13160,N_13362);
and U13588 (N_13588,N_12892,N_13259);
and U13589 (N_13589,N_12773,N_13020);
nand U13590 (N_13590,N_13488,N_13476);
nand U13591 (N_13591,N_12798,N_13030);
nand U13592 (N_13592,N_12809,N_13385);
xor U13593 (N_13593,N_13302,N_13282);
or U13594 (N_13594,N_13410,N_12968);
xnor U13595 (N_13595,N_13107,N_13395);
xor U13596 (N_13596,N_13361,N_12974);
nand U13597 (N_13597,N_13460,N_13262);
nor U13598 (N_13598,N_12879,N_12869);
xor U13599 (N_13599,N_13311,N_12965);
and U13600 (N_13600,N_13005,N_13462);
nand U13601 (N_13601,N_12804,N_13120);
or U13602 (N_13602,N_13360,N_13331);
nor U13603 (N_13603,N_12759,N_13204);
xor U13604 (N_13604,N_12937,N_13133);
nor U13605 (N_13605,N_12852,N_12956);
and U13606 (N_13606,N_13240,N_12854);
nand U13607 (N_13607,N_12925,N_13248);
or U13608 (N_13608,N_12877,N_12972);
nor U13609 (N_13609,N_12775,N_13253);
or U13610 (N_13610,N_13119,N_13113);
nor U13611 (N_13611,N_13415,N_12772);
xor U13612 (N_13612,N_12905,N_12878);
or U13613 (N_13613,N_12943,N_12907);
and U13614 (N_13614,N_12914,N_13214);
or U13615 (N_13615,N_12915,N_13367);
or U13616 (N_13616,N_13106,N_13371);
nor U13617 (N_13617,N_13211,N_13363);
nand U13618 (N_13618,N_12825,N_13484);
or U13619 (N_13619,N_12784,N_13437);
and U13620 (N_13620,N_13206,N_13124);
xnor U13621 (N_13621,N_12765,N_12936);
nor U13622 (N_13622,N_13357,N_12962);
xnor U13623 (N_13623,N_13296,N_13193);
xor U13624 (N_13624,N_12823,N_12888);
or U13625 (N_13625,N_13336,N_13150);
xor U13626 (N_13626,N_13380,N_12955);
nand U13627 (N_13627,N_13191,N_12839);
xor U13628 (N_13628,N_12884,N_13466);
and U13629 (N_13629,N_12806,N_13379);
nor U13630 (N_13630,N_13276,N_13482);
or U13631 (N_13631,N_12957,N_13241);
nor U13632 (N_13632,N_13097,N_12969);
xor U13633 (N_13633,N_13486,N_12891);
or U13634 (N_13634,N_13468,N_13422);
or U13635 (N_13635,N_13128,N_13252);
xnor U13636 (N_13636,N_13427,N_13327);
and U13637 (N_13637,N_13354,N_13186);
xor U13638 (N_13638,N_12849,N_13055);
nand U13639 (N_13639,N_13161,N_13234);
nand U13640 (N_13640,N_13060,N_12776);
or U13641 (N_13641,N_13008,N_13172);
and U13642 (N_13642,N_13413,N_13477);
xor U13643 (N_13643,N_12756,N_13231);
and U13644 (N_13644,N_13079,N_13286);
nand U13645 (N_13645,N_13404,N_13314);
nor U13646 (N_13646,N_12924,N_12977);
or U13647 (N_13647,N_13333,N_13173);
xor U13648 (N_13648,N_13047,N_12835);
and U13649 (N_13649,N_13381,N_13089);
and U13650 (N_13650,N_12896,N_13130);
nor U13651 (N_13651,N_13087,N_13353);
and U13652 (N_13652,N_13335,N_12882);
and U13653 (N_13653,N_12894,N_13074);
and U13654 (N_13654,N_13292,N_12950);
nor U13655 (N_13655,N_13043,N_13179);
or U13656 (N_13656,N_13245,N_13045);
nand U13657 (N_13657,N_13229,N_12779);
nand U13658 (N_13658,N_13077,N_12994);
xnor U13659 (N_13659,N_12829,N_13288);
and U13660 (N_13660,N_13220,N_13049);
and U13661 (N_13661,N_13356,N_13474);
and U13662 (N_13662,N_13393,N_13499);
xor U13663 (N_13663,N_13236,N_13062);
and U13664 (N_13664,N_13303,N_13465);
nor U13665 (N_13665,N_13121,N_12970);
xor U13666 (N_13666,N_12801,N_12958);
nor U13667 (N_13667,N_13319,N_13086);
and U13668 (N_13668,N_12959,N_13069);
and U13669 (N_13669,N_12862,N_13213);
and U13670 (N_13670,N_13337,N_13489);
nor U13671 (N_13671,N_12868,N_12946);
and U13672 (N_13672,N_13304,N_13271);
nand U13673 (N_13673,N_12911,N_12919);
xnor U13674 (N_13674,N_13050,N_13373);
xor U13675 (N_13675,N_13131,N_13290);
and U13676 (N_13676,N_13116,N_13028);
nand U13677 (N_13677,N_13382,N_13042);
and U13678 (N_13678,N_12799,N_12991);
and U13679 (N_13679,N_12922,N_12980);
and U13680 (N_13680,N_13143,N_13434);
and U13681 (N_13681,N_13254,N_12886);
and U13682 (N_13682,N_13080,N_12766);
or U13683 (N_13683,N_12912,N_13195);
nor U13684 (N_13684,N_12909,N_12858);
or U13685 (N_13685,N_13332,N_13199);
xnor U13686 (N_13686,N_12913,N_12881);
or U13687 (N_13687,N_12926,N_12808);
or U13688 (N_13688,N_13114,N_12810);
or U13689 (N_13689,N_13329,N_13149);
and U13690 (N_13690,N_12944,N_13343);
or U13691 (N_13691,N_13194,N_13136);
or U13692 (N_13692,N_13368,N_13175);
nand U13693 (N_13693,N_13090,N_13212);
or U13694 (N_13694,N_13221,N_12783);
nor U13695 (N_13695,N_13251,N_13467);
and U13696 (N_13696,N_13433,N_13472);
nor U13697 (N_13697,N_12999,N_12846);
nand U13698 (N_13698,N_13025,N_13325);
xnor U13699 (N_13699,N_12861,N_12934);
xnor U13700 (N_13700,N_13099,N_13481);
nand U13701 (N_13701,N_13301,N_13059);
or U13702 (N_13702,N_13438,N_12992);
xor U13703 (N_13703,N_13284,N_12751);
nand U13704 (N_13704,N_13330,N_12948);
nor U13705 (N_13705,N_13061,N_13483);
nand U13706 (N_13706,N_13166,N_13475);
and U13707 (N_13707,N_12976,N_12796);
nor U13708 (N_13708,N_12874,N_12795);
xnor U13709 (N_13709,N_12786,N_12935);
and U13710 (N_13710,N_13052,N_13485);
xnor U13711 (N_13711,N_12853,N_13323);
and U13712 (N_13712,N_12813,N_13281);
nand U13713 (N_13713,N_13135,N_13027);
xor U13714 (N_13714,N_13237,N_13320);
xor U13715 (N_13715,N_13402,N_13459);
nand U13716 (N_13716,N_13104,N_13024);
nor U13717 (N_13717,N_13294,N_13310);
nand U13718 (N_13718,N_13154,N_13033);
nor U13719 (N_13719,N_13036,N_13224);
nand U13720 (N_13720,N_13126,N_13015);
nor U13721 (N_13721,N_13228,N_13155);
and U13722 (N_13722,N_13197,N_13277);
and U13723 (N_13723,N_13058,N_13108);
and U13724 (N_13724,N_13287,N_13479);
xnor U13725 (N_13725,N_13246,N_13471);
xor U13726 (N_13726,N_13496,N_13494);
nor U13727 (N_13727,N_12814,N_12822);
and U13728 (N_13728,N_13366,N_13351);
xor U13729 (N_13729,N_13105,N_13418);
xnor U13730 (N_13730,N_12978,N_12782);
or U13731 (N_13731,N_12781,N_12865);
or U13732 (N_13732,N_13268,N_13181);
or U13733 (N_13733,N_13498,N_13265);
or U13734 (N_13734,N_13109,N_13280);
xor U13735 (N_13735,N_12979,N_13442);
xnor U13736 (N_13736,N_13044,N_12866);
or U13737 (N_13737,N_12908,N_13377);
nor U13738 (N_13738,N_13317,N_13196);
or U13739 (N_13739,N_13112,N_12855);
nor U13740 (N_13740,N_12777,N_12940);
or U13741 (N_13741,N_12921,N_13416);
nand U13742 (N_13742,N_12983,N_13152);
nor U13743 (N_13743,N_12845,N_12867);
and U13744 (N_13744,N_12831,N_12989);
or U13745 (N_13745,N_12785,N_12837);
nand U13746 (N_13746,N_12880,N_13283);
nand U13747 (N_13747,N_13142,N_13370);
or U13748 (N_13748,N_13269,N_12963);
nor U13749 (N_13749,N_13340,N_13176);
nand U13750 (N_13750,N_13358,N_12828);
or U13751 (N_13751,N_12763,N_13375);
or U13752 (N_13752,N_12997,N_13012);
nor U13753 (N_13753,N_13163,N_12764);
or U13754 (N_13754,N_13428,N_13334);
nor U13755 (N_13755,N_13100,N_13103);
nand U13756 (N_13756,N_12961,N_12818);
xor U13757 (N_13757,N_13068,N_13316);
xor U13758 (N_13758,N_13309,N_13026);
nand U13759 (N_13759,N_13315,N_13345);
and U13760 (N_13760,N_13313,N_13260);
and U13761 (N_13761,N_13170,N_13129);
nand U13762 (N_13762,N_13439,N_13095);
or U13763 (N_13763,N_12863,N_12952);
xnor U13764 (N_13764,N_13222,N_13347);
xor U13765 (N_13765,N_12803,N_13409);
or U13766 (N_13766,N_12780,N_13091);
nand U13767 (N_13767,N_13218,N_13192);
xor U13768 (N_13768,N_13398,N_12988);
xor U13769 (N_13769,N_12760,N_13307);
xnor U13770 (N_13770,N_12939,N_12841);
xnor U13771 (N_13771,N_12889,N_13070);
nor U13772 (N_13772,N_13293,N_13242);
nor U13773 (N_13773,N_13102,N_13169);
or U13774 (N_13774,N_13157,N_13305);
xor U13775 (N_13775,N_13289,N_13342);
nor U13776 (N_13776,N_12840,N_13185);
xnor U13777 (N_13777,N_13217,N_13038);
xor U13778 (N_13778,N_13075,N_13451);
xor U13779 (N_13779,N_13187,N_13078);
or U13780 (N_13780,N_13461,N_13134);
nor U13781 (N_13781,N_13396,N_13016);
and U13782 (N_13782,N_13064,N_13041);
nor U13783 (N_13783,N_12899,N_12857);
nand U13784 (N_13784,N_13403,N_13205);
nor U13785 (N_13785,N_12910,N_13400);
nand U13786 (N_13786,N_13318,N_12826);
or U13787 (N_13787,N_12815,N_12893);
nor U13788 (N_13788,N_13344,N_13390);
nor U13789 (N_13789,N_12856,N_13464);
nand U13790 (N_13790,N_13298,N_13184);
nand U13791 (N_13791,N_13445,N_13223);
and U13792 (N_13792,N_12923,N_12898);
and U13793 (N_13793,N_13441,N_13174);
nand U13794 (N_13794,N_13145,N_13401);
nor U13795 (N_13795,N_13374,N_13238);
nand U13796 (N_13796,N_12778,N_13388);
and U13797 (N_13797,N_13147,N_12906);
nor U13798 (N_13798,N_12942,N_13048);
xnor U13799 (N_13799,N_13225,N_12793);
nor U13800 (N_13800,N_13417,N_12945);
nor U13801 (N_13801,N_13137,N_13093);
xor U13802 (N_13802,N_13338,N_13180);
or U13803 (N_13803,N_13081,N_13053);
or U13804 (N_13804,N_12832,N_13249);
nor U13805 (N_13805,N_12932,N_13405);
or U13806 (N_13806,N_13376,N_13165);
and U13807 (N_13807,N_13412,N_13455);
and U13808 (N_13808,N_13350,N_13141);
or U13809 (N_13809,N_13306,N_13244);
nor U13810 (N_13810,N_12904,N_13122);
nor U13811 (N_13811,N_12800,N_12887);
nand U13812 (N_13812,N_12930,N_13207);
or U13813 (N_13813,N_13389,N_12990);
nor U13814 (N_13814,N_13010,N_13491);
and U13815 (N_13815,N_13056,N_12792);
xnor U13816 (N_13816,N_13443,N_13031);
or U13817 (N_13817,N_13423,N_13341);
nand U13818 (N_13818,N_12827,N_13138);
or U13819 (N_13819,N_13092,N_13431);
or U13820 (N_13820,N_13006,N_13009);
or U13821 (N_13821,N_13470,N_13312);
nand U13822 (N_13822,N_12838,N_12964);
nor U13823 (N_13823,N_13182,N_13297);
and U13824 (N_13824,N_13261,N_13203);
or U13825 (N_13825,N_12750,N_13034);
and U13826 (N_13826,N_12971,N_13273);
nor U13827 (N_13827,N_12761,N_13021);
and U13828 (N_13828,N_13039,N_12753);
nor U13829 (N_13829,N_13022,N_13085);
xor U13830 (N_13830,N_12797,N_12984);
xor U13831 (N_13831,N_12770,N_13430);
nand U13832 (N_13832,N_13115,N_13146);
nand U13833 (N_13833,N_13391,N_12774);
and U13834 (N_13834,N_12848,N_12824);
nand U13835 (N_13835,N_12768,N_12870);
nand U13836 (N_13836,N_13239,N_13232);
nor U13837 (N_13837,N_12771,N_12847);
xnor U13838 (N_13838,N_13063,N_12981);
or U13839 (N_13839,N_13407,N_13425);
nor U13840 (N_13840,N_12842,N_12757);
nor U13841 (N_13841,N_12833,N_12788);
xnor U13842 (N_13842,N_13118,N_12903);
nor U13843 (N_13843,N_13014,N_13352);
and U13844 (N_13844,N_12769,N_13365);
nor U13845 (N_13845,N_13378,N_12817);
xnor U13846 (N_13846,N_13094,N_13256);
nand U13847 (N_13847,N_12916,N_12975);
nor U13848 (N_13848,N_13326,N_13278);
xnor U13849 (N_13849,N_13258,N_13456);
xor U13850 (N_13850,N_12993,N_13057);
xor U13851 (N_13851,N_13153,N_12789);
or U13852 (N_13852,N_13071,N_13215);
nor U13853 (N_13853,N_12844,N_12933);
nand U13854 (N_13854,N_13372,N_13299);
xor U13855 (N_13855,N_13469,N_13397);
nand U13856 (N_13856,N_13151,N_13440);
nand U13857 (N_13857,N_12931,N_12998);
or U13858 (N_13858,N_13257,N_13399);
xnor U13859 (N_13859,N_13266,N_13051);
xor U13860 (N_13860,N_13463,N_13308);
nand U13861 (N_13861,N_13436,N_13110);
or U13862 (N_13862,N_13453,N_13339);
xor U13863 (N_13863,N_12900,N_12794);
xor U13864 (N_13864,N_13274,N_13392);
nand U13865 (N_13865,N_13226,N_12821);
nand U13866 (N_13866,N_12816,N_13140);
xnor U13867 (N_13867,N_12787,N_12967);
xnor U13868 (N_13868,N_13452,N_13183);
nand U13869 (N_13869,N_13066,N_12859);
nor U13870 (N_13870,N_12864,N_13098);
nand U13871 (N_13871,N_13201,N_13072);
xnor U13872 (N_13872,N_13435,N_12938);
nor U13873 (N_13873,N_13272,N_12902);
or U13874 (N_13874,N_13101,N_12973);
nand U13875 (N_13875,N_13403,N_13215);
nand U13876 (N_13876,N_13356,N_12768);
nand U13877 (N_13877,N_13197,N_12834);
xor U13878 (N_13878,N_12824,N_13364);
nor U13879 (N_13879,N_13309,N_13017);
nor U13880 (N_13880,N_12934,N_13320);
xor U13881 (N_13881,N_13066,N_13202);
and U13882 (N_13882,N_12961,N_13223);
xor U13883 (N_13883,N_12987,N_13047);
xor U13884 (N_13884,N_13249,N_13489);
nor U13885 (N_13885,N_13457,N_13076);
and U13886 (N_13886,N_12792,N_13234);
nand U13887 (N_13887,N_13401,N_13238);
xnor U13888 (N_13888,N_12777,N_13456);
or U13889 (N_13889,N_13163,N_13074);
nand U13890 (N_13890,N_13376,N_13239);
nor U13891 (N_13891,N_12798,N_13098);
nand U13892 (N_13892,N_12839,N_13300);
and U13893 (N_13893,N_13349,N_13442);
xor U13894 (N_13894,N_13173,N_13492);
xnor U13895 (N_13895,N_13089,N_13005);
xor U13896 (N_13896,N_12794,N_13387);
xnor U13897 (N_13897,N_13209,N_12933);
nor U13898 (N_13898,N_13080,N_12950);
and U13899 (N_13899,N_13301,N_12974);
xnor U13900 (N_13900,N_13182,N_13315);
and U13901 (N_13901,N_13137,N_12790);
xor U13902 (N_13902,N_12992,N_13369);
and U13903 (N_13903,N_12960,N_12929);
nor U13904 (N_13904,N_12762,N_12789);
xor U13905 (N_13905,N_13413,N_13281);
and U13906 (N_13906,N_12828,N_13399);
or U13907 (N_13907,N_13436,N_12918);
nand U13908 (N_13908,N_13006,N_13286);
nand U13909 (N_13909,N_12798,N_13188);
nand U13910 (N_13910,N_13209,N_13266);
and U13911 (N_13911,N_13421,N_13040);
nor U13912 (N_13912,N_13140,N_13276);
xnor U13913 (N_13913,N_13234,N_12955);
nand U13914 (N_13914,N_13194,N_13455);
xor U13915 (N_13915,N_12770,N_12906);
nand U13916 (N_13916,N_13302,N_13127);
and U13917 (N_13917,N_13221,N_13449);
nor U13918 (N_13918,N_13021,N_12899);
nand U13919 (N_13919,N_13496,N_13347);
and U13920 (N_13920,N_13273,N_12772);
nand U13921 (N_13921,N_12976,N_13371);
or U13922 (N_13922,N_12988,N_12817);
nand U13923 (N_13923,N_13392,N_13424);
xor U13924 (N_13924,N_13195,N_13446);
or U13925 (N_13925,N_13362,N_13207);
nor U13926 (N_13926,N_13207,N_13068);
nor U13927 (N_13927,N_13418,N_12822);
xor U13928 (N_13928,N_13349,N_12750);
or U13929 (N_13929,N_12851,N_13149);
xor U13930 (N_13930,N_13472,N_13115);
nand U13931 (N_13931,N_13323,N_12888);
and U13932 (N_13932,N_13455,N_13393);
and U13933 (N_13933,N_13083,N_12797);
and U13934 (N_13934,N_13201,N_13209);
xnor U13935 (N_13935,N_13155,N_13216);
nand U13936 (N_13936,N_13473,N_13054);
nor U13937 (N_13937,N_12863,N_13042);
and U13938 (N_13938,N_13100,N_12943);
nor U13939 (N_13939,N_12875,N_12983);
nor U13940 (N_13940,N_12824,N_13090);
and U13941 (N_13941,N_13085,N_13343);
or U13942 (N_13942,N_12884,N_12985);
nor U13943 (N_13943,N_13315,N_13467);
nand U13944 (N_13944,N_13457,N_13400);
xor U13945 (N_13945,N_13102,N_13377);
nor U13946 (N_13946,N_13126,N_13419);
or U13947 (N_13947,N_12961,N_13278);
xnor U13948 (N_13948,N_13262,N_13385);
or U13949 (N_13949,N_13224,N_12812);
and U13950 (N_13950,N_12979,N_13211);
nor U13951 (N_13951,N_12760,N_13255);
nand U13952 (N_13952,N_12870,N_13183);
or U13953 (N_13953,N_12833,N_12932);
xnor U13954 (N_13954,N_13257,N_13111);
nand U13955 (N_13955,N_13236,N_13247);
nand U13956 (N_13956,N_13251,N_12772);
xor U13957 (N_13957,N_13246,N_13133);
xnor U13958 (N_13958,N_12808,N_12834);
nand U13959 (N_13959,N_12789,N_13452);
and U13960 (N_13960,N_13132,N_13258);
nand U13961 (N_13961,N_13480,N_13039);
nand U13962 (N_13962,N_12956,N_13419);
xor U13963 (N_13963,N_13331,N_13057);
xnor U13964 (N_13964,N_13225,N_12953);
nand U13965 (N_13965,N_13135,N_13275);
nand U13966 (N_13966,N_13085,N_13154);
xor U13967 (N_13967,N_12851,N_13338);
nand U13968 (N_13968,N_13168,N_13226);
nor U13969 (N_13969,N_13256,N_13422);
nor U13970 (N_13970,N_13112,N_13136);
and U13971 (N_13971,N_13282,N_13185);
and U13972 (N_13972,N_13311,N_13429);
and U13973 (N_13973,N_13175,N_13327);
or U13974 (N_13974,N_12846,N_13478);
nor U13975 (N_13975,N_12804,N_12965);
and U13976 (N_13976,N_13484,N_13318);
and U13977 (N_13977,N_13078,N_13105);
xnor U13978 (N_13978,N_12778,N_13409);
and U13979 (N_13979,N_13396,N_12869);
and U13980 (N_13980,N_12780,N_13463);
xor U13981 (N_13981,N_13164,N_13074);
or U13982 (N_13982,N_13163,N_13227);
nand U13983 (N_13983,N_13357,N_12775);
nand U13984 (N_13984,N_12893,N_13219);
xor U13985 (N_13985,N_12906,N_13031);
or U13986 (N_13986,N_13445,N_12859);
nor U13987 (N_13987,N_13250,N_12911);
nand U13988 (N_13988,N_13220,N_12755);
nand U13989 (N_13989,N_12926,N_13102);
and U13990 (N_13990,N_13089,N_12870);
or U13991 (N_13991,N_12837,N_12833);
nor U13992 (N_13992,N_13412,N_12992);
nand U13993 (N_13993,N_12818,N_12907);
and U13994 (N_13994,N_13069,N_12892);
and U13995 (N_13995,N_13444,N_13049);
xor U13996 (N_13996,N_13010,N_13101);
or U13997 (N_13997,N_13451,N_13328);
nand U13998 (N_13998,N_12885,N_12783);
or U13999 (N_13999,N_12847,N_13279);
and U14000 (N_14000,N_13257,N_13218);
or U14001 (N_14001,N_12784,N_12965);
and U14002 (N_14002,N_13113,N_13174);
and U14003 (N_14003,N_13051,N_13355);
and U14004 (N_14004,N_13294,N_12846);
xor U14005 (N_14005,N_13196,N_13490);
or U14006 (N_14006,N_13456,N_13066);
and U14007 (N_14007,N_12914,N_13365);
nand U14008 (N_14008,N_13382,N_12939);
nor U14009 (N_14009,N_13163,N_13146);
nor U14010 (N_14010,N_13447,N_12841);
or U14011 (N_14011,N_13265,N_12885);
xnor U14012 (N_14012,N_13272,N_13311);
xnor U14013 (N_14013,N_12996,N_13129);
or U14014 (N_14014,N_13369,N_13156);
xor U14015 (N_14015,N_13291,N_13092);
or U14016 (N_14016,N_13406,N_13456);
or U14017 (N_14017,N_12941,N_13283);
and U14018 (N_14018,N_13444,N_13200);
xor U14019 (N_14019,N_13261,N_12919);
nor U14020 (N_14020,N_13462,N_13014);
or U14021 (N_14021,N_12960,N_12799);
xor U14022 (N_14022,N_12974,N_13496);
nor U14023 (N_14023,N_13021,N_12931);
and U14024 (N_14024,N_12941,N_13194);
and U14025 (N_14025,N_12754,N_12841);
and U14026 (N_14026,N_12803,N_13466);
and U14027 (N_14027,N_13117,N_12769);
or U14028 (N_14028,N_13400,N_13233);
nor U14029 (N_14029,N_12937,N_12868);
or U14030 (N_14030,N_13345,N_13323);
nand U14031 (N_14031,N_12997,N_13214);
nand U14032 (N_14032,N_12910,N_13139);
nor U14033 (N_14033,N_12776,N_13095);
xor U14034 (N_14034,N_13189,N_13349);
xor U14035 (N_14035,N_13487,N_13168);
and U14036 (N_14036,N_13318,N_13069);
or U14037 (N_14037,N_13143,N_13138);
and U14038 (N_14038,N_12960,N_12993);
nand U14039 (N_14039,N_13306,N_13372);
or U14040 (N_14040,N_13321,N_13111);
nand U14041 (N_14041,N_13445,N_13262);
and U14042 (N_14042,N_13191,N_13282);
xnor U14043 (N_14043,N_12843,N_13359);
nor U14044 (N_14044,N_13389,N_12856);
nand U14045 (N_14045,N_13400,N_13466);
and U14046 (N_14046,N_12792,N_13307);
or U14047 (N_14047,N_13377,N_13276);
and U14048 (N_14048,N_12778,N_13297);
nand U14049 (N_14049,N_12870,N_13279);
xor U14050 (N_14050,N_13361,N_13457);
nor U14051 (N_14051,N_13428,N_13155);
or U14052 (N_14052,N_13249,N_13335);
and U14053 (N_14053,N_12977,N_13111);
nand U14054 (N_14054,N_13190,N_13270);
nand U14055 (N_14055,N_13168,N_13290);
or U14056 (N_14056,N_12873,N_13448);
nand U14057 (N_14057,N_13438,N_13262);
nor U14058 (N_14058,N_12821,N_12950);
nand U14059 (N_14059,N_12889,N_13025);
nand U14060 (N_14060,N_12913,N_12865);
nand U14061 (N_14061,N_12987,N_13336);
xnor U14062 (N_14062,N_12955,N_13053);
xor U14063 (N_14063,N_12808,N_13107);
or U14064 (N_14064,N_13167,N_12913);
nand U14065 (N_14065,N_12793,N_13459);
nand U14066 (N_14066,N_13439,N_12903);
or U14067 (N_14067,N_13243,N_13418);
nand U14068 (N_14068,N_13065,N_13103);
or U14069 (N_14069,N_13292,N_13450);
and U14070 (N_14070,N_12945,N_13384);
nor U14071 (N_14071,N_13112,N_13359);
nor U14072 (N_14072,N_13312,N_13194);
or U14073 (N_14073,N_12804,N_13050);
nand U14074 (N_14074,N_13006,N_12858);
nand U14075 (N_14075,N_13288,N_13244);
xor U14076 (N_14076,N_13125,N_13303);
or U14077 (N_14077,N_13116,N_13330);
xor U14078 (N_14078,N_13293,N_13433);
or U14079 (N_14079,N_13279,N_12850);
and U14080 (N_14080,N_13211,N_13344);
nand U14081 (N_14081,N_13418,N_13063);
nor U14082 (N_14082,N_13084,N_12926);
or U14083 (N_14083,N_12903,N_13288);
nor U14084 (N_14084,N_13400,N_13096);
and U14085 (N_14085,N_13160,N_13167);
nand U14086 (N_14086,N_12833,N_12978);
and U14087 (N_14087,N_13383,N_13429);
nand U14088 (N_14088,N_13239,N_12821);
xor U14089 (N_14089,N_12912,N_12926);
nand U14090 (N_14090,N_12907,N_12946);
xnor U14091 (N_14091,N_13475,N_13222);
nand U14092 (N_14092,N_13315,N_13346);
and U14093 (N_14093,N_13383,N_12834);
or U14094 (N_14094,N_13330,N_13438);
nand U14095 (N_14095,N_13298,N_13466);
and U14096 (N_14096,N_13116,N_12869);
nand U14097 (N_14097,N_13091,N_12788);
or U14098 (N_14098,N_12922,N_13197);
nand U14099 (N_14099,N_13280,N_12936);
or U14100 (N_14100,N_13388,N_13202);
or U14101 (N_14101,N_12960,N_12911);
and U14102 (N_14102,N_13176,N_13109);
nand U14103 (N_14103,N_12896,N_13115);
nor U14104 (N_14104,N_13206,N_12968);
xnor U14105 (N_14105,N_13136,N_13275);
nand U14106 (N_14106,N_13498,N_12751);
or U14107 (N_14107,N_13303,N_12893);
nand U14108 (N_14108,N_13306,N_13260);
xnor U14109 (N_14109,N_12945,N_13416);
or U14110 (N_14110,N_13321,N_12965);
nor U14111 (N_14111,N_13478,N_12826);
or U14112 (N_14112,N_13004,N_13042);
xor U14113 (N_14113,N_13142,N_12843);
nor U14114 (N_14114,N_13038,N_13229);
or U14115 (N_14115,N_12825,N_12832);
or U14116 (N_14116,N_12795,N_13330);
nand U14117 (N_14117,N_13170,N_12770);
xnor U14118 (N_14118,N_13431,N_13241);
or U14119 (N_14119,N_12811,N_12844);
nor U14120 (N_14120,N_12796,N_12927);
or U14121 (N_14121,N_12925,N_13166);
or U14122 (N_14122,N_12957,N_12765);
or U14123 (N_14123,N_13353,N_12758);
nand U14124 (N_14124,N_13116,N_13040);
and U14125 (N_14125,N_13396,N_13444);
nand U14126 (N_14126,N_12859,N_13312);
xor U14127 (N_14127,N_13102,N_13361);
nor U14128 (N_14128,N_12983,N_13161);
or U14129 (N_14129,N_13389,N_13423);
xnor U14130 (N_14130,N_12824,N_12805);
nand U14131 (N_14131,N_13340,N_12860);
and U14132 (N_14132,N_13374,N_13491);
nand U14133 (N_14133,N_12833,N_13282);
or U14134 (N_14134,N_13015,N_12788);
nor U14135 (N_14135,N_13482,N_13468);
nand U14136 (N_14136,N_13233,N_13323);
nor U14137 (N_14137,N_13279,N_12954);
or U14138 (N_14138,N_13394,N_12774);
nor U14139 (N_14139,N_13395,N_13454);
and U14140 (N_14140,N_13101,N_13019);
xor U14141 (N_14141,N_13238,N_13037);
xnor U14142 (N_14142,N_13135,N_13293);
xnor U14143 (N_14143,N_13383,N_13173);
nor U14144 (N_14144,N_13053,N_13432);
and U14145 (N_14145,N_13373,N_13388);
xor U14146 (N_14146,N_13000,N_13417);
nor U14147 (N_14147,N_13080,N_13491);
xor U14148 (N_14148,N_13218,N_13438);
nand U14149 (N_14149,N_13063,N_13048);
nand U14150 (N_14150,N_13431,N_13009);
nand U14151 (N_14151,N_13053,N_13028);
or U14152 (N_14152,N_12792,N_13462);
nand U14153 (N_14153,N_12991,N_13045);
nand U14154 (N_14154,N_12849,N_13244);
or U14155 (N_14155,N_12763,N_12887);
nand U14156 (N_14156,N_13408,N_13132);
nor U14157 (N_14157,N_13277,N_12925);
nand U14158 (N_14158,N_13092,N_13221);
or U14159 (N_14159,N_13206,N_13465);
xnor U14160 (N_14160,N_12782,N_12923);
nand U14161 (N_14161,N_13446,N_12909);
or U14162 (N_14162,N_12915,N_13334);
and U14163 (N_14163,N_12763,N_13317);
nand U14164 (N_14164,N_13232,N_13171);
xnor U14165 (N_14165,N_12913,N_13199);
nor U14166 (N_14166,N_13422,N_13478);
and U14167 (N_14167,N_13027,N_12833);
nor U14168 (N_14168,N_13311,N_13019);
nand U14169 (N_14169,N_12960,N_13284);
or U14170 (N_14170,N_13041,N_12770);
or U14171 (N_14171,N_13051,N_12755);
nor U14172 (N_14172,N_13082,N_13467);
or U14173 (N_14173,N_13005,N_13418);
or U14174 (N_14174,N_13181,N_12776);
nor U14175 (N_14175,N_13216,N_13300);
nor U14176 (N_14176,N_12972,N_12836);
or U14177 (N_14177,N_13403,N_12938);
xor U14178 (N_14178,N_13176,N_13134);
nand U14179 (N_14179,N_12873,N_13034);
xnor U14180 (N_14180,N_13418,N_13109);
or U14181 (N_14181,N_12795,N_12797);
nor U14182 (N_14182,N_13200,N_13001);
nor U14183 (N_14183,N_12912,N_12815);
nand U14184 (N_14184,N_13456,N_12953);
or U14185 (N_14185,N_13459,N_12810);
xor U14186 (N_14186,N_12886,N_12855);
and U14187 (N_14187,N_13375,N_13343);
nor U14188 (N_14188,N_12960,N_13208);
and U14189 (N_14189,N_13330,N_12774);
nand U14190 (N_14190,N_13215,N_13247);
or U14191 (N_14191,N_13099,N_12836);
xor U14192 (N_14192,N_13011,N_12852);
nor U14193 (N_14193,N_13089,N_12878);
xnor U14194 (N_14194,N_13281,N_13147);
and U14195 (N_14195,N_12911,N_13474);
or U14196 (N_14196,N_12842,N_13242);
or U14197 (N_14197,N_12947,N_13339);
nor U14198 (N_14198,N_13216,N_13318);
nor U14199 (N_14199,N_13193,N_13047);
nor U14200 (N_14200,N_13388,N_13410);
xnor U14201 (N_14201,N_12906,N_13201);
nor U14202 (N_14202,N_12985,N_12868);
or U14203 (N_14203,N_13137,N_13230);
nor U14204 (N_14204,N_13353,N_13449);
and U14205 (N_14205,N_13143,N_12960);
or U14206 (N_14206,N_13277,N_13255);
nand U14207 (N_14207,N_13143,N_13441);
nor U14208 (N_14208,N_12887,N_12915);
nand U14209 (N_14209,N_13269,N_12771);
or U14210 (N_14210,N_13327,N_13252);
nor U14211 (N_14211,N_12809,N_12799);
nor U14212 (N_14212,N_13030,N_13181);
or U14213 (N_14213,N_12767,N_13329);
or U14214 (N_14214,N_12849,N_13085);
and U14215 (N_14215,N_12910,N_13286);
or U14216 (N_14216,N_12873,N_13495);
and U14217 (N_14217,N_12930,N_13201);
or U14218 (N_14218,N_13302,N_13297);
xnor U14219 (N_14219,N_13044,N_13449);
and U14220 (N_14220,N_13071,N_13218);
and U14221 (N_14221,N_13473,N_13260);
or U14222 (N_14222,N_13164,N_12830);
nand U14223 (N_14223,N_12903,N_13232);
nand U14224 (N_14224,N_12796,N_13047);
nand U14225 (N_14225,N_12984,N_13471);
nor U14226 (N_14226,N_12788,N_12946);
nand U14227 (N_14227,N_12859,N_12753);
nor U14228 (N_14228,N_13021,N_13382);
xnor U14229 (N_14229,N_13429,N_12866);
nor U14230 (N_14230,N_12865,N_13465);
xnor U14231 (N_14231,N_13228,N_12951);
nor U14232 (N_14232,N_13063,N_12860);
nand U14233 (N_14233,N_13117,N_13167);
or U14234 (N_14234,N_13126,N_13280);
nor U14235 (N_14235,N_12917,N_12786);
and U14236 (N_14236,N_13033,N_13053);
nand U14237 (N_14237,N_13125,N_12970);
xor U14238 (N_14238,N_13268,N_13464);
nor U14239 (N_14239,N_12776,N_12879);
xnor U14240 (N_14240,N_13150,N_13010);
xor U14241 (N_14241,N_12808,N_13143);
or U14242 (N_14242,N_13088,N_13137);
nor U14243 (N_14243,N_13026,N_12918);
or U14244 (N_14244,N_12923,N_13203);
nand U14245 (N_14245,N_13068,N_12978);
xnor U14246 (N_14246,N_13000,N_13077);
nor U14247 (N_14247,N_13099,N_13394);
or U14248 (N_14248,N_12920,N_12884);
xor U14249 (N_14249,N_12912,N_13132);
nand U14250 (N_14250,N_14033,N_13756);
xnor U14251 (N_14251,N_13532,N_13767);
xor U14252 (N_14252,N_13685,N_14091);
xor U14253 (N_14253,N_14174,N_13638);
nand U14254 (N_14254,N_13958,N_13772);
and U14255 (N_14255,N_14079,N_13779);
or U14256 (N_14256,N_14189,N_13785);
or U14257 (N_14257,N_13909,N_13898);
xor U14258 (N_14258,N_13748,N_14213);
nand U14259 (N_14259,N_13633,N_13952);
xnor U14260 (N_14260,N_13590,N_13837);
nand U14261 (N_14261,N_13819,N_13910);
nand U14262 (N_14262,N_14111,N_13709);
nand U14263 (N_14263,N_13630,N_13761);
xor U14264 (N_14264,N_14199,N_14121);
and U14265 (N_14265,N_13877,N_13614);
or U14266 (N_14266,N_13525,N_14103);
xnor U14267 (N_14267,N_13871,N_13731);
nor U14268 (N_14268,N_13987,N_14133);
or U14269 (N_14269,N_13777,N_14045);
and U14270 (N_14270,N_14218,N_13607);
nor U14271 (N_14271,N_13560,N_13594);
and U14272 (N_14272,N_13990,N_13942);
and U14273 (N_14273,N_14011,N_14143);
and U14274 (N_14274,N_13855,N_13551);
or U14275 (N_14275,N_13743,N_13730);
and U14276 (N_14276,N_14118,N_13860);
nand U14277 (N_14277,N_13567,N_13854);
xor U14278 (N_14278,N_13823,N_14196);
nor U14279 (N_14279,N_13572,N_13596);
or U14280 (N_14280,N_14206,N_14041);
xor U14281 (N_14281,N_14137,N_14031);
xor U14282 (N_14282,N_13912,N_14006);
nor U14283 (N_14283,N_13720,N_14126);
nor U14284 (N_14284,N_14120,N_13891);
or U14285 (N_14285,N_13674,N_13639);
or U14286 (N_14286,N_13671,N_13934);
xor U14287 (N_14287,N_13832,N_13751);
xnor U14288 (N_14288,N_14049,N_13565);
xnor U14289 (N_14289,N_13695,N_13876);
xnor U14290 (N_14290,N_13689,N_13644);
or U14291 (N_14291,N_13686,N_13542);
xnor U14292 (N_14292,N_14233,N_13875);
nor U14293 (N_14293,N_13889,N_14239);
xor U14294 (N_14294,N_13702,N_13788);
xor U14295 (N_14295,N_13935,N_13996);
nor U14296 (N_14296,N_13979,N_14180);
xnor U14297 (N_14297,N_14135,N_13853);
xor U14298 (N_14298,N_13859,N_13961);
xnor U14299 (N_14299,N_14238,N_13562);
and U14300 (N_14300,N_14013,N_13694);
nand U14301 (N_14301,N_13947,N_13547);
nor U14302 (N_14302,N_13956,N_13985);
xor U14303 (N_14303,N_13563,N_14172);
and U14304 (N_14304,N_13717,N_13553);
xor U14305 (N_14305,N_14227,N_13827);
or U14306 (N_14306,N_13949,N_14155);
or U14307 (N_14307,N_14003,N_14146);
and U14308 (N_14308,N_13518,N_13628);
nand U14309 (N_14309,N_13724,N_13882);
and U14310 (N_14310,N_13839,N_13757);
and U14311 (N_14311,N_13573,N_13955);
xor U14312 (N_14312,N_14212,N_13597);
nand U14313 (N_14313,N_13581,N_13840);
or U14314 (N_14314,N_13535,N_13737);
xnor U14315 (N_14315,N_14223,N_14047);
nand U14316 (N_14316,N_14202,N_13600);
xor U14317 (N_14317,N_14030,N_14070);
xor U14318 (N_14318,N_13744,N_13576);
nor U14319 (N_14319,N_13999,N_13514);
xnor U14320 (N_14320,N_13625,N_14123);
xnor U14321 (N_14321,N_13733,N_13601);
nor U14322 (N_14322,N_13842,N_14221);
or U14323 (N_14323,N_13826,N_13822);
and U14324 (N_14324,N_14021,N_13673);
or U14325 (N_14325,N_13536,N_13880);
xor U14326 (N_14326,N_13663,N_13977);
nor U14327 (N_14327,N_13810,N_13747);
nor U14328 (N_14328,N_13599,N_14089);
or U14329 (N_14329,N_14098,N_13554);
or U14330 (N_14330,N_13791,N_13787);
nand U14331 (N_14331,N_13591,N_13899);
xor U14332 (N_14332,N_14102,N_14176);
or U14333 (N_14333,N_13893,N_13660);
nand U14334 (N_14334,N_13746,N_13589);
and U14335 (N_14335,N_14169,N_13523);
and U14336 (N_14336,N_13897,N_14141);
nand U14337 (N_14337,N_14245,N_13764);
and U14338 (N_14338,N_14036,N_14088);
nand U14339 (N_14339,N_14232,N_13522);
xor U14340 (N_14340,N_13784,N_13510);
nor U14341 (N_14341,N_14086,N_13790);
nand U14342 (N_14342,N_13915,N_13896);
or U14343 (N_14343,N_13983,N_13656);
xnor U14344 (N_14344,N_13571,N_13556);
nand U14345 (N_14345,N_14226,N_13549);
or U14346 (N_14346,N_14188,N_13637);
nor U14347 (N_14347,N_14010,N_13558);
and U14348 (N_14348,N_13690,N_13856);
or U14349 (N_14349,N_14139,N_14096);
xnor U14350 (N_14350,N_13593,N_13980);
nand U14351 (N_14351,N_13742,N_13619);
xor U14352 (N_14352,N_14234,N_14197);
xor U14353 (N_14353,N_14005,N_14129);
nor U14354 (N_14354,N_13718,N_13966);
nor U14355 (N_14355,N_14183,N_14148);
nor U14356 (N_14356,N_13621,N_13833);
nand U14357 (N_14357,N_13907,N_13616);
nand U14358 (N_14358,N_13753,N_13651);
nor U14359 (N_14359,N_14162,N_13817);
nand U14360 (N_14360,N_13995,N_14019);
and U14361 (N_14361,N_13602,N_13623);
xor U14362 (N_14362,N_13729,N_14055);
nor U14363 (N_14363,N_13612,N_13771);
and U14364 (N_14364,N_13526,N_14128);
nand U14365 (N_14365,N_13994,N_14043);
nand U14366 (N_14366,N_14109,N_13850);
nor U14367 (N_14367,N_13750,N_13849);
and U14368 (N_14368,N_13680,N_14246);
and U14369 (N_14369,N_13603,N_14032);
xnor U14370 (N_14370,N_14097,N_13789);
nand U14371 (N_14371,N_13792,N_13675);
or U14372 (N_14372,N_13886,N_13858);
xor U14373 (N_14373,N_13939,N_14009);
or U14374 (N_14374,N_13968,N_14152);
nor U14375 (N_14375,N_13645,N_13710);
nand U14376 (N_14376,N_13626,N_14066);
and U14377 (N_14377,N_14080,N_13726);
xnor U14378 (N_14378,N_13502,N_13631);
and U14379 (N_14379,N_13964,N_13963);
nand U14380 (N_14380,N_13798,N_14192);
and U14381 (N_14381,N_13517,N_13975);
nor U14382 (N_14382,N_14171,N_13725);
xnor U14383 (N_14383,N_14076,N_13682);
and U14384 (N_14384,N_13931,N_13512);
nor U14385 (N_14385,N_13766,N_13878);
xor U14386 (N_14386,N_13927,N_13500);
xnor U14387 (N_14387,N_14000,N_14058);
nor U14388 (N_14388,N_14149,N_13611);
nand U14389 (N_14389,N_14165,N_13869);
and U14390 (N_14390,N_13847,N_13938);
nor U14391 (N_14391,N_13874,N_14007);
xor U14392 (N_14392,N_13799,N_13759);
nand U14393 (N_14393,N_13943,N_14104);
or U14394 (N_14394,N_13803,N_13648);
or U14395 (N_14395,N_14170,N_13890);
xor U14396 (N_14396,N_13884,N_14074);
nor U14397 (N_14397,N_13986,N_13866);
xor U14398 (N_14398,N_13804,N_13653);
xnor U14399 (N_14399,N_13794,N_13780);
and U14400 (N_14400,N_13960,N_13701);
nor U14401 (N_14401,N_14068,N_13754);
nand U14402 (N_14402,N_13579,N_14131);
and U14403 (N_14403,N_13984,N_13919);
or U14404 (N_14404,N_13598,N_14193);
or U14405 (N_14405,N_13678,N_13501);
nand U14406 (N_14406,N_13914,N_14144);
and U14407 (N_14407,N_14237,N_13800);
or U14408 (N_14408,N_13545,N_13716);
and U14409 (N_14409,N_13530,N_14130);
and U14410 (N_14410,N_13993,N_14012);
xor U14411 (N_14411,N_13580,N_13655);
nand U14412 (N_14412,N_13700,N_14230);
nor U14413 (N_14413,N_13795,N_13652);
and U14414 (N_14414,N_14201,N_13793);
xor U14415 (N_14415,N_13971,N_14248);
nor U14416 (N_14416,N_13913,N_13981);
xnor U14417 (N_14417,N_14210,N_13760);
and U14418 (N_14418,N_13516,N_13905);
xor U14419 (N_14419,N_14116,N_13688);
and U14420 (N_14420,N_13527,N_13959);
xnor U14421 (N_14421,N_14084,N_13998);
or U14422 (N_14422,N_13940,N_13515);
and U14423 (N_14423,N_13969,N_14101);
and U14424 (N_14424,N_13973,N_13774);
nand U14425 (N_14425,N_14225,N_13879);
and U14426 (N_14426,N_13807,N_14090);
nand U14427 (N_14427,N_13805,N_14028);
nand U14428 (N_14428,N_14067,N_14026);
xor U14429 (N_14429,N_13824,N_14077);
or U14430 (N_14430,N_13687,N_14053);
xor U14431 (N_14431,N_14185,N_13944);
xor U14432 (N_14432,N_13865,N_13714);
or U14433 (N_14433,N_14048,N_13740);
xor U14434 (N_14434,N_14136,N_13509);
nand U14435 (N_14435,N_13647,N_14020);
nor U14436 (N_14436,N_14163,N_14182);
and U14437 (N_14437,N_14219,N_13752);
or U14438 (N_14438,N_14108,N_13848);
nand U14439 (N_14439,N_14211,N_13967);
and U14440 (N_14440,N_13870,N_14075);
or U14441 (N_14441,N_13769,N_13681);
and U14442 (N_14442,N_13544,N_14017);
and U14443 (N_14443,N_13816,N_13814);
nand U14444 (N_14444,N_14214,N_13950);
xnor U14445 (N_14445,N_14140,N_13670);
or U14446 (N_14446,N_14069,N_13765);
or U14447 (N_14447,N_13796,N_14008);
nor U14448 (N_14448,N_14145,N_14179);
xnor U14449 (N_14449,N_13504,N_14110);
nor U14450 (N_14450,N_13519,N_14099);
nor U14451 (N_14451,N_14094,N_13829);
or U14452 (N_14452,N_13550,N_13811);
nor U14453 (N_14453,N_13908,N_13851);
and U14454 (N_14454,N_14134,N_14177);
and U14455 (N_14455,N_13520,N_14241);
nor U14456 (N_14456,N_14087,N_13592);
nor U14457 (N_14457,N_13929,N_13845);
and U14458 (N_14458,N_13922,N_13778);
xnor U14459 (N_14459,N_13584,N_13941);
nand U14460 (N_14460,N_13933,N_14247);
xnor U14461 (N_14461,N_14004,N_13894);
and U14462 (N_14462,N_13763,N_14157);
nand U14463 (N_14463,N_13538,N_14235);
xor U14464 (N_14464,N_14095,N_13782);
xnor U14465 (N_14465,N_13768,N_14166);
and U14466 (N_14466,N_13574,N_14125);
and U14467 (N_14467,N_13951,N_13861);
and U14468 (N_14468,N_13948,N_14178);
nor U14469 (N_14469,N_14002,N_13773);
nor U14470 (N_14470,N_14127,N_13524);
nand U14471 (N_14471,N_14132,N_13921);
xnor U14472 (N_14472,N_13801,N_13587);
nor U14473 (N_14473,N_14203,N_13617);
nor U14474 (N_14474,N_13945,N_13974);
or U14475 (N_14475,N_14156,N_13821);
and U14476 (N_14476,N_13722,N_14040);
nand U14477 (N_14477,N_14092,N_13528);
xnor U14478 (N_14478,N_13745,N_13885);
nor U14479 (N_14479,N_13721,N_14142);
or U14480 (N_14480,N_13582,N_14054);
nor U14481 (N_14481,N_13762,N_13978);
nor U14482 (N_14482,N_14207,N_13988);
nand U14483 (N_14483,N_13906,N_13711);
and U14484 (N_14484,N_13781,N_13642);
and U14485 (N_14485,N_14052,N_14208);
nor U14486 (N_14486,N_14194,N_13691);
nor U14487 (N_14487,N_13786,N_14059);
nor U14488 (N_14488,N_13972,N_14113);
and U14489 (N_14489,N_13734,N_13540);
nor U14490 (N_14490,N_14027,N_14035);
nor U14491 (N_14491,N_13615,N_13595);
nor U14492 (N_14492,N_14039,N_13583);
xor U14493 (N_14493,N_14173,N_13708);
xor U14494 (N_14494,N_13770,N_13677);
nor U14495 (N_14495,N_14138,N_14082);
nand U14496 (N_14496,N_14217,N_14195);
nor U14497 (N_14497,N_13669,N_13911);
and U14498 (N_14498,N_13723,N_13962);
and U14499 (N_14499,N_14244,N_13925);
and U14500 (N_14500,N_13577,N_13738);
xnor U14501 (N_14501,N_14100,N_14243);
or U14502 (N_14502,N_14001,N_13624);
nor U14503 (N_14503,N_13739,N_13627);
or U14504 (N_14504,N_13668,N_13991);
or U14505 (N_14505,N_14114,N_13634);
and U14506 (N_14506,N_13570,N_14119);
nor U14507 (N_14507,N_13641,N_13883);
and U14508 (N_14508,N_13683,N_13836);
and U14509 (N_14509,N_13643,N_13835);
and U14510 (N_14510,N_14107,N_14023);
or U14511 (N_14511,N_13719,N_13658);
nor U14512 (N_14512,N_13640,N_13531);
or U14513 (N_14513,N_14224,N_13902);
nand U14514 (N_14514,N_14093,N_14072);
xor U14515 (N_14515,N_13815,N_13957);
and U14516 (N_14516,N_13635,N_14071);
and U14517 (N_14517,N_13568,N_14198);
nand U14518 (N_14518,N_13546,N_13818);
nand U14519 (N_14519,N_13809,N_14167);
nand U14520 (N_14520,N_13873,N_14062);
or U14521 (N_14521,N_13704,N_13503);
nand U14522 (N_14522,N_13928,N_14181);
nor U14523 (N_14523,N_14184,N_13564);
and U14524 (N_14524,N_13569,N_14034);
or U14525 (N_14525,N_13953,N_14222);
xnor U14526 (N_14526,N_13982,N_13895);
and U14527 (N_14527,N_13812,N_14249);
nand U14528 (N_14528,N_13749,N_13863);
xnor U14529 (N_14529,N_13852,N_13622);
and U14530 (N_14530,N_13548,N_14124);
nand U14531 (N_14531,N_13808,N_14050);
nand U14532 (N_14532,N_13976,N_13900);
nor U14533 (N_14533,N_14115,N_13696);
or U14534 (N_14534,N_13825,N_14014);
and U14535 (N_14535,N_14236,N_13664);
nand U14536 (N_14536,N_14190,N_14158);
and U14537 (N_14537,N_14122,N_14215);
or U14538 (N_14538,N_13783,N_13507);
xnor U14539 (N_14539,N_13679,N_13555);
or U14540 (N_14540,N_14229,N_13705);
nor U14541 (N_14541,N_14063,N_14105);
and U14542 (N_14542,N_13693,N_13989);
nor U14543 (N_14543,N_14161,N_13684);
nor U14544 (N_14544,N_13736,N_13698);
nand U14545 (N_14545,N_14164,N_13888);
and U14546 (N_14546,N_13666,N_14117);
nor U14547 (N_14547,N_13926,N_13903);
xnor U14548 (N_14548,N_14046,N_13857);
nor U14549 (N_14549,N_13844,N_13838);
nor U14550 (N_14550,N_13657,N_14240);
xor U14551 (N_14551,N_13965,N_13586);
nand U14552 (N_14552,N_14216,N_13608);
xnor U14553 (N_14553,N_14200,N_13830);
nand U14554 (N_14554,N_13513,N_14044);
or U14555 (N_14555,N_14083,N_13662);
xor U14556 (N_14556,N_13713,N_13699);
nor U14557 (N_14557,N_13775,N_13506);
or U14558 (N_14558,N_13937,N_13557);
or U14559 (N_14559,N_13609,N_14220);
xor U14560 (N_14560,N_14015,N_13881);
nor U14561 (N_14561,N_13665,N_13636);
and U14562 (N_14562,N_13735,N_13578);
nor U14563 (N_14563,N_14159,N_14056);
and U14564 (N_14564,N_14022,N_13846);
nand U14565 (N_14565,N_13867,N_13534);
or U14566 (N_14566,N_14153,N_14038);
xor U14567 (N_14567,N_13727,N_13997);
nor U14568 (N_14568,N_13521,N_14112);
nand U14569 (N_14569,N_13632,N_13920);
or U14570 (N_14570,N_13936,N_13758);
nand U14571 (N_14571,N_13672,N_14191);
and U14572 (N_14572,N_13806,N_14064);
or U14573 (N_14573,N_14106,N_14154);
xor U14574 (N_14574,N_14078,N_14205);
nor U14575 (N_14575,N_14147,N_13649);
or U14576 (N_14576,N_13585,N_14231);
or U14577 (N_14577,N_13946,N_13892);
and U14578 (N_14578,N_14016,N_14168);
nand U14579 (N_14579,N_14018,N_13605);
xor U14580 (N_14580,N_14187,N_13924);
or U14581 (N_14581,N_13755,N_13629);
nor U14582 (N_14582,N_13697,N_13831);
or U14583 (N_14583,N_13970,N_14025);
nor U14584 (N_14584,N_13529,N_13654);
xnor U14585 (N_14585,N_13776,N_13588);
or U14586 (N_14586,N_13604,N_14150);
and U14587 (N_14587,N_13820,N_13901);
and U14588 (N_14588,N_13992,N_13618);
or U14589 (N_14589,N_14186,N_13620);
xor U14590 (N_14590,N_13954,N_13741);
nor U14591 (N_14591,N_13508,N_13930);
xnor U14592 (N_14592,N_13887,N_14060);
nand U14593 (N_14593,N_14242,N_13843);
or U14594 (N_14594,N_13715,N_14042);
and U14595 (N_14595,N_13613,N_13692);
xor U14596 (N_14596,N_13537,N_14057);
nand U14597 (N_14597,N_13646,N_13712);
nor U14598 (N_14598,N_14204,N_14051);
xnor U14599 (N_14599,N_14061,N_13552);
nand U14600 (N_14600,N_13862,N_14228);
or U14601 (N_14601,N_13904,N_13533);
nand U14602 (N_14602,N_13868,N_13918);
nor U14603 (N_14603,N_14029,N_13661);
or U14604 (N_14604,N_13676,N_13703);
and U14605 (N_14605,N_13864,N_13667);
nand U14606 (N_14606,N_14175,N_14151);
nand U14607 (N_14607,N_13559,N_13543);
and U14608 (N_14608,N_14065,N_13841);
xor U14609 (N_14609,N_14037,N_13916);
or U14610 (N_14610,N_14085,N_13650);
and U14611 (N_14611,N_14209,N_13541);
xnor U14612 (N_14612,N_13932,N_13834);
or U14613 (N_14613,N_13797,N_13732);
xor U14614 (N_14614,N_14073,N_13728);
nand U14615 (N_14615,N_13566,N_13802);
nand U14616 (N_14616,N_14160,N_13659);
xor U14617 (N_14617,N_13575,N_13511);
or U14618 (N_14618,N_13872,N_14081);
xnor U14619 (N_14619,N_13828,N_13606);
and U14620 (N_14620,N_13706,N_13707);
and U14621 (N_14621,N_14024,N_13917);
nor U14622 (N_14622,N_13610,N_13923);
nand U14623 (N_14623,N_13813,N_13561);
and U14624 (N_14624,N_13505,N_13539);
nand U14625 (N_14625,N_13750,N_14190);
and U14626 (N_14626,N_14040,N_13891);
or U14627 (N_14627,N_13563,N_14118);
and U14628 (N_14628,N_13652,N_14209);
nor U14629 (N_14629,N_13904,N_13795);
nor U14630 (N_14630,N_13633,N_14111);
nor U14631 (N_14631,N_13987,N_13656);
or U14632 (N_14632,N_14134,N_14069);
nand U14633 (N_14633,N_13742,N_14168);
nor U14634 (N_14634,N_14075,N_13873);
or U14635 (N_14635,N_14243,N_13910);
xnor U14636 (N_14636,N_14100,N_14125);
and U14637 (N_14637,N_13884,N_13933);
and U14638 (N_14638,N_13655,N_13592);
nor U14639 (N_14639,N_13630,N_13940);
and U14640 (N_14640,N_13814,N_13870);
and U14641 (N_14641,N_13813,N_13942);
xnor U14642 (N_14642,N_14215,N_13674);
and U14643 (N_14643,N_13616,N_13583);
nand U14644 (N_14644,N_14196,N_13925);
xnor U14645 (N_14645,N_14128,N_13845);
or U14646 (N_14646,N_13661,N_13957);
or U14647 (N_14647,N_13822,N_14228);
nand U14648 (N_14648,N_14135,N_13870);
and U14649 (N_14649,N_13834,N_13551);
xor U14650 (N_14650,N_13891,N_13814);
nand U14651 (N_14651,N_14205,N_14226);
nand U14652 (N_14652,N_13734,N_14050);
nor U14653 (N_14653,N_13542,N_13828);
xnor U14654 (N_14654,N_13838,N_14200);
and U14655 (N_14655,N_13571,N_14161);
xor U14656 (N_14656,N_13703,N_14245);
nand U14657 (N_14657,N_13839,N_13913);
nand U14658 (N_14658,N_13909,N_14129);
and U14659 (N_14659,N_14060,N_13825);
nand U14660 (N_14660,N_13684,N_13688);
xnor U14661 (N_14661,N_14229,N_13976);
and U14662 (N_14662,N_13573,N_13834);
nand U14663 (N_14663,N_13666,N_14168);
nand U14664 (N_14664,N_14119,N_13544);
nand U14665 (N_14665,N_13682,N_13633);
and U14666 (N_14666,N_14225,N_13810);
and U14667 (N_14667,N_13976,N_14076);
or U14668 (N_14668,N_13711,N_13825);
or U14669 (N_14669,N_14209,N_14082);
xor U14670 (N_14670,N_14239,N_13703);
xnor U14671 (N_14671,N_13895,N_14157);
nand U14672 (N_14672,N_14099,N_14230);
and U14673 (N_14673,N_14241,N_14055);
or U14674 (N_14674,N_13567,N_13721);
xnor U14675 (N_14675,N_13719,N_13915);
nor U14676 (N_14676,N_13535,N_14037);
nor U14677 (N_14677,N_13560,N_13993);
nor U14678 (N_14678,N_13722,N_13929);
nor U14679 (N_14679,N_13653,N_14124);
nand U14680 (N_14680,N_14242,N_13551);
and U14681 (N_14681,N_13769,N_13508);
xor U14682 (N_14682,N_14249,N_13663);
nand U14683 (N_14683,N_13926,N_14032);
nand U14684 (N_14684,N_14112,N_13575);
and U14685 (N_14685,N_14213,N_13825);
nand U14686 (N_14686,N_13943,N_13603);
xor U14687 (N_14687,N_14235,N_13511);
nor U14688 (N_14688,N_13521,N_14071);
xor U14689 (N_14689,N_13787,N_14100);
nor U14690 (N_14690,N_13998,N_14236);
or U14691 (N_14691,N_13948,N_14014);
xor U14692 (N_14692,N_14132,N_13743);
or U14693 (N_14693,N_14169,N_14040);
xor U14694 (N_14694,N_14203,N_13548);
nor U14695 (N_14695,N_13530,N_14218);
and U14696 (N_14696,N_13835,N_13594);
nor U14697 (N_14697,N_13551,N_13791);
xor U14698 (N_14698,N_13822,N_13554);
nor U14699 (N_14699,N_13668,N_14003);
nor U14700 (N_14700,N_14199,N_14196);
and U14701 (N_14701,N_13935,N_14011);
and U14702 (N_14702,N_13698,N_13594);
nand U14703 (N_14703,N_14148,N_13691);
and U14704 (N_14704,N_13855,N_13784);
and U14705 (N_14705,N_13957,N_14089);
or U14706 (N_14706,N_14165,N_14161);
xnor U14707 (N_14707,N_13677,N_14069);
nand U14708 (N_14708,N_14060,N_14142);
nand U14709 (N_14709,N_13779,N_13763);
nor U14710 (N_14710,N_13896,N_13603);
nor U14711 (N_14711,N_14186,N_13852);
xor U14712 (N_14712,N_14209,N_14056);
xnor U14713 (N_14713,N_14020,N_14214);
or U14714 (N_14714,N_13719,N_13801);
nand U14715 (N_14715,N_13584,N_13505);
or U14716 (N_14716,N_13835,N_13632);
and U14717 (N_14717,N_13743,N_13571);
xnor U14718 (N_14718,N_13706,N_14224);
nand U14719 (N_14719,N_14125,N_13983);
xor U14720 (N_14720,N_14221,N_13722);
nand U14721 (N_14721,N_13766,N_14078);
nor U14722 (N_14722,N_14019,N_13752);
nand U14723 (N_14723,N_13711,N_14174);
or U14724 (N_14724,N_13542,N_13505);
xor U14725 (N_14725,N_13503,N_13605);
or U14726 (N_14726,N_14236,N_13654);
nand U14727 (N_14727,N_14123,N_13934);
nor U14728 (N_14728,N_13926,N_13907);
nand U14729 (N_14729,N_13600,N_13659);
nor U14730 (N_14730,N_14117,N_14067);
and U14731 (N_14731,N_14126,N_13859);
nand U14732 (N_14732,N_13741,N_14228);
and U14733 (N_14733,N_14232,N_13809);
xnor U14734 (N_14734,N_14002,N_14025);
and U14735 (N_14735,N_14066,N_13621);
and U14736 (N_14736,N_13835,N_13874);
and U14737 (N_14737,N_13939,N_14035);
nor U14738 (N_14738,N_13956,N_14077);
xnor U14739 (N_14739,N_14059,N_13895);
and U14740 (N_14740,N_13556,N_13897);
nand U14741 (N_14741,N_13597,N_14159);
nand U14742 (N_14742,N_14144,N_14219);
or U14743 (N_14743,N_13771,N_13879);
or U14744 (N_14744,N_14149,N_13541);
xor U14745 (N_14745,N_13957,N_13534);
nor U14746 (N_14746,N_14196,N_13911);
or U14747 (N_14747,N_14189,N_14033);
and U14748 (N_14748,N_13769,N_13863);
xnor U14749 (N_14749,N_13955,N_13565);
and U14750 (N_14750,N_14024,N_13895);
or U14751 (N_14751,N_13776,N_14185);
nand U14752 (N_14752,N_13746,N_13710);
or U14753 (N_14753,N_14078,N_13761);
nand U14754 (N_14754,N_13980,N_13671);
nor U14755 (N_14755,N_13506,N_14157);
nor U14756 (N_14756,N_13520,N_14203);
nand U14757 (N_14757,N_14152,N_13574);
and U14758 (N_14758,N_14040,N_13520);
or U14759 (N_14759,N_13600,N_13547);
nand U14760 (N_14760,N_13793,N_13995);
and U14761 (N_14761,N_13947,N_14201);
nor U14762 (N_14762,N_13572,N_13617);
nand U14763 (N_14763,N_14128,N_13790);
xnor U14764 (N_14764,N_14074,N_13503);
nor U14765 (N_14765,N_13930,N_14106);
nand U14766 (N_14766,N_14151,N_13826);
or U14767 (N_14767,N_13638,N_14139);
and U14768 (N_14768,N_13640,N_14187);
nand U14769 (N_14769,N_13567,N_13703);
nor U14770 (N_14770,N_13521,N_13526);
nand U14771 (N_14771,N_14104,N_14172);
xnor U14772 (N_14772,N_13855,N_13617);
nor U14773 (N_14773,N_13544,N_14079);
nand U14774 (N_14774,N_13573,N_13789);
xor U14775 (N_14775,N_13662,N_13854);
nor U14776 (N_14776,N_13814,N_13899);
and U14777 (N_14777,N_14224,N_13589);
xor U14778 (N_14778,N_14037,N_13738);
nand U14779 (N_14779,N_13837,N_13690);
nand U14780 (N_14780,N_13829,N_13951);
nand U14781 (N_14781,N_13676,N_13526);
or U14782 (N_14782,N_13670,N_14084);
nand U14783 (N_14783,N_13544,N_14183);
and U14784 (N_14784,N_13942,N_13830);
and U14785 (N_14785,N_14104,N_13589);
nor U14786 (N_14786,N_13917,N_14230);
nand U14787 (N_14787,N_14178,N_13552);
xor U14788 (N_14788,N_14235,N_13912);
or U14789 (N_14789,N_13503,N_13765);
and U14790 (N_14790,N_13954,N_13763);
xnor U14791 (N_14791,N_13689,N_13755);
or U14792 (N_14792,N_13734,N_13985);
or U14793 (N_14793,N_13534,N_13820);
and U14794 (N_14794,N_13887,N_13911);
xor U14795 (N_14795,N_13656,N_13911);
xnor U14796 (N_14796,N_13752,N_14079);
or U14797 (N_14797,N_14214,N_13793);
xnor U14798 (N_14798,N_13807,N_13915);
and U14799 (N_14799,N_13532,N_13724);
xor U14800 (N_14800,N_13858,N_13801);
nor U14801 (N_14801,N_14149,N_14118);
nand U14802 (N_14802,N_13899,N_14232);
xor U14803 (N_14803,N_14044,N_13934);
or U14804 (N_14804,N_13640,N_13767);
or U14805 (N_14805,N_13569,N_14220);
or U14806 (N_14806,N_13522,N_13708);
or U14807 (N_14807,N_14021,N_13930);
and U14808 (N_14808,N_14041,N_13507);
nor U14809 (N_14809,N_13885,N_13732);
nor U14810 (N_14810,N_14002,N_13908);
nand U14811 (N_14811,N_13928,N_14133);
nor U14812 (N_14812,N_14111,N_13553);
and U14813 (N_14813,N_13845,N_13541);
and U14814 (N_14814,N_14033,N_14066);
nand U14815 (N_14815,N_13961,N_14248);
xor U14816 (N_14816,N_13980,N_13930);
nand U14817 (N_14817,N_13652,N_14194);
nor U14818 (N_14818,N_13966,N_13978);
nor U14819 (N_14819,N_14099,N_13993);
or U14820 (N_14820,N_13801,N_14036);
xnor U14821 (N_14821,N_14091,N_14169);
or U14822 (N_14822,N_14199,N_13910);
nor U14823 (N_14823,N_13814,N_13988);
and U14824 (N_14824,N_14053,N_13793);
and U14825 (N_14825,N_13680,N_14139);
nand U14826 (N_14826,N_13771,N_14191);
nand U14827 (N_14827,N_13925,N_13659);
or U14828 (N_14828,N_14055,N_13968);
xor U14829 (N_14829,N_13863,N_13952);
xor U14830 (N_14830,N_13885,N_13541);
nor U14831 (N_14831,N_13970,N_13557);
nand U14832 (N_14832,N_14054,N_13538);
xor U14833 (N_14833,N_13912,N_14051);
nand U14834 (N_14834,N_14054,N_14048);
xnor U14835 (N_14835,N_13580,N_13578);
nand U14836 (N_14836,N_13769,N_13909);
or U14837 (N_14837,N_14124,N_13557);
or U14838 (N_14838,N_14040,N_13973);
or U14839 (N_14839,N_13995,N_14025);
or U14840 (N_14840,N_13996,N_14158);
and U14841 (N_14841,N_13830,N_14077);
nand U14842 (N_14842,N_13850,N_13655);
nand U14843 (N_14843,N_13560,N_13861);
nor U14844 (N_14844,N_14002,N_14017);
nor U14845 (N_14845,N_13775,N_13816);
and U14846 (N_14846,N_13847,N_14223);
nand U14847 (N_14847,N_14148,N_13685);
nand U14848 (N_14848,N_13912,N_13974);
nor U14849 (N_14849,N_13846,N_14115);
nor U14850 (N_14850,N_13930,N_13848);
and U14851 (N_14851,N_13825,N_14146);
xnor U14852 (N_14852,N_14139,N_13541);
nor U14853 (N_14853,N_13942,N_13628);
nand U14854 (N_14854,N_13520,N_13511);
or U14855 (N_14855,N_14223,N_13964);
xor U14856 (N_14856,N_14247,N_13501);
nor U14857 (N_14857,N_13944,N_13587);
or U14858 (N_14858,N_13998,N_14192);
nand U14859 (N_14859,N_13522,N_13641);
xor U14860 (N_14860,N_14029,N_13727);
nor U14861 (N_14861,N_13634,N_14017);
and U14862 (N_14862,N_13715,N_14121);
xnor U14863 (N_14863,N_13779,N_13950);
xnor U14864 (N_14864,N_13544,N_13841);
and U14865 (N_14865,N_13684,N_13726);
and U14866 (N_14866,N_14004,N_13722);
and U14867 (N_14867,N_13997,N_13528);
or U14868 (N_14868,N_14012,N_13669);
nor U14869 (N_14869,N_14095,N_14229);
xnor U14870 (N_14870,N_14153,N_14098);
nor U14871 (N_14871,N_13849,N_13966);
xor U14872 (N_14872,N_13772,N_13594);
or U14873 (N_14873,N_13685,N_14064);
nor U14874 (N_14874,N_13513,N_14123);
or U14875 (N_14875,N_14116,N_13639);
and U14876 (N_14876,N_14102,N_13806);
nand U14877 (N_14877,N_13965,N_13837);
xor U14878 (N_14878,N_13722,N_13902);
nor U14879 (N_14879,N_14218,N_14075);
nand U14880 (N_14880,N_14220,N_13604);
xor U14881 (N_14881,N_13799,N_13664);
nor U14882 (N_14882,N_13618,N_13503);
or U14883 (N_14883,N_13760,N_13561);
or U14884 (N_14884,N_13878,N_13644);
xor U14885 (N_14885,N_14059,N_13834);
nand U14886 (N_14886,N_13725,N_13595);
and U14887 (N_14887,N_13635,N_13883);
xnor U14888 (N_14888,N_14027,N_14132);
xnor U14889 (N_14889,N_13669,N_13620);
nand U14890 (N_14890,N_13721,N_14244);
and U14891 (N_14891,N_13991,N_13768);
nand U14892 (N_14892,N_14216,N_14015);
and U14893 (N_14893,N_14081,N_14220);
and U14894 (N_14894,N_14161,N_13960);
nand U14895 (N_14895,N_13797,N_13762);
or U14896 (N_14896,N_13678,N_14188);
nand U14897 (N_14897,N_13677,N_14233);
and U14898 (N_14898,N_13595,N_13788);
nor U14899 (N_14899,N_14017,N_14086);
nand U14900 (N_14900,N_14187,N_13976);
nor U14901 (N_14901,N_13602,N_13868);
or U14902 (N_14902,N_13687,N_14051);
xnor U14903 (N_14903,N_13971,N_13792);
nor U14904 (N_14904,N_13972,N_13584);
xor U14905 (N_14905,N_14123,N_14008);
xnor U14906 (N_14906,N_14119,N_13657);
or U14907 (N_14907,N_13816,N_13502);
nand U14908 (N_14908,N_13998,N_13733);
nand U14909 (N_14909,N_14070,N_14224);
nand U14910 (N_14910,N_13738,N_14039);
nor U14911 (N_14911,N_13783,N_13853);
nor U14912 (N_14912,N_13821,N_13979);
xor U14913 (N_14913,N_13625,N_14121);
or U14914 (N_14914,N_13754,N_13694);
and U14915 (N_14915,N_13868,N_13669);
or U14916 (N_14916,N_14140,N_13776);
xor U14917 (N_14917,N_14135,N_13921);
xnor U14918 (N_14918,N_13828,N_14061);
nor U14919 (N_14919,N_13855,N_13520);
nor U14920 (N_14920,N_13854,N_14121);
or U14921 (N_14921,N_13874,N_14128);
and U14922 (N_14922,N_13726,N_14053);
or U14923 (N_14923,N_14032,N_13811);
and U14924 (N_14924,N_13869,N_13507);
and U14925 (N_14925,N_14066,N_13515);
nand U14926 (N_14926,N_14129,N_13861);
nand U14927 (N_14927,N_13812,N_14231);
nand U14928 (N_14928,N_14174,N_13730);
nor U14929 (N_14929,N_13732,N_14038);
nand U14930 (N_14930,N_14096,N_13574);
nor U14931 (N_14931,N_14077,N_14098);
nor U14932 (N_14932,N_14042,N_14244);
and U14933 (N_14933,N_13589,N_13914);
nor U14934 (N_14934,N_14206,N_14226);
nor U14935 (N_14935,N_13997,N_13753);
nor U14936 (N_14936,N_14148,N_13895);
nand U14937 (N_14937,N_14126,N_13502);
and U14938 (N_14938,N_13621,N_14229);
or U14939 (N_14939,N_14181,N_13722);
xnor U14940 (N_14940,N_13895,N_13502);
nor U14941 (N_14941,N_13650,N_13563);
xnor U14942 (N_14942,N_13926,N_13816);
nor U14943 (N_14943,N_13920,N_13627);
nor U14944 (N_14944,N_13799,N_14131);
and U14945 (N_14945,N_13688,N_13735);
nor U14946 (N_14946,N_13712,N_14207);
xor U14947 (N_14947,N_13627,N_13563);
or U14948 (N_14948,N_13728,N_13851);
and U14949 (N_14949,N_14028,N_14136);
and U14950 (N_14950,N_14081,N_13591);
and U14951 (N_14951,N_13808,N_13896);
nor U14952 (N_14952,N_14175,N_13968);
or U14953 (N_14953,N_13646,N_14045);
xnor U14954 (N_14954,N_13989,N_13574);
xnor U14955 (N_14955,N_14082,N_13825);
xnor U14956 (N_14956,N_13552,N_13624);
xor U14957 (N_14957,N_13535,N_13850);
and U14958 (N_14958,N_14104,N_14165);
nor U14959 (N_14959,N_13516,N_14218);
or U14960 (N_14960,N_13765,N_13568);
and U14961 (N_14961,N_13915,N_13868);
xor U14962 (N_14962,N_13966,N_14220);
and U14963 (N_14963,N_13530,N_13744);
xor U14964 (N_14964,N_13815,N_14157);
or U14965 (N_14965,N_13797,N_14135);
or U14966 (N_14966,N_14003,N_13967);
and U14967 (N_14967,N_13848,N_13949);
and U14968 (N_14968,N_13817,N_13977);
xor U14969 (N_14969,N_13568,N_14218);
nor U14970 (N_14970,N_13523,N_13794);
nor U14971 (N_14971,N_13974,N_13695);
and U14972 (N_14972,N_14117,N_13676);
nor U14973 (N_14973,N_13894,N_13885);
nor U14974 (N_14974,N_13756,N_13698);
xnor U14975 (N_14975,N_13742,N_13877);
nor U14976 (N_14976,N_14122,N_14216);
xnor U14977 (N_14977,N_13972,N_13718);
nand U14978 (N_14978,N_13571,N_13860);
xor U14979 (N_14979,N_13648,N_13751);
and U14980 (N_14980,N_13846,N_13925);
xor U14981 (N_14981,N_13713,N_13915);
nand U14982 (N_14982,N_14133,N_13743);
nand U14983 (N_14983,N_13963,N_14156);
and U14984 (N_14984,N_14229,N_13985);
xnor U14985 (N_14985,N_13878,N_13645);
and U14986 (N_14986,N_13891,N_13637);
nor U14987 (N_14987,N_13650,N_13785);
nand U14988 (N_14988,N_14086,N_13598);
nand U14989 (N_14989,N_14113,N_13822);
nand U14990 (N_14990,N_13798,N_13668);
and U14991 (N_14991,N_13892,N_13921);
xor U14992 (N_14992,N_13989,N_14006);
nand U14993 (N_14993,N_14205,N_13998);
xor U14994 (N_14994,N_13686,N_14209);
nor U14995 (N_14995,N_13534,N_14152);
nor U14996 (N_14996,N_14212,N_13908);
xnor U14997 (N_14997,N_14225,N_13760);
nand U14998 (N_14998,N_13511,N_13997);
or U14999 (N_14999,N_13974,N_13970);
xnor UO_0 (O_0,N_14773,N_14612);
nor UO_1 (O_1,N_14529,N_14671);
nand UO_2 (O_2,N_14829,N_14833);
or UO_3 (O_3,N_14939,N_14902);
nand UO_4 (O_4,N_14465,N_14459);
xor UO_5 (O_5,N_14848,N_14272);
xnor UO_6 (O_6,N_14283,N_14581);
xnor UO_7 (O_7,N_14933,N_14942);
and UO_8 (O_8,N_14991,N_14444);
nand UO_9 (O_9,N_14541,N_14821);
nor UO_10 (O_10,N_14972,N_14785);
nor UO_11 (O_11,N_14971,N_14817);
nor UO_12 (O_12,N_14864,N_14679);
or UO_13 (O_13,N_14310,N_14928);
or UO_14 (O_14,N_14711,N_14961);
nor UO_15 (O_15,N_14973,N_14966);
and UO_16 (O_16,N_14604,N_14960);
and UO_17 (O_17,N_14693,N_14446);
xor UO_18 (O_18,N_14329,N_14262);
or UO_19 (O_19,N_14984,N_14415);
xor UO_20 (O_20,N_14507,N_14631);
nor UO_21 (O_21,N_14878,N_14270);
xnor UO_22 (O_22,N_14330,N_14558);
nor UO_23 (O_23,N_14816,N_14700);
xor UO_24 (O_24,N_14783,N_14768);
nand UO_25 (O_25,N_14323,N_14941);
nand UO_26 (O_26,N_14646,N_14855);
and UO_27 (O_27,N_14709,N_14514);
xor UO_28 (O_28,N_14487,N_14666);
nor UO_29 (O_29,N_14999,N_14730);
or UO_30 (O_30,N_14766,N_14563);
xnor UO_31 (O_31,N_14919,N_14986);
xnor UO_32 (O_32,N_14936,N_14732);
nor UO_33 (O_33,N_14901,N_14682);
xnor UO_34 (O_34,N_14253,N_14691);
and UO_35 (O_35,N_14806,N_14910);
nand UO_36 (O_36,N_14412,N_14705);
nor UO_37 (O_37,N_14364,N_14717);
nand UO_38 (O_38,N_14657,N_14772);
or UO_39 (O_39,N_14726,N_14894);
or UO_40 (O_40,N_14553,N_14954);
and UO_41 (O_41,N_14265,N_14719);
nor UO_42 (O_42,N_14782,N_14510);
nor UO_43 (O_43,N_14505,N_14692);
xor UO_44 (O_44,N_14712,N_14259);
or UO_45 (O_45,N_14675,N_14303);
nand UO_46 (O_46,N_14276,N_14595);
nor UO_47 (O_47,N_14439,N_14771);
and UO_48 (O_48,N_14967,N_14292);
or UO_49 (O_49,N_14322,N_14668);
or UO_50 (O_50,N_14615,N_14610);
xor UO_51 (O_51,N_14792,N_14476);
or UO_52 (O_52,N_14392,N_14387);
nor UO_53 (O_53,N_14373,N_14371);
and UO_54 (O_54,N_14931,N_14331);
nand UO_55 (O_55,N_14361,N_14602);
nor UO_56 (O_56,N_14587,N_14836);
nor UO_57 (O_57,N_14865,N_14420);
nor UO_58 (O_58,N_14713,N_14900);
or UO_59 (O_59,N_14632,N_14530);
xor UO_60 (O_60,N_14449,N_14293);
xor UO_61 (O_61,N_14979,N_14251);
nor UO_62 (O_62,N_14795,N_14473);
nand UO_63 (O_63,N_14739,N_14983);
nand UO_64 (O_64,N_14353,N_14749);
nor UO_65 (O_65,N_14474,N_14334);
xnor UO_66 (O_66,N_14649,N_14533);
xor UO_67 (O_67,N_14764,N_14452);
nor UO_68 (O_68,N_14513,N_14951);
and UO_69 (O_69,N_14790,N_14450);
xnor UO_70 (O_70,N_14884,N_14582);
and UO_71 (O_71,N_14667,N_14736);
and UO_72 (O_72,N_14808,N_14565);
and UO_73 (O_73,N_14499,N_14949);
nor UO_74 (O_74,N_14492,N_14307);
nor UO_75 (O_75,N_14815,N_14740);
or UO_76 (O_76,N_14888,N_14289);
xnor UO_77 (O_77,N_14926,N_14267);
nor UO_78 (O_78,N_14280,N_14396);
nor UO_79 (O_79,N_14803,N_14407);
and UO_80 (O_80,N_14770,N_14639);
or UO_81 (O_81,N_14515,N_14596);
nor UO_82 (O_82,N_14897,N_14557);
and UO_83 (O_83,N_14852,N_14351);
or UO_84 (O_84,N_14588,N_14978);
nor UO_85 (O_85,N_14321,N_14315);
and UO_86 (O_86,N_14925,N_14309);
xor UO_87 (O_87,N_14355,N_14851);
or UO_88 (O_88,N_14826,N_14932);
nor UO_89 (O_89,N_14887,N_14468);
nand UO_90 (O_90,N_14707,N_14867);
or UO_91 (O_91,N_14332,N_14532);
and UO_92 (O_92,N_14422,N_14686);
nand UO_93 (O_93,N_14934,N_14592);
nand UO_94 (O_94,N_14943,N_14847);
and UO_95 (O_95,N_14818,N_14989);
or UO_96 (O_96,N_14413,N_14414);
nand UO_97 (O_97,N_14947,N_14920);
nor UO_98 (O_98,N_14964,N_14893);
and UO_99 (O_99,N_14752,N_14969);
and UO_100 (O_100,N_14814,N_14437);
nand UO_101 (O_101,N_14433,N_14625);
and UO_102 (O_102,N_14337,N_14774);
nor UO_103 (O_103,N_14389,N_14343);
and UO_104 (O_104,N_14540,N_14520);
or UO_105 (O_105,N_14708,N_14475);
or UO_106 (O_106,N_14737,N_14620);
or UO_107 (O_107,N_14921,N_14952);
and UO_108 (O_108,N_14432,N_14621);
and UO_109 (O_109,N_14630,N_14570);
nand UO_110 (O_110,N_14524,N_14341);
xnor UO_111 (O_111,N_14376,N_14429);
and UO_112 (O_112,N_14489,N_14794);
and UO_113 (O_113,N_14383,N_14655);
nand UO_114 (O_114,N_14410,N_14418);
nor UO_115 (O_115,N_14738,N_14491);
nor UO_116 (O_116,N_14349,N_14256);
or UO_117 (O_117,N_14759,N_14569);
nor UO_118 (O_118,N_14605,N_14512);
nand UO_119 (O_119,N_14835,N_14348);
xnor UO_120 (O_120,N_14299,N_14430);
xnor UO_121 (O_121,N_14627,N_14980);
nand UO_122 (O_122,N_14252,N_14832);
nor UO_123 (O_123,N_14757,N_14416);
or UO_124 (O_124,N_14377,N_14350);
nor UO_125 (O_125,N_14454,N_14765);
or UO_126 (O_126,N_14386,N_14805);
nor UO_127 (O_127,N_14899,N_14279);
xnor UO_128 (O_128,N_14269,N_14344);
or UO_129 (O_129,N_14600,N_14777);
xnor UO_130 (O_130,N_14417,N_14918);
nor UO_131 (O_131,N_14365,N_14311);
xor UO_132 (O_132,N_14635,N_14354);
or UO_133 (O_133,N_14304,N_14945);
and UO_134 (O_134,N_14527,N_14545);
nand UO_135 (O_135,N_14501,N_14706);
nor UO_136 (O_136,N_14963,N_14895);
and UO_137 (O_137,N_14519,N_14950);
and UO_138 (O_138,N_14486,N_14380);
nand UO_139 (O_139,N_14985,N_14975);
and UO_140 (O_140,N_14695,N_14687);
or UO_141 (O_141,N_14727,N_14990);
xnor UO_142 (O_142,N_14746,N_14658);
or UO_143 (O_143,N_14697,N_14731);
and UO_144 (O_144,N_14296,N_14591);
and UO_145 (O_145,N_14456,N_14339);
and UO_146 (O_146,N_14916,N_14479);
nor UO_147 (O_147,N_14576,N_14511);
or UO_148 (O_148,N_14968,N_14466);
nand UO_149 (O_149,N_14809,N_14500);
xnor UO_150 (O_150,N_14544,N_14388);
nor UO_151 (O_151,N_14250,N_14677);
and UO_152 (O_152,N_14426,N_14898);
or UO_153 (O_153,N_14325,N_14915);
nand UO_154 (O_154,N_14403,N_14518);
and UO_155 (O_155,N_14523,N_14779);
nand UO_156 (O_156,N_14427,N_14538);
nand UO_157 (O_157,N_14642,N_14965);
or UO_158 (O_158,N_14996,N_14616);
xor UO_159 (O_159,N_14406,N_14791);
and UO_160 (O_160,N_14882,N_14617);
xnor UO_161 (O_161,N_14756,N_14769);
nand UO_162 (O_162,N_14277,N_14647);
or UO_163 (O_163,N_14539,N_14335);
nor UO_164 (O_164,N_14393,N_14556);
and UO_165 (O_165,N_14799,N_14257);
nor UO_166 (O_166,N_14470,N_14760);
or UO_167 (O_167,N_14743,N_14734);
or UO_168 (O_168,N_14411,N_14670);
nand UO_169 (O_169,N_14913,N_14674);
nor UO_170 (O_170,N_14842,N_14589);
nor UO_171 (O_171,N_14750,N_14955);
xor UO_172 (O_172,N_14861,N_14645);
nand UO_173 (O_173,N_14398,N_14911);
or UO_174 (O_174,N_14301,N_14694);
or UO_175 (O_175,N_14298,N_14754);
xnor UO_176 (O_176,N_14652,N_14496);
xor UO_177 (O_177,N_14880,N_14534);
xor UO_178 (O_178,N_14813,N_14624);
nand UO_179 (O_179,N_14485,N_14892);
xnor UO_180 (O_180,N_14300,N_14297);
or UO_181 (O_181,N_14260,N_14609);
and UO_182 (O_182,N_14890,N_14326);
xnor UO_183 (O_183,N_14728,N_14696);
or UO_184 (O_184,N_14397,N_14502);
nor UO_185 (O_185,N_14603,N_14720);
and UO_186 (O_186,N_14665,N_14472);
or UO_187 (O_187,N_14729,N_14970);
or UO_188 (O_188,N_14281,N_14976);
and UO_189 (O_189,N_14856,N_14987);
or UO_190 (O_190,N_14903,N_14614);
nand UO_191 (O_191,N_14648,N_14327);
nand UO_192 (O_192,N_14555,N_14447);
or UO_193 (O_193,N_14497,N_14319);
nand UO_194 (O_194,N_14521,N_14715);
and UO_195 (O_195,N_14981,N_14352);
nor UO_196 (O_196,N_14345,N_14455);
and UO_197 (O_197,N_14995,N_14744);
nand UO_198 (O_198,N_14366,N_14929);
xnor UO_199 (O_199,N_14993,N_14287);
nand UO_200 (O_200,N_14956,N_14636);
or UO_201 (O_201,N_14896,N_14481);
nor UO_202 (O_202,N_14678,N_14577);
nor UO_203 (O_203,N_14275,N_14404);
and UO_204 (O_204,N_14324,N_14716);
and UO_205 (O_205,N_14844,N_14810);
and UO_206 (O_206,N_14912,N_14755);
or UO_207 (O_207,N_14255,N_14401);
nor UO_208 (O_208,N_14661,N_14723);
or UO_209 (O_209,N_14745,N_14643);
or UO_210 (O_210,N_14721,N_14982);
xor UO_211 (O_211,N_14284,N_14761);
or UO_212 (O_212,N_14690,N_14710);
xnor UO_213 (O_213,N_14735,N_14681);
nand UO_214 (O_214,N_14578,N_14571);
or UO_215 (O_215,N_14504,N_14843);
or UO_216 (O_216,N_14562,N_14458);
nor UO_217 (O_217,N_14837,N_14546);
nand UO_218 (O_218,N_14789,N_14333);
nor UO_219 (O_219,N_14493,N_14654);
nand UO_220 (O_220,N_14342,N_14435);
or UO_221 (O_221,N_14302,N_14689);
nand UO_222 (O_222,N_14846,N_14263);
xnor UO_223 (O_223,N_14428,N_14905);
xnor UO_224 (O_224,N_14360,N_14379);
or UO_225 (O_225,N_14751,N_14870);
and UO_226 (O_226,N_14282,N_14637);
nor UO_227 (O_227,N_14628,N_14575);
or UO_228 (O_228,N_14463,N_14471);
nand UO_229 (O_229,N_14683,N_14974);
xnor UO_230 (O_230,N_14409,N_14688);
nor UO_231 (O_231,N_14672,N_14480);
or UO_232 (O_232,N_14825,N_14607);
nand UO_233 (O_233,N_14914,N_14308);
and UO_234 (O_234,N_14525,N_14619);
or UO_235 (O_235,N_14306,N_14526);
nor UO_236 (O_236,N_14633,N_14359);
xor UO_237 (O_237,N_14725,N_14889);
nor UO_238 (O_238,N_14522,N_14800);
and UO_239 (O_239,N_14629,N_14651);
nor UO_240 (O_240,N_14781,N_14288);
nor UO_241 (O_241,N_14370,N_14274);
nor UO_242 (O_242,N_14859,N_14391);
or UO_243 (O_243,N_14722,N_14585);
nand UO_244 (O_244,N_14820,N_14927);
xnor UO_245 (O_245,N_14357,N_14811);
xor UO_246 (O_246,N_14611,N_14849);
or UO_247 (O_247,N_14369,N_14994);
nand UO_248 (O_248,N_14622,N_14704);
nor UO_249 (O_249,N_14598,N_14924);
and UO_250 (O_250,N_14566,N_14508);
nand UO_251 (O_251,N_14663,N_14358);
nor UO_252 (O_252,N_14548,N_14802);
or UO_253 (O_253,N_14273,N_14347);
or UO_254 (O_254,N_14823,N_14660);
xor UO_255 (O_255,N_14367,N_14786);
nand UO_256 (O_256,N_14599,N_14830);
nand UO_257 (O_257,N_14448,N_14988);
nand UO_258 (O_258,N_14885,N_14375);
nor UO_259 (O_259,N_14638,N_14494);
nand UO_260 (O_260,N_14372,N_14464);
and UO_261 (O_261,N_14363,N_14285);
and UO_262 (O_262,N_14659,N_14962);
nor UO_263 (O_263,N_14869,N_14268);
nor UO_264 (O_264,N_14295,N_14586);
or UO_265 (O_265,N_14702,N_14977);
nand UO_266 (O_266,N_14685,N_14703);
xnor UO_267 (O_267,N_14669,N_14488);
xnor UO_268 (O_268,N_14550,N_14374);
nor UO_269 (O_269,N_14460,N_14634);
or UO_270 (O_270,N_14753,N_14423);
nor UO_271 (O_271,N_14320,N_14857);
xor UO_272 (O_272,N_14640,N_14839);
nor UO_273 (O_273,N_14838,N_14390);
and UO_274 (O_274,N_14436,N_14935);
and UO_275 (O_275,N_14841,N_14767);
nand UO_276 (O_276,N_14294,N_14469);
nand UO_277 (O_277,N_14948,N_14385);
nand UO_278 (O_278,N_14457,N_14741);
nand UO_279 (O_279,N_14664,N_14421);
or UO_280 (O_280,N_14998,N_14762);
and UO_281 (O_281,N_14442,N_14537);
xnor UO_282 (O_282,N_14875,N_14891);
xor UO_283 (O_283,N_14547,N_14572);
or UO_284 (O_284,N_14382,N_14840);
nand UO_285 (O_285,N_14424,N_14938);
nand UO_286 (O_286,N_14946,N_14866);
or UO_287 (O_287,N_14580,N_14483);
and UO_288 (O_288,N_14787,N_14551);
and UO_289 (O_289,N_14775,N_14431);
or UO_290 (O_290,N_14845,N_14482);
nor UO_291 (O_291,N_14763,N_14579);
and UO_292 (O_292,N_14503,N_14362);
nor UO_293 (O_293,N_14405,N_14819);
and UO_294 (O_294,N_14758,N_14827);
nand UO_295 (O_295,N_14788,N_14590);
and UO_296 (O_296,N_14266,N_14796);
or UO_297 (O_297,N_14286,N_14395);
xnor UO_298 (O_298,N_14542,N_14854);
xnor UO_299 (O_299,N_14778,N_14626);
nor UO_300 (O_300,N_14724,N_14871);
nand UO_301 (O_301,N_14478,N_14742);
nand UO_302 (O_302,N_14879,N_14904);
or UO_303 (O_303,N_14881,N_14644);
or UO_304 (O_304,N_14714,N_14718);
xor UO_305 (O_305,N_14313,N_14340);
nor UO_306 (O_306,N_14594,N_14261);
nor UO_307 (O_307,N_14831,N_14543);
or UO_308 (O_308,N_14937,N_14923);
or UO_309 (O_309,N_14680,N_14822);
nor UO_310 (O_310,N_14930,N_14812);
or UO_311 (O_311,N_14873,N_14906);
or UO_312 (O_312,N_14801,N_14653);
nor UO_313 (O_313,N_14394,N_14290);
nor UO_314 (O_314,N_14399,N_14328);
or UO_315 (O_315,N_14314,N_14917);
nand UO_316 (O_316,N_14909,N_14384);
and UO_317 (O_317,N_14860,N_14528);
nor UO_318 (O_318,N_14509,N_14400);
xnor UO_319 (O_319,N_14506,N_14408);
nand UO_320 (O_320,N_14959,N_14997);
and UO_321 (O_321,N_14908,N_14608);
xnor UO_322 (O_322,N_14958,N_14944);
and UO_323 (O_323,N_14793,N_14650);
nor UO_324 (O_324,N_14443,N_14593);
or UO_325 (O_325,N_14560,N_14776);
nand UO_326 (O_326,N_14874,N_14317);
xnor UO_327 (O_327,N_14484,N_14356);
nand UO_328 (O_328,N_14346,N_14467);
xor UO_329 (O_329,N_14853,N_14858);
and UO_330 (O_330,N_14872,N_14568);
xor UO_331 (O_331,N_14549,N_14583);
xnor UO_332 (O_332,N_14517,N_14378);
or UO_333 (O_333,N_14561,N_14922);
and UO_334 (O_334,N_14883,N_14953);
nor UO_335 (O_335,N_14797,N_14368);
xor UO_336 (O_336,N_14490,N_14747);
xnor UO_337 (O_337,N_14613,N_14601);
or UO_338 (O_338,N_14451,N_14559);
nor UO_339 (O_339,N_14957,N_14305);
and UO_340 (O_340,N_14438,N_14264);
nand UO_341 (O_341,N_14453,N_14673);
xor UO_342 (O_342,N_14584,N_14574);
or UO_343 (O_343,N_14641,N_14606);
nor UO_344 (O_344,N_14564,N_14662);
or UO_345 (O_345,N_14597,N_14618);
and UO_346 (O_346,N_14862,N_14824);
nand UO_347 (O_347,N_14495,N_14699);
or UO_348 (O_348,N_14441,N_14434);
and UO_349 (O_349,N_14798,N_14316);
and UO_350 (O_350,N_14462,N_14940);
and UO_351 (O_351,N_14278,N_14318);
or UO_352 (O_352,N_14291,N_14834);
or UO_353 (O_353,N_14254,N_14780);
and UO_354 (O_354,N_14850,N_14567);
nor UO_355 (O_355,N_14684,N_14907);
nor UO_356 (O_356,N_14402,N_14656);
nand UO_357 (O_357,N_14701,N_14461);
nor UO_358 (O_358,N_14573,N_14886);
xnor UO_359 (O_359,N_14552,N_14498);
and UO_360 (O_360,N_14535,N_14445);
nor UO_361 (O_361,N_14863,N_14536);
xnor UO_362 (O_362,N_14312,N_14271);
or UO_363 (O_363,N_14804,N_14992);
xnor UO_364 (O_364,N_14868,N_14516);
and UO_365 (O_365,N_14440,N_14748);
and UO_366 (O_366,N_14531,N_14877);
nor UO_367 (O_367,N_14258,N_14876);
or UO_368 (O_368,N_14419,N_14623);
and UO_369 (O_369,N_14554,N_14807);
and UO_370 (O_370,N_14784,N_14477);
xor UO_371 (O_371,N_14381,N_14828);
nand UO_372 (O_372,N_14338,N_14676);
nor UO_373 (O_373,N_14698,N_14425);
nand UO_374 (O_374,N_14733,N_14336);
or UO_375 (O_375,N_14660,N_14446);
or UO_376 (O_376,N_14484,N_14474);
or UO_377 (O_377,N_14494,N_14348);
and UO_378 (O_378,N_14891,N_14451);
and UO_379 (O_379,N_14820,N_14320);
and UO_380 (O_380,N_14955,N_14491);
nand UO_381 (O_381,N_14802,N_14833);
nor UO_382 (O_382,N_14845,N_14349);
nand UO_383 (O_383,N_14969,N_14409);
and UO_384 (O_384,N_14799,N_14910);
xor UO_385 (O_385,N_14606,N_14823);
and UO_386 (O_386,N_14854,N_14525);
nor UO_387 (O_387,N_14367,N_14561);
nand UO_388 (O_388,N_14975,N_14291);
nor UO_389 (O_389,N_14936,N_14596);
nand UO_390 (O_390,N_14929,N_14437);
or UO_391 (O_391,N_14793,N_14402);
nand UO_392 (O_392,N_14273,N_14734);
nor UO_393 (O_393,N_14730,N_14388);
nor UO_394 (O_394,N_14591,N_14726);
xor UO_395 (O_395,N_14742,N_14995);
nand UO_396 (O_396,N_14592,N_14520);
and UO_397 (O_397,N_14587,N_14289);
and UO_398 (O_398,N_14289,N_14406);
nor UO_399 (O_399,N_14694,N_14430);
nor UO_400 (O_400,N_14548,N_14978);
or UO_401 (O_401,N_14316,N_14685);
or UO_402 (O_402,N_14779,N_14862);
nor UO_403 (O_403,N_14380,N_14743);
nor UO_404 (O_404,N_14286,N_14723);
nand UO_405 (O_405,N_14586,N_14617);
and UO_406 (O_406,N_14535,N_14540);
xnor UO_407 (O_407,N_14984,N_14590);
nor UO_408 (O_408,N_14636,N_14591);
nor UO_409 (O_409,N_14732,N_14767);
or UO_410 (O_410,N_14758,N_14399);
or UO_411 (O_411,N_14308,N_14390);
or UO_412 (O_412,N_14346,N_14998);
nand UO_413 (O_413,N_14363,N_14438);
nor UO_414 (O_414,N_14363,N_14540);
or UO_415 (O_415,N_14887,N_14375);
and UO_416 (O_416,N_14489,N_14464);
nor UO_417 (O_417,N_14613,N_14527);
or UO_418 (O_418,N_14562,N_14724);
or UO_419 (O_419,N_14359,N_14328);
or UO_420 (O_420,N_14574,N_14571);
nor UO_421 (O_421,N_14720,N_14571);
or UO_422 (O_422,N_14944,N_14291);
and UO_423 (O_423,N_14525,N_14676);
nor UO_424 (O_424,N_14760,N_14766);
xor UO_425 (O_425,N_14626,N_14358);
and UO_426 (O_426,N_14863,N_14387);
nand UO_427 (O_427,N_14856,N_14883);
nand UO_428 (O_428,N_14366,N_14361);
nand UO_429 (O_429,N_14530,N_14996);
xnor UO_430 (O_430,N_14790,N_14499);
nor UO_431 (O_431,N_14305,N_14465);
nand UO_432 (O_432,N_14633,N_14546);
and UO_433 (O_433,N_14515,N_14532);
xnor UO_434 (O_434,N_14940,N_14875);
or UO_435 (O_435,N_14295,N_14625);
nor UO_436 (O_436,N_14806,N_14999);
and UO_437 (O_437,N_14473,N_14325);
and UO_438 (O_438,N_14694,N_14982);
or UO_439 (O_439,N_14493,N_14725);
nand UO_440 (O_440,N_14906,N_14795);
xor UO_441 (O_441,N_14788,N_14976);
and UO_442 (O_442,N_14804,N_14887);
or UO_443 (O_443,N_14364,N_14456);
and UO_444 (O_444,N_14872,N_14911);
nand UO_445 (O_445,N_14412,N_14458);
nor UO_446 (O_446,N_14498,N_14281);
xor UO_447 (O_447,N_14979,N_14764);
and UO_448 (O_448,N_14717,N_14963);
xnor UO_449 (O_449,N_14634,N_14532);
nand UO_450 (O_450,N_14417,N_14281);
and UO_451 (O_451,N_14717,N_14285);
nand UO_452 (O_452,N_14599,N_14492);
xnor UO_453 (O_453,N_14293,N_14413);
xor UO_454 (O_454,N_14331,N_14620);
nand UO_455 (O_455,N_14724,N_14710);
nor UO_456 (O_456,N_14297,N_14496);
and UO_457 (O_457,N_14323,N_14464);
or UO_458 (O_458,N_14442,N_14554);
and UO_459 (O_459,N_14334,N_14988);
xnor UO_460 (O_460,N_14901,N_14737);
nor UO_461 (O_461,N_14292,N_14772);
or UO_462 (O_462,N_14661,N_14863);
nand UO_463 (O_463,N_14412,N_14774);
or UO_464 (O_464,N_14407,N_14946);
or UO_465 (O_465,N_14572,N_14908);
nor UO_466 (O_466,N_14760,N_14678);
xnor UO_467 (O_467,N_14657,N_14411);
nor UO_468 (O_468,N_14303,N_14495);
nand UO_469 (O_469,N_14941,N_14707);
nand UO_470 (O_470,N_14574,N_14914);
nor UO_471 (O_471,N_14723,N_14741);
xor UO_472 (O_472,N_14719,N_14261);
xor UO_473 (O_473,N_14776,N_14288);
xnor UO_474 (O_474,N_14635,N_14891);
nand UO_475 (O_475,N_14985,N_14485);
nand UO_476 (O_476,N_14569,N_14978);
or UO_477 (O_477,N_14531,N_14747);
and UO_478 (O_478,N_14944,N_14662);
and UO_479 (O_479,N_14757,N_14696);
and UO_480 (O_480,N_14843,N_14294);
or UO_481 (O_481,N_14610,N_14668);
or UO_482 (O_482,N_14787,N_14533);
or UO_483 (O_483,N_14259,N_14705);
or UO_484 (O_484,N_14820,N_14475);
or UO_485 (O_485,N_14796,N_14341);
and UO_486 (O_486,N_14713,N_14867);
xnor UO_487 (O_487,N_14580,N_14776);
or UO_488 (O_488,N_14916,N_14325);
nand UO_489 (O_489,N_14501,N_14395);
xor UO_490 (O_490,N_14437,N_14734);
xnor UO_491 (O_491,N_14588,N_14884);
nand UO_492 (O_492,N_14790,N_14422);
nor UO_493 (O_493,N_14345,N_14284);
nand UO_494 (O_494,N_14437,N_14865);
nor UO_495 (O_495,N_14513,N_14743);
xor UO_496 (O_496,N_14608,N_14870);
nor UO_497 (O_497,N_14398,N_14656);
nand UO_498 (O_498,N_14549,N_14604);
nor UO_499 (O_499,N_14652,N_14697);
and UO_500 (O_500,N_14397,N_14972);
nand UO_501 (O_501,N_14392,N_14282);
nor UO_502 (O_502,N_14390,N_14367);
or UO_503 (O_503,N_14417,N_14815);
and UO_504 (O_504,N_14718,N_14256);
or UO_505 (O_505,N_14829,N_14626);
nor UO_506 (O_506,N_14721,N_14562);
xnor UO_507 (O_507,N_14340,N_14480);
nand UO_508 (O_508,N_14815,N_14286);
or UO_509 (O_509,N_14540,N_14682);
nand UO_510 (O_510,N_14310,N_14411);
and UO_511 (O_511,N_14733,N_14847);
nand UO_512 (O_512,N_14485,N_14582);
or UO_513 (O_513,N_14694,N_14346);
and UO_514 (O_514,N_14765,N_14434);
or UO_515 (O_515,N_14367,N_14925);
nor UO_516 (O_516,N_14873,N_14377);
or UO_517 (O_517,N_14907,N_14539);
and UO_518 (O_518,N_14601,N_14709);
and UO_519 (O_519,N_14928,N_14866);
or UO_520 (O_520,N_14269,N_14274);
nor UO_521 (O_521,N_14827,N_14582);
xor UO_522 (O_522,N_14597,N_14499);
xnor UO_523 (O_523,N_14369,N_14564);
and UO_524 (O_524,N_14699,N_14569);
xnor UO_525 (O_525,N_14467,N_14713);
or UO_526 (O_526,N_14957,N_14789);
nor UO_527 (O_527,N_14925,N_14664);
xor UO_528 (O_528,N_14701,N_14911);
nand UO_529 (O_529,N_14574,N_14484);
nand UO_530 (O_530,N_14599,N_14936);
and UO_531 (O_531,N_14839,N_14742);
and UO_532 (O_532,N_14354,N_14985);
nor UO_533 (O_533,N_14420,N_14281);
nor UO_534 (O_534,N_14730,N_14762);
or UO_535 (O_535,N_14883,N_14919);
and UO_536 (O_536,N_14667,N_14830);
and UO_537 (O_537,N_14836,N_14305);
and UO_538 (O_538,N_14653,N_14871);
nor UO_539 (O_539,N_14656,N_14361);
or UO_540 (O_540,N_14460,N_14786);
nor UO_541 (O_541,N_14823,N_14263);
xor UO_542 (O_542,N_14703,N_14318);
or UO_543 (O_543,N_14384,N_14410);
and UO_544 (O_544,N_14267,N_14473);
nor UO_545 (O_545,N_14310,N_14904);
and UO_546 (O_546,N_14953,N_14738);
or UO_547 (O_547,N_14349,N_14852);
or UO_548 (O_548,N_14924,N_14885);
or UO_549 (O_549,N_14283,N_14517);
and UO_550 (O_550,N_14828,N_14406);
xnor UO_551 (O_551,N_14921,N_14258);
nor UO_552 (O_552,N_14252,N_14286);
nand UO_553 (O_553,N_14573,N_14785);
nor UO_554 (O_554,N_14929,N_14592);
nand UO_555 (O_555,N_14743,N_14343);
or UO_556 (O_556,N_14941,N_14899);
xnor UO_557 (O_557,N_14761,N_14276);
and UO_558 (O_558,N_14592,N_14795);
or UO_559 (O_559,N_14935,N_14597);
or UO_560 (O_560,N_14826,N_14280);
or UO_561 (O_561,N_14367,N_14834);
nand UO_562 (O_562,N_14403,N_14365);
xnor UO_563 (O_563,N_14529,N_14794);
xor UO_564 (O_564,N_14296,N_14916);
and UO_565 (O_565,N_14358,N_14907);
nor UO_566 (O_566,N_14312,N_14632);
xor UO_567 (O_567,N_14567,N_14994);
and UO_568 (O_568,N_14568,N_14347);
xnor UO_569 (O_569,N_14316,N_14450);
xor UO_570 (O_570,N_14778,N_14946);
or UO_571 (O_571,N_14707,N_14617);
nor UO_572 (O_572,N_14611,N_14375);
or UO_573 (O_573,N_14800,N_14985);
xor UO_574 (O_574,N_14650,N_14797);
and UO_575 (O_575,N_14403,N_14692);
or UO_576 (O_576,N_14945,N_14407);
and UO_577 (O_577,N_14948,N_14968);
nor UO_578 (O_578,N_14448,N_14803);
nand UO_579 (O_579,N_14667,N_14915);
nor UO_580 (O_580,N_14823,N_14557);
or UO_581 (O_581,N_14831,N_14710);
and UO_582 (O_582,N_14803,N_14455);
xor UO_583 (O_583,N_14647,N_14952);
xor UO_584 (O_584,N_14346,N_14959);
nand UO_585 (O_585,N_14369,N_14296);
xnor UO_586 (O_586,N_14687,N_14899);
xor UO_587 (O_587,N_14449,N_14866);
and UO_588 (O_588,N_14408,N_14776);
nand UO_589 (O_589,N_14506,N_14480);
or UO_590 (O_590,N_14892,N_14281);
xor UO_591 (O_591,N_14365,N_14697);
and UO_592 (O_592,N_14404,N_14548);
xor UO_593 (O_593,N_14381,N_14343);
nand UO_594 (O_594,N_14346,N_14256);
and UO_595 (O_595,N_14757,N_14672);
or UO_596 (O_596,N_14563,N_14329);
nor UO_597 (O_597,N_14357,N_14695);
nand UO_598 (O_598,N_14574,N_14599);
nor UO_599 (O_599,N_14850,N_14566);
nand UO_600 (O_600,N_14389,N_14487);
nand UO_601 (O_601,N_14733,N_14942);
and UO_602 (O_602,N_14346,N_14517);
and UO_603 (O_603,N_14368,N_14512);
nor UO_604 (O_604,N_14379,N_14517);
or UO_605 (O_605,N_14845,N_14855);
or UO_606 (O_606,N_14444,N_14468);
nor UO_607 (O_607,N_14313,N_14640);
or UO_608 (O_608,N_14633,N_14757);
xnor UO_609 (O_609,N_14777,N_14279);
or UO_610 (O_610,N_14393,N_14622);
and UO_611 (O_611,N_14686,N_14314);
nor UO_612 (O_612,N_14500,N_14436);
nor UO_613 (O_613,N_14422,N_14943);
xor UO_614 (O_614,N_14909,N_14537);
and UO_615 (O_615,N_14990,N_14531);
nand UO_616 (O_616,N_14402,N_14685);
nor UO_617 (O_617,N_14679,N_14455);
xnor UO_618 (O_618,N_14580,N_14602);
xor UO_619 (O_619,N_14661,N_14623);
nor UO_620 (O_620,N_14300,N_14817);
and UO_621 (O_621,N_14403,N_14302);
and UO_622 (O_622,N_14346,N_14995);
or UO_623 (O_623,N_14773,N_14923);
nor UO_624 (O_624,N_14257,N_14287);
nor UO_625 (O_625,N_14982,N_14977);
xnor UO_626 (O_626,N_14438,N_14511);
xor UO_627 (O_627,N_14763,N_14660);
xnor UO_628 (O_628,N_14599,N_14481);
or UO_629 (O_629,N_14261,N_14574);
nand UO_630 (O_630,N_14788,N_14999);
nor UO_631 (O_631,N_14501,N_14298);
nor UO_632 (O_632,N_14284,N_14288);
and UO_633 (O_633,N_14591,N_14759);
xor UO_634 (O_634,N_14328,N_14454);
nand UO_635 (O_635,N_14590,N_14586);
xnor UO_636 (O_636,N_14629,N_14744);
xor UO_637 (O_637,N_14345,N_14867);
and UO_638 (O_638,N_14561,N_14822);
nand UO_639 (O_639,N_14852,N_14729);
or UO_640 (O_640,N_14343,N_14832);
nor UO_641 (O_641,N_14433,N_14582);
nor UO_642 (O_642,N_14940,N_14290);
and UO_643 (O_643,N_14411,N_14575);
xor UO_644 (O_644,N_14594,N_14821);
nor UO_645 (O_645,N_14757,N_14725);
nor UO_646 (O_646,N_14816,N_14976);
xor UO_647 (O_647,N_14494,N_14761);
or UO_648 (O_648,N_14421,N_14529);
or UO_649 (O_649,N_14415,N_14469);
and UO_650 (O_650,N_14755,N_14705);
or UO_651 (O_651,N_14452,N_14957);
or UO_652 (O_652,N_14751,N_14739);
or UO_653 (O_653,N_14279,N_14787);
or UO_654 (O_654,N_14703,N_14297);
nand UO_655 (O_655,N_14711,N_14708);
xor UO_656 (O_656,N_14367,N_14892);
and UO_657 (O_657,N_14551,N_14595);
xnor UO_658 (O_658,N_14535,N_14572);
nand UO_659 (O_659,N_14932,N_14978);
nand UO_660 (O_660,N_14796,N_14989);
or UO_661 (O_661,N_14440,N_14751);
nor UO_662 (O_662,N_14494,N_14499);
nor UO_663 (O_663,N_14507,N_14267);
and UO_664 (O_664,N_14497,N_14313);
nor UO_665 (O_665,N_14254,N_14690);
xor UO_666 (O_666,N_14434,N_14784);
nand UO_667 (O_667,N_14591,N_14357);
nor UO_668 (O_668,N_14373,N_14825);
nand UO_669 (O_669,N_14694,N_14296);
or UO_670 (O_670,N_14472,N_14251);
and UO_671 (O_671,N_14766,N_14623);
and UO_672 (O_672,N_14672,N_14403);
xnor UO_673 (O_673,N_14365,N_14615);
nand UO_674 (O_674,N_14656,N_14362);
nor UO_675 (O_675,N_14390,N_14769);
xor UO_676 (O_676,N_14722,N_14327);
nor UO_677 (O_677,N_14526,N_14904);
and UO_678 (O_678,N_14346,N_14723);
xnor UO_679 (O_679,N_14639,N_14285);
xnor UO_680 (O_680,N_14855,N_14449);
and UO_681 (O_681,N_14962,N_14468);
nor UO_682 (O_682,N_14661,N_14855);
nor UO_683 (O_683,N_14302,N_14536);
nand UO_684 (O_684,N_14318,N_14833);
nor UO_685 (O_685,N_14850,N_14951);
nor UO_686 (O_686,N_14300,N_14364);
nand UO_687 (O_687,N_14342,N_14329);
xnor UO_688 (O_688,N_14408,N_14422);
or UO_689 (O_689,N_14382,N_14377);
and UO_690 (O_690,N_14330,N_14881);
nor UO_691 (O_691,N_14510,N_14896);
xnor UO_692 (O_692,N_14407,N_14930);
or UO_693 (O_693,N_14956,N_14865);
nand UO_694 (O_694,N_14855,N_14821);
and UO_695 (O_695,N_14483,N_14914);
or UO_696 (O_696,N_14639,N_14563);
nand UO_697 (O_697,N_14620,N_14459);
xor UO_698 (O_698,N_14856,N_14269);
or UO_699 (O_699,N_14524,N_14639);
nand UO_700 (O_700,N_14611,N_14914);
nor UO_701 (O_701,N_14850,N_14450);
or UO_702 (O_702,N_14682,N_14761);
and UO_703 (O_703,N_14556,N_14552);
xnor UO_704 (O_704,N_14430,N_14815);
and UO_705 (O_705,N_14320,N_14527);
nor UO_706 (O_706,N_14976,N_14566);
nor UO_707 (O_707,N_14655,N_14687);
or UO_708 (O_708,N_14788,N_14665);
xnor UO_709 (O_709,N_14655,N_14883);
nand UO_710 (O_710,N_14306,N_14820);
nand UO_711 (O_711,N_14466,N_14520);
and UO_712 (O_712,N_14540,N_14765);
nor UO_713 (O_713,N_14472,N_14706);
or UO_714 (O_714,N_14657,N_14739);
and UO_715 (O_715,N_14859,N_14285);
xnor UO_716 (O_716,N_14792,N_14650);
or UO_717 (O_717,N_14764,N_14362);
xor UO_718 (O_718,N_14416,N_14408);
nand UO_719 (O_719,N_14982,N_14510);
xnor UO_720 (O_720,N_14317,N_14836);
nand UO_721 (O_721,N_14460,N_14550);
nor UO_722 (O_722,N_14426,N_14728);
nand UO_723 (O_723,N_14786,N_14761);
nand UO_724 (O_724,N_14723,N_14868);
or UO_725 (O_725,N_14408,N_14472);
nor UO_726 (O_726,N_14432,N_14329);
nor UO_727 (O_727,N_14347,N_14933);
nor UO_728 (O_728,N_14456,N_14657);
nor UO_729 (O_729,N_14837,N_14708);
nor UO_730 (O_730,N_14915,N_14572);
nor UO_731 (O_731,N_14503,N_14590);
nor UO_732 (O_732,N_14530,N_14442);
nand UO_733 (O_733,N_14448,N_14944);
nor UO_734 (O_734,N_14300,N_14472);
nor UO_735 (O_735,N_14255,N_14373);
and UO_736 (O_736,N_14811,N_14548);
and UO_737 (O_737,N_14808,N_14769);
or UO_738 (O_738,N_14269,N_14972);
and UO_739 (O_739,N_14490,N_14604);
and UO_740 (O_740,N_14603,N_14296);
and UO_741 (O_741,N_14473,N_14758);
nand UO_742 (O_742,N_14283,N_14320);
nor UO_743 (O_743,N_14615,N_14578);
xnor UO_744 (O_744,N_14570,N_14763);
and UO_745 (O_745,N_14763,N_14295);
or UO_746 (O_746,N_14560,N_14936);
nand UO_747 (O_747,N_14735,N_14483);
or UO_748 (O_748,N_14585,N_14824);
nand UO_749 (O_749,N_14702,N_14307);
and UO_750 (O_750,N_14587,N_14334);
nand UO_751 (O_751,N_14622,N_14392);
nor UO_752 (O_752,N_14805,N_14934);
and UO_753 (O_753,N_14645,N_14379);
nand UO_754 (O_754,N_14293,N_14378);
nand UO_755 (O_755,N_14356,N_14554);
nand UO_756 (O_756,N_14393,N_14903);
xnor UO_757 (O_757,N_14565,N_14791);
nor UO_758 (O_758,N_14256,N_14403);
or UO_759 (O_759,N_14306,N_14268);
and UO_760 (O_760,N_14352,N_14783);
or UO_761 (O_761,N_14959,N_14721);
xnor UO_762 (O_762,N_14435,N_14820);
xnor UO_763 (O_763,N_14657,N_14914);
xnor UO_764 (O_764,N_14650,N_14569);
and UO_765 (O_765,N_14293,N_14843);
nand UO_766 (O_766,N_14867,N_14856);
xor UO_767 (O_767,N_14921,N_14607);
nor UO_768 (O_768,N_14346,N_14971);
and UO_769 (O_769,N_14409,N_14748);
xnor UO_770 (O_770,N_14983,N_14911);
xor UO_771 (O_771,N_14467,N_14839);
or UO_772 (O_772,N_14819,N_14739);
nand UO_773 (O_773,N_14873,N_14539);
or UO_774 (O_774,N_14587,N_14367);
nand UO_775 (O_775,N_14979,N_14717);
nand UO_776 (O_776,N_14924,N_14477);
nand UO_777 (O_777,N_14768,N_14700);
and UO_778 (O_778,N_14452,N_14457);
and UO_779 (O_779,N_14861,N_14867);
and UO_780 (O_780,N_14886,N_14695);
and UO_781 (O_781,N_14876,N_14415);
xor UO_782 (O_782,N_14835,N_14616);
or UO_783 (O_783,N_14250,N_14681);
xor UO_784 (O_784,N_14485,N_14942);
or UO_785 (O_785,N_14768,N_14877);
nor UO_786 (O_786,N_14756,N_14935);
xnor UO_787 (O_787,N_14652,N_14545);
xor UO_788 (O_788,N_14917,N_14291);
xor UO_789 (O_789,N_14981,N_14772);
nor UO_790 (O_790,N_14434,N_14658);
xor UO_791 (O_791,N_14744,N_14336);
nand UO_792 (O_792,N_14504,N_14934);
xor UO_793 (O_793,N_14472,N_14926);
xor UO_794 (O_794,N_14490,N_14468);
nand UO_795 (O_795,N_14515,N_14505);
nor UO_796 (O_796,N_14968,N_14857);
or UO_797 (O_797,N_14669,N_14922);
and UO_798 (O_798,N_14606,N_14872);
xnor UO_799 (O_799,N_14332,N_14959);
or UO_800 (O_800,N_14658,N_14527);
and UO_801 (O_801,N_14449,N_14603);
or UO_802 (O_802,N_14584,N_14272);
nand UO_803 (O_803,N_14471,N_14595);
nand UO_804 (O_804,N_14503,N_14535);
nand UO_805 (O_805,N_14969,N_14371);
or UO_806 (O_806,N_14476,N_14418);
or UO_807 (O_807,N_14786,N_14440);
and UO_808 (O_808,N_14351,N_14719);
nand UO_809 (O_809,N_14667,N_14749);
xnor UO_810 (O_810,N_14463,N_14457);
nor UO_811 (O_811,N_14761,N_14411);
and UO_812 (O_812,N_14923,N_14544);
nand UO_813 (O_813,N_14354,N_14404);
nand UO_814 (O_814,N_14952,N_14966);
or UO_815 (O_815,N_14787,N_14393);
nand UO_816 (O_816,N_14526,N_14578);
and UO_817 (O_817,N_14700,N_14486);
nand UO_818 (O_818,N_14353,N_14577);
xor UO_819 (O_819,N_14804,N_14916);
nand UO_820 (O_820,N_14838,N_14362);
nor UO_821 (O_821,N_14377,N_14522);
nor UO_822 (O_822,N_14390,N_14283);
and UO_823 (O_823,N_14917,N_14469);
nor UO_824 (O_824,N_14726,N_14829);
or UO_825 (O_825,N_14644,N_14276);
and UO_826 (O_826,N_14393,N_14992);
nand UO_827 (O_827,N_14780,N_14377);
xnor UO_828 (O_828,N_14301,N_14394);
xor UO_829 (O_829,N_14863,N_14888);
nor UO_830 (O_830,N_14578,N_14762);
nor UO_831 (O_831,N_14413,N_14960);
or UO_832 (O_832,N_14282,N_14803);
nor UO_833 (O_833,N_14804,N_14302);
xnor UO_834 (O_834,N_14669,N_14905);
nor UO_835 (O_835,N_14369,N_14849);
nor UO_836 (O_836,N_14583,N_14432);
or UO_837 (O_837,N_14300,N_14679);
nand UO_838 (O_838,N_14725,N_14774);
or UO_839 (O_839,N_14316,N_14502);
nor UO_840 (O_840,N_14872,N_14481);
and UO_841 (O_841,N_14407,N_14526);
nor UO_842 (O_842,N_14389,N_14558);
or UO_843 (O_843,N_14843,N_14862);
or UO_844 (O_844,N_14518,N_14788);
nor UO_845 (O_845,N_14787,N_14749);
xnor UO_846 (O_846,N_14659,N_14474);
nor UO_847 (O_847,N_14391,N_14251);
and UO_848 (O_848,N_14815,N_14914);
nor UO_849 (O_849,N_14624,N_14351);
nand UO_850 (O_850,N_14921,N_14651);
or UO_851 (O_851,N_14656,N_14390);
nand UO_852 (O_852,N_14355,N_14572);
or UO_853 (O_853,N_14319,N_14367);
nand UO_854 (O_854,N_14789,N_14304);
xnor UO_855 (O_855,N_14944,N_14526);
nor UO_856 (O_856,N_14350,N_14333);
xor UO_857 (O_857,N_14417,N_14252);
nor UO_858 (O_858,N_14826,N_14437);
and UO_859 (O_859,N_14498,N_14410);
xnor UO_860 (O_860,N_14894,N_14768);
and UO_861 (O_861,N_14501,N_14487);
nor UO_862 (O_862,N_14668,N_14678);
xor UO_863 (O_863,N_14809,N_14892);
or UO_864 (O_864,N_14983,N_14267);
nand UO_865 (O_865,N_14449,N_14459);
nand UO_866 (O_866,N_14924,N_14428);
or UO_867 (O_867,N_14631,N_14418);
or UO_868 (O_868,N_14385,N_14837);
and UO_869 (O_869,N_14438,N_14611);
nand UO_870 (O_870,N_14590,N_14598);
or UO_871 (O_871,N_14912,N_14823);
xor UO_872 (O_872,N_14997,N_14413);
nor UO_873 (O_873,N_14967,N_14605);
nand UO_874 (O_874,N_14818,N_14843);
nor UO_875 (O_875,N_14626,N_14951);
or UO_876 (O_876,N_14603,N_14827);
nand UO_877 (O_877,N_14375,N_14331);
and UO_878 (O_878,N_14544,N_14982);
and UO_879 (O_879,N_14395,N_14410);
and UO_880 (O_880,N_14838,N_14896);
nor UO_881 (O_881,N_14371,N_14381);
nand UO_882 (O_882,N_14601,N_14616);
nand UO_883 (O_883,N_14678,N_14348);
nand UO_884 (O_884,N_14695,N_14410);
nand UO_885 (O_885,N_14635,N_14446);
or UO_886 (O_886,N_14510,N_14903);
nand UO_887 (O_887,N_14824,N_14326);
or UO_888 (O_888,N_14987,N_14461);
xnor UO_889 (O_889,N_14658,N_14358);
nand UO_890 (O_890,N_14775,N_14614);
and UO_891 (O_891,N_14483,N_14949);
nor UO_892 (O_892,N_14275,N_14880);
or UO_893 (O_893,N_14615,N_14775);
nor UO_894 (O_894,N_14460,N_14454);
nand UO_895 (O_895,N_14359,N_14961);
or UO_896 (O_896,N_14641,N_14741);
nand UO_897 (O_897,N_14452,N_14775);
and UO_898 (O_898,N_14427,N_14932);
and UO_899 (O_899,N_14926,N_14716);
or UO_900 (O_900,N_14914,N_14390);
or UO_901 (O_901,N_14828,N_14310);
nor UO_902 (O_902,N_14628,N_14784);
nor UO_903 (O_903,N_14557,N_14359);
and UO_904 (O_904,N_14450,N_14910);
or UO_905 (O_905,N_14358,N_14364);
nand UO_906 (O_906,N_14412,N_14276);
xnor UO_907 (O_907,N_14453,N_14910);
nand UO_908 (O_908,N_14837,N_14654);
or UO_909 (O_909,N_14882,N_14444);
or UO_910 (O_910,N_14696,N_14598);
or UO_911 (O_911,N_14581,N_14740);
or UO_912 (O_912,N_14313,N_14563);
nand UO_913 (O_913,N_14370,N_14458);
xnor UO_914 (O_914,N_14308,N_14619);
nand UO_915 (O_915,N_14292,N_14715);
or UO_916 (O_916,N_14375,N_14953);
xnor UO_917 (O_917,N_14949,N_14416);
nand UO_918 (O_918,N_14416,N_14366);
or UO_919 (O_919,N_14876,N_14836);
and UO_920 (O_920,N_14276,N_14504);
nand UO_921 (O_921,N_14773,N_14557);
nand UO_922 (O_922,N_14676,N_14910);
nor UO_923 (O_923,N_14743,N_14725);
and UO_924 (O_924,N_14357,N_14937);
xnor UO_925 (O_925,N_14628,N_14288);
nand UO_926 (O_926,N_14784,N_14902);
or UO_927 (O_927,N_14354,N_14628);
or UO_928 (O_928,N_14799,N_14947);
nor UO_929 (O_929,N_14536,N_14514);
or UO_930 (O_930,N_14570,N_14820);
and UO_931 (O_931,N_14442,N_14570);
nor UO_932 (O_932,N_14969,N_14612);
and UO_933 (O_933,N_14737,N_14385);
or UO_934 (O_934,N_14428,N_14559);
nand UO_935 (O_935,N_14404,N_14927);
and UO_936 (O_936,N_14290,N_14625);
nor UO_937 (O_937,N_14947,N_14364);
xnor UO_938 (O_938,N_14613,N_14947);
nor UO_939 (O_939,N_14435,N_14441);
and UO_940 (O_940,N_14427,N_14675);
xor UO_941 (O_941,N_14670,N_14447);
nor UO_942 (O_942,N_14905,N_14527);
nand UO_943 (O_943,N_14867,N_14384);
nor UO_944 (O_944,N_14646,N_14969);
nand UO_945 (O_945,N_14367,N_14933);
or UO_946 (O_946,N_14265,N_14286);
nand UO_947 (O_947,N_14779,N_14869);
or UO_948 (O_948,N_14779,N_14974);
xnor UO_949 (O_949,N_14691,N_14810);
nor UO_950 (O_950,N_14332,N_14927);
or UO_951 (O_951,N_14994,N_14467);
xnor UO_952 (O_952,N_14395,N_14265);
or UO_953 (O_953,N_14311,N_14333);
nand UO_954 (O_954,N_14502,N_14755);
nor UO_955 (O_955,N_14779,N_14795);
nand UO_956 (O_956,N_14441,N_14554);
nand UO_957 (O_957,N_14424,N_14847);
nand UO_958 (O_958,N_14280,N_14554);
and UO_959 (O_959,N_14661,N_14944);
nor UO_960 (O_960,N_14345,N_14397);
and UO_961 (O_961,N_14842,N_14334);
xor UO_962 (O_962,N_14863,N_14703);
xor UO_963 (O_963,N_14355,N_14663);
nand UO_964 (O_964,N_14254,N_14565);
xnor UO_965 (O_965,N_14438,N_14967);
or UO_966 (O_966,N_14883,N_14961);
nand UO_967 (O_967,N_14320,N_14753);
or UO_968 (O_968,N_14478,N_14806);
nor UO_969 (O_969,N_14562,N_14626);
nor UO_970 (O_970,N_14720,N_14819);
xnor UO_971 (O_971,N_14435,N_14614);
and UO_972 (O_972,N_14288,N_14399);
or UO_973 (O_973,N_14808,N_14891);
xnor UO_974 (O_974,N_14901,N_14579);
and UO_975 (O_975,N_14273,N_14578);
and UO_976 (O_976,N_14334,N_14637);
nand UO_977 (O_977,N_14256,N_14741);
and UO_978 (O_978,N_14502,N_14741);
or UO_979 (O_979,N_14470,N_14966);
nor UO_980 (O_980,N_14661,N_14305);
xor UO_981 (O_981,N_14579,N_14606);
xnor UO_982 (O_982,N_14400,N_14367);
and UO_983 (O_983,N_14638,N_14711);
nor UO_984 (O_984,N_14716,N_14859);
and UO_985 (O_985,N_14970,N_14829);
or UO_986 (O_986,N_14792,N_14643);
nand UO_987 (O_987,N_14318,N_14602);
nor UO_988 (O_988,N_14921,N_14499);
nand UO_989 (O_989,N_14756,N_14985);
or UO_990 (O_990,N_14466,N_14897);
nor UO_991 (O_991,N_14886,N_14412);
nor UO_992 (O_992,N_14397,N_14646);
or UO_993 (O_993,N_14923,N_14822);
or UO_994 (O_994,N_14669,N_14908);
xor UO_995 (O_995,N_14636,N_14424);
xnor UO_996 (O_996,N_14633,N_14331);
xor UO_997 (O_997,N_14842,N_14498);
or UO_998 (O_998,N_14457,N_14764);
and UO_999 (O_999,N_14850,N_14691);
or UO_1000 (O_1000,N_14694,N_14550);
xnor UO_1001 (O_1001,N_14786,N_14827);
nor UO_1002 (O_1002,N_14255,N_14689);
xor UO_1003 (O_1003,N_14642,N_14805);
nor UO_1004 (O_1004,N_14372,N_14625);
xnor UO_1005 (O_1005,N_14515,N_14663);
nand UO_1006 (O_1006,N_14732,N_14612);
or UO_1007 (O_1007,N_14563,N_14304);
or UO_1008 (O_1008,N_14835,N_14699);
or UO_1009 (O_1009,N_14687,N_14820);
or UO_1010 (O_1010,N_14552,N_14470);
or UO_1011 (O_1011,N_14410,N_14340);
nand UO_1012 (O_1012,N_14363,N_14576);
nor UO_1013 (O_1013,N_14644,N_14490);
or UO_1014 (O_1014,N_14944,N_14287);
or UO_1015 (O_1015,N_14701,N_14449);
or UO_1016 (O_1016,N_14967,N_14409);
nand UO_1017 (O_1017,N_14865,N_14965);
or UO_1018 (O_1018,N_14633,N_14387);
xnor UO_1019 (O_1019,N_14507,N_14324);
nand UO_1020 (O_1020,N_14250,N_14465);
nand UO_1021 (O_1021,N_14383,N_14254);
and UO_1022 (O_1022,N_14934,N_14273);
and UO_1023 (O_1023,N_14372,N_14481);
xnor UO_1024 (O_1024,N_14482,N_14252);
and UO_1025 (O_1025,N_14891,N_14834);
nor UO_1026 (O_1026,N_14342,N_14917);
xor UO_1027 (O_1027,N_14886,N_14481);
xor UO_1028 (O_1028,N_14377,N_14417);
and UO_1029 (O_1029,N_14315,N_14480);
xor UO_1030 (O_1030,N_14755,N_14916);
or UO_1031 (O_1031,N_14354,N_14489);
or UO_1032 (O_1032,N_14719,N_14754);
or UO_1033 (O_1033,N_14620,N_14869);
xnor UO_1034 (O_1034,N_14439,N_14664);
nand UO_1035 (O_1035,N_14627,N_14961);
or UO_1036 (O_1036,N_14375,N_14928);
xor UO_1037 (O_1037,N_14485,N_14393);
or UO_1038 (O_1038,N_14821,N_14494);
nor UO_1039 (O_1039,N_14719,N_14608);
nor UO_1040 (O_1040,N_14740,N_14416);
nand UO_1041 (O_1041,N_14644,N_14282);
nand UO_1042 (O_1042,N_14529,N_14322);
nor UO_1043 (O_1043,N_14579,N_14799);
or UO_1044 (O_1044,N_14861,N_14692);
and UO_1045 (O_1045,N_14349,N_14607);
nor UO_1046 (O_1046,N_14824,N_14397);
and UO_1047 (O_1047,N_14927,N_14298);
nand UO_1048 (O_1048,N_14397,N_14914);
xnor UO_1049 (O_1049,N_14278,N_14664);
and UO_1050 (O_1050,N_14293,N_14445);
xor UO_1051 (O_1051,N_14722,N_14658);
and UO_1052 (O_1052,N_14323,N_14777);
nor UO_1053 (O_1053,N_14371,N_14307);
and UO_1054 (O_1054,N_14389,N_14876);
nand UO_1055 (O_1055,N_14662,N_14996);
nor UO_1056 (O_1056,N_14407,N_14908);
or UO_1057 (O_1057,N_14842,N_14328);
or UO_1058 (O_1058,N_14775,N_14355);
nor UO_1059 (O_1059,N_14373,N_14385);
xnor UO_1060 (O_1060,N_14405,N_14372);
or UO_1061 (O_1061,N_14509,N_14868);
nor UO_1062 (O_1062,N_14730,N_14849);
and UO_1063 (O_1063,N_14543,N_14695);
nor UO_1064 (O_1064,N_14589,N_14638);
or UO_1065 (O_1065,N_14617,N_14303);
nand UO_1066 (O_1066,N_14272,N_14687);
nand UO_1067 (O_1067,N_14764,N_14637);
xnor UO_1068 (O_1068,N_14652,N_14904);
nor UO_1069 (O_1069,N_14263,N_14397);
xnor UO_1070 (O_1070,N_14764,N_14880);
and UO_1071 (O_1071,N_14963,N_14701);
nand UO_1072 (O_1072,N_14647,N_14281);
nand UO_1073 (O_1073,N_14302,N_14966);
or UO_1074 (O_1074,N_14909,N_14407);
nor UO_1075 (O_1075,N_14787,N_14836);
or UO_1076 (O_1076,N_14408,N_14366);
and UO_1077 (O_1077,N_14681,N_14879);
nand UO_1078 (O_1078,N_14282,N_14826);
or UO_1079 (O_1079,N_14706,N_14307);
or UO_1080 (O_1080,N_14896,N_14738);
nor UO_1081 (O_1081,N_14865,N_14689);
and UO_1082 (O_1082,N_14948,N_14854);
nand UO_1083 (O_1083,N_14748,N_14451);
xor UO_1084 (O_1084,N_14390,N_14808);
nor UO_1085 (O_1085,N_14544,N_14661);
nand UO_1086 (O_1086,N_14975,N_14263);
xor UO_1087 (O_1087,N_14966,N_14776);
or UO_1088 (O_1088,N_14612,N_14666);
or UO_1089 (O_1089,N_14654,N_14563);
xnor UO_1090 (O_1090,N_14601,N_14531);
xnor UO_1091 (O_1091,N_14504,N_14445);
or UO_1092 (O_1092,N_14501,N_14598);
and UO_1093 (O_1093,N_14563,N_14807);
xor UO_1094 (O_1094,N_14435,N_14751);
and UO_1095 (O_1095,N_14812,N_14385);
and UO_1096 (O_1096,N_14282,N_14846);
nand UO_1097 (O_1097,N_14782,N_14481);
nand UO_1098 (O_1098,N_14952,N_14308);
nor UO_1099 (O_1099,N_14572,N_14631);
nand UO_1100 (O_1100,N_14437,N_14481);
nand UO_1101 (O_1101,N_14337,N_14779);
xor UO_1102 (O_1102,N_14563,N_14550);
nor UO_1103 (O_1103,N_14659,N_14327);
nor UO_1104 (O_1104,N_14641,N_14721);
nand UO_1105 (O_1105,N_14476,N_14569);
and UO_1106 (O_1106,N_14322,N_14301);
and UO_1107 (O_1107,N_14379,N_14339);
nor UO_1108 (O_1108,N_14786,N_14933);
nor UO_1109 (O_1109,N_14390,N_14500);
nand UO_1110 (O_1110,N_14813,N_14887);
xnor UO_1111 (O_1111,N_14791,N_14993);
nand UO_1112 (O_1112,N_14556,N_14701);
and UO_1113 (O_1113,N_14348,N_14338);
or UO_1114 (O_1114,N_14986,N_14263);
nor UO_1115 (O_1115,N_14990,N_14675);
or UO_1116 (O_1116,N_14292,N_14880);
xor UO_1117 (O_1117,N_14573,N_14423);
xnor UO_1118 (O_1118,N_14715,N_14330);
or UO_1119 (O_1119,N_14541,N_14620);
or UO_1120 (O_1120,N_14722,N_14422);
and UO_1121 (O_1121,N_14287,N_14488);
or UO_1122 (O_1122,N_14519,N_14430);
nand UO_1123 (O_1123,N_14847,N_14578);
and UO_1124 (O_1124,N_14510,N_14702);
and UO_1125 (O_1125,N_14749,N_14925);
and UO_1126 (O_1126,N_14401,N_14952);
and UO_1127 (O_1127,N_14734,N_14372);
nor UO_1128 (O_1128,N_14947,N_14952);
or UO_1129 (O_1129,N_14886,N_14782);
xnor UO_1130 (O_1130,N_14589,N_14660);
and UO_1131 (O_1131,N_14393,N_14510);
nor UO_1132 (O_1132,N_14681,N_14425);
nand UO_1133 (O_1133,N_14278,N_14454);
or UO_1134 (O_1134,N_14578,N_14963);
nand UO_1135 (O_1135,N_14794,N_14978);
xnor UO_1136 (O_1136,N_14709,N_14928);
xnor UO_1137 (O_1137,N_14558,N_14896);
xnor UO_1138 (O_1138,N_14610,N_14819);
or UO_1139 (O_1139,N_14857,N_14439);
xor UO_1140 (O_1140,N_14290,N_14917);
xnor UO_1141 (O_1141,N_14660,N_14455);
and UO_1142 (O_1142,N_14323,N_14867);
and UO_1143 (O_1143,N_14365,N_14489);
or UO_1144 (O_1144,N_14524,N_14872);
xor UO_1145 (O_1145,N_14553,N_14600);
nor UO_1146 (O_1146,N_14923,N_14642);
or UO_1147 (O_1147,N_14621,N_14744);
nand UO_1148 (O_1148,N_14895,N_14655);
xnor UO_1149 (O_1149,N_14433,N_14410);
nor UO_1150 (O_1150,N_14759,N_14576);
xnor UO_1151 (O_1151,N_14573,N_14354);
xor UO_1152 (O_1152,N_14275,N_14913);
xnor UO_1153 (O_1153,N_14762,N_14556);
xnor UO_1154 (O_1154,N_14397,N_14366);
or UO_1155 (O_1155,N_14434,N_14743);
and UO_1156 (O_1156,N_14680,N_14832);
nand UO_1157 (O_1157,N_14546,N_14367);
nand UO_1158 (O_1158,N_14311,N_14617);
and UO_1159 (O_1159,N_14318,N_14779);
or UO_1160 (O_1160,N_14605,N_14961);
and UO_1161 (O_1161,N_14400,N_14968);
and UO_1162 (O_1162,N_14821,N_14272);
nor UO_1163 (O_1163,N_14702,N_14301);
or UO_1164 (O_1164,N_14892,N_14255);
and UO_1165 (O_1165,N_14857,N_14745);
nor UO_1166 (O_1166,N_14340,N_14326);
xor UO_1167 (O_1167,N_14624,N_14969);
nand UO_1168 (O_1168,N_14862,N_14372);
nor UO_1169 (O_1169,N_14935,N_14703);
or UO_1170 (O_1170,N_14926,N_14274);
xnor UO_1171 (O_1171,N_14628,N_14867);
nand UO_1172 (O_1172,N_14586,N_14929);
nand UO_1173 (O_1173,N_14318,N_14518);
xor UO_1174 (O_1174,N_14781,N_14889);
or UO_1175 (O_1175,N_14516,N_14360);
nand UO_1176 (O_1176,N_14677,N_14568);
nor UO_1177 (O_1177,N_14720,N_14702);
nand UO_1178 (O_1178,N_14721,N_14498);
and UO_1179 (O_1179,N_14884,N_14262);
nand UO_1180 (O_1180,N_14842,N_14641);
or UO_1181 (O_1181,N_14279,N_14997);
nor UO_1182 (O_1182,N_14357,N_14584);
nor UO_1183 (O_1183,N_14964,N_14651);
nand UO_1184 (O_1184,N_14553,N_14407);
xor UO_1185 (O_1185,N_14276,N_14291);
nand UO_1186 (O_1186,N_14934,N_14890);
nand UO_1187 (O_1187,N_14918,N_14590);
or UO_1188 (O_1188,N_14923,N_14761);
nand UO_1189 (O_1189,N_14672,N_14807);
nor UO_1190 (O_1190,N_14261,N_14689);
or UO_1191 (O_1191,N_14969,N_14337);
nand UO_1192 (O_1192,N_14903,N_14279);
xor UO_1193 (O_1193,N_14374,N_14485);
or UO_1194 (O_1194,N_14584,N_14359);
or UO_1195 (O_1195,N_14991,N_14535);
and UO_1196 (O_1196,N_14412,N_14536);
and UO_1197 (O_1197,N_14886,N_14641);
nor UO_1198 (O_1198,N_14919,N_14753);
nor UO_1199 (O_1199,N_14323,N_14918);
and UO_1200 (O_1200,N_14416,N_14895);
xor UO_1201 (O_1201,N_14864,N_14469);
nand UO_1202 (O_1202,N_14532,N_14566);
nor UO_1203 (O_1203,N_14359,N_14653);
nand UO_1204 (O_1204,N_14581,N_14377);
and UO_1205 (O_1205,N_14874,N_14318);
nand UO_1206 (O_1206,N_14661,N_14368);
nand UO_1207 (O_1207,N_14486,N_14361);
nor UO_1208 (O_1208,N_14326,N_14899);
or UO_1209 (O_1209,N_14283,N_14305);
nor UO_1210 (O_1210,N_14600,N_14978);
xnor UO_1211 (O_1211,N_14290,N_14611);
nor UO_1212 (O_1212,N_14859,N_14880);
xnor UO_1213 (O_1213,N_14328,N_14680);
nor UO_1214 (O_1214,N_14739,N_14865);
nand UO_1215 (O_1215,N_14997,N_14442);
xor UO_1216 (O_1216,N_14683,N_14822);
and UO_1217 (O_1217,N_14482,N_14389);
nand UO_1218 (O_1218,N_14957,N_14402);
or UO_1219 (O_1219,N_14548,N_14798);
nor UO_1220 (O_1220,N_14786,N_14940);
nor UO_1221 (O_1221,N_14856,N_14587);
nand UO_1222 (O_1222,N_14723,N_14310);
nor UO_1223 (O_1223,N_14273,N_14303);
or UO_1224 (O_1224,N_14775,N_14316);
and UO_1225 (O_1225,N_14444,N_14525);
nor UO_1226 (O_1226,N_14762,N_14281);
or UO_1227 (O_1227,N_14788,N_14779);
xnor UO_1228 (O_1228,N_14279,N_14515);
or UO_1229 (O_1229,N_14420,N_14789);
nand UO_1230 (O_1230,N_14747,N_14858);
nand UO_1231 (O_1231,N_14777,N_14366);
nand UO_1232 (O_1232,N_14586,N_14959);
nor UO_1233 (O_1233,N_14859,N_14439);
nor UO_1234 (O_1234,N_14846,N_14829);
and UO_1235 (O_1235,N_14596,N_14893);
and UO_1236 (O_1236,N_14802,N_14942);
nand UO_1237 (O_1237,N_14511,N_14491);
and UO_1238 (O_1238,N_14403,N_14324);
nand UO_1239 (O_1239,N_14521,N_14419);
and UO_1240 (O_1240,N_14900,N_14652);
or UO_1241 (O_1241,N_14356,N_14940);
xor UO_1242 (O_1242,N_14511,N_14396);
nor UO_1243 (O_1243,N_14927,N_14556);
or UO_1244 (O_1244,N_14639,N_14437);
nor UO_1245 (O_1245,N_14466,N_14406);
or UO_1246 (O_1246,N_14269,N_14535);
or UO_1247 (O_1247,N_14754,N_14566);
nand UO_1248 (O_1248,N_14990,N_14487);
nor UO_1249 (O_1249,N_14629,N_14466);
nor UO_1250 (O_1250,N_14588,N_14425);
xor UO_1251 (O_1251,N_14727,N_14338);
xor UO_1252 (O_1252,N_14528,N_14904);
and UO_1253 (O_1253,N_14762,N_14708);
nor UO_1254 (O_1254,N_14904,N_14998);
xor UO_1255 (O_1255,N_14251,N_14729);
nand UO_1256 (O_1256,N_14949,N_14598);
and UO_1257 (O_1257,N_14451,N_14862);
or UO_1258 (O_1258,N_14696,N_14467);
xor UO_1259 (O_1259,N_14417,N_14881);
nor UO_1260 (O_1260,N_14633,N_14472);
nand UO_1261 (O_1261,N_14358,N_14420);
or UO_1262 (O_1262,N_14741,N_14569);
xnor UO_1263 (O_1263,N_14413,N_14329);
xor UO_1264 (O_1264,N_14971,N_14311);
or UO_1265 (O_1265,N_14793,N_14625);
xor UO_1266 (O_1266,N_14465,N_14682);
xor UO_1267 (O_1267,N_14947,N_14401);
nor UO_1268 (O_1268,N_14363,N_14902);
nand UO_1269 (O_1269,N_14355,N_14356);
nor UO_1270 (O_1270,N_14442,N_14326);
nand UO_1271 (O_1271,N_14565,N_14547);
xor UO_1272 (O_1272,N_14732,N_14921);
nand UO_1273 (O_1273,N_14903,N_14806);
and UO_1274 (O_1274,N_14443,N_14460);
and UO_1275 (O_1275,N_14948,N_14927);
xor UO_1276 (O_1276,N_14438,N_14643);
nand UO_1277 (O_1277,N_14556,N_14982);
and UO_1278 (O_1278,N_14703,N_14654);
or UO_1279 (O_1279,N_14799,N_14509);
xor UO_1280 (O_1280,N_14981,N_14379);
and UO_1281 (O_1281,N_14812,N_14479);
or UO_1282 (O_1282,N_14296,N_14400);
or UO_1283 (O_1283,N_14588,N_14489);
or UO_1284 (O_1284,N_14300,N_14838);
nand UO_1285 (O_1285,N_14382,N_14458);
nand UO_1286 (O_1286,N_14448,N_14829);
nor UO_1287 (O_1287,N_14904,N_14927);
or UO_1288 (O_1288,N_14486,N_14988);
nor UO_1289 (O_1289,N_14821,N_14644);
nand UO_1290 (O_1290,N_14680,N_14375);
nand UO_1291 (O_1291,N_14840,N_14293);
and UO_1292 (O_1292,N_14955,N_14928);
nor UO_1293 (O_1293,N_14913,N_14673);
nor UO_1294 (O_1294,N_14509,N_14983);
nand UO_1295 (O_1295,N_14497,N_14406);
nor UO_1296 (O_1296,N_14915,N_14737);
and UO_1297 (O_1297,N_14991,N_14493);
or UO_1298 (O_1298,N_14298,N_14442);
xnor UO_1299 (O_1299,N_14719,N_14262);
nor UO_1300 (O_1300,N_14639,N_14855);
nor UO_1301 (O_1301,N_14350,N_14768);
or UO_1302 (O_1302,N_14302,N_14984);
xor UO_1303 (O_1303,N_14472,N_14930);
and UO_1304 (O_1304,N_14968,N_14616);
nand UO_1305 (O_1305,N_14640,N_14554);
nor UO_1306 (O_1306,N_14547,N_14357);
or UO_1307 (O_1307,N_14775,N_14721);
and UO_1308 (O_1308,N_14945,N_14375);
or UO_1309 (O_1309,N_14850,N_14893);
nand UO_1310 (O_1310,N_14845,N_14408);
xor UO_1311 (O_1311,N_14288,N_14499);
or UO_1312 (O_1312,N_14444,N_14867);
or UO_1313 (O_1313,N_14798,N_14919);
xnor UO_1314 (O_1314,N_14506,N_14280);
and UO_1315 (O_1315,N_14356,N_14551);
nor UO_1316 (O_1316,N_14366,N_14409);
or UO_1317 (O_1317,N_14291,N_14613);
nor UO_1318 (O_1318,N_14358,N_14896);
nor UO_1319 (O_1319,N_14896,N_14699);
nand UO_1320 (O_1320,N_14619,N_14635);
nand UO_1321 (O_1321,N_14433,N_14338);
xnor UO_1322 (O_1322,N_14532,N_14452);
or UO_1323 (O_1323,N_14878,N_14592);
nand UO_1324 (O_1324,N_14804,N_14958);
and UO_1325 (O_1325,N_14365,N_14285);
xor UO_1326 (O_1326,N_14401,N_14682);
nand UO_1327 (O_1327,N_14851,N_14517);
nand UO_1328 (O_1328,N_14392,N_14838);
nand UO_1329 (O_1329,N_14414,N_14421);
nor UO_1330 (O_1330,N_14321,N_14317);
or UO_1331 (O_1331,N_14735,N_14626);
xor UO_1332 (O_1332,N_14696,N_14393);
nor UO_1333 (O_1333,N_14338,N_14580);
nand UO_1334 (O_1334,N_14581,N_14776);
xor UO_1335 (O_1335,N_14422,N_14475);
nor UO_1336 (O_1336,N_14962,N_14882);
nand UO_1337 (O_1337,N_14639,N_14712);
nor UO_1338 (O_1338,N_14373,N_14391);
and UO_1339 (O_1339,N_14341,N_14657);
nor UO_1340 (O_1340,N_14382,N_14579);
or UO_1341 (O_1341,N_14449,N_14370);
xor UO_1342 (O_1342,N_14509,N_14431);
or UO_1343 (O_1343,N_14416,N_14346);
or UO_1344 (O_1344,N_14922,N_14897);
nor UO_1345 (O_1345,N_14252,N_14887);
nand UO_1346 (O_1346,N_14626,N_14921);
xor UO_1347 (O_1347,N_14366,N_14539);
nor UO_1348 (O_1348,N_14666,N_14782);
nor UO_1349 (O_1349,N_14912,N_14768);
or UO_1350 (O_1350,N_14515,N_14802);
and UO_1351 (O_1351,N_14967,N_14963);
nand UO_1352 (O_1352,N_14522,N_14893);
nor UO_1353 (O_1353,N_14280,N_14624);
nand UO_1354 (O_1354,N_14931,N_14510);
xnor UO_1355 (O_1355,N_14324,N_14634);
and UO_1356 (O_1356,N_14814,N_14641);
xnor UO_1357 (O_1357,N_14708,N_14254);
or UO_1358 (O_1358,N_14562,N_14437);
and UO_1359 (O_1359,N_14692,N_14572);
nor UO_1360 (O_1360,N_14413,N_14578);
nor UO_1361 (O_1361,N_14991,N_14421);
nand UO_1362 (O_1362,N_14768,N_14786);
nand UO_1363 (O_1363,N_14471,N_14796);
and UO_1364 (O_1364,N_14833,N_14630);
and UO_1365 (O_1365,N_14662,N_14749);
or UO_1366 (O_1366,N_14270,N_14597);
nor UO_1367 (O_1367,N_14775,N_14535);
or UO_1368 (O_1368,N_14515,N_14936);
xor UO_1369 (O_1369,N_14588,N_14930);
xnor UO_1370 (O_1370,N_14652,N_14301);
nand UO_1371 (O_1371,N_14499,N_14573);
nor UO_1372 (O_1372,N_14895,N_14445);
or UO_1373 (O_1373,N_14507,N_14687);
xnor UO_1374 (O_1374,N_14533,N_14994);
and UO_1375 (O_1375,N_14914,N_14709);
and UO_1376 (O_1376,N_14840,N_14267);
xnor UO_1377 (O_1377,N_14668,N_14348);
xnor UO_1378 (O_1378,N_14321,N_14442);
and UO_1379 (O_1379,N_14446,N_14908);
xor UO_1380 (O_1380,N_14743,N_14876);
xor UO_1381 (O_1381,N_14263,N_14500);
and UO_1382 (O_1382,N_14575,N_14554);
xor UO_1383 (O_1383,N_14478,N_14553);
nor UO_1384 (O_1384,N_14744,N_14647);
and UO_1385 (O_1385,N_14308,N_14295);
xnor UO_1386 (O_1386,N_14758,N_14737);
and UO_1387 (O_1387,N_14266,N_14678);
nand UO_1388 (O_1388,N_14808,N_14780);
or UO_1389 (O_1389,N_14855,N_14996);
xnor UO_1390 (O_1390,N_14724,N_14835);
xor UO_1391 (O_1391,N_14763,N_14985);
xnor UO_1392 (O_1392,N_14600,N_14664);
or UO_1393 (O_1393,N_14904,N_14436);
nor UO_1394 (O_1394,N_14367,N_14886);
nor UO_1395 (O_1395,N_14879,N_14455);
nand UO_1396 (O_1396,N_14378,N_14777);
xnor UO_1397 (O_1397,N_14471,N_14528);
nor UO_1398 (O_1398,N_14447,N_14310);
and UO_1399 (O_1399,N_14350,N_14575);
or UO_1400 (O_1400,N_14494,N_14370);
nand UO_1401 (O_1401,N_14537,N_14559);
or UO_1402 (O_1402,N_14690,N_14475);
or UO_1403 (O_1403,N_14435,N_14302);
xnor UO_1404 (O_1404,N_14888,N_14342);
nor UO_1405 (O_1405,N_14553,N_14422);
nor UO_1406 (O_1406,N_14923,N_14400);
and UO_1407 (O_1407,N_14452,N_14250);
or UO_1408 (O_1408,N_14483,N_14376);
nor UO_1409 (O_1409,N_14391,N_14393);
nor UO_1410 (O_1410,N_14858,N_14538);
or UO_1411 (O_1411,N_14363,N_14979);
nand UO_1412 (O_1412,N_14792,N_14484);
and UO_1413 (O_1413,N_14267,N_14496);
nor UO_1414 (O_1414,N_14996,N_14440);
and UO_1415 (O_1415,N_14967,N_14906);
nand UO_1416 (O_1416,N_14318,N_14912);
or UO_1417 (O_1417,N_14300,N_14702);
nor UO_1418 (O_1418,N_14988,N_14259);
xnor UO_1419 (O_1419,N_14559,N_14330);
and UO_1420 (O_1420,N_14399,N_14281);
xor UO_1421 (O_1421,N_14617,N_14480);
nand UO_1422 (O_1422,N_14470,N_14584);
and UO_1423 (O_1423,N_14613,N_14345);
or UO_1424 (O_1424,N_14336,N_14840);
or UO_1425 (O_1425,N_14629,N_14269);
nand UO_1426 (O_1426,N_14633,N_14460);
or UO_1427 (O_1427,N_14789,N_14502);
nor UO_1428 (O_1428,N_14801,N_14484);
nor UO_1429 (O_1429,N_14841,N_14827);
nand UO_1430 (O_1430,N_14570,N_14477);
or UO_1431 (O_1431,N_14596,N_14739);
and UO_1432 (O_1432,N_14308,N_14449);
nand UO_1433 (O_1433,N_14585,N_14667);
and UO_1434 (O_1434,N_14566,N_14369);
and UO_1435 (O_1435,N_14665,N_14443);
nor UO_1436 (O_1436,N_14628,N_14623);
nor UO_1437 (O_1437,N_14470,N_14733);
nor UO_1438 (O_1438,N_14316,N_14916);
and UO_1439 (O_1439,N_14540,N_14707);
nand UO_1440 (O_1440,N_14911,N_14431);
and UO_1441 (O_1441,N_14319,N_14661);
xor UO_1442 (O_1442,N_14861,N_14250);
and UO_1443 (O_1443,N_14357,N_14626);
xnor UO_1444 (O_1444,N_14458,N_14378);
nor UO_1445 (O_1445,N_14329,N_14403);
nor UO_1446 (O_1446,N_14909,N_14261);
xor UO_1447 (O_1447,N_14267,N_14495);
and UO_1448 (O_1448,N_14513,N_14328);
nand UO_1449 (O_1449,N_14358,N_14329);
nor UO_1450 (O_1450,N_14736,N_14938);
or UO_1451 (O_1451,N_14632,N_14423);
nor UO_1452 (O_1452,N_14497,N_14325);
and UO_1453 (O_1453,N_14861,N_14750);
xor UO_1454 (O_1454,N_14593,N_14751);
xnor UO_1455 (O_1455,N_14647,N_14434);
nor UO_1456 (O_1456,N_14671,N_14286);
xor UO_1457 (O_1457,N_14629,N_14579);
xor UO_1458 (O_1458,N_14328,N_14777);
and UO_1459 (O_1459,N_14408,N_14355);
nor UO_1460 (O_1460,N_14981,N_14408);
nor UO_1461 (O_1461,N_14508,N_14541);
nor UO_1462 (O_1462,N_14426,N_14455);
nand UO_1463 (O_1463,N_14826,N_14308);
nand UO_1464 (O_1464,N_14981,N_14254);
nand UO_1465 (O_1465,N_14964,N_14454);
and UO_1466 (O_1466,N_14822,N_14498);
and UO_1467 (O_1467,N_14567,N_14849);
nor UO_1468 (O_1468,N_14516,N_14666);
nand UO_1469 (O_1469,N_14255,N_14618);
nor UO_1470 (O_1470,N_14817,N_14618);
or UO_1471 (O_1471,N_14490,N_14498);
and UO_1472 (O_1472,N_14831,N_14708);
nand UO_1473 (O_1473,N_14316,N_14792);
nand UO_1474 (O_1474,N_14383,N_14584);
or UO_1475 (O_1475,N_14277,N_14593);
nand UO_1476 (O_1476,N_14645,N_14542);
and UO_1477 (O_1477,N_14584,N_14260);
nor UO_1478 (O_1478,N_14271,N_14790);
xnor UO_1479 (O_1479,N_14623,N_14723);
or UO_1480 (O_1480,N_14891,N_14616);
xor UO_1481 (O_1481,N_14344,N_14297);
nand UO_1482 (O_1482,N_14751,N_14761);
nor UO_1483 (O_1483,N_14847,N_14588);
nand UO_1484 (O_1484,N_14670,N_14606);
nand UO_1485 (O_1485,N_14749,N_14251);
nand UO_1486 (O_1486,N_14391,N_14797);
or UO_1487 (O_1487,N_14661,N_14410);
or UO_1488 (O_1488,N_14468,N_14975);
nor UO_1489 (O_1489,N_14668,N_14755);
and UO_1490 (O_1490,N_14647,N_14856);
xnor UO_1491 (O_1491,N_14832,N_14560);
and UO_1492 (O_1492,N_14258,N_14518);
or UO_1493 (O_1493,N_14372,N_14547);
nor UO_1494 (O_1494,N_14633,N_14532);
nand UO_1495 (O_1495,N_14618,N_14507);
and UO_1496 (O_1496,N_14978,N_14871);
and UO_1497 (O_1497,N_14923,N_14630);
or UO_1498 (O_1498,N_14837,N_14553);
nand UO_1499 (O_1499,N_14561,N_14776);
or UO_1500 (O_1500,N_14939,N_14983);
nand UO_1501 (O_1501,N_14776,N_14559);
and UO_1502 (O_1502,N_14929,N_14568);
nor UO_1503 (O_1503,N_14448,N_14781);
xnor UO_1504 (O_1504,N_14391,N_14779);
or UO_1505 (O_1505,N_14527,N_14677);
xnor UO_1506 (O_1506,N_14887,N_14406);
and UO_1507 (O_1507,N_14574,N_14820);
and UO_1508 (O_1508,N_14920,N_14926);
or UO_1509 (O_1509,N_14559,N_14873);
or UO_1510 (O_1510,N_14984,N_14695);
nor UO_1511 (O_1511,N_14376,N_14706);
or UO_1512 (O_1512,N_14449,N_14884);
nor UO_1513 (O_1513,N_14589,N_14446);
or UO_1514 (O_1514,N_14634,N_14786);
and UO_1515 (O_1515,N_14294,N_14949);
and UO_1516 (O_1516,N_14502,N_14582);
or UO_1517 (O_1517,N_14419,N_14935);
nor UO_1518 (O_1518,N_14685,N_14822);
nor UO_1519 (O_1519,N_14540,N_14498);
xnor UO_1520 (O_1520,N_14497,N_14779);
nand UO_1521 (O_1521,N_14842,N_14920);
or UO_1522 (O_1522,N_14921,N_14745);
or UO_1523 (O_1523,N_14967,N_14819);
nand UO_1524 (O_1524,N_14861,N_14329);
xnor UO_1525 (O_1525,N_14304,N_14600);
nor UO_1526 (O_1526,N_14655,N_14675);
and UO_1527 (O_1527,N_14741,N_14766);
or UO_1528 (O_1528,N_14985,N_14317);
nand UO_1529 (O_1529,N_14428,N_14583);
xnor UO_1530 (O_1530,N_14675,N_14769);
and UO_1531 (O_1531,N_14974,N_14945);
nor UO_1532 (O_1532,N_14885,N_14423);
and UO_1533 (O_1533,N_14686,N_14650);
nand UO_1534 (O_1534,N_14528,N_14550);
and UO_1535 (O_1535,N_14409,N_14626);
xor UO_1536 (O_1536,N_14626,N_14400);
and UO_1537 (O_1537,N_14564,N_14741);
nand UO_1538 (O_1538,N_14389,N_14809);
nand UO_1539 (O_1539,N_14320,N_14376);
and UO_1540 (O_1540,N_14575,N_14367);
nand UO_1541 (O_1541,N_14378,N_14871);
or UO_1542 (O_1542,N_14494,N_14307);
or UO_1543 (O_1543,N_14997,N_14328);
and UO_1544 (O_1544,N_14286,N_14543);
nor UO_1545 (O_1545,N_14805,N_14350);
xor UO_1546 (O_1546,N_14433,N_14800);
nand UO_1547 (O_1547,N_14776,N_14550);
nor UO_1548 (O_1548,N_14415,N_14366);
or UO_1549 (O_1549,N_14288,N_14578);
and UO_1550 (O_1550,N_14880,N_14912);
or UO_1551 (O_1551,N_14542,N_14813);
nand UO_1552 (O_1552,N_14284,N_14727);
and UO_1553 (O_1553,N_14905,N_14447);
nand UO_1554 (O_1554,N_14583,N_14729);
xnor UO_1555 (O_1555,N_14489,N_14857);
and UO_1556 (O_1556,N_14263,N_14556);
or UO_1557 (O_1557,N_14495,N_14911);
or UO_1558 (O_1558,N_14615,N_14316);
xnor UO_1559 (O_1559,N_14721,N_14369);
or UO_1560 (O_1560,N_14727,N_14425);
nand UO_1561 (O_1561,N_14676,N_14351);
and UO_1562 (O_1562,N_14849,N_14571);
xnor UO_1563 (O_1563,N_14437,N_14740);
xnor UO_1564 (O_1564,N_14773,N_14390);
nand UO_1565 (O_1565,N_14531,N_14845);
nand UO_1566 (O_1566,N_14714,N_14750);
or UO_1567 (O_1567,N_14821,N_14992);
xnor UO_1568 (O_1568,N_14923,N_14769);
xnor UO_1569 (O_1569,N_14687,N_14506);
nor UO_1570 (O_1570,N_14476,N_14350);
and UO_1571 (O_1571,N_14885,N_14437);
nor UO_1572 (O_1572,N_14588,N_14502);
and UO_1573 (O_1573,N_14672,N_14569);
xnor UO_1574 (O_1574,N_14980,N_14495);
and UO_1575 (O_1575,N_14741,N_14254);
nor UO_1576 (O_1576,N_14684,N_14606);
and UO_1577 (O_1577,N_14286,N_14426);
and UO_1578 (O_1578,N_14428,N_14946);
or UO_1579 (O_1579,N_14612,N_14261);
and UO_1580 (O_1580,N_14885,N_14793);
and UO_1581 (O_1581,N_14936,N_14368);
nor UO_1582 (O_1582,N_14638,N_14509);
nand UO_1583 (O_1583,N_14881,N_14694);
nor UO_1584 (O_1584,N_14798,N_14991);
nand UO_1585 (O_1585,N_14583,N_14790);
nor UO_1586 (O_1586,N_14825,N_14856);
nand UO_1587 (O_1587,N_14760,N_14876);
and UO_1588 (O_1588,N_14520,N_14702);
and UO_1589 (O_1589,N_14353,N_14813);
and UO_1590 (O_1590,N_14869,N_14388);
or UO_1591 (O_1591,N_14895,N_14743);
or UO_1592 (O_1592,N_14368,N_14721);
nor UO_1593 (O_1593,N_14819,N_14490);
xnor UO_1594 (O_1594,N_14555,N_14534);
xor UO_1595 (O_1595,N_14526,N_14342);
and UO_1596 (O_1596,N_14895,N_14425);
or UO_1597 (O_1597,N_14521,N_14454);
or UO_1598 (O_1598,N_14648,N_14681);
nand UO_1599 (O_1599,N_14296,N_14953);
or UO_1600 (O_1600,N_14931,N_14462);
xnor UO_1601 (O_1601,N_14834,N_14419);
nor UO_1602 (O_1602,N_14695,N_14546);
xor UO_1603 (O_1603,N_14849,N_14827);
nand UO_1604 (O_1604,N_14453,N_14300);
and UO_1605 (O_1605,N_14806,N_14556);
nand UO_1606 (O_1606,N_14834,N_14828);
nand UO_1607 (O_1607,N_14793,N_14990);
and UO_1608 (O_1608,N_14649,N_14899);
nand UO_1609 (O_1609,N_14473,N_14607);
nor UO_1610 (O_1610,N_14844,N_14322);
and UO_1611 (O_1611,N_14521,N_14313);
xor UO_1612 (O_1612,N_14370,N_14415);
or UO_1613 (O_1613,N_14520,N_14372);
nand UO_1614 (O_1614,N_14894,N_14959);
nand UO_1615 (O_1615,N_14341,N_14941);
or UO_1616 (O_1616,N_14740,N_14381);
or UO_1617 (O_1617,N_14821,N_14250);
and UO_1618 (O_1618,N_14842,N_14861);
and UO_1619 (O_1619,N_14754,N_14328);
and UO_1620 (O_1620,N_14845,N_14342);
and UO_1621 (O_1621,N_14475,N_14411);
or UO_1622 (O_1622,N_14616,N_14422);
and UO_1623 (O_1623,N_14645,N_14950);
or UO_1624 (O_1624,N_14377,N_14269);
nor UO_1625 (O_1625,N_14851,N_14803);
nor UO_1626 (O_1626,N_14537,N_14273);
nor UO_1627 (O_1627,N_14349,N_14436);
and UO_1628 (O_1628,N_14283,N_14425);
nor UO_1629 (O_1629,N_14922,N_14652);
nand UO_1630 (O_1630,N_14330,N_14279);
nand UO_1631 (O_1631,N_14814,N_14444);
xnor UO_1632 (O_1632,N_14328,N_14323);
nor UO_1633 (O_1633,N_14622,N_14875);
xnor UO_1634 (O_1634,N_14522,N_14274);
xnor UO_1635 (O_1635,N_14438,N_14494);
or UO_1636 (O_1636,N_14672,N_14349);
or UO_1637 (O_1637,N_14780,N_14441);
nand UO_1638 (O_1638,N_14663,N_14364);
nor UO_1639 (O_1639,N_14465,N_14828);
nor UO_1640 (O_1640,N_14690,N_14640);
nor UO_1641 (O_1641,N_14996,N_14814);
xor UO_1642 (O_1642,N_14629,N_14587);
xor UO_1643 (O_1643,N_14521,N_14446);
nor UO_1644 (O_1644,N_14792,N_14685);
xnor UO_1645 (O_1645,N_14525,N_14359);
or UO_1646 (O_1646,N_14910,N_14287);
or UO_1647 (O_1647,N_14592,N_14337);
xor UO_1648 (O_1648,N_14972,N_14879);
and UO_1649 (O_1649,N_14697,N_14644);
or UO_1650 (O_1650,N_14271,N_14407);
nand UO_1651 (O_1651,N_14484,N_14889);
nand UO_1652 (O_1652,N_14873,N_14602);
or UO_1653 (O_1653,N_14487,N_14255);
xor UO_1654 (O_1654,N_14870,N_14352);
nand UO_1655 (O_1655,N_14371,N_14869);
or UO_1656 (O_1656,N_14336,N_14596);
nand UO_1657 (O_1657,N_14728,N_14775);
xnor UO_1658 (O_1658,N_14920,N_14748);
xnor UO_1659 (O_1659,N_14252,N_14618);
nand UO_1660 (O_1660,N_14963,N_14281);
and UO_1661 (O_1661,N_14751,N_14324);
and UO_1662 (O_1662,N_14594,N_14775);
nor UO_1663 (O_1663,N_14423,N_14898);
or UO_1664 (O_1664,N_14594,N_14370);
nor UO_1665 (O_1665,N_14614,N_14308);
nand UO_1666 (O_1666,N_14937,N_14835);
nand UO_1667 (O_1667,N_14345,N_14671);
or UO_1668 (O_1668,N_14317,N_14508);
or UO_1669 (O_1669,N_14630,N_14418);
nor UO_1670 (O_1670,N_14779,N_14842);
nand UO_1671 (O_1671,N_14725,N_14265);
nand UO_1672 (O_1672,N_14693,N_14618);
nor UO_1673 (O_1673,N_14307,N_14824);
nand UO_1674 (O_1674,N_14772,N_14866);
xor UO_1675 (O_1675,N_14674,N_14412);
and UO_1676 (O_1676,N_14691,N_14274);
or UO_1677 (O_1677,N_14383,N_14753);
nor UO_1678 (O_1678,N_14527,N_14524);
and UO_1679 (O_1679,N_14709,N_14602);
xor UO_1680 (O_1680,N_14262,N_14827);
or UO_1681 (O_1681,N_14870,N_14300);
xnor UO_1682 (O_1682,N_14501,N_14325);
nor UO_1683 (O_1683,N_14459,N_14353);
nand UO_1684 (O_1684,N_14660,N_14850);
and UO_1685 (O_1685,N_14483,N_14336);
nand UO_1686 (O_1686,N_14661,N_14725);
or UO_1687 (O_1687,N_14553,N_14396);
and UO_1688 (O_1688,N_14461,N_14990);
xor UO_1689 (O_1689,N_14767,N_14726);
xnor UO_1690 (O_1690,N_14346,N_14890);
xnor UO_1691 (O_1691,N_14996,N_14283);
xnor UO_1692 (O_1692,N_14301,N_14970);
xor UO_1693 (O_1693,N_14655,N_14587);
nor UO_1694 (O_1694,N_14253,N_14538);
and UO_1695 (O_1695,N_14843,N_14430);
or UO_1696 (O_1696,N_14582,N_14497);
xnor UO_1697 (O_1697,N_14314,N_14739);
and UO_1698 (O_1698,N_14875,N_14499);
or UO_1699 (O_1699,N_14985,N_14833);
or UO_1700 (O_1700,N_14762,N_14282);
and UO_1701 (O_1701,N_14459,N_14612);
or UO_1702 (O_1702,N_14314,N_14963);
xor UO_1703 (O_1703,N_14327,N_14999);
nand UO_1704 (O_1704,N_14963,N_14928);
nand UO_1705 (O_1705,N_14260,N_14952);
or UO_1706 (O_1706,N_14629,N_14442);
or UO_1707 (O_1707,N_14277,N_14694);
nor UO_1708 (O_1708,N_14751,N_14504);
xor UO_1709 (O_1709,N_14943,N_14989);
xor UO_1710 (O_1710,N_14405,N_14393);
nor UO_1711 (O_1711,N_14995,N_14455);
nor UO_1712 (O_1712,N_14860,N_14268);
and UO_1713 (O_1713,N_14740,N_14858);
xor UO_1714 (O_1714,N_14724,N_14985);
or UO_1715 (O_1715,N_14957,N_14929);
nand UO_1716 (O_1716,N_14327,N_14548);
and UO_1717 (O_1717,N_14601,N_14807);
or UO_1718 (O_1718,N_14693,N_14701);
xnor UO_1719 (O_1719,N_14742,N_14303);
nor UO_1720 (O_1720,N_14929,N_14347);
xnor UO_1721 (O_1721,N_14833,N_14263);
or UO_1722 (O_1722,N_14913,N_14406);
nand UO_1723 (O_1723,N_14824,N_14896);
or UO_1724 (O_1724,N_14664,N_14928);
xor UO_1725 (O_1725,N_14717,N_14267);
and UO_1726 (O_1726,N_14681,N_14586);
and UO_1727 (O_1727,N_14309,N_14680);
xnor UO_1728 (O_1728,N_14899,N_14252);
nand UO_1729 (O_1729,N_14443,N_14543);
nand UO_1730 (O_1730,N_14387,N_14704);
xnor UO_1731 (O_1731,N_14469,N_14408);
xor UO_1732 (O_1732,N_14455,N_14816);
xnor UO_1733 (O_1733,N_14637,N_14781);
nor UO_1734 (O_1734,N_14685,N_14288);
or UO_1735 (O_1735,N_14543,N_14465);
and UO_1736 (O_1736,N_14729,N_14958);
and UO_1737 (O_1737,N_14332,N_14364);
xor UO_1738 (O_1738,N_14477,N_14610);
nor UO_1739 (O_1739,N_14485,N_14936);
or UO_1740 (O_1740,N_14619,N_14891);
nand UO_1741 (O_1741,N_14510,N_14670);
and UO_1742 (O_1742,N_14331,N_14676);
nor UO_1743 (O_1743,N_14507,N_14995);
nand UO_1744 (O_1744,N_14380,N_14962);
and UO_1745 (O_1745,N_14624,N_14773);
xor UO_1746 (O_1746,N_14785,N_14258);
and UO_1747 (O_1747,N_14795,N_14638);
nand UO_1748 (O_1748,N_14742,N_14648);
and UO_1749 (O_1749,N_14260,N_14366);
or UO_1750 (O_1750,N_14366,N_14372);
and UO_1751 (O_1751,N_14284,N_14467);
or UO_1752 (O_1752,N_14442,N_14604);
xnor UO_1753 (O_1753,N_14685,N_14250);
nand UO_1754 (O_1754,N_14464,N_14589);
and UO_1755 (O_1755,N_14405,N_14374);
xor UO_1756 (O_1756,N_14486,N_14538);
nor UO_1757 (O_1757,N_14820,N_14733);
xnor UO_1758 (O_1758,N_14608,N_14613);
or UO_1759 (O_1759,N_14546,N_14607);
nor UO_1760 (O_1760,N_14925,N_14800);
and UO_1761 (O_1761,N_14291,N_14503);
nor UO_1762 (O_1762,N_14700,N_14252);
xor UO_1763 (O_1763,N_14812,N_14473);
or UO_1764 (O_1764,N_14439,N_14695);
nand UO_1765 (O_1765,N_14590,N_14495);
and UO_1766 (O_1766,N_14314,N_14879);
nand UO_1767 (O_1767,N_14897,N_14675);
nor UO_1768 (O_1768,N_14557,N_14351);
xor UO_1769 (O_1769,N_14334,N_14782);
xor UO_1770 (O_1770,N_14888,N_14275);
or UO_1771 (O_1771,N_14506,N_14349);
nor UO_1772 (O_1772,N_14498,N_14774);
or UO_1773 (O_1773,N_14275,N_14778);
nand UO_1774 (O_1774,N_14592,N_14585);
xor UO_1775 (O_1775,N_14653,N_14875);
nor UO_1776 (O_1776,N_14678,N_14688);
xnor UO_1777 (O_1777,N_14647,N_14460);
nor UO_1778 (O_1778,N_14528,N_14775);
or UO_1779 (O_1779,N_14410,N_14746);
and UO_1780 (O_1780,N_14408,N_14735);
or UO_1781 (O_1781,N_14587,N_14498);
or UO_1782 (O_1782,N_14340,N_14544);
or UO_1783 (O_1783,N_14478,N_14847);
or UO_1784 (O_1784,N_14306,N_14711);
and UO_1785 (O_1785,N_14458,N_14978);
nor UO_1786 (O_1786,N_14583,N_14984);
and UO_1787 (O_1787,N_14595,N_14312);
xor UO_1788 (O_1788,N_14566,N_14466);
nor UO_1789 (O_1789,N_14666,N_14756);
and UO_1790 (O_1790,N_14332,N_14998);
and UO_1791 (O_1791,N_14578,N_14600);
nor UO_1792 (O_1792,N_14844,N_14740);
nand UO_1793 (O_1793,N_14728,N_14644);
and UO_1794 (O_1794,N_14579,N_14345);
or UO_1795 (O_1795,N_14527,N_14440);
nor UO_1796 (O_1796,N_14312,N_14579);
and UO_1797 (O_1797,N_14399,N_14690);
or UO_1798 (O_1798,N_14288,N_14461);
and UO_1799 (O_1799,N_14647,N_14596);
and UO_1800 (O_1800,N_14327,N_14394);
nor UO_1801 (O_1801,N_14464,N_14340);
nand UO_1802 (O_1802,N_14820,N_14934);
nor UO_1803 (O_1803,N_14922,N_14999);
or UO_1804 (O_1804,N_14654,N_14657);
nand UO_1805 (O_1805,N_14600,N_14447);
xor UO_1806 (O_1806,N_14700,N_14551);
or UO_1807 (O_1807,N_14808,N_14759);
and UO_1808 (O_1808,N_14731,N_14709);
nand UO_1809 (O_1809,N_14601,N_14720);
nand UO_1810 (O_1810,N_14839,N_14307);
and UO_1811 (O_1811,N_14986,N_14916);
xor UO_1812 (O_1812,N_14366,N_14993);
nor UO_1813 (O_1813,N_14561,N_14707);
nor UO_1814 (O_1814,N_14348,N_14286);
xor UO_1815 (O_1815,N_14311,N_14967);
and UO_1816 (O_1816,N_14499,N_14519);
xnor UO_1817 (O_1817,N_14721,N_14818);
nor UO_1818 (O_1818,N_14714,N_14536);
xnor UO_1819 (O_1819,N_14790,N_14648);
nor UO_1820 (O_1820,N_14293,N_14447);
xnor UO_1821 (O_1821,N_14628,N_14542);
xnor UO_1822 (O_1822,N_14979,N_14526);
nor UO_1823 (O_1823,N_14441,N_14926);
nor UO_1824 (O_1824,N_14770,N_14896);
xor UO_1825 (O_1825,N_14696,N_14982);
xor UO_1826 (O_1826,N_14266,N_14646);
and UO_1827 (O_1827,N_14655,N_14943);
or UO_1828 (O_1828,N_14816,N_14826);
and UO_1829 (O_1829,N_14655,N_14782);
xnor UO_1830 (O_1830,N_14720,N_14269);
and UO_1831 (O_1831,N_14969,N_14341);
nand UO_1832 (O_1832,N_14543,N_14818);
nand UO_1833 (O_1833,N_14593,N_14737);
nand UO_1834 (O_1834,N_14270,N_14324);
nor UO_1835 (O_1835,N_14785,N_14468);
and UO_1836 (O_1836,N_14858,N_14890);
nand UO_1837 (O_1837,N_14445,N_14261);
xor UO_1838 (O_1838,N_14517,N_14893);
xor UO_1839 (O_1839,N_14386,N_14412);
nor UO_1840 (O_1840,N_14927,N_14393);
or UO_1841 (O_1841,N_14798,N_14476);
xnor UO_1842 (O_1842,N_14947,N_14429);
and UO_1843 (O_1843,N_14392,N_14341);
xor UO_1844 (O_1844,N_14933,N_14737);
nor UO_1845 (O_1845,N_14561,N_14288);
xor UO_1846 (O_1846,N_14901,N_14380);
and UO_1847 (O_1847,N_14543,N_14283);
or UO_1848 (O_1848,N_14349,N_14802);
nor UO_1849 (O_1849,N_14462,N_14512);
nor UO_1850 (O_1850,N_14286,N_14615);
xor UO_1851 (O_1851,N_14769,N_14990);
and UO_1852 (O_1852,N_14455,N_14443);
xnor UO_1853 (O_1853,N_14997,N_14681);
and UO_1854 (O_1854,N_14722,N_14457);
nand UO_1855 (O_1855,N_14559,N_14969);
nand UO_1856 (O_1856,N_14416,N_14435);
xor UO_1857 (O_1857,N_14738,N_14826);
and UO_1858 (O_1858,N_14374,N_14939);
xor UO_1859 (O_1859,N_14395,N_14477);
or UO_1860 (O_1860,N_14434,N_14901);
or UO_1861 (O_1861,N_14785,N_14250);
or UO_1862 (O_1862,N_14602,N_14733);
nor UO_1863 (O_1863,N_14477,N_14846);
and UO_1864 (O_1864,N_14587,N_14934);
nand UO_1865 (O_1865,N_14536,N_14638);
or UO_1866 (O_1866,N_14721,N_14252);
and UO_1867 (O_1867,N_14903,N_14816);
or UO_1868 (O_1868,N_14447,N_14836);
or UO_1869 (O_1869,N_14440,N_14870);
and UO_1870 (O_1870,N_14761,N_14585);
xor UO_1871 (O_1871,N_14992,N_14579);
or UO_1872 (O_1872,N_14557,N_14802);
xnor UO_1873 (O_1873,N_14979,N_14814);
xor UO_1874 (O_1874,N_14910,N_14581);
or UO_1875 (O_1875,N_14744,N_14523);
or UO_1876 (O_1876,N_14955,N_14733);
nor UO_1877 (O_1877,N_14442,N_14452);
or UO_1878 (O_1878,N_14574,N_14878);
and UO_1879 (O_1879,N_14364,N_14963);
nand UO_1880 (O_1880,N_14971,N_14994);
nor UO_1881 (O_1881,N_14364,N_14366);
and UO_1882 (O_1882,N_14625,N_14430);
or UO_1883 (O_1883,N_14584,N_14841);
nand UO_1884 (O_1884,N_14508,N_14418);
nand UO_1885 (O_1885,N_14786,N_14469);
or UO_1886 (O_1886,N_14681,N_14289);
and UO_1887 (O_1887,N_14980,N_14731);
nand UO_1888 (O_1888,N_14859,N_14270);
nand UO_1889 (O_1889,N_14596,N_14620);
nand UO_1890 (O_1890,N_14822,N_14434);
or UO_1891 (O_1891,N_14266,N_14653);
nand UO_1892 (O_1892,N_14996,N_14735);
nor UO_1893 (O_1893,N_14330,N_14960);
nand UO_1894 (O_1894,N_14789,N_14694);
xnor UO_1895 (O_1895,N_14443,N_14879);
nor UO_1896 (O_1896,N_14609,N_14781);
xnor UO_1897 (O_1897,N_14870,N_14691);
xor UO_1898 (O_1898,N_14513,N_14467);
nor UO_1899 (O_1899,N_14946,N_14847);
nor UO_1900 (O_1900,N_14338,N_14894);
nor UO_1901 (O_1901,N_14747,N_14576);
nor UO_1902 (O_1902,N_14654,N_14924);
or UO_1903 (O_1903,N_14729,N_14754);
nand UO_1904 (O_1904,N_14684,N_14666);
nor UO_1905 (O_1905,N_14366,N_14916);
nor UO_1906 (O_1906,N_14521,N_14609);
nor UO_1907 (O_1907,N_14396,N_14787);
nor UO_1908 (O_1908,N_14579,N_14406);
nor UO_1909 (O_1909,N_14877,N_14365);
or UO_1910 (O_1910,N_14750,N_14978);
or UO_1911 (O_1911,N_14321,N_14810);
or UO_1912 (O_1912,N_14462,N_14421);
nor UO_1913 (O_1913,N_14461,N_14473);
nor UO_1914 (O_1914,N_14655,N_14920);
nor UO_1915 (O_1915,N_14528,N_14903);
xor UO_1916 (O_1916,N_14796,N_14553);
nor UO_1917 (O_1917,N_14590,N_14605);
xor UO_1918 (O_1918,N_14868,N_14551);
and UO_1919 (O_1919,N_14442,N_14505);
and UO_1920 (O_1920,N_14571,N_14696);
or UO_1921 (O_1921,N_14664,N_14808);
nand UO_1922 (O_1922,N_14636,N_14617);
nor UO_1923 (O_1923,N_14388,N_14550);
or UO_1924 (O_1924,N_14637,N_14354);
xor UO_1925 (O_1925,N_14950,N_14935);
and UO_1926 (O_1926,N_14799,N_14311);
xor UO_1927 (O_1927,N_14491,N_14559);
or UO_1928 (O_1928,N_14498,N_14760);
or UO_1929 (O_1929,N_14721,N_14348);
xnor UO_1930 (O_1930,N_14527,N_14380);
nand UO_1931 (O_1931,N_14842,N_14864);
and UO_1932 (O_1932,N_14917,N_14798);
xor UO_1933 (O_1933,N_14614,N_14549);
or UO_1934 (O_1934,N_14972,N_14412);
or UO_1935 (O_1935,N_14462,N_14802);
or UO_1936 (O_1936,N_14766,N_14693);
xor UO_1937 (O_1937,N_14832,N_14261);
xor UO_1938 (O_1938,N_14568,N_14722);
nand UO_1939 (O_1939,N_14638,N_14356);
nor UO_1940 (O_1940,N_14969,N_14711);
nor UO_1941 (O_1941,N_14850,N_14959);
or UO_1942 (O_1942,N_14352,N_14454);
nand UO_1943 (O_1943,N_14805,N_14534);
xnor UO_1944 (O_1944,N_14331,N_14833);
nand UO_1945 (O_1945,N_14292,N_14931);
and UO_1946 (O_1946,N_14555,N_14891);
and UO_1947 (O_1947,N_14747,N_14891);
and UO_1948 (O_1948,N_14984,N_14886);
nand UO_1949 (O_1949,N_14866,N_14766);
and UO_1950 (O_1950,N_14590,N_14530);
nand UO_1951 (O_1951,N_14367,N_14620);
or UO_1952 (O_1952,N_14895,N_14354);
or UO_1953 (O_1953,N_14707,N_14803);
or UO_1954 (O_1954,N_14744,N_14254);
or UO_1955 (O_1955,N_14532,N_14619);
nor UO_1956 (O_1956,N_14400,N_14711);
xor UO_1957 (O_1957,N_14535,N_14934);
or UO_1958 (O_1958,N_14912,N_14826);
xor UO_1959 (O_1959,N_14474,N_14513);
xor UO_1960 (O_1960,N_14889,N_14362);
and UO_1961 (O_1961,N_14571,N_14388);
xor UO_1962 (O_1962,N_14760,N_14835);
nor UO_1963 (O_1963,N_14619,N_14731);
nand UO_1964 (O_1964,N_14999,N_14759);
or UO_1965 (O_1965,N_14617,N_14619);
nor UO_1966 (O_1966,N_14877,N_14767);
or UO_1967 (O_1967,N_14332,N_14287);
xnor UO_1968 (O_1968,N_14776,N_14902);
nand UO_1969 (O_1969,N_14975,N_14700);
or UO_1970 (O_1970,N_14252,N_14349);
xnor UO_1971 (O_1971,N_14722,N_14439);
xor UO_1972 (O_1972,N_14893,N_14311);
and UO_1973 (O_1973,N_14275,N_14307);
nand UO_1974 (O_1974,N_14415,N_14665);
xor UO_1975 (O_1975,N_14488,N_14855);
xor UO_1976 (O_1976,N_14964,N_14363);
or UO_1977 (O_1977,N_14344,N_14555);
nand UO_1978 (O_1978,N_14497,N_14673);
xnor UO_1979 (O_1979,N_14522,N_14790);
nor UO_1980 (O_1980,N_14954,N_14951);
nand UO_1981 (O_1981,N_14498,N_14903);
xnor UO_1982 (O_1982,N_14343,N_14839);
nor UO_1983 (O_1983,N_14499,N_14357);
or UO_1984 (O_1984,N_14525,N_14351);
xor UO_1985 (O_1985,N_14675,N_14436);
xor UO_1986 (O_1986,N_14279,N_14491);
nand UO_1987 (O_1987,N_14316,N_14730);
and UO_1988 (O_1988,N_14693,N_14316);
xor UO_1989 (O_1989,N_14834,N_14528);
nand UO_1990 (O_1990,N_14685,N_14483);
or UO_1991 (O_1991,N_14339,N_14833);
xnor UO_1992 (O_1992,N_14479,N_14767);
or UO_1993 (O_1993,N_14909,N_14987);
or UO_1994 (O_1994,N_14259,N_14817);
nor UO_1995 (O_1995,N_14411,N_14975);
or UO_1996 (O_1996,N_14593,N_14351);
nand UO_1997 (O_1997,N_14660,N_14918);
nor UO_1998 (O_1998,N_14253,N_14659);
and UO_1999 (O_1999,N_14419,N_14687);
endmodule