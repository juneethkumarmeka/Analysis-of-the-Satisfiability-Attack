module basic_2000_20000_2500_5_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1279,In_505);
and U1 (N_1,In_1717,In_533);
nor U2 (N_2,In_419,In_1915);
and U3 (N_3,In_23,In_887);
xor U4 (N_4,In_34,In_1436);
xor U5 (N_5,In_640,In_1596);
xnor U6 (N_6,In_1158,In_649);
nor U7 (N_7,In_1002,In_607);
or U8 (N_8,In_216,In_1393);
nand U9 (N_9,In_1300,In_1824);
nor U10 (N_10,In_827,In_790);
and U11 (N_11,In_412,In_314);
nor U12 (N_12,In_1130,In_58);
nor U13 (N_13,In_681,In_1573);
or U14 (N_14,In_331,In_896);
and U15 (N_15,In_266,In_1327);
nand U16 (N_16,In_1498,In_1391);
and U17 (N_17,In_1024,In_1248);
xnor U18 (N_18,In_1359,In_694);
and U19 (N_19,In_89,In_559);
nand U20 (N_20,In_56,In_1131);
nor U21 (N_21,In_853,In_1445);
nor U22 (N_22,In_516,In_1291);
nand U23 (N_23,In_162,In_1946);
nor U24 (N_24,In_252,In_1532);
xnor U25 (N_25,In_1956,In_1213);
nand U26 (N_26,In_1141,In_1677);
xor U27 (N_27,In_1053,In_1030);
nand U28 (N_28,In_821,In_1838);
and U29 (N_29,In_203,In_699);
and U30 (N_30,In_1776,In_297);
or U31 (N_31,In_95,In_1608);
nor U32 (N_32,In_91,In_1365);
nor U33 (N_33,In_1404,In_1802);
or U34 (N_34,In_1278,In_1952);
nand U35 (N_35,In_1982,In_1834);
or U36 (N_36,In_974,In_1363);
or U37 (N_37,In_679,In_1550);
xnor U38 (N_38,In_1620,In_723);
nand U39 (N_39,In_773,In_213);
and U40 (N_40,In_918,In_447);
and U41 (N_41,In_1925,In_1991);
or U42 (N_42,In_1678,In_262);
and U43 (N_43,In_995,In_595);
or U44 (N_44,In_772,In_1630);
nor U45 (N_45,In_124,In_770);
and U46 (N_46,In_558,In_459);
nor U47 (N_47,In_1521,In_1716);
and U48 (N_48,In_1818,In_479);
or U49 (N_49,In_1435,In_1453);
nand U50 (N_50,In_1253,In_1829);
and U51 (N_51,In_917,In_734);
nor U52 (N_52,In_1633,In_1562);
nand U53 (N_53,In_754,In_1303);
and U54 (N_54,In_486,In_1176);
or U55 (N_55,In_1961,In_1013);
and U56 (N_56,In_1512,In_243);
or U57 (N_57,In_219,In_1302);
nand U58 (N_58,In_1627,In_1821);
or U59 (N_59,In_635,In_322);
nand U60 (N_60,In_1696,In_1509);
nand U61 (N_61,In_633,In_1665);
or U62 (N_62,In_903,In_687);
or U63 (N_63,In_902,In_1764);
and U64 (N_64,In_490,In_1746);
nand U65 (N_65,In_1661,In_296);
nand U66 (N_66,In_581,In_1820);
nand U67 (N_67,In_254,In_1258);
nor U68 (N_68,In_1273,In_820);
xor U69 (N_69,In_1595,In_66);
nand U70 (N_70,In_183,In_1170);
or U71 (N_71,In_1421,In_863);
xnor U72 (N_72,In_404,In_340);
xor U73 (N_73,In_1728,In_550);
nand U74 (N_74,In_763,In_776);
or U75 (N_75,In_1179,In_920);
nor U76 (N_76,In_1823,In_192);
xnor U77 (N_77,In_1756,In_1115);
xnor U78 (N_78,In_1741,In_532);
or U79 (N_79,In_703,In_40);
nor U80 (N_80,In_1180,In_1038);
nor U81 (N_81,In_562,In_286);
xor U82 (N_82,In_1760,In_1736);
or U83 (N_83,In_1351,In_1969);
nand U84 (N_84,In_281,In_657);
nand U85 (N_85,In_292,In_55);
and U86 (N_86,In_242,In_1408);
nor U87 (N_87,In_1772,In_28);
or U88 (N_88,In_1744,In_232);
nor U89 (N_89,In_1243,In_1223);
xor U90 (N_90,In_85,In_1767);
or U91 (N_91,In_1538,In_816);
xor U92 (N_92,In_1047,In_676);
nor U93 (N_93,In_1462,In_1916);
and U94 (N_94,In_1191,In_1774);
nor U95 (N_95,In_1282,In_453);
nand U96 (N_96,In_1255,In_950);
nor U97 (N_97,In_1718,In_466);
and U98 (N_98,In_1088,In_991);
nand U99 (N_99,In_1528,In_919);
or U100 (N_100,In_425,In_1603);
nor U101 (N_101,In_1800,In_1315);
and U102 (N_102,In_683,In_1794);
xnor U103 (N_103,In_1139,In_1529);
xor U104 (N_104,In_1742,In_193);
or U105 (N_105,In_282,In_1655);
nand U106 (N_106,In_1073,In_1947);
xor U107 (N_107,In_938,In_1670);
or U108 (N_108,In_874,In_915);
or U109 (N_109,In_573,In_1567);
nand U110 (N_110,In_18,In_1936);
nand U111 (N_111,In_1753,In_717);
and U112 (N_112,In_1428,In_599);
and U113 (N_113,In_1525,In_1890);
xor U114 (N_114,In_1578,In_1340);
nand U115 (N_115,In_546,In_794);
nor U116 (N_116,In_619,In_841);
nor U117 (N_117,In_1322,In_988);
and U118 (N_118,In_985,In_336);
and U119 (N_119,In_1241,In_1084);
nand U120 (N_120,In_1975,In_103);
xor U121 (N_121,In_1960,In_906);
nand U122 (N_122,In_1636,In_202);
nor U123 (N_123,In_1726,In_1334);
nor U124 (N_124,In_1685,In_366);
xnor U125 (N_125,In_1424,In_872);
nand U126 (N_126,In_1389,In_571);
nor U127 (N_127,In_527,In_1967);
and U128 (N_128,In_87,In_365);
nor U129 (N_129,In_48,In_1246);
xnor U130 (N_130,In_467,In_442);
and U131 (N_131,In_1054,In_1125);
nand U132 (N_132,In_511,In_1019);
nor U133 (N_133,In_200,In_739);
nand U134 (N_134,In_628,In_38);
or U135 (N_135,In_1264,In_519);
and U136 (N_136,In_39,In_1866);
nand U137 (N_137,In_730,In_1527);
and U138 (N_138,In_960,In_1508);
xor U139 (N_139,In_310,In_1150);
or U140 (N_140,In_1092,In_1239);
nand U141 (N_141,In_492,In_673);
xor U142 (N_142,In_777,In_413);
and U143 (N_143,In_1537,In_1720);
nor U144 (N_144,In_343,In_1924);
xor U145 (N_145,In_1839,In_1474);
nand U146 (N_146,In_1863,In_1667);
nand U147 (N_147,In_1173,In_1730);
and U148 (N_148,In_789,In_1362);
and U149 (N_149,In_1690,In_708);
nand U150 (N_150,In_588,In_871);
xnor U151 (N_151,In_1888,In_1051);
nand U152 (N_152,In_450,In_346);
or U153 (N_153,In_1260,In_733);
and U154 (N_154,In_62,In_1872);
and U155 (N_155,In_823,In_1556);
nand U156 (N_156,In_1122,In_1461);
or U157 (N_157,In_1162,In_1154);
xnor U158 (N_158,In_631,In_160);
or U159 (N_159,In_877,In_291);
and U160 (N_160,In_1657,In_568);
or U161 (N_161,In_1885,In_1438);
or U162 (N_162,In_1601,In_614);
nor U163 (N_163,In_1681,In_484);
or U164 (N_164,In_1459,In_1989);
and U165 (N_165,In_370,In_1713);
or U166 (N_166,In_940,In_376);
and U167 (N_167,In_120,In_197);
or U168 (N_168,In_1877,In_181);
nor U169 (N_169,In_256,In_1927);
xnor U170 (N_170,In_510,In_131);
xor U171 (N_171,In_1894,In_1926);
xnor U172 (N_172,In_133,In_755);
nand U173 (N_173,In_1647,In_438);
xnor U174 (N_174,In_1933,In_1939);
nand U175 (N_175,In_441,In_552);
xor U176 (N_176,In_1352,In_861);
nor U177 (N_177,In_651,In_199);
or U178 (N_178,In_826,In_566);
nor U179 (N_179,In_500,In_1049);
nand U180 (N_180,In_353,In_639);
or U181 (N_181,In_1524,In_1400);
or U182 (N_182,In_383,In_899);
nand U183 (N_183,In_1990,In_1324);
or U184 (N_184,In_241,In_774);
xor U185 (N_185,In_721,In_1074);
or U186 (N_186,In_1777,In_260);
nand U187 (N_187,In_1920,In_692);
or U188 (N_188,In_767,In_1797);
nor U189 (N_189,In_585,In_361);
xor U190 (N_190,In_1367,In_107);
nand U191 (N_191,In_1914,In_1022);
and U192 (N_192,In_410,In_1177);
xnor U193 (N_193,In_72,In_1199);
or U194 (N_194,In_1228,In_1395);
nor U195 (N_195,In_185,In_1999);
and U196 (N_196,In_76,In_32);
or U197 (N_197,In_1549,In_956);
xor U198 (N_198,In_650,In_1068);
or U199 (N_199,In_1923,In_443);
xnor U200 (N_200,In_518,In_1148);
xnor U201 (N_201,In_10,In_688);
nor U202 (N_202,In_892,In_1867);
nand U203 (N_203,In_1370,In_1574);
and U204 (N_204,In_1114,In_667);
nor U205 (N_205,In_1195,In_1959);
and U206 (N_206,In_210,In_1346);
nand U207 (N_207,In_436,In_1515);
nor U208 (N_208,In_1862,In_1345);
or U209 (N_209,In_168,In_283);
nor U210 (N_210,In_1161,In_724);
and U211 (N_211,In_1376,In_1789);
nor U212 (N_212,In_464,In_358);
xor U213 (N_213,In_525,In_1500);
nor U214 (N_214,In_304,In_476);
and U215 (N_215,In_1166,In_944);
or U216 (N_216,In_886,In_775);
nor U217 (N_217,In_801,In_324);
nor U218 (N_218,In_71,In_967);
nor U219 (N_219,In_587,In_1263);
or U220 (N_220,In_839,In_1472);
nor U221 (N_221,In_803,In_1714);
or U222 (N_222,In_371,In_1479);
nor U223 (N_223,In_514,In_380);
or U224 (N_224,In_257,In_1548);
or U225 (N_225,In_395,In_482);
or U226 (N_226,In_1725,In_251);
nor U227 (N_227,In_1640,In_608);
nand U228 (N_228,In_287,In_1251);
and U229 (N_229,In_24,In_1676);
xnor U230 (N_230,In_136,In_1105);
nor U231 (N_231,In_646,In_98);
nor U232 (N_232,In_992,In_1159);
or U233 (N_233,In_1869,In_384);
nand U234 (N_234,In_350,In_1897);
xnor U235 (N_235,In_207,In_972);
xor U236 (N_236,In_1828,In_642);
and U237 (N_237,In_970,In_1378);
nand U238 (N_238,In_196,In_272);
or U239 (N_239,In_1443,In_311);
xnor U240 (N_240,In_1257,In_362);
nor U241 (N_241,In_134,In_109);
nand U242 (N_242,In_147,In_223);
nand U243 (N_243,In_644,In_420);
nor U244 (N_244,In_700,In_1165);
and U245 (N_245,In_1672,In_893);
nand U246 (N_246,In_1427,In_165);
nand U247 (N_247,In_578,In_1819);
nor U248 (N_248,In_1503,In_746);
or U249 (N_249,In_1795,In_1413);
nor U250 (N_250,In_1792,In_1788);
or U251 (N_251,In_1942,In_1856);
nand U252 (N_252,In_1487,In_1910);
or U253 (N_253,In_549,In_1859);
xor U254 (N_254,In_1769,In_8);
and U255 (N_255,In_1481,In_1875);
xnor U256 (N_256,In_153,In_1850);
and U257 (N_257,In_1368,In_655);
and U258 (N_258,In_1467,In_1913);
or U259 (N_259,In_1695,In_69);
nand U260 (N_260,In_1851,In_1106);
or U261 (N_261,In_689,In_130);
or U262 (N_262,In_851,In_212);
or U263 (N_263,In_1815,In_318);
nand U264 (N_264,In_285,In_1575);
and U265 (N_265,In_1662,In_1360);
or U266 (N_266,In_1204,In_811);
nand U267 (N_267,In_647,In_1848);
and U268 (N_268,In_706,In_1476);
or U269 (N_269,In_1379,In_1041);
nand U270 (N_270,In_1212,In_271);
nand U271 (N_271,In_537,In_885);
or U272 (N_272,In_1766,In_378);
nor U273 (N_273,In_515,In_1009);
xnor U274 (N_274,In_480,In_1171);
nor U275 (N_275,In_1809,In_1634);
and U276 (N_276,In_570,In_865);
nor U277 (N_277,In_1194,In_1683);
or U278 (N_278,In_1921,In_855);
and U279 (N_279,In_665,In_491);
xor U280 (N_280,In_809,In_854);
xor U281 (N_281,In_1722,In_1617);
and U282 (N_282,In_1120,In_907);
or U283 (N_283,In_1941,In_1135);
nor U284 (N_284,In_526,In_959);
and U285 (N_285,In_799,In_173);
and U286 (N_286,In_1733,In_215);
nor U287 (N_287,In_1289,In_586);
or U288 (N_288,In_1895,In_1691);
nand U289 (N_289,In_668,In_154);
xor U290 (N_290,In_830,In_387);
xnor U291 (N_291,In_53,In_1584);
nor U292 (N_292,In_806,In_461);
xor U293 (N_293,In_1387,In_392);
and U294 (N_294,In_1687,In_979);
xor U295 (N_295,In_836,In_513);
or U296 (N_296,In_81,In_315);
nor U297 (N_297,In_1423,In_1025);
or U298 (N_298,In_9,In_1896);
and U299 (N_299,In_334,In_1099);
or U300 (N_300,In_463,In_1882);
or U301 (N_301,In_1905,In_389);
nor U302 (N_302,In_188,In_1048);
nand U303 (N_303,In_309,In_895);
and U304 (N_304,In_954,In_849);
nand U305 (N_305,In_337,In_1534);
nand U306 (N_306,In_0,In_1645);
xor U307 (N_307,In_374,In_764);
nor U308 (N_308,In_422,In_1276);
or U309 (N_309,In_1621,In_101);
nand U310 (N_310,In_696,In_1321);
nor U311 (N_311,In_1197,In_911);
and U312 (N_312,In_320,In_49);
nand U313 (N_313,In_1401,In_548);
nor U314 (N_314,In_1259,In_1310);
or U315 (N_315,In_295,In_1232);
and U316 (N_316,In_1734,In_391);
and U317 (N_317,In_544,In_267);
nand U318 (N_318,In_489,In_1477);
nor U319 (N_319,In_1101,In_971);
xor U320 (N_320,In_308,In_1689);
or U321 (N_321,In_127,In_345);
nand U322 (N_322,In_517,In_837);
and U323 (N_323,In_1210,In_198);
and U324 (N_324,In_1016,In_1307);
or U325 (N_325,In_278,In_729);
nor U326 (N_326,In_329,In_1786);
nand U327 (N_327,In_1565,In_1268);
and U328 (N_328,In_1996,In_728);
nand U329 (N_329,In_1485,In_225);
xor U330 (N_330,In_140,In_142);
and U331 (N_331,In_44,In_1205);
and U332 (N_332,In_1704,In_1441);
nand U333 (N_333,In_1446,In_669);
and U334 (N_334,In_1870,In_230);
nand U335 (N_335,In_67,In_132);
and U336 (N_336,In_355,In_590);
and U337 (N_337,In_235,In_424);
xor U338 (N_338,In_110,In_1117);
or U339 (N_339,In_1412,In_1275);
and U340 (N_340,In_645,In_701);
or U341 (N_341,In_1032,In_1847);
nand U342 (N_342,In_744,In_743);
xor U343 (N_343,In_75,In_888);
or U344 (N_344,In_1316,In_949);
or U345 (N_345,In_189,In_1182);
nand U346 (N_346,In_236,In_786);
xor U347 (N_347,In_1514,In_713);
xnor U348 (N_348,In_434,In_1660);
and U349 (N_349,In_1699,In_156);
xnor U350 (N_350,In_298,In_35);
xnor U351 (N_351,In_509,In_3);
and U352 (N_352,In_1879,In_521);
and U353 (N_353,In_1825,In_1118);
nor U354 (N_354,In_661,In_1229);
nand U355 (N_355,In_167,In_280);
or U356 (N_356,In_686,In_1187);
or U357 (N_357,In_125,In_1271);
or U358 (N_358,In_916,In_1974);
and U359 (N_359,In_1891,In_625);
xor U360 (N_360,In_1478,In_555);
and U361 (N_361,In_884,In_363);
nand U362 (N_362,In_209,In_469);
xnor U363 (N_363,In_1035,In_752);
nand U364 (N_364,In_1039,In_714);
and U365 (N_365,In_576,In_575);
and U366 (N_366,In_1664,In_1331);
nand U367 (N_367,In_1526,In_1849);
and U368 (N_368,In_1325,In_265);
or U369 (N_369,In_1308,In_65);
nor U370 (N_370,In_1604,In_1277);
or U371 (N_371,In_704,In_214);
and U372 (N_372,In_819,In_1113);
or U373 (N_373,In_718,In_300);
or U374 (N_374,In_1439,In_1116);
xnor U375 (N_375,In_293,In_274);
and U376 (N_376,In_538,In_709);
xor U377 (N_377,In_656,In_1296);
or U378 (N_378,In_951,In_1666);
xnor U379 (N_379,In_1066,In_1398);
and U380 (N_380,In_386,In_1385);
nor U381 (N_381,In_897,In_1200);
or U382 (N_382,In_155,In_1012);
or U383 (N_383,In_802,In_1993);
nand U384 (N_384,In_1708,In_41);
nand U385 (N_385,In_1873,In_828);
nand U386 (N_386,In_1855,In_1475);
or U387 (N_387,In_246,In_941);
and U388 (N_388,In_317,In_580);
or U389 (N_389,In_128,In_627);
xor U390 (N_390,In_449,In_1571);
or U391 (N_391,In_494,In_59);
nor U392 (N_392,In_341,In_456);
or U393 (N_393,In_1163,In_942);
and U394 (N_394,In_1483,In_602);
or U395 (N_395,In_1312,In_748);
xnor U396 (N_396,In_1626,In_1755);
nand U397 (N_397,In_149,In_1480);
or U398 (N_398,In_11,In_1738);
xnor U399 (N_399,In_1495,In_407);
nor U400 (N_400,In_778,In_1752);
or U401 (N_401,In_624,In_445);
or U402 (N_402,In_927,In_1231);
nor U403 (N_403,In_399,In_868);
or U404 (N_404,In_21,In_997);
xnor U405 (N_405,In_975,In_15);
nand U406 (N_406,In_454,In_1256);
and U407 (N_407,In_622,In_832);
xnor U408 (N_408,In_962,In_187);
nand U409 (N_409,In_990,In_1288);
or U410 (N_410,In_1014,In_175);
xor U411 (N_411,In_1629,In_1206);
or U412 (N_412,In_1426,In_1545);
nor U413 (N_413,In_301,In_584);
nand U414 (N_414,In_1970,In_842);
nor U415 (N_415,In_1332,In_910);
or U416 (N_416,In_810,In_118);
nor U417 (N_417,In_1065,In_270);
or U418 (N_418,In_1469,In_620);
or U419 (N_419,In_791,In_1059);
or U420 (N_420,In_618,In_90);
xor U421 (N_421,In_859,In_1323);
nand U422 (N_422,In_751,In_1631);
and U423 (N_423,In_1304,In_348);
or U424 (N_424,In_247,In_1132);
and U425 (N_425,In_1816,In_1757);
nand U426 (N_426,In_659,In_1386);
or U427 (N_427,In_290,In_1912);
nor U428 (N_428,In_883,In_535);
or U429 (N_429,In_817,In_379);
nor U430 (N_430,In_1997,In_561);
or U431 (N_431,In_63,In_1488);
or U432 (N_432,In_1096,In_1076);
nand U433 (N_433,In_1390,In_978);
xor U434 (N_434,In_1056,In_1236);
nor U435 (N_435,In_1419,In_637);
and U436 (N_436,In_1031,In_937);
and U437 (N_437,In_1175,In_451);
nand U438 (N_438,In_418,In_1082);
nor U439 (N_439,In_1440,In_1811);
xor U440 (N_440,In_333,In_1020);
or U441 (N_441,In_597,In_1599);
or U442 (N_442,In_1922,In_846);
and U443 (N_443,In_1669,In_1637);
nor U444 (N_444,In_163,In_1420);
nand U445 (N_445,In_394,In_1593);
xor U446 (N_446,In_102,In_195);
xnor U447 (N_447,In_2,In_936);
or U448 (N_448,In_731,In_1272);
xor U449 (N_449,In_437,In_478);
nand U450 (N_450,In_176,In_1406);
xnor U451 (N_451,In_1383,In_357);
xor U452 (N_452,In_626,In_1147);
xnor U453 (N_453,In_229,In_1977);
xnor U454 (N_454,In_1465,In_1919);
xor U455 (N_455,In_1558,In_1411);
and U456 (N_456,In_1265,In_758);
or U457 (N_457,In_1779,In_1706);
and U458 (N_458,In_1652,In_1618);
xnor U459 (N_459,In_682,In_779);
xnor U460 (N_460,In_1235,In_998);
and U461 (N_461,In_1778,In_1140);
and U462 (N_462,In_1790,In_1763);
nand U463 (N_463,In_603,In_1871);
nor U464 (N_464,In_512,In_536);
xnor U465 (N_465,In_1954,In_1622);
xnor U466 (N_466,In_1731,In_37);
or U467 (N_467,In_1417,In_1301);
and U468 (N_468,In_780,In_1358);
xor U469 (N_469,In_493,In_1902);
nor U470 (N_470,In_1058,In_572);
nor U471 (N_471,In_306,In_1157);
and U472 (N_472,In_1785,In_398);
and U473 (N_473,In_660,In_73);
and U474 (N_474,In_6,In_403);
and U475 (N_475,In_850,In_460);
nor U476 (N_476,In_1858,In_600);
nand U477 (N_477,In_13,In_139);
nand U478 (N_478,In_574,In_609);
nor U479 (N_479,In_857,In_1998);
or U480 (N_480,In_901,In_191);
xnor U481 (N_481,In_1414,In_1486);
nand U482 (N_482,In_1840,In_77);
xnor U483 (N_483,In_1313,In_1727);
nand U484 (N_484,In_814,In_598);
nor U485 (N_485,In_1579,In_1262);
nand U486 (N_486,In_1112,In_556);
xor U487 (N_487,In_1893,In_1384);
or U488 (N_488,In_158,In_1610);
or U489 (N_489,In_690,In_1748);
and U490 (N_490,In_354,In_1454);
and U491 (N_491,In_1090,In_994);
xnor U492 (N_492,In_534,In_756);
and U493 (N_493,In_1951,In_258);
nor U494 (N_494,In_1463,In_1184);
and U495 (N_495,In_636,In_1380);
nor U496 (N_496,In_50,In_813);
xnor U497 (N_497,In_12,In_1111);
or U498 (N_498,In_965,In_615);
and U499 (N_499,In_1222,In_727);
nor U500 (N_500,In_1298,In_435);
and U501 (N_501,In_1188,In_1473);
nand U502 (N_502,In_986,In_1671);
or U503 (N_503,In_1144,In_1309);
nand U504 (N_504,In_1,In_319);
xnor U505 (N_505,In_1928,In_1693);
or U506 (N_506,In_1217,In_638);
or U507 (N_507,In_472,In_1250);
xor U508 (N_508,In_1684,In_481);
xnor U509 (N_509,In_205,In_352);
or U510 (N_510,In_431,In_1702);
nor U511 (N_511,In_1590,In_1172);
and U512 (N_512,In_159,In_800);
and U513 (N_513,In_402,In_1771);
or U514 (N_514,In_1045,In_1397);
or U515 (N_515,In_1451,In_629);
nand U516 (N_516,In_1089,In_169);
nor U517 (N_517,In_1522,In_80);
nor U518 (N_518,In_1602,In_579);
or U519 (N_519,In_1900,In_946);
and U520 (N_520,In_503,In_428);
nor U521 (N_521,In_1129,In_1865);
nand U522 (N_522,In_1831,In_1710);
nor U523 (N_523,In_1805,In_1539);
nor U524 (N_524,In_1496,In_847);
or U525 (N_525,In_934,In_1531);
nor U526 (N_526,In_397,In_47);
xor U527 (N_527,In_186,In_226);
and U528 (N_528,In_373,In_496);
nor U529 (N_529,In_1552,In_1592);
or U530 (N_530,In_935,In_483);
and U531 (N_531,In_1218,In_439);
xor U532 (N_532,In_923,In_577);
nor U533 (N_533,In_468,In_843);
nand U534 (N_534,In_1973,In_1055);
and U535 (N_535,In_1761,In_444);
xnor U536 (N_536,In_1709,In_952);
xor U537 (N_537,In_742,In_1980);
xnor U538 (N_538,In_1018,In_1589);
nor U539 (N_539,In_249,In_838);
xor U540 (N_540,In_1028,In_1729);
and U541 (N_541,In_864,In_889);
and U542 (N_542,In_1934,In_144);
xor U543 (N_543,In_621,In_1501);
nor U544 (N_544,In_1224,In_675);
xor U545 (N_545,In_617,In_1987);
and U546 (N_546,In_1208,In_875);
xnor U547 (N_547,In_1804,In_415);
xnor U548 (N_548,In_1072,In_1765);
nor U549 (N_549,In_740,In_42);
and U550 (N_550,In_129,In_539);
nor U551 (N_551,In_1432,In_1192);
nand U552 (N_552,In_1864,In_1654);
nand U553 (N_553,In_43,In_1523);
xnor U554 (N_554,In_1470,In_610);
or U555 (N_555,In_771,In_1546);
nor U556 (N_556,In_833,In_244);
nand U557 (N_557,In_981,In_1768);
or U558 (N_558,In_1650,In_16);
and U559 (N_559,In_1227,In_1458);
nor U560 (N_560,In_1635,In_239);
nand U561 (N_561,In_1095,In_596);
and U562 (N_562,In_1564,In_1433);
nand U563 (N_563,In_501,In_719);
nor U564 (N_564,In_1280,In_1553);
nand U565 (N_565,In_1103,In_741);
xnor U566 (N_566,In_522,In_217);
nand U567 (N_567,In_1929,In_808);
nand U568 (N_568,In_452,In_929);
or U569 (N_569,In_498,In_1688);
nand U570 (N_570,In_1949,In_1560);
xnor U571 (N_571,In_641,In_1787);
or U572 (N_572,In_338,In_1557);
nor U573 (N_573,In_697,In_1673);
and U574 (N_574,In_1422,In_1945);
and U575 (N_575,In_1281,In_57);
and U576 (N_576,In_912,In_1046);
xor U577 (N_577,In_488,In_1686);
and U578 (N_578,In_122,In_368);
nor U579 (N_579,In_330,In_1201);
nor U580 (N_580,In_1214,In_1083);
xnor U581 (N_581,In_963,In_508);
and U582 (N_582,In_798,In_54);
nand U583 (N_583,In_1675,In_592);
and U584 (N_584,In_1707,In_31);
xnor U585 (N_585,In_1126,In_1202);
or U586 (N_586,In_261,In_349);
xor U587 (N_587,In_82,In_1530);
xnor U588 (N_588,In_612,In_966);
xnor U589 (N_589,In_792,In_1773);
and U590 (N_590,In_870,In_1447);
xnor U591 (N_591,In_1061,In_1086);
or U592 (N_592,In_1356,In_1211);
nor U593 (N_593,In_264,In_1868);
nand U594 (N_594,In_135,In_807);
or U595 (N_595,In_1405,In_1881);
xnor U596 (N_596,In_1817,In_1242);
and U597 (N_597,In_964,In_1448);
xor U598 (N_598,In_1156,In_1085);
and U599 (N_599,In_928,In_1554);
xor U600 (N_600,In_1963,In_1430);
xnor U601 (N_601,In_1606,In_369);
nand U602 (N_602,In_499,In_1536);
nor U603 (N_603,In_240,In_5);
or U604 (N_604,In_1979,In_1649);
nand U605 (N_605,In_1299,In_1425);
nand U606 (N_606,In_433,In_805);
or U607 (N_607,In_1155,In_1283);
xor U608 (N_608,In_1029,In_86);
or U609 (N_609,In_845,In_1335);
nand U610 (N_610,In_1006,In_1328);
nand U611 (N_611,In_1452,In_1418);
or U612 (N_612,In_359,In_237);
nand U613 (N_613,In_666,In_74);
nor U614 (N_614,In_1121,In_245);
and U615 (N_615,In_1287,In_1219);
or U616 (N_616,In_1247,In_385);
nand U617 (N_617,In_1842,In_396);
or U618 (N_618,In_211,In_111);
and U619 (N_619,In_1966,In_921);
xnor U620 (N_620,In_268,In_787);
nand U621 (N_621,In_922,In_1723);
nand U622 (N_622,In_194,In_1489);
nor U623 (N_623,In_541,In_455);
or U624 (N_624,In_1266,In_145);
or U625 (N_625,In_1641,In_1780);
nor U626 (N_626,In_1449,In_969);
nor U627 (N_627,In_325,In_528);
and U628 (N_628,In_1782,In_761);
nand U629 (N_629,In_344,In_406);
and U630 (N_630,In_1775,In_430);
nand U631 (N_631,In_797,In_465);
nand U632 (N_632,In_1510,In_1889);
or U633 (N_633,In_1918,In_531);
xor U634 (N_634,In_1290,In_1369);
xnor U635 (N_635,In_1884,In_1409);
or U636 (N_636,In_753,In_22);
and U637 (N_637,In_939,In_277);
nand U638 (N_638,In_1494,In_984);
nand U639 (N_639,In_1471,In_1931);
nand U640 (N_640,In_726,In_1330);
nor U641 (N_641,In_393,In_914);
nor U642 (N_642,In_1429,In_1682);
nor U643 (N_643,In_106,In_417);
xor U644 (N_644,In_1835,In_1762);
xnor U645 (N_645,In_999,In_1252);
or U646 (N_646,In_114,In_1513);
or U647 (N_647,In_1899,In_1381);
and U648 (N_648,In_1193,In_151);
nor U649 (N_649,In_327,In_1388);
or U650 (N_650,In_1274,In_1361);
nor U651 (N_651,In_1585,In_1992);
or U652 (N_652,In_1146,In_1535);
and U653 (N_653,In_1832,In_105);
or U654 (N_654,In_382,In_178);
nor U655 (N_655,In_1044,In_852);
nand U656 (N_656,In_1908,In_1355);
nor U657 (N_657,In_1442,In_1607);
nor U658 (N_658,In_543,In_1903);
or U659 (N_659,In_1735,In_1050);
or U660 (N_660,In_924,In_1098);
nor U661 (N_661,In_523,In_747);
nor U662 (N_662,In_1017,In_1540);
or U663 (N_663,In_1254,In_137);
nor U664 (N_664,In_487,In_64);
nor U665 (N_665,In_94,In_1067);
xnor U666 (N_666,In_108,In_275);
or U667 (N_667,In_1783,In_1077);
or U668 (N_668,In_1955,In_208);
nor U669 (N_669,In_1070,In_1745);
nor U670 (N_670,In_674,In_594);
nand U671 (N_671,In_234,In_250);
xor U672 (N_672,In_1069,In_1541);
and U673 (N_673,In_1415,In_957);
and U674 (N_674,In_759,In_1806);
nor U675 (N_675,In_1583,In_930);
or U676 (N_676,In_1234,In_989);
nor U677 (N_677,In_218,In_475);
or U678 (N_678,In_1705,In_25);
or U679 (N_679,In_1183,In_1830);
nand U680 (N_680,In_1052,In_652);
xnor U681 (N_681,In_27,In_1492);
nor U682 (N_682,In_1062,In_339);
and U683 (N_683,In_1911,In_848);
and U684 (N_684,In_530,In_423);
or U685 (N_685,In_1668,In_769);
xor U686 (N_686,In_663,In_1700);
and U687 (N_687,In_554,In_473);
xnor U688 (N_688,In_1003,In_1724);
and U689 (N_689,In_1493,In_497);
and U690 (N_690,In_356,In_613);
or U691 (N_691,In_1504,In_831);
and U692 (N_692,In_1643,In_1883);
or U693 (N_693,In_1852,In_97);
nor U694 (N_694,In_1001,In_45);
nor U695 (N_695,In_1907,In_968);
nor U696 (N_696,In_1759,In_448);
nor U697 (N_697,In_1075,In_303);
and U698 (N_698,In_835,In_1588);
nand U699 (N_699,In_1845,In_1983);
or U700 (N_700,In_1134,In_1826);
and U701 (N_701,In_1249,In_1813);
nor U702 (N_702,In_695,In_1174);
xnor U703 (N_703,In_1642,In_1339);
or U704 (N_704,In_1233,In_567);
xor U705 (N_705,In_171,In_1833);
nor U706 (N_706,In_1519,In_302);
nor U707 (N_707,In_678,In_347);
nor U708 (N_708,In_1747,In_737);
nor U709 (N_709,In_1810,In_1071);
or U710 (N_710,In_702,In_1547);
nor U711 (N_711,In_1796,In_1225);
xor U712 (N_712,In_931,In_1591);
or U713 (N_713,In_1857,In_1109);
nand U714 (N_714,In_908,In_1632);
xor U715 (N_715,In_1292,In_1674);
or U716 (N_716,In_143,In_1468);
xnor U717 (N_717,In_1119,In_524);
nand U718 (N_718,In_1466,In_1751);
nor U719 (N_719,In_977,In_1357);
nand U720 (N_720,In_1036,In_1758);
nor U721 (N_721,In_440,In_520);
and U722 (N_722,In_1008,In_471);
and U723 (N_723,In_1703,In_1568);
xor U724 (N_724,In_1311,In_1007);
and U725 (N_725,In_166,In_1372);
and U726 (N_726,In_1943,In_829);
xnor U727 (N_727,In_1326,In_900);
xor U728 (N_728,In_1732,In_1337);
nand U729 (N_729,In_858,In_1027);
and U730 (N_730,In_1457,In_1822);
and U731 (N_731,In_184,In_1484);
xor U732 (N_732,In_1793,In_982);
or U733 (N_733,In_1798,In_563);
and U734 (N_734,In_1057,In_170);
and U735 (N_735,In_477,In_1561);
and U736 (N_736,In_1861,In_547);
and U737 (N_737,In_1807,In_316);
or U738 (N_738,In_1658,In_1968);
nor U739 (N_739,In_248,In_1181);
or U740 (N_740,In_1853,In_1042);
or U741 (N_741,In_1784,In_890);
nand U742 (N_742,In_542,In_589);
or U743 (N_743,In_557,In_222);
or U744 (N_744,In_1906,In_1149);
nor U745 (N_745,In_1267,In_1739);
nand U746 (N_746,In_1026,In_782);
nor U747 (N_747,In_680,In_793);
and U748 (N_748,In_1497,In_14);
nor U749 (N_749,In_495,In_736);
xor U750 (N_750,In_1697,In_1226);
xor U751 (N_751,In_905,In_1133);
or U752 (N_752,In_866,In_326);
or U753 (N_753,In_409,In_1063);
and U754 (N_754,In_948,In_1416);
or U755 (N_755,In_342,In_1295);
xor U756 (N_756,In_351,In_372);
nand U757 (N_757,In_757,In_1382);
and U758 (N_758,In_99,In_1944);
or U759 (N_759,In_684,In_141);
nand U760 (N_760,In_1081,In_377);
xnor U761 (N_761,In_117,In_1570);
nor U762 (N_762,In_1694,In_1638);
xor U763 (N_763,In_1207,In_1455);
nand U764 (N_764,In_788,In_405);
and U765 (N_765,In_4,In_93);
xnor U766 (N_766,In_1994,In_30);
nor U767 (N_767,In_1491,In_711);
or U768 (N_768,In_1245,In_1803);
xor U769 (N_769,In_1623,In_1965);
xor U770 (N_770,In_591,In_1097);
and U771 (N_771,In_1093,In_1005);
nor U772 (N_772,In_1353,In_1663);
and U773 (N_773,In_862,In_426);
nor U774 (N_774,In_1995,In_818);
or U775 (N_775,In_161,In_1948);
or U776 (N_776,In_1371,In_593);
or U777 (N_777,In_46,In_485);
and U778 (N_778,In_1612,In_1107);
nor U779 (N_779,In_1347,In_328);
and U780 (N_780,In_904,In_1544);
xnor U781 (N_781,In_560,In_1653);
nor U782 (N_782,In_1209,In_1812);
xnor U783 (N_783,In_1964,In_1836);
xnor U784 (N_784,In_429,In_1377);
or U785 (N_785,In_1619,In_947);
nor U786 (N_786,In_955,In_1123);
xor U787 (N_787,In_749,In_1185);
nand U788 (N_788,In_1011,In_1594);
nand U789 (N_789,In_1152,In_1692);
xnor U790 (N_790,In_231,In_1102);
or U791 (N_791,In_201,In_664);
or U792 (N_792,In_712,In_1957);
nand U793 (N_793,In_432,In_881);
or U794 (N_794,In_112,In_1507);
nand U795 (N_795,In_289,In_364);
nand U796 (N_796,In_305,In_987);
nor U797 (N_797,In_390,In_958);
nand U798 (N_798,In_909,In_1198);
nor U799 (N_799,In_1880,In_29);
nand U800 (N_800,In_1917,In_1986);
nor U801 (N_801,In_146,In_925);
nand U802 (N_802,In_1261,In_1613);
or U803 (N_803,In_1542,In_1801);
nor U804 (N_804,In_1104,In_564);
and U805 (N_805,In_565,In_332);
xor U806 (N_806,In_1164,In_1244);
xor U807 (N_807,In_1127,In_233);
nor U808 (N_808,In_1043,In_654);
nand U809 (N_809,In_844,In_119);
or U810 (N_810,In_1392,In_1886);
xnor U811 (N_811,In_507,In_7);
nand U812 (N_812,In_1100,In_299);
nand U813 (N_813,In_1976,In_1294);
xnor U814 (N_814,In_1305,In_880);
nand U815 (N_815,In_750,In_321);
nor U816 (N_816,In_1962,In_174);
xnor U817 (N_817,In_1344,In_148);
and U818 (N_818,In_1932,In_1314);
and U819 (N_819,In_1841,In_1582);
nor U820 (N_820,In_1559,In_604);
or U821 (N_821,In_401,In_79);
nand U822 (N_822,In_983,In_873);
nand U823 (N_823,In_1269,In_1712);
or U824 (N_824,In_1000,In_606);
nand U825 (N_825,In_738,In_1010);
xor U826 (N_826,In_92,In_1935);
nand U827 (N_827,In_1080,In_677);
and U828 (N_828,In_1137,In_768);
and U829 (N_829,In_259,In_840);
nand U830 (N_830,In_1566,In_172);
xnor U831 (N_831,In_1754,In_1876);
and U832 (N_832,In_1329,In_1285);
xor U833 (N_833,In_1023,In_1940);
nand U834 (N_834,In_1456,In_1799);
nor U835 (N_835,In_375,In_1737);
and U836 (N_836,In_506,In_1399);
nand U837 (N_837,In_427,In_1517);
nand U838 (N_838,In_1701,In_1160);
or U839 (N_839,In_36,In_1605);
or U840 (N_840,In_529,In_313);
nor U841 (N_841,In_1319,In_882);
xor U842 (N_842,In_891,In_60);
and U843 (N_843,In_312,In_1124);
xor U844 (N_844,In_1586,In_1644);
or U845 (N_845,In_913,In_1108);
xor U846 (N_846,In_1033,In_204);
xnor U847 (N_847,In_1721,In_1953);
and U848 (N_848,In_1659,In_943);
xnor U849 (N_849,In_1844,In_164);
nor U850 (N_850,In_825,In_1190);
or U851 (N_851,In_1698,In_1189);
nand U852 (N_852,In_540,In_1136);
nor U853 (N_853,In_1958,In_953);
nand U854 (N_854,In_1837,In_551);
nand U855 (N_855,In_121,In_1040);
and U856 (N_856,In_1781,In_1597);
nand U857 (N_857,In_1854,In_898);
and U858 (N_858,In_1402,In_1286);
or U859 (N_859,In_732,In_1037);
or U860 (N_860,In_115,In_705);
or U861 (N_861,In_1151,In_933);
or U862 (N_862,In_1516,In_1348);
xor U863 (N_863,In_294,In_1350);
or U864 (N_864,In_1297,In_1651);
and U865 (N_865,In_1898,In_182);
nand U866 (N_866,In_1238,In_1985);
and U867 (N_867,In_867,In_414);
nor U868 (N_868,In_150,In_1981);
and U869 (N_869,In_710,In_1598);
xnor U870 (N_870,In_1646,In_288);
and U871 (N_871,In_116,In_996);
nor U872 (N_872,In_1215,In_1972);
nor U873 (N_873,In_1284,In_1615);
and U874 (N_874,In_228,In_367);
nor U875 (N_875,In_1366,In_569);
xnor U876 (N_876,In_360,In_1364);
and U877 (N_877,In_1950,In_253);
or U878 (N_878,In_126,In_458);
and U879 (N_879,In_1518,In_745);
and U880 (N_880,In_255,In_623);
xor U881 (N_881,In_945,In_1138);
and U882 (N_882,In_263,In_856);
xor U883 (N_883,In_1434,In_1015);
nand U884 (N_884,In_1221,In_1342);
xor U885 (N_885,In_1930,In_671);
xor U886 (N_886,In_1770,In_123);
nand U887 (N_887,In_1091,In_932);
nand U888 (N_888,In_1719,In_1984);
nand U889 (N_889,In_1349,In_1410);
xor U890 (N_890,In_1431,In_765);
and U891 (N_891,In_1060,In_973);
xnor U892 (N_892,In_400,In_1087);
xor U893 (N_893,In_605,In_1110);
or U894 (N_894,In_19,In_1656);
or U895 (N_895,In_1374,In_1711);
nor U896 (N_896,In_470,In_1403);
nor U897 (N_897,In_51,In_1679);
xnor U898 (N_898,In_88,In_582);
nand U899 (N_899,In_179,In_860);
nand U900 (N_900,In_1064,In_1142);
xor U901 (N_901,In_284,In_381);
or U902 (N_902,In_1614,In_1394);
or U903 (N_903,In_279,In_276);
xnor U904 (N_904,In_474,In_20);
or U905 (N_905,In_1715,In_411);
xnor U906 (N_906,In_416,In_707);
nor U907 (N_907,In_113,In_190);
xnor U908 (N_908,In_1320,In_504);
nand U909 (N_909,In_722,In_643);
xnor U910 (N_910,In_1230,In_273);
or U911 (N_911,In_961,In_894);
nor U912 (N_912,In_1569,In_783);
nand U913 (N_913,In_812,In_693);
nand U914 (N_914,In_1460,In_177);
and U915 (N_915,In_878,In_1520);
nand U916 (N_916,In_1354,In_720);
and U917 (N_917,In_735,In_1543);
nand U918 (N_918,In_1196,In_1396);
or U919 (N_919,In_583,In_1078);
xor U920 (N_920,In_1341,In_1482);
nor U921 (N_921,In_1909,In_658);
nand U922 (N_922,In_1572,In_1580);
or U923 (N_923,In_1293,In_1034);
xor U924 (N_924,In_1971,In_1577);
xnor U925 (N_925,In_1609,In_1576);
nor U926 (N_926,In_876,In_1336);
or U927 (N_927,In_1343,In_269);
nand U928 (N_928,In_1153,In_1464);
or U929 (N_929,In_670,In_760);
or U930 (N_930,In_766,In_1407);
and U931 (N_931,In_180,In_61);
or U932 (N_932,In_157,In_1167);
and U933 (N_933,In_84,In_1551);
xor U934 (N_934,In_83,In_104);
nor U935 (N_935,In_1079,In_672);
or U936 (N_936,In_1600,In_1499);
or U937 (N_937,In_1237,In_815);
xnor U938 (N_938,In_1750,In_388);
xor U939 (N_939,In_1938,In_634);
or U940 (N_940,In_1444,In_784);
nor U941 (N_941,In_980,In_795);
nor U942 (N_942,In_1306,In_648);
and U943 (N_943,In_206,In_1375);
nor U944 (N_944,In_698,In_796);
and U945 (N_945,In_691,In_879);
or U946 (N_946,In_1505,In_1740);
xor U947 (N_947,In_822,In_1216);
nor U948 (N_948,In_1860,In_68);
or U949 (N_949,In_462,In_1220);
and U950 (N_950,In_1628,In_716);
xnor U951 (N_951,In_1878,In_662);
or U952 (N_952,In_1901,In_804);
nand U953 (N_953,In_993,In_52);
and U954 (N_954,In_785,In_611);
and U955 (N_955,In_1827,In_138);
xnor U956 (N_956,In_1937,In_1587);
nand U957 (N_957,In_408,In_220);
nor U958 (N_958,In_1680,In_1490);
or U959 (N_959,In_1555,In_1887);
or U960 (N_960,In_221,In_1874);
or U961 (N_961,In_1318,In_1317);
nor U962 (N_962,In_1843,In_1270);
or U963 (N_963,In_1743,In_1004);
nor U964 (N_964,In_26,In_1648);
and U965 (N_965,In_601,In_17);
or U966 (N_966,In_33,In_1581);
nor U967 (N_967,In_1178,In_630);
nor U968 (N_968,In_1168,In_1338);
nand U969 (N_969,In_781,In_1169);
nor U970 (N_970,In_926,In_616);
nand U971 (N_971,In_1904,In_824);
nand U972 (N_972,In_1094,In_70);
or U973 (N_973,In_1791,In_1625);
nand U974 (N_974,In_446,In_421);
xor U975 (N_975,In_152,In_307);
xor U976 (N_976,In_96,In_1978);
nor U977 (N_977,In_78,In_553);
nor U978 (N_978,In_715,In_1749);
nor U979 (N_979,In_1502,In_1240);
xor U980 (N_980,In_1814,In_1616);
nand U981 (N_981,In_545,In_869);
nor U982 (N_982,In_1506,In_1892);
or U983 (N_983,In_323,In_1145);
xnor U984 (N_984,In_1143,In_100);
nor U985 (N_985,In_335,In_1186);
and U986 (N_986,In_632,In_224);
and U987 (N_987,In_685,In_238);
nand U988 (N_988,In_653,In_227);
nor U989 (N_989,In_1450,In_1533);
nor U990 (N_990,In_762,In_1808);
xor U991 (N_991,In_976,In_1437);
or U992 (N_992,In_1511,In_1611);
nor U993 (N_993,In_1021,In_1203);
or U994 (N_994,In_1846,In_725);
xnor U995 (N_995,In_1624,In_834);
xnor U996 (N_996,In_1373,In_1128);
nand U997 (N_997,In_1333,In_502);
nor U998 (N_998,In_1639,In_457);
or U999 (N_999,In_1988,In_1563);
xor U1000 (N_1000,In_308,In_1793);
nand U1001 (N_1001,In_865,In_1380);
nor U1002 (N_1002,In_295,In_1470);
or U1003 (N_1003,In_715,In_1224);
nor U1004 (N_1004,In_251,In_1768);
xor U1005 (N_1005,In_1695,In_1759);
or U1006 (N_1006,In_1969,In_433);
xor U1007 (N_1007,In_805,In_116);
xor U1008 (N_1008,In_1870,In_1604);
or U1009 (N_1009,In_646,In_1933);
nor U1010 (N_1010,In_128,In_607);
and U1011 (N_1011,In_1403,In_983);
and U1012 (N_1012,In_1904,In_1333);
nor U1013 (N_1013,In_1914,In_1527);
nor U1014 (N_1014,In_1775,In_215);
or U1015 (N_1015,In_884,In_1343);
xnor U1016 (N_1016,In_1168,In_1763);
and U1017 (N_1017,In_1417,In_1494);
or U1018 (N_1018,In_1580,In_906);
xor U1019 (N_1019,In_38,In_1596);
nor U1020 (N_1020,In_51,In_952);
or U1021 (N_1021,In_1760,In_704);
xnor U1022 (N_1022,In_1881,In_673);
nor U1023 (N_1023,In_700,In_311);
nor U1024 (N_1024,In_952,In_1645);
and U1025 (N_1025,In_239,In_46);
and U1026 (N_1026,In_1109,In_1044);
nand U1027 (N_1027,In_667,In_1927);
nor U1028 (N_1028,In_1988,In_448);
or U1029 (N_1029,In_290,In_960);
xor U1030 (N_1030,In_774,In_372);
and U1031 (N_1031,In_268,In_1290);
and U1032 (N_1032,In_1157,In_948);
or U1033 (N_1033,In_1473,In_1115);
nor U1034 (N_1034,In_1152,In_647);
xnor U1035 (N_1035,In_1105,In_394);
and U1036 (N_1036,In_1068,In_828);
and U1037 (N_1037,In_1033,In_1030);
nor U1038 (N_1038,In_1852,In_1148);
nand U1039 (N_1039,In_1437,In_276);
and U1040 (N_1040,In_855,In_1140);
nor U1041 (N_1041,In_702,In_469);
and U1042 (N_1042,In_1305,In_331);
and U1043 (N_1043,In_1056,In_551);
nand U1044 (N_1044,In_883,In_1874);
nand U1045 (N_1045,In_789,In_1571);
or U1046 (N_1046,In_1754,In_879);
xnor U1047 (N_1047,In_107,In_767);
nor U1048 (N_1048,In_37,In_277);
and U1049 (N_1049,In_1865,In_1215);
or U1050 (N_1050,In_1278,In_510);
and U1051 (N_1051,In_33,In_1482);
or U1052 (N_1052,In_88,In_1860);
xor U1053 (N_1053,In_1217,In_1397);
and U1054 (N_1054,In_1581,In_1472);
and U1055 (N_1055,In_1135,In_163);
nand U1056 (N_1056,In_316,In_1684);
nor U1057 (N_1057,In_1784,In_1301);
xor U1058 (N_1058,In_1998,In_336);
nor U1059 (N_1059,In_327,In_297);
nand U1060 (N_1060,In_767,In_552);
or U1061 (N_1061,In_1818,In_529);
xnor U1062 (N_1062,In_719,In_1186);
nor U1063 (N_1063,In_1784,In_1015);
xnor U1064 (N_1064,In_1557,In_151);
nor U1065 (N_1065,In_1039,In_830);
xnor U1066 (N_1066,In_1436,In_756);
nand U1067 (N_1067,In_1727,In_595);
xnor U1068 (N_1068,In_1920,In_1561);
nand U1069 (N_1069,In_1076,In_857);
xnor U1070 (N_1070,In_929,In_736);
nand U1071 (N_1071,In_1507,In_1125);
and U1072 (N_1072,In_817,In_330);
xor U1073 (N_1073,In_416,In_858);
xor U1074 (N_1074,In_1277,In_465);
and U1075 (N_1075,In_1920,In_1900);
nor U1076 (N_1076,In_640,In_1541);
xnor U1077 (N_1077,In_142,In_1943);
xor U1078 (N_1078,In_1929,In_1105);
xor U1079 (N_1079,In_1819,In_1427);
nor U1080 (N_1080,In_1855,In_1002);
xor U1081 (N_1081,In_782,In_10);
or U1082 (N_1082,In_1975,In_1424);
nor U1083 (N_1083,In_736,In_1551);
or U1084 (N_1084,In_317,In_1701);
or U1085 (N_1085,In_1564,In_788);
and U1086 (N_1086,In_1790,In_1767);
nor U1087 (N_1087,In_1298,In_1444);
and U1088 (N_1088,In_569,In_856);
or U1089 (N_1089,In_1156,In_989);
xnor U1090 (N_1090,In_1326,In_173);
nor U1091 (N_1091,In_1798,In_1963);
nand U1092 (N_1092,In_387,In_1782);
nand U1093 (N_1093,In_1867,In_1549);
or U1094 (N_1094,In_1108,In_70);
xor U1095 (N_1095,In_1832,In_1450);
or U1096 (N_1096,In_435,In_181);
nand U1097 (N_1097,In_878,In_1480);
xnor U1098 (N_1098,In_545,In_565);
xor U1099 (N_1099,In_1552,In_1176);
xor U1100 (N_1100,In_1734,In_1145);
or U1101 (N_1101,In_1552,In_102);
xnor U1102 (N_1102,In_728,In_1810);
nor U1103 (N_1103,In_1757,In_773);
or U1104 (N_1104,In_1820,In_222);
nand U1105 (N_1105,In_1119,In_914);
nand U1106 (N_1106,In_202,In_288);
or U1107 (N_1107,In_1683,In_1609);
xnor U1108 (N_1108,In_1638,In_1438);
nor U1109 (N_1109,In_1827,In_975);
xor U1110 (N_1110,In_933,In_1638);
and U1111 (N_1111,In_123,In_1893);
xor U1112 (N_1112,In_1944,In_713);
nor U1113 (N_1113,In_736,In_1756);
and U1114 (N_1114,In_1076,In_1907);
nand U1115 (N_1115,In_792,In_378);
or U1116 (N_1116,In_1826,In_1278);
and U1117 (N_1117,In_762,In_1120);
nand U1118 (N_1118,In_1300,In_955);
xor U1119 (N_1119,In_1331,In_1155);
or U1120 (N_1120,In_1451,In_1573);
xor U1121 (N_1121,In_1943,In_254);
nand U1122 (N_1122,In_1601,In_1067);
xor U1123 (N_1123,In_354,In_1113);
or U1124 (N_1124,In_1349,In_438);
and U1125 (N_1125,In_986,In_1231);
or U1126 (N_1126,In_1051,In_1343);
xor U1127 (N_1127,In_197,In_827);
nor U1128 (N_1128,In_1554,In_873);
nor U1129 (N_1129,In_789,In_800);
and U1130 (N_1130,In_404,In_475);
xor U1131 (N_1131,In_613,In_1191);
and U1132 (N_1132,In_1296,In_381);
or U1133 (N_1133,In_1135,In_336);
nand U1134 (N_1134,In_151,In_870);
or U1135 (N_1135,In_168,In_608);
or U1136 (N_1136,In_1049,In_85);
nand U1137 (N_1137,In_1429,In_271);
and U1138 (N_1138,In_1447,In_320);
nand U1139 (N_1139,In_679,In_233);
nor U1140 (N_1140,In_685,In_782);
and U1141 (N_1141,In_1071,In_402);
or U1142 (N_1142,In_1779,In_936);
and U1143 (N_1143,In_1915,In_448);
or U1144 (N_1144,In_656,In_62);
nor U1145 (N_1145,In_783,In_760);
nor U1146 (N_1146,In_908,In_1387);
and U1147 (N_1147,In_647,In_1128);
and U1148 (N_1148,In_1805,In_270);
and U1149 (N_1149,In_212,In_1961);
nand U1150 (N_1150,In_320,In_1395);
and U1151 (N_1151,In_1094,In_1604);
nand U1152 (N_1152,In_1130,In_1013);
xnor U1153 (N_1153,In_217,In_590);
or U1154 (N_1154,In_1064,In_1491);
nor U1155 (N_1155,In_419,In_1829);
or U1156 (N_1156,In_1487,In_1861);
nand U1157 (N_1157,In_436,In_1277);
and U1158 (N_1158,In_1033,In_1011);
and U1159 (N_1159,In_1893,In_651);
nand U1160 (N_1160,In_1900,In_1936);
nor U1161 (N_1161,In_347,In_777);
nor U1162 (N_1162,In_1423,In_144);
or U1163 (N_1163,In_1936,In_1274);
nand U1164 (N_1164,In_1319,In_489);
nand U1165 (N_1165,In_1973,In_173);
nor U1166 (N_1166,In_968,In_946);
nor U1167 (N_1167,In_1277,In_1078);
or U1168 (N_1168,In_243,In_436);
nor U1169 (N_1169,In_1555,In_1599);
nand U1170 (N_1170,In_435,In_1040);
and U1171 (N_1171,In_197,In_1208);
nor U1172 (N_1172,In_1175,In_720);
and U1173 (N_1173,In_903,In_178);
and U1174 (N_1174,In_521,In_81);
and U1175 (N_1175,In_379,In_22);
and U1176 (N_1176,In_1639,In_1076);
and U1177 (N_1177,In_1130,In_1774);
and U1178 (N_1178,In_549,In_875);
and U1179 (N_1179,In_738,In_1464);
or U1180 (N_1180,In_117,In_1178);
nor U1181 (N_1181,In_699,In_467);
or U1182 (N_1182,In_11,In_895);
and U1183 (N_1183,In_1812,In_797);
nand U1184 (N_1184,In_1601,In_711);
xnor U1185 (N_1185,In_427,In_1613);
nand U1186 (N_1186,In_763,In_1358);
and U1187 (N_1187,In_169,In_675);
xor U1188 (N_1188,In_291,In_450);
xnor U1189 (N_1189,In_1138,In_1794);
and U1190 (N_1190,In_448,In_685);
nor U1191 (N_1191,In_1289,In_554);
and U1192 (N_1192,In_9,In_153);
or U1193 (N_1193,In_1820,In_124);
nand U1194 (N_1194,In_1673,In_1029);
and U1195 (N_1195,In_443,In_1698);
nand U1196 (N_1196,In_1446,In_507);
and U1197 (N_1197,In_1005,In_742);
nand U1198 (N_1198,In_207,In_1480);
xor U1199 (N_1199,In_751,In_294);
nor U1200 (N_1200,In_49,In_1653);
nand U1201 (N_1201,In_190,In_43);
nand U1202 (N_1202,In_590,In_1354);
nor U1203 (N_1203,In_841,In_1138);
or U1204 (N_1204,In_891,In_539);
nand U1205 (N_1205,In_1250,In_1635);
and U1206 (N_1206,In_1465,In_1740);
xor U1207 (N_1207,In_929,In_3);
and U1208 (N_1208,In_925,In_1460);
xor U1209 (N_1209,In_900,In_295);
and U1210 (N_1210,In_868,In_82);
xor U1211 (N_1211,In_1790,In_1461);
or U1212 (N_1212,In_376,In_1533);
nand U1213 (N_1213,In_1729,In_729);
nand U1214 (N_1214,In_487,In_828);
xor U1215 (N_1215,In_1266,In_1982);
and U1216 (N_1216,In_1238,In_1787);
nand U1217 (N_1217,In_748,In_1201);
and U1218 (N_1218,In_242,In_1292);
and U1219 (N_1219,In_1584,In_1813);
and U1220 (N_1220,In_1271,In_926);
and U1221 (N_1221,In_1448,In_1162);
nand U1222 (N_1222,In_1648,In_873);
xnor U1223 (N_1223,In_1870,In_1186);
xnor U1224 (N_1224,In_1515,In_1464);
xor U1225 (N_1225,In_356,In_1061);
xor U1226 (N_1226,In_1622,In_680);
xor U1227 (N_1227,In_1492,In_1333);
or U1228 (N_1228,In_1801,In_54);
nor U1229 (N_1229,In_1268,In_483);
and U1230 (N_1230,In_1040,In_597);
nand U1231 (N_1231,In_1851,In_71);
or U1232 (N_1232,In_595,In_577);
nor U1233 (N_1233,In_62,In_542);
nor U1234 (N_1234,In_1509,In_225);
nor U1235 (N_1235,In_539,In_1341);
and U1236 (N_1236,In_516,In_1993);
nor U1237 (N_1237,In_866,In_1083);
nor U1238 (N_1238,In_1863,In_1636);
or U1239 (N_1239,In_942,In_99);
xnor U1240 (N_1240,In_927,In_1113);
xnor U1241 (N_1241,In_1744,In_607);
nor U1242 (N_1242,In_1081,In_783);
nand U1243 (N_1243,In_1524,In_441);
or U1244 (N_1244,In_184,In_780);
nor U1245 (N_1245,In_1169,In_970);
and U1246 (N_1246,In_61,In_906);
and U1247 (N_1247,In_1548,In_625);
or U1248 (N_1248,In_1809,In_1662);
and U1249 (N_1249,In_51,In_1321);
nand U1250 (N_1250,In_1584,In_387);
nand U1251 (N_1251,In_1446,In_1293);
nand U1252 (N_1252,In_746,In_1363);
and U1253 (N_1253,In_1279,In_153);
nand U1254 (N_1254,In_1042,In_1924);
or U1255 (N_1255,In_307,In_547);
and U1256 (N_1256,In_1424,In_619);
nor U1257 (N_1257,In_1828,In_261);
and U1258 (N_1258,In_256,In_1653);
nand U1259 (N_1259,In_722,In_884);
or U1260 (N_1260,In_297,In_614);
or U1261 (N_1261,In_1645,In_1232);
xor U1262 (N_1262,In_536,In_1454);
nor U1263 (N_1263,In_736,In_1484);
and U1264 (N_1264,In_363,In_513);
xnor U1265 (N_1265,In_59,In_1773);
or U1266 (N_1266,In_783,In_364);
nand U1267 (N_1267,In_1203,In_248);
xor U1268 (N_1268,In_549,In_909);
nand U1269 (N_1269,In_805,In_115);
xnor U1270 (N_1270,In_1484,In_1374);
nor U1271 (N_1271,In_742,In_1349);
and U1272 (N_1272,In_228,In_745);
and U1273 (N_1273,In_163,In_1486);
nor U1274 (N_1274,In_987,In_1435);
xnor U1275 (N_1275,In_1323,In_1561);
xor U1276 (N_1276,In_578,In_178);
or U1277 (N_1277,In_1218,In_633);
nor U1278 (N_1278,In_670,In_1754);
or U1279 (N_1279,In_582,In_1050);
xor U1280 (N_1280,In_949,In_571);
or U1281 (N_1281,In_675,In_1836);
nand U1282 (N_1282,In_1029,In_78);
and U1283 (N_1283,In_171,In_635);
or U1284 (N_1284,In_1697,In_710);
nor U1285 (N_1285,In_1365,In_143);
nand U1286 (N_1286,In_1378,In_795);
xnor U1287 (N_1287,In_1094,In_944);
or U1288 (N_1288,In_923,In_710);
or U1289 (N_1289,In_1603,In_1192);
nor U1290 (N_1290,In_46,In_1119);
nor U1291 (N_1291,In_750,In_1742);
nand U1292 (N_1292,In_81,In_1543);
and U1293 (N_1293,In_381,In_1687);
xor U1294 (N_1294,In_179,In_1284);
nand U1295 (N_1295,In_509,In_373);
nor U1296 (N_1296,In_518,In_1191);
or U1297 (N_1297,In_935,In_388);
xor U1298 (N_1298,In_1534,In_610);
nor U1299 (N_1299,In_1737,In_1324);
nor U1300 (N_1300,In_1050,In_1325);
or U1301 (N_1301,In_1128,In_626);
xnor U1302 (N_1302,In_1742,In_432);
or U1303 (N_1303,In_1578,In_1727);
nand U1304 (N_1304,In_202,In_378);
nand U1305 (N_1305,In_400,In_44);
or U1306 (N_1306,In_1211,In_499);
and U1307 (N_1307,In_1111,In_1499);
nor U1308 (N_1308,In_1154,In_1218);
or U1309 (N_1309,In_532,In_831);
xnor U1310 (N_1310,In_1036,In_1756);
or U1311 (N_1311,In_1565,In_315);
or U1312 (N_1312,In_842,In_697);
and U1313 (N_1313,In_967,In_296);
and U1314 (N_1314,In_169,In_193);
and U1315 (N_1315,In_1706,In_1225);
and U1316 (N_1316,In_1152,In_651);
nor U1317 (N_1317,In_585,In_1373);
nand U1318 (N_1318,In_63,In_1961);
nand U1319 (N_1319,In_824,In_1968);
and U1320 (N_1320,In_1816,In_1975);
nor U1321 (N_1321,In_238,In_1853);
or U1322 (N_1322,In_872,In_1982);
and U1323 (N_1323,In_1383,In_263);
xnor U1324 (N_1324,In_1490,In_49);
xor U1325 (N_1325,In_679,In_610);
and U1326 (N_1326,In_1389,In_824);
nand U1327 (N_1327,In_1517,In_357);
and U1328 (N_1328,In_287,In_483);
and U1329 (N_1329,In_317,In_1246);
xor U1330 (N_1330,In_1830,In_925);
or U1331 (N_1331,In_678,In_1827);
and U1332 (N_1332,In_1935,In_1153);
and U1333 (N_1333,In_1294,In_261);
and U1334 (N_1334,In_1854,In_479);
xor U1335 (N_1335,In_756,In_746);
xnor U1336 (N_1336,In_1420,In_210);
xor U1337 (N_1337,In_1328,In_1121);
xnor U1338 (N_1338,In_1418,In_1833);
nor U1339 (N_1339,In_1879,In_602);
nand U1340 (N_1340,In_1391,In_1395);
nand U1341 (N_1341,In_1048,In_991);
nor U1342 (N_1342,In_1827,In_1258);
and U1343 (N_1343,In_715,In_647);
xor U1344 (N_1344,In_584,In_1638);
nor U1345 (N_1345,In_1237,In_827);
or U1346 (N_1346,In_194,In_1502);
or U1347 (N_1347,In_745,In_1927);
or U1348 (N_1348,In_1906,In_1478);
xor U1349 (N_1349,In_1586,In_1001);
nand U1350 (N_1350,In_846,In_1046);
xnor U1351 (N_1351,In_1292,In_732);
nor U1352 (N_1352,In_1704,In_84);
nand U1353 (N_1353,In_954,In_1609);
or U1354 (N_1354,In_617,In_1428);
or U1355 (N_1355,In_1053,In_466);
and U1356 (N_1356,In_215,In_599);
or U1357 (N_1357,In_1640,In_1988);
or U1358 (N_1358,In_1850,In_1642);
nor U1359 (N_1359,In_1706,In_1041);
and U1360 (N_1360,In_1830,In_176);
or U1361 (N_1361,In_101,In_1543);
or U1362 (N_1362,In_838,In_1119);
and U1363 (N_1363,In_901,In_528);
nand U1364 (N_1364,In_192,In_1567);
and U1365 (N_1365,In_142,In_1676);
or U1366 (N_1366,In_1568,In_403);
and U1367 (N_1367,In_1418,In_1168);
nor U1368 (N_1368,In_1475,In_215);
nor U1369 (N_1369,In_303,In_565);
and U1370 (N_1370,In_1552,In_507);
xor U1371 (N_1371,In_1211,In_1924);
xnor U1372 (N_1372,In_1254,In_858);
or U1373 (N_1373,In_407,In_467);
xnor U1374 (N_1374,In_494,In_851);
xor U1375 (N_1375,In_1525,In_1227);
nand U1376 (N_1376,In_898,In_1059);
or U1377 (N_1377,In_1526,In_473);
nor U1378 (N_1378,In_1774,In_356);
nor U1379 (N_1379,In_1568,In_1827);
xor U1380 (N_1380,In_675,In_1903);
nor U1381 (N_1381,In_1287,In_338);
and U1382 (N_1382,In_1343,In_955);
and U1383 (N_1383,In_1541,In_1337);
or U1384 (N_1384,In_927,In_1317);
nor U1385 (N_1385,In_362,In_1839);
and U1386 (N_1386,In_1846,In_1788);
xnor U1387 (N_1387,In_1164,In_1249);
xnor U1388 (N_1388,In_1668,In_1925);
xnor U1389 (N_1389,In_939,In_1599);
nor U1390 (N_1390,In_1185,In_231);
or U1391 (N_1391,In_207,In_1772);
nand U1392 (N_1392,In_845,In_1127);
nand U1393 (N_1393,In_1830,In_191);
xnor U1394 (N_1394,In_545,In_442);
or U1395 (N_1395,In_1568,In_957);
or U1396 (N_1396,In_204,In_851);
xnor U1397 (N_1397,In_1602,In_1687);
and U1398 (N_1398,In_1079,In_140);
or U1399 (N_1399,In_1468,In_790);
nand U1400 (N_1400,In_63,In_758);
or U1401 (N_1401,In_793,In_1704);
xor U1402 (N_1402,In_1728,In_1611);
or U1403 (N_1403,In_1058,In_102);
nor U1404 (N_1404,In_1842,In_1185);
nand U1405 (N_1405,In_353,In_1514);
or U1406 (N_1406,In_799,In_1878);
and U1407 (N_1407,In_1419,In_212);
nor U1408 (N_1408,In_1913,In_1045);
nand U1409 (N_1409,In_1906,In_662);
nand U1410 (N_1410,In_1075,In_1552);
and U1411 (N_1411,In_766,In_1092);
and U1412 (N_1412,In_1687,In_1043);
nor U1413 (N_1413,In_431,In_601);
nand U1414 (N_1414,In_897,In_116);
and U1415 (N_1415,In_558,In_424);
and U1416 (N_1416,In_1034,In_325);
xnor U1417 (N_1417,In_1800,In_84);
or U1418 (N_1418,In_1744,In_507);
and U1419 (N_1419,In_1866,In_1357);
or U1420 (N_1420,In_220,In_914);
nand U1421 (N_1421,In_667,In_283);
and U1422 (N_1422,In_1624,In_1054);
xnor U1423 (N_1423,In_704,In_419);
xor U1424 (N_1424,In_1143,In_358);
and U1425 (N_1425,In_1995,In_1767);
nand U1426 (N_1426,In_846,In_1847);
nand U1427 (N_1427,In_54,In_1405);
and U1428 (N_1428,In_1366,In_1705);
xor U1429 (N_1429,In_811,In_655);
and U1430 (N_1430,In_221,In_1645);
and U1431 (N_1431,In_1650,In_1752);
or U1432 (N_1432,In_628,In_1302);
or U1433 (N_1433,In_410,In_1267);
and U1434 (N_1434,In_1912,In_978);
and U1435 (N_1435,In_1993,In_1484);
or U1436 (N_1436,In_1168,In_615);
nor U1437 (N_1437,In_1532,In_842);
and U1438 (N_1438,In_1669,In_530);
nor U1439 (N_1439,In_1505,In_1259);
xor U1440 (N_1440,In_287,In_648);
nand U1441 (N_1441,In_1287,In_224);
xnor U1442 (N_1442,In_1060,In_1382);
nor U1443 (N_1443,In_715,In_749);
or U1444 (N_1444,In_322,In_1633);
nand U1445 (N_1445,In_1395,In_1613);
nand U1446 (N_1446,In_3,In_332);
xnor U1447 (N_1447,In_994,In_1364);
nor U1448 (N_1448,In_1811,In_593);
or U1449 (N_1449,In_1577,In_1908);
nor U1450 (N_1450,In_357,In_431);
or U1451 (N_1451,In_1073,In_534);
nor U1452 (N_1452,In_608,In_1163);
nor U1453 (N_1453,In_948,In_338);
and U1454 (N_1454,In_492,In_792);
or U1455 (N_1455,In_822,In_111);
and U1456 (N_1456,In_175,In_344);
or U1457 (N_1457,In_697,In_1043);
nand U1458 (N_1458,In_1473,In_359);
or U1459 (N_1459,In_786,In_1800);
nand U1460 (N_1460,In_471,In_285);
xor U1461 (N_1461,In_1662,In_1386);
nand U1462 (N_1462,In_1804,In_1403);
or U1463 (N_1463,In_130,In_466);
nand U1464 (N_1464,In_1428,In_244);
xor U1465 (N_1465,In_8,In_1451);
and U1466 (N_1466,In_1914,In_212);
or U1467 (N_1467,In_1660,In_802);
and U1468 (N_1468,In_652,In_420);
xor U1469 (N_1469,In_1816,In_242);
nor U1470 (N_1470,In_1888,In_368);
or U1471 (N_1471,In_1809,In_143);
nor U1472 (N_1472,In_1469,In_1272);
and U1473 (N_1473,In_837,In_328);
or U1474 (N_1474,In_1085,In_1606);
xnor U1475 (N_1475,In_445,In_668);
nor U1476 (N_1476,In_185,In_978);
or U1477 (N_1477,In_1315,In_1638);
or U1478 (N_1478,In_333,In_1852);
and U1479 (N_1479,In_1497,In_1485);
xnor U1480 (N_1480,In_1734,In_1767);
or U1481 (N_1481,In_102,In_221);
and U1482 (N_1482,In_1985,In_1219);
or U1483 (N_1483,In_1410,In_886);
nor U1484 (N_1484,In_149,In_636);
nor U1485 (N_1485,In_553,In_1840);
xor U1486 (N_1486,In_1026,In_1546);
nand U1487 (N_1487,In_1331,In_1421);
xor U1488 (N_1488,In_482,In_1843);
or U1489 (N_1489,In_1265,In_612);
nor U1490 (N_1490,In_266,In_505);
xor U1491 (N_1491,In_713,In_1171);
or U1492 (N_1492,In_1070,In_1342);
or U1493 (N_1493,In_1650,In_1479);
or U1494 (N_1494,In_159,In_843);
xnor U1495 (N_1495,In_1557,In_311);
nor U1496 (N_1496,In_47,In_74);
nor U1497 (N_1497,In_1079,In_1497);
or U1498 (N_1498,In_1483,In_1118);
and U1499 (N_1499,In_723,In_354);
nand U1500 (N_1500,In_1445,In_1227);
nor U1501 (N_1501,In_224,In_973);
nand U1502 (N_1502,In_290,In_1150);
xnor U1503 (N_1503,In_194,In_508);
nor U1504 (N_1504,In_181,In_373);
nor U1505 (N_1505,In_1742,In_1566);
and U1506 (N_1506,In_1551,In_241);
and U1507 (N_1507,In_376,In_1962);
nor U1508 (N_1508,In_756,In_431);
nand U1509 (N_1509,In_395,In_396);
or U1510 (N_1510,In_616,In_1583);
xor U1511 (N_1511,In_1447,In_1498);
and U1512 (N_1512,In_988,In_1750);
xor U1513 (N_1513,In_1483,In_20);
or U1514 (N_1514,In_935,In_1262);
nand U1515 (N_1515,In_617,In_344);
and U1516 (N_1516,In_1687,In_1576);
xor U1517 (N_1517,In_1705,In_740);
and U1518 (N_1518,In_1083,In_1653);
nand U1519 (N_1519,In_994,In_151);
and U1520 (N_1520,In_1219,In_1946);
nand U1521 (N_1521,In_1386,In_1680);
and U1522 (N_1522,In_1929,In_1883);
and U1523 (N_1523,In_88,In_778);
or U1524 (N_1524,In_1353,In_1931);
nor U1525 (N_1525,In_28,In_728);
and U1526 (N_1526,In_1159,In_908);
or U1527 (N_1527,In_221,In_428);
or U1528 (N_1528,In_519,In_1079);
xor U1529 (N_1529,In_1880,In_459);
and U1530 (N_1530,In_1184,In_1303);
and U1531 (N_1531,In_1259,In_223);
xor U1532 (N_1532,In_1210,In_1736);
xor U1533 (N_1533,In_1530,In_628);
and U1534 (N_1534,In_484,In_4);
or U1535 (N_1535,In_896,In_709);
nand U1536 (N_1536,In_1668,In_916);
or U1537 (N_1537,In_1576,In_333);
xor U1538 (N_1538,In_518,In_1385);
and U1539 (N_1539,In_1328,In_777);
and U1540 (N_1540,In_222,In_517);
nor U1541 (N_1541,In_270,In_564);
xnor U1542 (N_1542,In_383,In_1772);
nor U1543 (N_1543,In_1725,In_792);
nor U1544 (N_1544,In_1381,In_750);
nand U1545 (N_1545,In_1836,In_479);
and U1546 (N_1546,In_1455,In_875);
xor U1547 (N_1547,In_756,In_862);
xor U1548 (N_1548,In_612,In_740);
nand U1549 (N_1549,In_1062,In_1686);
nand U1550 (N_1550,In_483,In_1041);
nor U1551 (N_1551,In_1840,In_860);
nand U1552 (N_1552,In_1329,In_1532);
or U1553 (N_1553,In_198,In_1700);
and U1554 (N_1554,In_1069,In_1719);
nand U1555 (N_1555,In_761,In_267);
and U1556 (N_1556,In_1827,In_698);
nand U1557 (N_1557,In_1526,In_1678);
and U1558 (N_1558,In_3,In_138);
or U1559 (N_1559,In_1951,In_828);
xnor U1560 (N_1560,In_1425,In_1498);
or U1561 (N_1561,In_1524,In_1433);
nand U1562 (N_1562,In_603,In_825);
and U1563 (N_1563,In_1722,In_1783);
or U1564 (N_1564,In_445,In_184);
and U1565 (N_1565,In_96,In_25);
nand U1566 (N_1566,In_1679,In_239);
and U1567 (N_1567,In_86,In_1579);
and U1568 (N_1568,In_1056,In_861);
nor U1569 (N_1569,In_32,In_968);
xnor U1570 (N_1570,In_1038,In_1285);
and U1571 (N_1571,In_1012,In_1900);
nand U1572 (N_1572,In_1841,In_324);
nand U1573 (N_1573,In_1763,In_1623);
nor U1574 (N_1574,In_1707,In_913);
or U1575 (N_1575,In_429,In_1789);
nor U1576 (N_1576,In_282,In_1661);
and U1577 (N_1577,In_1435,In_1522);
and U1578 (N_1578,In_1423,In_780);
nand U1579 (N_1579,In_424,In_1506);
or U1580 (N_1580,In_1943,In_1526);
nor U1581 (N_1581,In_1541,In_1175);
xor U1582 (N_1582,In_1625,In_244);
nor U1583 (N_1583,In_797,In_45);
xor U1584 (N_1584,In_1492,In_611);
and U1585 (N_1585,In_185,In_516);
nand U1586 (N_1586,In_345,In_1823);
nand U1587 (N_1587,In_1692,In_444);
nor U1588 (N_1588,In_1785,In_339);
and U1589 (N_1589,In_564,In_664);
and U1590 (N_1590,In_1076,In_1046);
and U1591 (N_1591,In_1069,In_322);
nor U1592 (N_1592,In_1352,In_693);
xor U1593 (N_1593,In_636,In_902);
xnor U1594 (N_1594,In_1192,In_1341);
or U1595 (N_1595,In_1224,In_1100);
xor U1596 (N_1596,In_1262,In_1594);
or U1597 (N_1597,In_1981,In_848);
or U1598 (N_1598,In_316,In_824);
and U1599 (N_1599,In_838,In_1207);
or U1600 (N_1600,In_628,In_1432);
xor U1601 (N_1601,In_1716,In_1435);
and U1602 (N_1602,In_1246,In_1733);
or U1603 (N_1603,In_1210,In_1059);
and U1604 (N_1604,In_1101,In_422);
or U1605 (N_1605,In_1574,In_1647);
xor U1606 (N_1606,In_559,In_1032);
nor U1607 (N_1607,In_1273,In_1155);
or U1608 (N_1608,In_1172,In_1940);
nand U1609 (N_1609,In_1791,In_64);
nand U1610 (N_1610,In_1536,In_37);
or U1611 (N_1611,In_1301,In_1178);
nor U1612 (N_1612,In_59,In_1102);
nand U1613 (N_1613,In_38,In_1131);
xnor U1614 (N_1614,In_1398,In_1792);
xor U1615 (N_1615,In_94,In_511);
nand U1616 (N_1616,In_1014,In_1041);
or U1617 (N_1617,In_1578,In_1415);
and U1618 (N_1618,In_944,In_1482);
or U1619 (N_1619,In_1337,In_29);
nor U1620 (N_1620,In_834,In_340);
nand U1621 (N_1621,In_215,In_670);
nor U1622 (N_1622,In_1440,In_1837);
xnor U1623 (N_1623,In_1919,In_859);
nand U1624 (N_1624,In_1995,In_749);
nor U1625 (N_1625,In_983,In_544);
nor U1626 (N_1626,In_1387,In_133);
and U1627 (N_1627,In_434,In_1940);
or U1628 (N_1628,In_689,In_1820);
nand U1629 (N_1629,In_23,In_1450);
and U1630 (N_1630,In_1041,In_1104);
nand U1631 (N_1631,In_279,In_1886);
nor U1632 (N_1632,In_963,In_1969);
or U1633 (N_1633,In_484,In_1132);
and U1634 (N_1634,In_1540,In_1738);
and U1635 (N_1635,In_1328,In_1129);
xor U1636 (N_1636,In_1560,In_133);
nand U1637 (N_1637,In_147,In_1278);
nand U1638 (N_1638,In_762,In_146);
and U1639 (N_1639,In_491,In_348);
nand U1640 (N_1640,In_867,In_1533);
and U1641 (N_1641,In_406,In_929);
xor U1642 (N_1642,In_1255,In_337);
and U1643 (N_1643,In_616,In_373);
xnor U1644 (N_1644,In_329,In_1608);
or U1645 (N_1645,In_1993,In_212);
or U1646 (N_1646,In_1089,In_614);
and U1647 (N_1647,In_241,In_629);
or U1648 (N_1648,In_484,In_228);
and U1649 (N_1649,In_394,In_1399);
or U1650 (N_1650,In_1599,In_1721);
and U1651 (N_1651,In_1139,In_1276);
or U1652 (N_1652,In_859,In_1946);
and U1653 (N_1653,In_1701,In_578);
and U1654 (N_1654,In_1020,In_661);
nand U1655 (N_1655,In_699,In_1989);
xnor U1656 (N_1656,In_1736,In_271);
nand U1657 (N_1657,In_1188,In_1093);
or U1658 (N_1658,In_497,In_157);
xor U1659 (N_1659,In_714,In_532);
nand U1660 (N_1660,In_673,In_1720);
and U1661 (N_1661,In_1986,In_205);
nor U1662 (N_1662,In_41,In_376);
nor U1663 (N_1663,In_433,In_203);
xor U1664 (N_1664,In_1716,In_625);
xnor U1665 (N_1665,In_1768,In_1378);
nand U1666 (N_1666,In_1451,In_732);
and U1667 (N_1667,In_80,In_375);
nand U1668 (N_1668,In_1210,In_1546);
xor U1669 (N_1669,In_1084,In_922);
nor U1670 (N_1670,In_1336,In_435);
nor U1671 (N_1671,In_1750,In_1870);
nor U1672 (N_1672,In_1924,In_27);
xnor U1673 (N_1673,In_1987,In_1845);
xor U1674 (N_1674,In_1077,In_1035);
or U1675 (N_1675,In_1586,In_179);
nand U1676 (N_1676,In_719,In_113);
nand U1677 (N_1677,In_1756,In_1801);
nand U1678 (N_1678,In_781,In_145);
and U1679 (N_1679,In_932,In_1771);
xnor U1680 (N_1680,In_814,In_1015);
and U1681 (N_1681,In_1765,In_1666);
nand U1682 (N_1682,In_1819,In_1080);
nand U1683 (N_1683,In_308,In_83);
and U1684 (N_1684,In_1076,In_1103);
and U1685 (N_1685,In_681,In_928);
nor U1686 (N_1686,In_1771,In_1209);
or U1687 (N_1687,In_431,In_1832);
nand U1688 (N_1688,In_675,In_1134);
xnor U1689 (N_1689,In_1543,In_541);
nor U1690 (N_1690,In_1699,In_111);
nand U1691 (N_1691,In_109,In_980);
or U1692 (N_1692,In_1,In_681);
or U1693 (N_1693,In_250,In_191);
nand U1694 (N_1694,In_1485,In_1054);
and U1695 (N_1695,In_1763,In_1794);
or U1696 (N_1696,In_983,In_1354);
nand U1697 (N_1697,In_965,In_879);
xnor U1698 (N_1698,In_685,In_793);
nor U1699 (N_1699,In_631,In_961);
xor U1700 (N_1700,In_1552,In_561);
or U1701 (N_1701,In_646,In_288);
nor U1702 (N_1702,In_1766,In_632);
and U1703 (N_1703,In_1623,In_157);
xor U1704 (N_1704,In_1651,In_1554);
xnor U1705 (N_1705,In_1359,In_1936);
xnor U1706 (N_1706,In_1341,In_723);
or U1707 (N_1707,In_1170,In_96);
or U1708 (N_1708,In_803,In_1822);
nand U1709 (N_1709,In_1140,In_1938);
xnor U1710 (N_1710,In_1445,In_920);
xor U1711 (N_1711,In_585,In_1043);
nand U1712 (N_1712,In_328,In_318);
nor U1713 (N_1713,In_1987,In_1288);
nor U1714 (N_1714,In_583,In_1499);
xnor U1715 (N_1715,In_676,In_1631);
and U1716 (N_1716,In_1,In_525);
and U1717 (N_1717,In_975,In_1352);
nor U1718 (N_1718,In_845,In_1436);
xor U1719 (N_1719,In_1222,In_1297);
xor U1720 (N_1720,In_96,In_1095);
and U1721 (N_1721,In_1094,In_1758);
nor U1722 (N_1722,In_28,In_1087);
xnor U1723 (N_1723,In_83,In_835);
and U1724 (N_1724,In_555,In_203);
nor U1725 (N_1725,In_623,In_785);
and U1726 (N_1726,In_391,In_1457);
or U1727 (N_1727,In_783,In_220);
xor U1728 (N_1728,In_99,In_1682);
nand U1729 (N_1729,In_857,In_0);
or U1730 (N_1730,In_777,In_1233);
or U1731 (N_1731,In_249,In_1085);
nor U1732 (N_1732,In_437,In_1673);
xnor U1733 (N_1733,In_1499,In_1626);
or U1734 (N_1734,In_801,In_1561);
and U1735 (N_1735,In_785,In_698);
nor U1736 (N_1736,In_1187,In_852);
and U1737 (N_1737,In_137,In_1614);
xor U1738 (N_1738,In_413,In_874);
and U1739 (N_1739,In_82,In_1691);
or U1740 (N_1740,In_1321,In_1253);
xor U1741 (N_1741,In_1663,In_1103);
and U1742 (N_1742,In_1087,In_1826);
and U1743 (N_1743,In_1417,In_716);
or U1744 (N_1744,In_928,In_1444);
and U1745 (N_1745,In_555,In_1942);
nand U1746 (N_1746,In_25,In_1614);
xor U1747 (N_1747,In_1280,In_1384);
nand U1748 (N_1748,In_1649,In_1413);
xor U1749 (N_1749,In_1967,In_578);
nand U1750 (N_1750,In_231,In_1998);
xnor U1751 (N_1751,In_1122,In_951);
and U1752 (N_1752,In_1515,In_612);
or U1753 (N_1753,In_735,In_154);
or U1754 (N_1754,In_958,In_1098);
nand U1755 (N_1755,In_442,In_956);
xnor U1756 (N_1756,In_1727,In_1460);
nor U1757 (N_1757,In_733,In_877);
xnor U1758 (N_1758,In_1868,In_1864);
and U1759 (N_1759,In_1848,In_1765);
or U1760 (N_1760,In_1254,In_319);
xor U1761 (N_1761,In_900,In_1917);
nand U1762 (N_1762,In_1555,In_894);
nor U1763 (N_1763,In_1466,In_555);
nand U1764 (N_1764,In_1911,In_1916);
nor U1765 (N_1765,In_1613,In_1922);
or U1766 (N_1766,In_860,In_1124);
and U1767 (N_1767,In_81,In_1814);
and U1768 (N_1768,In_1580,In_515);
and U1769 (N_1769,In_747,In_41);
and U1770 (N_1770,In_425,In_1306);
or U1771 (N_1771,In_286,In_82);
nand U1772 (N_1772,In_757,In_1318);
or U1773 (N_1773,In_315,In_616);
xnor U1774 (N_1774,In_867,In_1882);
and U1775 (N_1775,In_1269,In_51);
nand U1776 (N_1776,In_1120,In_1760);
and U1777 (N_1777,In_1662,In_343);
xor U1778 (N_1778,In_1028,In_1933);
xor U1779 (N_1779,In_1871,In_893);
nor U1780 (N_1780,In_1656,In_276);
and U1781 (N_1781,In_327,In_1331);
nand U1782 (N_1782,In_1408,In_1677);
or U1783 (N_1783,In_954,In_348);
nor U1784 (N_1784,In_1560,In_1431);
xor U1785 (N_1785,In_1792,In_1752);
nor U1786 (N_1786,In_1209,In_1024);
and U1787 (N_1787,In_805,In_125);
and U1788 (N_1788,In_172,In_1970);
xnor U1789 (N_1789,In_1039,In_143);
xor U1790 (N_1790,In_1433,In_1655);
or U1791 (N_1791,In_19,In_1826);
nor U1792 (N_1792,In_1114,In_837);
nor U1793 (N_1793,In_941,In_252);
nand U1794 (N_1794,In_579,In_1485);
nor U1795 (N_1795,In_957,In_1445);
xnor U1796 (N_1796,In_318,In_44);
or U1797 (N_1797,In_1013,In_405);
or U1798 (N_1798,In_1032,In_184);
or U1799 (N_1799,In_277,In_737);
or U1800 (N_1800,In_948,In_618);
nand U1801 (N_1801,In_994,In_1081);
nor U1802 (N_1802,In_170,In_856);
or U1803 (N_1803,In_816,In_973);
nand U1804 (N_1804,In_299,In_1519);
nor U1805 (N_1805,In_437,In_1282);
and U1806 (N_1806,In_49,In_1745);
xor U1807 (N_1807,In_195,In_1073);
and U1808 (N_1808,In_1721,In_1737);
xnor U1809 (N_1809,In_454,In_585);
nand U1810 (N_1810,In_1862,In_898);
nor U1811 (N_1811,In_1124,In_1457);
nand U1812 (N_1812,In_745,In_503);
nand U1813 (N_1813,In_298,In_572);
or U1814 (N_1814,In_1838,In_21);
nand U1815 (N_1815,In_1203,In_836);
nand U1816 (N_1816,In_71,In_943);
or U1817 (N_1817,In_410,In_854);
nand U1818 (N_1818,In_674,In_1590);
or U1819 (N_1819,In_1133,In_1388);
or U1820 (N_1820,In_1187,In_143);
nor U1821 (N_1821,In_1734,In_618);
or U1822 (N_1822,In_1830,In_1080);
xor U1823 (N_1823,In_1136,In_299);
nand U1824 (N_1824,In_1344,In_1355);
xor U1825 (N_1825,In_597,In_181);
nand U1826 (N_1826,In_1055,In_1406);
nand U1827 (N_1827,In_658,In_659);
nor U1828 (N_1828,In_627,In_408);
nor U1829 (N_1829,In_1167,In_146);
and U1830 (N_1830,In_1490,In_1719);
xnor U1831 (N_1831,In_6,In_1120);
xor U1832 (N_1832,In_1327,In_1306);
nor U1833 (N_1833,In_1906,In_1050);
xor U1834 (N_1834,In_143,In_1222);
nor U1835 (N_1835,In_584,In_155);
nor U1836 (N_1836,In_702,In_1314);
xor U1837 (N_1837,In_965,In_1515);
nand U1838 (N_1838,In_144,In_521);
xor U1839 (N_1839,In_1532,In_44);
nand U1840 (N_1840,In_1397,In_1926);
nor U1841 (N_1841,In_1325,In_863);
or U1842 (N_1842,In_1609,In_1165);
xnor U1843 (N_1843,In_1117,In_281);
xor U1844 (N_1844,In_468,In_1511);
nand U1845 (N_1845,In_1237,In_302);
and U1846 (N_1846,In_1388,In_1966);
and U1847 (N_1847,In_1403,In_1021);
nor U1848 (N_1848,In_748,In_474);
xnor U1849 (N_1849,In_1968,In_146);
nor U1850 (N_1850,In_1296,In_1637);
nor U1851 (N_1851,In_1146,In_773);
nand U1852 (N_1852,In_305,In_194);
and U1853 (N_1853,In_1320,In_1147);
and U1854 (N_1854,In_723,In_353);
nor U1855 (N_1855,In_1461,In_13);
nand U1856 (N_1856,In_1670,In_480);
xor U1857 (N_1857,In_488,In_341);
nand U1858 (N_1858,In_1661,In_647);
nor U1859 (N_1859,In_904,In_1379);
or U1860 (N_1860,In_1627,In_1610);
or U1861 (N_1861,In_1079,In_1887);
or U1862 (N_1862,In_826,In_936);
nand U1863 (N_1863,In_1235,In_816);
and U1864 (N_1864,In_281,In_1916);
xor U1865 (N_1865,In_31,In_310);
nand U1866 (N_1866,In_1964,In_1971);
xnor U1867 (N_1867,In_1907,In_348);
nor U1868 (N_1868,In_1369,In_931);
xnor U1869 (N_1869,In_267,In_1898);
and U1870 (N_1870,In_1970,In_826);
nor U1871 (N_1871,In_1880,In_1876);
or U1872 (N_1872,In_1982,In_982);
or U1873 (N_1873,In_1275,In_853);
and U1874 (N_1874,In_1551,In_844);
nor U1875 (N_1875,In_54,In_1585);
nand U1876 (N_1876,In_889,In_195);
and U1877 (N_1877,In_1680,In_1172);
or U1878 (N_1878,In_1170,In_1706);
or U1879 (N_1879,In_251,In_1577);
nand U1880 (N_1880,In_1932,In_894);
nor U1881 (N_1881,In_1015,In_677);
xnor U1882 (N_1882,In_1338,In_476);
nand U1883 (N_1883,In_1824,In_245);
nor U1884 (N_1884,In_781,In_1316);
and U1885 (N_1885,In_505,In_490);
or U1886 (N_1886,In_1766,In_148);
or U1887 (N_1887,In_188,In_153);
xor U1888 (N_1888,In_1834,In_1604);
xnor U1889 (N_1889,In_1613,In_1385);
nor U1890 (N_1890,In_363,In_1111);
xnor U1891 (N_1891,In_172,In_150);
or U1892 (N_1892,In_86,In_192);
or U1893 (N_1893,In_1840,In_288);
and U1894 (N_1894,In_980,In_140);
nand U1895 (N_1895,In_696,In_385);
xor U1896 (N_1896,In_1621,In_634);
or U1897 (N_1897,In_916,In_1300);
and U1898 (N_1898,In_1989,In_1131);
or U1899 (N_1899,In_835,In_1367);
and U1900 (N_1900,In_1495,In_1767);
or U1901 (N_1901,In_1206,In_113);
nand U1902 (N_1902,In_1225,In_1462);
nor U1903 (N_1903,In_518,In_607);
or U1904 (N_1904,In_812,In_669);
xnor U1905 (N_1905,In_671,In_1682);
nor U1906 (N_1906,In_1480,In_271);
nand U1907 (N_1907,In_1163,In_460);
xnor U1908 (N_1908,In_257,In_432);
nand U1909 (N_1909,In_607,In_1289);
xor U1910 (N_1910,In_1672,In_544);
xor U1911 (N_1911,In_1715,In_634);
nand U1912 (N_1912,In_1915,In_1067);
or U1913 (N_1913,In_797,In_260);
nand U1914 (N_1914,In_1757,In_1893);
and U1915 (N_1915,In_545,In_1142);
nor U1916 (N_1916,In_1489,In_828);
xnor U1917 (N_1917,In_1097,In_1938);
and U1918 (N_1918,In_1244,In_227);
nor U1919 (N_1919,In_1696,In_1096);
and U1920 (N_1920,In_711,In_1023);
xor U1921 (N_1921,In_278,In_1213);
nand U1922 (N_1922,In_358,In_937);
or U1923 (N_1923,In_1584,In_1066);
or U1924 (N_1924,In_1750,In_809);
and U1925 (N_1925,In_1126,In_95);
and U1926 (N_1926,In_156,In_1871);
or U1927 (N_1927,In_1875,In_859);
and U1928 (N_1928,In_1990,In_1349);
or U1929 (N_1929,In_58,In_1509);
nor U1930 (N_1930,In_49,In_1262);
or U1931 (N_1931,In_1666,In_1239);
nand U1932 (N_1932,In_1338,In_236);
xnor U1933 (N_1933,In_1688,In_108);
xor U1934 (N_1934,In_1673,In_1360);
nand U1935 (N_1935,In_739,In_70);
nor U1936 (N_1936,In_1438,In_1674);
nand U1937 (N_1937,In_1073,In_1097);
nand U1938 (N_1938,In_318,In_1084);
xnor U1939 (N_1939,In_404,In_1360);
and U1940 (N_1940,In_1640,In_43);
and U1941 (N_1941,In_1848,In_362);
or U1942 (N_1942,In_1335,In_376);
nand U1943 (N_1943,In_1438,In_1282);
and U1944 (N_1944,In_1925,In_1557);
or U1945 (N_1945,In_1509,In_763);
nor U1946 (N_1946,In_603,In_1000);
xor U1947 (N_1947,In_808,In_679);
nor U1948 (N_1948,In_1772,In_255);
nand U1949 (N_1949,In_1068,In_144);
nor U1950 (N_1950,In_639,In_1466);
nor U1951 (N_1951,In_1301,In_1699);
xnor U1952 (N_1952,In_1844,In_1874);
nand U1953 (N_1953,In_1744,In_332);
nand U1954 (N_1954,In_7,In_1607);
nand U1955 (N_1955,In_1403,In_1437);
nand U1956 (N_1956,In_1158,In_752);
nand U1957 (N_1957,In_206,In_1729);
nor U1958 (N_1958,In_1749,In_36);
nand U1959 (N_1959,In_1354,In_214);
nor U1960 (N_1960,In_1201,In_387);
nor U1961 (N_1961,In_34,In_686);
or U1962 (N_1962,In_502,In_1391);
or U1963 (N_1963,In_1413,In_1014);
and U1964 (N_1964,In_1507,In_726);
or U1965 (N_1965,In_986,In_1382);
nand U1966 (N_1966,In_174,In_1700);
nand U1967 (N_1967,In_266,In_715);
and U1968 (N_1968,In_1693,In_1704);
xnor U1969 (N_1969,In_773,In_1582);
nor U1970 (N_1970,In_1360,In_1945);
and U1971 (N_1971,In_1399,In_1587);
xor U1972 (N_1972,In_108,In_1611);
nand U1973 (N_1973,In_50,In_432);
and U1974 (N_1974,In_1398,In_1236);
or U1975 (N_1975,In_581,In_1599);
and U1976 (N_1976,In_1114,In_901);
xor U1977 (N_1977,In_616,In_410);
nand U1978 (N_1978,In_415,In_1416);
xor U1979 (N_1979,In_521,In_1222);
xnor U1980 (N_1980,In_48,In_258);
nor U1981 (N_1981,In_1704,In_1585);
xnor U1982 (N_1982,In_220,In_400);
or U1983 (N_1983,In_114,In_1288);
or U1984 (N_1984,In_1458,In_462);
nor U1985 (N_1985,In_59,In_1436);
nand U1986 (N_1986,In_410,In_1625);
nand U1987 (N_1987,In_195,In_1318);
nor U1988 (N_1988,In_650,In_1427);
nor U1989 (N_1989,In_1622,In_1841);
xnor U1990 (N_1990,In_107,In_1818);
or U1991 (N_1991,In_1839,In_1786);
nor U1992 (N_1992,In_862,In_1473);
nand U1993 (N_1993,In_1771,In_876);
or U1994 (N_1994,In_953,In_1982);
nor U1995 (N_1995,In_1521,In_982);
and U1996 (N_1996,In_784,In_1513);
nand U1997 (N_1997,In_1380,In_536);
or U1998 (N_1998,In_850,In_747);
and U1999 (N_1999,In_725,In_149);
or U2000 (N_2000,In_1263,In_611);
nor U2001 (N_2001,In_839,In_129);
and U2002 (N_2002,In_363,In_1769);
nor U2003 (N_2003,In_836,In_102);
nor U2004 (N_2004,In_1557,In_1240);
and U2005 (N_2005,In_1054,In_612);
nand U2006 (N_2006,In_171,In_1404);
or U2007 (N_2007,In_289,In_721);
or U2008 (N_2008,In_818,In_1539);
and U2009 (N_2009,In_1930,In_1851);
nor U2010 (N_2010,In_815,In_1156);
and U2011 (N_2011,In_1436,In_1597);
nand U2012 (N_2012,In_646,In_1083);
nor U2013 (N_2013,In_1591,In_916);
xnor U2014 (N_2014,In_71,In_1872);
or U2015 (N_2015,In_1856,In_1272);
or U2016 (N_2016,In_1336,In_655);
or U2017 (N_2017,In_90,In_1527);
or U2018 (N_2018,In_1284,In_1630);
xnor U2019 (N_2019,In_26,In_1777);
xnor U2020 (N_2020,In_1742,In_483);
nor U2021 (N_2021,In_1788,In_1980);
nor U2022 (N_2022,In_460,In_1373);
xnor U2023 (N_2023,In_136,In_687);
nor U2024 (N_2024,In_1791,In_763);
xnor U2025 (N_2025,In_777,In_778);
or U2026 (N_2026,In_37,In_1336);
or U2027 (N_2027,In_1746,In_1895);
or U2028 (N_2028,In_536,In_1410);
nand U2029 (N_2029,In_368,In_200);
xor U2030 (N_2030,In_1737,In_1352);
nor U2031 (N_2031,In_869,In_843);
and U2032 (N_2032,In_226,In_1926);
or U2033 (N_2033,In_12,In_1109);
nand U2034 (N_2034,In_1567,In_1446);
nor U2035 (N_2035,In_473,In_1361);
xor U2036 (N_2036,In_201,In_1583);
xor U2037 (N_2037,In_1897,In_1516);
xnor U2038 (N_2038,In_67,In_1022);
nand U2039 (N_2039,In_1045,In_1287);
nor U2040 (N_2040,In_420,In_264);
nand U2041 (N_2041,In_1928,In_758);
and U2042 (N_2042,In_1151,In_1756);
and U2043 (N_2043,In_226,In_222);
and U2044 (N_2044,In_157,In_328);
and U2045 (N_2045,In_193,In_1543);
nand U2046 (N_2046,In_845,In_1027);
and U2047 (N_2047,In_1135,In_650);
nor U2048 (N_2048,In_228,In_196);
and U2049 (N_2049,In_503,In_432);
and U2050 (N_2050,In_57,In_1549);
and U2051 (N_2051,In_626,In_477);
nand U2052 (N_2052,In_1092,In_950);
xnor U2053 (N_2053,In_1304,In_663);
nor U2054 (N_2054,In_1531,In_1827);
xnor U2055 (N_2055,In_356,In_385);
nor U2056 (N_2056,In_328,In_885);
xnor U2057 (N_2057,In_856,In_517);
and U2058 (N_2058,In_452,In_1774);
and U2059 (N_2059,In_1134,In_1528);
and U2060 (N_2060,In_253,In_1263);
xnor U2061 (N_2061,In_1122,In_975);
nand U2062 (N_2062,In_1038,In_1613);
and U2063 (N_2063,In_1212,In_1513);
or U2064 (N_2064,In_693,In_249);
nor U2065 (N_2065,In_518,In_1289);
xor U2066 (N_2066,In_1249,In_1974);
xor U2067 (N_2067,In_1460,In_1323);
xor U2068 (N_2068,In_102,In_814);
xnor U2069 (N_2069,In_1270,In_364);
or U2070 (N_2070,In_611,In_1467);
or U2071 (N_2071,In_1038,In_1828);
or U2072 (N_2072,In_1618,In_1779);
and U2073 (N_2073,In_1181,In_1610);
nand U2074 (N_2074,In_1750,In_1964);
xor U2075 (N_2075,In_398,In_322);
xnor U2076 (N_2076,In_1009,In_3);
xor U2077 (N_2077,In_1656,In_1002);
xnor U2078 (N_2078,In_621,In_1943);
nor U2079 (N_2079,In_200,In_1440);
nor U2080 (N_2080,In_1166,In_1314);
or U2081 (N_2081,In_183,In_725);
nand U2082 (N_2082,In_1391,In_1896);
nand U2083 (N_2083,In_1992,In_1477);
or U2084 (N_2084,In_1974,In_1609);
xor U2085 (N_2085,In_1918,In_172);
or U2086 (N_2086,In_735,In_1645);
xnor U2087 (N_2087,In_1860,In_979);
and U2088 (N_2088,In_1011,In_194);
xor U2089 (N_2089,In_1195,In_1440);
and U2090 (N_2090,In_276,In_824);
and U2091 (N_2091,In_865,In_1221);
or U2092 (N_2092,In_1218,In_1293);
nor U2093 (N_2093,In_1748,In_488);
nor U2094 (N_2094,In_177,In_1049);
nor U2095 (N_2095,In_1410,In_695);
and U2096 (N_2096,In_1366,In_511);
nand U2097 (N_2097,In_1312,In_36);
or U2098 (N_2098,In_635,In_1084);
or U2099 (N_2099,In_83,In_1794);
nand U2100 (N_2100,In_34,In_1250);
xnor U2101 (N_2101,In_1614,In_385);
nor U2102 (N_2102,In_1353,In_1907);
and U2103 (N_2103,In_1154,In_97);
xor U2104 (N_2104,In_660,In_1093);
xor U2105 (N_2105,In_1716,In_862);
nand U2106 (N_2106,In_233,In_1193);
xor U2107 (N_2107,In_610,In_153);
or U2108 (N_2108,In_801,In_436);
and U2109 (N_2109,In_363,In_77);
and U2110 (N_2110,In_2,In_190);
nor U2111 (N_2111,In_588,In_806);
and U2112 (N_2112,In_1106,In_672);
and U2113 (N_2113,In_1182,In_373);
or U2114 (N_2114,In_1781,In_170);
and U2115 (N_2115,In_691,In_932);
and U2116 (N_2116,In_658,In_1900);
nand U2117 (N_2117,In_1400,In_1451);
nor U2118 (N_2118,In_560,In_587);
nor U2119 (N_2119,In_406,In_49);
or U2120 (N_2120,In_675,In_1471);
or U2121 (N_2121,In_1876,In_1530);
xnor U2122 (N_2122,In_298,In_711);
and U2123 (N_2123,In_1160,In_845);
and U2124 (N_2124,In_540,In_1707);
xor U2125 (N_2125,In_941,In_1878);
xor U2126 (N_2126,In_614,In_832);
and U2127 (N_2127,In_1076,In_590);
and U2128 (N_2128,In_1613,In_1608);
xnor U2129 (N_2129,In_1316,In_1124);
or U2130 (N_2130,In_1762,In_1691);
or U2131 (N_2131,In_1020,In_1866);
nor U2132 (N_2132,In_581,In_946);
xnor U2133 (N_2133,In_290,In_1506);
and U2134 (N_2134,In_1348,In_1780);
xnor U2135 (N_2135,In_1148,In_1678);
nor U2136 (N_2136,In_615,In_443);
xor U2137 (N_2137,In_114,In_1903);
and U2138 (N_2138,In_622,In_1691);
xnor U2139 (N_2139,In_1656,In_267);
and U2140 (N_2140,In_92,In_69);
and U2141 (N_2141,In_1952,In_88);
xor U2142 (N_2142,In_1034,In_1450);
or U2143 (N_2143,In_63,In_639);
nand U2144 (N_2144,In_1670,In_377);
nand U2145 (N_2145,In_26,In_1368);
nor U2146 (N_2146,In_572,In_831);
xor U2147 (N_2147,In_744,In_474);
or U2148 (N_2148,In_97,In_1839);
nor U2149 (N_2149,In_1248,In_334);
nand U2150 (N_2150,In_430,In_452);
and U2151 (N_2151,In_1655,In_1178);
and U2152 (N_2152,In_1308,In_933);
or U2153 (N_2153,In_187,In_1372);
and U2154 (N_2154,In_556,In_237);
nor U2155 (N_2155,In_1794,In_1948);
nand U2156 (N_2156,In_731,In_919);
nor U2157 (N_2157,In_469,In_393);
and U2158 (N_2158,In_910,In_476);
nor U2159 (N_2159,In_860,In_1026);
and U2160 (N_2160,In_1069,In_785);
nor U2161 (N_2161,In_361,In_144);
or U2162 (N_2162,In_1417,In_1565);
nor U2163 (N_2163,In_1306,In_1467);
nor U2164 (N_2164,In_1069,In_653);
xnor U2165 (N_2165,In_839,In_1721);
or U2166 (N_2166,In_1458,In_1391);
and U2167 (N_2167,In_289,In_251);
nand U2168 (N_2168,In_436,In_479);
nor U2169 (N_2169,In_1458,In_449);
or U2170 (N_2170,In_1202,In_1456);
and U2171 (N_2171,In_1719,In_538);
nand U2172 (N_2172,In_246,In_1325);
xor U2173 (N_2173,In_1291,In_271);
nor U2174 (N_2174,In_920,In_776);
or U2175 (N_2175,In_1690,In_995);
xor U2176 (N_2176,In_1812,In_738);
and U2177 (N_2177,In_270,In_927);
and U2178 (N_2178,In_1852,In_1701);
xnor U2179 (N_2179,In_832,In_571);
nand U2180 (N_2180,In_1027,In_442);
nor U2181 (N_2181,In_429,In_430);
xnor U2182 (N_2182,In_759,In_699);
nand U2183 (N_2183,In_1569,In_886);
or U2184 (N_2184,In_1587,In_628);
or U2185 (N_2185,In_88,In_953);
and U2186 (N_2186,In_71,In_1291);
and U2187 (N_2187,In_1456,In_1223);
nand U2188 (N_2188,In_402,In_4);
nand U2189 (N_2189,In_1699,In_422);
and U2190 (N_2190,In_546,In_1480);
nor U2191 (N_2191,In_367,In_647);
or U2192 (N_2192,In_590,In_861);
and U2193 (N_2193,In_1987,In_1146);
nor U2194 (N_2194,In_339,In_1078);
xnor U2195 (N_2195,In_1305,In_1422);
nand U2196 (N_2196,In_578,In_79);
and U2197 (N_2197,In_1329,In_985);
and U2198 (N_2198,In_647,In_1408);
or U2199 (N_2199,In_699,In_1669);
nand U2200 (N_2200,In_385,In_100);
and U2201 (N_2201,In_1279,In_481);
and U2202 (N_2202,In_1700,In_1032);
xnor U2203 (N_2203,In_1363,In_738);
xor U2204 (N_2204,In_1714,In_301);
nor U2205 (N_2205,In_1110,In_1580);
nor U2206 (N_2206,In_1876,In_1757);
xnor U2207 (N_2207,In_24,In_910);
or U2208 (N_2208,In_269,In_372);
nor U2209 (N_2209,In_1607,In_1536);
xnor U2210 (N_2210,In_1230,In_1333);
nor U2211 (N_2211,In_1817,In_64);
nand U2212 (N_2212,In_1787,In_554);
or U2213 (N_2213,In_191,In_674);
xnor U2214 (N_2214,In_464,In_1622);
nor U2215 (N_2215,In_1342,In_403);
and U2216 (N_2216,In_535,In_850);
nand U2217 (N_2217,In_438,In_1392);
xnor U2218 (N_2218,In_1145,In_369);
nand U2219 (N_2219,In_1565,In_625);
or U2220 (N_2220,In_864,In_1496);
or U2221 (N_2221,In_1070,In_588);
or U2222 (N_2222,In_246,In_230);
nand U2223 (N_2223,In_1349,In_1434);
xor U2224 (N_2224,In_692,In_346);
nand U2225 (N_2225,In_1885,In_201);
xor U2226 (N_2226,In_683,In_342);
nand U2227 (N_2227,In_857,In_875);
nand U2228 (N_2228,In_1785,In_1997);
xnor U2229 (N_2229,In_1723,In_971);
nor U2230 (N_2230,In_468,In_1684);
and U2231 (N_2231,In_1446,In_85);
nand U2232 (N_2232,In_252,In_709);
or U2233 (N_2233,In_819,In_503);
nor U2234 (N_2234,In_485,In_346);
and U2235 (N_2235,In_400,In_374);
or U2236 (N_2236,In_1476,In_1364);
and U2237 (N_2237,In_1463,In_1581);
xor U2238 (N_2238,In_915,In_1764);
and U2239 (N_2239,In_1972,In_762);
or U2240 (N_2240,In_59,In_1154);
or U2241 (N_2241,In_959,In_317);
and U2242 (N_2242,In_1348,In_571);
xor U2243 (N_2243,In_564,In_309);
or U2244 (N_2244,In_1799,In_1254);
xnor U2245 (N_2245,In_1081,In_1284);
and U2246 (N_2246,In_1124,In_403);
and U2247 (N_2247,In_146,In_1662);
nand U2248 (N_2248,In_1108,In_822);
nor U2249 (N_2249,In_1623,In_1860);
or U2250 (N_2250,In_1464,In_859);
xnor U2251 (N_2251,In_1442,In_12);
or U2252 (N_2252,In_1492,In_1389);
and U2253 (N_2253,In_1249,In_1368);
xnor U2254 (N_2254,In_1347,In_1229);
nor U2255 (N_2255,In_1081,In_1339);
or U2256 (N_2256,In_353,In_1651);
nor U2257 (N_2257,In_354,In_1513);
and U2258 (N_2258,In_191,In_1973);
nand U2259 (N_2259,In_1448,In_1776);
xnor U2260 (N_2260,In_78,In_149);
nand U2261 (N_2261,In_1543,In_1810);
and U2262 (N_2262,In_853,In_1115);
nor U2263 (N_2263,In_1477,In_1298);
xnor U2264 (N_2264,In_1115,In_1140);
or U2265 (N_2265,In_1896,In_1439);
nor U2266 (N_2266,In_1049,In_397);
or U2267 (N_2267,In_283,In_527);
xor U2268 (N_2268,In_1401,In_602);
xnor U2269 (N_2269,In_1907,In_1477);
xor U2270 (N_2270,In_3,In_50);
or U2271 (N_2271,In_1787,In_373);
and U2272 (N_2272,In_1255,In_268);
nand U2273 (N_2273,In_824,In_632);
or U2274 (N_2274,In_254,In_1883);
nand U2275 (N_2275,In_983,In_1515);
xor U2276 (N_2276,In_1488,In_314);
xor U2277 (N_2277,In_1427,In_1082);
and U2278 (N_2278,In_1146,In_847);
xor U2279 (N_2279,In_437,In_1154);
and U2280 (N_2280,In_52,In_1415);
nor U2281 (N_2281,In_1065,In_311);
nor U2282 (N_2282,In_1517,In_1885);
or U2283 (N_2283,In_1628,In_735);
nand U2284 (N_2284,In_1990,In_1476);
nor U2285 (N_2285,In_322,In_1248);
xnor U2286 (N_2286,In_214,In_131);
and U2287 (N_2287,In_1506,In_814);
nand U2288 (N_2288,In_461,In_48);
xnor U2289 (N_2289,In_383,In_87);
xor U2290 (N_2290,In_659,In_1587);
nand U2291 (N_2291,In_1766,In_1429);
and U2292 (N_2292,In_1777,In_1264);
nand U2293 (N_2293,In_1968,In_1927);
or U2294 (N_2294,In_1119,In_1215);
and U2295 (N_2295,In_78,In_1162);
nor U2296 (N_2296,In_876,In_1562);
nand U2297 (N_2297,In_1846,In_1938);
nand U2298 (N_2298,In_1590,In_1078);
xor U2299 (N_2299,In_1684,In_1351);
xor U2300 (N_2300,In_565,In_56);
and U2301 (N_2301,In_1519,In_767);
nor U2302 (N_2302,In_614,In_548);
or U2303 (N_2303,In_940,In_965);
xnor U2304 (N_2304,In_82,In_751);
or U2305 (N_2305,In_1812,In_829);
or U2306 (N_2306,In_252,In_831);
nand U2307 (N_2307,In_851,In_1423);
xor U2308 (N_2308,In_1381,In_1528);
and U2309 (N_2309,In_446,In_472);
and U2310 (N_2310,In_1471,In_1617);
and U2311 (N_2311,In_9,In_642);
nor U2312 (N_2312,In_1169,In_837);
xor U2313 (N_2313,In_1256,In_1556);
nand U2314 (N_2314,In_1445,In_1340);
or U2315 (N_2315,In_1028,In_1730);
nor U2316 (N_2316,In_1808,In_200);
xnor U2317 (N_2317,In_548,In_1794);
and U2318 (N_2318,In_938,In_89);
xor U2319 (N_2319,In_946,In_1799);
nor U2320 (N_2320,In_1011,In_808);
xor U2321 (N_2321,In_1623,In_663);
or U2322 (N_2322,In_150,In_88);
xor U2323 (N_2323,In_438,In_182);
xor U2324 (N_2324,In_205,In_1481);
and U2325 (N_2325,In_590,In_1573);
nand U2326 (N_2326,In_395,In_840);
nor U2327 (N_2327,In_725,In_1260);
xnor U2328 (N_2328,In_1417,In_1574);
and U2329 (N_2329,In_914,In_427);
and U2330 (N_2330,In_1283,In_1430);
or U2331 (N_2331,In_242,In_1216);
nand U2332 (N_2332,In_1435,In_1301);
and U2333 (N_2333,In_482,In_1678);
nand U2334 (N_2334,In_1395,In_1192);
and U2335 (N_2335,In_1712,In_469);
nor U2336 (N_2336,In_993,In_1384);
xnor U2337 (N_2337,In_680,In_370);
or U2338 (N_2338,In_476,In_127);
nand U2339 (N_2339,In_644,In_159);
nor U2340 (N_2340,In_538,In_1239);
nor U2341 (N_2341,In_1265,In_1310);
and U2342 (N_2342,In_711,In_1506);
nand U2343 (N_2343,In_961,In_1598);
or U2344 (N_2344,In_261,In_1384);
nor U2345 (N_2345,In_339,In_1289);
nor U2346 (N_2346,In_1540,In_1533);
xor U2347 (N_2347,In_858,In_332);
nor U2348 (N_2348,In_119,In_8);
nor U2349 (N_2349,In_500,In_1711);
or U2350 (N_2350,In_225,In_559);
xnor U2351 (N_2351,In_1464,In_470);
nor U2352 (N_2352,In_1116,In_270);
nor U2353 (N_2353,In_92,In_1849);
xnor U2354 (N_2354,In_752,In_1176);
nor U2355 (N_2355,In_573,In_154);
and U2356 (N_2356,In_839,In_1524);
nor U2357 (N_2357,In_110,In_347);
xnor U2358 (N_2358,In_505,In_1759);
nand U2359 (N_2359,In_300,In_233);
xnor U2360 (N_2360,In_1489,In_1265);
xor U2361 (N_2361,In_670,In_1096);
nand U2362 (N_2362,In_495,In_180);
or U2363 (N_2363,In_722,In_1980);
nor U2364 (N_2364,In_1793,In_1384);
nor U2365 (N_2365,In_1747,In_152);
and U2366 (N_2366,In_565,In_304);
and U2367 (N_2367,In_1399,In_1533);
and U2368 (N_2368,In_1337,In_147);
or U2369 (N_2369,In_397,In_610);
and U2370 (N_2370,In_594,In_1902);
and U2371 (N_2371,In_820,In_1420);
nand U2372 (N_2372,In_766,In_1813);
nand U2373 (N_2373,In_1019,In_1702);
and U2374 (N_2374,In_588,In_1712);
nand U2375 (N_2375,In_491,In_433);
and U2376 (N_2376,In_1623,In_1939);
xor U2377 (N_2377,In_815,In_1667);
xnor U2378 (N_2378,In_1618,In_1292);
nor U2379 (N_2379,In_403,In_1837);
xnor U2380 (N_2380,In_1245,In_1405);
nor U2381 (N_2381,In_1448,In_1541);
nor U2382 (N_2382,In_537,In_366);
nor U2383 (N_2383,In_816,In_1960);
and U2384 (N_2384,In_421,In_429);
nor U2385 (N_2385,In_1975,In_923);
and U2386 (N_2386,In_900,In_884);
xnor U2387 (N_2387,In_1651,In_1115);
or U2388 (N_2388,In_659,In_1193);
and U2389 (N_2389,In_792,In_943);
nor U2390 (N_2390,In_1836,In_892);
or U2391 (N_2391,In_1681,In_434);
nand U2392 (N_2392,In_1276,In_1596);
and U2393 (N_2393,In_1615,In_1207);
xor U2394 (N_2394,In_668,In_202);
xor U2395 (N_2395,In_261,In_917);
and U2396 (N_2396,In_1352,In_1402);
or U2397 (N_2397,In_661,In_1001);
nand U2398 (N_2398,In_417,In_1637);
or U2399 (N_2399,In_1948,In_592);
or U2400 (N_2400,In_1426,In_1666);
nor U2401 (N_2401,In_424,In_1139);
xor U2402 (N_2402,In_757,In_1575);
or U2403 (N_2403,In_1800,In_852);
or U2404 (N_2404,In_1080,In_920);
or U2405 (N_2405,In_1545,In_1496);
and U2406 (N_2406,In_1174,In_528);
nor U2407 (N_2407,In_731,In_969);
or U2408 (N_2408,In_1896,In_216);
or U2409 (N_2409,In_1942,In_738);
or U2410 (N_2410,In_511,In_764);
and U2411 (N_2411,In_144,In_394);
xnor U2412 (N_2412,In_856,In_1833);
xor U2413 (N_2413,In_1190,In_1140);
or U2414 (N_2414,In_387,In_1049);
nor U2415 (N_2415,In_1986,In_242);
or U2416 (N_2416,In_1878,In_209);
and U2417 (N_2417,In_1995,In_1079);
or U2418 (N_2418,In_1004,In_1995);
and U2419 (N_2419,In_34,In_1776);
xnor U2420 (N_2420,In_1256,In_127);
nor U2421 (N_2421,In_1881,In_1672);
nor U2422 (N_2422,In_410,In_1314);
or U2423 (N_2423,In_1970,In_477);
or U2424 (N_2424,In_1922,In_916);
or U2425 (N_2425,In_271,In_106);
or U2426 (N_2426,In_150,In_1068);
or U2427 (N_2427,In_292,In_1384);
nand U2428 (N_2428,In_1408,In_817);
and U2429 (N_2429,In_1583,In_1276);
or U2430 (N_2430,In_301,In_1474);
nor U2431 (N_2431,In_1354,In_1818);
nor U2432 (N_2432,In_986,In_1769);
or U2433 (N_2433,In_1530,In_620);
xnor U2434 (N_2434,In_17,In_1872);
and U2435 (N_2435,In_1937,In_1413);
nand U2436 (N_2436,In_710,In_1918);
and U2437 (N_2437,In_996,In_1298);
and U2438 (N_2438,In_712,In_1736);
nor U2439 (N_2439,In_159,In_1817);
nor U2440 (N_2440,In_1473,In_785);
and U2441 (N_2441,In_1606,In_1536);
nand U2442 (N_2442,In_784,In_1644);
xnor U2443 (N_2443,In_1875,In_1844);
or U2444 (N_2444,In_1739,In_1868);
nor U2445 (N_2445,In_1343,In_1145);
and U2446 (N_2446,In_208,In_1959);
nor U2447 (N_2447,In_793,In_735);
and U2448 (N_2448,In_346,In_1136);
xor U2449 (N_2449,In_116,In_663);
nand U2450 (N_2450,In_915,In_1994);
or U2451 (N_2451,In_1313,In_1271);
nor U2452 (N_2452,In_1985,In_115);
xnor U2453 (N_2453,In_208,In_1786);
nand U2454 (N_2454,In_1107,In_1168);
nor U2455 (N_2455,In_803,In_597);
and U2456 (N_2456,In_1284,In_1101);
nor U2457 (N_2457,In_421,In_339);
xnor U2458 (N_2458,In_1253,In_648);
nand U2459 (N_2459,In_1742,In_459);
and U2460 (N_2460,In_498,In_581);
nor U2461 (N_2461,In_156,In_785);
or U2462 (N_2462,In_227,In_137);
and U2463 (N_2463,In_1255,In_520);
or U2464 (N_2464,In_846,In_1355);
nand U2465 (N_2465,In_1398,In_1905);
and U2466 (N_2466,In_1536,In_815);
and U2467 (N_2467,In_1502,In_519);
nor U2468 (N_2468,In_1508,In_484);
or U2469 (N_2469,In_1985,In_1866);
nor U2470 (N_2470,In_22,In_856);
nor U2471 (N_2471,In_1720,In_763);
xnor U2472 (N_2472,In_1913,In_959);
nand U2473 (N_2473,In_685,In_673);
and U2474 (N_2474,In_1323,In_711);
nand U2475 (N_2475,In_1534,In_36);
or U2476 (N_2476,In_74,In_769);
nor U2477 (N_2477,In_1916,In_1518);
xor U2478 (N_2478,In_1592,In_1934);
nand U2479 (N_2479,In_271,In_890);
nor U2480 (N_2480,In_1305,In_893);
and U2481 (N_2481,In_488,In_1179);
or U2482 (N_2482,In_194,In_764);
nor U2483 (N_2483,In_314,In_1823);
nand U2484 (N_2484,In_1524,In_656);
nand U2485 (N_2485,In_899,In_919);
or U2486 (N_2486,In_632,In_942);
nor U2487 (N_2487,In_741,In_597);
and U2488 (N_2488,In_1250,In_656);
and U2489 (N_2489,In_1675,In_1128);
xor U2490 (N_2490,In_585,In_884);
xnor U2491 (N_2491,In_1191,In_116);
nor U2492 (N_2492,In_5,In_1309);
and U2493 (N_2493,In_1189,In_359);
nor U2494 (N_2494,In_1618,In_7);
xnor U2495 (N_2495,In_397,In_882);
and U2496 (N_2496,In_959,In_1716);
nand U2497 (N_2497,In_915,In_1305);
nand U2498 (N_2498,In_1720,In_117);
nor U2499 (N_2499,In_1269,In_501);
nand U2500 (N_2500,In_13,In_1131);
nand U2501 (N_2501,In_186,In_283);
or U2502 (N_2502,In_1966,In_1067);
nand U2503 (N_2503,In_963,In_1455);
nor U2504 (N_2504,In_1106,In_1422);
or U2505 (N_2505,In_124,In_1236);
and U2506 (N_2506,In_326,In_1367);
or U2507 (N_2507,In_1441,In_365);
xor U2508 (N_2508,In_1996,In_1366);
and U2509 (N_2509,In_1358,In_808);
or U2510 (N_2510,In_452,In_835);
nor U2511 (N_2511,In_1875,In_992);
xor U2512 (N_2512,In_1711,In_810);
nor U2513 (N_2513,In_1113,In_178);
or U2514 (N_2514,In_1069,In_1143);
nor U2515 (N_2515,In_1238,In_1929);
or U2516 (N_2516,In_1423,In_1993);
xnor U2517 (N_2517,In_1074,In_1274);
or U2518 (N_2518,In_1139,In_868);
nor U2519 (N_2519,In_1063,In_1728);
nand U2520 (N_2520,In_77,In_744);
nand U2521 (N_2521,In_1424,In_1514);
nor U2522 (N_2522,In_1212,In_1840);
xor U2523 (N_2523,In_1435,In_886);
nand U2524 (N_2524,In_1990,In_1673);
nor U2525 (N_2525,In_489,In_883);
and U2526 (N_2526,In_72,In_753);
xor U2527 (N_2527,In_348,In_807);
nand U2528 (N_2528,In_468,In_875);
xor U2529 (N_2529,In_97,In_711);
xor U2530 (N_2530,In_816,In_666);
nand U2531 (N_2531,In_970,In_1903);
or U2532 (N_2532,In_316,In_1534);
or U2533 (N_2533,In_750,In_1264);
xnor U2534 (N_2534,In_1562,In_1677);
nor U2535 (N_2535,In_358,In_628);
nor U2536 (N_2536,In_795,In_94);
nor U2537 (N_2537,In_1690,In_1413);
or U2538 (N_2538,In_582,In_9);
and U2539 (N_2539,In_806,In_1292);
and U2540 (N_2540,In_839,In_667);
or U2541 (N_2541,In_1378,In_1868);
xnor U2542 (N_2542,In_1131,In_1706);
xnor U2543 (N_2543,In_1241,In_1052);
nor U2544 (N_2544,In_1079,In_700);
nand U2545 (N_2545,In_823,In_321);
nor U2546 (N_2546,In_244,In_1787);
xnor U2547 (N_2547,In_1626,In_1864);
and U2548 (N_2548,In_1819,In_294);
or U2549 (N_2549,In_759,In_1510);
xor U2550 (N_2550,In_743,In_1136);
nand U2551 (N_2551,In_329,In_1577);
nand U2552 (N_2552,In_921,In_1627);
nor U2553 (N_2553,In_312,In_140);
xnor U2554 (N_2554,In_1229,In_1306);
and U2555 (N_2555,In_747,In_1205);
nor U2556 (N_2556,In_1927,In_1738);
and U2557 (N_2557,In_1725,In_1524);
and U2558 (N_2558,In_633,In_650);
nor U2559 (N_2559,In_1835,In_1756);
or U2560 (N_2560,In_1440,In_859);
nor U2561 (N_2561,In_1583,In_1220);
nor U2562 (N_2562,In_1776,In_176);
and U2563 (N_2563,In_1333,In_1190);
and U2564 (N_2564,In_754,In_967);
nand U2565 (N_2565,In_1339,In_1567);
and U2566 (N_2566,In_93,In_1311);
nor U2567 (N_2567,In_910,In_724);
and U2568 (N_2568,In_1619,In_1658);
nand U2569 (N_2569,In_1246,In_151);
xnor U2570 (N_2570,In_1994,In_186);
and U2571 (N_2571,In_1784,In_996);
xnor U2572 (N_2572,In_337,In_1894);
xor U2573 (N_2573,In_276,In_673);
nor U2574 (N_2574,In_384,In_79);
nand U2575 (N_2575,In_1766,In_1229);
nand U2576 (N_2576,In_1925,In_1464);
and U2577 (N_2577,In_181,In_1536);
and U2578 (N_2578,In_1375,In_744);
nor U2579 (N_2579,In_996,In_1455);
nand U2580 (N_2580,In_1956,In_517);
nor U2581 (N_2581,In_298,In_617);
nor U2582 (N_2582,In_197,In_169);
and U2583 (N_2583,In_1146,In_323);
nor U2584 (N_2584,In_696,In_411);
nor U2585 (N_2585,In_574,In_307);
and U2586 (N_2586,In_817,In_1503);
nand U2587 (N_2587,In_106,In_1212);
nand U2588 (N_2588,In_814,In_1768);
and U2589 (N_2589,In_581,In_941);
and U2590 (N_2590,In_1224,In_1826);
and U2591 (N_2591,In_1602,In_1865);
nand U2592 (N_2592,In_195,In_1484);
and U2593 (N_2593,In_839,In_994);
nand U2594 (N_2594,In_1629,In_594);
nand U2595 (N_2595,In_468,In_298);
and U2596 (N_2596,In_1009,In_1513);
nor U2597 (N_2597,In_1821,In_278);
nor U2598 (N_2598,In_1746,In_161);
xnor U2599 (N_2599,In_172,In_925);
nor U2600 (N_2600,In_776,In_1232);
nor U2601 (N_2601,In_904,In_1402);
and U2602 (N_2602,In_32,In_465);
xor U2603 (N_2603,In_1122,In_347);
xor U2604 (N_2604,In_805,In_646);
xnor U2605 (N_2605,In_634,In_589);
or U2606 (N_2606,In_764,In_457);
nand U2607 (N_2607,In_1560,In_730);
and U2608 (N_2608,In_1452,In_468);
nand U2609 (N_2609,In_1461,In_1551);
nor U2610 (N_2610,In_1887,In_394);
and U2611 (N_2611,In_290,In_159);
or U2612 (N_2612,In_1772,In_537);
or U2613 (N_2613,In_1815,In_701);
nor U2614 (N_2614,In_93,In_1966);
and U2615 (N_2615,In_618,In_244);
xor U2616 (N_2616,In_408,In_799);
xor U2617 (N_2617,In_1452,In_1020);
nor U2618 (N_2618,In_1698,In_613);
and U2619 (N_2619,In_404,In_1072);
nor U2620 (N_2620,In_1181,In_839);
and U2621 (N_2621,In_98,In_680);
or U2622 (N_2622,In_1953,In_750);
xnor U2623 (N_2623,In_1575,In_1012);
and U2624 (N_2624,In_869,In_1212);
xnor U2625 (N_2625,In_394,In_1303);
nand U2626 (N_2626,In_104,In_1625);
xnor U2627 (N_2627,In_1067,In_1398);
nor U2628 (N_2628,In_1451,In_1664);
nand U2629 (N_2629,In_1299,In_717);
xor U2630 (N_2630,In_1775,In_1916);
or U2631 (N_2631,In_1710,In_280);
nor U2632 (N_2632,In_611,In_1439);
nor U2633 (N_2633,In_640,In_695);
and U2634 (N_2634,In_1112,In_340);
nor U2635 (N_2635,In_1578,In_599);
and U2636 (N_2636,In_1310,In_739);
nor U2637 (N_2637,In_6,In_173);
nor U2638 (N_2638,In_132,In_1759);
nand U2639 (N_2639,In_754,In_1870);
and U2640 (N_2640,In_1902,In_862);
xnor U2641 (N_2641,In_1507,In_247);
or U2642 (N_2642,In_610,In_551);
nor U2643 (N_2643,In_1148,In_50);
or U2644 (N_2644,In_1426,In_1506);
and U2645 (N_2645,In_825,In_1238);
nand U2646 (N_2646,In_259,In_1011);
and U2647 (N_2647,In_229,In_348);
xnor U2648 (N_2648,In_1144,In_391);
nor U2649 (N_2649,In_1662,In_1585);
nand U2650 (N_2650,In_1609,In_188);
nand U2651 (N_2651,In_63,In_1299);
and U2652 (N_2652,In_1918,In_1503);
and U2653 (N_2653,In_372,In_415);
nand U2654 (N_2654,In_1286,In_1597);
nor U2655 (N_2655,In_879,In_1502);
nand U2656 (N_2656,In_1478,In_1592);
and U2657 (N_2657,In_1382,In_170);
nand U2658 (N_2658,In_1793,In_589);
and U2659 (N_2659,In_1568,In_871);
nor U2660 (N_2660,In_1359,In_372);
and U2661 (N_2661,In_1044,In_68);
nand U2662 (N_2662,In_1730,In_1045);
or U2663 (N_2663,In_339,In_177);
and U2664 (N_2664,In_379,In_1184);
nor U2665 (N_2665,In_406,In_934);
nand U2666 (N_2666,In_353,In_703);
xnor U2667 (N_2667,In_552,In_1984);
nand U2668 (N_2668,In_433,In_1213);
or U2669 (N_2669,In_688,In_199);
and U2670 (N_2670,In_352,In_1501);
nand U2671 (N_2671,In_566,In_1264);
nand U2672 (N_2672,In_1508,In_1567);
nor U2673 (N_2673,In_1786,In_256);
xor U2674 (N_2674,In_833,In_199);
xor U2675 (N_2675,In_266,In_1568);
and U2676 (N_2676,In_603,In_1003);
and U2677 (N_2677,In_1573,In_1989);
nand U2678 (N_2678,In_47,In_1279);
nor U2679 (N_2679,In_547,In_1047);
or U2680 (N_2680,In_1799,In_1156);
xor U2681 (N_2681,In_1726,In_1216);
nand U2682 (N_2682,In_1750,In_1602);
xnor U2683 (N_2683,In_518,In_1921);
nor U2684 (N_2684,In_130,In_1206);
and U2685 (N_2685,In_465,In_1);
nand U2686 (N_2686,In_1319,In_1396);
xnor U2687 (N_2687,In_275,In_1370);
or U2688 (N_2688,In_1189,In_176);
nor U2689 (N_2689,In_1397,In_120);
xor U2690 (N_2690,In_823,In_1426);
and U2691 (N_2691,In_505,In_184);
xor U2692 (N_2692,In_1072,In_387);
nor U2693 (N_2693,In_1506,In_119);
nor U2694 (N_2694,In_1288,In_502);
or U2695 (N_2695,In_1809,In_818);
or U2696 (N_2696,In_1447,In_385);
nor U2697 (N_2697,In_1149,In_1237);
nand U2698 (N_2698,In_1732,In_366);
nor U2699 (N_2699,In_392,In_572);
or U2700 (N_2700,In_598,In_1987);
and U2701 (N_2701,In_474,In_632);
xor U2702 (N_2702,In_1197,In_877);
or U2703 (N_2703,In_723,In_1134);
nor U2704 (N_2704,In_254,In_117);
nor U2705 (N_2705,In_906,In_1178);
and U2706 (N_2706,In_1937,In_1690);
nor U2707 (N_2707,In_642,In_786);
nor U2708 (N_2708,In_1560,In_604);
and U2709 (N_2709,In_1593,In_263);
nor U2710 (N_2710,In_535,In_1765);
or U2711 (N_2711,In_1705,In_672);
and U2712 (N_2712,In_996,In_922);
or U2713 (N_2713,In_76,In_457);
and U2714 (N_2714,In_1714,In_598);
nand U2715 (N_2715,In_400,In_942);
nand U2716 (N_2716,In_1536,In_732);
nor U2717 (N_2717,In_280,In_1372);
nand U2718 (N_2718,In_648,In_13);
xnor U2719 (N_2719,In_86,In_1064);
nor U2720 (N_2720,In_1585,In_1188);
or U2721 (N_2721,In_1420,In_500);
xnor U2722 (N_2722,In_1146,In_373);
xor U2723 (N_2723,In_157,In_1708);
xor U2724 (N_2724,In_827,In_1268);
nand U2725 (N_2725,In_452,In_1369);
nor U2726 (N_2726,In_410,In_738);
or U2727 (N_2727,In_1483,In_464);
nor U2728 (N_2728,In_1662,In_1094);
xnor U2729 (N_2729,In_1841,In_152);
nor U2730 (N_2730,In_1024,In_1122);
nor U2731 (N_2731,In_1809,In_1547);
nand U2732 (N_2732,In_503,In_1720);
xor U2733 (N_2733,In_418,In_948);
nand U2734 (N_2734,In_514,In_1556);
nor U2735 (N_2735,In_558,In_1769);
nand U2736 (N_2736,In_1795,In_23);
or U2737 (N_2737,In_1496,In_550);
nand U2738 (N_2738,In_1445,In_1098);
xnor U2739 (N_2739,In_117,In_384);
nand U2740 (N_2740,In_485,In_1696);
nor U2741 (N_2741,In_11,In_719);
nand U2742 (N_2742,In_287,In_1983);
nand U2743 (N_2743,In_1891,In_544);
xnor U2744 (N_2744,In_841,In_317);
nand U2745 (N_2745,In_705,In_1294);
and U2746 (N_2746,In_1272,In_1154);
and U2747 (N_2747,In_1531,In_539);
nand U2748 (N_2748,In_1032,In_1399);
and U2749 (N_2749,In_168,In_1470);
or U2750 (N_2750,In_1130,In_694);
nor U2751 (N_2751,In_698,In_1466);
nand U2752 (N_2752,In_1451,In_1441);
xnor U2753 (N_2753,In_1671,In_1640);
or U2754 (N_2754,In_1273,In_384);
nand U2755 (N_2755,In_1967,In_1633);
xnor U2756 (N_2756,In_427,In_468);
xor U2757 (N_2757,In_1653,In_1270);
nand U2758 (N_2758,In_1588,In_1636);
and U2759 (N_2759,In_90,In_224);
nor U2760 (N_2760,In_1379,In_1229);
nand U2761 (N_2761,In_1908,In_181);
or U2762 (N_2762,In_316,In_185);
xor U2763 (N_2763,In_391,In_1086);
nand U2764 (N_2764,In_1420,In_883);
nand U2765 (N_2765,In_1702,In_17);
nand U2766 (N_2766,In_806,In_1747);
nor U2767 (N_2767,In_1255,In_1466);
xnor U2768 (N_2768,In_1543,In_1036);
nand U2769 (N_2769,In_63,In_154);
nand U2770 (N_2770,In_136,In_1423);
nand U2771 (N_2771,In_421,In_573);
or U2772 (N_2772,In_862,In_276);
xor U2773 (N_2773,In_1121,In_1885);
xor U2774 (N_2774,In_1966,In_718);
nor U2775 (N_2775,In_1172,In_1215);
and U2776 (N_2776,In_1116,In_1338);
xnor U2777 (N_2777,In_23,In_859);
nand U2778 (N_2778,In_1599,In_171);
and U2779 (N_2779,In_154,In_721);
xor U2780 (N_2780,In_496,In_1712);
and U2781 (N_2781,In_701,In_1805);
xor U2782 (N_2782,In_541,In_41);
nand U2783 (N_2783,In_1838,In_1388);
nand U2784 (N_2784,In_1917,In_1388);
nor U2785 (N_2785,In_1170,In_920);
or U2786 (N_2786,In_1368,In_1145);
xnor U2787 (N_2787,In_16,In_1913);
or U2788 (N_2788,In_1341,In_753);
and U2789 (N_2789,In_284,In_176);
and U2790 (N_2790,In_623,In_818);
nor U2791 (N_2791,In_1253,In_233);
xor U2792 (N_2792,In_1624,In_1061);
or U2793 (N_2793,In_104,In_289);
xnor U2794 (N_2794,In_14,In_1047);
nand U2795 (N_2795,In_1361,In_310);
or U2796 (N_2796,In_571,In_1081);
nor U2797 (N_2797,In_747,In_1567);
nand U2798 (N_2798,In_514,In_525);
nor U2799 (N_2799,In_560,In_1093);
nor U2800 (N_2800,In_779,In_209);
xor U2801 (N_2801,In_1208,In_328);
or U2802 (N_2802,In_186,In_892);
nand U2803 (N_2803,In_254,In_1800);
xor U2804 (N_2804,In_1126,In_1452);
nand U2805 (N_2805,In_1829,In_1589);
or U2806 (N_2806,In_790,In_788);
and U2807 (N_2807,In_1987,In_1655);
nor U2808 (N_2808,In_1378,In_130);
nor U2809 (N_2809,In_1001,In_529);
nor U2810 (N_2810,In_1867,In_730);
xnor U2811 (N_2811,In_1828,In_716);
and U2812 (N_2812,In_186,In_811);
nand U2813 (N_2813,In_1474,In_1628);
and U2814 (N_2814,In_372,In_1947);
and U2815 (N_2815,In_287,In_1515);
nor U2816 (N_2816,In_936,In_680);
and U2817 (N_2817,In_408,In_183);
nand U2818 (N_2818,In_761,In_1125);
xnor U2819 (N_2819,In_1320,In_1109);
and U2820 (N_2820,In_1339,In_1778);
nand U2821 (N_2821,In_669,In_1800);
xnor U2822 (N_2822,In_311,In_1935);
and U2823 (N_2823,In_428,In_1748);
and U2824 (N_2824,In_737,In_1575);
nor U2825 (N_2825,In_248,In_757);
nor U2826 (N_2826,In_1910,In_1187);
or U2827 (N_2827,In_1901,In_858);
nor U2828 (N_2828,In_467,In_1962);
nand U2829 (N_2829,In_683,In_686);
xnor U2830 (N_2830,In_507,In_977);
xnor U2831 (N_2831,In_343,In_1706);
xor U2832 (N_2832,In_1173,In_1590);
nor U2833 (N_2833,In_721,In_1311);
or U2834 (N_2834,In_45,In_1187);
nand U2835 (N_2835,In_1496,In_360);
nand U2836 (N_2836,In_341,In_245);
nor U2837 (N_2837,In_1916,In_1864);
nor U2838 (N_2838,In_552,In_451);
nor U2839 (N_2839,In_946,In_1144);
or U2840 (N_2840,In_352,In_288);
or U2841 (N_2841,In_959,In_1672);
and U2842 (N_2842,In_397,In_1551);
and U2843 (N_2843,In_1017,In_1585);
or U2844 (N_2844,In_213,In_1414);
and U2845 (N_2845,In_161,In_1661);
or U2846 (N_2846,In_151,In_1395);
xor U2847 (N_2847,In_1017,In_296);
nor U2848 (N_2848,In_1007,In_1491);
nand U2849 (N_2849,In_1877,In_1276);
nor U2850 (N_2850,In_1293,In_498);
or U2851 (N_2851,In_1062,In_444);
and U2852 (N_2852,In_1148,In_1403);
and U2853 (N_2853,In_1134,In_524);
nand U2854 (N_2854,In_1686,In_1345);
or U2855 (N_2855,In_1718,In_1996);
and U2856 (N_2856,In_210,In_1704);
and U2857 (N_2857,In_1267,In_53);
nor U2858 (N_2858,In_586,In_101);
nand U2859 (N_2859,In_900,In_1166);
and U2860 (N_2860,In_1203,In_1760);
nor U2861 (N_2861,In_1966,In_350);
and U2862 (N_2862,In_108,In_926);
xor U2863 (N_2863,In_1104,In_1166);
xnor U2864 (N_2864,In_193,In_638);
xnor U2865 (N_2865,In_244,In_1968);
nand U2866 (N_2866,In_1525,In_1671);
xor U2867 (N_2867,In_1233,In_1007);
or U2868 (N_2868,In_179,In_1473);
nand U2869 (N_2869,In_1817,In_134);
xnor U2870 (N_2870,In_33,In_1205);
nor U2871 (N_2871,In_1022,In_1718);
and U2872 (N_2872,In_1641,In_413);
xnor U2873 (N_2873,In_1183,In_1103);
nand U2874 (N_2874,In_925,In_438);
nand U2875 (N_2875,In_323,In_269);
or U2876 (N_2876,In_462,In_597);
xor U2877 (N_2877,In_1283,In_1095);
nor U2878 (N_2878,In_1260,In_1478);
and U2879 (N_2879,In_1938,In_1572);
nand U2880 (N_2880,In_1742,In_1014);
or U2881 (N_2881,In_1033,In_1062);
or U2882 (N_2882,In_773,In_1349);
xnor U2883 (N_2883,In_1653,In_440);
nor U2884 (N_2884,In_1434,In_1047);
nor U2885 (N_2885,In_711,In_620);
xnor U2886 (N_2886,In_829,In_481);
and U2887 (N_2887,In_658,In_752);
nand U2888 (N_2888,In_1265,In_583);
xor U2889 (N_2889,In_1973,In_258);
and U2890 (N_2890,In_560,In_751);
nor U2891 (N_2891,In_474,In_1045);
nand U2892 (N_2892,In_1034,In_1869);
xnor U2893 (N_2893,In_142,In_861);
nor U2894 (N_2894,In_1893,In_692);
and U2895 (N_2895,In_1282,In_1867);
nor U2896 (N_2896,In_1503,In_1618);
xor U2897 (N_2897,In_1983,In_63);
and U2898 (N_2898,In_517,In_148);
xnor U2899 (N_2899,In_70,In_286);
xor U2900 (N_2900,In_1824,In_463);
nor U2901 (N_2901,In_1157,In_1169);
nor U2902 (N_2902,In_917,In_1037);
xnor U2903 (N_2903,In_559,In_1705);
and U2904 (N_2904,In_1461,In_561);
nand U2905 (N_2905,In_889,In_1380);
nand U2906 (N_2906,In_914,In_1573);
nor U2907 (N_2907,In_1520,In_1686);
xnor U2908 (N_2908,In_1567,In_628);
nor U2909 (N_2909,In_1978,In_449);
or U2910 (N_2910,In_1283,In_1934);
nor U2911 (N_2911,In_1974,In_1175);
or U2912 (N_2912,In_748,In_810);
xnor U2913 (N_2913,In_497,In_535);
or U2914 (N_2914,In_1398,In_573);
nor U2915 (N_2915,In_1657,In_1963);
xnor U2916 (N_2916,In_1284,In_1248);
xor U2917 (N_2917,In_605,In_416);
nor U2918 (N_2918,In_706,In_1411);
nor U2919 (N_2919,In_1714,In_984);
and U2920 (N_2920,In_1474,In_527);
xor U2921 (N_2921,In_170,In_1931);
and U2922 (N_2922,In_69,In_538);
or U2923 (N_2923,In_1734,In_258);
or U2924 (N_2924,In_1067,In_513);
and U2925 (N_2925,In_1948,In_960);
xnor U2926 (N_2926,In_998,In_477);
and U2927 (N_2927,In_1896,In_447);
nor U2928 (N_2928,In_1148,In_843);
and U2929 (N_2929,In_161,In_1760);
nand U2930 (N_2930,In_694,In_1376);
nor U2931 (N_2931,In_116,In_1199);
xor U2932 (N_2932,In_625,In_1024);
or U2933 (N_2933,In_1820,In_1406);
xor U2934 (N_2934,In_571,In_1199);
and U2935 (N_2935,In_623,In_1638);
nor U2936 (N_2936,In_1177,In_983);
nor U2937 (N_2937,In_1966,In_1486);
nand U2938 (N_2938,In_503,In_255);
xnor U2939 (N_2939,In_41,In_431);
or U2940 (N_2940,In_743,In_1491);
or U2941 (N_2941,In_1782,In_1324);
nor U2942 (N_2942,In_1295,In_1233);
or U2943 (N_2943,In_535,In_1906);
and U2944 (N_2944,In_1516,In_1909);
xnor U2945 (N_2945,In_1823,In_1908);
nor U2946 (N_2946,In_462,In_179);
nand U2947 (N_2947,In_1865,In_1272);
and U2948 (N_2948,In_1240,In_92);
nor U2949 (N_2949,In_396,In_103);
and U2950 (N_2950,In_1709,In_184);
nor U2951 (N_2951,In_65,In_1445);
and U2952 (N_2952,In_482,In_521);
nor U2953 (N_2953,In_416,In_946);
and U2954 (N_2954,In_654,In_959);
xnor U2955 (N_2955,In_1708,In_937);
nor U2956 (N_2956,In_353,In_364);
nor U2957 (N_2957,In_1437,In_709);
nand U2958 (N_2958,In_237,In_1840);
nor U2959 (N_2959,In_1051,In_1812);
or U2960 (N_2960,In_758,In_210);
nor U2961 (N_2961,In_384,In_1270);
and U2962 (N_2962,In_1910,In_596);
nand U2963 (N_2963,In_1568,In_256);
or U2964 (N_2964,In_636,In_1381);
nor U2965 (N_2965,In_484,In_54);
xnor U2966 (N_2966,In_563,In_697);
xor U2967 (N_2967,In_1877,In_1288);
or U2968 (N_2968,In_1438,In_238);
nor U2969 (N_2969,In_352,In_1682);
and U2970 (N_2970,In_959,In_927);
nor U2971 (N_2971,In_538,In_1567);
nand U2972 (N_2972,In_791,In_1323);
xor U2973 (N_2973,In_797,In_1678);
nor U2974 (N_2974,In_944,In_134);
and U2975 (N_2975,In_934,In_984);
xor U2976 (N_2976,In_1931,In_909);
and U2977 (N_2977,In_450,In_939);
or U2978 (N_2978,In_1177,In_1695);
or U2979 (N_2979,In_594,In_294);
nor U2980 (N_2980,In_1617,In_1006);
or U2981 (N_2981,In_1883,In_184);
or U2982 (N_2982,In_1156,In_641);
xnor U2983 (N_2983,In_1217,In_1458);
nand U2984 (N_2984,In_1916,In_714);
xnor U2985 (N_2985,In_636,In_1703);
nand U2986 (N_2986,In_802,In_888);
and U2987 (N_2987,In_966,In_1400);
nand U2988 (N_2988,In_302,In_278);
and U2989 (N_2989,In_837,In_1135);
or U2990 (N_2990,In_201,In_1529);
or U2991 (N_2991,In_345,In_1970);
and U2992 (N_2992,In_1035,In_689);
nand U2993 (N_2993,In_1552,In_15);
or U2994 (N_2994,In_190,In_776);
xnor U2995 (N_2995,In_1981,In_442);
nand U2996 (N_2996,In_1461,In_635);
or U2997 (N_2997,In_1651,In_1170);
nand U2998 (N_2998,In_702,In_55);
nor U2999 (N_2999,In_1901,In_365);
xor U3000 (N_3000,In_1101,In_1332);
or U3001 (N_3001,In_506,In_337);
and U3002 (N_3002,In_1486,In_113);
or U3003 (N_3003,In_155,In_1682);
xnor U3004 (N_3004,In_139,In_1575);
xor U3005 (N_3005,In_1868,In_617);
nand U3006 (N_3006,In_1773,In_192);
nand U3007 (N_3007,In_1696,In_743);
or U3008 (N_3008,In_1890,In_1513);
or U3009 (N_3009,In_1324,In_557);
and U3010 (N_3010,In_854,In_541);
xor U3011 (N_3011,In_190,In_1156);
nand U3012 (N_3012,In_1350,In_1196);
xor U3013 (N_3013,In_1085,In_163);
xnor U3014 (N_3014,In_87,In_499);
or U3015 (N_3015,In_1253,In_1665);
xnor U3016 (N_3016,In_1664,In_492);
xnor U3017 (N_3017,In_1363,In_1050);
and U3018 (N_3018,In_1543,In_152);
and U3019 (N_3019,In_1364,In_1219);
nand U3020 (N_3020,In_1578,In_1984);
and U3021 (N_3021,In_1927,In_1720);
nor U3022 (N_3022,In_881,In_1016);
xnor U3023 (N_3023,In_852,In_1786);
or U3024 (N_3024,In_738,In_1241);
xor U3025 (N_3025,In_543,In_611);
or U3026 (N_3026,In_1339,In_886);
or U3027 (N_3027,In_733,In_1981);
xor U3028 (N_3028,In_1417,In_939);
xnor U3029 (N_3029,In_1097,In_447);
nand U3030 (N_3030,In_621,In_178);
xnor U3031 (N_3031,In_1690,In_1316);
or U3032 (N_3032,In_1707,In_42);
nand U3033 (N_3033,In_1595,In_776);
nor U3034 (N_3034,In_25,In_1568);
or U3035 (N_3035,In_1366,In_809);
nand U3036 (N_3036,In_1811,In_1925);
or U3037 (N_3037,In_40,In_1382);
nand U3038 (N_3038,In_1521,In_1124);
and U3039 (N_3039,In_1926,In_1633);
xnor U3040 (N_3040,In_1951,In_559);
and U3041 (N_3041,In_609,In_992);
nand U3042 (N_3042,In_1482,In_558);
and U3043 (N_3043,In_337,In_245);
and U3044 (N_3044,In_453,In_555);
nand U3045 (N_3045,In_1406,In_1732);
or U3046 (N_3046,In_1920,In_1930);
nor U3047 (N_3047,In_1262,In_1450);
or U3048 (N_3048,In_349,In_657);
nand U3049 (N_3049,In_646,In_684);
and U3050 (N_3050,In_1131,In_1579);
and U3051 (N_3051,In_1228,In_1896);
nor U3052 (N_3052,In_1916,In_660);
nor U3053 (N_3053,In_191,In_1212);
nor U3054 (N_3054,In_1776,In_783);
xor U3055 (N_3055,In_999,In_799);
nand U3056 (N_3056,In_822,In_1911);
nand U3057 (N_3057,In_1581,In_416);
xor U3058 (N_3058,In_624,In_887);
nand U3059 (N_3059,In_1107,In_1149);
nand U3060 (N_3060,In_1297,In_929);
nor U3061 (N_3061,In_472,In_1074);
or U3062 (N_3062,In_1954,In_1839);
xnor U3063 (N_3063,In_927,In_723);
xor U3064 (N_3064,In_1502,In_1280);
nor U3065 (N_3065,In_244,In_651);
or U3066 (N_3066,In_524,In_164);
and U3067 (N_3067,In_396,In_862);
nand U3068 (N_3068,In_556,In_395);
nand U3069 (N_3069,In_1003,In_1873);
and U3070 (N_3070,In_641,In_703);
xnor U3071 (N_3071,In_1745,In_1272);
nor U3072 (N_3072,In_470,In_970);
nand U3073 (N_3073,In_903,In_1440);
or U3074 (N_3074,In_475,In_914);
nand U3075 (N_3075,In_1817,In_1767);
xnor U3076 (N_3076,In_64,In_285);
and U3077 (N_3077,In_943,In_168);
nor U3078 (N_3078,In_1786,In_1692);
or U3079 (N_3079,In_507,In_1135);
nor U3080 (N_3080,In_570,In_1288);
xnor U3081 (N_3081,In_1336,In_946);
xnor U3082 (N_3082,In_216,In_1346);
nand U3083 (N_3083,In_971,In_269);
nand U3084 (N_3084,In_948,In_643);
nor U3085 (N_3085,In_1463,In_1825);
nor U3086 (N_3086,In_1240,In_924);
nand U3087 (N_3087,In_1229,In_1407);
xor U3088 (N_3088,In_1422,In_1300);
and U3089 (N_3089,In_579,In_1598);
or U3090 (N_3090,In_392,In_602);
xor U3091 (N_3091,In_1802,In_1907);
and U3092 (N_3092,In_438,In_1731);
nor U3093 (N_3093,In_937,In_1730);
xnor U3094 (N_3094,In_480,In_364);
nor U3095 (N_3095,In_1249,In_186);
nor U3096 (N_3096,In_1266,In_1595);
and U3097 (N_3097,In_1725,In_889);
xor U3098 (N_3098,In_416,In_1557);
or U3099 (N_3099,In_1188,In_445);
xor U3100 (N_3100,In_1869,In_1434);
or U3101 (N_3101,In_712,In_1642);
nor U3102 (N_3102,In_1741,In_14);
and U3103 (N_3103,In_1735,In_1053);
nand U3104 (N_3104,In_972,In_791);
nor U3105 (N_3105,In_1303,In_1364);
xnor U3106 (N_3106,In_519,In_657);
nand U3107 (N_3107,In_213,In_915);
nand U3108 (N_3108,In_769,In_721);
nand U3109 (N_3109,In_952,In_1977);
or U3110 (N_3110,In_560,In_261);
or U3111 (N_3111,In_364,In_1478);
nor U3112 (N_3112,In_242,In_127);
and U3113 (N_3113,In_117,In_1295);
nand U3114 (N_3114,In_797,In_1499);
and U3115 (N_3115,In_1272,In_1549);
nand U3116 (N_3116,In_294,In_954);
or U3117 (N_3117,In_1466,In_889);
or U3118 (N_3118,In_1892,In_699);
and U3119 (N_3119,In_253,In_1782);
or U3120 (N_3120,In_1161,In_868);
nand U3121 (N_3121,In_314,In_128);
xor U3122 (N_3122,In_1714,In_140);
and U3123 (N_3123,In_1434,In_1296);
and U3124 (N_3124,In_823,In_364);
nand U3125 (N_3125,In_1086,In_332);
nor U3126 (N_3126,In_1970,In_1177);
and U3127 (N_3127,In_1199,In_584);
xnor U3128 (N_3128,In_983,In_1460);
nand U3129 (N_3129,In_1462,In_1035);
or U3130 (N_3130,In_509,In_1429);
or U3131 (N_3131,In_997,In_248);
nand U3132 (N_3132,In_1161,In_407);
xnor U3133 (N_3133,In_986,In_345);
nor U3134 (N_3134,In_1032,In_1924);
xnor U3135 (N_3135,In_1132,In_323);
nor U3136 (N_3136,In_1378,In_1991);
nand U3137 (N_3137,In_100,In_792);
and U3138 (N_3138,In_892,In_469);
and U3139 (N_3139,In_1781,In_1272);
xnor U3140 (N_3140,In_1605,In_468);
nand U3141 (N_3141,In_538,In_1771);
xor U3142 (N_3142,In_305,In_990);
nor U3143 (N_3143,In_841,In_1685);
nor U3144 (N_3144,In_1275,In_1863);
xnor U3145 (N_3145,In_1535,In_955);
nor U3146 (N_3146,In_1308,In_494);
nand U3147 (N_3147,In_521,In_1865);
nor U3148 (N_3148,In_1692,In_381);
nand U3149 (N_3149,In_379,In_1914);
nand U3150 (N_3150,In_263,In_1359);
or U3151 (N_3151,In_1347,In_965);
nand U3152 (N_3152,In_1992,In_29);
and U3153 (N_3153,In_1856,In_106);
nor U3154 (N_3154,In_613,In_1487);
nor U3155 (N_3155,In_1441,In_672);
nand U3156 (N_3156,In_98,In_1364);
xor U3157 (N_3157,In_188,In_1897);
xor U3158 (N_3158,In_1331,In_1753);
nand U3159 (N_3159,In_581,In_146);
or U3160 (N_3160,In_922,In_422);
nand U3161 (N_3161,In_660,In_1507);
or U3162 (N_3162,In_7,In_569);
nor U3163 (N_3163,In_321,In_1080);
xnor U3164 (N_3164,In_1018,In_151);
or U3165 (N_3165,In_676,In_65);
xnor U3166 (N_3166,In_1119,In_872);
and U3167 (N_3167,In_1332,In_438);
nand U3168 (N_3168,In_86,In_1271);
and U3169 (N_3169,In_222,In_898);
nand U3170 (N_3170,In_809,In_24);
nand U3171 (N_3171,In_1232,In_674);
and U3172 (N_3172,In_607,In_371);
xnor U3173 (N_3173,In_1856,In_1990);
and U3174 (N_3174,In_1119,In_1984);
or U3175 (N_3175,In_571,In_116);
xnor U3176 (N_3176,In_793,In_1888);
nand U3177 (N_3177,In_1604,In_1038);
or U3178 (N_3178,In_596,In_1854);
nand U3179 (N_3179,In_629,In_810);
or U3180 (N_3180,In_1618,In_1690);
xnor U3181 (N_3181,In_980,In_1254);
nor U3182 (N_3182,In_1167,In_1126);
nand U3183 (N_3183,In_418,In_681);
or U3184 (N_3184,In_1274,In_84);
xnor U3185 (N_3185,In_1929,In_71);
xnor U3186 (N_3186,In_481,In_708);
nand U3187 (N_3187,In_306,In_1484);
xnor U3188 (N_3188,In_361,In_1364);
xor U3189 (N_3189,In_213,In_1193);
or U3190 (N_3190,In_1150,In_1652);
nand U3191 (N_3191,In_639,In_1073);
or U3192 (N_3192,In_601,In_790);
and U3193 (N_3193,In_1100,In_1545);
or U3194 (N_3194,In_1763,In_262);
xnor U3195 (N_3195,In_1631,In_314);
nor U3196 (N_3196,In_38,In_847);
nand U3197 (N_3197,In_330,In_1663);
and U3198 (N_3198,In_1188,In_1227);
xor U3199 (N_3199,In_639,In_588);
and U3200 (N_3200,In_681,In_1680);
nor U3201 (N_3201,In_7,In_677);
or U3202 (N_3202,In_1834,In_103);
nand U3203 (N_3203,In_32,In_59);
nand U3204 (N_3204,In_525,In_1688);
nor U3205 (N_3205,In_452,In_666);
nand U3206 (N_3206,In_1063,In_1272);
nor U3207 (N_3207,In_21,In_1878);
or U3208 (N_3208,In_284,In_125);
or U3209 (N_3209,In_1180,In_1848);
nand U3210 (N_3210,In_386,In_105);
or U3211 (N_3211,In_890,In_564);
and U3212 (N_3212,In_755,In_273);
nand U3213 (N_3213,In_1159,In_802);
xnor U3214 (N_3214,In_397,In_1651);
and U3215 (N_3215,In_1395,In_213);
and U3216 (N_3216,In_440,In_1675);
nand U3217 (N_3217,In_1571,In_927);
nand U3218 (N_3218,In_1123,In_345);
or U3219 (N_3219,In_434,In_1472);
nor U3220 (N_3220,In_305,In_1837);
nor U3221 (N_3221,In_1952,In_251);
nand U3222 (N_3222,In_1777,In_589);
nand U3223 (N_3223,In_130,In_593);
nand U3224 (N_3224,In_348,In_1504);
nor U3225 (N_3225,In_505,In_125);
xnor U3226 (N_3226,In_1976,In_703);
nor U3227 (N_3227,In_475,In_178);
and U3228 (N_3228,In_1398,In_1553);
or U3229 (N_3229,In_1780,In_1185);
nor U3230 (N_3230,In_1495,In_87);
or U3231 (N_3231,In_134,In_627);
nor U3232 (N_3232,In_1714,In_1376);
and U3233 (N_3233,In_1989,In_1125);
nor U3234 (N_3234,In_751,In_908);
or U3235 (N_3235,In_552,In_96);
or U3236 (N_3236,In_379,In_319);
nand U3237 (N_3237,In_1345,In_1793);
nand U3238 (N_3238,In_1891,In_352);
and U3239 (N_3239,In_474,In_1379);
nand U3240 (N_3240,In_1140,In_1452);
or U3241 (N_3241,In_953,In_236);
or U3242 (N_3242,In_1846,In_646);
nor U3243 (N_3243,In_926,In_1413);
nand U3244 (N_3244,In_1509,In_534);
nand U3245 (N_3245,In_1704,In_553);
and U3246 (N_3246,In_69,In_1211);
and U3247 (N_3247,In_817,In_352);
or U3248 (N_3248,In_203,In_40);
nor U3249 (N_3249,In_476,In_588);
or U3250 (N_3250,In_659,In_1840);
xor U3251 (N_3251,In_959,In_1630);
nor U3252 (N_3252,In_903,In_1121);
and U3253 (N_3253,In_112,In_633);
nand U3254 (N_3254,In_909,In_673);
nand U3255 (N_3255,In_1148,In_475);
nand U3256 (N_3256,In_1149,In_898);
nand U3257 (N_3257,In_1798,In_1198);
nand U3258 (N_3258,In_1732,In_1669);
or U3259 (N_3259,In_157,In_242);
nand U3260 (N_3260,In_237,In_534);
and U3261 (N_3261,In_1362,In_590);
nor U3262 (N_3262,In_251,In_1541);
xor U3263 (N_3263,In_1423,In_1404);
and U3264 (N_3264,In_92,In_538);
nand U3265 (N_3265,In_497,In_1630);
nor U3266 (N_3266,In_1972,In_1889);
and U3267 (N_3267,In_549,In_121);
nor U3268 (N_3268,In_1243,In_1331);
or U3269 (N_3269,In_951,In_1037);
nor U3270 (N_3270,In_572,In_1311);
nand U3271 (N_3271,In_549,In_64);
and U3272 (N_3272,In_368,In_1301);
nor U3273 (N_3273,In_184,In_543);
nor U3274 (N_3274,In_817,In_162);
nor U3275 (N_3275,In_169,In_1749);
nand U3276 (N_3276,In_822,In_1102);
or U3277 (N_3277,In_1314,In_721);
or U3278 (N_3278,In_1274,In_894);
nor U3279 (N_3279,In_1160,In_413);
and U3280 (N_3280,In_748,In_1639);
xnor U3281 (N_3281,In_230,In_356);
xor U3282 (N_3282,In_462,In_1272);
nor U3283 (N_3283,In_1822,In_1193);
nor U3284 (N_3284,In_1934,In_1742);
xor U3285 (N_3285,In_103,In_1158);
xor U3286 (N_3286,In_1955,In_61);
nand U3287 (N_3287,In_959,In_392);
nor U3288 (N_3288,In_344,In_786);
and U3289 (N_3289,In_461,In_790);
or U3290 (N_3290,In_1763,In_38);
xor U3291 (N_3291,In_1632,In_1303);
or U3292 (N_3292,In_1965,In_442);
nand U3293 (N_3293,In_234,In_1500);
and U3294 (N_3294,In_1681,In_97);
or U3295 (N_3295,In_1285,In_1576);
xor U3296 (N_3296,In_1192,In_1321);
or U3297 (N_3297,In_884,In_1176);
xor U3298 (N_3298,In_1801,In_330);
xor U3299 (N_3299,In_1907,In_177);
xor U3300 (N_3300,In_1220,In_152);
and U3301 (N_3301,In_848,In_350);
or U3302 (N_3302,In_42,In_824);
nand U3303 (N_3303,In_364,In_1548);
nand U3304 (N_3304,In_1150,In_901);
and U3305 (N_3305,In_1695,In_1411);
xnor U3306 (N_3306,In_798,In_1587);
or U3307 (N_3307,In_834,In_786);
xor U3308 (N_3308,In_262,In_512);
or U3309 (N_3309,In_403,In_1565);
nor U3310 (N_3310,In_1516,In_723);
or U3311 (N_3311,In_29,In_1584);
nor U3312 (N_3312,In_33,In_479);
or U3313 (N_3313,In_1943,In_1449);
and U3314 (N_3314,In_1807,In_8);
nand U3315 (N_3315,In_1486,In_1208);
nand U3316 (N_3316,In_771,In_1683);
and U3317 (N_3317,In_1069,In_1608);
nand U3318 (N_3318,In_717,In_648);
or U3319 (N_3319,In_956,In_1149);
nor U3320 (N_3320,In_526,In_1689);
and U3321 (N_3321,In_1920,In_1686);
and U3322 (N_3322,In_1711,In_516);
xnor U3323 (N_3323,In_1323,In_1879);
xor U3324 (N_3324,In_942,In_848);
xor U3325 (N_3325,In_1923,In_1900);
nor U3326 (N_3326,In_1793,In_1708);
xor U3327 (N_3327,In_1752,In_1325);
nor U3328 (N_3328,In_1962,In_33);
nor U3329 (N_3329,In_213,In_1129);
xor U3330 (N_3330,In_728,In_647);
nand U3331 (N_3331,In_1117,In_1636);
nor U3332 (N_3332,In_26,In_1463);
nand U3333 (N_3333,In_302,In_831);
xor U3334 (N_3334,In_1586,In_151);
xnor U3335 (N_3335,In_1378,In_1879);
nand U3336 (N_3336,In_1885,In_230);
or U3337 (N_3337,In_1238,In_1887);
nand U3338 (N_3338,In_1521,In_1990);
nor U3339 (N_3339,In_1269,In_249);
nand U3340 (N_3340,In_1079,In_722);
xor U3341 (N_3341,In_1054,In_789);
or U3342 (N_3342,In_1840,In_497);
and U3343 (N_3343,In_283,In_916);
nand U3344 (N_3344,In_726,In_554);
xnor U3345 (N_3345,In_221,In_1996);
xor U3346 (N_3346,In_945,In_359);
and U3347 (N_3347,In_748,In_1090);
and U3348 (N_3348,In_249,In_935);
and U3349 (N_3349,In_803,In_54);
or U3350 (N_3350,In_1004,In_1247);
or U3351 (N_3351,In_1210,In_1556);
or U3352 (N_3352,In_322,In_652);
xnor U3353 (N_3353,In_1346,In_538);
and U3354 (N_3354,In_972,In_918);
or U3355 (N_3355,In_77,In_1083);
and U3356 (N_3356,In_1441,In_819);
nand U3357 (N_3357,In_936,In_51);
and U3358 (N_3358,In_1682,In_1019);
nand U3359 (N_3359,In_744,In_1661);
xnor U3360 (N_3360,In_441,In_1766);
nand U3361 (N_3361,In_1024,In_368);
xnor U3362 (N_3362,In_1174,In_1392);
nor U3363 (N_3363,In_155,In_560);
nor U3364 (N_3364,In_1391,In_1936);
nand U3365 (N_3365,In_1424,In_1323);
xnor U3366 (N_3366,In_433,In_1617);
and U3367 (N_3367,In_1905,In_1108);
and U3368 (N_3368,In_1435,In_1421);
and U3369 (N_3369,In_1297,In_498);
and U3370 (N_3370,In_1810,In_215);
xnor U3371 (N_3371,In_51,In_978);
nor U3372 (N_3372,In_380,In_1317);
and U3373 (N_3373,In_577,In_746);
xnor U3374 (N_3374,In_615,In_321);
and U3375 (N_3375,In_614,In_473);
xor U3376 (N_3376,In_323,In_145);
or U3377 (N_3377,In_525,In_27);
xor U3378 (N_3378,In_1135,In_1777);
or U3379 (N_3379,In_1724,In_1567);
and U3380 (N_3380,In_843,In_1169);
xor U3381 (N_3381,In_1817,In_158);
nor U3382 (N_3382,In_595,In_1654);
nand U3383 (N_3383,In_1704,In_712);
nor U3384 (N_3384,In_1175,In_561);
and U3385 (N_3385,In_1849,In_917);
xor U3386 (N_3386,In_1607,In_1037);
nor U3387 (N_3387,In_584,In_705);
nand U3388 (N_3388,In_72,In_1186);
xor U3389 (N_3389,In_1065,In_319);
xnor U3390 (N_3390,In_1380,In_485);
xor U3391 (N_3391,In_1386,In_858);
and U3392 (N_3392,In_28,In_1788);
nor U3393 (N_3393,In_1588,In_1950);
or U3394 (N_3394,In_816,In_1645);
nor U3395 (N_3395,In_1955,In_1666);
xor U3396 (N_3396,In_1951,In_1846);
or U3397 (N_3397,In_1683,In_335);
nand U3398 (N_3398,In_399,In_474);
and U3399 (N_3399,In_1549,In_1466);
nor U3400 (N_3400,In_984,In_1809);
nand U3401 (N_3401,In_1643,In_746);
nor U3402 (N_3402,In_1089,In_1720);
or U3403 (N_3403,In_86,In_1935);
nand U3404 (N_3404,In_877,In_1504);
nand U3405 (N_3405,In_1386,In_293);
xor U3406 (N_3406,In_1471,In_1666);
nand U3407 (N_3407,In_777,In_318);
nand U3408 (N_3408,In_932,In_1798);
and U3409 (N_3409,In_1440,In_1494);
nand U3410 (N_3410,In_1267,In_1197);
or U3411 (N_3411,In_331,In_1747);
nand U3412 (N_3412,In_791,In_1042);
and U3413 (N_3413,In_1306,In_1445);
nand U3414 (N_3414,In_1543,In_112);
nor U3415 (N_3415,In_1974,In_1032);
nand U3416 (N_3416,In_727,In_1941);
or U3417 (N_3417,In_766,In_1381);
or U3418 (N_3418,In_1393,In_1461);
or U3419 (N_3419,In_781,In_454);
nand U3420 (N_3420,In_1187,In_1589);
nand U3421 (N_3421,In_954,In_1760);
xor U3422 (N_3422,In_811,In_585);
nor U3423 (N_3423,In_1319,In_1301);
or U3424 (N_3424,In_353,In_1708);
and U3425 (N_3425,In_1807,In_1871);
nand U3426 (N_3426,In_388,In_1053);
and U3427 (N_3427,In_987,In_66);
nor U3428 (N_3428,In_1300,In_7);
or U3429 (N_3429,In_126,In_1396);
xor U3430 (N_3430,In_1063,In_1978);
xor U3431 (N_3431,In_1308,In_279);
or U3432 (N_3432,In_701,In_277);
xor U3433 (N_3433,In_1995,In_889);
and U3434 (N_3434,In_1195,In_1462);
nand U3435 (N_3435,In_1640,In_171);
nand U3436 (N_3436,In_636,In_1523);
nor U3437 (N_3437,In_440,In_1017);
xor U3438 (N_3438,In_1226,In_1021);
xnor U3439 (N_3439,In_1677,In_4);
xnor U3440 (N_3440,In_758,In_544);
nand U3441 (N_3441,In_1679,In_1778);
or U3442 (N_3442,In_548,In_467);
or U3443 (N_3443,In_1433,In_1078);
or U3444 (N_3444,In_757,In_935);
nor U3445 (N_3445,In_1446,In_563);
and U3446 (N_3446,In_1925,In_1538);
nor U3447 (N_3447,In_1662,In_324);
and U3448 (N_3448,In_1955,In_970);
nand U3449 (N_3449,In_132,In_1140);
xor U3450 (N_3450,In_790,In_1297);
nand U3451 (N_3451,In_265,In_70);
nor U3452 (N_3452,In_1818,In_717);
and U3453 (N_3453,In_922,In_586);
xor U3454 (N_3454,In_1195,In_1365);
xnor U3455 (N_3455,In_59,In_90);
nand U3456 (N_3456,In_1837,In_1679);
nor U3457 (N_3457,In_1618,In_642);
and U3458 (N_3458,In_562,In_376);
and U3459 (N_3459,In_660,In_938);
nor U3460 (N_3460,In_805,In_780);
nor U3461 (N_3461,In_1745,In_692);
nor U3462 (N_3462,In_654,In_1451);
nand U3463 (N_3463,In_462,In_696);
and U3464 (N_3464,In_1892,In_1785);
nand U3465 (N_3465,In_463,In_848);
nand U3466 (N_3466,In_654,In_513);
xor U3467 (N_3467,In_1907,In_599);
and U3468 (N_3468,In_206,In_1214);
nor U3469 (N_3469,In_1532,In_900);
nor U3470 (N_3470,In_984,In_1187);
nand U3471 (N_3471,In_1128,In_430);
nor U3472 (N_3472,In_1549,In_97);
and U3473 (N_3473,In_830,In_1302);
or U3474 (N_3474,In_708,In_67);
nor U3475 (N_3475,In_91,In_165);
xnor U3476 (N_3476,In_617,In_1678);
xor U3477 (N_3477,In_1593,In_482);
and U3478 (N_3478,In_1324,In_707);
nor U3479 (N_3479,In_1944,In_950);
nand U3480 (N_3480,In_1654,In_96);
nand U3481 (N_3481,In_476,In_1847);
or U3482 (N_3482,In_1179,In_1389);
nand U3483 (N_3483,In_1582,In_1672);
xor U3484 (N_3484,In_919,In_590);
nor U3485 (N_3485,In_123,In_1256);
xor U3486 (N_3486,In_96,In_925);
or U3487 (N_3487,In_1038,In_1774);
or U3488 (N_3488,In_1110,In_27);
and U3489 (N_3489,In_422,In_318);
nor U3490 (N_3490,In_540,In_970);
and U3491 (N_3491,In_1719,In_1590);
nand U3492 (N_3492,In_146,In_116);
nor U3493 (N_3493,In_1876,In_0);
and U3494 (N_3494,In_1846,In_1752);
nor U3495 (N_3495,In_84,In_879);
and U3496 (N_3496,In_275,In_1301);
or U3497 (N_3497,In_454,In_971);
xor U3498 (N_3498,In_803,In_1243);
or U3499 (N_3499,In_1103,In_1518);
nand U3500 (N_3500,In_1664,In_1560);
xor U3501 (N_3501,In_1106,In_1509);
and U3502 (N_3502,In_383,In_1253);
and U3503 (N_3503,In_1323,In_434);
nand U3504 (N_3504,In_86,In_1971);
or U3505 (N_3505,In_1117,In_899);
and U3506 (N_3506,In_132,In_63);
nor U3507 (N_3507,In_839,In_330);
nor U3508 (N_3508,In_1950,In_1366);
or U3509 (N_3509,In_465,In_173);
nand U3510 (N_3510,In_1222,In_1056);
nand U3511 (N_3511,In_1503,In_1787);
nand U3512 (N_3512,In_764,In_454);
or U3513 (N_3513,In_1864,In_533);
nor U3514 (N_3514,In_1194,In_1700);
and U3515 (N_3515,In_1794,In_681);
and U3516 (N_3516,In_759,In_988);
nand U3517 (N_3517,In_1953,In_1784);
xor U3518 (N_3518,In_1944,In_1323);
or U3519 (N_3519,In_840,In_1057);
and U3520 (N_3520,In_509,In_575);
or U3521 (N_3521,In_1082,In_109);
nand U3522 (N_3522,In_415,In_624);
xor U3523 (N_3523,In_1835,In_845);
nand U3524 (N_3524,In_916,In_734);
nor U3525 (N_3525,In_1348,In_1961);
nand U3526 (N_3526,In_233,In_1687);
and U3527 (N_3527,In_379,In_1853);
nor U3528 (N_3528,In_1034,In_133);
nor U3529 (N_3529,In_555,In_899);
and U3530 (N_3530,In_550,In_928);
xnor U3531 (N_3531,In_1504,In_1674);
nand U3532 (N_3532,In_1799,In_1466);
xnor U3533 (N_3533,In_327,In_1487);
or U3534 (N_3534,In_971,In_1809);
nor U3535 (N_3535,In_287,In_76);
and U3536 (N_3536,In_1539,In_1689);
or U3537 (N_3537,In_599,In_104);
nor U3538 (N_3538,In_1422,In_133);
nor U3539 (N_3539,In_1702,In_367);
nor U3540 (N_3540,In_1728,In_1537);
xor U3541 (N_3541,In_1170,In_1239);
nor U3542 (N_3542,In_1648,In_1723);
and U3543 (N_3543,In_1121,In_325);
and U3544 (N_3544,In_1238,In_1545);
nand U3545 (N_3545,In_1483,In_410);
or U3546 (N_3546,In_1691,In_995);
and U3547 (N_3547,In_1976,In_885);
nand U3548 (N_3548,In_1889,In_1182);
nand U3549 (N_3549,In_274,In_573);
and U3550 (N_3550,In_1716,In_1907);
and U3551 (N_3551,In_74,In_1154);
nand U3552 (N_3552,In_1486,In_1114);
and U3553 (N_3553,In_1269,In_1101);
nand U3554 (N_3554,In_1457,In_455);
or U3555 (N_3555,In_826,In_1672);
and U3556 (N_3556,In_1305,In_1594);
nand U3557 (N_3557,In_1350,In_834);
and U3558 (N_3558,In_709,In_1426);
nand U3559 (N_3559,In_559,In_384);
nand U3560 (N_3560,In_1875,In_1980);
and U3561 (N_3561,In_534,In_311);
or U3562 (N_3562,In_603,In_463);
nor U3563 (N_3563,In_1763,In_1407);
or U3564 (N_3564,In_1438,In_1979);
nand U3565 (N_3565,In_495,In_612);
xnor U3566 (N_3566,In_1081,In_897);
nand U3567 (N_3567,In_714,In_203);
or U3568 (N_3568,In_883,In_867);
or U3569 (N_3569,In_1364,In_433);
nor U3570 (N_3570,In_1057,In_1441);
or U3571 (N_3571,In_905,In_1161);
nor U3572 (N_3572,In_235,In_150);
nor U3573 (N_3573,In_1350,In_724);
xnor U3574 (N_3574,In_293,In_783);
nor U3575 (N_3575,In_686,In_329);
and U3576 (N_3576,In_455,In_1905);
nand U3577 (N_3577,In_311,In_413);
or U3578 (N_3578,In_1925,In_674);
and U3579 (N_3579,In_131,In_1188);
nand U3580 (N_3580,In_95,In_1264);
and U3581 (N_3581,In_1874,In_275);
xnor U3582 (N_3582,In_291,In_444);
and U3583 (N_3583,In_1596,In_848);
xor U3584 (N_3584,In_1101,In_301);
and U3585 (N_3585,In_1662,In_1308);
nand U3586 (N_3586,In_385,In_1959);
and U3587 (N_3587,In_561,In_1737);
xor U3588 (N_3588,In_213,In_1668);
and U3589 (N_3589,In_1980,In_1940);
nor U3590 (N_3590,In_1424,In_406);
nand U3591 (N_3591,In_1237,In_1385);
and U3592 (N_3592,In_399,In_208);
nor U3593 (N_3593,In_307,In_438);
nand U3594 (N_3594,In_1752,In_1968);
nor U3595 (N_3595,In_167,In_1028);
and U3596 (N_3596,In_1959,In_1815);
nand U3597 (N_3597,In_804,In_1253);
xor U3598 (N_3598,In_1105,In_3);
and U3599 (N_3599,In_1421,In_1723);
xor U3600 (N_3600,In_1394,In_700);
and U3601 (N_3601,In_273,In_1448);
nor U3602 (N_3602,In_1759,In_1477);
nand U3603 (N_3603,In_1827,In_366);
xor U3604 (N_3604,In_1703,In_345);
nand U3605 (N_3605,In_1954,In_1472);
or U3606 (N_3606,In_1115,In_898);
nor U3607 (N_3607,In_1594,In_1332);
nor U3608 (N_3608,In_1134,In_1736);
or U3609 (N_3609,In_1903,In_1046);
nor U3610 (N_3610,In_75,In_1139);
nand U3611 (N_3611,In_1996,In_1922);
or U3612 (N_3612,In_1141,In_1972);
nand U3613 (N_3613,In_973,In_340);
nor U3614 (N_3614,In_146,In_1624);
or U3615 (N_3615,In_96,In_562);
nor U3616 (N_3616,In_149,In_58);
and U3617 (N_3617,In_334,In_1168);
and U3618 (N_3618,In_1272,In_845);
nor U3619 (N_3619,In_867,In_1357);
nor U3620 (N_3620,In_1923,In_1290);
xor U3621 (N_3621,In_1285,In_845);
xor U3622 (N_3622,In_357,In_915);
nor U3623 (N_3623,In_275,In_862);
and U3624 (N_3624,In_110,In_648);
nand U3625 (N_3625,In_685,In_1503);
xnor U3626 (N_3626,In_309,In_1396);
and U3627 (N_3627,In_450,In_1452);
nand U3628 (N_3628,In_849,In_1533);
and U3629 (N_3629,In_1451,In_1856);
or U3630 (N_3630,In_173,In_379);
nand U3631 (N_3631,In_1451,In_105);
or U3632 (N_3632,In_216,In_344);
xnor U3633 (N_3633,In_15,In_1019);
xnor U3634 (N_3634,In_365,In_1616);
or U3635 (N_3635,In_1349,In_1831);
or U3636 (N_3636,In_547,In_1964);
xnor U3637 (N_3637,In_724,In_1466);
xnor U3638 (N_3638,In_10,In_796);
nor U3639 (N_3639,In_1571,In_1406);
xor U3640 (N_3640,In_1470,In_243);
and U3641 (N_3641,In_28,In_1194);
and U3642 (N_3642,In_1364,In_1759);
and U3643 (N_3643,In_510,In_1346);
nand U3644 (N_3644,In_1907,In_113);
or U3645 (N_3645,In_1188,In_395);
xnor U3646 (N_3646,In_1364,In_887);
xnor U3647 (N_3647,In_845,In_710);
or U3648 (N_3648,In_1152,In_622);
nor U3649 (N_3649,In_495,In_1317);
nand U3650 (N_3650,In_1027,In_148);
and U3651 (N_3651,In_109,In_207);
xnor U3652 (N_3652,In_983,In_1347);
nand U3653 (N_3653,In_655,In_772);
xor U3654 (N_3654,In_1760,In_1109);
and U3655 (N_3655,In_427,In_527);
or U3656 (N_3656,In_27,In_933);
xnor U3657 (N_3657,In_1997,In_807);
and U3658 (N_3658,In_616,In_1514);
xor U3659 (N_3659,In_147,In_62);
or U3660 (N_3660,In_1526,In_327);
or U3661 (N_3661,In_61,In_1429);
nand U3662 (N_3662,In_1009,In_546);
nor U3663 (N_3663,In_284,In_626);
nor U3664 (N_3664,In_850,In_1121);
xnor U3665 (N_3665,In_258,In_643);
xor U3666 (N_3666,In_242,In_1529);
or U3667 (N_3667,In_116,In_783);
and U3668 (N_3668,In_348,In_936);
nand U3669 (N_3669,In_1984,In_748);
and U3670 (N_3670,In_645,In_1490);
and U3671 (N_3671,In_375,In_349);
or U3672 (N_3672,In_1821,In_571);
xor U3673 (N_3673,In_1331,In_1263);
nand U3674 (N_3674,In_63,In_1517);
nand U3675 (N_3675,In_155,In_1740);
or U3676 (N_3676,In_724,In_1117);
and U3677 (N_3677,In_1684,In_445);
nand U3678 (N_3678,In_1904,In_22);
and U3679 (N_3679,In_184,In_589);
nand U3680 (N_3680,In_1003,In_1462);
nand U3681 (N_3681,In_210,In_902);
nand U3682 (N_3682,In_876,In_671);
and U3683 (N_3683,In_1790,In_1424);
xnor U3684 (N_3684,In_1180,In_1275);
or U3685 (N_3685,In_924,In_1456);
or U3686 (N_3686,In_674,In_1089);
nand U3687 (N_3687,In_1727,In_1587);
nand U3688 (N_3688,In_1616,In_168);
and U3689 (N_3689,In_1183,In_477);
and U3690 (N_3690,In_1332,In_597);
nand U3691 (N_3691,In_1899,In_1286);
nor U3692 (N_3692,In_1208,In_1755);
nand U3693 (N_3693,In_1280,In_1126);
and U3694 (N_3694,In_840,In_468);
xor U3695 (N_3695,In_1186,In_1124);
xor U3696 (N_3696,In_129,In_1698);
and U3697 (N_3697,In_350,In_1854);
and U3698 (N_3698,In_1721,In_1776);
and U3699 (N_3699,In_589,In_1669);
xor U3700 (N_3700,In_70,In_804);
nand U3701 (N_3701,In_707,In_318);
or U3702 (N_3702,In_520,In_302);
xor U3703 (N_3703,In_9,In_1463);
and U3704 (N_3704,In_1435,In_511);
nand U3705 (N_3705,In_636,In_1081);
or U3706 (N_3706,In_1442,In_1528);
and U3707 (N_3707,In_1077,In_225);
nand U3708 (N_3708,In_1766,In_1876);
and U3709 (N_3709,In_355,In_1012);
xnor U3710 (N_3710,In_1118,In_712);
and U3711 (N_3711,In_1769,In_1558);
and U3712 (N_3712,In_1039,In_970);
nor U3713 (N_3713,In_1397,In_440);
and U3714 (N_3714,In_1517,In_1745);
nand U3715 (N_3715,In_149,In_231);
nand U3716 (N_3716,In_1080,In_1702);
and U3717 (N_3717,In_1602,In_473);
nor U3718 (N_3718,In_894,In_915);
or U3719 (N_3719,In_1863,In_1289);
nor U3720 (N_3720,In_446,In_1601);
or U3721 (N_3721,In_356,In_1376);
or U3722 (N_3722,In_759,In_1301);
nand U3723 (N_3723,In_1210,In_1800);
nor U3724 (N_3724,In_1465,In_1056);
nor U3725 (N_3725,In_1997,In_282);
xor U3726 (N_3726,In_640,In_692);
nand U3727 (N_3727,In_428,In_1752);
nor U3728 (N_3728,In_663,In_527);
nor U3729 (N_3729,In_520,In_160);
or U3730 (N_3730,In_379,In_1421);
nor U3731 (N_3731,In_997,In_1634);
or U3732 (N_3732,In_888,In_684);
nor U3733 (N_3733,In_337,In_948);
or U3734 (N_3734,In_1376,In_891);
or U3735 (N_3735,In_718,In_1280);
or U3736 (N_3736,In_1868,In_506);
and U3737 (N_3737,In_1518,In_464);
nor U3738 (N_3738,In_705,In_1137);
xnor U3739 (N_3739,In_388,In_470);
and U3740 (N_3740,In_281,In_241);
or U3741 (N_3741,In_223,In_1190);
xor U3742 (N_3742,In_149,In_43);
nand U3743 (N_3743,In_1559,In_1838);
or U3744 (N_3744,In_1148,In_972);
nor U3745 (N_3745,In_136,In_1170);
nor U3746 (N_3746,In_1942,In_1173);
nor U3747 (N_3747,In_1809,In_737);
nor U3748 (N_3748,In_920,In_229);
nand U3749 (N_3749,In_1912,In_1245);
xnor U3750 (N_3750,In_677,In_1426);
and U3751 (N_3751,In_506,In_944);
xnor U3752 (N_3752,In_980,In_719);
nor U3753 (N_3753,In_1776,In_824);
or U3754 (N_3754,In_372,In_736);
xor U3755 (N_3755,In_875,In_394);
and U3756 (N_3756,In_894,In_1594);
or U3757 (N_3757,In_185,In_1872);
or U3758 (N_3758,In_1816,In_367);
xor U3759 (N_3759,In_1979,In_1200);
xnor U3760 (N_3760,In_709,In_1036);
or U3761 (N_3761,In_1280,In_882);
nand U3762 (N_3762,In_1639,In_566);
nand U3763 (N_3763,In_1863,In_932);
nor U3764 (N_3764,In_754,In_1302);
nand U3765 (N_3765,In_949,In_651);
nand U3766 (N_3766,In_261,In_403);
xnor U3767 (N_3767,In_1360,In_1001);
nand U3768 (N_3768,In_1110,In_1374);
nand U3769 (N_3769,In_173,In_962);
xnor U3770 (N_3770,In_92,In_1387);
or U3771 (N_3771,In_1430,In_133);
or U3772 (N_3772,In_192,In_1081);
nor U3773 (N_3773,In_1834,In_1576);
xnor U3774 (N_3774,In_1561,In_796);
nor U3775 (N_3775,In_1987,In_1460);
xnor U3776 (N_3776,In_677,In_904);
or U3777 (N_3777,In_89,In_894);
or U3778 (N_3778,In_844,In_1948);
nor U3779 (N_3779,In_1427,In_243);
xnor U3780 (N_3780,In_558,In_736);
or U3781 (N_3781,In_1543,In_550);
and U3782 (N_3782,In_1457,In_1543);
and U3783 (N_3783,In_735,In_1387);
nor U3784 (N_3784,In_1422,In_315);
xor U3785 (N_3785,In_999,In_610);
xor U3786 (N_3786,In_1887,In_420);
nand U3787 (N_3787,In_709,In_1766);
nor U3788 (N_3788,In_369,In_583);
nand U3789 (N_3789,In_1215,In_761);
and U3790 (N_3790,In_142,In_1458);
or U3791 (N_3791,In_1831,In_1447);
xor U3792 (N_3792,In_1985,In_25);
nand U3793 (N_3793,In_280,In_466);
nand U3794 (N_3794,In_126,In_1089);
nor U3795 (N_3795,In_373,In_1320);
nor U3796 (N_3796,In_1846,In_589);
or U3797 (N_3797,In_1809,In_804);
or U3798 (N_3798,In_1924,In_1887);
nand U3799 (N_3799,In_752,In_206);
or U3800 (N_3800,In_87,In_868);
nor U3801 (N_3801,In_1678,In_740);
and U3802 (N_3802,In_1185,In_1028);
nand U3803 (N_3803,In_553,In_1516);
and U3804 (N_3804,In_548,In_608);
nor U3805 (N_3805,In_1401,In_462);
nor U3806 (N_3806,In_776,In_84);
nor U3807 (N_3807,In_823,In_1852);
and U3808 (N_3808,In_1349,In_1927);
nor U3809 (N_3809,In_804,In_313);
or U3810 (N_3810,In_1095,In_14);
nor U3811 (N_3811,In_874,In_1517);
nand U3812 (N_3812,In_1627,In_1943);
or U3813 (N_3813,In_309,In_1383);
and U3814 (N_3814,In_757,In_698);
nor U3815 (N_3815,In_1434,In_1555);
nand U3816 (N_3816,In_1807,In_1090);
nand U3817 (N_3817,In_1900,In_194);
or U3818 (N_3818,In_903,In_74);
and U3819 (N_3819,In_1704,In_680);
xor U3820 (N_3820,In_1559,In_779);
nor U3821 (N_3821,In_425,In_1628);
or U3822 (N_3822,In_196,In_1711);
nand U3823 (N_3823,In_513,In_1541);
or U3824 (N_3824,In_981,In_550);
nor U3825 (N_3825,In_1025,In_1263);
or U3826 (N_3826,In_1573,In_984);
or U3827 (N_3827,In_475,In_1719);
xor U3828 (N_3828,In_610,In_947);
xor U3829 (N_3829,In_69,In_1044);
nor U3830 (N_3830,In_1852,In_441);
nand U3831 (N_3831,In_1483,In_1172);
or U3832 (N_3832,In_482,In_869);
or U3833 (N_3833,In_990,In_1062);
xor U3834 (N_3834,In_1201,In_661);
xnor U3835 (N_3835,In_1550,In_520);
xor U3836 (N_3836,In_855,In_285);
or U3837 (N_3837,In_185,In_963);
xnor U3838 (N_3838,In_561,In_1674);
xnor U3839 (N_3839,In_1621,In_1310);
or U3840 (N_3840,In_635,In_701);
nor U3841 (N_3841,In_1717,In_1788);
nor U3842 (N_3842,In_1659,In_1986);
xor U3843 (N_3843,In_775,In_720);
xor U3844 (N_3844,In_62,In_1496);
and U3845 (N_3845,In_505,In_608);
and U3846 (N_3846,In_681,In_1463);
or U3847 (N_3847,In_1140,In_1241);
xor U3848 (N_3848,In_949,In_1447);
and U3849 (N_3849,In_1414,In_410);
nand U3850 (N_3850,In_370,In_44);
nor U3851 (N_3851,In_1237,In_327);
xnor U3852 (N_3852,In_1458,In_1642);
nand U3853 (N_3853,In_432,In_1440);
xnor U3854 (N_3854,In_126,In_20);
nor U3855 (N_3855,In_1609,In_426);
or U3856 (N_3856,In_1201,In_1103);
or U3857 (N_3857,In_398,In_1201);
nand U3858 (N_3858,In_742,In_853);
and U3859 (N_3859,In_1985,In_1687);
xnor U3860 (N_3860,In_967,In_581);
or U3861 (N_3861,In_1558,In_173);
and U3862 (N_3862,In_483,In_635);
and U3863 (N_3863,In_1140,In_1245);
or U3864 (N_3864,In_291,In_1510);
xnor U3865 (N_3865,In_540,In_188);
nor U3866 (N_3866,In_1064,In_1009);
or U3867 (N_3867,In_1536,In_1925);
nand U3868 (N_3868,In_1267,In_485);
xnor U3869 (N_3869,In_1327,In_1735);
nor U3870 (N_3870,In_1274,In_8);
and U3871 (N_3871,In_1344,In_1243);
or U3872 (N_3872,In_722,In_51);
xor U3873 (N_3873,In_738,In_1333);
nand U3874 (N_3874,In_1866,In_1683);
nand U3875 (N_3875,In_1416,In_978);
nand U3876 (N_3876,In_323,In_1983);
nand U3877 (N_3877,In_1328,In_1530);
and U3878 (N_3878,In_861,In_1683);
or U3879 (N_3879,In_617,In_1655);
nor U3880 (N_3880,In_1002,In_1281);
xor U3881 (N_3881,In_1045,In_1311);
xnor U3882 (N_3882,In_1719,In_75);
and U3883 (N_3883,In_345,In_948);
nand U3884 (N_3884,In_22,In_1509);
nand U3885 (N_3885,In_964,In_1505);
and U3886 (N_3886,In_696,In_417);
nand U3887 (N_3887,In_1080,In_78);
or U3888 (N_3888,In_525,In_1499);
or U3889 (N_3889,In_796,In_1461);
xnor U3890 (N_3890,In_1737,In_1029);
xor U3891 (N_3891,In_1163,In_879);
xor U3892 (N_3892,In_30,In_1578);
xor U3893 (N_3893,In_1792,In_449);
or U3894 (N_3894,In_594,In_1728);
xnor U3895 (N_3895,In_544,In_1904);
nor U3896 (N_3896,In_1119,In_284);
nand U3897 (N_3897,In_1220,In_1438);
or U3898 (N_3898,In_504,In_1053);
nor U3899 (N_3899,In_1237,In_460);
or U3900 (N_3900,In_1089,In_1108);
xor U3901 (N_3901,In_951,In_332);
and U3902 (N_3902,In_50,In_1822);
nand U3903 (N_3903,In_1351,In_665);
and U3904 (N_3904,In_1577,In_248);
nand U3905 (N_3905,In_1402,In_70);
or U3906 (N_3906,In_915,In_762);
nor U3907 (N_3907,In_230,In_1695);
and U3908 (N_3908,In_297,In_594);
and U3909 (N_3909,In_447,In_362);
nand U3910 (N_3910,In_1070,In_1290);
or U3911 (N_3911,In_411,In_1791);
xnor U3912 (N_3912,In_1346,In_914);
or U3913 (N_3913,In_1958,In_872);
or U3914 (N_3914,In_202,In_1971);
nor U3915 (N_3915,In_814,In_596);
nand U3916 (N_3916,In_827,In_17);
nor U3917 (N_3917,In_1286,In_764);
and U3918 (N_3918,In_104,In_1503);
nor U3919 (N_3919,In_562,In_754);
and U3920 (N_3920,In_765,In_932);
and U3921 (N_3921,In_1634,In_562);
nor U3922 (N_3922,In_1574,In_1863);
and U3923 (N_3923,In_701,In_929);
nor U3924 (N_3924,In_1375,In_371);
xnor U3925 (N_3925,In_1671,In_1456);
nand U3926 (N_3926,In_1604,In_771);
xor U3927 (N_3927,In_1898,In_1419);
xor U3928 (N_3928,In_1807,In_96);
nor U3929 (N_3929,In_1585,In_209);
and U3930 (N_3930,In_1150,In_1700);
xor U3931 (N_3931,In_233,In_1285);
nand U3932 (N_3932,In_982,In_251);
or U3933 (N_3933,In_960,In_1600);
and U3934 (N_3934,In_412,In_1354);
nor U3935 (N_3935,In_1466,In_1578);
nand U3936 (N_3936,In_1150,In_1157);
xnor U3937 (N_3937,In_1477,In_1721);
nor U3938 (N_3938,In_807,In_1968);
and U3939 (N_3939,In_1477,In_1740);
nand U3940 (N_3940,In_121,In_451);
nor U3941 (N_3941,In_1370,In_289);
nor U3942 (N_3942,In_1482,In_1993);
and U3943 (N_3943,In_1358,In_1630);
xnor U3944 (N_3944,In_1553,In_1378);
nand U3945 (N_3945,In_1989,In_981);
xnor U3946 (N_3946,In_181,In_1690);
xor U3947 (N_3947,In_862,In_264);
nand U3948 (N_3948,In_942,In_487);
xor U3949 (N_3949,In_690,In_596);
nor U3950 (N_3950,In_755,In_270);
nor U3951 (N_3951,In_623,In_296);
and U3952 (N_3952,In_676,In_547);
and U3953 (N_3953,In_558,In_403);
and U3954 (N_3954,In_169,In_602);
nand U3955 (N_3955,In_1304,In_1297);
nor U3956 (N_3956,In_1522,In_1658);
nand U3957 (N_3957,In_1177,In_1002);
or U3958 (N_3958,In_472,In_1287);
or U3959 (N_3959,In_1707,In_1877);
xnor U3960 (N_3960,In_948,In_1126);
nand U3961 (N_3961,In_1218,In_1245);
or U3962 (N_3962,In_1940,In_1366);
and U3963 (N_3963,In_162,In_955);
xnor U3964 (N_3964,In_1369,In_1639);
and U3965 (N_3965,In_239,In_855);
nor U3966 (N_3966,In_439,In_638);
and U3967 (N_3967,In_1743,In_1307);
nand U3968 (N_3968,In_750,In_1768);
nor U3969 (N_3969,In_1140,In_342);
or U3970 (N_3970,In_810,In_93);
xor U3971 (N_3971,In_1141,In_51);
and U3972 (N_3972,In_658,In_555);
xnor U3973 (N_3973,In_1432,In_371);
or U3974 (N_3974,In_1973,In_1428);
nand U3975 (N_3975,In_523,In_846);
xnor U3976 (N_3976,In_1222,In_804);
nor U3977 (N_3977,In_1882,In_1326);
nand U3978 (N_3978,In_382,In_968);
nand U3979 (N_3979,In_1561,In_1396);
and U3980 (N_3980,In_432,In_705);
or U3981 (N_3981,In_747,In_1839);
xnor U3982 (N_3982,In_1200,In_1167);
nand U3983 (N_3983,In_88,In_547);
nor U3984 (N_3984,In_1861,In_1637);
nand U3985 (N_3985,In_391,In_1);
and U3986 (N_3986,In_1300,In_288);
or U3987 (N_3987,In_929,In_1580);
and U3988 (N_3988,In_591,In_572);
nand U3989 (N_3989,In_1509,In_1314);
nand U3990 (N_3990,In_1854,In_772);
or U3991 (N_3991,In_1572,In_758);
and U3992 (N_3992,In_1985,In_1009);
nand U3993 (N_3993,In_639,In_785);
or U3994 (N_3994,In_165,In_1599);
and U3995 (N_3995,In_92,In_659);
nand U3996 (N_3996,In_1796,In_1281);
xnor U3997 (N_3997,In_1750,In_1773);
nor U3998 (N_3998,In_293,In_709);
xnor U3999 (N_3999,In_1217,In_668);
nand U4000 (N_4000,N_2202,N_1763);
nor U4001 (N_4001,N_3820,N_3481);
nor U4002 (N_4002,N_48,N_2314);
nand U4003 (N_4003,N_3065,N_3279);
nand U4004 (N_4004,N_2976,N_1233);
and U4005 (N_4005,N_1511,N_3423);
nand U4006 (N_4006,N_555,N_1813);
nand U4007 (N_4007,N_2626,N_136);
xnor U4008 (N_4008,N_3497,N_3074);
nand U4009 (N_4009,N_3232,N_1135);
xnor U4010 (N_4010,N_2258,N_2718);
nand U4011 (N_4011,N_2520,N_1873);
xor U4012 (N_4012,N_3957,N_3321);
xor U4013 (N_4013,N_91,N_2483);
or U4014 (N_4014,N_1319,N_1426);
nor U4015 (N_4015,N_1288,N_1333);
nor U4016 (N_4016,N_2195,N_353);
or U4017 (N_4017,N_3499,N_2814);
and U4018 (N_4018,N_179,N_776);
xnor U4019 (N_4019,N_2201,N_1057);
nor U4020 (N_4020,N_1651,N_2822);
nor U4021 (N_4021,N_1356,N_2405);
nand U4022 (N_4022,N_3688,N_2186);
nor U4023 (N_4023,N_3454,N_2431);
nor U4024 (N_4024,N_1568,N_2940);
nand U4025 (N_4025,N_721,N_3160);
xor U4026 (N_4026,N_1263,N_3652);
or U4027 (N_4027,N_676,N_1852);
xor U4028 (N_4028,N_2671,N_2500);
nor U4029 (N_4029,N_1343,N_838);
xor U4030 (N_4030,N_2825,N_12);
and U4031 (N_4031,N_1876,N_1848);
xor U4032 (N_4032,N_273,N_380);
or U4033 (N_4033,N_3048,N_2459);
nor U4034 (N_4034,N_1614,N_2119);
or U4035 (N_4035,N_3143,N_1454);
xor U4036 (N_4036,N_115,N_3381);
xnor U4037 (N_4037,N_3139,N_3432);
nor U4038 (N_4038,N_3185,N_3617);
and U4039 (N_4039,N_2886,N_1579);
nor U4040 (N_4040,N_3811,N_531);
nor U4041 (N_4041,N_3162,N_149);
nand U4042 (N_4042,N_1087,N_469);
xor U4043 (N_4043,N_3534,N_1912);
and U4044 (N_4044,N_3782,N_228);
and U4045 (N_4045,N_2853,N_2439);
xnor U4046 (N_4046,N_2658,N_2245);
nand U4047 (N_4047,N_2710,N_3612);
xnor U4048 (N_4048,N_1108,N_794);
xor U4049 (N_4049,N_2582,N_3325);
nor U4050 (N_4050,N_3387,N_2329);
and U4051 (N_4051,N_2029,N_1257);
nand U4052 (N_4052,N_1727,N_29);
xnor U4053 (N_4053,N_3603,N_382);
nor U4054 (N_4054,N_967,N_1332);
xnor U4055 (N_4055,N_683,N_1141);
or U4056 (N_4056,N_3997,N_1715);
nand U4057 (N_4057,N_3837,N_3710);
nand U4058 (N_4058,N_2112,N_309);
xnor U4059 (N_4059,N_3177,N_522);
or U4060 (N_4060,N_3706,N_3707);
or U4061 (N_4061,N_537,N_597);
nor U4062 (N_4062,N_2184,N_1884);
and U4063 (N_4063,N_3470,N_2028);
nor U4064 (N_4064,N_2270,N_185);
nand U4065 (N_4065,N_3885,N_3240);
nor U4066 (N_4066,N_599,N_1311);
nand U4067 (N_4067,N_1793,N_3389);
xnor U4068 (N_4068,N_434,N_1053);
and U4069 (N_4069,N_2730,N_3701);
xnor U4070 (N_4070,N_3189,N_2930);
nor U4071 (N_4071,N_8,N_2999);
and U4072 (N_4072,N_2126,N_3463);
and U4073 (N_4073,N_411,N_2278);
nand U4074 (N_4074,N_884,N_1149);
nand U4075 (N_4075,N_548,N_880);
xnor U4076 (N_4076,N_1205,N_2952);
or U4077 (N_4077,N_3511,N_3646);
xnor U4078 (N_4078,N_253,N_231);
or U4079 (N_4079,N_1166,N_1880);
and U4080 (N_4080,N_2975,N_3639);
nor U4081 (N_4081,N_865,N_1939);
or U4082 (N_4082,N_644,N_3327);
xnor U4083 (N_4083,N_1812,N_2370);
nand U4084 (N_4084,N_2285,N_225);
and U4085 (N_4085,N_2792,N_1392);
nor U4086 (N_4086,N_515,N_367);
and U4087 (N_4087,N_3464,N_1637);
nand U4088 (N_4088,N_1602,N_3214);
or U4089 (N_4089,N_1353,N_1190);
nand U4090 (N_4090,N_337,N_1776);
and U4091 (N_4091,N_1713,N_874);
or U4092 (N_4092,N_2210,N_1497);
or U4093 (N_4093,N_2102,N_1393);
xnor U4094 (N_4094,N_685,N_2947);
nor U4095 (N_4095,N_1990,N_3451);
and U4096 (N_4096,N_10,N_1015);
nand U4097 (N_4097,N_1917,N_3097);
nor U4098 (N_4098,N_3219,N_2025);
and U4099 (N_4099,N_94,N_3952);
and U4100 (N_4100,N_453,N_2908);
or U4101 (N_4101,N_1847,N_361);
nor U4102 (N_4102,N_3072,N_1785);
nor U4103 (N_4103,N_2051,N_2824);
and U4104 (N_4104,N_3150,N_2239);
nand U4105 (N_4105,N_2386,N_3939);
nor U4106 (N_4106,N_412,N_3988);
nor U4107 (N_4107,N_2181,N_3248);
nor U4108 (N_4108,N_1951,N_2173);
nand U4109 (N_4109,N_1494,N_2523);
or U4110 (N_4110,N_1596,N_3153);
nand U4111 (N_4111,N_928,N_425);
nor U4112 (N_4112,N_3404,N_1611);
or U4113 (N_4113,N_2008,N_363);
xnor U4114 (N_4114,N_1978,N_2770);
or U4115 (N_4115,N_516,N_3204);
nand U4116 (N_4116,N_2113,N_2388);
nand U4117 (N_4117,N_1640,N_2951);
xnor U4118 (N_4118,N_197,N_1060);
nand U4119 (N_4119,N_2687,N_474);
nor U4120 (N_4120,N_3108,N_2396);
nor U4121 (N_4121,N_691,N_2701);
or U4122 (N_4122,N_2869,N_3426);
and U4123 (N_4123,N_1030,N_1928);
nor U4124 (N_4124,N_3370,N_593);
and U4125 (N_4125,N_3130,N_889);
nor U4126 (N_4126,N_1226,N_974);
nand U4127 (N_4127,N_3797,N_2636);
xnor U4128 (N_4128,N_3763,N_780);
xor U4129 (N_4129,N_2410,N_1883);
and U4130 (N_4130,N_1676,N_99);
nand U4131 (N_4131,N_2544,N_3880);
and U4132 (N_4132,N_965,N_3504);
xor U4133 (N_4133,N_2810,N_343);
and U4134 (N_4134,N_3604,N_1737);
nand U4135 (N_4135,N_362,N_2041);
xor U4136 (N_4136,N_3073,N_3347);
xnor U4137 (N_4137,N_3635,N_1164);
and U4138 (N_4138,N_3424,N_598);
xor U4139 (N_4139,N_3491,N_284);
and U4140 (N_4140,N_2514,N_752);
xor U4141 (N_4141,N_699,N_1224);
nand U4142 (N_4142,N_872,N_1790);
nor U4143 (N_4143,N_1496,N_2616);
xnor U4144 (N_4144,N_402,N_2859);
and U4145 (N_4145,N_3449,N_232);
or U4146 (N_4146,N_2489,N_3476);
and U4147 (N_4147,N_1133,N_1483);
or U4148 (N_4148,N_2120,N_1677);
nand U4149 (N_4149,N_1477,N_1758);
nor U4150 (N_4150,N_972,N_1703);
and U4151 (N_4151,N_1625,N_514);
xor U4152 (N_4152,N_2702,N_2358);
xnor U4153 (N_4153,N_1692,N_2654);
nor U4154 (N_4154,N_1368,N_3802);
nand U4155 (N_4155,N_3700,N_3902);
xnor U4156 (N_4156,N_1414,N_1932);
nor U4157 (N_4157,N_2958,N_1527);
and U4158 (N_4158,N_3538,N_1519);
xor U4159 (N_4159,N_1088,N_162);
nand U4160 (N_4160,N_2040,N_3188);
nor U4161 (N_4161,N_2602,N_3319);
and U4162 (N_4162,N_3758,N_1396);
nand U4163 (N_4163,N_3954,N_1449);
and U4164 (N_4164,N_3698,N_558);
or U4165 (N_4165,N_1838,N_3580);
and U4166 (N_4166,N_817,N_2033);
or U4167 (N_4167,N_1699,N_2921);
nor U4168 (N_4168,N_3228,N_366);
xnor U4169 (N_4169,N_1961,N_3658);
xnor U4170 (N_4170,N_1736,N_3172);
and U4171 (N_4171,N_1730,N_2129);
or U4172 (N_4172,N_619,N_881);
xor U4173 (N_4173,N_2594,N_244);
nand U4174 (N_4174,N_2457,N_1968);
nand U4175 (N_4175,N_1777,N_3436);
xor U4176 (N_4176,N_2864,N_2843);
or U4177 (N_4177,N_3391,N_415);
nor U4178 (N_4178,N_109,N_792);
xnor U4179 (N_4179,N_3402,N_1595);
xor U4180 (N_4180,N_2540,N_2623);
and U4181 (N_4181,N_3754,N_1992);
xnor U4182 (N_4182,N_2277,N_1362);
and U4183 (N_4183,N_3917,N_964);
xnor U4184 (N_4184,N_2346,N_3661);
and U4185 (N_4185,N_1706,N_1290);
and U4186 (N_4186,N_1276,N_523);
and U4187 (N_4187,N_3961,N_2093);
nand U4188 (N_4188,N_1977,N_3283);
nand U4189 (N_4189,N_499,N_3374);
xor U4190 (N_4190,N_2624,N_3779);
nand U4191 (N_4191,N_1336,N_845);
xor U4192 (N_4192,N_2024,N_2490);
nand U4193 (N_4193,N_3884,N_1153);
nand U4194 (N_4194,N_3765,N_3545);
and U4195 (N_4195,N_740,N_579);
xnor U4196 (N_4196,N_2087,N_525);
or U4197 (N_4197,N_2089,N_44);
and U4198 (N_4198,N_692,N_3574);
and U4199 (N_4199,N_3227,N_2234);
and U4200 (N_4200,N_1745,N_1533);
nand U4201 (N_4201,N_3618,N_1284);
and U4202 (N_4202,N_520,N_66);
nor U4203 (N_4203,N_1212,N_3846);
and U4204 (N_4204,N_132,N_2144);
nor U4205 (N_4205,N_782,N_2242);
nand U4206 (N_4206,N_1560,N_2746);
xnor U4207 (N_4207,N_2812,N_7);
nand U4208 (N_4208,N_121,N_3873);
xor U4209 (N_4209,N_1085,N_860);
and U4210 (N_4210,N_3577,N_1955);
xnor U4211 (N_4211,N_1804,N_941);
nand U4212 (N_4212,N_583,N_2620);
or U4213 (N_4213,N_2494,N_513);
or U4214 (N_4214,N_203,N_2989);
and U4215 (N_4215,N_1842,N_3103);
and U4216 (N_4216,N_496,N_2892);
or U4217 (N_4217,N_2456,N_639);
nand U4218 (N_4218,N_2121,N_1881);
nand U4219 (N_4219,N_2496,N_533);
nand U4220 (N_4220,N_1324,N_1514);
or U4221 (N_4221,N_2703,N_3082);
nand U4222 (N_4222,N_3662,N_3888);
or U4223 (N_4223,N_1856,N_870);
or U4224 (N_4224,N_1456,N_3516);
nand U4225 (N_4225,N_3026,N_2527);
xor U4226 (N_4226,N_2154,N_2114);
or U4227 (N_4227,N_2080,N_2668);
or U4228 (N_4228,N_1230,N_1757);
or U4229 (N_4229,N_3959,N_2414);
or U4230 (N_4230,N_3126,N_862);
xor U4231 (N_4231,N_191,N_171);
xnor U4232 (N_4232,N_3894,N_393);
nor U4233 (N_4233,N_3183,N_3443);
xnor U4234 (N_4234,N_1559,N_2092);
xnor U4235 (N_4235,N_3334,N_1399);
nor U4236 (N_4236,N_1517,N_1024);
xnor U4237 (N_4237,N_761,N_3627);
and U4238 (N_4238,N_71,N_1654);
nand U4239 (N_4239,N_2170,N_1075);
or U4240 (N_4240,N_2452,N_1582);
or U4241 (N_4241,N_3469,N_3487);
xor U4242 (N_4242,N_3774,N_113);
and U4243 (N_4243,N_3715,N_1524);
nor U4244 (N_4244,N_3909,N_604);
xnor U4245 (N_4245,N_1258,N_3863);
nand U4246 (N_4246,N_1644,N_2555);
nor U4247 (N_4247,N_2541,N_1780);
nand U4248 (N_4248,N_2798,N_3361);
and U4249 (N_4249,N_1464,N_3013);
xor U4250 (N_4250,N_1575,N_1033);
or U4251 (N_4251,N_2992,N_3777);
xnor U4252 (N_4252,N_2493,N_3025);
nor U4253 (N_4253,N_2592,N_3142);
or U4254 (N_4254,N_830,N_293);
and U4255 (N_4255,N_1253,N_1208);
nand U4256 (N_4256,N_1971,N_3019);
xor U4257 (N_4257,N_3290,N_1993);
nand U4258 (N_4258,N_1126,N_1427);
or U4259 (N_4259,N_3783,N_1753);
nor U4260 (N_4260,N_3507,N_1983);
nand U4261 (N_4261,N_2534,N_2529);
xor U4262 (N_4262,N_385,N_416);
xnor U4263 (N_4263,N_1283,N_317);
nand U4264 (N_4264,N_3216,N_128);
and U4265 (N_4265,N_748,N_760);
nand U4266 (N_4266,N_3641,N_1280);
nor U4267 (N_4267,N_652,N_1512);
nand U4268 (N_4268,N_2428,N_2614);
nor U4269 (N_4269,N_1416,N_3887);
nor U4270 (N_4270,N_2223,N_995);
or U4271 (N_4271,N_2364,N_950);
and U4272 (N_4272,N_2966,N_2572);
xor U4273 (N_4273,N_700,N_2505);
or U4274 (N_4274,N_1620,N_1530);
or U4275 (N_4275,N_694,N_485);
nand U4276 (N_4276,N_444,N_512);
nor U4277 (N_4277,N_3044,N_114);
nor U4278 (N_4278,N_1549,N_3995);
or U4279 (N_4279,N_569,N_247);
xor U4280 (N_4280,N_2332,N_3716);
nand U4281 (N_4281,N_3611,N_1980);
xnor U4282 (N_4282,N_1055,N_3889);
and U4283 (N_4283,N_3131,N_1443);
nand U4284 (N_4284,N_3000,N_14);
or U4285 (N_4285,N_1171,N_3007);
or U4286 (N_4286,N_1987,N_1272);
xnor U4287 (N_4287,N_2971,N_373);
xor U4288 (N_4288,N_1684,N_1781);
and U4289 (N_4289,N_2183,N_3831);
or U4290 (N_4290,N_511,N_1635);
nand U4291 (N_4291,N_2785,N_65);
nor U4292 (N_4292,N_2900,N_1342);
xor U4293 (N_4293,N_495,N_467);
xor U4294 (N_4294,N_3191,N_784);
xnor U4295 (N_4295,N_3137,N_357);
nand U4296 (N_4296,N_3704,N_1735);
nand U4297 (N_4297,N_3819,N_1120);
nor U4298 (N_4298,N_815,N_3650);
nor U4299 (N_4299,N_1448,N_2338);
or U4300 (N_4300,N_256,N_1937);
or U4301 (N_4301,N_3903,N_2235);
xor U4302 (N_4302,N_2969,N_2461);
and U4303 (N_4303,N_355,N_3647);
nor U4304 (N_4304,N_387,N_1236);
or U4305 (N_4305,N_3827,N_1066);
nor U4306 (N_4306,N_3259,N_3590);
nor U4307 (N_4307,N_725,N_3791);
nand U4308 (N_4308,N_3541,N_3182);
xor U4309 (N_4309,N_869,N_430);
and U4310 (N_4310,N_1222,N_1460);
or U4311 (N_4311,N_2495,N_2189);
or U4312 (N_4312,N_2728,N_1964);
xnor U4313 (N_4313,N_2401,N_1632);
xor U4314 (N_4314,N_3798,N_3267);
xnor U4315 (N_4315,N_996,N_897);
nor U4316 (N_4316,N_1282,N_2857);
and U4317 (N_4317,N_1437,N_1119);
or U4318 (N_4318,N_1587,N_111);
nand U4319 (N_4319,N_1138,N_2968);
nor U4320 (N_4320,N_3268,N_3942);
nand U4321 (N_4321,N_1307,N_1320);
xor U4322 (N_4322,N_2561,N_3586);
and U4323 (N_4323,N_2590,N_3023);
and U4324 (N_4324,N_2964,N_38);
and U4325 (N_4325,N_3212,N_2954);
nand U4326 (N_4326,N_3483,N_3292);
and U4327 (N_4327,N_2176,N_2330);
xnor U4328 (N_4328,N_1213,N_2221);
and U4329 (N_4329,N_803,N_1963);
nand U4330 (N_4330,N_1686,N_508);
nor U4331 (N_4331,N_539,N_2241);
xnor U4332 (N_4332,N_3123,N_1178);
nand U4333 (N_4333,N_647,N_2589);
nor U4334 (N_4334,N_2931,N_1092);
xnor U4335 (N_4335,N_648,N_3157);
nor U4336 (N_4336,N_606,N_2765);
xor U4337 (N_4337,N_1438,N_2497);
nand U4338 (N_4338,N_2054,N_1039);
or U4339 (N_4339,N_3333,N_768);
or U4340 (N_4340,N_313,N_535);
and U4341 (N_4341,N_2331,N_1729);
nor U4342 (N_4342,N_3466,N_820);
nand U4343 (N_4343,N_557,N_3281);
or U4344 (N_4344,N_46,N_751);
nor U4345 (N_4345,N_3064,N_1020);
nor U4346 (N_4346,N_2115,N_2509);
nand U4347 (N_4347,N_1982,N_2784);
xor U4348 (N_4348,N_876,N_1806);
nand U4349 (N_4349,N_1599,N_2984);
or U4350 (N_4350,N_3421,N_1146);
xor U4351 (N_4351,N_2191,N_3236);
nor U4352 (N_4352,N_1962,N_2586);
xnor U4353 (N_4353,N_2336,N_1931);
xnor U4354 (N_4354,N_167,N_2635);
and U4355 (N_4355,N_673,N_3061);
nand U4356 (N_4356,N_3757,N_1655);
nand U4357 (N_4357,N_3186,N_2284);
or U4358 (N_4358,N_476,N_1633);
and U4359 (N_4359,N_2875,N_1225);
nor U4360 (N_4360,N_2633,N_2848);
xor U4361 (N_4361,N_1136,N_1889);
xnor U4362 (N_4362,N_3824,N_1869);
and U4363 (N_4363,N_887,N_2665);
or U4364 (N_4364,N_2216,N_1503);
or U4365 (N_4365,N_2521,N_1664);
nand U4366 (N_4366,N_1246,N_1774);
nor U4367 (N_4367,N_1663,N_449);
or U4368 (N_4368,N_3736,N_1360);
and U4369 (N_4369,N_3723,N_1761);
nand U4370 (N_4370,N_566,N_3332);
nor U4371 (N_4371,N_1795,N_3645);
xor U4372 (N_4372,N_1026,N_33);
and U4373 (N_4373,N_3833,N_2103);
nor U4374 (N_4374,N_2829,N_3830);
nand U4375 (N_4375,N_2070,N_1613);
nor U4376 (N_4376,N_282,N_788);
and U4377 (N_4377,N_773,N_3572);
or U4378 (N_4378,N_427,N_505);
and U4379 (N_4379,N_1529,N_2874);
xor U4380 (N_4380,N_3222,N_1605);
xnor U4381 (N_4381,N_3242,N_1007);
and U4382 (N_4382,N_3843,N_2359);
nor U4383 (N_4383,N_3922,N_2741);
and U4384 (N_4384,N_1034,N_2383);
nand U4385 (N_4385,N_2427,N_369);
or U4386 (N_4386,N_438,N_3747);
or U4387 (N_4387,N_3835,N_3148);
xor U4388 (N_4388,N_728,N_3168);
nand U4389 (N_4389,N_1380,N_1771);
or U4390 (N_4390,N_2877,N_2532);
nand U4391 (N_4391,N_2168,N_2570);
nor U4392 (N_4392,N_1754,N_826);
nand U4393 (N_4393,N_2652,N_446);
and U4394 (N_4394,N_2716,N_3442);
nor U4395 (N_4395,N_3581,N_354);
and U4396 (N_4396,N_1447,N_85);
or U4397 (N_4397,N_3510,N_2122);
and U4398 (N_4398,N_2994,N_1124);
nor U4399 (N_4399,N_3394,N_1563);
or U4400 (N_4400,N_3866,N_3090);
nor U4401 (N_4401,N_1996,N_2982);
nor U4402 (N_4402,N_1834,N_3860);
nor U4403 (N_4403,N_1071,N_2946);
xnor U4404 (N_4404,N_359,N_3951);
xnor U4405 (N_4405,N_3050,N_473);
and U4406 (N_4406,N_2655,N_76);
and U4407 (N_4407,N_1310,N_1067);
xnor U4408 (N_4408,N_3931,N_3803);
or U4409 (N_4409,N_923,N_3339);
nor U4410 (N_4410,N_1418,N_223);
nor U4411 (N_4411,N_1286,N_2842);
xor U4412 (N_4412,N_3610,N_856);
xor U4413 (N_4413,N_2110,N_2883);
xor U4414 (N_4414,N_2898,N_3159);
or U4415 (N_4415,N_2981,N_1446);
and U4416 (N_4416,N_1231,N_1803);
xor U4417 (N_4417,N_3138,N_2904);
nand U4418 (N_4418,N_465,N_2193);
or U4419 (N_4419,N_3342,N_3468);
and U4420 (N_4420,N_3169,N_2916);
and U4421 (N_4421,N_1920,N_381);
or U4422 (N_4422,N_3392,N_3815);
and U4423 (N_4423,N_3982,N_2794);
or U4424 (N_4424,N_2253,N_2583);
or U4425 (N_4425,N_3264,N_1421);
or U4426 (N_4426,N_248,N_2065);
or U4427 (N_4427,N_3,N_1256);
xnor U4428 (N_4428,N_3203,N_49);
or U4429 (N_4429,N_568,N_534);
nor U4430 (N_4430,N_3233,N_3949);
nor U4431 (N_4431,N_1617,N_2302);
nand U4432 (N_4432,N_312,N_1478);
nor U4433 (N_4433,N_1097,N_3358);
and U4434 (N_4434,N_1616,N_1194);
or U4435 (N_4435,N_1875,N_590);
xnor U4436 (N_4436,N_2140,N_2693);
nand U4437 (N_4437,N_3795,N_1227);
and U4438 (N_4438,N_3626,N_13);
or U4439 (N_4439,N_2747,N_3258);
or U4440 (N_4440,N_707,N_2852);
or U4441 (N_4441,N_710,N_1081);
and U4442 (N_4442,N_2977,N_1576);
or U4443 (N_4443,N_3799,N_2604);
xnor U4444 (N_4444,N_2552,N_1317);
nand U4445 (N_4445,N_2268,N_5);
xnor U4446 (N_4446,N_1808,N_2448);
nor U4447 (N_4447,N_2545,N_1100);
xor U4448 (N_4448,N_3492,N_2726);
xor U4449 (N_4449,N_3947,N_795);
nand U4450 (N_4450,N_666,N_1997);
xnor U4451 (N_4451,N_1316,N_3225);
and U4452 (N_4452,N_213,N_3271);
nor U4453 (N_4453,N_2360,N_2763);
nand U4454 (N_4454,N_2888,N_112);
and U4455 (N_4455,N_1289,N_1441);
nor U4456 (N_4456,N_1440,N_3030);
nand U4457 (N_4457,N_1434,N_3431);
or U4458 (N_4458,N_252,N_52);
or U4459 (N_4459,N_591,N_2547);
and U4460 (N_4460,N_1510,N_161);
nor U4461 (N_4461,N_3813,N_3014);
xor U4462 (N_4462,N_87,N_2803);
and U4463 (N_4463,N_1469,N_2071);
or U4464 (N_4464,N_2651,N_1241);
or U4465 (N_4465,N_571,N_1406);
nand U4466 (N_4466,N_3685,N_1009);
nand U4467 (N_4467,N_2757,N_399);
or U4468 (N_4468,N_3398,N_2709);
or U4469 (N_4469,N_3051,N_1318);
or U4470 (N_4470,N_352,N_2854);
and U4471 (N_4471,N_2862,N_741);
nand U4472 (N_4472,N_1351,N_1429);
nor U4473 (N_4473,N_2714,N_1255);
nand U4474 (N_4474,N_3360,N_96);
and U4475 (N_4475,N_3550,N_3643);
and U4476 (N_4476,N_3656,N_1409);
xnor U4477 (N_4477,N_1601,N_3067);
xnor U4478 (N_4478,N_1784,N_1608);
or U4479 (N_4479,N_3127,N_799);
and U4480 (N_4480,N_307,N_2890);
nor U4481 (N_4481,N_2808,N_2599);
or U4482 (N_4482,N_1536,N_772);
xnor U4483 (N_4483,N_1643,N_285);
nand U4484 (N_4484,N_3748,N_1339);
nor U4485 (N_4485,N_1174,N_140);
nand U4486 (N_4486,N_2434,N_2771);
or U4487 (N_4487,N_1183,N_3865);
or U4488 (N_4488,N_2639,N_2618);
nand U4489 (N_4489,N_686,N_3056);
xor U4490 (N_4490,N_2725,N_1712);
nor U4491 (N_4491,N_1470,N_813);
and U4492 (N_4492,N_1861,N_2453);
xor U4493 (N_4493,N_3286,N_3839);
nor U4494 (N_4494,N_2030,N_3953);
nand U4495 (N_4495,N_565,N_3195);
and U4496 (N_4496,N_3848,N_3628);
xor U4497 (N_4497,N_1093,N_3599);
xnor U4498 (N_4498,N_567,N_2157);
nand U4499 (N_4499,N_186,N_2006);
nor U4500 (N_4500,N_1755,N_435);
or U4501 (N_4501,N_3665,N_1902);
or U4502 (N_4502,N_1700,N_702);
nor U4503 (N_4503,N_1267,N_2696);
nand U4504 (N_4504,N_241,N_3806);
nor U4505 (N_4505,N_3505,N_3911);
nand U4506 (N_4506,N_833,N_1435);
and U4507 (N_4507,N_3549,N_3093);
xnor U4508 (N_4508,N_1589,N_2203);
nand U4509 (N_4509,N_2190,N_2525);
xor U4510 (N_4510,N_960,N_1879);
or U4511 (N_4511,N_917,N_2537);
nand U4512 (N_4512,N_3414,N_2913);
xnor U4513 (N_4513,N_308,N_1821);
or U4514 (N_4514,N_2603,N_235);
nand U4515 (N_4515,N_2048,N_2867);
nand U4516 (N_4516,N_2516,N_2788);
nand U4517 (N_4517,N_1714,N_1590);
and U4518 (N_4518,N_612,N_1238);
and U4519 (N_4519,N_2485,N_3722);
or U4520 (N_4520,N_1132,N_914);
or U4521 (N_4521,N_3407,N_2860);
xnor U4522 (N_4522,N_1352,N_2729);
or U4523 (N_4523,N_3415,N_2713);
xor U4524 (N_4524,N_547,N_1006);
nand U4525 (N_4525,N_3828,N_407);
or U4526 (N_4526,N_1505,N_3684);
nor U4527 (N_4527,N_3496,N_374);
or U4528 (N_4528,N_1583,N_1184);
nand U4529 (N_4529,N_3540,N_1032);
or U4530 (N_4530,N_916,N_375);
nor U4531 (N_4531,N_480,N_3304);
xor U4532 (N_4532,N_3714,N_2596);
and U4533 (N_4533,N_1104,N_1245);
nand U4534 (N_4534,N_1830,N_3477);
nand U4535 (N_4535,N_2536,N_545);
nor U4536 (N_4536,N_464,N_1693);
nand U4537 (N_4537,N_2909,N_727);
nand U4538 (N_4538,N_669,N_3871);
nand U4539 (N_4539,N_3859,N_1110);
nor U4540 (N_4540,N_3529,N_2722);
xor U4541 (N_4541,N_2690,N_1726);
or U4542 (N_4542,N_3238,N_3932);
and U4543 (N_4543,N_124,N_3670);
xnor U4544 (N_4544,N_1553,N_431);
or U4545 (N_4545,N_100,N_2588);
nand U4546 (N_4546,N_587,N_2038);
nand U4547 (N_4547,N_3689,N_3767);
or U4548 (N_4548,N_1304,N_3733);
and U4549 (N_4549,N_2175,N_1944);
xnor U4550 (N_4550,N_3792,N_1775);
nor U4551 (N_4551,N_2571,N_278);
nand U4552 (N_4552,N_954,N_2096);
and U4553 (N_4553,N_1232,N_3338);
xor U4554 (N_4554,N_2685,N_2422);
nor U4555 (N_4555,N_180,N_1091);
and U4556 (N_4556,N_461,N_3602);
xnor U4557 (N_4557,N_3291,N_2901);
nor U4558 (N_4558,N_1407,N_3786);
and U4559 (N_4559,N_2720,N_1891);
or U4560 (N_4560,N_2645,N_251);
or U4561 (N_4561,N_1957,N_2988);
xor U4562 (N_4562,N_2082,N_613);
nand U4563 (N_4563,N_3176,N_3948);
or U4564 (N_4564,N_2809,N_3544);
or U4565 (N_4565,N_3691,N_2465);
nor U4566 (N_4566,N_3681,N_2831);
nor U4567 (N_4567,N_929,N_3768);
nor U4568 (N_4568,N_3457,N_3045);
or U4569 (N_4569,N_2441,N_2800);
nor U4570 (N_4570,N_2476,N_2367);
nand U4571 (N_4571,N_2879,N_97);
xnor U4572 (N_4572,N_300,N_3596);
nor U4573 (N_4573,N_3519,N_466);
nor U4574 (N_4574,N_452,N_1237);
and U4575 (N_4575,N_3087,N_2398);
nor U4576 (N_4576,N_871,N_2281);
nand U4577 (N_4577,N_2118,N_717);
and U4578 (N_4578,N_314,N_2625);
xnor U4579 (N_4579,N_3814,N_585);
or U4580 (N_4580,N_3003,N_1363);
xnor U4581 (N_4581,N_1683,N_703);
and U4582 (N_4582,N_2158,N_2263);
xor U4583 (N_4583,N_1082,N_774);
or U4584 (N_4584,N_2044,N_390);
and U4585 (N_4585,N_3060,N_2847);
and U4586 (N_4586,N_1106,N_3117);
nor U4587 (N_4587,N_2020,N_631);
xor U4588 (N_4588,N_3459,N_1005);
and U4589 (N_4589,N_324,N_2098);
or U4590 (N_4590,N_3619,N_389);
nand U4591 (N_4591,N_3525,N_47);
nor U4592 (N_4592,N_2791,N_1899);
nor U4593 (N_4593,N_2629,N_2256);
and U4594 (N_4594,N_2743,N_2403);
xor U4595 (N_4595,N_1765,N_269);
nand U4596 (N_4596,N_219,N_1489);
xnor U4597 (N_4597,N_2228,N_532);
nor U4598 (N_4598,N_2100,N_767);
and U4599 (N_4599,N_2463,N_106);
or U4600 (N_4600,N_3687,N_2744);
and U4601 (N_4601,N_1783,N_2326);
nand U4602 (N_4602,N_556,N_1016);
or U4603 (N_4603,N_2937,N_45);
nor U4604 (N_4604,N_3512,N_800);
xor U4605 (N_4605,N_1667,N_3523);
nand U4606 (N_4606,N_2849,N_1155);
or U4607 (N_4607,N_3136,N_3642);
xnor U4608 (N_4608,N_240,N_3104);
nor U4609 (N_4609,N_3410,N_1139);
xnor U4610 (N_4610,N_2085,N_518);
xor U4611 (N_4611,N_1308,N_1886);
or U4612 (N_4612,N_50,N_1819);
nand U4613 (N_4613,N_3052,N_2074);
nor U4614 (N_4614,N_1170,N_3140);
nand U4615 (N_4615,N_1264,N_1114);
nand U4616 (N_4616,N_383,N_836);
and U4617 (N_4617,N_3241,N_1002);
xnor U4618 (N_4618,N_580,N_663);
xor U4619 (N_4619,N_2679,N_450);
nand U4620 (N_4620,N_747,N_3625);
or U4621 (N_4621,N_3343,N_1791);
nand U4622 (N_4622,N_2464,N_336);
or U4623 (N_4623,N_915,N_3475);
nand U4624 (N_4624,N_1382,N_658);
and U4625 (N_4625,N_1922,N_3840);
or U4626 (N_4626,N_2715,N_1506);
and U4627 (N_4627,N_3536,N_1622);
nor U4628 (N_4628,N_3832,N_3116);
and U4629 (N_4629,N_2733,N_712);
nor U4630 (N_4630,N_259,N_2451);
nand U4631 (N_4631,N_2295,N_2577);
and U4632 (N_4632,N_2475,N_360);
and U4633 (N_4633,N_3311,N_2447);
nor U4634 (N_4634,N_3564,N_3135);
or U4635 (N_4635,N_2257,N_384);
xnor U4636 (N_4636,N_3718,N_3929);
nor U4637 (N_4637,N_2185,N_3278);
xnor U4638 (N_4638,N_1619,N_2939);
and U4639 (N_4639,N_1105,N_2214);
or U4640 (N_4640,N_1665,N_816);
nor U4641 (N_4641,N_679,N_2294);
nor U4642 (N_4642,N_2311,N_2279);
nor U4643 (N_4643,N_3297,N_2298);
or U4644 (N_4644,N_1154,N_1722);
xnor U4645 (N_4645,N_1564,N_3196);
xnor U4646 (N_4646,N_3977,N_3376);
nand U4647 (N_4647,N_2469,N_1586);
or U4648 (N_4648,N_212,N_2745);
nor U4649 (N_4649,N_3447,N_623);
and U4650 (N_4650,N_1728,N_447);
and U4651 (N_4651,N_1028,N_1656);
xnor U4652 (N_4652,N_624,N_3844);
xor U4653 (N_4653,N_1720,N_3772);
and U4654 (N_4654,N_1465,N_3462);
nand U4655 (N_4655,N_1833,N_3027);
nand U4656 (N_4656,N_730,N_3930);
nor U4657 (N_4657,N_3900,N_1732);
nor U4658 (N_4658,N_2777,N_1198);
nor U4659 (N_4659,N_634,N_2099);
nand U4660 (N_4660,N_3296,N_1628);
xor U4661 (N_4661,N_3197,N_1528);
or U4662 (N_4662,N_3883,N_3941);
xor U4663 (N_4663,N_3673,N_2661);
or U4664 (N_4664,N_1479,N_1648);
or U4665 (N_4665,N_116,N_1305);
and U4666 (N_4666,N_159,N_3908);
and U4667 (N_4667,N_3029,N_3439);
nor U4668 (N_4668,N_428,N_778);
nor U4669 (N_4669,N_3059,N_2492);
nand U4670 (N_4670,N_3648,N_423);
nor U4671 (N_4671,N_1216,N_1853);
xnor U4672 (N_4672,N_1562,N_549);
nor U4673 (N_4673,N_1457,N_2608);
and U4674 (N_4674,N_35,N_1481);
and U4675 (N_4675,N_943,N_2305);
or U4676 (N_4676,N_320,N_848);
or U4677 (N_4677,N_2292,N_135);
nor U4678 (N_4678,N_1531,N_1278);
nand U4679 (N_4679,N_1017,N_3926);
nor U4680 (N_4680,N_2799,N_3276);
nor U4681 (N_4681,N_1935,N_234);
or U4682 (N_4682,N_3766,N_779);
xnor U4683 (N_4683,N_3825,N_1865);
xnor U4684 (N_4684,N_2177,N_3434);
nor U4685 (N_4685,N_3913,N_1298);
nor U4686 (N_4686,N_864,N_454);
nand U4687 (N_4687,N_2557,N_3015);
and U4688 (N_4688,N_3406,N_2775);
xor U4689 (N_4689,N_1988,N_2553);
and U4690 (N_4690,N_3762,N_2086);
and U4691 (N_4691,N_470,N_992);
xor U4692 (N_4692,N_2751,N_2786);
nand U4693 (N_4693,N_83,N_230);
and U4694 (N_4694,N_3621,N_922);
nor U4695 (N_4695,N_3937,N_2621);
nand U4696 (N_4696,N_1394,N_3046);
xnor U4697 (N_4697,N_319,N_3429);
nor U4698 (N_4698,N_654,N_1953);
or U4699 (N_4699,N_577,N_2683);
nor U4700 (N_4700,N_3605,N_1041);
nand U4701 (N_4701,N_2344,N_2050);
nor U4702 (N_4702,N_2826,N_1334);
nand U4703 (N_4703,N_2147,N_2046);
xnor U4704 (N_4704,N_2163,N_3220);
nor U4705 (N_4705,N_1537,N_2217);
nor U4706 (N_4706,N_701,N_1878);
nand U4707 (N_4707,N_2827,N_2944);
or U4708 (N_4708,N_997,N_620);
or U4709 (N_4709,N_2761,N_1782);
nor U4710 (N_4710,N_3978,N_2225);
and U4711 (N_4711,N_722,N_805);
or U4712 (N_4712,N_3344,N_2443);
or U4713 (N_4713,N_1569,N_146);
xnor U4714 (N_4714,N_2605,N_2778);
nand U4715 (N_4715,N_56,N_63);
or U4716 (N_4716,N_2432,N_1359);
nand U4717 (N_4717,N_3301,N_2019);
and U4718 (N_4718,N_2251,N_1040);
nand U4719 (N_4719,N_2850,N_2205);
nor U4720 (N_4720,N_3193,N_2932);
nor U4721 (N_4721,N_2416,N_956);
nand U4722 (N_4722,N_1065,N_3274);
nand U4723 (N_4723,N_1668,N_2573);
or U4724 (N_4724,N_2865,N_2042);
nor U4725 (N_4725,N_3102,N_1666);
nand U4726 (N_4726,N_2057,N_413);
and U4727 (N_4727,N_1670,N_3365);
or U4728 (N_4728,N_2950,N_1452);
nor U4729 (N_4729,N_1636,N_655);
nand U4730 (N_4730,N_1102,N_1043);
nand U4731 (N_4731,N_1175,N_2133);
and U4732 (N_4732,N_946,N_554);
nand U4733 (N_4733,N_1173,N_2627);
xor U4734 (N_4734,N_3877,N_688);
nor U4735 (N_4735,N_2845,N_3266);
xor U4736 (N_4736,N_1816,N_3713);
nor U4737 (N_4737,N_1492,N_723);
xor U4738 (N_4738,N_3719,N_3237);
or U4739 (N_4739,N_18,N_2882);
or U4740 (N_4740,N_1914,N_2262);
and U4741 (N_4741,N_2721,N_1261);
xnor U4742 (N_4742,N_3034,N_3823);
nor U4743 (N_4743,N_1064,N_249);
xor U4744 (N_4744,N_414,N_786);
or U4745 (N_4745,N_3210,N_789);
nor U4746 (N_4746,N_32,N_2789);
nand U4747 (N_4747,N_1045,N_3672);
nor U4748 (N_4748,N_2334,N_616);
xor U4749 (N_4749,N_2748,N_769);
xnor U4750 (N_4750,N_3310,N_2617);
nand U4751 (N_4751,N_1348,N_1858);
or U4752 (N_4752,N_2870,N_726);
and U4753 (N_4753,N_110,N_506);
or U4754 (N_4754,N_1244,N_1936);
and U4755 (N_4755,N_3472,N_1927);
nand U4756 (N_4756,N_1285,N_2817);
or U4757 (N_4757,N_1260,N_1972);
xor U4758 (N_4758,N_1523,N_878);
or U4759 (N_4759,N_3356,N_1079);
nor U4760 (N_4760,N_3960,N_1172);
nand U4761 (N_4761,N_2580,N_2395);
or U4762 (N_4762,N_3836,N_2754);
or U4763 (N_4763,N_3039,N_2739);
nor U4764 (N_4764,N_1828,N_3962);
nand U4765 (N_4765,N_2047,N_1711);
xnor U4766 (N_4766,N_1376,N_1561);
and U4767 (N_4767,N_2707,N_2004);
xor U4768 (N_4768,N_190,N_3369);
nor U4769 (N_4769,N_3517,N_2468);
xnor U4770 (N_4770,N_3756,N_3318);
and U4771 (N_4771,N_3841,N_157);
and U4772 (N_4772,N_1943,N_2838);
nor U4773 (N_4773,N_1509,N_3055);
nand U4774 (N_4774,N_460,N_1725);
nor U4775 (N_4775,N_1857,N_408);
xnor U4776 (N_4776,N_2986,N_3260);
and U4777 (N_4777,N_117,N_479);
or U4778 (N_4778,N_1814,N_2056);
xnor U4779 (N_4779,N_552,N_2136);
xor U4780 (N_4780,N_1384,N_2011);
nand U4781 (N_4781,N_1734,N_999);
and U4782 (N_4782,N_156,N_1960);
or U4783 (N_4783,N_3445,N_2546);
or U4784 (N_4784,N_3740,N_3566);
or U4785 (N_4785,N_2873,N_3801);
nor U4786 (N_4786,N_2955,N_3340);
nand U4787 (N_4787,N_1574,N_1604);
and U4788 (N_4788,N_1372,N_2015);
xnor U4789 (N_4789,N_1408,N_3155);
nand U4790 (N_4790,N_3915,N_1818);
xor U4791 (N_4791,N_1107,N_2309);
nor U4792 (N_4792,N_783,N_1069);
nand U4793 (N_4793,N_3111,N_1789);
nand U4794 (N_4794,N_1023,N_2942);
and U4795 (N_4795,N_2643,N_1450);
or U4796 (N_4796,N_1634,N_621);
or U4797 (N_4797,N_3273,N_1022);
or U4798 (N_4798,N_3983,N_2619);
nand U4799 (N_4799,N_2924,N_1704);
nand U4800 (N_4800,N_3289,N_849);
or U4801 (N_4801,N_1411,N_174);
nand U4802 (N_4802,N_1086,N_3500);
and U4803 (N_4803,N_863,N_2402);
nor U4804 (N_4804,N_3294,N_1369);
or U4805 (N_4805,N_1101,N_82);
or U4806 (N_4806,N_30,N_3211);
or U4807 (N_4807,N_797,N_23);
nand U4808 (N_4808,N_2980,N_1572);
nand U4809 (N_4809,N_3458,N_104);
nand U4810 (N_4810,N_3555,N_1518);
or U4811 (N_4811,N_1262,N_3263);
nand U4812 (N_4812,N_386,N_3096);
and U4813 (N_4813,N_1598,N_2768);
or U4814 (N_4814,N_1580,N_1547);
and U4815 (N_4815,N_968,N_1946);
nand U4816 (N_4816,N_2660,N_1089);
or U4817 (N_4817,N_3405,N_3194);
nand U4818 (N_4818,N_2699,N_2538);
and U4819 (N_4819,N_2264,N_503);
and U4820 (N_4820,N_3649,N_3620);
and U4821 (N_4821,N_429,N_455);
or U4822 (N_4822,N_3471,N_1292);
nand U4823 (N_4823,N_2591,N_2723);
xnor U4824 (N_4824,N_3058,N_148);
and U4825 (N_4825,N_1025,N_2631);
nor U4826 (N_4826,N_502,N_2209);
and U4827 (N_4827,N_2156,N_1901);
nor U4828 (N_4828,N_510,N_2948);
nand U4829 (N_4829,N_3371,N_2426);
xnor U4830 (N_4830,N_2659,N_873);
nand U4831 (N_4831,N_607,N_1959);
xnor U4832 (N_4832,N_350,N_1799);
xnor U4833 (N_4833,N_829,N_1490);
or U4834 (N_4834,N_665,N_3964);
nand U4835 (N_4835,N_3038,N_73);
nor U4836 (N_4836,N_2990,N_823);
xor U4837 (N_4837,N_1941,N_2128);
nor U4838 (N_4838,N_2756,N_2379);
nor U4839 (N_4839,N_3353,N_442);
nand U4840 (N_4840,N_3910,N_1621);
and U4841 (N_4841,N_3226,N_1892);
xnor U4842 (N_4842,N_3601,N_306);
and U4843 (N_4843,N_2407,N_1269);
nor U4844 (N_4844,N_925,N_218);
nor U4845 (N_4845,N_318,N_3752);
or U4846 (N_4846,N_2823,N_3363);
xnor U4847 (N_4847,N_298,N_1809);
xnor U4848 (N_4848,N_1868,N_2444);
and U4849 (N_4849,N_1169,N_376);
nor U4850 (N_4850,N_1610,N_2910);
and U4851 (N_4851,N_3109,N_3923);
xnor U4852 (N_4852,N_250,N_1176);
or U4853 (N_4853,N_2454,N_2013);
or U4854 (N_4854,N_1247,N_3769);
xnor U4855 (N_4855,N_134,N_3147);
and U4856 (N_4856,N_2151,N_20);
xor U4857 (N_4857,N_1760,N_1118);
nor U4858 (N_4858,N_989,N_1095);
and U4859 (N_4859,N_37,N_2058);
nor U4860 (N_4860,N_1129,N_1315);
or U4861 (N_4861,N_1068,N_837);
xor U4862 (N_4862,N_754,N_2353);
or U4863 (N_4863,N_2061,N_1300);
and U4864 (N_4864,N_2734,N_3667);
nand U4865 (N_4865,N_2563,N_2208);
and U4866 (N_4866,N_656,N_1862);
or U4867 (N_4867,N_1798,N_3528);
nor U4868 (N_4868,N_3584,N_2167);
nor U4869 (N_4869,N_2155,N_3958);
or U4870 (N_4870,N_1099,N_2526);
or U4871 (N_4871,N_847,N_608);
xnor U4872 (N_4872,N_2139,N_2127);
nand U4873 (N_4873,N_3727,N_541);
xnor U4874 (N_4874,N_1820,N_2380);
or U4875 (N_4875,N_790,N_632);
or U4876 (N_4876,N_3397,N_2912);
nor U4877 (N_4877,N_105,N_1480);
and U4878 (N_4878,N_660,N_2200);
or U4879 (N_4879,N_2097,N_3531);
and U4880 (N_4880,N_934,N_1877);
or U4881 (N_4881,N_1504,N_198);
and U4882 (N_4882,N_130,N_3452);
nand U4883 (N_4883,N_3565,N_377);
xnor U4884 (N_4884,N_1314,N_178);
and U4885 (N_4885,N_1425,N_1672);
xnor U4886 (N_4886,N_729,N_3972);
and U4887 (N_4887,N_3856,N_2108);
and U4888 (N_4888,N_1895,N_3372);
xnor U4889 (N_4889,N_3348,N_3368);
and U4890 (N_4890,N_3486,N_2271);
nand U4891 (N_4891,N_1131,N_1748);
nand U4892 (N_4892,N_3380,N_2945);
nor U4893 (N_4893,N_1430,N_3901);
or U4894 (N_4894,N_1641,N_3838);
nand U4895 (N_4895,N_436,N_378);
xnor U4896 (N_4896,N_749,N_2418);
xor U4897 (N_4897,N_3257,N_292);
xnor U4898 (N_4898,N_3146,N_3980);
xor U4899 (N_4899,N_1463,N_295);
xnor U4900 (N_4900,N_3578,N_276);
or U4901 (N_4901,N_1148,N_3568);
and U4902 (N_4902,N_226,N_2357);
xnor U4903 (N_4903,N_1591,N_1851);
or U4904 (N_4904,N_1287,N_2063);
nor U4905 (N_4905,N_935,N_1924);
nor U4906 (N_4906,N_526,N_1270);
xnor U4907 (N_4907,N_1723,N_919);
nor U4908 (N_4908,N_2535,N_3933);
xor U4909 (N_4909,N_101,N_28);
nor U4910 (N_4910,N_283,N_3760);
or U4911 (N_4911,N_1541,N_2837);
nand U4912 (N_4912,N_2881,N_2389);
xnor U4913 (N_4913,N_2349,N_2413);
or U4914 (N_4914,N_1248,N_2480);
nand U4915 (N_4915,N_1741,N_294);
or U4916 (N_4916,N_901,N_3616);
and U4917 (N_4917,N_1934,N_1433);
and U4918 (N_4918,N_3623,N_2356);
xnor U4919 (N_4919,N_3412,N_1973);
nor U4920 (N_4920,N_3631,N_501);
and U4921 (N_4921,N_2764,N_182);
or U4922 (N_4922,N_42,N_2037);
and U4923 (N_4923,N_2088,N_1849);
nor U4924 (N_4924,N_911,N_538);
and U4925 (N_4925,N_611,N_1888);
nor U4926 (N_4926,N_2880,N_2501);
nor U4927 (N_4927,N_1746,N_2406);
or U4928 (N_4928,N_2286,N_1827);
or U4929 (N_4929,N_302,N_888);
nand U4930 (N_4930,N_1905,N_3202);
or U4931 (N_4931,N_1475,N_1221);
and U4932 (N_4932,N_1044,N_277);
nor U4933 (N_4933,N_3390,N_3235);
or U4934 (N_4934,N_1841,N_1415);
xnor U4935 (N_4935,N_3992,N_1488);
xor U4936 (N_4936,N_595,N_1013);
nand U4937 (N_4937,N_483,N_1903);
nor U4938 (N_4938,N_2731,N_2960);
nor U4939 (N_4939,N_347,N_1716);
and U4940 (N_4940,N_3024,N_422);
xor U4941 (N_4941,N_2851,N_2566);
xor U4942 (N_4942,N_3323,N_1907);
xor U4943 (N_4943,N_2844,N_2222);
or U4944 (N_4944,N_3053,N_1952);
nor U4945 (N_4945,N_1165,N_3598);
nor U4946 (N_4946,N_1516,N_1297);
xor U4947 (N_4947,N_2124,N_3918);
nand U4948 (N_4948,N_2165,N_2408);
nor U4949 (N_4949,N_16,N_1484);
or U4950 (N_4950,N_2821,N_1570);
nor U4951 (N_4951,N_2512,N_1035);
nor U4952 (N_4952,N_2308,N_2484);
or U4953 (N_4953,N_3987,N_1597);
nor U4954 (N_4954,N_3732,N_340);
nand U4955 (N_4955,N_2642,N_3473);
nand U4956 (N_4956,N_3637,N_370);
nor U4957 (N_4957,N_3515,N_2212);
and U4958 (N_4958,N_1196,N_3697);
nand U4959 (N_4959,N_739,N_3247);
or U4960 (N_4960,N_3671,N_2499);
nor U4961 (N_4961,N_3252,N_1431);
xor U4962 (N_4962,N_2146,N_3254);
or U4963 (N_4963,N_891,N_633);
and U4964 (N_4964,N_391,N_1773);
or U4965 (N_4965,N_2676,N_279);
nand U4966 (N_4966,N_93,N_2440);
nand U4967 (N_4967,N_1918,N_2669);
nor U4968 (N_4968,N_2260,N_3530);
nor U4969 (N_4969,N_433,N_275);
or U4970 (N_4970,N_3316,N_2646);
or U4971 (N_4971,N_1404,N_1717);
nor U4972 (N_4972,N_2564,N_3742);
or U4973 (N_4973,N_1778,N_1462);
or U4974 (N_4974,N_855,N_2760);
nor U4975 (N_4975,N_2255,N_993);
and U4976 (N_4976,N_64,N_2587);
and U4977 (N_4977,N_2962,N_3057);
or U4978 (N_4978,N_3805,N_618);
nor U4979 (N_4979,N_3589,N_2872);
or U4980 (N_4980,N_2010,N_2307);
or U4981 (N_4981,N_609,N_1501);
xnor U4982 (N_4982,N_194,N_2724);
nand U4983 (N_4983,N_3809,N_15);
and U4984 (N_4984,N_3277,N_1037);
xnor U4985 (N_4985,N_2700,N_3474);
and U4986 (N_4986,N_3654,N_742);
nand U4987 (N_4987,N_3993,N_3943);
xnor U4988 (N_4988,N_3506,N_2003);
or U4989 (N_4989,N_1268,N_2363);
or U4990 (N_4990,N_2031,N_1223);
nand U4991 (N_4991,N_3230,N_625);
and U4992 (N_4992,N_3686,N_2104);
and U4993 (N_4993,N_1401,N_424);
nand U4994 (N_4994,N_3213,N_2755);
nand U4995 (N_4995,N_3676,N_3776);
and U4996 (N_4996,N_1367,N_3354);
xor U4997 (N_4997,N_2769,N_1979);
xor U4998 (N_4998,N_53,N_675);
and U4999 (N_4999,N_88,N_3891);
nor U5000 (N_5000,N_1271,N_432);
xnor U5001 (N_5001,N_98,N_3299);
and U5002 (N_5002,N_392,N_1239);
nand U5003 (N_5003,N_546,N_1669);
xnor U5004 (N_5004,N_281,N_1103);
nand U5005 (N_5005,N_574,N_200);
xnor U5006 (N_5006,N_2911,N_2244);
nor U5007 (N_5007,N_1398,N_1731);
xnor U5008 (N_5008,N_1189,N_3101);
xor U5009 (N_5009,N_3696,N_948);
nor U5010 (N_5010,N_6,N_976);
nor U5011 (N_5011,N_3543,N_1163);
xor U5012 (N_5012,N_563,N_3313);
or U5013 (N_5013,N_3180,N_603);
nor U5014 (N_5014,N_2362,N_2510);
xor U5015 (N_5015,N_681,N_1548);
or U5016 (N_5016,N_3190,N_978);
nand U5017 (N_5017,N_1312,N_2179);
and U5018 (N_5018,N_1294,N_3850);
xor U5019 (N_5019,N_3853,N_165);
nor U5020 (N_5020,N_1615,N_238);
or U5021 (N_5021,N_441,N_3063);
xor U5022 (N_5022,N_1555,N_3562);
or U5023 (N_5023,N_1801,N_1365);
or U5024 (N_5024,N_3875,N_2069);
nor U5025 (N_5025,N_3171,N_653);
or U5026 (N_5026,N_3609,N_1958);
or U5027 (N_5027,N_3855,N_488);
and U5028 (N_5028,N_2312,N_143);
nor U5029 (N_5029,N_3440,N_1832);
nor U5030 (N_5030,N_918,N_1768);
nor U5031 (N_5031,N_1839,N_1626);
nand U5032 (N_5032,N_41,N_2012);
or U5033 (N_5033,N_2273,N_777);
or U5034 (N_5034,N_3563,N_2076);
nor U5035 (N_5035,N_1486,N_311);
nand U5036 (N_5036,N_3062,N_1998);
or U5037 (N_5037,N_1800,N_3444);
nand U5038 (N_5038,N_3357,N_3399);
or U5039 (N_5039,N_2543,N_1950);
or U5040 (N_5040,N_962,N_288);
or U5041 (N_5041,N_3669,N_1249);
nand U5042 (N_5042,N_659,N_1217);
or U5043 (N_5043,N_1985,N_3085);
xor U5044 (N_5044,N_1387,N_419);
xor U5045 (N_5045,N_3113,N_55);
or U5046 (N_5046,N_2369,N_890);
nand U5047 (N_5047,N_979,N_758);
and U5048 (N_5048,N_3006,N_2918);
or U5049 (N_5049,N_2376,N_1999);
or U5050 (N_5050,N_1817,N_341);
and U5051 (N_5051,N_2927,N_2123);
nand U5052 (N_5052,N_2023,N_958);
xor U5053 (N_5053,N_600,N_3307);
and U5054 (N_5054,N_2248,N_1389);
xor U5055 (N_5055,N_1061,N_81);
nor U5056 (N_5056,N_2753,N_902);
nand U5057 (N_5057,N_490,N_2568);
xor U5058 (N_5058,N_3816,N_1345);
xnor U5059 (N_5059,N_629,N_2300);
nand U5060 (N_5060,N_245,N_2301);
xor U5061 (N_5061,N_139,N_371);
or U5062 (N_5062,N_2199,N_236);
and U5063 (N_5063,N_1051,N_2793);
xor U5064 (N_5064,N_1439,N_851);
and U5065 (N_5065,N_2866,N_2491);
nand U5066 (N_5066,N_3975,N_2956);
and U5067 (N_5067,N_3106,N_3455);
nand U5068 (N_5068,N_1843,N_1592);
nand U5069 (N_5069,N_1823,N_2670);
nand U5070 (N_5070,N_2996,N_207);
and U5071 (N_5071,N_3624,N_3524);
xnor U5072 (N_5072,N_299,N_401);
or U5073 (N_5073,N_2897,N_2045);
or U5074 (N_5074,N_2027,N_1325);
xor U5075 (N_5075,N_1864,N_3336);
nor U5076 (N_5076,N_822,N_3804);
nand U5077 (N_5077,N_1707,N_1558);
nand U5078 (N_5078,N_2073,N_3761);
and U5079 (N_5079,N_1254,N_977);
nand U5080 (N_5080,N_1293,N_3759);
xnor U5081 (N_5081,N_2653,N_268);
or U5082 (N_5082,N_3864,N_2220);
nor U5083 (N_5083,N_2970,N_2567);
nor U5084 (N_5084,N_3465,N_1162);
or U5085 (N_5085,N_2736,N_3091);
nand U5086 (N_5086,N_735,N_2425);
nand U5087 (N_5087,N_2161,N_1358);
and U5088 (N_5088,N_1738,N_332);
nand U5089 (N_5089,N_3121,N_2732);
nand U5090 (N_5090,N_233,N_2384);
nor U5091 (N_5091,N_2423,N_2657);
nor U5092 (N_5092,N_642,N_983);
or U5093 (N_5093,N_1680,N_2417);
and U5094 (N_5094,N_1161,N_866);
or U5095 (N_5095,N_2481,N_147);
nor U5096 (N_5096,N_1357,N_2885);
nor U5097 (N_5097,N_2833,N_481);
xnor U5098 (N_5098,N_2610,N_3229);
or U5099 (N_5099,N_3388,N_266);
nor U5100 (N_5100,N_2397,N_2348);
and U5101 (N_5101,N_346,N_1646);
nand U5102 (N_5102,N_3845,N_3973);
nor U5103 (N_5103,N_2899,N_1756);
nand U5104 (N_5104,N_744,N_3857);
nor U5105 (N_5105,N_1870,N_1228);
and U5106 (N_5106,N_103,N_1191);
nand U5107 (N_5107,N_3427,N_2280);
nor U5108 (N_5108,N_910,N_2781);
xnor U5109 (N_5109,N_3251,N_3567);
or U5110 (N_5110,N_896,N_3393);
and U5111 (N_5111,N_491,N_947);
nand U5112 (N_5112,N_1412,N_793);
nor U5113 (N_5113,N_3200,N_1989);
nor U5114 (N_5114,N_3998,N_1181);
nor U5115 (N_5115,N_2055,N_3256);
or U5116 (N_5116,N_1525,N_2316);
nand U5117 (N_5117,N_1606,N_1658);
nand U5118 (N_5118,N_457,N_2409);
nand U5119 (N_5119,N_2022,N_909);
or U5120 (N_5120,N_1377,N_3377);
nor U5121 (N_5121,N_2868,N_1251);
and U5122 (N_5122,N_1585,N_1507);
or U5123 (N_5123,N_1893,N_3272);
and U5124 (N_5124,N_1096,N_3309);
or U5125 (N_5125,N_500,N_877);
nor U5126 (N_5126,N_1395,N_1473);
or U5127 (N_5127,N_3640,N_2446);
and U5128 (N_5128,N_963,N_2717);
xnor U5129 (N_5129,N_1386,N_3032);
or U5130 (N_5130,N_3818,N_1014);
nor U5131 (N_5131,N_2293,N_3575);
and U5132 (N_5132,N_2762,N_3907);
xor U5133 (N_5133,N_664,N_3675);
xor U5134 (N_5134,N_630,N_1214);
or U5135 (N_5135,N_1046,N_1894);
and U5136 (N_5136,N_1295,N_1145);
nand U5137 (N_5137,N_3033,N_1898);
and U5138 (N_5138,N_1860,N_1442);
or U5139 (N_5139,N_1649,N_192);
nand U5140 (N_5140,N_2839,N_835);
and U5141 (N_5141,N_224,N_193);
xnor U5142 (N_5142,N_3968,N_263);
or U5143 (N_5143,N_1687,N_142);
nor U5144 (N_5144,N_2524,N_544);
nor U5145 (N_5145,N_2034,N_3367);
xnor U5146 (N_5146,N_2105,N_542);
and U5147 (N_5147,N_1593,N_1874);
or U5148 (N_5148,N_2974,N_3858);
nand U5149 (N_5149,N_1413,N_1128);
xnor U5150 (N_5150,N_67,N_141);
xnor U5151 (N_5151,N_3021,N_3778);
and U5152 (N_5152,N_2289,N_3285);
nor U5153 (N_5153,N_2664,N_560);
and U5154 (N_5154,N_3702,N_1805);
nor U5155 (N_5155,N_1887,N_3651);
xnor U5156 (N_5156,N_3099,N_1445);
and U5157 (N_5157,N_1259,N_1059);
nor U5158 (N_5158,N_766,N_3011);
nor U5159 (N_5159,N_1180,N_2231);
or U5160 (N_5160,N_801,N_892);
and U5161 (N_5161,N_2606,N_1520);
xor U5162 (N_5162,N_1049,N_2894);
and U5163 (N_5163,N_2698,N_315);
nor U5164 (N_5164,N_3078,N_475);
nor U5165 (N_5165,N_133,N_2072);
xor U5166 (N_5166,N_2997,N_3364);
xor U5167 (N_5167,N_271,N_2324);
nor U5168 (N_5168,N_2153,N_3999);
or U5169 (N_5169,N_3699,N_635);
or U5170 (N_5170,N_188,N_1826);
nor U5171 (N_5171,N_2575,N_3709);
xnor U5172 (N_5172,N_345,N_2656);
nand U5173 (N_5173,N_3302,N_406);
and U5174 (N_5174,N_2742,N_3784);
nor U5175 (N_5175,N_1150,N_843);
and U5176 (N_5176,N_3622,N_1152);
nand U5177 (N_5177,N_2049,N_3881);
or U5178 (N_5178,N_921,N_2782);
and U5179 (N_5179,N_90,N_3284);
xor U5180 (N_5180,N_409,N_2985);
nor U5181 (N_5181,N_2018,N_684);
nand U5182 (N_5182,N_3337,N_3955);
and U5183 (N_5183,N_463,N_418);
or U5184 (N_5184,N_2925,N_3110);
nand U5185 (N_5185,N_839,N_379);
nor U5186 (N_5186,N_2884,N_3737);
xor U5187 (N_5187,N_3914,N_3547);
nand U5188 (N_5188,N_3614,N_1385);
xor U5189 (N_5189,N_2318,N_671);
or U5190 (N_5190,N_3928,N_3826);
nand U5191 (N_5191,N_2517,N_1701);
or U5192 (N_5192,N_152,N_2043);
xnor U5193 (N_5193,N_832,N_2667);
nor U5194 (N_5194,N_677,N_1);
or U5195 (N_5195,N_2207,N_1432);
or U5196 (N_5196,N_325,N_2554);
and U5197 (N_5197,N_637,N_196);
or U5198 (N_5198,N_1631,N_3842);
or U5199 (N_5199,N_920,N_3851);
or U5200 (N_5200,N_2333,N_2101);
and U5201 (N_5201,N_2674,N_3746);
xor U5202 (N_5202,N_903,N_693);
xor U5203 (N_5203,N_3419,N_2148);
and U5204 (N_5204,N_806,N_2581);
nand U5205 (N_5205,N_3904,N_1422);
or U5206 (N_5206,N_1420,N_3944);
nor U5207 (N_5207,N_711,N_3979);
xor U5208 (N_5208,N_2987,N_559);
and U5209 (N_5209,N_51,N_1911);
nand U5210 (N_5210,N_738,N_1942);
nor U5211 (N_5211,N_3834,N_714);
nor U5212 (N_5212,N_696,N_825);
or U5213 (N_5213,N_1337,N_1885);
and U5214 (N_5214,N_1710,N_86);
and U5215 (N_5215,N_2392,N_1378);
or U5216 (N_5216,N_1209,N_3217);
xnor U5217 (N_5217,N_3775,N_2365);
nor U5218 (N_5218,N_1499,N_1513);
xnor U5219 (N_5219,N_3868,N_1010);
nand U5220 (N_5220,N_2953,N_2374);
or U5221 (N_5221,N_1762,N_1158);
and U5222 (N_5222,N_3435,N_1074);
or U5223 (N_5223,N_3028,N_321);
or U5224 (N_5224,N_2673,N_3245);
and U5225 (N_5225,N_3729,N_3724);
xor U5226 (N_5226,N_1029,N_708);
nor U5227 (N_5227,N_137,N_959);
and U5228 (N_5228,N_2531,N_3438);
nand U5229 (N_5229,N_3869,N_3731);
xnor U5230 (N_5230,N_1355,N_220);
nor U5231 (N_5231,N_2780,N_2783);
nand U5232 (N_5232,N_3969,N_2983);
and U5233 (N_5233,N_2276,N_906);
xnor U5234 (N_5234,N_2246,N_2522);
or U5235 (N_5235,N_3098,N_3780);
nand U5236 (N_5236,N_1419,N_2064);
and U5237 (N_5237,N_2283,N_1410);
nand U5238 (N_5238,N_2515,N_1056);
xnor U5239 (N_5239,N_3209,N_2922);
nand U5240 (N_5240,N_297,N_827);
or U5241 (N_5241,N_2919,N_3054);
nor U5242 (N_5242,N_2805,N_564);
and U5243 (N_5243,N_2196,N_2162);
xnor U5244 (N_5244,N_2215,N_4);
or U5245 (N_5245,N_3070,N_3378);
and U5246 (N_5246,N_3249,N_3680);
nand U5247 (N_5247,N_3553,N_3847);
xor U5248 (N_5248,N_2091,N_3583);
nor U5249 (N_5249,N_3532,N_2915);
and U5250 (N_5250,N_1600,N_3080);
xor U5251 (N_5251,N_1675,N_697);
and U5252 (N_5252,N_1691,N_857);
or U5253 (N_5253,N_1361,N_2466);
xnor U5254 (N_5254,N_3738,N_1112);
nor U5255 (N_5255,N_1080,N_2371);
xnor U5256 (N_5256,N_2001,N_706);
nand U5257 (N_5257,N_1328,N_1301);
xnor U5258 (N_5258,N_3068,N_2419);
nor U5259 (N_5259,N_1266,N_1047);
nand U5260 (N_5260,N_3144,N_627);
or U5261 (N_5261,N_421,N_1193);
nand U5262 (N_5262,N_1482,N_3122);
nor U5263 (N_5263,N_2275,N_1157);
and U5264 (N_5264,N_3158,N_304);
nor U5265 (N_5265,N_1724,N_3558);
nor U5266 (N_5266,N_1976,N_2174);
nand U5267 (N_5267,N_214,N_39);
nor U5268 (N_5268,N_2706,N_1984);
nand U5269 (N_5269,N_2036,N_2479);
nor U5270 (N_5270,N_924,N_810);
nand U5271 (N_5271,N_3322,N_316);
nor U5272 (N_5272,N_27,N_957);
or U5273 (N_5273,N_961,N_3790);
nor U5274 (N_5274,N_3636,N_3996);
or U5275 (N_5275,N_594,N_1203);
nand U5276 (N_5276,N_971,N_1671);
nor U5277 (N_5277,N_581,N_217);
nor U5278 (N_5278,N_1050,N_3261);
xor U5279 (N_5279,N_394,N_819);
nand U5280 (N_5280,N_1472,N_602);
and U5281 (N_5281,N_169,N_3692);
or U5282 (N_5282,N_1273,N_3205);
nand U5283 (N_5283,N_2306,N_2445);
or U5284 (N_5284,N_824,N_2508);
nor U5285 (N_5285,N_3269,N_397);
nand U5286 (N_5286,N_1688,N_1965);
xor U5287 (N_5287,N_26,N_2166);
or U5288 (N_5288,N_944,N_3861);
nor U5289 (N_5289,N_1845,N_3441);
xnor U5290 (N_5290,N_2740,N_2787);
nor U5291 (N_5291,N_2790,N_3595);
nand U5292 (N_5292,N_3739,N_2662);
and U5293 (N_5293,N_420,N_2327);
xor U5294 (N_5294,N_1567,N_638);
or U5295 (N_5295,N_2556,N_2160);
nor U5296 (N_5296,N_2130,N_2759);
or U5297 (N_5297,N_2801,N_3270);
xnor U5298 (N_5298,N_3695,N_3349);
or U5299 (N_5299,N_1967,N_1697);
xor U5300 (N_5300,N_205,N_2337);
or U5301 (N_5301,N_1695,N_1906);
and U5302 (N_5302,N_3721,N_3416);
and U5303 (N_5303,N_254,N_1896);
nor U5304 (N_5304,N_1063,N_2551);
or U5305 (N_5305,N_1556,N_3049);
xnor U5306 (N_5306,N_2498,N_57);
and U5307 (N_5307,N_1682,N_183);
and U5308 (N_5308,N_1544,N_1142);
xor U5309 (N_5309,N_3066,N_2504);
xor U5310 (N_5310,N_1364,N_2579);
and U5311 (N_5311,N_1344,N_3588);
and U5312 (N_5312,N_3341,N_645);
nand U5313 (N_5313,N_3546,N_3295);
nand U5314 (N_5314,N_1846,N_2682);
and U5315 (N_5315,N_2917,N_3280);
xor U5316 (N_5316,N_3559,N_265);
and U5317 (N_5317,N_530,N_2957);
xnor U5318 (N_5318,N_3331,N_1933);
and U5319 (N_5319,N_2259,N_781);
nand U5320 (N_5320,N_326,N_2000);
xor U5321 (N_5321,N_1908,N_2094);
or U5322 (N_5322,N_3417,N_1373);
nor U5323 (N_5323,N_3788,N_3409);
and U5324 (N_5324,N_715,N_1077);
nor U5325 (N_5325,N_3966,N_3905);
and U5326 (N_5326,N_1769,N_716);
and U5327 (N_5327,N_3115,N_31);
nor U5328 (N_5328,N_2021,N_1639);
and U5329 (N_5329,N_2858,N_3069);
or U5330 (N_5330,N_1185,N_1975);
nor U5331 (N_5331,N_358,N_3151);
nor U5332 (N_5332,N_1326,N_2449);
or U5333 (N_5333,N_3509,N_3829);
xor U5334 (N_5334,N_3298,N_1296);
nand U5335 (N_5335,N_2026,N_1179);
nand U5336 (N_5336,N_517,N_1151);
or U5337 (N_5337,N_689,N_272);
or U5338 (N_5338,N_3537,N_737);
xor U5339 (N_5339,N_842,N_239);
nor U5340 (N_5340,N_3287,N_662);
or U5341 (N_5341,N_1038,N_898);
and U5342 (N_5342,N_927,N_651);
or U5343 (N_5343,N_2878,N_2644);
and U5344 (N_5344,N_2437,N_2795);
and U5345 (N_5345,N_3047,N_3974);
nand U5346 (N_5346,N_509,N_3036);
nor U5347 (N_5347,N_1546,N_640);
and U5348 (N_5348,N_3787,N_2035);
nor U5349 (N_5349,N_1379,N_709);
nor U5350 (N_5350,N_1011,N_3502);
or U5351 (N_5351,N_482,N_524);
xor U5352 (N_5352,N_553,N_3490);
or U5353 (N_5353,N_596,N_1323);
and U5354 (N_5354,N_858,N_875);
nor U5355 (N_5355,N_628,N_2320);
and U5356 (N_5356,N_3355,N_3450);
or U5357 (N_5357,N_1949,N_3382);
and U5358 (N_5358,N_617,N_1788);
or U5359 (N_5359,N_3031,N_1471);
and U5360 (N_5360,N_3867,N_3239);
xor U5361 (N_5361,N_3329,N_3720);
nand U5362 (N_5362,N_1837,N_3886);
and U5363 (N_5363,N_926,N_2039);
nand U5364 (N_5364,N_1111,N_3461);
nor U5365 (N_5365,N_2368,N_497);
xor U5366 (N_5366,N_3149,N_3352);
nor U5367 (N_5367,N_227,N_2896);
nor U5368 (N_5368,N_1822,N_2436);
xnor U5369 (N_5369,N_1660,N_2310);
xor U5370 (N_5370,N_1739,N_1125);
or U5371 (N_5371,N_2321,N_753);
xor U5372 (N_5372,N_2229,N_2684);
nor U5373 (N_5373,N_3892,N_1134);
or U5374 (N_5374,N_2607,N_3346);
or U5375 (N_5375,N_2943,N_2304);
and U5376 (N_5376,N_3174,N_3037);
nand U5377 (N_5377,N_575,N_456);
xnor U5378 (N_5378,N_704,N_2836);
and U5379 (N_5379,N_3965,N_22);
nor U5380 (N_5380,N_1275,N_2666);
or U5381 (N_5381,N_2488,N_3215);
nand U5382 (N_5382,N_2562,N_1991);
and U5383 (N_5383,N_3484,N_1083);
or U5384 (N_5384,N_404,N_2749);
or U5385 (N_5385,N_3924,N_1052);
nor U5386 (N_5386,N_3010,N_61);
nor U5387 (N_5387,N_2005,N_2672);
or U5388 (N_5388,N_2236,N_1436);
nand U5389 (N_5389,N_2111,N_3479);
or U5390 (N_5390,N_3872,N_1187);
or U5391 (N_5391,N_1624,N_3300);
and U5392 (N_5392,N_3478,N_3181);
nor U5393 (N_5393,N_2641,N_3420);
and U5394 (N_5394,N_1200,N_144);
nor U5395 (N_5395,N_536,N_1058);
xnor U5396 (N_5396,N_3173,N_3771);
and U5397 (N_5397,N_242,N_2238);
and U5398 (N_5398,N_2638,N_2060);
nand U5399 (N_5399,N_1938,N_2648);
and U5400 (N_5400,N_2697,N_2213);
nor U5401 (N_5401,N_2613,N_3935);
nand U5402 (N_5402,N_3489,N_1532);
nor U5403 (N_5403,N_364,N_610);
nand U5404 (N_5404,N_102,N_1919);
nand U5405 (N_5405,N_3548,N_1084);
and U5406 (N_5406,N_2066,N_1274);
nand U5407 (N_5407,N_1277,N_3120);
and U5408 (N_5408,N_1612,N_2067);
xor U5409 (N_5409,N_3981,N_846);
and U5410 (N_5410,N_2686,N_2230);
and U5411 (N_5411,N_998,N_1455);
xnor U5412 (N_5412,N_3022,N_3936);
or U5413 (N_5413,N_2680,N_1986);
or U5414 (N_5414,N_410,N_990);
and U5415 (N_5415,N_2933,N_1201);
nand U5416 (N_5416,N_351,N_3615);
nand U5417 (N_5417,N_2429,N_969);
nor U5418 (N_5418,N_3940,N_323);
nand U5419 (N_5419,N_3114,N_949);
nor U5420 (N_5420,N_601,N_3950);
xor U5421 (N_5421,N_750,N_3508);
or U5422 (N_5422,N_1661,N_187);
or U5423 (N_5423,N_3585,N_2772);
and U5424 (N_5424,N_1444,N_695);
xnor U5425 (N_5425,N_970,N_841);
and U5426 (N_5426,N_2090,N_2341);
xnor U5427 (N_5427,N_3579,N_1866);
nor U5428 (N_5428,N_3366,N_3317);
nand U5429 (N_5429,N_3184,N_344);
nor U5430 (N_5430,N_3041,N_3630);
nand U5431 (N_5431,N_2187,N_1689);
and U5432 (N_5432,N_2528,N_986);
nand U5433 (N_5433,N_2774,N_2347);
nor U5434 (N_5434,N_216,N_1577);
or U5435 (N_5435,N_2164,N_1925);
or U5436 (N_5436,N_3986,N_75);
xnor U5437 (N_5437,N_25,N_861);
nor U5438 (N_5438,N_2704,N_3607);
and U5439 (N_5439,N_895,N_853);
nand U5440 (N_5440,N_3482,N_2816);
or U5441 (N_5441,N_1836,N_2095);
nor U5442 (N_5442,N_1630,N_3882);
nor U5443 (N_5443,N_3849,N_1054);
nand U5444 (N_5444,N_1346,N_2649);
nand U5445 (N_5445,N_588,N_2630);
nor U5446 (N_5446,N_2470,N_2628);
xor U5447 (N_5447,N_3593,N_3112);
nand U5448 (N_5448,N_1603,N_3418);
or U5449 (N_5449,N_356,N_1698);
nor U5450 (N_5450,N_1904,N_3495);
or U5451 (N_5451,N_2149,N_2539);
nor U5452 (N_5452,N_3682,N_1550);
or U5453 (N_5453,N_2226,N_72);
nor U5454 (N_5454,N_2585,N_2125);
and U5455 (N_5455,N_2972,N_2378);
or U5456 (N_5456,N_2297,N_2188);
nor U5457 (N_5457,N_1202,N_698);
nor U5458 (N_5458,N_1747,N_3413);
and U5459 (N_5459,N_2559,N_3561);
or U5460 (N_5460,N_2352,N_2998);
or U5461 (N_5461,N_3925,N_1341);
xor U5462 (N_5462,N_3556,N_687);
and U5463 (N_5463,N_1195,N_211);
nor U5464 (N_5464,N_886,N_2959);
nand U5465 (N_5465,N_3890,N_2681);
xnor U5466 (N_5466,N_3725,N_2841);
and U5467 (N_5467,N_2211,N_2738);
and U5468 (N_5468,N_2237,N_3644);
or U5469 (N_5469,N_2609,N_3608);
or U5470 (N_5470,N_2375,N_1122);
xnor U5471 (N_5471,N_2109,N_3638);
or U5472 (N_5472,N_3218,N_2967);
nand U5473 (N_5473,N_1787,N_3199);
and U5474 (N_5474,N_1584,N_3100);
nor U5475 (N_5475,N_1383,N_303);
nand U5476 (N_5476,N_1127,N_955);
or U5477 (N_5477,N_930,N_3351);
nand U5478 (N_5478,N_1335,N_3383);
nand U5479 (N_5479,N_2317,N_764);
xor U5480 (N_5480,N_2804,N_2905);
xnor U5481 (N_5481,N_417,N_3745);
or U5482 (N_5482,N_3128,N_3198);
nand U5483 (N_5483,N_2773,N_2303);
nand U5484 (N_5484,N_1331,N_1500);
nor U5485 (N_5485,N_3971,N_108);
and U5486 (N_5486,N_2576,N_785);
xor U5487 (N_5487,N_2142,N_3433);
or U5488 (N_5488,N_1018,N_1578);
nor U5489 (N_5489,N_2243,N_2694);
nand U5490 (N_5490,N_1685,N_1374);
and U5491 (N_5491,N_770,N_1647);
nand U5492 (N_5492,N_589,N_1115);
xnor U5493 (N_5493,N_3659,N_1802);
nor U5494 (N_5494,N_3730,N_3012);
or U5495 (N_5495,N_3001,N_3223);
and U5496 (N_5496,N_3897,N_2650);
and U5497 (N_5497,N_657,N_2695);
nor U5498 (N_5498,N_2806,N_335);
and U5499 (N_5499,N_1391,N_2995);
and U5500 (N_5500,N_388,N_1229);
xnor U5501 (N_5501,N_809,N_2863);
xnor U5502 (N_5502,N_3422,N_2296);
and U5503 (N_5503,N_131,N_2632);
nand U5504 (N_5504,N_3493,N_1743);
and U5505 (N_5505,N_3967,N_1327);
nand U5506 (N_5506,N_668,N_988);
or U5507 (N_5507,N_2382,N_2601);
nor U5508 (N_5508,N_994,N_3634);
nand U5509 (N_5509,N_2077,N_3207);
xor U5510 (N_5510,N_1981,N_2455);
xnor U5511 (N_5511,N_494,N_3460);
xor U5512 (N_5512,N_21,N_222);
and U5513 (N_5513,N_540,N_762);
xor U5514 (N_5514,N_78,N_528);
xor U5515 (N_5515,N_2471,N_2415);
nand U5516 (N_5516,N_1543,N_3822);
or U5517 (N_5517,N_255,N_1495);
nor U5518 (N_5518,N_1767,N_286);
xor U5519 (N_5519,N_1073,N_1375);
or U5520 (N_5520,N_2486,N_3514);
and U5521 (N_5521,N_1538,N_868);
nand U5522 (N_5522,N_398,N_2565);
and U5523 (N_5523,N_1390,N_1031);
nand U5524 (N_5524,N_181,N_3912);
and U5525 (N_5525,N_2400,N_3005);
nor U5526 (N_5526,N_173,N_118);
and U5527 (N_5527,N_3385,N_3994);
or U5528 (N_5528,N_2315,N_3711);
and U5529 (N_5529,N_1123,N_940);
and U5530 (N_5530,N_2269,N_3751);
nor U5531 (N_5531,N_1424,N_3498);
or U5532 (N_5532,N_626,N_3288);
or U5533 (N_5533,N_1607,N_1109);
xnor U5534 (N_5534,N_733,N_1371);
nor U5535 (N_5535,N_982,N_59);
nor U5536 (N_5536,N_2265,N_3265);
nor U5537 (N_5537,N_472,N_1542);
xnor U5538 (N_5538,N_92,N_1766);
and U5539 (N_5539,N_3535,N_331);
and U5540 (N_5540,N_3201,N_1235);
nor U5541 (N_5541,N_2232,N_2169);
xnor U5542 (N_5542,N_2796,N_3705);
nor U5543 (N_5543,N_720,N_3899);
nand U5544 (N_5544,N_3934,N_2675);
nor U5545 (N_5545,N_731,N_678);
nand U5546 (N_5546,N_3326,N_3456);
xnor U5547 (N_5547,N_1182,N_1705);
and U5548 (N_5548,N_3386,N_3165);
or U5549 (N_5549,N_3016,N_3075);
and U5550 (N_5550,N_2963,N_899);
nand U5551 (N_5551,N_543,N_2240);
and U5552 (N_5552,N_1770,N_1829);
nor U5553 (N_5553,N_2595,N_2462);
nor U5554 (N_5554,N_1167,N_2828);
or U5555 (N_5555,N_462,N_1003);
or U5556 (N_5556,N_3020,N_3674);
nor U5557 (N_5557,N_3876,N_3708);
xor U5558 (N_5558,N_1974,N_3320);
or U5559 (N_5559,N_3324,N_3134);
nor U5560 (N_5560,N_2929,N_301);
and U5561 (N_5561,N_2542,N_458);
nor U5562 (N_5562,N_19,N_1871);
xnor U5563 (N_5563,N_2131,N_3094);
nor U5564 (N_5564,N_2487,N_439);
xnor U5565 (N_5565,N_60,N_3916);
nand U5566 (N_5566,N_1001,N_2914);
xor U5567 (N_5567,N_478,N_2247);
xor U5568 (N_5568,N_818,N_1926);
nand U5569 (N_5569,N_264,N_2361);
nor U5570 (N_5570,N_1042,N_3035);
or U5571 (N_5571,N_1265,N_2835);
or U5572 (N_5572,N_551,N_2053);
xnor U5573 (N_5573,N_2615,N_1076);
nand U5574 (N_5574,N_2965,N_127);
nand U5575 (N_5575,N_3303,N_3009);
nand U5576 (N_5576,N_2218,N_1340);
xor U5577 (N_5577,N_2979,N_2062);
or U5578 (N_5578,N_2290,N_3250);
and U5579 (N_5579,N_339,N_3750);
xnor U5580 (N_5580,N_3312,N_2530);
or U5581 (N_5581,N_202,N_2634);
and U5582 (N_5582,N_287,N_1772);
nand U5583 (N_5583,N_2926,N_682);
nor U5584 (N_5584,N_2319,N_2350);
and U5585 (N_5585,N_2117,N_166);
or U5586 (N_5586,N_1160,N_643);
nand U5587 (N_5587,N_3989,N_1815);
nor U5588 (N_5588,N_199,N_550);
and U5589 (N_5589,N_1540,N_125);
xnor U5590 (N_5590,N_2766,N_1674);
or U5591 (N_5591,N_3976,N_54);
nor U5592 (N_5592,N_2876,N_489);
xor U5593 (N_5593,N_2282,N_3521);
and U5594 (N_5594,N_322,N_2598);
nor U5595 (N_5595,N_3430,N_2640);
xor U5596 (N_5596,N_3694,N_808);
or U5597 (N_5597,N_1708,N_1388);
xnor U5598 (N_5598,N_622,N_3597);
nand U5599 (N_5599,N_3741,N_289);
xnor U5600 (N_5600,N_1890,N_951);
or U5601 (N_5601,N_3118,N_2941);
and U5602 (N_5602,N_3305,N_151);
nor U5603 (N_5603,N_3898,N_2506);
nor U5604 (N_5604,N_486,N_3789);
nor U5605 (N_5605,N_1797,N_1653);
and U5606 (N_5606,N_3453,N_69);
and U5607 (N_5607,N_426,N_2339);
and U5608 (N_5608,N_1709,N_3735);
or U5609 (N_5609,N_1749,N_1370);
and U5610 (N_5610,N_3411,N_2192);
and U5611 (N_5611,N_2776,N_3306);
or U5612 (N_5612,N_1459,N_3896);
nand U5613 (N_5613,N_893,N_2387);
xnor U5614 (N_5614,N_274,N_468);
and U5615 (N_5615,N_3770,N_1645);
xnor U5616 (N_5616,N_221,N_991);
nand U5617 (N_5617,N_498,N_2978);
xor U5618 (N_5618,N_2502,N_690);
and U5619 (N_5619,N_1493,N_3606);
nand U5620 (N_5620,N_2438,N_1243);
xnor U5621 (N_5621,N_3569,N_1618);
or U5622 (N_5622,N_2482,N_1810);
nor U5623 (N_5623,N_980,N_1070);
nor U5624 (N_5624,N_641,N_2993);
nand U5625 (N_5625,N_2840,N_3946);
nand U5626 (N_5626,N_3282,N_3800);
nand U5627 (N_5627,N_119,N_1219);
nor U5628 (N_5628,N_719,N_1428);
nand U5629 (N_5629,N_3042,N_811);
and U5630 (N_5630,N_3125,N_2372);
nor U5631 (N_5631,N_3906,N_1638);
nor U5632 (N_5632,N_2752,N_3335);
or U5633 (N_5633,N_2597,N_584);
nor U5634 (N_5634,N_3518,N_189);
and U5635 (N_5635,N_3314,N_2299);
xnor U5636 (N_5636,N_945,N_3253);
nor U5637 (N_5637,N_3573,N_2084);
nand U5638 (N_5638,N_2267,N_3077);
nand U5639 (N_5639,N_1321,N_243);
xor U5640 (N_5640,N_1526,N_2719);
or U5641 (N_5641,N_3141,N_3076);
or U5642 (N_5642,N_1915,N_765);
xnor U5643 (N_5643,N_812,N_1750);
or U5644 (N_5644,N_1240,N_2399);
and U5645 (N_5645,N_3690,N_3156);
nand U5646 (N_5646,N_3088,N_43);
nand U5647 (N_5647,N_807,N_787);
and U5648 (N_5648,N_3002,N_1381);
xor U5649 (N_5649,N_1291,N_3919);
and U5650 (N_5650,N_2708,N_3668);
nand U5651 (N_5651,N_966,N_3350);
nand U5652 (N_5652,N_1476,N_2622);
nand U5653 (N_5653,N_3362,N_260);
nand U5654 (N_5654,N_756,N_905);
nor U5655 (N_5655,N_3105,N_2834);
or U5656 (N_5656,N_1000,N_1309);
and U5657 (N_5657,N_1008,N_3591);
nand U5658 (N_5658,N_981,N_1423);
nand U5659 (N_5659,N_310,N_2991);
or U5660 (N_5660,N_614,N_975);
nor U5661 (N_5661,N_3480,N_1521);
and U5662 (N_5662,N_3040,N_1872);
nand U5663 (N_5663,N_2032,N_561);
or U5664 (N_5664,N_1956,N_867);
nand U5665 (N_5665,N_0,N_3527);
or U5666 (N_5666,N_477,N_3991);
or U5667 (N_5667,N_1945,N_2366);
nand U5668 (N_5668,N_3592,N_3170);
nand U5669 (N_5669,N_2291,N_734);
nor U5670 (N_5670,N_3542,N_3166);
and U5671 (N_5671,N_2152,N_80);
or U5672 (N_5672,N_2083,N_1485);
or U5673 (N_5673,N_89,N_1552);
and U5674 (N_5674,N_2180,N_2578);
and U5675 (N_5675,N_680,N_759);
nor U5676 (N_5676,N_2735,N_1588);
xor U5677 (N_5677,N_1302,N_2711);
and U5678 (N_5678,N_1186,N_2612);
xor U5679 (N_5679,N_852,N_126);
and U5680 (N_5680,N_17,N_1306);
and U5681 (N_5681,N_3359,N_3175);
xnor U5682 (N_5682,N_527,N_2391);
nor U5683 (N_5683,N_395,N_984);
nor U5684 (N_5684,N_2503,N_440);
or U5685 (N_5685,N_1811,N_2861);
xor U5686 (N_5686,N_2569,N_2855);
nor U5687 (N_5687,N_3956,N_3192);
xnor U5688 (N_5688,N_1642,N_2159);
xnor U5689 (N_5689,N_3683,N_2961);
or U5690 (N_5690,N_3328,N_912);
and U5691 (N_5691,N_160,N_3081);
and U5692 (N_5692,N_348,N_123);
nor U5693 (N_5693,N_1650,N_2274);
nand U5694 (N_5694,N_1366,N_328);
and U5695 (N_5695,N_2474,N_3970);
xnor U5696 (N_5696,N_1863,N_2107);
nand U5697 (N_5697,N_3315,N_70);
nor U5698 (N_5698,N_2381,N_3255);
nor U5699 (N_5699,N_3666,N_746);
nor U5700 (N_5700,N_206,N_802);
nor U5701 (N_5701,N_3743,N_2549);
or U5702 (N_5702,N_3379,N_2871);
nor U5703 (N_5703,N_2889,N_1679);
or U5704 (N_5704,N_3551,N_1554);
or U5705 (N_5705,N_400,N_2249);
or U5706 (N_5706,N_796,N_1994);
or U5707 (N_5707,N_1759,N_3437);
nand U5708 (N_5708,N_2250,N_484);
xnor U5709 (N_5709,N_3092,N_3129);
and U5710 (N_5710,N_3533,N_487);
nand U5711 (N_5711,N_3945,N_62);
nor U5712 (N_5712,N_1740,N_3554);
xor U5713 (N_5713,N_3921,N_2272);
nor U5714 (N_5714,N_3862,N_1143);
nand U5715 (N_5715,N_1474,N_667);
or U5716 (N_5716,N_1400,N_493);
and U5717 (N_5717,N_68,N_168);
nor U5718 (N_5718,N_2390,N_1491);
or U5719 (N_5719,N_1350,N_2737);
nand U5720 (N_5720,N_3330,N_2830);
or U5721 (N_5721,N_562,N_1299);
nor U5722 (N_5722,N_507,N_3243);
and U5723 (N_5723,N_985,N_2574);
nand U5724 (N_5724,N_1144,N_672);
nor U5725 (N_5725,N_649,N_1786);
nand U5726 (N_5726,N_2145,N_1468);
and U5727 (N_5727,N_3043,N_3086);
or U5728 (N_5728,N_2478,N_492);
xnor U5729 (N_5729,N_2807,N_1347);
and U5730 (N_5730,N_828,N_267);
nor U5731 (N_5731,N_334,N_952);
nand U5732 (N_5732,N_2377,N_2637);
nor U5733 (N_5733,N_296,N_58);
xnor U5734 (N_5734,N_2548,N_3084);
nor U5735 (N_5735,N_3520,N_933);
nor U5736 (N_5736,N_3660,N_1349);
nor U5737 (N_5737,N_2691,N_3785);
xor U5738 (N_5738,N_1859,N_3817);
nand U5739 (N_5739,N_2197,N_1882);
nor U5740 (N_5740,N_1694,N_615);
xor U5741 (N_5741,N_2758,N_2287);
and U5742 (N_5742,N_755,N_3793);
nor U5743 (N_5743,N_2815,N_2472);
nor U5744 (N_5744,N_2261,N_138);
xnor U5745 (N_5745,N_3246,N_3448);
and U5746 (N_5746,N_3262,N_2204);
or U5747 (N_5747,N_2811,N_129);
or U5748 (N_5748,N_1751,N_3167);
nand U5749 (N_5749,N_1192,N_2007);
nand U5750 (N_5750,N_3893,N_2511);
or U5751 (N_5751,N_3345,N_3655);
xor U5752 (N_5752,N_2106,N_2182);
and U5753 (N_5753,N_1211,N_1652);
and U5754 (N_5754,N_745,N_1508);
and U5755 (N_5755,N_1947,N_3089);
and U5756 (N_5756,N_1721,N_2558);
and U5757 (N_5757,N_2002,N_743);
xnor U5758 (N_5758,N_570,N_246);
nor U5759 (N_5759,N_3224,N_3781);
or U5760 (N_5760,N_2533,N_3576);
nand U5761 (N_5761,N_349,N_939);
or U5762 (N_5762,N_1921,N_661);
nor U5763 (N_5763,N_1929,N_257);
or U5764 (N_5764,N_1673,N_3145);
nor U5765 (N_5765,N_1197,N_1403);
nand U5766 (N_5766,N_3526,N_372);
nor U5767 (N_5767,N_3004,N_215);
nand U5768 (N_5768,N_2797,N_3124);
or U5769 (N_5769,N_3494,N_840);
and U5770 (N_5770,N_1969,N_3985);
xnor U5771 (N_5771,N_2420,N_1623);
nand U5772 (N_5772,N_2079,N_3234);
and U5773 (N_5773,N_36,N_2219);
and U5774 (N_5774,N_1338,N_1234);
xnor U5775 (N_5775,N_1930,N_3513);
xor U5776 (N_5776,N_175,N_1027);
nand U5777 (N_5777,N_150,N_2172);
nand U5778 (N_5778,N_2178,N_1742);
and U5779 (N_5779,N_2518,N_3984);
nand U5780 (N_5780,N_2052,N_2767);
or U5781 (N_5781,N_3071,N_894);
nand U5782 (N_5782,N_2936,N_771);
and U5783 (N_5783,N_2677,N_1702);
nand U5784 (N_5784,N_2373,N_1831);
nand U5785 (N_5785,N_1461,N_3632);
nand U5786 (N_5786,N_2477,N_3895);
and U5787 (N_5787,N_2600,N_831);
and U5788 (N_5788,N_368,N_2750);
xor U5789 (N_5789,N_1113,N_258);
nor U5790 (N_5790,N_3179,N_261);
and U5791 (N_5791,N_1910,N_2891);
and U5792 (N_5792,N_2433,N_3467);
xnor U5793 (N_5793,N_804,N_3396);
nor U5794 (N_5794,N_2411,N_2393);
nand U5795 (N_5795,N_2450,N_3852);
or U5796 (N_5796,N_176,N_172);
nand U5797 (N_5797,N_1215,N_365);
nand U5798 (N_5798,N_3821,N_907);
or U5799 (N_5799,N_636,N_2288);
or U5800 (N_5800,N_2354,N_1329);
nand U5801 (N_5801,N_122,N_3503);
or U5802 (N_5802,N_3107,N_519);
nor U5803 (N_5803,N_1451,N_3764);
or U5804 (N_5804,N_3557,N_3373);
or U5805 (N_5805,N_445,N_2460);
xor U5806 (N_5806,N_329,N_3152);
nand U5807 (N_5807,N_2893,N_2802);
nand U5808 (N_5808,N_2923,N_1733);
nor U5809 (N_5809,N_2689,N_3703);
nor U5810 (N_5810,N_2820,N_3594);
nand U5811 (N_5811,N_1539,N_2442);
xnor U5812 (N_5812,N_1824,N_1690);
xnor U5813 (N_5813,N_724,N_2404);
or U5814 (N_5814,N_3187,N_2132);
nand U5815 (N_5815,N_573,N_2143);
nand U5816 (N_5816,N_1844,N_1629);
and U5817 (N_5817,N_3657,N_2325);
or U5818 (N_5818,N_1147,N_3600);
xor U5819 (N_5819,N_913,N_95);
and U5820 (N_5820,N_2813,N_936);
nor U5821 (N_5821,N_3208,N_3677);
and U5822 (N_5822,N_973,N_1867);
nand U5823 (N_5823,N_237,N_3679);
or U5824 (N_5824,N_120,N_1168);
or U5825 (N_5825,N_2078,N_3018);
nand U5826 (N_5826,N_1594,N_1522);
or U5827 (N_5827,N_3870,N_1923);
nor U5828 (N_5828,N_2903,N_448);
or U5829 (N_5829,N_1220,N_2150);
nor U5830 (N_5830,N_953,N_908);
and U5831 (N_5831,N_1354,N_1417);
and U5832 (N_5832,N_1779,N_3749);
nand U5833 (N_5833,N_3633,N_2688);
or U5834 (N_5834,N_1840,N_1140);
nor U5835 (N_5835,N_3629,N_650);
and U5836 (N_5836,N_1322,N_1681);
nand U5837 (N_5837,N_2116,N_3308);
xor U5838 (N_5838,N_270,N_3161);
or U5839 (N_5839,N_2342,N_775);
and U5840 (N_5840,N_814,N_3133);
nand U5841 (N_5841,N_1850,N_291);
or U5842 (N_5842,N_1458,N_1210);
or U5843 (N_5843,N_1502,N_1752);
and U5844 (N_5844,N_3963,N_718);
nor U5845 (N_5845,N_882,N_2907);
xnor U5846 (N_5846,N_1252,N_1279);
nor U5847 (N_5847,N_904,N_674);
nor U5848 (N_5848,N_3231,N_3395);
and U5849 (N_5849,N_2227,N_3570);
nand U5850 (N_5850,N_11,N_9);
or U5851 (N_5851,N_3400,N_2424);
or U5852 (N_5852,N_2009,N_1177);
nor U5853 (N_5853,N_201,N_1627);
xnor U5854 (N_5854,N_2435,N_3571);
and U5855 (N_5855,N_937,N_3017);
nor U5856 (N_5856,N_155,N_844);
or U5857 (N_5857,N_1565,N_3008);
or U5858 (N_5858,N_582,N_713);
nor U5859 (N_5859,N_1807,N_2412);
and U5860 (N_5860,N_229,N_3384);
nand U5861 (N_5861,N_330,N_883);
nand U5862 (N_5862,N_1764,N_1313);
xor U5863 (N_5863,N_1498,N_605);
or U5864 (N_5864,N_1206,N_3717);
nor U5865 (N_5865,N_1019,N_791);
xor U5866 (N_5866,N_3163,N_2856);
nand U5867 (N_5867,N_1078,N_3582);
or U5868 (N_5868,N_1855,N_576);
nor U5869 (N_5869,N_2194,N_2678);
or U5870 (N_5870,N_1021,N_1913);
and U5871 (N_5871,N_1250,N_1696);
xor U5872 (N_5872,N_987,N_732);
xnor U5873 (N_5873,N_1121,N_572);
nor U5874 (N_5874,N_3794,N_2712);
or U5875 (N_5875,N_3874,N_2137);
nor U5876 (N_5876,N_1199,N_3178);
xnor U5877 (N_5877,N_2171,N_1573);
and U5878 (N_5878,N_3425,N_153);
nand U5879 (N_5879,N_3678,N_3164);
xor U5880 (N_5880,N_3728,N_2663);
nor U5881 (N_5881,N_2935,N_2);
nand U5882 (N_5882,N_2394,N_1916);
and U5883 (N_5883,N_3938,N_885);
nand U5884 (N_5884,N_34,N_1062);
or U5885 (N_5885,N_2059,N_1453);
nand U5886 (N_5886,N_1072,N_3501);
or U5887 (N_5887,N_3920,N_2550);
or U5888 (N_5888,N_1534,N_209);
xor U5889 (N_5889,N_1909,N_195);
and U5890 (N_5890,N_1098,N_3653);
nor U5891 (N_5891,N_451,N_3275);
xnor U5892 (N_5892,N_1566,N_3293);
or U5893 (N_5893,N_1466,N_3206);
nor U5894 (N_5894,N_2224,N_2647);
and U5895 (N_5895,N_437,N_2351);
nor U5896 (N_5896,N_942,N_3812);
and U5897 (N_5897,N_2075,N_3990);
nand U5898 (N_5898,N_1330,N_177);
nand U5899 (N_5899,N_2819,N_2895);
and U5900 (N_5900,N_1835,N_280);
xnor U5901 (N_5901,N_900,N_443);
nor U5902 (N_5902,N_3095,N_1303);
or U5903 (N_5903,N_1137,N_2430);
and U5904 (N_5904,N_1659,N_2340);
and U5905 (N_5905,N_163,N_164);
nand U5906 (N_5906,N_578,N_3132);
or U5907 (N_5907,N_79,N_170);
nor U5908 (N_5908,N_3810,N_3808);
nand U5909 (N_5909,N_3244,N_3664);
or U5910 (N_5910,N_1662,N_2938);
or U5911 (N_5911,N_2949,N_2014);
and U5912 (N_5912,N_1970,N_2973);
nor U5913 (N_5913,N_1571,N_262);
nand U5914 (N_5914,N_3613,N_184);
nor U5915 (N_5915,N_2902,N_145);
xnor U5916 (N_5916,N_2345,N_3587);
or U5917 (N_5917,N_3154,N_3854);
xor U5918 (N_5918,N_1094,N_107);
and U5919 (N_5919,N_1188,N_1156);
xor U5920 (N_5920,N_705,N_3663);
and U5921 (N_5921,N_2467,N_592);
xor U5922 (N_5922,N_2328,N_938);
nand U5923 (N_5923,N_2560,N_1405);
or U5924 (N_5924,N_2068,N_1854);
nand U5925 (N_5925,N_1954,N_1281);
or U5926 (N_5926,N_3552,N_1204);
nor U5927 (N_5927,N_2343,N_586);
xor U5928 (N_5928,N_798,N_1004);
nand U5929 (N_5929,N_3079,N_1609);
and U5930 (N_5930,N_1719,N_3744);
and U5931 (N_5931,N_2507,N_1467);
or U5932 (N_5932,N_854,N_1012);
xor U5933 (N_5933,N_3401,N_2832);
nand U5934 (N_5934,N_2138,N_2355);
and U5935 (N_5935,N_2335,N_2519);
xor U5936 (N_5936,N_204,N_1036);
and U5937 (N_5937,N_1796,N_2081);
nor U5938 (N_5938,N_3693,N_2593);
nor U5939 (N_5939,N_1940,N_2611);
xnor U5940 (N_5940,N_1657,N_1545);
xor U5941 (N_5941,N_2705,N_1718);
xor U5942 (N_5942,N_1397,N_504);
and U5943 (N_5943,N_3446,N_2584);
or U5944 (N_5944,N_1535,N_1948);
and U5945 (N_5945,N_1825,N_2385);
or U5946 (N_5946,N_74,N_154);
and U5947 (N_5947,N_1402,N_2323);
nand U5948 (N_5948,N_2421,N_40);
and U5949 (N_5949,N_931,N_3560);
or U5950 (N_5950,N_1897,N_2198);
nand U5951 (N_5951,N_3539,N_1794);
nor U5952 (N_5952,N_850,N_3807);
xor U5953 (N_5953,N_3221,N_2692);
and U5954 (N_5954,N_396,N_879);
nand U5955 (N_5955,N_763,N_3428);
and U5956 (N_5956,N_333,N_3734);
xor U5957 (N_5957,N_2252,N_3119);
nand U5958 (N_5958,N_208,N_305);
xor U5959 (N_5959,N_2206,N_2458);
nand U5960 (N_5960,N_24,N_77);
xor U5961 (N_5961,N_3408,N_210);
or U5962 (N_5962,N_3522,N_529);
or U5963 (N_5963,N_405,N_2266);
or U5964 (N_5964,N_3375,N_1218);
or U5965 (N_5965,N_342,N_521);
xnor U5966 (N_5966,N_1487,N_2313);
nand U5967 (N_5967,N_3753,N_736);
nand U5968 (N_5968,N_1557,N_3726);
xor U5969 (N_5969,N_1117,N_2135);
and U5970 (N_5970,N_2233,N_2016);
or U5971 (N_5971,N_3485,N_158);
xnor U5972 (N_5972,N_932,N_471);
or U5973 (N_5973,N_1581,N_2727);
nor U5974 (N_5974,N_2906,N_2779);
nand U5975 (N_5975,N_3488,N_2934);
or U5976 (N_5976,N_1995,N_2818);
and U5977 (N_5977,N_3773,N_2513);
and U5978 (N_5978,N_3755,N_3403);
xor U5979 (N_5979,N_1159,N_327);
xor U5980 (N_5980,N_3083,N_2928);
xor U5981 (N_5981,N_3879,N_1744);
xor U5982 (N_5982,N_290,N_670);
and U5983 (N_5983,N_1966,N_1116);
xnor U5984 (N_5984,N_834,N_1900);
nor U5985 (N_5985,N_2322,N_1048);
nor U5986 (N_5986,N_2887,N_821);
nor U5987 (N_5987,N_2846,N_1515);
nand U5988 (N_5988,N_646,N_3796);
or U5989 (N_5989,N_859,N_2254);
nand U5990 (N_5990,N_1551,N_84);
nor U5991 (N_5991,N_459,N_2141);
or U5992 (N_5992,N_1792,N_3878);
xor U5993 (N_5993,N_338,N_1207);
and U5994 (N_5994,N_1090,N_3927);
or U5995 (N_5995,N_757,N_403);
xor U5996 (N_5996,N_3712,N_1130);
nand U5997 (N_5997,N_1678,N_2473);
xnor U5998 (N_5998,N_2017,N_2134);
xor U5999 (N_5999,N_1242,N_2920);
xnor U6000 (N_6000,N_1825,N_1005);
and U6001 (N_6001,N_1238,N_3601);
or U6002 (N_6002,N_712,N_884);
xnor U6003 (N_6003,N_2805,N_2165);
or U6004 (N_6004,N_3344,N_1727);
nor U6005 (N_6005,N_153,N_3726);
nor U6006 (N_6006,N_3775,N_3965);
xor U6007 (N_6007,N_36,N_841);
nand U6008 (N_6008,N_3968,N_1686);
and U6009 (N_6009,N_657,N_1148);
or U6010 (N_6010,N_3945,N_3169);
or U6011 (N_6011,N_1751,N_2921);
or U6012 (N_6012,N_3045,N_2929);
xnor U6013 (N_6013,N_221,N_2388);
nor U6014 (N_6014,N_1377,N_2778);
xnor U6015 (N_6015,N_1650,N_3264);
or U6016 (N_6016,N_1350,N_2136);
xor U6017 (N_6017,N_1106,N_2230);
and U6018 (N_6018,N_2528,N_2065);
xnor U6019 (N_6019,N_704,N_3177);
and U6020 (N_6020,N_3636,N_3396);
nor U6021 (N_6021,N_2264,N_581);
or U6022 (N_6022,N_3930,N_1526);
and U6023 (N_6023,N_125,N_127);
nand U6024 (N_6024,N_3571,N_988);
and U6025 (N_6025,N_1260,N_6);
and U6026 (N_6026,N_1002,N_2851);
nand U6027 (N_6027,N_2695,N_111);
or U6028 (N_6028,N_1988,N_1886);
nor U6029 (N_6029,N_164,N_760);
and U6030 (N_6030,N_3391,N_1925);
nand U6031 (N_6031,N_1471,N_2232);
xnor U6032 (N_6032,N_667,N_3391);
nand U6033 (N_6033,N_1475,N_2999);
or U6034 (N_6034,N_495,N_3872);
nor U6035 (N_6035,N_2073,N_276);
xnor U6036 (N_6036,N_143,N_3305);
or U6037 (N_6037,N_207,N_836);
nand U6038 (N_6038,N_3993,N_742);
and U6039 (N_6039,N_3454,N_293);
and U6040 (N_6040,N_575,N_366);
xor U6041 (N_6041,N_1406,N_2636);
xnor U6042 (N_6042,N_2389,N_3776);
nor U6043 (N_6043,N_2012,N_2774);
and U6044 (N_6044,N_1016,N_3972);
xnor U6045 (N_6045,N_3858,N_626);
and U6046 (N_6046,N_3998,N_3836);
nor U6047 (N_6047,N_1172,N_2995);
xor U6048 (N_6048,N_3116,N_1349);
or U6049 (N_6049,N_3084,N_2056);
and U6050 (N_6050,N_2803,N_779);
and U6051 (N_6051,N_3082,N_1377);
and U6052 (N_6052,N_1779,N_2467);
and U6053 (N_6053,N_941,N_2064);
and U6054 (N_6054,N_552,N_240);
xor U6055 (N_6055,N_3341,N_2612);
nor U6056 (N_6056,N_1764,N_2360);
nor U6057 (N_6057,N_1724,N_2238);
nand U6058 (N_6058,N_2403,N_1068);
nor U6059 (N_6059,N_637,N_1815);
nand U6060 (N_6060,N_2563,N_688);
nor U6061 (N_6061,N_3650,N_2199);
or U6062 (N_6062,N_2908,N_1991);
nand U6063 (N_6063,N_2998,N_3602);
nand U6064 (N_6064,N_3622,N_3753);
nand U6065 (N_6065,N_3844,N_3815);
nor U6066 (N_6066,N_3831,N_2352);
or U6067 (N_6067,N_919,N_59);
xnor U6068 (N_6068,N_1267,N_356);
or U6069 (N_6069,N_3632,N_1151);
or U6070 (N_6070,N_1267,N_1203);
xor U6071 (N_6071,N_371,N_34);
nor U6072 (N_6072,N_1605,N_3866);
nand U6073 (N_6073,N_3988,N_2113);
and U6074 (N_6074,N_3858,N_1363);
nor U6075 (N_6075,N_823,N_3467);
xnor U6076 (N_6076,N_2696,N_2620);
xor U6077 (N_6077,N_1347,N_3674);
nand U6078 (N_6078,N_2878,N_2271);
and U6079 (N_6079,N_3822,N_179);
or U6080 (N_6080,N_600,N_125);
xnor U6081 (N_6081,N_3316,N_88);
or U6082 (N_6082,N_1641,N_2608);
xor U6083 (N_6083,N_293,N_3685);
xnor U6084 (N_6084,N_3612,N_3328);
xnor U6085 (N_6085,N_1262,N_3741);
nor U6086 (N_6086,N_2678,N_1225);
xor U6087 (N_6087,N_3843,N_2767);
or U6088 (N_6088,N_676,N_2917);
xor U6089 (N_6089,N_1557,N_67);
xor U6090 (N_6090,N_2382,N_1883);
and U6091 (N_6091,N_217,N_3445);
or U6092 (N_6092,N_2323,N_1045);
and U6093 (N_6093,N_3164,N_110);
nand U6094 (N_6094,N_3367,N_2555);
or U6095 (N_6095,N_1205,N_1025);
and U6096 (N_6096,N_1318,N_2549);
nor U6097 (N_6097,N_316,N_1116);
nor U6098 (N_6098,N_3817,N_3978);
and U6099 (N_6099,N_190,N_2160);
or U6100 (N_6100,N_3781,N_1404);
nand U6101 (N_6101,N_1378,N_685);
xnor U6102 (N_6102,N_213,N_3261);
xnor U6103 (N_6103,N_144,N_1343);
xor U6104 (N_6104,N_3,N_151);
or U6105 (N_6105,N_1661,N_2014);
nand U6106 (N_6106,N_1197,N_3129);
and U6107 (N_6107,N_830,N_815);
or U6108 (N_6108,N_2307,N_1748);
and U6109 (N_6109,N_3654,N_354);
and U6110 (N_6110,N_1111,N_3942);
and U6111 (N_6111,N_2184,N_682);
or U6112 (N_6112,N_640,N_1642);
or U6113 (N_6113,N_3018,N_2121);
nand U6114 (N_6114,N_3771,N_360);
xor U6115 (N_6115,N_1258,N_2399);
nor U6116 (N_6116,N_1596,N_2392);
nor U6117 (N_6117,N_152,N_3219);
xor U6118 (N_6118,N_1972,N_2318);
or U6119 (N_6119,N_2258,N_1002);
xor U6120 (N_6120,N_2468,N_2076);
and U6121 (N_6121,N_476,N_3085);
nor U6122 (N_6122,N_1984,N_895);
nor U6123 (N_6123,N_949,N_3438);
or U6124 (N_6124,N_2910,N_3669);
or U6125 (N_6125,N_1503,N_1799);
and U6126 (N_6126,N_1351,N_2068);
and U6127 (N_6127,N_199,N_1629);
xnor U6128 (N_6128,N_630,N_2083);
or U6129 (N_6129,N_576,N_2239);
or U6130 (N_6130,N_3400,N_676);
nor U6131 (N_6131,N_219,N_2703);
or U6132 (N_6132,N_3159,N_835);
or U6133 (N_6133,N_2696,N_919);
nand U6134 (N_6134,N_3827,N_3536);
nor U6135 (N_6135,N_2666,N_1901);
or U6136 (N_6136,N_1702,N_3897);
nand U6137 (N_6137,N_1845,N_3638);
or U6138 (N_6138,N_337,N_1790);
nand U6139 (N_6139,N_187,N_3520);
and U6140 (N_6140,N_3757,N_583);
xor U6141 (N_6141,N_195,N_2480);
or U6142 (N_6142,N_2932,N_666);
or U6143 (N_6143,N_2470,N_2575);
nor U6144 (N_6144,N_1991,N_713);
or U6145 (N_6145,N_1564,N_1415);
or U6146 (N_6146,N_351,N_227);
nand U6147 (N_6147,N_641,N_2154);
nand U6148 (N_6148,N_3389,N_3270);
nand U6149 (N_6149,N_2322,N_1209);
nor U6150 (N_6150,N_2993,N_1942);
nor U6151 (N_6151,N_576,N_212);
xnor U6152 (N_6152,N_3540,N_927);
nor U6153 (N_6153,N_2484,N_12);
and U6154 (N_6154,N_3662,N_1701);
and U6155 (N_6155,N_1789,N_1753);
nor U6156 (N_6156,N_1292,N_3764);
and U6157 (N_6157,N_3790,N_3034);
and U6158 (N_6158,N_2738,N_2866);
nor U6159 (N_6159,N_1230,N_333);
and U6160 (N_6160,N_1259,N_2424);
or U6161 (N_6161,N_2343,N_423);
nor U6162 (N_6162,N_2576,N_720);
and U6163 (N_6163,N_1270,N_372);
or U6164 (N_6164,N_326,N_1907);
nand U6165 (N_6165,N_788,N_2944);
xnor U6166 (N_6166,N_136,N_1532);
or U6167 (N_6167,N_1224,N_1532);
or U6168 (N_6168,N_2920,N_1937);
and U6169 (N_6169,N_1462,N_2134);
nor U6170 (N_6170,N_2424,N_1918);
and U6171 (N_6171,N_1041,N_3375);
xnor U6172 (N_6172,N_83,N_2557);
nand U6173 (N_6173,N_1436,N_1200);
xnor U6174 (N_6174,N_2446,N_583);
or U6175 (N_6175,N_3876,N_1974);
and U6176 (N_6176,N_2652,N_3642);
nand U6177 (N_6177,N_2603,N_2542);
nor U6178 (N_6178,N_2072,N_280);
xnor U6179 (N_6179,N_2390,N_236);
nor U6180 (N_6180,N_2436,N_1580);
nor U6181 (N_6181,N_3040,N_2715);
or U6182 (N_6182,N_847,N_1246);
nor U6183 (N_6183,N_2298,N_2730);
nor U6184 (N_6184,N_3039,N_2978);
xnor U6185 (N_6185,N_3100,N_1334);
nor U6186 (N_6186,N_2014,N_3863);
nand U6187 (N_6187,N_1814,N_1200);
xor U6188 (N_6188,N_1650,N_1250);
or U6189 (N_6189,N_1211,N_530);
xnor U6190 (N_6190,N_3081,N_3528);
and U6191 (N_6191,N_3529,N_3552);
xor U6192 (N_6192,N_3818,N_2198);
or U6193 (N_6193,N_1239,N_58);
nor U6194 (N_6194,N_2626,N_3641);
and U6195 (N_6195,N_2118,N_859);
nor U6196 (N_6196,N_1038,N_3761);
nor U6197 (N_6197,N_1833,N_3615);
nor U6198 (N_6198,N_1353,N_2862);
nor U6199 (N_6199,N_2872,N_2346);
and U6200 (N_6200,N_2758,N_805);
nand U6201 (N_6201,N_829,N_3979);
nand U6202 (N_6202,N_1176,N_3461);
or U6203 (N_6203,N_3979,N_3748);
xor U6204 (N_6204,N_865,N_1926);
nor U6205 (N_6205,N_681,N_341);
nand U6206 (N_6206,N_2321,N_222);
nand U6207 (N_6207,N_193,N_3872);
nor U6208 (N_6208,N_1775,N_1233);
or U6209 (N_6209,N_1939,N_3817);
xnor U6210 (N_6210,N_187,N_3780);
nor U6211 (N_6211,N_3303,N_1740);
nor U6212 (N_6212,N_1731,N_1379);
nand U6213 (N_6213,N_983,N_2803);
nor U6214 (N_6214,N_962,N_3595);
xnor U6215 (N_6215,N_3623,N_3205);
nor U6216 (N_6216,N_2253,N_3746);
nand U6217 (N_6217,N_1377,N_2923);
xor U6218 (N_6218,N_3174,N_1610);
nor U6219 (N_6219,N_1370,N_1755);
nand U6220 (N_6220,N_1252,N_824);
xnor U6221 (N_6221,N_1599,N_3952);
nor U6222 (N_6222,N_2918,N_2885);
or U6223 (N_6223,N_131,N_1666);
nor U6224 (N_6224,N_2412,N_1800);
or U6225 (N_6225,N_390,N_1327);
xnor U6226 (N_6226,N_528,N_818);
nand U6227 (N_6227,N_912,N_3212);
and U6228 (N_6228,N_1118,N_3855);
or U6229 (N_6229,N_3755,N_174);
and U6230 (N_6230,N_2637,N_379);
xor U6231 (N_6231,N_2393,N_2571);
nor U6232 (N_6232,N_1561,N_3750);
and U6233 (N_6233,N_832,N_156);
xor U6234 (N_6234,N_981,N_1281);
xor U6235 (N_6235,N_2703,N_3766);
nand U6236 (N_6236,N_2068,N_3563);
and U6237 (N_6237,N_1716,N_1897);
xor U6238 (N_6238,N_560,N_1712);
and U6239 (N_6239,N_3074,N_3655);
xor U6240 (N_6240,N_1019,N_1124);
xnor U6241 (N_6241,N_3679,N_933);
or U6242 (N_6242,N_2273,N_3758);
or U6243 (N_6243,N_452,N_2191);
nor U6244 (N_6244,N_3410,N_492);
nor U6245 (N_6245,N_3841,N_2602);
and U6246 (N_6246,N_2073,N_2201);
nand U6247 (N_6247,N_2530,N_1437);
nor U6248 (N_6248,N_2301,N_2871);
nand U6249 (N_6249,N_3342,N_3558);
or U6250 (N_6250,N_1681,N_1617);
xnor U6251 (N_6251,N_2380,N_991);
nor U6252 (N_6252,N_1210,N_2141);
xor U6253 (N_6253,N_2429,N_3959);
nor U6254 (N_6254,N_3076,N_894);
and U6255 (N_6255,N_2941,N_1680);
and U6256 (N_6256,N_726,N_3587);
nor U6257 (N_6257,N_1179,N_1255);
xnor U6258 (N_6258,N_739,N_201);
nor U6259 (N_6259,N_190,N_3434);
nor U6260 (N_6260,N_853,N_2630);
or U6261 (N_6261,N_1216,N_3310);
nor U6262 (N_6262,N_3697,N_1855);
nor U6263 (N_6263,N_2894,N_3961);
nand U6264 (N_6264,N_980,N_227);
and U6265 (N_6265,N_2866,N_140);
and U6266 (N_6266,N_2281,N_505);
xnor U6267 (N_6267,N_218,N_1613);
nor U6268 (N_6268,N_3516,N_160);
xnor U6269 (N_6269,N_2053,N_799);
nor U6270 (N_6270,N_1910,N_1195);
nor U6271 (N_6271,N_3236,N_3355);
nor U6272 (N_6272,N_3241,N_1388);
xnor U6273 (N_6273,N_711,N_1707);
or U6274 (N_6274,N_1615,N_185);
or U6275 (N_6275,N_3837,N_892);
or U6276 (N_6276,N_2,N_1777);
xnor U6277 (N_6277,N_148,N_2729);
nand U6278 (N_6278,N_1350,N_2345);
xnor U6279 (N_6279,N_2876,N_1877);
and U6280 (N_6280,N_1102,N_3859);
xor U6281 (N_6281,N_1184,N_69);
nor U6282 (N_6282,N_3021,N_1084);
nand U6283 (N_6283,N_3092,N_3108);
or U6284 (N_6284,N_561,N_937);
and U6285 (N_6285,N_2549,N_181);
nor U6286 (N_6286,N_2754,N_1459);
xor U6287 (N_6287,N_2180,N_941);
nor U6288 (N_6288,N_3004,N_2204);
xor U6289 (N_6289,N_3445,N_1965);
nor U6290 (N_6290,N_562,N_1167);
xnor U6291 (N_6291,N_3053,N_579);
or U6292 (N_6292,N_2323,N_1129);
and U6293 (N_6293,N_1074,N_472);
nand U6294 (N_6294,N_1299,N_1719);
nand U6295 (N_6295,N_2200,N_920);
and U6296 (N_6296,N_464,N_1194);
xnor U6297 (N_6297,N_1208,N_708);
nand U6298 (N_6298,N_3848,N_3529);
xor U6299 (N_6299,N_3077,N_3328);
xor U6300 (N_6300,N_962,N_1630);
or U6301 (N_6301,N_3253,N_1004);
nand U6302 (N_6302,N_620,N_1211);
nand U6303 (N_6303,N_1674,N_1331);
nor U6304 (N_6304,N_2543,N_3067);
nand U6305 (N_6305,N_3756,N_455);
or U6306 (N_6306,N_1579,N_637);
nor U6307 (N_6307,N_572,N_1152);
nand U6308 (N_6308,N_2614,N_664);
xnor U6309 (N_6309,N_3660,N_988);
nor U6310 (N_6310,N_1654,N_3586);
xor U6311 (N_6311,N_3131,N_537);
or U6312 (N_6312,N_3799,N_1736);
and U6313 (N_6313,N_1821,N_1874);
xnor U6314 (N_6314,N_756,N_3380);
or U6315 (N_6315,N_1994,N_2916);
nand U6316 (N_6316,N_1365,N_2327);
or U6317 (N_6317,N_2084,N_2073);
xnor U6318 (N_6318,N_1682,N_2901);
or U6319 (N_6319,N_797,N_1070);
nor U6320 (N_6320,N_3904,N_3589);
nor U6321 (N_6321,N_1480,N_2743);
nand U6322 (N_6322,N_3717,N_666);
xor U6323 (N_6323,N_2373,N_2527);
and U6324 (N_6324,N_3359,N_971);
or U6325 (N_6325,N_1595,N_1406);
xnor U6326 (N_6326,N_3860,N_1457);
or U6327 (N_6327,N_3979,N_2330);
xor U6328 (N_6328,N_1713,N_858);
or U6329 (N_6329,N_2509,N_3655);
nand U6330 (N_6330,N_3335,N_1406);
nor U6331 (N_6331,N_2054,N_3714);
nor U6332 (N_6332,N_3012,N_3454);
nand U6333 (N_6333,N_3491,N_837);
and U6334 (N_6334,N_550,N_3412);
or U6335 (N_6335,N_3539,N_3615);
or U6336 (N_6336,N_1076,N_2543);
xor U6337 (N_6337,N_49,N_1706);
or U6338 (N_6338,N_55,N_769);
and U6339 (N_6339,N_785,N_462);
and U6340 (N_6340,N_1476,N_2337);
or U6341 (N_6341,N_648,N_299);
xnor U6342 (N_6342,N_1121,N_1079);
nand U6343 (N_6343,N_3445,N_1212);
or U6344 (N_6344,N_3510,N_1221);
nand U6345 (N_6345,N_1710,N_2257);
nand U6346 (N_6346,N_2186,N_3230);
nand U6347 (N_6347,N_1519,N_3268);
xnor U6348 (N_6348,N_192,N_2120);
nand U6349 (N_6349,N_131,N_673);
nand U6350 (N_6350,N_1159,N_3649);
or U6351 (N_6351,N_532,N_3971);
nand U6352 (N_6352,N_3683,N_2099);
or U6353 (N_6353,N_532,N_1986);
nor U6354 (N_6354,N_3286,N_3538);
xnor U6355 (N_6355,N_3366,N_3101);
and U6356 (N_6356,N_2381,N_3948);
or U6357 (N_6357,N_1658,N_175);
nor U6358 (N_6358,N_3659,N_3370);
or U6359 (N_6359,N_3970,N_3402);
and U6360 (N_6360,N_984,N_454);
or U6361 (N_6361,N_3892,N_3670);
and U6362 (N_6362,N_3450,N_2382);
xor U6363 (N_6363,N_1336,N_1364);
or U6364 (N_6364,N_2014,N_3700);
xnor U6365 (N_6365,N_1611,N_3036);
nor U6366 (N_6366,N_1132,N_517);
or U6367 (N_6367,N_1508,N_2315);
nor U6368 (N_6368,N_3116,N_1035);
nor U6369 (N_6369,N_1284,N_415);
nand U6370 (N_6370,N_3503,N_3972);
and U6371 (N_6371,N_684,N_2100);
nor U6372 (N_6372,N_1238,N_3998);
and U6373 (N_6373,N_2854,N_812);
nand U6374 (N_6374,N_985,N_2895);
nor U6375 (N_6375,N_117,N_1636);
or U6376 (N_6376,N_1619,N_1331);
xor U6377 (N_6377,N_713,N_135);
nand U6378 (N_6378,N_841,N_1295);
nand U6379 (N_6379,N_70,N_2307);
or U6380 (N_6380,N_2257,N_1735);
nand U6381 (N_6381,N_2730,N_1543);
and U6382 (N_6382,N_1179,N_1877);
nor U6383 (N_6383,N_1359,N_293);
nor U6384 (N_6384,N_2119,N_2779);
xnor U6385 (N_6385,N_1456,N_1600);
xnor U6386 (N_6386,N_1587,N_1919);
nor U6387 (N_6387,N_2501,N_3930);
xor U6388 (N_6388,N_3279,N_1180);
and U6389 (N_6389,N_728,N_3092);
nor U6390 (N_6390,N_3599,N_926);
and U6391 (N_6391,N_2666,N_3549);
xnor U6392 (N_6392,N_978,N_1932);
and U6393 (N_6393,N_2949,N_1397);
nand U6394 (N_6394,N_523,N_321);
or U6395 (N_6395,N_906,N_2150);
nor U6396 (N_6396,N_2782,N_3818);
xnor U6397 (N_6397,N_3077,N_230);
xnor U6398 (N_6398,N_1940,N_2928);
xnor U6399 (N_6399,N_777,N_1392);
nor U6400 (N_6400,N_3405,N_1162);
nor U6401 (N_6401,N_2320,N_884);
nand U6402 (N_6402,N_2859,N_32);
nand U6403 (N_6403,N_338,N_656);
and U6404 (N_6404,N_2049,N_555);
nor U6405 (N_6405,N_1907,N_3352);
and U6406 (N_6406,N_3860,N_2006);
nor U6407 (N_6407,N_1219,N_1293);
nor U6408 (N_6408,N_556,N_1870);
and U6409 (N_6409,N_3691,N_1692);
and U6410 (N_6410,N_2499,N_2004);
or U6411 (N_6411,N_3358,N_3902);
xor U6412 (N_6412,N_578,N_1693);
or U6413 (N_6413,N_1437,N_357);
nand U6414 (N_6414,N_2180,N_2298);
nor U6415 (N_6415,N_142,N_399);
or U6416 (N_6416,N_3695,N_3850);
or U6417 (N_6417,N_2133,N_2895);
nand U6418 (N_6418,N_2884,N_1802);
or U6419 (N_6419,N_294,N_3422);
nor U6420 (N_6420,N_265,N_2321);
nor U6421 (N_6421,N_1821,N_2608);
and U6422 (N_6422,N_2159,N_3377);
and U6423 (N_6423,N_3994,N_258);
xor U6424 (N_6424,N_3373,N_3354);
xnor U6425 (N_6425,N_293,N_301);
nand U6426 (N_6426,N_1360,N_2980);
nor U6427 (N_6427,N_1629,N_140);
nand U6428 (N_6428,N_3437,N_3120);
nand U6429 (N_6429,N_1066,N_2183);
xnor U6430 (N_6430,N_763,N_824);
and U6431 (N_6431,N_2255,N_119);
nand U6432 (N_6432,N_3042,N_2037);
nor U6433 (N_6433,N_3465,N_3124);
or U6434 (N_6434,N_1985,N_499);
or U6435 (N_6435,N_1984,N_1004);
or U6436 (N_6436,N_3239,N_3475);
nor U6437 (N_6437,N_427,N_13);
or U6438 (N_6438,N_3895,N_3622);
nor U6439 (N_6439,N_857,N_2620);
nand U6440 (N_6440,N_2355,N_756);
and U6441 (N_6441,N_105,N_2742);
or U6442 (N_6442,N_3232,N_3926);
or U6443 (N_6443,N_893,N_2222);
nor U6444 (N_6444,N_3051,N_2406);
or U6445 (N_6445,N_3858,N_1588);
or U6446 (N_6446,N_3517,N_3333);
nand U6447 (N_6447,N_1946,N_2150);
nor U6448 (N_6448,N_3776,N_2535);
and U6449 (N_6449,N_54,N_2329);
and U6450 (N_6450,N_3141,N_528);
and U6451 (N_6451,N_3967,N_1693);
or U6452 (N_6452,N_169,N_1974);
nand U6453 (N_6453,N_966,N_1384);
xor U6454 (N_6454,N_1558,N_1018);
and U6455 (N_6455,N_1496,N_1595);
nand U6456 (N_6456,N_3113,N_2921);
nand U6457 (N_6457,N_3822,N_1945);
nand U6458 (N_6458,N_3010,N_2181);
nor U6459 (N_6459,N_150,N_7);
or U6460 (N_6460,N_266,N_1336);
and U6461 (N_6461,N_3277,N_1214);
and U6462 (N_6462,N_809,N_391);
nand U6463 (N_6463,N_3212,N_124);
or U6464 (N_6464,N_3037,N_3664);
and U6465 (N_6465,N_523,N_3406);
nor U6466 (N_6466,N_2059,N_3854);
nor U6467 (N_6467,N_3084,N_532);
and U6468 (N_6468,N_2815,N_1421);
xor U6469 (N_6469,N_507,N_3545);
or U6470 (N_6470,N_1254,N_3600);
nor U6471 (N_6471,N_1486,N_452);
nor U6472 (N_6472,N_3922,N_713);
nor U6473 (N_6473,N_324,N_3199);
and U6474 (N_6474,N_3486,N_3234);
or U6475 (N_6475,N_2686,N_408);
and U6476 (N_6476,N_2106,N_1712);
xor U6477 (N_6477,N_3236,N_3836);
xnor U6478 (N_6478,N_2855,N_2291);
or U6479 (N_6479,N_3074,N_3985);
nor U6480 (N_6480,N_1718,N_1865);
or U6481 (N_6481,N_2197,N_1921);
nor U6482 (N_6482,N_2625,N_240);
and U6483 (N_6483,N_1334,N_569);
and U6484 (N_6484,N_2799,N_3302);
nand U6485 (N_6485,N_1684,N_2158);
nor U6486 (N_6486,N_471,N_345);
nor U6487 (N_6487,N_3009,N_3117);
or U6488 (N_6488,N_3533,N_110);
or U6489 (N_6489,N_920,N_820);
or U6490 (N_6490,N_3484,N_3227);
xnor U6491 (N_6491,N_613,N_1622);
nand U6492 (N_6492,N_2217,N_3254);
xor U6493 (N_6493,N_65,N_2276);
nand U6494 (N_6494,N_319,N_3907);
xor U6495 (N_6495,N_2490,N_2014);
or U6496 (N_6496,N_2447,N_903);
nor U6497 (N_6497,N_667,N_3249);
nor U6498 (N_6498,N_3713,N_1108);
or U6499 (N_6499,N_3755,N_2250);
and U6500 (N_6500,N_3299,N_1522);
nor U6501 (N_6501,N_2983,N_289);
xor U6502 (N_6502,N_954,N_685);
nand U6503 (N_6503,N_2693,N_1599);
nor U6504 (N_6504,N_3938,N_480);
or U6505 (N_6505,N_223,N_3346);
xnor U6506 (N_6506,N_1032,N_576);
xnor U6507 (N_6507,N_1497,N_242);
nand U6508 (N_6508,N_353,N_2387);
nor U6509 (N_6509,N_3480,N_1795);
and U6510 (N_6510,N_1001,N_399);
nor U6511 (N_6511,N_2374,N_1244);
xnor U6512 (N_6512,N_2013,N_3434);
xnor U6513 (N_6513,N_3181,N_1128);
and U6514 (N_6514,N_1377,N_2591);
nor U6515 (N_6515,N_2256,N_3057);
nand U6516 (N_6516,N_2249,N_1770);
nor U6517 (N_6517,N_2638,N_1626);
nand U6518 (N_6518,N_3281,N_1189);
and U6519 (N_6519,N_2117,N_3835);
nor U6520 (N_6520,N_1136,N_3986);
nor U6521 (N_6521,N_1467,N_759);
xnor U6522 (N_6522,N_1945,N_2178);
nand U6523 (N_6523,N_2762,N_2480);
nor U6524 (N_6524,N_3529,N_216);
nor U6525 (N_6525,N_1002,N_366);
nor U6526 (N_6526,N_2628,N_1594);
nand U6527 (N_6527,N_139,N_669);
or U6528 (N_6528,N_3679,N_3588);
nor U6529 (N_6529,N_1580,N_2629);
nor U6530 (N_6530,N_384,N_2151);
nor U6531 (N_6531,N_1420,N_688);
nor U6532 (N_6532,N_1903,N_1958);
xnor U6533 (N_6533,N_1499,N_3301);
or U6534 (N_6534,N_1218,N_2883);
and U6535 (N_6535,N_1801,N_3328);
xnor U6536 (N_6536,N_675,N_390);
nand U6537 (N_6537,N_735,N_2843);
nor U6538 (N_6538,N_3938,N_3647);
and U6539 (N_6539,N_762,N_1255);
nor U6540 (N_6540,N_2417,N_443);
nand U6541 (N_6541,N_1350,N_1556);
xnor U6542 (N_6542,N_2412,N_3027);
nor U6543 (N_6543,N_687,N_2275);
and U6544 (N_6544,N_1019,N_1041);
and U6545 (N_6545,N_2117,N_1293);
nand U6546 (N_6546,N_1747,N_528);
nand U6547 (N_6547,N_140,N_3710);
and U6548 (N_6548,N_2325,N_3546);
nor U6549 (N_6549,N_3374,N_3018);
or U6550 (N_6550,N_1004,N_1357);
xnor U6551 (N_6551,N_2077,N_1019);
nand U6552 (N_6552,N_889,N_717);
nand U6553 (N_6553,N_1233,N_3137);
nand U6554 (N_6554,N_3433,N_1509);
or U6555 (N_6555,N_2296,N_1391);
or U6556 (N_6556,N_2777,N_3663);
nand U6557 (N_6557,N_1245,N_671);
xnor U6558 (N_6558,N_2283,N_137);
nor U6559 (N_6559,N_1609,N_535);
or U6560 (N_6560,N_2663,N_3286);
xor U6561 (N_6561,N_276,N_621);
or U6562 (N_6562,N_1531,N_552);
and U6563 (N_6563,N_3523,N_3079);
or U6564 (N_6564,N_81,N_1055);
xnor U6565 (N_6565,N_2060,N_2334);
nand U6566 (N_6566,N_376,N_1854);
or U6567 (N_6567,N_2755,N_1149);
xor U6568 (N_6568,N_523,N_532);
xnor U6569 (N_6569,N_930,N_176);
xnor U6570 (N_6570,N_12,N_500);
nor U6571 (N_6571,N_1294,N_3251);
and U6572 (N_6572,N_3184,N_2799);
nor U6573 (N_6573,N_1746,N_2408);
or U6574 (N_6574,N_1309,N_1715);
or U6575 (N_6575,N_3786,N_2678);
nand U6576 (N_6576,N_582,N_3848);
or U6577 (N_6577,N_447,N_3349);
and U6578 (N_6578,N_2688,N_2654);
xor U6579 (N_6579,N_72,N_1736);
or U6580 (N_6580,N_251,N_608);
nor U6581 (N_6581,N_3515,N_1231);
xnor U6582 (N_6582,N_1449,N_46);
nand U6583 (N_6583,N_3559,N_1733);
nand U6584 (N_6584,N_1311,N_3154);
or U6585 (N_6585,N_2319,N_2065);
nor U6586 (N_6586,N_2658,N_2061);
or U6587 (N_6587,N_2963,N_1944);
or U6588 (N_6588,N_3035,N_3040);
nand U6589 (N_6589,N_1879,N_1220);
or U6590 (N_6590,N_2358,N_152);
or U6591 (N_6591,N_1012,N_2640);
and U6592 (N_6592,N_1911,N_3210);
nor U6593 (N_6593,N_1065,N_2916);
xnor U6594 (N_6594,N_217,N_2388);
nor U6595 (N_6595,N_1174,N_2679);
nor U6596 (N_6596,N_3548,N_3813);
nor U6597 (N_6597,N_1213,N_3054);
xnor U6598 (N_6598,N_1771,N_3142);
nand U6599 (N_6599,N_2365,N_2268);
nand U6600 (N_6600,N_1360,N_2131);
or U6601 (N_6601,N_3790,N_87);
and U6602 (N_6602,N_476,N_3359);
and U6603 (N_6603,N_1446,N_2308);
or U6604 (N_6604,N_689,N_730);
nor U6605 (N_6605,N_3182,N_1027);
xor U6606 (N_6606,N_3480,N_1182);
or U6607 (N_6607,N_2209,N_1336);
xnor U6608 (N_6608,N_1491,N_498);
nand U6609 (N_6609,N_3001,N_3732);
xnor U6610 (N_6610,N_3079,N_1793);
and U6611 (N_6611,N_3536,N_2066);
nand U6612 (N_6612,N_1039,N_1106);
or U6613 (N_6613,N_2025,N_408);
or U6614 (N_6614,N_2213,N_554);
or U6615 (N_6615,N_2267,N_3353);
xnor U6616 (N_6616,N_2896,N_3841);
nand U6617 (N_6617,N_295,N_3648);
nor U6618 (N_6618,N_230,N_3924);
or U6619 (N_6619,N_750,N_1786);
and U6620 (N_6620,N_566,N_697);
xnor U6621 (N_6621,N_730,N_480);
nor U6622 (N_6622,N_3779,N_2704);
or U6623 (N_6623,N_1190,N_3149);
or U6624 (N_6624,N_3276,N_1111);
and U6625 (N_6625,N_1356,N_2248);
xnor U6626 (N_6626,N_1002,N_1996);
or U6627 (N_6627,N_3351,N_126);
and U6628 (N_6628,N_3198,N_1827);
or U6629 (N_6629,N_2813,N_2451);
nand U6630 (N_6630,N_3114,N_2697);
or U6631 (N_6631,N_2647,N_1675);
nor U6632 (N_6632,N_688,N_3055);
nand U6633 (N_6633,N_3353,N_3955);
or U6634 (N_6634,N_1959,N_61);
and U6635 (N_6635,N_2478,N_910);
and U6636 (N_6636,N_1648,N_255);
nor U6637 (N_6637,N_3313,N_1113);
nand U6638 (N_6638,N_38,N_988);
nand U6639 (N_6639,N_1672,N_467);
xor U6640 (N_6640,N_3497,N_650);
nor U6641 (N_6641,N_3572,N_1456);
nand U6642 (N_6642,N_1500,N_2620);
and U6643 (N_6643,N_401,N_1471);
or U6644 (N_6644,N_3684,N_549);
nand U6645 (N_6645,N_1361,N_3678);
xor U6646 (N_6646,N_3368,N_1942);
nor U6647 (N_6647,N_3710,N_2826);
xor U6648 (N_6648,N_2975,N_325);
or U6649 (N_6649,N_2393,N_1174);
nand U6650 (N_6650,N_329,N_1753);
nand U6651 (N_6651,N_1327,N_737);
xor U6652 (N_6652,N_584,N_1225);
or U6653 (N_6653,N_3,N_2820);
nand U6654 (N_6654,N_3583,N_831);
and U6655 (N_6655,N_3082,N_2122);
or U6656 (N_6656,N_2613,N_1268);
and U6657 (N_6657,N_1180,N_3558);
nand U6658 (N_6658,N_139,N_175);
nor U6659 (N_6659,N_467,N_217);
xnor U6660 (N_6660,N_1799,N_1913);
or U6661 (N_6661,N_3355,N_1135);
nand U6662 (N_6662,N_1322,N_1976);
nand U6663 (N_6663,N_3870,N_2211);
or U6664 (N_6664,N_1732,N_2546);
and U6665 (N_6665,N_1003,N_96);
or U6666 (N_6666,N_3939,N_564);
xnor U6667 (N_6667,N_809,N_1642);
and U6668 (N_6668,N_2871,N_2798);
or U6669 (N_6669,N_134,N_2802);
nand U6670 (N_6670,N_2665,N_3828);
or U6671 (N_6671,N_702,N_3690);
nor U6672 (N_6672,N_2380,N_3032);
or U6673 (N_6673,N_2737,N_1696);
nand U6674 (N_6674,N_2575,N_1729);
and U6675 (N_6675,N_812,N_3767);
or U6676 (N_6676,N_565,N_2815);
nor U6677 (N_6677,N_2018,N_308);
nor U6678 (N_6678,N_1372,N_156);
or U6679 (N_6679,N_1566,N_2846);
or U6680 (N_6680,N_962,N_3117);
nand U6681 (N_6681,N_1684,N_2338);
or U6682 (N_6682,N_2994,N_3082);
and U6683 (N_6683,N_1030,N_3839);
xnor U6684 (N_6684,N_1484,N_188);
xor U6685 (N_6685,N_3213,N_1561);
or U6686 (N_6686,N_2909,N_2357);
and U6687 (N_6687,N_1416,N_681);
nand U6688 (N_6688,N_757,N_321);
nor U6689 (N_6689,N_384,N_1474);
nand U6690 (N_6690,N_3815,N_1773);
xor U6691 (N_6691,N_5,N_2370);
xor U6692 (N_6692,N_1757,N_532);
and U6693 (N_6693,N_967,N_3889);
nor U6694 (N_6694,N_1597,N_2607);
and U6695 (N_6695,N_3565,N_2484);
and U6696 (N_6696,N_2913,N_765);
and U6697 (N_6697,N_470,N_2517);
nor U6698 (N_6698,N_359,N_1198);
nand U6699 (N_6699,N_3324,N_2740);
xnor U6700 (N_6700,N_3958,N_2674);
nor U6701 (N_6701,N_824,N_3667);
nor U6702 (N_6702,N_3380,N_2922);
nand U6703 (N_6703,N_1550,N_1466);
and U6704 (N_6704,N_2249,N_2504);
nor U6705 (N_6705,N_2715,N_1761);
and U6706 (N_6706,N_1696,N_1794);
nand U6707 (N_6707,N_84,N_3230);
xor U6708 (N_6708,N_198,N_3502);
or U6709 (N_6709,N_738,N_1430);
and U6710 (N_6710,N_1954,N_3637);
nand U6711 (N_6711,N_3862,N_1500);
xnor U6712 (N_6712,N_3127,N_83);
or U6713 (N_6713,N_969,N_3192);
and U6714 (N_6714,N_3282,N_919);
nor U6715 (N_6715,N_170,N_1627);
or U6716 (N_6716,N_99,N_3391);
nand U6717 (N_6717,N_44,N_1138);
nand U6718 (N_6718,N_1013,N_1382);
nor U6719 (N_6719,N_3337,N_3303);
nand U6720 (N_6720,N_2005,N_1877);
nand U6721 (N_6721,N_2429,N_547);
nand U6722 (N_6722,N_534,N_2708);
nor U6723 (N_6723,N_3136,N_2691);
nand U6724 (N_6724,N_1366,N_485);
or U6725 (N_6725,N_1270,N_1893);
and U6726 (N_6726,N_2252,N_3838);
nor U6727 (N_6727,N_376,N_2834);
and U6728 (N_6728,N_1392,N_2539);
and U6729 (N_6729,N_2459,N_2390);
xnor U6730 (N_6730,N_3377,N_3549);
and U6731 (N_6731,N_3686,N_2814);
nor U6732 (N_6732,N_579,N_1024);
nand U6733 (N_6733,N_1515,N_3074);
xor U6734 (N_6734,N_2987,N_97);
and U6735 (N_6735,N_2537,N_2759);
nor U6736 (N_6736,N_1786,N_1560);
or U6737 (N_6737,N_670,N_3840);
or U6738 (N_6738,N_2644,N_134);
nor U6739 (N_6739,N_3784,N_493);
or U6740 (N_6740,N_2018,N_846);
nand U6741 (N_6741,N_798,N_3052);
nor U6742 (N_6742,N_1886,N_2889);
or U6743 (N_6743,N_3674,N_2794);
nor U6744 (N_6744,N_3241,N_2992);
or U6745 (N_6745,N_1457,N_2653);
and U6746 (N_6746,N_3994,N_3923);
xor U6747 (N_6747,N_2427,N_904);
nand U6748 (N_6748,N_3926,N_958);
nor U6749 (N_6749,N_1619,N_1627);
and U6750 (N_6750,N_3667,N_2320);
or U6751 (N_6751,N_1909,N_605);
or U6752 (N_6752,N_1002,N_3203);
nand U6753 (N_6753,N_3551,N_2049);
xor U6754 (N_6754,N_13,N_3517);
and U6755 (N_6755,N_545,N_614);
nand U6756 (N_6756,N_1135,N_2914);
nor U6757 (N_6757,N_3172,N_1609);
nand U6758 (N_6758,N_1477,N_240);
nor U6759 (N_6759,N_198,N_2067);
nand U6760 (N_6760,N_2414,N_743);
nor U6761 (N_6761,N_2505,N_1823);
nor U6762 (N_6762,N_865,N_3053);
and U6763 (N_6763,N_1263,N_1153);
xnor U6764 (N_6764,N_3573,N_263);
nor U6765 (N_6765,N_2855,N_11);
nand U6766 (N_6766,N_3474,N_1265);
nand U6767 (N_6767,N_233,N_2279);
nand U6768 (N_6768,N_1110,N_974);
xor U6769 (N_6769,N_623,N_3948);
nand U6770 (N_6770,N_3266,N_901);
xnor U6771 (N_6771,N_1708,N_694);
and U6772 (N_6772,N_2892,N_253);
nor U6773 (N_6773,N_3781,N_49);
xnor U6774 (N_6774,N_3396,N_1599);
and U6775 (N_6775,N_3321,N_2832);
and U6776 (N_6776,N_672,N_3862);
xor U6777 (N_6777,N_3862,N_2764);
nand U6778 (N_6778,N_642,N_2944);
nor U6779 (N_6779,N_3120,N_2085);
nand U6780 (N_6780,N_936,N_383);
nor U6781 (N_6781,N_336,N_939);
nand U6782 (N_6782,N_1394,N_286);
nor U6783 (N_6783,N_2577,N_1244);
nand U6784 (N_6784,N_3605,N_2194);
nand U6785 (N_6785,N_2852,N_2326);
and U6786 (N_6786,N_1937,N_3078);
nor U6787 (N_6787,N_408,N_245);
nand U6788 (N_6788,N_2037,N_949);
or U6789 (N_6789,N_371,N_88);
nor U6790 (N_6790,N_3935,N_140);
and U6791 (N_6791,N_273,N_3181);
nor U6792 (N_6792,N_2177,N_3978);
or U6793 (N_6793,N_2137,N_298);
and U6794 (N_6794,N_1923,N_1473);
and U6795 (N_6795,N_1907,N_1218);
or U6796 (N_6796,N_3297,N_1939);
nor U6797 (N_6797,N_36,N_2249);
xnor U6798 (N_6798,N_1820,N_1589);
and U6799 (N_6799,N_330,N_1805);
and U6800 (N_6800,N_2867,N_783);
nand U6801 (N_6801,N_1704,N_2398);
and U6802 (N_6802,N_1083,N_1530);
or U6803 (N_6803,N_2497,N_3590);
xor U6804 (N_6804,N_3148,N_2972);
nor U6805 (N_6805,N_2329,N_3751);
nand U6806 (N_6806,N_1941,N_109);
or U6807 (N_6807,N_1389,N_3172);
nor U6808 (N_6808,N_156,N_2446);
or U6809 (N_6809,N_1349,N_3062);
and U6810 (N_6810,N_3077,N_516);
or U6811 (N_6811,N_3156,N_3181);
and U6812 (N_6812,N_3977,N_3447);
nand U6813 (N_6813,N_3752,N_1792);
and U6814 (N_6814,N_3511,N_371);
nand U6815 (N_6815,N_647,N_3724);
nor U6816 (N_6816,N_570,N_3269);
nand U6817 (N_6817,N_3176,N_1913);
xnor U6818 (N_6818,N_1568,N_1169);
and U6819 (N_6819,N_1061,N_552);
xor U6820 (N_6820,N_3906,N_3888);
and U6821 (N_6821,N_1656,N_1278);
nand U6822 (N_6822,N_1200,N_1668);
xor U6823 (N_6823,N_2124,N_2149);
or U6824 (N_6824,N_250,N_3392);
nor U6825 (N_6825,N_754,N_1921);
xor U6826 (N_6826,N_1157,N_2394);
nand U6827 (N_6827,N_2279,N_2293);
nor U6828 (N_6828,N_3249,N_979);
nand U6829 (N_6829,N_1743,N_48);
and U6830 (N_6830,N_1431,N_1757);
nand U6831 (N_6831,N_457,N_2282);
nor U6832 (N_6832,N_3485,N_1999);
and U6833 (N_6833,N_3396,N_667);
nand U6834 (N_6834,N_2231,N_2355);
nor U6835 (N_6835,N_1880,N_222);
nor U6836 (N_6836,N_696,N_1177);
xnor U6837 (N_6837,N_3945,N_3196);
or U6838 (N_6838,N_3065,N_1051);
and U6839 (N_6839,N_1110,N_1313);
nand U6840 (N_6840,N_1903,N_466);
and U6841 (N_6841,N_3449,N_815);
and U6842 (N_6842,N_2709,N_1624);
or U6843 (N_6843,N_3352,N_3255);
nand U6844 (N_6844,N_2490,N_2771);
nand U6845 (N_6845,N_3031,N_301);
or U6846 (N_6846,N_1284,N_1673);
and U6847 (N_6847,N_3005,N_847);
or U6848 (N_6848,N_2752,N_3898);
and U6849 (N_6849,N_1138,N_1040);
and U6850 (N_6850,N_885,N_3941);
nand U6851 (N_6851,N_2810,N_3936);
and U6852 (N_6852,N_19,N_865);
nor U6853 (N_6853,N_358,N_598);
or U6854 (N_6854,N_939,N_1160);
and U6855 (N_6855,N_2253,N_2318);
and U6856 (N_6856,N_687,N_612);
xor U6857 (N_6857,N_3456,N_550);
nor U6858 (N_6858,N_1899,N_2129);
nor U6859 (N_6859,N_2892,N_3602);
or U6860 (N_6860,N_527,N_1913);
or U6861 (N_6861,N_3215,N_3210);
nor U6862 (N_6862,N_232,N_2655);
nand U6863 (N_6863,N_2624,N_2247);
or U6864 (N_6864,N_100,N_2569);
or U6865 (N_6865,N_329,N_953);
nor U6866 (N_6866,N_2,N_2681);
xor U6867 (N_6867,N_1858,N_2862);
xnor U6868 (N_6868,N_3226,N_350);
nor U6869 (N_6869,N_3922,N_2549);
xnor U6870 (N_6870,N_3229,N_19);
xor U6871 (N_6871,N_1578,N_3784);
or U6872 (N_6872,N_1976,N_2346);
xor U6873 (N_6873,N_2289,N_3676);
or U6874 (N_6874,N_3556,N_2833);
and U6875 (N_6875,N_2215,N_3092);
or U6876 (N_6876,N_2180,N_3882);
xor U6877 (N_6877,N_2023,N_1217);
nor U6878 (N_6878,N_3999,N_3041);
nand U6879 (N_6879,N_834,N_3190);
or U6880 (N_6880,N_2693,N_3255);
nand U6881 (N_6881,N_2360,N_3121);
and U6882 (N_6882,N_3932,N_2256);
nor U6883 (N_6883,N_2226,N_1448);
and U6884 (N_6884,N_1029,N_1994);
and U6885 (N_6885,N_1736,N_3129);
and U6886 (N_6886,N_3138,N_858);
xor U6887 (N_6887,N_1551,N_847);
nand U6888 (N_6888,N_2242,N_3219);
and U6889 (N_6889,N_3311,N_2585);
nor U6890 (N_6890,N_3770,N_2184);
and U6891 (N_6891,N_3550,N_2761);
or U6892 (N_6892,N_3553,N_1327);
nand U6893 (N_6893,N_3935,N_478);
xor U6894 (N_6894,N_1503,N_2169);
nor U6895 (N_6895,N_1327,N_3044);
nand U6896 (N_6896,N_848,N_3116);
or U6897 (N_6897,N_317,N_1831);
nand U6898 (N_6898,N_3964,N_3144);
nor U6899 (N_6899,N_1185,N_3876);
xnor U6900 (N_6900,N_628,N_1986);
nand U6901 (N_6901,N_3354,N_393);
xor U6902 (N_6902,N_3427,N_2419);
and U6903 (N_6903,N_3108,N_177);
or U6904 (N_6904,N_1462,N_3229);
xor U6905 (N_6905,N_874,N_222);
nand U6906 (N_6906,N_2735,N_1548);
nand U6907 (N_6907,N_719,N_2748);
xnor U6908 (N_6908,N_3417,N_880);
nand U6909 (N_6909,N_2362,N_3572);
xor U6910 (N_6910,N_2657,N_811);
xor U6911 (N_6911,N_2340,N_2974);
xor U6912 (N_6912,N_2180,N_572);
and U6913 (N_6913,N_1403,N_1740);
nand U6914 (N_6914,N_2281,N_473);
or U6915 (N_6915,N_2928,N_2503);
and U6916 (N_6916,N_981,N_2351);
xnor U6917 (N_6917,N_3561,N_3020);
and U6918 (N_6918,N_3071,N_1930);
and U6919 (N_6919,N_1078,N_3123);
nor U6920 (N_6920,N_314,N_1083);
nor U6921 (N_6921,N_1263,N_904);
xor U6922 (N_6922,N_3825,N_488);
xnor U6923 (N_6923,N_1055,N_315);
and U6924 (N_6924,N_2205,N_412);
xnor U6925 (N_6925,N_2906,N_338);
and U6926 (N_6926,N_2540,N_557);
and U6927 (N_6927,N_686,N_3554);
nor U6928 (N_6928,N_560,N_1414);
nor U6929 (N_6929,N_2977,N_1421);
or U6930 (N_6930,N_1227,N_930);
and U6931 (N_6931,N_562,N_1859);
or U6932 (N_6932,N_654,N_3131);
and U6933 (N_6933,N_1827,N_596);
and U6934 (N_6934,N_3446,N_2375);
nor U6935 (N_6935,N_3539,N_2674);
nor U6936 (N_6936,N_1735,N_1221);
or U6937 (N_6937,N_3616,N_1547);
xor U6938 (N_6938,N_884,N_2804);
nor U6939 (N_6939,N_3195,N_2077);
nor U6940 (N_6940,N_2533,N_2934);
or U6941 (N_6941,N_3255,N_3565);
nor U6942 (N_6942,N_3996,N_1452);
nand U6943 (N_6943,N_3220,N_3929);
or U6944 (N_6944,N_597,N_1238);
xnor U6945 (N_6945,N_2230,N_3052);
xor U6946 (N_6946,N_2492,N_156);
and U6947 (N_6947,N_3987,N_758);
nor U6948 (N_6948,N_1551,N_1273);
nand U6949 (N_6949,N_2700,N_1547);
nand U6950 (N_6950,N_3692,N_1449);
xor U6951 (N_6951,N_2967,N_3063);
nor U6952 (N_6952,N_2712,N_2632);
and U6953 (N_6953,N_1600,N_2781);
nand U6954 (N_6954,N_431,N_3611);
nor U6955 (N_6955,N_2921,N_1931);
or U6956 (N_6956,N_1755,N_3393);
or U6957 (N_6957,N_88,N_3825);
xnor U6958 (N_6958,N_2174,N_2857);
nor U6959 (N_6959,N_1598,N_3029);
nor U6960 (N_6960,N_1367,N_461);
nand U6961 (N_6961,N_1790,N_1384);
or U6962 (N_6962,N_869,N_3986);
xor U6963 (N_6963,N_1848,N_2369);
nor U6964 (N_6964,N_1316,N_3611);
nor U6965 (N_6965,N_3569,N_907);
nor U6966 (N_6966,N_569,N_3830);
nand U6967 (N_6967,N_762,N_1957);
nand U6968 (N_6968,N_1044,N_3709);
nand U6969 (N_6969,N_1525,N_1323);
xnor U6970 (N_6970,N_3868,N_2956);
nand U6971 (N_6971,N_1082,N_819);
xnor U6972 (N_6972,N_3789,N_3460);
nor U6973 (N_6973,N_1949,N_363);
and U6974 (N_6974,N_3986,N_3545);
nor U6975 (N_6975,N_2996,N_1832);
or U6976 (N_6976,N_901,N_3967);
nand U6977 (N_6977,N_3128,N_753);
nor U6978 (N_6978,N_501,N_1689);
xnor U6979 (N_6979,N_1285,N_1526);
nor U6980 (N_6980,N_1707,N_3134);
or U6981 (N_6981,N_3899,N_988);
and U6982 (N_6982,N_3403,N_3901);
nand U6983 (N_6983,N_3434,N_1640);
nand U6984 (N_6984,N_1817,N_1616);
or U6985 (N_6985,N_2254,N_2321);
xnor U6986 (N_6986,N_3114,N_1542);
and U6987 (N_6987,N_1088,N_1528);
or U6988 (N_6988,N_109,N_315);
nand U6989 (N_6989,N_698,N_1726);
xnor U6990 (N_6990,N_3923,N_3765);
or U6991 (N_6991,N_1010,N_2666);
and U6992 (N_6992,N_3502,N_3017);
nand U6993 (N_6993,N_3283,N_844);
and U6994 (N_6994,N_3847,N_2817);
or U6995 (N_6995,N_236,N_343);
nand U6996 (N_6996,N_684,N_1233);
xnor U6997 (N_6997,N_2702,N_1913);
nor U6998 (N_6998,N_1087,N_573);
or U6999 (N_6999,N_2011,N_116);
nor U7000 (N_7000,N_1870,N_3578);
nand U7001 (N_7001,N_2481,N_3636);
nor U7002 (N_7002,N_1070,N_1676);
or U7003 (N_7003,N_670,N_3128);
or U7004 (N_7004,N_3175,N_3270);
or U7005 (N_7005,N_2421,N_2426);
nor U7006 (N_7006,N_906,N_1206);
nand U7007 (N_7007,N_1465,N_1678);
or U7008 (N_7008,N_1790,N_1742);
nand U7009 (N_7009,N_3797,N_388);
xor U7010 (N_7010,N_1072,N_2790);
xnor U7011 (N_7011,N_950,N_3965);
or U7012 (N_7012,N_2745,N_1742);
or U7013 (N_7013,N_3329,N_3156);
xnor U7014 (N_7014,N_334,N_1009);
nand U7015 (N_7015,N_44,N_2842);
and U7016 (N_7016,N_912,N_793);
xor U7017 (N_7017,N_2693,N_2614);
nor U7018 (N_7018,N_2214,N_331);
xor U7019 (N_7019,N_2750,N_1685);
xnor U7020 (N_7020,N_3113,N_3859);
and U7021 (N_7021,N_160,N_2122);
nor U7022 (N_7022,N_3354,N_3632);
xor U7023 (N_7023,N_1272,N_3689);
xor U7024 (N_7024,N_3287,N_1782);
xor U7025 (N_7025,N_825,N_767);
and U7026 (N_7026,N_3466,N_330);
nor U7027 (N_7027,N_3146,N_296);
nor U7028 (N_7028,N_3080,N_2955);
nor U7029 (N_7029,N_3044,N_3549);
and U7030 (N_7030,N_3564,N_694);
nor U7031 (N_7031,N_1828,N_677);
xor U7032 (N_7032,N_3041,N_1840);
nor U7033 (N_7033,N_2154,N_1612);
nand U7034 (N_7034,N_187,N_1416);
and U7035 (N_7035,N_868,N_2035);
or U7036 (N_7036,N_459,N_430);
xor U7037 (N_7037,N_225,N_271);
xnor U7038 (N_7038,N_2706,N_701);
nor U7039 (N_7039,N_3782,N_777);
and U7040 (N_7040,N_686,N_700);
xnor U7041 (N_7041,N_772,N_3263);
nor U7042 (N_7042,N_1895,N_3146);
xor U7043 (N_7043,N_2802,N_938);
and U7044 (N_7044,N_2050,N_1333);
xnor U7045 (N_7045,N_1609,N_2376);
or U7046 (N_7046,N_1432,N_788);
nand U7047 (N_7047,N_1437,N_2670);
nor U7048 (N_7048,N_2560,N_645);
nand U7049 (N_7049,N_699,N_2759);
or U7050 (N_7050,N_103,N_3860);
nor U7051 (N_7051,N_1472,N_3552);
or U7052 (N_7052,N_2208,N_1117);
and U7053 (N_7053,N_1592,N_2776);
xnor U7054 (N_7054,N_2908,N_2903);
nand U7055 (N_7055,N_1859,N_3643);
xor U7056 (N_7056,N_1152,N_873);
or U7057 (N_7057,N_2867,N_3759);
or U7058 (N_7058,N_1750,N_1997);
and U7059 (N_7059,N_586,N_1728);
xnor U7060 (N_7060,N_3051,N_804);
nand U7061 (N_7061,N_3177,N_918);
xor U7062 (N_7062,N_1931,N_888);
xnor U7063 (N_7063,N_2306,N_2474);
xnor U7064 (N_7064,N_732,N_2799);
xor U7065 (N_7065,N_1913,N_2927);
nand U7066 (N_7066,N_2821,N_196);
nor U7067 (N_7067,N_1057,N_580);
and U7068 (N_7068,N_219,N_3342);
and U7069 (N_7069,N_2794,N_1539);
and U7070 (N_7070,N_3700,N_3978);
and U7071 (N_7071,N_317,N_322);
nor U7072 (N_7072,N_2025,N_3748);
or U7073 (N_7073,N_2656,N_162);
nand U7074 (N_7074,N_3173,N_3195);
and U7075 (N_7075,N_2648,N_1215);
and U7076 (N_7076,N_2282,N_253);
xnor U7077 (N_7077,N_1852,N_1280);
or U7078 (N_7078,N_1083,N_2489);
or U7079 (N_7079,N_547,N_1426);
nor U7080 (N_7080,N_1323,N_3486);
or U7081 (N_7081,N_1852,N_3389);
nor U7082 (N_7082,N_3017,N_671);
xor U7083 (N_7083,N_2815,N_3276);
or U7084 (N_7084,N_3698,N_3093);
xnor U7085 (N_7085,N_262,N_1167);
xor U7086 (N_7086,N_2728,N_118);
nand U7087 (N_7087,N_2297,N_643);
or U7088 (N_7088,N_2498,N_3950);
nor U7089 (N_7089,N_3114,N_2522);
and U7090 (N_7090,N_795,N_750);
and U7091 (N_7091,N_3484,N_1423);
or U7092 (N_7092,N_1049,N_147);
xor U7093 (N_7093,N_226,N_2063);
nor U7094 (N_7094,N_1975,N_413);
or U7095 (N_7095,N_3569,N_471);
nor U7096 (N_7096,N_3821,N_2752);
nand U7097 (N_7097,N_3957,N_3165);
and U7098 (N_7098,N_2827,N_2326);
or U7099 (N_7099,N_2782,N_1615);
xor U7100 (N_7100,N_2612,N_3320);
nor U7101 (N_7101,N_85,N_3168);
nor U7102 (N_7102,N_1248,N_2741);
and U7103 (N_7103,N_2478,N_3470);
xor U7104 (N_7104,N_170,N_2707);
nor U7105 (N_7105,N_687,N_2059);
xnor U7106 (N_7106,N_2457,N_1947);
or U7107 (N_7107,N_2537,N_2505);
and U7108 (N_7108,N_554,N_54);
nand U7109 (N_7109,N_949,N_3151);
and U7110 (N_7110,N_2627,N_3100);
or U7111 (N_7111,N_3869,N_1076);
nand U7112 (N_7112,N_437,N_3792);
or U7113 (N_7113,N_1349,N_1211);
or U7114 (N_7114,N_1717,N_1737);
nand U7115 (N_7115,N_1840,N_3556);
and U7116 (N_7116,N_2185,N_3534);
nand U7117 (N_7117,N_3031,N_1148);
and U7118 (N_7118,N_2919,N_3677);
nand U7119 (N_7119,N_158,N_1585);
xor U7120 (N_7120,N_333,N_3174);
and U7121 (N_7121,N_2140,N_139);
and U7122 (N_7122,N_3743,N_2599);
nand U7123 (N_7123,N_3450,N_282);
or U7124 (N_7124,N_3286,N_2139);
nand U7125 (N_7125,N_2990,N_3781);
nor U7126 (N_7126,N_131,N_2109);
or U7127 (N_7127,N_1009,N_1486);
nor U7128 (N_7128,N_1676,N_3699);
and U7129 (N_7129,N_2604,N_121);
nor U7130 (N_7130,N_3764,N_2645);
nand U7131 (N_7131,N_2499,N_3430);
xnor U7132 (N_7132,N_500,N_1596);
or U7133 (N_7133,N_2427,N_3311);
or U7134 (N_7134,N_1145,N_1647);
nand U7135 (N_7135,N_472,N_3335);
or U7136 (N_7136,N_1985,N_2925);
and U7137 (N_7137,N_2051,N_2024);
or U7138 (N_7138,N_3662,N_620);
nor U7139 (N_7139,N_3738,N_2959);
nor U7140 (N_7140,N_1782,N_3885);
or U7141 (N_7141,N_3482,N_559);
and U7142 (N_7142,N_3169,N_2179);
or U7143 (N_7143,N_2086,N_261);
and U7144 (N_7144,N_229,N_1804);
and U7145 (N_7145,N_2449,N_1293);
nand U7146 (N_7146,N_1252,N_2811);
or U7147 (N_7147,N_880,N_633);
or U7148 (N_7148,N_3604,N_3493);
xnor U7149 (N_7149,N_925,N_3845);
or U7150 (N_7150,N_1297,N_545);
or U7151 (N_7151,N_3272,N_3943);
nand U7152 (N_7152,N_2593,N_889);
nor U7153 (N_7153,N_247,N_780);
nor U7154 (N_7154,N_3127,N_554);
or U7155 (N_7155,N_2693,N_3658);
xnor U7156 (N_7156,N_2151,N_3407);
xor U7157 (N_7157,N_3085,N_2412);
nor U7158 (N_7158,N_1762,N_1205);
xor U7159 (N_7159,N_3355,N_2207);
xnor U7160 (N_7160,N_637,N_3242);
nor U7161 (N_7161,N_3852,N_788);
and U7162 (N_7162,N_2840,N_396);
and U7163 (N_7163,N_3272,N_2451);
nor U7164 (N_7164,N_2391,N_1658);
xor U7165 (N_7165,N_2971,N_2912);
nor U7166 (N_7166,N_2551,N_1430);
xnor U7167 (N_7167,N_3765,N_786);
nor U7168 (N_7168,N_517,N_857);
or U7169 (N_7169,N_2436,N_289);
and U7170 (N_7170,N_570,N_1339);
or U7171 (N_7171,N_461,N_761);
and U7172 (N_7172,N_422,N_2797);
and U7173 (N_7173,N_1649,N_757);
xor U7174 (N_7174,N_521,N_3727);
nand U7175 (N_7175,N_1252,N_3815);
xor U7176 (N_7176,N_2166,N_2231);
nor U7177 (N_7177,N_953,N_1820);
or U7178 (N_7178,N_986,N_1454);
nand U7179 (N_7179,N_3048,N_1719);
nor U7180 (N_7180,N_1727,N_607);
xnor U7181 (N_7181,N_2597,N_1742);
or U7182 (N_7182,N_1189,N_305);
nor U7183 (N_7183,N_559,N_2461);
nor U7184 (N_7184,N_3251,N_3131);
nor U7185 (N_7185,N_3562,N_2826);
xor U7186 (N_7186,N_2793,N_3716);
nor U7187 (N_7187,N_3587,N_2398);
or U7188 (N_7188,N_2685,N_3121);
nand U7189 (N_7189,N_3353,N_2939);
xor U7190 (N_7190,N_3480,N_374);
or U7191 (N_7191,N_1051,N_3949);
and U7192 (N_7192,N_2025,N_258);
nor U7193 (N_7193,N_1536,N_79);
nand U7194 (N_7194,N_501,N_3925);
nand U7195 (N_7195,N_2277,N_762);
xor U7196 (N_7196,N_3366,N_802);
and U7197 (N_7197,N_1443,N_1783);
nor U7198 (N_7198,N_934,N_1781);
xor U7199 (N_7199,N_412,N_1158);
nand U7200 (N_7200,N_3837,N_334);
and U7201 (N_7201,N_2404,N_128);
and U7202 (N_7202,N_373,N_3038);
xor U7203 (N_7203,N_3152,N_133);
nor U7204 (N_7204,N_1309,N_588);
nand U7205 (N_7205,N_2560,N_519);
or U7206 (N_7206,N_293,N_3814);
xor U7207 (N_7207,N_2448,N_1434);
or U7208 (N_7208,N_2747,N_712);
xnor U7209 (N_7209,N_1334,N_561);
nor U7210 (N_7210,N_3139,N_2534);
or U7211 (N_7211,N_3244,N_3245);
nand U7212 (N_7212,N_914,N_2333);
or U7213 (N_7213,N_1840,N_3578);
nand U7214 (N_7214,N_2737,N_877);
xnor U7215 (N_7215,N_1392,N_1100);
nand U7216 (N_7216,N_82,N_1446);
nor U7217 (N_7217,N_3842,N_3079);
or U7218 (N_7218,N_1006,N_3433);
xnor U7219 (N_7219,N_1596,N_3886);
and U7220 (N_7220,N_2527,N_704);
and U7221 (N_7221,N_1252,N_1028);
nor U7222 (N_7222,N_2190,N_1940);
nor U7223 (N_7223,N_3021,N_1522);
nor U7224 (N_7224,N_1612,N_233);
nand U7225 (N_7225,N_2837,N_2108);
nor U7226 (N_7226,N_2263,N_2318);
or U7227 (N_7227,N_1791,N_3733);
xnor U7228 (N_7228,N_3030,N_744);
nand U7229 (N_7229,N_31,N_3254);
and U7230 (N_7230,N_3993,N_1032);
or U7231 (N_7231,N_3947,N_2413);
or U7232 (N_7232,N_3088,N_34);
or U7233 (N_7233,N_1262,N_2190);
nand U7234 (N_7234,N_3408,N_3921);
or U7235 (N_7235,N_3509,N_1305);
xor U7236 (N_7236,N_1793,N_2848);
nor U7237 (N_7237,N_3519,N_3598);
or U7238 (N_7238,N_1610,N_2056);
nand U7239 (N_7239,N_3065,N_3094);
xnor U7240 (N_7240,N_3139,N_1019);
and U7241 (N_7241,N_1904,N_3351);
xor U7242 (N_7242,N_1780,N_2331);
nand U7243 (N_7243,N_3856,N_3681);
nand U7244 (N_7244,N_188,N_1117);
xnor U7245 (N_7245,N_2698,N_2580);
and U7246 (N_7246,N_1876,N_97);
xor U7247 (N_7247,N_1300,N_92);
nand U7248 (N_7248,N_674,N_330);
nand U7249 (N_7249,N_3195,N_3798);
xor U7250 (N_7250,N_3197,N_778);
and U7251 (N_7251,N_3460,N_805);
and U7252 (N_7252,N_179,N_2273);
nor U7253 (N_7253,N_3894,N_1900);
and U7254 (N_7254,N_2658,N_314);
or U7255 (N_7255,N_3920,N_1683);
or U7256 (N_7256,N_2782,N_1299);
nand U7257 (N_7257,N_2911,N_3670);
nor U7258 (N_7258,N_1617,N_1652);
nor U7259 (N_7259,N_3192,N_2091);
nor U7260 (N_7260,N_278,N_3265);
or U7261 (N_7261,N_1396,N_2357);
or U7262 (N_7262,N_1204,N_2519);
nand U7263 (N_7263,N_3300,N_1768);
nand U7264 (N_7264,N_2181,N_390);
or U7265 (N_7265,N_3722,N_3114);
nand U7266 (N_7266,N_1993,N_2103);
xor U7267 (N_7267,N_3,N_3049);
xor U7268 (N_7268,N_2394,N_1092);
xnor U7269 (N_7269,N_2203,N_532);
or U7270 (N_7270,N_1740,N_1414);
xnor U7271 (N_7271,N_1160,N_2256);
nand U7272 (N_7272,N_3063,N_2499);
and U7273 (N_7273,N_845,N_1409);
or U7274 (N_7274,N_2548,N_958);
nand U7275 (N_7275,N_3017,N_492);
nand U7276 (N_7276,N_1910,N_2150);
nand U7277 (N_7277,N_2647,N_1964);
or U7278 (N_7278,N_1119,N_3693);
or U7279 (N_7279,N_2731,N_2555);
nor U7280 (N_7280,N_67,N_3515);
nor U7281 (N_7281,N_3544,N_3750);
xor U7282 (N_7282,N_866,N_1241);
xnor U7283 (N_7283,N_662,N_3107);
nand U7284 (N_7284,N_3304,N_1754);
nand U7285 (N_7285,N_1780,N_3325);
and U7286 (N_7286,N_2827,N_2221);
nor U7287 (N_7287,N_1505,N_1782);
nand U7288 (N_7288,N_3330,N_1032);
nor U7289 (N_7289,N_3201,N_2266);
or U7290 (N_7290,N_3080,N_3172);
nand U7291 (N_7291,N_2517,N_407);
xor U7292 (N_7292,N_1842,N_3169);
nand U7293 (N_7293,N_2128,N_1684);
or U7294 (N_7294,N_172,N_2461);
or U7295 (N_7295,N_909,N_2135);
xor U7296 (N_7296,N_1344,N_2853);
or U7297 (N_7297,N_1593,N_643);
or U7298 (N_7298,N_574,N_1231);
or U7299 (N_7299,N_1884,N_444);
nand U7300 (N_7300,N_2866,N_1133);
or U7301 (N_7301,N_2299,N_3670);
nand U7302 (N_7302,N_2762,N_2270);
nor U7303 (N_7303,N_1435,N_1531);
nor U7304 (N_7304,N_2149,N_1335);
xor U7305 (N_7305,N_1893,N_1101);
and U7306 (N_7306,N_1955,N_2297);
nor U7307 (N_7307,N_1479,N_3843);
or U7308 (N_7308,N_2056,N_3692);
nand U7309 (N_7309,N_2238,N_285);
and U7310 (N_7310,N_275,N_2144);
nand U7311 (N_7311,N_586,N_2961);
nor U7312 (N_7312,N_196,N_2178);
or U7313 (N_7313,N_72,N_924);
nand U7314 (N_7314,N_1242,N_3854);
nand U7315 (N_7315,N_3411,N_979);
or U7316 (N_7316,N_2033,N_352);
nand U7317 (N_7317,N_1007,N_3804);
nand U7318 (N_7318,N_3813,N_440);
xnor U7319 (N_7319,N_422,N_1519);
nand U7320 (N_7320,N_2740,N_1944);
nand U7321 (N_7321,N_2065,N_3630);
and U7322 (N_7322,N_1955,N_2701);
xnor U7323 (N_7323,N_1549,N_3365);
or U7324 (N_7324,N_2111,N_3726);
or U7325 (N_7325,N_2508,N_1467);
nand U7326 (N_7326,N_3882,N_2444);
nor U7327 (N_7327,N_3223,N_3813);
nand U7328 (N_7328,N_1361,N_985);
nor U7329 (N_7329,N_2895,N_2598);
xor U7330 (N_7330,N_2680,N_2757);
and U7331 (N_7331,N_3902,N_3206);
nor U7332 (N_7332,N_465,N_1055);
xor U7333 (N_7333,N_3461,N_2072);
xor U7334 (N_7334,N_1971,N_2960);
or U7335 (N_7335,N_2697,N_2155);
xor U7336 (N_7336,N_1104,N_2887);
nor U7337 (N_7337,N_1809,N_325);
nand U7338 (N_7338,N_180,N_3379);
xor U7339 (N_7339,N_3928,N_2284);
xor U7340 (N_7340,N_2586,N_1772);
nand U7341 (N_7341,N_3162,N_712);
nor U7342 (N_7342,N_2541,N_603);
nor U7343 (N_7343,N_2277,N_2098);
or U7344 (N_7344,N_2027,N_2540);
nand U7345 (N_7345,N_2957,N_2264);
nor U7346 (N_7346,N_40,N_763);
or U7347 (N_7347,N_2791,N_69);
nand U7348 (N_7348,N_3893,N_3243);
xnor U7349 (N_7349,N_584,N_1429);
and U7350 (N_7350,N_1134,N_3905);
or U7351 (N_7351,N_2668,N_2994);
nor U7352 (N_7352,N_2214,N_2893);
and U7353 (N_7353,N_1395,N_408);
nand U7354 (N_7354,N_2889,N_3297);
or U7355 (N_7355,N_1809,N_636);
and U7356 (N_7356,N_1912,N_1231);
nor U7357 (N_7357,N_2680,N_3735);
nor U7358 (N_7358,N_2548,N_2266);
or U7359 (N_7359,N_3108,N_3193);
and U7360 (N_7360,N_1909,N_1037);
or U7361 (N_7361,N_135,N_3509);
nor U7362 (N_7362,N_1275,N_126);
nor U7363 (N_7363,N_3598,N_457);
and U7364 (N_7364,N_1302,N_2059);
nor U7365 (N_7365,N_2996,N_2418);
or U7366 (N_7366,N_274,N_3729);
nand U7367 (N_7367,N_3417,N_2197);
nand U7368 (N_7368,N_2787,N_2789);
xor U7369 (N_7369,N_3907,N_3314);
nand U7370 (N_7370,N_3483,N_1104);
and U7371 (N_7371,N_1753,N_2344);
nor U7372 (N_7372,N_2545,N_2709);
and U7373 (N_7373,N_921,N_2719);
nand U7374 (N_7374,N_2801,N_3722);
or U7375 (N_7375,N_2523,N_449);
and U7376 (N_7376,N_3830,N_3887);
or U7377 (N_7377,N_3136,N_3109);
and U7378 (N_7378,N_178,N_1937);
nor U7379 (N_7379,N_3613,N_1756);
and U7380 (N_7380,N_3282,N_1805);
nor U7381 (N_7381,N_3442,N_619);
nand U7382 (N_7382,N_3642,N_3141);
nor U7383 (N_7383,N_2324,N_2898);
or U7384 (N_7384,N_750,N_2010);
nor U7385 (N_7385,N_3215,N_3406);
nor U7386 (N_7386,N_1319,N_1713);
nand U7387 (N_7387,N_3783,N_3054);
xor U7388 (N_7388,N_2810,N_1177);
or U7389 (N_7389,N_2342,N_2116);
xnor U7390 (N_7390,N_2955,N_1454);
nor U7391 (N_7391,N_3879,N_2451);
nor U7392 (N_7392,N_27,N_1286);
xnor U7393 (N_7393,N_2873,N_451);
or U7394 (N_7394,N_1668,N_3999);
nand U7395 (N_7395,N_205,N_866);
nor U7396 (N_7396,N_1533,N_3436);
nand U7397 (N_7397,N_3113,N_3598);
or U7398 (N_7398,N_3728,N_3164);
xor U7399 (N_7399,N_377,N_228);
nor U7400 (N_7400,N_367,N_627);
or U7401 (N_7401,N_1068,N_449);
nor U7402 (N_7402,N_196,N_1393);
xnor U7403 (N_7403,N_1716,N_2574);
xnor U7404 (N_7404,N_728,N_3031);
or U7405 (N_7405,N_3731,N_1949);
and U7406 (N_7406,N_507,N_3633);
and U7407 (N_7407,N_3582,N_1037);
or U7408 (N_7408,N_505,N_2482);
xor U7409 (N_7409,N_984,N_2837);
or U7410 (N_7410,N_3032,N_229);
and U7411 (N_7411,N_2608,N_3542);
nand U7412 (N_7412,N_3954,N_1844);
xor U7413 (N_7413,N_573,N_1189);
and U7414 (N_7414,N_3532,N_2029);
nand U7415 (N_7415,N_1888,N_1936);
xnor U7416 (N_7416,N_1175,N_618);
nor U7417 (N_7417,N_1217,N_263);
nand U7418 (N_7418,N_3671,N_356);
or U7419 (N_7419,N_1633,N_2630);
and U7420 (N_7420,N_1957,N_711);
xnor U7421 (N_7421,N_838,N_2451);
nand U7422 (N_7422,N_1320,N_2711);
and U7423 (N_7423,N_2721,N_547);
nand U7424 (N_7424,N_3321,N_1880);
or U7425 (N_7425,N_298,N_1247);
nor U7426 (N_7426,N_1314,N_1384);
nand U7427 (N_7427,N_2468,N_349);
and U7428 (N_7428,N_3967,N_31);
or U7429 (N_7429,N_3336,N_1707);
or U7430 (N_7430,N_838,N_2005);
xor U7431 (N_7431,N_3191,N_3853);
or U7432 (N_7432,N_2568,N_2574);
or U7433 (N_7433,N_2026,N_3718);
or U7434 (N_7434,N_593,N_3683);
or U7435 (N_7435,N_515,N_740);
nor U7436 (N_7436,N_2885,N_199);
nor U7437 (N_7437,N_2084,N_3803);
and U7438 (N_7438,N_1875,N_1389);
and U7439 (N_7439,N_32,N_1873);
or U7440 (N_7440,N_765,N_3720);
and U7441 (N_7441,N_3379,N_2383);
nor U7442 (N_7442,N_3561,N_2982);
nand U7443 (N_7443,N_2031,N_3024);
xnor U7444 (N_7444,N_2330,N_1844);
nand U7445 (N_7445,N_811,N_1286);
nand U7446 (N_7446,N_1798,N_256);
xnor U7447 (N_7447,N_1395,N_1096);
and U7448 (N_7448,N_266,N_3564);
nor U7449 (N_7449,N_1439,N_3280);
nor U7450 (N_7450,N_1227,N_793);
xnor U7451 (N_7451,N_417,N_2222);
or U7452 (N_7452,N_3126,N_1240);
and U7453 (N_7453,N_2237,N_744);
nor U7454 (N_7454,N_2210,N_2974);
nand U7455 (N_7455,N_3851,N_2338);
nor U7456 (N_7456,N_2611,N_2579);
xor U7457 (N_7457,N_2173,N_1264);
and U7458 (N_7458,N_1714,N_636);
xnor U7459 (N_7459,N_2703,N_1554);
and U7460 (N_7460,N_2013,N_1231);
or U7461 (N_7461,N_2677,N_2310);
xnor U7462 (N_7462,N_3591,N_2793);
and U7463 (N_7463,N_181,N_1210);
xnor U7464 (N_7464,N_2587,N_2444);
and U7465 (N_7465,N_2100,N_2909);
or U7466 (N_7466,N_1967,N_3505);
xnor U7467 (N_7467,N_2549,N_2708);
or U7468 (N_7468,N_3675,N_3658);
or U7469 (N_7469,N_3002,N_1897);
xnor U7470 (N_7470,N_2000,N_215);
xnor U7471 (N_7471,N_1755,N_784);
or U7472 (N_7472,N_3473,N_572);
nand U7473 (N_7473,N_3485,N_3746);
nor U7474 (N_7474,N_2488,N_2831);
and U7475 (N_7475,N_2864,N_2236);
and U7476 (N_7476,N_3591,N_2116);
xnor U7477 (N_7477,N_1311,N_487);
nor U7478 (N_7478,N_2093,N_724);
and U7479 (N_7479,N_3338,N_1255);
nor U7480 (N_7480,N_3842,N_2208);
nand U7481 (N_7481,N_1097,N_1251);
nand U7482 (N_7482,N_2363,N_962);
nand U7483 (N_7483,N_939,N_2070);
and U7484 (N_7484,N_2653,N_3182);
and U7485 (N_7485,N_358,N_124);
or U7486 (N_7486,N_1475,N_1314);
nor U7487 (N_7487,N_1710,N_2421);
xnor U7488 (N_7488,N_863,N_988);
xnor U7489 (N_7489,N_1802,N_1520);
or U7490 (N_7490,N_1012,N_2204);
and U7491 (N_7491,N_2717,N_3981);
and U7492 (N_7492,N_1392,N_1632);
xor U7493 (N_7493,N_3320,N_2126);
and U7494 (N_7494,N_772,N_3319);
xor U7495 (N_7495,N_2971,N_1825);
nor U7496 (N_7496,N_1963,N_262);
xnor U7497 (N_7497,N_325,N_3625);
nand U7498 (N_7498,N_3664,N_2524);
nand U7499 (N_7499,N_1807,N_276);
nand U7500 (N_7500,N_3145,N_3848);
xor U7501 (N_7501,N_1403,N_3832);
and U7502 (N_7502,N_834,N_901);
and U7503 (N_7503,N_82,N_2509);
and U7504 (N_7504,N_1255,N_3837);
xnor U7505 (N_7505,N_2873,N_2742);
nor U7506 (N_7506,N_194,N_173);
xor U7507 (N_7507,N_54,N_3158);
nor U7508 (N_7508,N_1957,N_2737);
nor U7509 (N_7509,N_3525,N_2496);
and U7510 (N_7510,N_126,N_1474);
or U7511 (N_7511,N_1749,N_812);
or U7512 (N_7512,N_271,N_3961);
xor U7513 (N_7513,N_265,N_139);
and U7514 (N_7514,N_1753,N_357);
xnor U7515 (N_7515,N_3938,N_1104);
and U7516 (N_7516,N_846,N_1844);
xnor U7517 (N_7517,N_184,N_3928);
nand U7518 (N_7518,N_3534,N_1615);
nor U7519 (N_7519,N_1486,N_2028);
or U7520 (N_7520,N_754,N_1754);
and U7521 (N_7521,N_3398,N_738);
xor U7522 (N_7522,N_2086,N_2699);
or U7523 (N_7523,N_1715,N_3586);
nand U7524 (N_7524,N_2116,N_3584);
and U7525 (N_7525,N_3191,N_849);
xnor U7526 (N_7526,N_572,N_3588);
xor U7527 (N_7527,N_2512,N_2788);
xnor U7528 (N_7528,N_240,N_132);
or U7529 (N_7529,N_3540,N_2773);
and U7530 (N_7530,N_3405,N_3313);
xnor U7531 (N_7531,N_2545,N_3418);
and U7532 (N_7532,N_682,N_2754);
nor U7533 (N_7533,N_35,N_729);
nand U7534 (N_7534,N_2384,N_743);
nand U7535 (N_7535,N_605,N_538);
or U7536 (N_7536,N_1432,N_3714);
xor U7537 (N_7537,N_218,N_3852);
nor U7538 (N_7538,N_82,N_2728);
xnor U7539 (N_7539,N_1148,N_3273);
or U7540 (N_7540,N_1690,N_537);
or U7541 (N_7541,N_1303,N_1472);
xor U7542 (N_7542,N_2029,N_1207);
nor U7543 (N_7543,N_3949,N_3977);
xnor U7544 (N_7544,N_3375,N_3036);
nand U7545 (N_7545,N_1938,N_3762);
xnor U7546 (N_7546,N_422,N_1972);
or U7547 (N_7547,N_3072,N_221);
and U7548 (N_7548,N_3651,N_375);
xor U7549 (N_7549,N_1716,N_3287);
or U7550 (N_7550,N_1552,N_1155);
nor U7551 (N_7551,N_1287,N_1122);
and U7552 (N_7552,N_1819,N_450);
or U7553 (N_7553,N_741,N_3933);
nor U7554 (N_7554,N_3119,N_95);
or U7555 (N_7555,N_3411,N_915);
and U7556 (N_7556,N_2641,N_321);
nand U7557 (N_7557,N_3285,N_1345);
nand U7558 (N_7558,N_1398,N_2923);
nor U7559 (N_7559,N_955,N_1915);
or U7560 (N_7560,N_3748,N_704);
nand U7561 (N_7561,N_3755,N_2959);
nor U7562 (N_7562,N_1746,N_1516);
nor U7563 (N_7563,N_1053,N_1675);
or U7564 (N_7564,N_1160,N_1461);
and U7565 (N_7565,N_3481,N_2897);
nand U7566 (N_7566,N_1532,N_94);
nand U7567 (N_7567,N_1084,N_480);
or U7568 (N_7568,N_1015,N_3129);
nand U7569 (N_7569,N_77,N_553);
nor U7570 (N_7570,N_2855,N_1915);
nand U7571 (N_7571,N_1760,N_1847);
or U7572 (N_7572,N_3142,N_2091);
and U7573 (N_7573,N_2942,N_3798);
xnor U7574 (N_7574,N_2243,N_1390);
xor U7575 (N_7575,N_2822,N_535);
and U7576 (N_7576,N_3247,N_841);
or U7577 (N_7577,N_2662,N_3697);
or U7578 (N_7578,N_2649,N_3316);
xnor U7579 (N_7579,N_811,N_123);
xnor U7580 (N_7580,N_1276,N_495);
xnor U7581 (N_7581,N_3131,N_1048);
nor U7582 (N_7582,N_3804,N_2601);
or U7583 (N_7583,N_3607,N_2111);
xnor U7584 (N_7584,N_3404,N_2483);
xnor U7585 (N_7585,N_2394,N_1845);
or U7586 (N_7586,N_3326,N_1371);
nor U7587 (N_7587,N_2856,N_902);
xnor U7588 (N_7588,N_3829,N_3260);
and U7589 (N_7589,N_3911,N_105);
or U7590 (N_7590,N_2326,N_1356);
xor U7591 (N_7591,N_77,N_278);
and U7592 (N_7592,N_3127,N_3459);
nor U7593 (N_7593,N_2803,N_959);
or U7594 (N_7594,N_2926,N_2054);
nand U7595 (N_7595,N_211,N_2985);
xnor U7596 (N_7596,N_845,N_2485);
nor U7597 (N_7597,N_858,N_2805);
or U7598 (N_7598,N_1785,N_1481);
nand U7599 (N_7599,N_1117,N_3933);
and U7600 (N_7600,N_2968,N_3189);
nor U7601 (N_7601,N_1645,N_338);
nor U7602 (N_7602,N_829,N_843);
or U7603 (N_7603,N_1267,N_1839);
and U7604 (N_7604,N_575,N_3622);
and U7605 (N_7605,N_3030,N_2089);
nor U7606 (N_7606,N_2736,N_3747);
and U7607 (N_7607,N_3062,N_2254);
or U7608 (N_7608,N_2556,N_3213);
nor U7609 (N_7609,N_2671,N_3233);
nand U7610 (N_7610,N_3915,N_3363);
or U7611 (N_7611,N_1441,N_2537);
or U7612 (N_7612,N_2593,N_3449);
and U7613 (N_7613,N_3117,N_3134);
nor U7614 (N_7614,N_456,N_921);
xor U7615 (N_7615,N_3800,N_2224);
nand U7616 (N_7616,N_3611,N_3679);
and U7617 (N_7617,N_2011,N_2043);
xor U7618 (N_7618,N_279,N_2491);
or U7619 (N_7619,N_2917,N_2037);
nand U7620 (N_7620,N_2050,N_3156);
or U7621 (N_7621,N_1645,N_2631);
or U7622 (N_7622,N_932,N_39);
nand U7623 (N_7623,N_3057,N_2316);
and U7624 (N_7624,N_3617,N_513);
nor U7625 (N_7625,N_828,N_375);
nor U7626 (N_7626,N_1330,N_1124);
nor U7627 (N_7627,N_45,N_3097);
xor U7628 (N_7628,N_3109,N_977);
and U7629 (N_7629,N_2505,N_1365);
xnor U7630 (N_7630,N_1081,N_2483);
nor U7631 (N_7631,N_1663,N_2901);
nor U7632 (N_7632,N_1794,N_643);
nor U7633 (N_7633,N_298,N_3857);
nor U7634 (N_7634,N_1033,N_479);
xnor U7635 (N_7635,N_3065,N_1541);
and U7636 (N_7636,N_3876,N_702);
xor U7637 (N_7637,N_3148,N_516);
or U7638 (N_7638,N_1859,N_2142);
and U7639 (N_7639,N_404,N_1004);
and U7640 (N_7640,N_1567,N_1715);
nand U7641 (N_7641,N_2363,N_2932);
and U7642 (N_7642,N_2221,N_1490);
nand U7643 (N_7643,N_3766,N_3747);
nor U7644 (N_7644,N_827,N_1179);
nor U7645 (N_7645,N_1928,N_1263);
or U7646 (N_7646,N_246,N_3398);
and U7647 (N_7647,N_1029,N_767);
xor U7648 (N_7648,N_2682,N_530);
and U7649 (N_7649,N_1995,N_712);
xor U7650 (N_7650,N_2299,N_2520);
nand U7651 (N_7651,N_1494,N_2916);
nor U7652 (N_7652,N_3092,N_1328);
and U7653 (N_7653,N_2073,N_3459);
nand U7654 (N_7654,N_3065,N_2892);
nor U7655 (N_7655,N_3471,N_214);
xnor U7656 (N_7656,N_1033,N_2780);
nand U7657 (N_7657,N_2106,N_768);
nand U7658 (N_7658,N_2556,N_1984);
nand U7659 (N_7659,N_2768,N_2316);
or U7660 (N_7660,N_645,N_1079);
and U7661 (N_7661,N_3349,N_2400);
and U7662 (N_7662,N_2301,N_1778);
xor U7663 (N_7663,N_3717,N_829);
and U7664 (N_7664,N_2475,N_2964);
or U7665 (N_7665,N_949,N_2524);
or U7666 (N_7666,N_898,N_753);
nor U7667 (N_7667,N_3036,N_732);
nor U7668 (N_7668,N_66,N_3272);
nand U7669 (N_7669,N_247,N_1931);
nand U7670 (N_7670,N_1682,N_3602);
nand U7671 (N_7671,N_2141,N_3077);
or U7672 (N_7672,N_26,N_2435);
nor U7673 (N_7673,N_1800,N_2448);
and U7674 (N_7674,N_1438,N_522);
or U7675 (N_7675,N_2131,N_649);
xnor U7676 (N_7676,N_3323,N_1402);
or U7677 (N_7677,N_287,N_2414);
and U7678 (N_7678,N_952,N_1424);
and U7679 (N_7679,N_2647,N_1651);
nand U7680 (N_7680,N_1500,N_3998);
and U7681 (N_7681,N_3935,N_1571);
or U7682 (N_7682,N_3576,N_1840);
xor U7683 (N_7683,N_3629,N_3713);
nand U7684 (N_7684,N_2707,N_2365);
nor U7685 (N_7685,N_2969,N_785);
nand U7686 (N_7686,N_163,N_2947);
xnor U7687 (N_7687,N_2486,N_2455);
nor U7688 (N_7688,N_930,N_1498);
xor U7689 (N_7689,N_2923,N_3933);
and U7690 (N_7690,N_277,N_3987);
nor U7691 (N_7691,N_2872,N_2343);
nor U7692 (N_7692,N_91,N_3039);
nand U7693 (N_7693,N_1440,N_3917);
xnor U7694 (N_7694,N_2673,N_3482);
nor U7695 (N_7695,N_1568,N_3048);
xor U7696 (N_7696,N_3328,N_236);
nand U7697 (N_7697,N_865,N_1434);
and U7698 (N_7698,N_3022,N_745);
xnor U7699 (N_7699,N_3314,N_2663);
nand U7700 (N_7700,N_1400,N_2303);
and U7701 (N_7701,N_3742,N_3340);
and U7702 (N_7702,N_2448,N_3094);
nor U7703 (N_7703,N_947,N_1376);
nor U7704 (N_7704,N_3583,N_3384);
xor U7705 (N_7705,N_935,N_189);
xor U7706 (N_7706,N_3714,N_3123);
xnor U7707 (N_7707,N_3023,N_1387);
xor U7708 (N_7708,N_330,N_1861);
or U7709 (N_7709,N_150,N_2000);
nor U7710 (N_7710,N_18,N_3055);
or U7711 (N_7711,N_2401,N_1489);
xor U7712 (N_7712,N_3625,N_3841);
or U7713 (N_7713,N_2134,N_3343);
xnor U7714 (N_7714,N_152,N_1439);
or U7715 (N_7715,N_977,N_300);
and U7716 (N_7716,N_1286,N_3600);
nor U7717 (N_7717,N_1623,N_2475);
nor U7718 (N_7718,N_1256,N_2498);
and U7719 (N_7719,N_2724,N_1092);
nand U7720 (N_7720,N_488,N_1935);
nand U7721 (N_7721,N_1374,N_3660);
xor U7722 (N_7722,N_2955,N_346);
xnor U7723 (N_7723,N_3372,N_784);
nand U7724 (N_7724,N_3408,N_2729);
or U7725 (N_7725,N_3597,N_1196);
nor U7726 (N_7726,N_3372,N_1519);
nand U7727 (N_7727,N_3836,N_504);
nand U7728 (N_7728,N_3213,N_857);
or U7729 (N_7729,N_1743,N_374);
nand U7730 (N_7730,N_3042,N_813);
and U7731 (N_7731,N_179,N_2825);
and U7732 (N_7732,N_2719,N_2829);
xor U7733 (N_7733,N_873,N_3077);
xor U7734 (N_7734,N_184,N_3725);
or U7735 (N_7735,N_1293,N_1116);
nand U7736 (N_7736,N_638,N_1857);
and U7737 (N_7737,N_891,N_1495);
nor U7738 (N_7738,N_617,N_41);
or U7739 (N_7739,N_75,N_3406);
nand U7740 (N_7740,N_3800,N_343);
and U7741 (N_7741,N_3890,N_2511);
or U7742 (N_7742,N_2633,N_3516);
nand U7743 (N_7743,N_864,N_3318);
or U7744 (N_7744,N_1002,N_1380);
xnor U7745 (N_7745,N_1740,N_136);
nor U7746 (N_7746,N_397,N_2205);
nor U7747 (N_7747,N_1640,N_3347);
nand U7748 (N_7748,N_646,N_1921);
nand U7749 (N_7749,N_2051,N_430);
nor U7750 (N_7750,N_2653,N_3466);
or U7751 (N_7751,N_1185,N_2159);
xor U7752 (N_7752,N_3994,N_1224);
and U7753 (N_7753,N_902,N_1972);
or U7754 (N_7754,N_3707,N_852);
nand U7755 (N_7755,N_3649,N_2982);
or U7756 (N_7756,N_1149,N_542);
nand U7757 (N_7757,N_2834,N_3645);
xnor U7758 (N_7758,N_1024,N_1945);
nor U7759 (N_7759,N_2109,N_2565);
nand U7760 (N_7760,N_2466,N_581);
or U7761 (N_7761,N_405,N_1705);
nor U7762 (N_7762,N_898,N_1272);
nand U7763 (N_7763,N_1000,N_190);
nand U7764 (N_7764,N_1428,N_1627);
and U7765 (N_7765,N_3491,N_586);
or U7766 (N_7766,N_1312,N_766);
nor U7767 (N_7767,N_1420,N_1206);
nand U7768 (N_7768,N_547,N_2049);
or U7769 (N_7769,N_422,N_13);
and U7770 (N_7770,N_2025,N_3953);
or U7771 (N_7771,N_3132,N_2350);
or U7772 (N_7772,N_203,N_3290);
nor U7773 (N_7773,N_2121,N_1420);
and U7774 (N_7774,N_31,N_3821);
and U7775 (N_7775,N_1457,N_3853);
and U7776 (N_7776,N_3974,N_105);
nand U7777 (N_7777,N_2582,N_1966);
or U7778 (N_7778,N_2555,N_693);
nand U7779 (N_7779,N_3284,N_2097);
or U7780 (N_7780,N_756,N_3604);
nor U7781 (N_7781,N_720,N_3847);
xnor U7782 (N_7782,N_93,N_3598);
xor U7783 (N_7783,N_3572,N_557);
or U7784 (N_7784,N_364,N_2986);
and U7785 (N_7785,N_3900,N_2919);
and U7786 (N_7786,N_3808,N_3978);
and U7787 (N_7787,N_3544,N_426);
or U7788 (N_7788,N_3915,N_2276);
nor U7789 (N_7789,N_2764,N_131);
xor U7790 (N_7790,N_3332,N_137);
or U7791 (N_7791,N_3274,N_2585);
xor U7792 (N_7792,N_2162,N_3186);
and U7793 (N_7793,N_3879,N_966);
nand U7794 (N_7794,N_1386,N_2539);
or U7795 (N_7795,N_1498,N_845);
xnor U7796 (N_7796,N_2039,N_660);
nand U7797 (N_7797,N_294,N_1201);
xor U7798 (N_7798,N_83,N_3412);
and U7799 (N_7799,N_3907,N_3965);
and U7800 (N_7800,N_12,N_1733);
or U7801 (N_7801,N_3512,N_181);
nor U7802 (N_7802,N_3323,N_1437);
and U7803 (N_7803,N_219,N_515);
and U7804 (N_7804,N_3757,N_2860);
nor U7805 (N_7805,N_2953,N_3167);
nor U7806 (N_7806,N_1190,N_712);
or U7807 (N_7807,N_540,N_3646);
and U7808 (N_7808,N_891,N_3223);
nand U7809 (N_7809,N_982,N_1521);
or U7810 (N_7810,N_3680,N_3162);
nand U7811 (N_7811,N_2488,N_3935);
and U7812 (N_7812,N_2426,N_2498);
xor U7813 (N_7813,N_183,N_2775);
nand U7814 (N_7814,N_1126,N_2284);
and U7815 (N_7815,N_1963,N_338);
and U7816 (N_7816,N_1683,N_1571);
nand U7817 (N_7817,N_3856,N_1886);
nand U7818 (N_7818,N_68,N_1813);
nor U7819 (N_7819,N_2343,N_1178);
or U7820 (N_7820,N_1796,N_1573);
xnor U7821 (N_7821,N_3687,N_1691);
nand U7822 (N_7822,N_769,N_2367);
nor U7823 (N_7823,N_3982,N_3764);
or U7824 (N_7824,N_2696,N_2706);
xnor U7825 (N_7825,N_2449,N_2359);
xnor U7826 (N_7826,N_1245,N_174);
nor U7827 (N_7827,N_3545,N_2916);
nor U7828 (N_7828,N_475,N_3168);
nand U7829 (N_7829,N_798,N_1130);
or U7830 (N_7830,N_2097,N_793);
xor U7831 (N_7831,N_3393,N_1221);
xor U7832 (N_7832,N_361,N_3);
nor U7833 (N_7833,N_3715,N_1495);
nor U7834 (N_7834,N_3755,N_2104);
xnor U7835 (N_7835,N_310,N_503);
and U7836 (N_7836,N_455,N_2487);
or U7837 (N_7837,N_524,N_2663);
xor U7838 (N_7838,N_3936,N_34);
nor U7839 (N_7839,N_686,N_3674);
or U7840 (N_7840,N_1465,N_3474);
nor U7841 (N_7841,N_3217,N_2477);
and U7842 (N_7842,N_2085,N_3333);
xor U7843 (N_7843,N_3801,N_1675);
nor U7844 (N_7844,N_3298,N_3503);
or U7845 (N_7845,N_2939,N_3583);
xnor U7846 (N_7846,N_2876,N_3135);
and U7847 (N_7847,N_2804,N_1027);
nand U7848 (N_7848,N_1965,N_3149);
nor U7849 (N_7849,N_1030,N_655);
nand U7850 (N_7850,N_3869,N_3938);
nand U7851 (N_7851,N_2587,N_3562);
or U7852 (N_7852,N_1738,N_2627);
and U7853 (N_7853,N_3680,N_343);
or U7854 (N_7854,N_310,N_2868);
xnor U7855 (N_7855,N_3236,N_2105);
or U7856 (N_7856,N_918,N_2686);
xnor U7857 (N_7857,N_2079,N_3795);
or U7858 (N_7858,N_148,N_323);
xnor U7859 (N_7859,N_852,N_3104);
xor U7860 (N_7860,N_2940,N_3764);
nand U7861 (N_7861,N_1196,N_205);
xor U7862 (N_7862,N_3452,N_3449);
or U7863 (N_7863,N_3691,N_2855);
or U7864 (N_7864,N_2090,N_945);
nand U7865 (N_7865,N_3640,N_2077);
or U7866 (N_7866,N_2410,N_2432);
nand U7867 (N_7867,N_312,N_1818);
and U7868 (N_7868,N_3181,N_2918);
or U7869 (N_7869,N_973,N_3994);
or U7870 (N_7870,N_250,N_972);
nor U7871 (N_7871,N_763,N_3587);
and U7872 (N_7872,N_3415,N_3691);
and U7873 (N_7873,N_21,N_3575);
nand U7874 (N_7874,N_937,N_2037);
nor U7875 (N_7875,N_371,N_2856);
nand U7876 (N_7876,N_3081,N_3220);
xor U7877 (N_7877,N_1614,N_1517);
or U7878 (N_7878,N_2658,N_3979);
nor U7879 (N_7879,N_2656,N_3334);
nand U7880 (N_7880,N_2626,N_1697);
nand U7881 (N_7881,N_3964,N_2887);
nand U7882 (N_7882,N_2434,N_951);
xnor U7883 (N_7883,N_725,N_3286);
nand U7884 (N_7884,N_1629,N_2780);
nor U7885 (N_7885,N_1766,N_1506);
and U7886 (N_7886,N_1347,N_1164);
and U7887 (N_7887,N_941,N_2690);
nand U7888 (N_7888,N_3638,N_2599);
nand U7889 (N_7889,N_2508,N_3369);
or U7890 (N_7890,N_2364,N_2927);
or U7891 (N_7891,N_2531,N_3978);
nand U7892 (N_7892,N_827,N_1320);
and U7893 (N_7893,N_2518,N_1170);
nand U7894 (N_7894,N_865,N_661);
nor U7895 (N_7895,N_2255,N_1841);
or U7896 (N_7896,N_1761,N_940);
xnor U7897 (N_7897,N_2099,N_3325);
nor U7898 (N_7898,N_2372,N_3678);
xor U7899 (N_7899,N_3918,N_1416);
nor U7900 (N_7900,N_2204,N_1208);
nor U7901 (N_7901,N_3158,N_3608);
xor U7902 (N_7902,N_1038,N_2083);
and U7903 (N_7903,N_1241,N_10);
and U7904 (N_7904,N_1425,N_3113);
or U7905 (N_7905,N_903,N_1773);
and U7906 (N_7906,N_1672,N_1762);
and U7907 (N_7907,N_1370,N_2871);
nor U7908 (N_7908,N_1887,N_3305);
and U7909 (N_7909,N_608,N_2416);
nand U7910 (N_7910,N_283,N_1197);
and U7911 (N_7911,N_1563,N_3865);
nor U7912 (N_7912,N_2097,N_869);
and U7913 (N_7913,N_3168,N_1380);
nand U7914 (N_7914,N_44,N_26);
nand U7915 (N_7915,N_1402,N_588);
nand U7916 (N_7916,N_2511,N_803);
xor U7917 (N_7917,N_2159,N_1053);
nand U7918 (N_7918,N_3358,N_2738);
and U7919 (N_7919,N_3576,N_2978);
or U7920 (N_7920,N_3100,N_2360);
nand U7921 (N_7921,N_1957,N_1995);
nor U7922 (N_7922,N_694,N_3019);
nand U7923 (N_7923,N_2396,N_1193);
nand U7924 (N_7924,N_2763,N_1016);
nand U7925 (N_7925,N_3774,N_536);
or U7926 (N_7926,N_2810,N_1470);
and U7927 (N_7927,N_384,N_3396);
nor U7928 (N_7928,N_3275,N_540);
xor U7929 (N_7929,N_152,N_2002);
xor U7930 (N_7930,N_2667,N_2805);
or U7931 (N_7931,N_3715,N_3546);
or U7932 (N_7932,N_3648,N_961);
nor U7933 (N_7933,N_395,N_931);
and U7934 (N_7934,N_2057,N_2141);
or U7935 (N_7935,N_2475,N_3783);
nand U7936 (N_7936,N_959,N_2787);
nor U7937 (N_7937,N_3882,N_1479);
and U7938 (N_7938,N_2577,N_290);
nand U7939 (N_7939,N_2777,N_1573);
or U7940 (N_7940,N_2733,N_831);
or U7941 (N_7941,N_2274,N_1964);
nand U7942 (N_7942,N_1201,N_972);
nor U7943 (N_7943,N_1605,N_2554);
xor U7944 (N_7944,N_3507,N_835);
or U7945 (N_7945,N_1667,N_1169);
and U7946 (N_7946,N_404,N_2136);
or U7947 (N_7947,N_1843,N_2836);
xnor U7948 (N_7948,N_3451,N_3600);
nor U7949 (N_7949,N_1236,N_1247);
nor U7950 (N_7950,N_931,N_3076);
xor U7951 (N_7951,N_3857,N_2298);
nor U7952 (N_7952,N_1836,N_2953);
nor U7953 (N_7953,N_1249,N_2928);
xor U7954 (N_7954,N_3922,N_1867);
or U7955 (N_7955,N_65,N_989);
xnor U7956 (N_7956,N_3521,N_623);
or U7957 (N_7957,N_2842,N_929);
and U7958 (N_7958,N_3383,N_113);
or U7959 (N_7959,N_12,N_2476);
nand U7960 (N_7960,N_293,N_2172);
or U7961 (N_7961,N_3452,N_3955);
and U7962 (N_7962,N_168,N_2111);
and U7963 (N_7963,N_713,N_1089);
nor U7964 (N_7964,N_1752,N_2056);
nand U7965 (N_7965,N_920,N_846);
or U7966 (N_7966,N_324,N_400);
and U7967 (N_7967,N_914,N_3027);
and U7968 (N_7968,N_1131,N_1178);
nand U7969 (N_7969,N_3090,N_3256);
nor U7970 (N_7970,N_549,N_1927);
xnor U7971 (N_7971,N_3716,N_1074);
nand U7972 (N_7972,N_2664,N_3350);
or U7973 (N_7973,N_3675,N_1158);
nand U7974 (N_7974,N_2634,N_475);
or U7975 (N_7975,N_741,N_3002);
nand U7976 (N_7976,N_876,N_1765);
nor U7977 (N_7977,N_278,N_963);
and U7978 (N_7978,N_958,N_3388);
nand U7979 (N_7979,N_2098,N_3315);
nand U7980 (N_7980,N_2147,N_2474);
and U7981 (N_7981,N_15,N_1690);
nor U7982 (N_7982,N_1687,N_2253);
nor U7983 (N_7983,N_2129,N_2667);
nand U7984 (N_7984,N_1969,N_3657);
nand U7985 (N_7985,N_81,N_3993);
and U7986 (N_7986,N_80,N_2965);
xor U7987 (N_7987,N_1482,N_2298);
and U7988 (N_7988,N_3710,N_78);
nor U7989 (N_7989,N_2832,N_1543);
or U7990 (N_7990,N_3695,N_1029);
and U7991 (N_7991,N_2696,N_1578);
nand U7992 (N_7992,N_255,N_2175);
nor U7993 (N_7993,N_1590,N_1757);
and U7994 (N_7994,N_615,N_1458);
nand U7995 (N_7995,N_2600,N_2798);
nand U7996 (N_7996,N_1310,N_566);
or U7997 (N_7997,N_3026,N_847);
and U7998 (N_7998,N_1566,N_2117);
nand U7999 (N_7999,N_1871,N_249);
and U8000 (N_8000,N_5011,N_4026);
xnor U8001 (N_8001,N_6488,N_4333);
nor U8002 (N_8002,N_4299,N_7135);
nand U8003 (N_8003,N_5015,N_5110);
nand U8004 (N_8004,N_4501,N_5808);
and U8005 (N_8005,N_4843,N_7730);
nor U8006 (N_8006,N_4669,N_7616);
nand U8007 (N_8007,N_4628,N_5669);
nor U8008 (N_8008,N_4246,N_4869);
or U8009 (N_8009,N_5656,N_5544);
nor U8010 (N_8010,N_5214,N_5264);
nor U8011 (N_8011,N_6332,N_6453);
nor U8012 (N_8012,N_4516,N_6907);
or U8013 (N_8013,N_7691,N_7658);
nor U8014 (N_8014,N_6195,N_5225);
nor U8015 (N_8015,N_4047,N_7073);
and U8016 (N_8016,N_7092,N_5397);
and U8017 (N_8017,N_7447,N_6759);
or U8018 (N_8018,N_5887,N_6828);
or U8019 (N_8019,N_4506,N_5112);
nor U8020 (N_8020,N_5921,N_4830);
or U8021 (N_8021,N_5687,N_4155);
xnor U8022 (N_8022,N_4953,N_5806);
and U8023 (N_8023,N_4563,N_5106);
xnor U8024 (N_8024,N_7442,N_6309);
nand U8025 (N_8025,N_7376,N_6266);
and U8026 (N_8026,N_6871,N_6348);
xnor U8027 (N_8027,N_7938,N_6702);
and U8028 (N_8028,N_7881,N_7731);
or U8029 (N_8029,N_7665,N_7509);
xnor U8030 (N_8030,N_5568,N_7986);
nor U8031 (N_8031,N_4507,N_6933);
xor U8032 (N_8032,N_5021,N_4440);
or U8033 (N_8033,N_6654,N_6604);
xnor U8034 (N_8034,N_6032,N_6710);
nor U8035 (N_8035,N_4379,N_4231);
nand U8036 (N_8036,N_7241,N_6399);
and U8037 (N_8037,N_6910,N_5729);
and U8038 (N_8038,N_5027,N_5467);
or U8039 (N_8039,N_4374,N_4559);
xnor U8040 (N_8040,N_6324,N_4193);
nand U8041 (N_8041,N_5678,N_4046);
and U8042 (N_8042,N_5444,N_4300);
and U8043 (N_8043,N_5658,N_5240);
xor U8044 (N_8044,N_4122,N_6406);
or U8045 (N_8045,N_7670,N_7985);
xor U8046 (N_8046,N_4050,N_7928);
nor U8047 (N_8047,N_4138,N_4065);
or U8048 (N_8048,N_6262,N_4557);
xor U8049 (N_8049,N_4127,N_4357);
nor U8050 (N_8050,N_7176,N_5630);
nand U8051 (N_8051,N_6043,N_6184);
nand U8052 (N_8052,N_6113,N_4492);
xnor U8053 (N_8053,N_5255,N_6967);
nor U8054 (N_8054,N_4130,N_5781);
nand U8055 (N_8055,N_5171,N_5952);
or U8056 (N_8056,N_7811,N_5280);
or U8057 (N_8057,N_6872,N_5035);
xor U8058 (N_8058,N_7686,N_5212);
and U8059 (N_8059,N_5742,N_6561);
and U8060 (N_8060,N_6424,N_4799);
xnor U8061 (N_8061,N_7266,N_5968);
nor U8062 (N_8062,N_5030,N_5843);
xnor U8063 (N_8063,N_6592,N_5004);
nand U8064 (N_8064,N_6006,N_5946);
nand U8065 (N_8065,N_6436,N_5713);
or U8066 (N_8066,N_5067,N_6943);
nand U8067 (N_8067,N_7210,N_6499);
xor U8068 (N_8068,N_7931,N_6473);
or U8069 (N_8069,N_6186,N_5470);
nor U8070 (N_8070,N_7402,N_6882);
or U8071 (N_8071,N_7059,N_7606);
nand U8072 (N_8072,N_7747,N_5538);
nor U8073 (N_8073,N_7152,N_4608);
or U8074 (N_8074,N_6680,N_7309);
xnor U8075 (N_8075,N_5517,N_5271);
and U8076 (N_8076,N_7288,N_6439);
nand U8077 (N_8077,N_4917,N_4933);
nor U8078 (N_8078,N_6743,N_5247);
xnor U8079 (N_8079,N_7192,N_6272);
nand U8080 (N_8080,N_5790,N_7901);
or U8081 (N_8081,N_6832,N_7111);
nand U8082 (N_8082,N_4409,N_5681);
and U8083 (N_8083,N_4522,N_4739);
or U8084 (N_8084,N_5583,N_7307);
nand U8085 (N_8085,N_4405,N_4326);
or U8086 (N_8086,N_7071,N_4452);
and U8087 (N_8087,N_6545,N_5262);
and U8088 (N_8088,N_5132,N_7050);
and U8089 (N_8089,N_5433,N_5780);
nand U8090 (N_8090,N_4024,N_6254);
and U8091 (N_8091,N_4717,N_5490);
xor U8092 (N_8092,N_5496,N_5267);
xor U8093 (N_8093,N_6117,N_6143);
nand U8094 (N_8094,N_7108,N_4632);
nor U8095 (N_8095,N_6288,N_4599);
or U8096 (N_8096,N_6377,N_7429);
and U8097 (N_8097,N_4412,N_4012);
nand U8098 (N_8098,N_5390,N_7704);
nand U8099 (N_8099,N_5498,N_4881);
nand U8100 (N_8100,N_4825,N_7661);
nand U8101 (N_8101,N_6628,N_4515);
and U8102 (N_8102,N_5291,N_7409);
nor U8103 (N_8103,N_4081,N_5322);
or U8104 (N_8104,N_5674,N_5492);
xor U8105 (N_8105,N_6596,N_6625);
xor U8106 (N_8106,N_5315,N_4797);
nand U8107 (N_8107,N_4631,N_4644);
xor U8108 (N_8108,N_4248,N_5254);
xor U8109 (N_8109,N_5393,N_6898);
xor U8110 (N_8110,N_6648,N_7721);
and U8111 (N_8111,N_6397,N_6347);
xor U8112 (N_8112,N_7656,N_6569);
nor U8113 (N_8113,N_5596,N_6552);
xnor U8114 (N_8114,N_4304,N_7366);
nand U8115 (N_8115,N_6790,N_7400);
nor U8116 (N_8116,N_6979,N_4359);
or U8117 (N_8117,N_4441,N_7741);
or U8118 (N_8118,N_6445,N_7879);
and U8119 (N_8119,N_6753,N_4150);
xor U8120 (N_8120,N_4167,N_7662);
or U8121 (N_8121,N_6082,N_6854);
and U8122 (N_8122,N_6926,N_5976);
xor U8123 (N_8123,N_7281,N_6106);
and U8124 (N_8124,N_7696,N_5890);
nand U8125 (N_8125,N_4884,N_6206);
or U8126 (N_8126,N_5526,N_6644);
nand U8127 (N_8127,N_4156,N_5119);
and U8128 (N_8128,N_7086,N_5978);
nor U8129 (N_8129,N_6181,N_5204);
xor U8130 (N_8130,N_5605,N_4879);
nor U8131 (N_8131,N_4232,N_7875);
or U8132 (N_8132,N_7773,N_5823);
or U8133 (N_8133,N_4927,N_5775);
xnor U8134 (N_8134,N_7983,N_6835);
nand U8135 (N_8135,N_4703,N_4419);
xnor U8136 (N_8136,N_5885,N_5032);
nor U8137 (N_8137,N_7461,N_6142);
nor U8138 (N_8138,N_4236,N_5524);
nor U8139 (N_8139,N_5279,N_5845);
nand U8140 (N_8140,N_4479,N_6018);
and U8141 (N_8141,N_7479,N_6825);
nor U8142 (N_8142,N_5772,N_6598);
and U8143 (N_8143,N_5536,N_4991);
xor U8144 (N_8144,N_5796,N_7069);
and U8145 (N_8145,N_5344,N_5288);
or U8146 (N_8146,N_6443,N_5940);
xnor U8147 (N_8147,N_5202,N_7531);
nor U8148 (N_8148,N_7585,N_6541);
or U8149 (N_8149,N_6720,N_4311);
xor U8150 (N_8150,N_6161,N_4029);
xnor U8151 (N_8151,N_7627,N_5017);
nand U8152 (N_8152,N_7868,N_5882);
or U8153 (N_8153,N_4380,N_6028);
or U8154 (N_8154,N_4905,N_5399);
nand U8155 (N_8155,N_7379,N_7638);
and U8156 (N_8156,N_5599,N_6593);
or U8157 (N_8157,N_4275,N_5158);
nor U8158 (N_8158,N_4614,N_6237);
and U8159 (N_8159,N_7488,N_6489);
nor U8160 (N_8160,N_6256,N_7882);
and U8161 (N_8161,N_4609,N_7935);
nor U8162 (N_8162,N_7578,N_4903);
xnor U8163 (N_8163,N_6997,N_7280);
xor U8164 (N_8164,N_6877,N_6883);
and U8165 (N_8165,N_4158,N_6211);
nand U8166 (N_8166,N_5215,N_7269);
and U8167 (N_8167,N_6233,N_7300);
xor U8168 (N_8168,N_6135,N_6989);
nand U8169 (N_8169,N_7399,N_6159);
and U8170 (N_8170,N_7864,N_4372);
nand U8171 (N_8171,N_4861,N_6626);
xor U8172 (N_8172,N_7748,N_7386);
or U8173 (N_8173,N_5146,N_4640);
or U8174 (N_8174,N_5220,N_4673);
nor U8175 (N_8175,N_4698,N_4543);
nor U8176 (N_8176,N_7609,N_7457);
xnor U8177 (N_8177,N_5121,N_6846);
or U8178 (N_8178,N_7951,N_5539);
nor U8179 (N_8179,N_6641,N_6158);
xor U8180 (N_8180,N_4654,N_7624);
nand U8181 (N_8181,N_7746,N_6634);
xor U8182 (N_8182,N_4104,N_6605);
or U8183 (N_8183,N_4023,N_6026);
nand U8184 (N_8184,N_4320,N_6708);
and U8185 (N_8185,N_6789,N_6056);
nor U8186 (N_8186,N_5797,N_6468);
or U8187 (N_8187,N_7452,N_4641);
xnor U8188 (N_8188,N_7497,N_6966);
xor U8189 (N_8189,N_7714,N_6418);
or U8190 (N_8190,N_4438,N_4459);
nand U8191 (N_8191,N_5786,N_7889);
nand U8192 (N_8192,N_5038,N_7233);
and U8193 (N_8193,N_7297,N_5779);
nand U8194 (N_8194,N_4367,N_6948);
nor U8195 (N_8195,N_6707,N_6880);
nand U8196 (N_8196,N_4291,N_7956);
nand U8197 (N_8197,N_6820,N_6518);
nand U8198 (N_8198,N_4085,N_4755);
and U8199 (N_8199,N_6071,N_5556);
xor U8200 (N_8200,N_7754,N_7100);
and U8201 (N_8201,N_5703,N_4356);
nand U8202 (N_8202,N_4472,N_5062);
nor U8203 (N_8203,N_6420,N_6294);
xnor U8204 (N_8204,N_6160,N_7155);
nor U8205 (N_8205,N_6042,N_6075);
xnor U8206 (N_8206,N_7989,N_7795);
nand U8207 (N_8207,N_6601,N_5512);
or U8208 (N_8208,N_5275,N_6249);
nor U8209 (N_8209,N_7924,N_4593);
xor U8210 (N_8210,N_5403,N_6778);
or U8211 (N_8211,N_6293,N_4022);
nor U8212 (N_8212,N_7012,N_7314);
or U8213 (N_8213,N_4382,N_6289);
and U8214 (N_8214,N_5977,N_5396);
xor U8215 (N_8215,N_4317,N_6922);
or U8216 (N_8216,N_7343,N_7642);
nand U8217 (N_8217,N_4341,N_6532);
and U8218 (N_8218,N_6386,N_6960);
nand U8219 (N_8219,N_5651,N_4836);
nand U8220 (N_8220,N_7356,N_4396);
xor U8221 (N_8221,N_6565,N_4094);
and U8222 (N_8222,N_7854,N_6187);
xnor U8223 (N_8223,N_4048,N_5418);
xor U8224 (N_8224,N_6769,N_6834);
nand U8225 (N_8225,N_4141,N_4213);
nand U8226 (N_8226,N_7674,N_7319);
nor U8227 (N_8227,N_6435,N_5653);
or U8228 (N_8228,N_6996,N_7637);
or U8229 (N_8229,N_5206,N_7903);
xor U8230 (N_8230,N_7002,N_7843);
or U8231 (N_8231,N_6061,N_6542);
nand U8232 (N_8232,N_4277,N_5289);
or U8233 (N_8233,N_6889,N_6422);
and U8234 (N_8234,N_5569,N_4980);
nor U8235 (N_8235,N_4073,N_7040);
or U8236 (N_8236,N_6809,N_7412);
or U8237 (N_8237,N_5350,N_4388);
nand U8238 (N_8238,N_7713,N_6354);
xor U8239 (N_8239,N_5364,N_4194);
xnor U8240 (N_8240,N_4037,N_5691);
nand U8241 (N_8241,N_5353,N_6353);
nor U8242 (N_8242,N_4763,N_6325);
and U8243 (N_8243,N_6315,N_4265);
and U8244 (N_8244,N_7772,N_5666);
and U8245 (N_8245,N_5499,N_7635);
and U8246 (N_8246,N_5413,N_5239);
nand U8247 (N_8247,N_4790,N_4660);
nor U8248 (N_8248,N_6686,N_5566);
and U8249 (N_8249,N_6972,N_6307);
nand U8250 (N_8250,N_5545,N_5486);
xor U8251 (N_8251,N_6652,N_6805);
or U8252 (N_8252,N_7774,N_5114);
nor U8253 (N_8253,N_5075,N_4488);
nor U8254 (N_8254,N_7743,N_7087);
nor U8255 (N_8255,N_4421,N_5714);
and U8256 (N_8256,N_6793,N_5912);
xor U8257 (N_8257,N_7380,N_6658);
or U8258 (N_8258,N_5815,N_5902);
nor U8259 (N_8259,N_7188,N_7478);
xnor U8260 (N_8260,N_4181,N_6303);
or U8261 (N_8261,N_6058,N_5056);
xnor U8262 (N_8262,N_4298,N_6137);
nor U8263 (N_8263,N_6215,N_7676);
nor U8264 (N_8264,N_4993,N_6934);
nor U8265 (N_8265,N_7337,N_6306);
or U8266 (N_8266,N_6537,N_4571);
nand U8267 (N_8267,N_5466,N_5865);
nor U8268 (N_8268,N_6494,N_6388);
xor U8269 (N_8269,N_4596,N_6697);
xnor U8270 (N_8270,N_6801,N_4397);
nor U8271 (N_8271,N_6799,N_7855);
and U8272 (N_8272,N_5919,N_6768);
and U8273 (N_8273,N_5861,N_5179);
xor U8274 (N_8274,N_5161,N_6337);
xor U8275 (N_8275,N_4491,N_5031);
and U8276 (N_8276,N_7137,N_6166);
nand U8277 (N_8277,N_6699,N_4895);
and U8278 (N_8278,N_7758,N_7377);
or U8279 (N_8279,N_4948,N_7945);
and U8280 (N_8280,N_4683,N_6078);
xnor U8281 (N_8281,N_4649,N_4365);
xor U8282 (N_8282,N_5810,N_6393);
xnor U8283 (N_8283,N_6385,N_6150);
nor U8284 (N_8284,N_6069,N_5620);
nor U8285 (N_8285,N_6946,N_5229);
xnor U8286 (N_8286,N_4994,N_5740);
or U8287 (N_8287,N_7278,N_5276);
nand U8288 (N_8288,N_7853,N_4377);
or U8289 (N_8289,N_7990,N_5708);
and U8290 (N_8290,N_6915,N_6346);
nor U8291 (N_8291,N_5553,N_6767);
or U8292 (N_8292,N_6570,N_7055);
nand U8293 (N_8293,N_4885,N_7567);
nand U8294 (N_8294,N_6030,N_7859);
or U8295 (N_8295,N_7098,N_4972);
nand U8296 (N_8296,N_7798,N_7061);
nor U8297 (N_8297,N_7183,N_5250);
and U8298 (N_8298,N_6020,N_5047);
nand U8299 (N_8299,N_5287,N_7886);
and U8300 (N_8300,N_4757,N_7866);
nor U8301 (N_8301,N_5881,N_4659);
and U8302 (N_8302,N_7202,N_6819);
nand U8303 (N_8303,N_4692,N_5958);
xor U8304 (N_8304,N_5257,N_5515);
or U8305 (N_8305,N_5311,N_4893);
xnor U8306 (N_8306,N_7425,N_4618);
xor U8307 (N_8307,N_6705,N_4486);
nor U8308 (N_8308,N_5195,N_6450);
nand U8309 (N_8309,N_6007,N_4096);
nand U8310 (N_8310,N_4108,N_6665);
or U8311 (N_8311,N_5480,N_6119);
xnor U8312 (N_8312,N_5489,N_5677);
or U8313 (N_8313,N_6299,N_5246);
nand U8314 (N_8314,N_7724,N_4661);
nor U8315 (N_8315,N_5870,N_7024);
nor U8316 (N_8316,N_4575,N_6320);
xnor U8317 (N_8317,N_7821,N_7131);
or U8318 (N_8318,N_5048,N_7367);
and U8319 (N_8319,N_6088,N_5685);
xor U8320 (N_8320,N_4935,N_6437);
nor U8321 (N_8321,N_6923,N_7545);
or U8322 (N_8322,N_4307,N_5154);
nand U8323 (N_8323,N_7922,N_4016);
nand U8324 (N_8324,N_4959,N_7562);
nand U8325 (N_8325,N_7148,N_7296);
nand U8326 (N_8326,N_7602,N_6602);
or U8327 (N_8327,N_7783,N_7787);
or U8328 (N_8328,N_4222,N_6065);
nor U8329 (N_8329,N_5847,N_7660);
xnor U8330 (N_8330,N_5901,N_6275);
and U8331 (N_8331,N_6177,N_6099);
xnor U8332 (N_8332,N_5231,N_7801);
and U8333 (N_8333,N_6752,N_6991);
and U8334 (N_8334,N_5458,N_6362);
or U8335 (N_8335,N_4762,N_4498);
nand U8336 (N_8336,N_7967,N_5338);
nand U8337 (N_8337,N_4818,N_7358);
and U8338 (N_8338,N_6505,N_6496);
nor U8339 (N_8339,N_6140,N_6970);
xnor U8340 (N_8340,N_5943,N_4053);
xor U8341 (N_8341,N_4204,N_4574);
nand U8342 (N_8342,N_7178,N_6920);
nand U8343 (N_8343,N_7632,N_4713);
nand U8344 (N_8344,N_7083,N_6958);
nor U8345 (N_8345,N_4091,N_7958);
or U8346 (N_8346,N_5629,N_5707);
nor U8347 (N_8347,N_5970,N_7294);
nand U8348 (N_8348,N_7852,N_7397);
nand U8349 (N_8349,N_6380,N_4215);
xor U8350 (N_8350,N_6156,N_7819);
xor U8351 (N_8351,N_5003,N_7739);
nor U8352 (N_8352,N_7907,N_6701);
nor U8353 (N_8353,N_6528,N_4615);
nor U8354 (N_8354,N_7289,N_5582);
and U8355 (N_8355,N_4592,N_7825);
or U8356 (N_8356,N_4667,N_7978);
nor U8357 (N_8357,N_6929,N_6531);
nand U8358 (N_8358,N_6067,N_6090);
or U8359 (N_8359,N_6227,N_7926);
or U8360 (N_8360,N_5145,N_5180);
and U8361 (N_8361,N_6257,N_7459);
nand U8362 (N_8362,N_4961,N_6433);
or U8363 (N_8363,N_7211,N_7162);
nand U8364 (N_8364,N_5755,N_7937);
or U8365 (N_8365,N_6214,N_6739);
nor U8366 (N_8366,N_5826,N_7678);
xor U8367 (N_8367,N_7502,N_6260);
nand U8368 (N_8368,N_5571,N_4852);
xor U8369 (N_8369,N_6270,N_5450);
and U8370 (N_8370,N_4199,N_6683);
or U8371 (N_8371,N_7027,N_7503);
nand U8372 (N_8372,N_5717,N_7416);
xnor U8373 (N_8373,N_6218,N_6999);
nand U8374 (N_8374,N_5210,N_5337);
xor U8375 (N_8375,N_5739,N_5925);
xnor U8376 (N_8376,N_5648,N_7483);
nand U8377 (N_8377,N_6642,N_6956);
or U8378 (N_8378,N_7433,N_6807);
nor U8379 (N_8379,N_4846,N_5420);
xor U8380 (N_8380,N_7372,N_7778);
or U8381 (N_8381,N_5473,N_4312);
and U8382 (N_8382,N_4912,N_4146);
nand U8383 (N_8383,N_7293,N_6931);
or U8384 (N_8384,N_6118,N_4476);
xnor U8385 (N_8385,N_4803,N_4378);
nand U8386 (N_8386,N_6107,N_4495);
and U8387 (N_8387,N_4366,N_7733);
nor U8388 (N_8388,N_7789,N_7756);
or U8389 (N_8389,N_7341,N_6977);
xor U8390 (N_8390,N_4785,N_5323);
or U8391 (N_8391,N_7598,N_4144);
nor U8392 (N_8392,N_5643,N_7918);
xnor U8393 (N_8393,N_7501,N_6583);
nand U8394 (N_8394,N_5265,N_4671);
xnor U8395 (N_8395,N_6250,N_7646);
nor U8396 (N_8396,N_7641,N_4975);
or U8397 (N_8397,N_5842,N_6857);
nor U8398 (N_8398,N_5252,N_4160);
xnor U8399 (N_8399,N_4668,N_4678);
xor U8400 (N_8400,N_6190,N_5563);
and U8401 (N_8401,N_7818,N_7890);
xor U8402 (N_8402,N_5966,N_7534);
and U8403 (N_8403,N_5661,N_4734);
nor U8404 (N_8404,N_7446,N_6247);
nand U8405 (N_8405,N_4514,N_5369);
and U8406 (N_8406,N_7109,N_7649);
nand U8407 (N_8407,N_6426,N_6917);
xnor U8408 (N_8408,N_7988,N_5532);
nor U8409 (N_8409,N_6452,N_6229);
nor U8410 (N_8410,N_6341,N_5734);
or U8411 (N_8411,N_4925,N_4627);
or U8412 (N_8412,N_7207,N_6533);
or U8413 (N_8413,N_4430,N_6163);
xnor U8414 (N_8414,N_5937,N_6639);
xnor U8415 (N_8415,N_4114,N_5672);
xor U8416 (N_8416,N_4701,N_7608);
xor U8417 (N_8417,N_7243,N_6414);
and U8418 (N_8418,N_5875,N_6251);
xnor U8419 (N_8419,N_7332,N_7516);
nor U8420 (N_8420,N_6339,N_4942);
and U8421 (N_8421,N_6285,N_6754);
nor U8422 (N_8422,N_4107,N_7512);
and U8423 (N_8423,N_5342,N_6925);
and U8424 (N_8424,N_6615,N_4340);
and U8425 (N_8425,N_5948,N_6438);
nand U8426 (N_8426,N_4496,N_5346);
xor U8427 (N_8427,N_6231,N_6838);
xnor U8428 (N_8428,N_4511,N_7753);
xnor U8429 (N_8429,N_7657,N_7260);
or U8430 (N_8430,N_4560,N_6133);
or U8431 (N_8431,N_4630,N_6062);
nand U8432 (N_8432,N_5793,N_7742);
xnor U8433 (N_8433,N_5655,N_4664);
nor U8434 (N_8434,N_7060,N_7831);
xor U8435 (N_8435,N_6109,N_4247);
or U8436 (N_8436,N_6447,N_6130);
xnor U8437 (N_8437,N_6671,N_5888);
and U8438 (N_8438,N_7541,N_7264);
or U8439 (N_8439,N_5654,N_7408);
xor U8440 (N_8440,N_5401,N_4982);
or U8441 (N_8441,N_5310,N_7568);
nand U8442 (N_8442,N_5422,N_4779);
or U8443 (N_8443,N_4658,N_6813);
xnor U8444 (N_8444,N_7695,N_6046);
or U8445 (N_8445,N_5900,N_4418);
nor U8446 (N_8446,N_7103,N_4148);
or U8447 (N_8447,N_4605,N_7075);
nand U8448 (N_8448,N_6148,N_6896);
nand U8449 (N_8449,N_4996,N_4190);
or U8450 (N_8450,N_6548,N_5631);
and U8451 (N_8451,N_5169,N_6207);
and U8452 (N_8452,N_4898,N_5432);
nor U8453 (N_8453,N_6389,N_7485);
nand U8454 (N_8454,N_5095,N_5495);
xnor U8455 (N_8455,N_4188,N_4460);
nand U8456 (N_8456,N_4075,N_6350);
and U8457 (N_8457,N_5407,N_7577);
or U8458 (N_8458,N_6985,N_4240);
xnor U8459 (N_8459,N_5384,N_5872);
nand U8460 (N_8460,N_5748,N_7239);
xor U8461 (N_8461,N_5947,N_7230);
or U8462 (N_8462,N_5136,N_4139);
nor U8463 (N_8463,N_5022,N_7047);
nand U8464 (N_8464,N_5663,N_7364);
nor U8465 (N_8465,N_6517,N_7450);
nor U8466 (N_8466,N_5664,N_7844);
or U8467 (N_8467,N_5211,N_6559);
xnor U8468 (N_8468,N_5196,N_5528);
xor U8469 (N_8469,N_4261,N_5012);
and U8470 (N_8470,N_5971,N_4976);
xnor U8471 (N_8471,N_7303,N_5628);
xor U8472 (N_8472,N_4577,N_4196);
and U8473 (N_8473,N_6573,N_7138);
nor U8474 (N_8474,N_4842,N_7735);
nand U8475 (N_8475,N_5621,N_7121);
nor U8476 (N_8476,N_7267,N_4095);
nand U8477 (N_8477,N_4788,N_7850);
and U8478 (N_8478,N_5501,N_4694);
nor U8479 (N_8479,N_4131,N_4348);
nor U8480 (N_8480,N_7328,N_4760);
xor U8481 (N_8481,N_5477,N_5676);
or U8482 (N_8482,N_4786,N_6607);
or U8483 (N_8483,N_6971,N_6624);
xnor U8484 (N_8484,N_5541,N_6802);
nand U8485 (N_8485,N_5419,N_4854);
and U8486 (N_8486,N_7929,N_6564);
xnor U8487 (N_8487,N_7342,N_7044);
or U8488 (N_8488,N_5670,N_5789);
and U8489 (N_8489,N_6305,N_5002);
and U8490 (N_8490,N_4233,N_6198);
xnor U8491 (N_8491,N_5294,N_5982);
xor U8492 (N_8492,N_5704,N_5581);
xor U8493 (N_8493,N_6597,N_6038);
nand U8494 (N_8494,N_4212,N_6226);
xor U8495 (N_8495,N_5094,N_6423);
or U8496 (N_8496,N_4071,N_4088);
xnor U8497 (N_8497,N_4334,N_7569);
nor U8498 (N_8498,N_4454,N_7771);
nand U8499 (N_8499,N_7845,N_4705);
or U8500 (N_8500,N_4391,N_5368);
or U8501 (N_8501,N_7791,N_5990);
xor U8502 (N_8502,N_6578,N_7981);
and U8503 (N_8503,N_5509,N_7345);
nor U8504 (N_8504,N_4413,N_4239);
nand U8505 (N_8505,N_4921,N_6125);
or U8506 (N_8506,N_6715,N_7949);
or U8507 (N_8507,N_5984,N_5956);
nor U8508 (N_8508,N_6012,N_4999);
nand U8509 (N_8509,N_6566,N_4688);
nor U8510 (N_8510,N_7639,N_7145);
and U8511 (N_8511,N_4038,N_7349);
xor U8512 (N_8512,N_5879,N_6120);
or U8513 (N_8513,N_6902,N_6224);
and U8514 (N_8514,N_6964,N_7565);
or U8515 (N_8515,N_7458,N_4197);
xnor U8516 (N_8516,N_7102,N_7240);
xor U8517 (N_8517,N_7816,N_5903);
or U8518 (N_8518,N_6913,N_5423);
and U8519 (N_8519,N_5743,N_5756);
and U8520 (N_8520,N_7499,N_4633);
nor U8521 (N_8521,N_6180,N_6893);
xnor U8522 (N_8522,N_5117,N_7370);
or U8523 (N_8523,N_4226,N_5414);
and U8524 (N_8524,N_5375,N_6342);
nand U8525 (N_8525,N_5869,N_6208);
xnor U8526 (N_8526,N_7994,N_4255);
or U8527 (N_8527,N_5128,N_4297);
and U8528 (N_8528,N_7263,N_4635);
nand U8529 (N_8529,N_6308,N_7781);
xnor U8530 (N_8530,N_6129,N_6110);
and U8531 (N_8531,N_5312,N_6791);
and U8532 (N_8532,N_7813,N_7703);
nand U8533 (N_8533,N_6390,N_4979);
or U8534 (N_8534,N_4693,N_5431);
nor U8535 (N_8535,N_5593,N_6076);
xnor U8536 (N_8536,N_7315,N_6629);
or U8537 (N_8537,N_6905,N_7736);
or U8538 (N_8538,N_7869,N_6023);
or U8539 (N_8539,N_5427,N_5615);
and U8540 (N_8540,N_5720,N_7236);
nor U8541 (N_8541,N_4989,N_5300);
nand U8542 (N_8542,N_6482,N_6126);
or U8543 (N_8543,N_7547,N_7225);
and U8544 (N_8544,N_4858,N_6022);
or U8545 (N_8545,N_6982,N_7043);
nand U8546 (N_8546,N_7838,N_7827);
and U8547 (N_8547,N_4890,N_6973);
and U8548 (N_8548,N_6193,N_5933);
and U8549 (N_8549,N_4267,N_4736);
nand U8550 (N_8550,N_6974,N_5728);
and U8551 (N_8551,N_7707,N_4220);
or U8552 (N_8552,N_5771,N_4118);
nand U8553 (N_8553,N_7941,N_5928);
xor U8554 (N_8554,N_5485,N_4331);
xnor U8555 (N_8555,N_4973,N_4957);
and U8556 (N_8556,N_6580,N_4759);
nor U8557 (N_8557,N_7035,N_6553);
nand U8558 (N_8558,N_6009,N_4234);
nor U8559 (N_8559,N_5634,N_5584);
or U8560 (N_8560,N_6606,N_7158);
nand U8561 (N_8561,N_5440,N_4054);
nand U8562 (N_8562,N_4264,N_7053);
or U8563 (N_8563,N_4477,N_4590);
or U8564 (N_8564,N_4662,N_7728);
and U8565 (N_8565,N_5608,N_5142);
nor U8566 (N_8566,N_5805,N_6381);
nand U8567 (N_8567,N_7588,N_5218);
nand U8568 (N_8568,N_5764,N_6279);
and U8569 (N_8569,N_7976,N_5361);
xnor U8570 (N_8570,N_4532,N_6631);
xnor U8571 (N_8571,N_4035,N_7418);
nand U8572 (N_8572,N_7000,N_5235);
and U8573 (N_8573,N_5377,N_6987);
nand U8574 (N_8574,N_5107,N_7510);
nor U8575 (N_8575,N_7504,N_5345);
xor U8576 (N_8576,N_5472,N_6456);
nor U8577 (N_8577,N_7745,N_6219);
and U8578 (N_8578,N_6689,N_4256);
nor U8579 (N_8579,N_7486,N_5054);
xor U8580 (N_8580,N_7543,N_7597);
nor U8581 (N_8581,N_5647,N_5574);
nor U8582 (N_8582,N_6535,N_7391);
nor U8583 (N_8583,N_4562,N_4944);
nor U8584 (N_8584,N_6576,N_4295);
and U8585 (N_8585,N_7081,N_7519);
xor U8586 (N_8586,N_6498,N_4422);
nand U8587 (N_8587,N_4203,N_6096);
nand U8588 (N_8588,N_6124,N_5570);
xor U8589 (N_8589,N_6944,N_6830);
nor U8590 (N_8590,N_6365,N_6291);
xor U8591 (N_8591,N_7760,N_6314);
nor U8592 (N_8592,N_5695,N_7214);
and U8593 (N_8593,N_6503,N_4787);
and U8594 (N_8594,N_4823,N_4178);
and U8595 (N_8595,N_7355,N_5932);
xnor U8596 (N_8596,N_5320,N_4816);
nor U8597 (N_8597,N_4500,N_6036);
nor U8598 (N_8598,N_5455,N_4362);
nand U8599 (N_8599,N_4329,N_5731);
or U8600 (N_8600,N_4238,N_7550);
and U8601 (N_8601,N_4242,N_5060);
nand U8602 (N_8602,N_4530,N_7298);
nor U8603 (N_8603,N_4154,N_4952);
nor U8604 (N_8604,N_7208,N_7222);
nor U8605 (N_8605,N_6138,N_4283);
nand U8606 (N_8606,N_4346,N_4009);
nand U8607 (N_8607,N_5511,N_4536);
xnor U8608 (N_8608,N_6068,N_7815);
and U8609 (N_8609,N_4849,N_6673);
or U8610 (N_8610,N_4856,N_7310);
xnor U8611 (N_8611,N_6500,N_5540);
and U8612 (N_8612,N_5679,N_7029);
nand U8613 (N_8613,N_5358,N_6000);
xor U8614 (N_8614,N_5809,N_5349);
xnor U8615 (N_8615,N_5891,N_4914);
nand U8616 (N_8616,N_5803,N_6839);
or U8617 (N_8617,N_4013,N_6264);
nor U8618 (N_8618,N_4850,N_7699);
xnor U8619 (N_8619,N_5580,N_6713);
or U8620 (N_8620,N_5160,N_4244);
xor U8621 (N_8621,N_4014,N_4510);
or U8622 (N_8622,N_6083,N_7273);
nand U8623 (N_8623,N_5383,N_4449);
nor U8624 (N_8624,N_6441,N_6204);
and U8625 (N_8625,N_5617,N_4558);
or U8626 (N_8626,N_5352,N_7718);
and U8627 (N_8627,N_6092,N_4882);
or U8628 (N_8628,N_4273,N_4315);
xnor U8629 (N_8629,N_7335,N_4503);
xnor U8630 (N_8630,N_6909,N_5659);
or U8631 (N_8631,N_6525,N_4744);
xnor U8632 (N_8632,N_6609,N_7766);
and U8633 (N_8633,N_6691,N_4335);
xor U8634 (N_8634,N_4845,N_7823);
and U8635 (N_8635,N_6168,N_5381);
or U8636 (N_8636,N_7169,N_4301);
and U8637 (N_8637,N_7573,N_7561);
xnor U8638 (N_8638,N_5573,N_7576);
or U8639 (N_8639,N_6189,N_5821);
and U8640 (N_8640,N_5248,N_4001);
xnor U8641 (N_8641,N_4336,N_6474);
nor U8642 (N_8642,N_6906,N_4909);
or U8643 (N_8643,N_5927,N_5757);
and U8644 (N_8644,N_5446,N_5270);
or U8645 (N_8645,N_7968,N_7134);
nand U8646 (N_8646,N_7659,N_6998);
nor U8647 (N_8647,N_5127,N_4580);
xor U8648 (N_8648,N_6412,N_4392);
or U8649 (N_8649,N_4918,N_5827);
nand U8650 (N_8650,N_7524,N_6127);
nor U8651 (N_8651,N_4539,N_4185);
xnor U8652 (N_8652,N_4978,N_6721);
and U8653 (N_8653,N_4863,N_7533);
xnor U8654 (N_8654,N_4735,N_4908);
or U8655 (N_8655,N_7995,N_7506);
nor U8656 (N_8656,N_4271,N_7817);
nand U8657 (N_8657,N_7302,N_5951);
or U8658 (N_8658,N_7799,N_7586);
and U8659 (N_8659,N_6371,N_7552);
nor U8660 (N_8660,N_5627,N_6886);
nor U8661 (N_8661,N_6620,N_6486);
xor U8662 (N_8662,N_7902,N_6661);
and U8663 (N_8663,N_7435,N_5864);
nor U8664 (N_8664,N_5644,N_5321);
and U8665 (N_8665,N_7532,N_4617);
and U8666 (N_8666,N_7846,N_4083);
nand U8667 (N_8667,N_4084,N_7164);
nor U8668 (N_8668,N_7877,N_7206);
and U8669 (N_8669,N_5281,N_5084);
nor U8670 (N_8670,N_6228,N_6014);
nand U8671 (N_8671,N_6995,N_7768);
xnor U8672 (N_8672,N_6766,N_6611);
nand U8673 (N_8673,N_7339,N_6055);
or U8674 (N_8674,N_5476,N_7891);
nand U8675 (N_8675,N_5851,N_6234);
or U8676 (N_8676,N_4920,N_4132);
xnor U8677 (N_8677,N_6959,N_6879);
nor U8678 (N_8678,N_4517,N_4195);
nor U8679 (N_8679,N_5591,N_7039);
nand U8680 (N_8680,N_4519,N_5832);
or U8681 (N_8681,N_7362,N_6428);
nand U8682 (N_8682,N_5899,N_7226);
and U8683 (N_8683,N_7394,N_7738);
nor U8684 (N_8684,N_5760,N_4099);
and U8685 (N_8685,N_5625,N_4166);
or U8686 (N_8686,N_6066,N_7078);
or U8687 (N_8687,N_4010,N_5001);
xor U8688 (N_8688,N_5518,N_4752);
nor U8689 (N_8689,N_4296,N_7256);
nand U8690 (N_8690,N_6323,N_6434);
xor U8691 (N_8691,N_4028,N_5961);
nor U8692 (N_8692,N_7865,N_7923);
nand U8693 (N_8693,N_7481,N_4481);
or U8694 (N_8694,N_7221,N_4395);
xor U8695 (N_8695,N_5735,N_5645);
and U8696 (N_8696,N_5996,N_7381);
nand U8697 (N_8697,N_4955,N_6112);
or U8698 (N_8698,N_7915,N_6461);
and U8699 (N_8699,N_5430,N_6049);
nor U8700 (N_8700,N_7253,N_4900);
nor U8701 (N_8701,N_7205,N_5061);
and U8702 (N_8702,N_7195,N_7539);
or U8703 (N_8703,N_5914,N_5208);
xnor U8704 (N_8704,N_4260,N_5304);
nand U8705 (N_8705,N_7700,N_5699);
nand U8706 (N_8706,N_6737,N_6884);
nor U8707 (N_8707,N_6514,N_6005);
xnor U8708 (N_8708,N_7009,N_4177);
xnor U8709 (N_8709,N_6455,N_4783);
and U8710 (N_8710,N_6327,N_4444);
and U8711 (N_8711,N_5614,N_6961);
and U8712 (N_8712,N_6955,N_5336);
nor U8713 (N_8713,N_7849,N_5464);
nor U8714 (N_8714,N_7384,N_7407);
nand U8715 (N_8715,N_6064,N_5269);
or U8716 (N_8716,N_4970,N_5134);
or U8717 (N_8717,N_5639,N_5163);
nand U8718 (N_8718,N_4512,N_7276);
or U8719 (N_8719,N_4210,N_7689);
xor U8720 (N_8720,N_7830,N_4116);
nand U8721 (N_8721,N_6379,N_4871);
nand U8722 (N_8722,N_6919,N_5590);
or U8723 (N_8723,N_4465,N_6374);
xor U8724 (N_8724,N_5802,N_6849);
nand U8725 (N_8725,N_7187,N_6507);
nand U8726 (N_8726,N_6824,N_5831);
nor U8727 (N_8727,N_7560,N_7648);
and U8728 (N_8728,N_7036,N_4737);
and U8729 (N_8729,N_6976,N_6045);
nand U8730 (N_8730,N_7669,N_5758);
xnor U8731 (N_8731,N_6495,N_5533);
or U8732 (N_8732,N_5082,N_4838);
nand U8733 (N_8733,N_4289,N_7076);
xor U8734 (N_8734,N_7475,N_6688);
nor U8735 (N_8735,N_5356,N_6928);
nor U8736 (N_8736,N_5326,N_4164);
xor U8737 (N_8737,N_7403,N_4111);
xnor U8738 (N_8738,N_5715,N_4092);
nand U8739 (N_8739,N_6888,N_4358);
nor U8740 (N_8740,N_5069,N_4773);
nor U8741 (N_8741,N_5016,N_7065);
nor U8742 (N_8742,N_7872,N_6044);
nor U8743 (N_8743,N_5025,N_5791);
nor U8744 (N_8744,N_7594,N_6039);
or U8745 (N_8745,N_5935,N_7701);
xnor U8746 (N_8746,N_4940,N_6274);
nor U8747 (N_8747,N_7354,N_7644);
nor U8748 (N_8748,N_6859,N_6940);
or U8749 (N_8749,N_4080,N_4294);
or U8750 (N_8750,N_6122,N_4272);
nor U8751 (N_8751,N_6662,N_6269);
and U8752 (N_8752,N_5380,N_6930);
nor U8753 (N_8753,N_5409,N_6164);
nor U8754 (N_8754,N_4910,N_5165);
or U8755 (N_8755,N_6035,N_7242);
xnor U8756 (N_8756,N_7974,N_4314);
nor U8757 (N_8757,N_7847,N_6993);
and U8758 (N_8758,N_4645,N_7074);
and U8759 (N_8759,N_5979,N_5607);
or U8760 (N_8760,N_6100,N_6949);
nand U8761 (N_8761,N_6774,N_6729);
xnor U8762 (N_8762,N_6344,N_4995);
or U8763 (N_8763,N_6284,N_7279);
and U8764 (N_8764,N_4966,N_4913);
xnor U8765 (N_8765,N_4322,N_5113);
or U8766 (N_8766,N_7715,N_5190);
xnor U8767 (N_8767,N_5986,N_6440);
nor U8768 (N_8768,N_6780,N_7993);
nand U8769 (N_8769,N_6287,N_6183);
or U8770 (N_8770,N_4990,N_7017);
xor U8771 (N_8771,N_6636,N_4262);
nor U8772 (N_8772,N_6782,N_7472);
xor U8773 (N_8773,N_7038,N_5386);
or U8774 (N_8774,N_7477,N_6410);
nand U8775 (N_8775,N_4963,N_6115);
nor U8776 (N_8776,N_6034,N_4874);
xor U8777 (N_8777,N_5456,N_6772);
nand U8778 (N_8778,N_4201,N_5074);
nor U8779 (N_8779,N_6259,N_6747);
and U8780 (N_8780,N_5878,N_4404);
xor U8781 (N_8781,N_5076,N_4061);
nor U8782 (N_8782,N_5398,N_6776);
nor U8783 (N_8783,N_4363,N_7025);
nand U8784 (N_8784,N_4706,N_4021);
nand U8785 (N_8785,N_4259,N_6304);
or U8786 (N_8786,N_6722,N_4709);
and U8787 (N_8787,N_6340,N_7605);
xnor U8788 (N_8788,N_4343,N_5080);
or U8789 (N_8789,N_5156,N_4834);
xnor U8790 (N_8790,N_5007,N_7191);
nor U8791 (N_8791,N_4126,N_6575);
nand U8792 (N_8792,N_6382,N_6085);
xnor U8793 (N_8793,N_5768,N_4872);
nand U8794 (N_8794,N_6093,N_6493);
nand U8795 (N_8795,N_6684,N_4984);
or U8796 (N_8796,N_7023,N_6470);
and U8797 (N_8797,N_6816,N_4451);
nor U8798 (N_8798,N_4258,N_7911);
or U8799 (N_8799,N_6939,N_7320);
nand U8800 (N_8800,N_4864,N_4112);
nand U8801 (N_8801,N_5867,N_4008);
or U8802 (N_8802,N_7962,N_5497);
xor U8803 (N_8803,N_7710,N_4527);
nor U8804 (N_8804,N_7603,N_6788);
or U8805 (N_8805,N_5598,N_6063);
and U8806 (N_8806,N_7369,N_5578);
and U8807 (N_8807,N_6663,N_7175);
nor U8808 (N_8808,N_4988,N_5118);
or U8809 (N_8809,N_5153,N_5228);
xnor U8810 (N_8810,N_4768,N_5690);
nand U8811 (N_8811,N_4687,N_7572);
and U8812 (N_8812,N_5752,N_5692);
and U8813 (N_8813,N_5597,N_4450);
nand U8814 (N_8814,N_4967,N_4589);
xor U8815 (N_8815,N_5261,N_5981);
xnor U8816 (N_8816,N_5066,N_5883);
or U8817 (N_8817,N_4812,N_5711);
and U8818 (N_8818,N_4653,N_6173);
nand U8819 (N_8819,N_4548,N_5051);
nand U8820 (N_8820,N_5957,N_5534);
or U8821 (N_8821,N_5077,N_6679);
and U8822 (N_8822,N_6185,N_7003);
or U8823 (N_8823,N_4003,N_6073);
and U8824 (N_8824,N_6236,N_5335);
xnor U8825 (N_8825,N_6988,N_4386);
xor U8826 (N_8826,N_4149,N_5343);
nor U8827 (N_8827,N_4005,N_5245);
xor U8828 (N_8828,N_5362,N_4525);
and U8829 (N_8829,N_5026,N_6579);
xor U8830 (N_8830,N_4179,N_6577);
xnor U8831 (N_8831,N_4821,N_7062);
or U8832 (N_8832,N_4133,N_4862);
nor U8833 (N_8833,N_4676,N_4721);
nand U8834 (N_8834,N_4426,N_7385);
and U8835 (N_8835,N_4423,N_7997);
xor U8836 (N_8836,N_4011,N_5317);
nor U8837 (N_8837,N_4915,N_4928);
or U8838 (N_8838,N_5613,N_4742);
xor U8839 (N_8839,N_5998,N_6313);
and U8840 (N_8840,N_6822,N_7119);
nand U8841 (N_8841,N_5818,N_5955);
nand U8842 (N_8842,N_7908,N_7917);
nor U8843 (N_8843,N_7143,N_5462);
or U8844 (N_8844,N_7151,N_7963);
nand U8845 (N_8845,N_7518,N_4410);
or U8846 (N_8846,N_5668,N_5862);
nor U8847 (N_8847,N_4089,N_6328);
xor U8848 (N_8848,N_7106,N_6847);
or U8849 (N_8849,N_4235,N_7085);
or U8850 (N_8850,N_6311,N_4373);
nand U8851 (N_8851,N_5049,N_7507);
xor U8852 (N_8852,N_7808,N_4537);
nand U8853 (N_8853,N_4873,N_6714);
nor U8854 (N_8854,N_6852,N_5959);
xnor U8855 (N_8855,N_7204,N_5855);
xor U8856 (N_8856,N_4603,N_4564);
nor U8857 (N_8857,N_6912,N_6199);
or U8858 (N_8858,N_6105,N_5594);
xnor U8859 (N_8859,N_7037,N_6836);
and U8860 (N_8860,N_7999,N_6398);
and U8861 (N_8861,N_6610,N_7757);
xnor U8862 (N_8862,N_4470,N_4529);
or U8863 (N_8863,N_7014,N_6540);
and U8864 (N_8864,N_4145,N_4499);
nor U8865 (N_8865,N_7809,N_5745);
and U8866 (N_8866,N_7013,N_7800);
and U8867 (N_8867,N_4591,N_7542);
nand U8868 (N_8868,N_4464,N_6811);
nand U8869 (N_8869,N_6155,N_7094);
and U8870 (N_8870,N_7146,N_5370);
xnor U8871 (N_8871,N_6154,N_6111);
nor U8872 (N_8872,N_4648,N_7415);
or U8873 (N_8873,N_7708,N_4594);
and U8874 (N_8874,N_7784,N_7655);
nor U8875 (N_8875,N_5296,N_6429);
nor U8876 (N_8876,N_5922,N_4180);
or U8877 (N_8877,N_4796,N_5085);
nor U8878 (N_8878,N_5896,N_6329);
nor U8879 (N_8879,N_4302,N_7245);
and U8880 (N_8880,N_7057,N_5604);
xor U8881 (N_8881,N_5277,N_7805);
or U8882 (N_8882,N_7904,N_5194);
nor U8883 (N_8883,N_7957,N_4288);
nor U8884 (N_8884,N_5151,N_6319);
xnor U8885 (N_8885,N_7471,N_4685);
and U8886 (N_8886,N_7513,N_4526);
nand U8887 (N_8887,N_7517,N_7591);
and U8888 (N_8888,N_6258,N_6724);
or U8889 (N_8889,N_5736,N_4403);
and U8890 (N_8890,N_5841,N_6355);
nand U8891 (N_8891,N_7998,N_4069);
xnor U8892 (N_8892,N_5055,N_5576);
xor U8893 (N_8893,N_4714,N_5817);
xor U8894 (N_8894,N_7666,N_4308);
nor U8895 (N_8895,N_6856,N_7255);
and U8896 (N_8896,N_4293,N_4198);
nand U8897 (N_8897,N_6001,N_5686);
nand U8898 (N_8898,N_7688,N_4716);
or U8899 (N_8899,N_6808,N_7897);
xor U8900 (N_8900,N_5727,N_5893);
nor U8901 (N_8901,N_7558,N_7031);
xor U8902 (N_8902,N_5493,N_5293);
or U8903 (N_8903,N_6205,N_6770);
and U8904 (N_8904,N_5989,N_5033);
nand U8905 (N_8905,N_7104,N_6664);
nand U8906 (N_8906,N_4087,N_7227);
nand U8907 (N_8907,N_7373,N_6666);
nor U8908 (N_8908,N_5230,N_5747);
or U8909 (N_8909,N_5642,N_6677);
and U8910 (N_8910,N_6763,N_6885);
nor U8911 (N_8911,N_7867,N_7672);
or U8912 (N_8912,N_4478,N_6950);
nand U8913 (N_8913,N_7788,N_6152);
nor U8914 (N_8914,N_5402,N_4082);
nand U8915 (N_8915,N_6239,N_5997);
and U8916 (N_8916,N_7420,N_7934);
or U8917 (N_8917,N_5040,N_6360);
nor U8918 (N_8918,N_5172,N_6727);
nor U8919 (N_8919,N_4534,N_5207);
xor U8920 (N_8920,N_5008,N_6376);
or U8921 (N_8921,N_4528,N_4901);
and U8922 (N_8922,N_7898,N_4542);
and U8923 (N_8923,N_7436,N_4162);
nor U8924 (N_8924,N_5366,N_7785);
or U8925 (N_8925,N_7180,N_5301);
nor U8926 (N_8926,N_7905,N_7709);
xor U8927 (N_8927,N_5812,N_5983);
xor U8928 (N_8928,N_5483,N_6927);
or U8929 (N_8929,N_7258,N_4802);
xnor U8930 (N_8930,N_4184,N_5778);
nor U8931 (N_8931,N_7113,N_7080);
xor U8932 (N_8932,N_4602,N_4473);
nand U8933 (N_8933,N_4280,N_6040);
or U8934 (N_8934,N_5514,N_6196);
xnor U8935 (N_8935,N_6735,N_5712);
or U8936 (N_8936,N_6848,N_4696);
or U8937 (N_8937,N_7163,N_4490);
and U8938 (N_8938,N_7600,N_7615);
and U8939 (N_8939,N_6765,N_7828);
or U8940 (N_8940,N_4828,N_6268);
or U8941 (N_8941,N_6512,N_4625);
or U8942 (N_8942,N_5014,N_7224);
nand U8943 (N_8943,N_5611,N_4457);
and U8944 (N_8944,N_4202,N_5297);
or U8945 (N_8945,N_4217,N_7250);
and U8946 (N_8946,N_5777,N_5649);
nor U8947 (N_8947,N_5500,N_4351);
nand U8948 (N_8948,N_5359,N_6192);
nand U8949 (N_8949,N_7019,N_4584);
nand U8950 (N_8950,N_4467,N_7953);
nand U8951 (N_8951,N_4620,N_6756);
nor U8952 (N_8952,N_6230,N_7620);
and U8953 (N_8953,N_4877,N_6102);
nand U8954 (N_8954,N_6052,N_5457);
nand U8955 (N_8955,N_5609,N_5622);
nor U8956 (N_8956,N_4286,N_4943);
nor U8957 (N_8957,N_4187,N_5537);
nand U8958 (N_8958,N_7032,N_6942);
nor U8959 (N_8959,N_5941,N_6617);
and U8960 (N_8960,N_6868,N_6352);
nor U8961 (N_8961,N_4892,N_7182);
xnor U8962 (N_8962,N_7702,N_5588);
or U8963 (N_8963,N_7640,N_6843);
or U8964 (N_8964,N_7170,N_6899);
nand U8965 (N_8965,N_4585,N_7045);
nand U8966 (N_8966,N_6792,N_4936);
or U8967 (N_8967,N_7398,N_4700);
nor U8968 (N_8968,N_5071,N_5917);
nor U8969 (N_8969,N_5960,N_5299);
nor U8970 (N_8970,N_7463,N_4686);
or U8971 (N_8971,N_4567,N_7130);
nor U8972 (N_8972,N_5479,N_7285);
nor U8973 (N_8973,N_6712,N_5314);
or U8974 (N_8974,N_5181,N_4431);
or U8975 (N_8975,N_5527,N_4129);
and U8976 (N_8976,N_6829,N_6373);
nor U8977 (N_8977,N_5776,N_7698);
or U8978 (N_8978,N_4652,N_7737);
xnor U8979 (N_8979,N_6405,N_4253);
and U8980 (N_8980,N_5141,N_4657);
nand U8981 (N_8981,N_4062,N_5129);
nor U8982 (N_8982,N_6136,N_5334);
nand U8983 (N_8983,N_6777,N_4339);
xor U8984 (N_8984,N_7546,N_5999);
nand U8985 (N_8985,N_6524,N_5081);
and U8986 (N_8986,N_5673,N_4777);
nand U8987 (N_8987,N_5282,N_5371);
xnor U8988 (N_8988,N_5863,N_4337);
xor U8989 (N_8989,N_7883,N_6711);
nor U8990 (N_8990,N_6471,N_4566);
xnor U8991 (N_8991,N_4690,N_4971);
xnor U8992 (N_8992,N_7535,N_6442);
xnor U8993 (N_8993,N_4266,N_4274);
nand U8994 (N_8994,N_5525,N_5660);
xor U8995 (N_8995,N_4429,N_5292);
and U8996 (N_8996,N_6718,N_7909);
or U8997 (N_8997,N_7361,N_6527);
xor U8998 (N_8998,N_6941,N_4110);
xor U8999 (N_8999,N_7114,N_7824);
nand U9000 (N_9000,N_6243,N_7832);
xor U9001 (N_9001,N_4036,N_7647);
or U9002 (N_9002,N_4360,N_6733);
nor U9003 (N_9003,N_6002,N_7251);
nand U9004 (N_9004,N_6011,N_5606);
and U9005 (N_9005,N_6432,N_4218);
and U9006 (N_9006,N_6656,N_6400);
xor U9007 (N_9007,N_6123,N_4833);
or U9008 (N_9008,N_5624,N_5633);
xnor U9009 (N_9009,N_5555,N_6402);
nand U9010 (N_9010,N_4626,N_4583);
xor U9011 (N_9011,N_5123,N_5944);
or U9012 (N_9012,N_4025,N_6866);
and U9013 (N_9013,N_5637,N_7177);
xor U9014 (N_9014,N_5765,N_5435);
or U9015 (N_9015,N_7257,N_6375);
nor U9016 (N_9016,N_4613,N_5018);
nor U9017 (N_9017,N_6855,N_6087);
or U9018 (N_9018,N_4610,N_7806);
xnor U9019 (N_9019,N_4052,N_7124);
and U9020 (N_9020,N_6630,N_7282);
and U9021 (N_9021,N_7498,N_7357);
or U9022 (N_9022,N_6842,N_7112);
xnor U9023 (N_9023,N_6458,N_4876);
xor U9024 (N_9024,N_5461,N_5020);
or U9025 (N_9025,N_5295,N_6562);
nor U9026 (N_9026,N_4309,N_5429);
xor U9027 (N_9027,N_5950,N_6744);
nand U9028 (N_9028,N_5652,N_6290);
nand U9029 (N_9029,N_6312,N_7201);
and U9030 (N_9030,N_7168,N_6582);
nand U9031 (N_9031,N_7969,N_7070);
nor U9032 (N_9032,N_6543,N_4804);
and U9033 (N_9033,N_7144,N_5372);
nor U9034 (N_9034,N_6153,N_5305);
or U9035 (N_9035,N_4436,N_7117);
nor U9036 (N_9036,N_4891,N_5303);
nor U9037 (N_9037,N_5097,N_6516);
or U9038 (N_9038,N_5554,N_7105);
or U9039 (N_9039,N_7860,N_6396);
and U9040 (N_9040,N_7066,N_6016);
nor U9041 (N_9041,N_4161,N_4043);
and U9042 (N_9042,N_4764,N_4031);
and U9043 (N_9043,N_6059,N_6276);
and U9044 (N_9044,N_6084,N_4044);
nor U9045 (N_9045,N_4809,N_4552);
nand U9046 (N_9046,N_5562,N_5694);
and U9047 (N_9047,N_6216,N_5188);
or U9048 (N_9048,N_4547,N_7740);
nor U9049 (N_9049,N_4819,N_5939);
nand U9050 (N_9050,N_4619,N_7271);
nand U9051 (N_9051,N_4387,N_6485);
nor U9052 (N_9052,N_4851,N_6556);
nand U9053 (N_9053,N_7571,N_5072);
nor U9054 (N_9054,N_6672,N_6932);
or U9055 (N_9055,N_7623,N_6574);
and U9056 (N_9056,N_5693,N_5186);
xor U9057 (N_9057,N_7209,N_6041);
and U9058 (N_9058,N_4060,N_7939);
or U9059 (N_9059,N_6283,N_4565);
nand U9060 (N_9060,N_5671,N_6370);
xor U9061 (N_9061,N_5242,N_5897);
nor U9062 (N_9062,N_5357,N_4923);
xnor U9063 (N_9063,N_5421,N_4810);
xnor U9064 (N_9064,N_6921,N_4406);
nand U9065 (N_9065,N_6861,N_7599);
xor U9066 (N_9066,N_6869,N_5238);
nand U9067 (N_9067,N_7413,N_6139);
xnor U9068 (N_9068,N_4587,N_6567);
xnor U9069 (N_9069,N_6336,N_5434);
or U9070 (N_9070,N_6716,N_6448);
nor U9071 (N_9071,N_5360,N_4746);
xnor U9072 (N_9072,N_7022,N_4119);
nand U9073 (N_9073,N_7093,N_4466);
nor U9074 (N_9074,N_4829,N_5042);
nor U9075 (N_9075,N_4672,N_5560);
xor U9076 (N_9076,N_7947,N_4986);
or U9077 (N_9077,N_5449,N_6741);
nor U9078 (N_9078,N_5037,N_6378);
nand U9079 (N_9079,N_5138,N_4776);
nand U9080 (N_9080,N_5058,N_4798);
nand U9081 (N_9081,N_4806,N_5769);
xnor U9082 (N_9082,N_5665,N_4433);
nor U9083 (N_9083,N_7091,N_6594);
or U9084 (N_9084,N_4946,N_4579);
nor U9085 (N_9085,N_4338,N_5219);
or U9086 (N_9086,N_5750,N_7326);
nor U9087 (N_9087,N_7492,N_5612);
or U9088 (N_9088,N_5962,N_6281);
xor U9089 (N_9089,N_7287,N_5391);
or U9090 (N_9090,N_6627,N_6924);
xnor U9091 (N_9091,N_5873,N_4434);
and U9092 (N_9092,N_7556,N_7755);
nor U9093 (N_9093,N_5258,N_4000);
or U9094 (N_9094,N_4448,N_5243);
and U9095 (N_9095,N_5972,N_6506);
and U9096 (N_9096,N_4582,N_6821);
or U9097 (N_9097,N_7527,N_6409);
nor U9098 (N_9098,N_4077,N_7618);
and U9099 (N_9099,N_6277,N_5632);
nand U9100 (N_9100,N_5993,N_5319);
nor U9101 (N_9101,N_4353,N_6764);
xnor U9102 (N_9102,N_4292,N_4730);
nand U9103 (N_9103,N_7523,N_5884);
and U9104 (N_9104,N_7580,N_5102);
nor U9105 (N_9105,N_4839,N_4097);
nand U9106 (N_9106,N_4848,N_4720);
nand U9107 (N_9107,N_5109,N_7538);
or U9108 (N_9108,N_7274,N_6563);
xor U9109 (N_9109,N_6761,N_5041);
or U9110 (N_9110,N_6330,N_4115);
nand U9111 (N_9111,N_7460,N_6242);
xor U9112 (N_9112,N_6171,N_4040);
nor U9113 (N_9113,N_6201,N_7858);
nand U9114 (N_9114,N_6757,N_4896);
nand U9115 (N_9115,N_4754,N_5404);
and U9116 (N_9116,N_6191,N_4604);
nor U9117 (N_9117,N_5623,N_7213);
nand U9118 (N_9118,N_5619,N_5744);
nand U9119 (N_9119,N_6484,N_7589);
and U9120 (N_9120,N_6145,N_6300);
and U9121 (N_9121,N_6367,N_6787);
nor U9122 (N_9122,N_7374,N_6621);
nand U9123 (N_9123,N_5602,N_5722);
nor U9124 (N_9124,N_7153,N_5452);
or U9125 (N_9125,N_7697,N_6167);
nand U9126 (N_9126,N_4934,N_5408);
or U9127 (N_9127,N_7596,N_4432);
and U9128 (N_9128,N_6392,N_4769);
xnor U9129 (N_9129,N_6873,N_6700);
nand U9130 (N_9130,N_7020,N_4588);
and U9131 (N_9131,N_6692,N_6024);
xor U9132 (N_9132,N_6748,N_6908);
xnor U9133 (N_9133,N_6326,N_4157);
nor U9134 (N_9134,N_5491,N_7575);
nor U9135 (N_9135,N_7462,N_4125);
xor U9136 (N_9136,N_7663,N_5000);
and U9137 (N_9137,N_6349,N_7982);
and U9138 (N_9138,N_5130,N_7943);
and U9139 (N_9139,N_6646,N_7984);
xor U9140 (N_9140,N_7127,N_6003);
xor U9141 (N_9141,N_4612,N_7290);
nand U9142 (N_9142,N_6990,N_6008);
and U9143 (N_9143,N_4551,N_7001);
nor U9144 (N_9144,N_6244,N_5233);
nor U9145 (N_9145,N_4105,N_5412);
xor U9146 (N_9146,N_4058,N_4134);
and U9147 (N_9147,N_4347,N_7125);
or U9148 (N_9148,N_7996,N_5994);
or U9149 (N_9149,N_4880,N_6551);
or U9150 (N_9150,N_6415,N_5098);
xor U9151 (N_9151,N_5494,N_7063);
or U9152 (N_9152,N_7765,N_5365);
or U9153 (N_9153,N_7894,N_4749);
and U9154 (N_9154,N_7284,N_5909);
nand U9155 (N_9155,N_6401,N_4949);
nor U9156 (N_9156,N_7181,N_5967);
nand U9157 (N_9157,N_6775,N_4956);
nand U9158 (N_9158,N_7247,N_7028);
xnor U9159 (N_9159,N_6321,N_6612);
and U9160 (N_9160,N_7338,N_4352);
and U9161 (N_9161,N_4428,N_7167);
and U9162 (N_9162,N_7004,N_6521);
nand U9163 (N_9163,N_4342,N_7223);
and U9164 (N_9164,N_7021,N_5753);
nand U9165 (N_9165,N_6749,N_6221);
nand U9166 (N_9166,N_7252,N_5988);
nor U9167 (N_9167,N_4886,N_7313);
nor U9168 (N_9168,N_7383,N_5086);
nand U9169 (N_9169,N_4600,N_4684);
nand U9170 (N_9170,N_6812,N_5859);
nand U9171 (N_9171,N_5895,N_4555);
xor U9172 (N_9172,N_4541,N_6529);
nand U9173 (N_9173,N_6074,N_4782);
and U9174 (N_9174,N_7810,N_4425);
nor U9175 (N_9175,N_5232,N_4817);
and U9176 (N_9176,N_5148,N_6523);
or U9177 (N_9177,N_5638,N_6253);
nor U9178 (N_9178,N_7682,N_5746);
nand U9179 (N_9179,N_4414,N_7174);
and U9180 (N_9180,N_4894,N_6571);
xor U9181 (N_9181,N_5059,N_7862);
xnor U9182 (N_9182,N_7884,N_6687);
and U9183 (N_9183,N_6760,N_6841);
xor U9184 (N_9184,N_7333,N_7234);
or U9185 (N_9185,N_7566,N_7650);
xor U9186 (N_9186,N_5226,N_6918);
nor U9187 (N_9187,N_7980,N_4435);
xor U9188 (N_9188,N_6526,N_6298);
or U9189 (N_9189,N_4727,N_5507);
and U9190 (N_9190,N_5565,N_6608);
nand U9191 (N_9191,N_7675,N_7767);
xor U9192 (N_9192,N_4159,N_4878);
and U9193 (N_9193,N_6292,N_5730);
nand U9194 (N_9194,N_4761,N_7880);
xnor U9195 (N_9195,N_7438,N_5741);
xor U9196 (N_9196,N_4544,N_6509);
nor U9197 (N_9197,N_4556,N_7196);
or U9198 (N_9198,N_7693,N_5915);
nor U9199 (N_9199,N_4616,N_7814);
nand U9200 (N_9200,N_6202,N_4607);
xor U9201 (N_9201,N_7761,N_6019);
and U9202 (N_9202,N_6951,N_7405);
xnor U9203 (N_9203,N_5273,N_4455);
nand U9204 (N_9204,N_7752,N_6870);
nand U9205 (N_9205,N_6660,N_5641);
nand U9206 (N_9206,N_5618,N_5236);
and U9207 (N_9207,N_7317,N_6858);
and U9208 (N_9208,N_7190,N_4174);
nand U9209 (N_9209,N_7068,N_6176);
nor U9210 (N_9210,N_4595,N_4784);
nand U9211 (N_9211,N_4330,N_4056);
or U9212 (N_9212,N_7197,N_5610);
nor U9213 (N_9213,N_6149,N_7631);
xor U9214 (N_9214,N_5199,N_5546);
or U9215 (N_9215,N_5592,N_7514);
and U9216 (N_9216,N_7629,N_5726);
nand U9217 (N_9217,N_7272,N_6318);
nor U9218 (N_9218,N_6368,N_7839);
nand U9219 (N_9219,N_7979,N_5868);
xor U9220 (N_9220,N_6785,N_6773);
xnor U9221 (N_9221,N_4229,N_6017);
or U9222 (N_9222,N_6723,N_6653);
xnor U9223 (N_9223,N_4546,N_4553);
or U9224 (N_9224,N_4461,N_5837);
nor U9225 (N_9225,N_5379,N_5087);
nand U9226 (N_9226,N_4237,N_7007);
or U9227 (N_9227,N_4906,N_7652);
nand U9228 (N_9228,N_6817,N_5487);
nand U9229 (N_9229,N_4550,N_7216);
and U9230 (N_9230,N_7212,N_4670);
xnor U9231 (N_9231,N_6417,N_4163);
and U9232 (N_9232,N_7930,N_4447);
nor U9233 (N_9233,N_6459,N_6659);
nand U9234 (N_9234,N_4808,N_4325);
or U9235 (N_9235,N_5389,N_6616);
nand U9236 (N_9236,N_7421,N_5835);
or U9237 (N_9237,N_5834,N_5176);
xnor U9238 (N_9238,N_5877,N_5683);
nor U9239 (N_9239,N_4324,N_5339);
or U9240 (N_9240,N_5125,N_6121);
nor U9241 (N_9241,N_5963,N_6364);
nor U9242 (N_9242,N_7136,N_7360);
xor U9243 (N_9243,N_5424,N_7149);
xnor U9244 (N_9244,N_7874,N_4168);
or U9245 (N_9245,N_5131,N_5200);
xnor U9246 (N_9246,N_6586,N_4487);
nor U9247 (N_9247,N_7977,N_5006);
and U9248 (N_9248,N_5330,N_4729);
xnor U9249 (N_9249,N_5820,N_6255);
or U9250 (N_9250,N_5448,N_4269);
or U9251 (N_9251,N_5991,N_5437);
or U9252 (N_9252,N_7837,N_4427);
or U9253 (N_9253,N_6837,N_7363);
and U9254 (N_9254,N_5926,N_6675);
or U9255 (N_9255,N_7126,N_6698);
xor U9256 (N_9256,N_4747,N_5460);
nor U9257 (N_9257,N_5385,N_4400);
xor U9258 (N_9258,N_5521,N_5530);
and U9259 (N_9259,N_4355,N_6408);
and U9260 (N_9260,N_7836,N_5259);
and U9261 (N_9261,N_7607,N_7563);
or U9262 (N_9262,N_5965,N_5159);
xor U9263 (N_9263,N_4183,N_4070);
or U9264 (N_9264,N_4932,N_5137);
xnor U9265 (N_9265,N_6351,N_4919);
nand U9266 (N_9266,N_5949,N_5341);
nor U9267 (N_9267,N_6430,N_6416);
or U9268 (N_9268,N_6246,N_6280);
and U9269 (N_9269,N_6860,N_7966);
or U9270 (N_9270,N_5616,N_6048);
nor U9271 (N_9271,N_5987,N_4707);
or U9272 (N_9272,N_6750,N_4937);
nor U9273 (N_9273,N_7323,N_7154);
nand U9274 (N_9274,N_4677,N_5144);
nor U9275 (N_9275,N_6174,N_7590);
xor U9276 (N_9276,N_4800,N_5589);
or U9277 (N_9277,N_5023,N_7536);
nand U9278 (N_9278,N_5108,N_7763);
nand U9279 (N_9279,N_6645,N_5719);
xor U9280 (N_9280,N_5969,N_5564);
and U9281 (N_9281,N_6572,N_7653);
or U9282 (N_9282,N_6203,N_7095);
xor U9283 (N_9283,N_5814,N_5975);
and U9284 (N_9284,N_4969,N_4538);
nand U9285 (N_9285,N_4855,N_5503);
nor U9286 (N_9286,N_7932,N_7353);
nand U9287 (N_9287,N_4983,N_4811);
nand U9288 (N_9288,N_6965,N_4889);
or U9289 (N_9289,N_4279,N_6317);
nor U9290 (N_9290,N_5738,N_7330);
and U9291 (N_9291,N_7726,N_5441);
xor U9292 (N_9292,N_4922,N_4926);
or U9293 (N_9293,N_6728,N_4715);
nor U9294 (N_9294,N_4189,N_4545);
xor U9295 (N_9295,N_4093,N_5122);
nand U9296 (N_9296,N_4245,N_6027);
and U9297 (N_9297,N_7612,N_6874);
nand U9298 (N_9298,N_5203,N_4221);
nand U9299 (N_9299,N_5415,N_7793);
nor U9300 (N_9300,N_4987,N_7634);
nand U9301 (N_9301,N_7681,N_6649);
nor U9302 (N_9302,N_7026,N_4227);
xnor U9303 (N_9303,N_7992,N_4725);
and U9304 (N_9304,N_5829,N_4192);
and U9305 (N_9305,N_5505,N_4822);
and U9306 (N_9306,N_5083,N_6851);
nor U9307 (N_9307,N_5451,N_4076);
nor U9308 (N_9308,N_5954,N_6981);
nand U9309 (N_9309,N_6238,N_5822);
xor U9310 (N_9310,N_5481,N_5773);
or U9311 (N_9311,N_7916,N_5454);
nand U9312 (N_9312,N_4369,N_4282);
nor U9313 (N_9313,N_6235,N_7107);
or U9314 (N_9314,N_7173,N_7684);
nor U9315 (N_9315,N_5600,N_5351);
nor U9316 (N_9316,N_7564,N_5662);
xor U9317 (N_9317,N_4650,N_4958);
nor U9318 (N_9318,N_5475,N_6369);
or U9319 (N_9319,N_7432,N_7101);
and U9320 (N_9320,N_5177,N_7762);
or U9321 (N_9321,N_7959,N_6876);
nor U9322 (N_9322,N_4057,N_4100);
or U9323 (N_9323,N_4902,N_4767);
and U9324 (N_9324,N_7325,N_7440);
nand U9325 (N_9325,N_5698,N_7090);
xnor U9326 (N_9326,N_5725,N_4497);
nor U9327 (N_9327,N_6413,N_7097);
nor U9328 (N_9328,N_5502,N_5189);
and U9329 (N_9329,N_4305,N_6395);
nand U9330 (N_9330,N_6978,N_6103);
and U9331 (N_9331,N_7474,N_4636);
and U9332 (N_9332,N_5438,N_6681);
and U9333 (N_9333,N_5348,N_7404);
nor U9334 (N_9334,N_4899,N_5550);
or U9335 (N_9335,N_5100,N_7249);
nor U9336 (N_9336,N_7491,N_6054);
and U9337 (N_9337,N_7217,N_4361);
and U9338 (N_9338,N_7365,N_5754);
nor U9339 (N_9339,N_6169,N_5043);
or U9340 (N_9340,N_4327,N_5308);
or U9341 (N_9341,N_4389,N_4143);
nand U9342 (N_9342,N_7306,N_6827);
xor U9343 (N_9343,N_7885,N_4985);
nor U9344 (N_9344,N_5073,N_7324);
or U9345 (N_9345,N_6783,N_4938);
xor U9346 (N_9346,N_4795,N_6655);
xnor U9347 (N_9347,N_5388,N_5111);
nand U9348 (N_9348,N_7079,N_6947);
xor U9349 (N_9349,N_5376,N_4771);
and U9350 (N_9350,N_7444,N_6460);
and U9351 (N_9351,N_4276,N_4907);
nor U9352 (N_9352,N_6050,N_6831);
nand U9353 (N_9353,N_4208,N_6968);
xor U9354 (N_9354,N_5680,N_4859);
nand U9355 (N_9355,N_7525,N_5149);
nand U9356 (N_9356,N_6676,N_5973);
or U9357 (N_9357,N_5173,N_6751);
nand U9358 (N_9358,N_7744,N_5795);
nand U9359 (N_9359,N_7179,N_4954);
nand U9360 (N_9360,N_4303,N_4442);
nand U9361 (N_9361,N_6635,N_4814);
xnor U9362 (N_9362,N_7476,N_4865);
nand U9363 (N_9363,N_7914,N_4135);
nand U9364 (N_9364,N_5938,N_5241);
or U9365 (N_9365,N_7712,N_4622);
xnor U9366 (N_9366,N_4109,N_5904);
or U9367 (N_9367,N_4250,N_5572);
nand U9368 (N_9368,N_6322,N_6213);
xor U9369 (N_9369,N_4634,N_4520);
nand U9370 (N_9370,N_7218,N_4756);
xnor U9371 (N_9371,N_5702,N_7537);
or U9372 (N_9372,N_5036,N_5465);
and U9373 (N_9373,N_7776,N_7470);
nand U9374 (N_9374,N_4576,N_5063);
or U9375 (N_9375,N_6962,N_7705);
and U9376 (N_9376,N_5093,N_5635);
xnor U9377 (N_9377,N_4774,N_7008);
or U9378 (N_9378,N_7848,N_7322);
and U9379 (N_9379,N_6804,N_6480);
or U9380 (N_9380,N_5044,N_6850);
nor U9381 (N_9381,N_7308,N_7613);
nor U9382 (N_9382,N_7797,N_7775);
nand U9383 (N_9383,N_6265,N_6887);
nor U9384 (N_9384,N_6384,N_6147);
and U9385 (N_9385,N_5586,N_6945);
or U9386 (N_9386,N_4504,N_6179);
nand U9387 (N_9387,N_6481,N_6963);
nand U9388 (N_9388,N_7010,N_6004);
nor U9389 (N_9389,N_6131,N_7268);
or U9390 (N_9390,N_4643,N_6310);
and U9391 (N_9391,N_7454,N_5906);
nand U9392 (N_9392,N_4826,N_7423);
and U9393 (N_9393,N_4586,N_6222);
xnor U9394 (N_9394,N_6372,N_6864);
nand U9395 (N_9395,N_4027,N_4870);
nor U9396 (N_9396,N_5936,N_5840);
or U9397 (N_9397,N_4666,N_4408);
nand U9398 (N_9398,N_7975,N_4837);
and U9399 (N_9399,N_7445,N_7643);
nand U9400 (N_9400,N_5516,N_6538);
and U9401 (N_9401,N_4176,N_7925);
nor U9402 (N_9402,N_7056,N_7448);
xor U9403 (N_9403,N_6755,N_4831);
nor U9404 (N_9404,N_5510,N_7910);
nand U9405 (N_9405,N_7551,N_7803);
nand U9406 (N_9406,N_6051,N_5090);
xnor U9407 (N_9407,N_5306,N_4313);
nand U9408 (N_9408,N_6719,N_5700);
nor U9409 (N_9409,N_6431,N_7329);
nor U9410 (N_9410,N_6953,N_4844);
nand U9411 (N_9411,N_6795,N_5543);
or U9412 (N_9412,N_7084,N_7439);
xnor U9413 (N_9413,N_6025,N_7387);
xor U9414 (N_9414,N_5482,N_5164);
nand U9415 (N_9415,N_4318,N_5116);
nor U9416 (N_9416,N_5929,N_4748);
nor U9417 (N_9417,N_7292,N_6508);
xnor U9418 (N_9418,N_4965,N_6786);
and U9419 (N_9419,N_6547,N_6361);
nand U9420 (N_9420,N_6053,N_7835);
or U9421 (N_9421,N_4384,N_4041);
nand U9422 (N_9422,N_5911,N_6335);
or U9423 (N_9423,N_7172,N_7099);
or U9424 (N_9424,N_5889,N_5830);
xnor U9425 (N_9425,N_5167,N_6638);
nand U9426 (N_9426,N_6897,N_5824);
xnor U9427 (N_9427,N_6273,N_7729);
and U9428 (N_9428,N_4738,N_5213);
nor U9429 (N_9429,N_7683,N_6797);
xnor U9430 (N_9430,N_4524,N_7786);
nor U9431 (N_9431,N_7139,N_6404);
and U9432 (N_9432,N_5332,N_4241);
and U9433 (N_9433,N_7270,N_6446);
nor U9434 (N_9434,N_4875,N_6091);
xnor U9435 (N_9435,N_4402,N_4508);
nor U9436 (N_9436,N_7417,N_6491);
and U9437 (N_9437,N_5646,N_5224);
or U9438 (N_9438,N_7892,N_7350);
xnor U9439 (N_9439,N_7352,N_6810);
and U9440 (N_9440,N_7128,N_6853);
nand U9441 (N_9441,N_4743,N_5701);
and U9442 (N_9442,N_7312,N_5459);
nand U9443 (N_9443,N_5088,N_7895);
xnor U9444 (N_9444,N_4191,N_7262);
and U9445 (N_9445,N_4469,N_5836);
or U9446 (N_9446,N_4997,N_7334);
nor U9447 (N_9447,N_6425,N_4841);
nor U9448 (N_9448,N_6613,N_5417);
or U9449 (N_9449,N_7203,N_7351);
and U9450 (N_9450,N_4117,N_4569);
or U9451 (N_9451,N_6165,N_5221);
nor U9452 (N_9452,N_6465,N_7961);
xnor U9453 (N_9453,N_7295,N_6892);
nor U9454 (N_9454,N_6550,N_6297);
nand U9455 (N_9455,N_4034,N_7857);
or U9456 (N_9456,N_5174,N_7487);
xor U9457 (N_9457,N_6241,N_5819);
nor U9458 (N_9458,N_7617,N_5101);
nand U9459 (N_9459,N_5065,N_4068);
nor U9460 (N_9460,N_4789,N_6674);
and U9461 (N_9461,N_5716,N_5150);
nor U9462 (N_9462,N_5547,N_6454);
nand U9463 (N_9463,N_5825,N_5354);
or U9464 (N_9464,N_6762,N_5667);
xor U9465 (N_9465,N_4689,N_7780);
nor U9466 (N_9466,N_4765,N_4475);
and U9467 (N_9467,N_6282,N_5684);
xnor U9468 (N_9468,N_6444,N_5029);
nor U9469 (N_9469,N_5682,N_7521);
or U9470 (N_9470,N_6732,N_4055);
nand U9471 (N_9471,N_7157,N_7764);
or U9472 (N_9472,N_6622,N_6271);
xnor U9473 (N_9473,N_5266,N_4780);
or U9474 (N_9474,N_4170,N_7722);
nand U9475 (N_9475,N_4710,N_6994);
nand U9476 (N_9476,N_7842,N_6515);
xor U9477 (N_9477,N_4206,N_7244);
or U9478 (N_9478,N_5559,N_6333);
xor U9479 (N_9479,N_5217,N_4805);
and U9480 (N_9480,N_7955,N_7382);
xnor U9481 (N_9481,N_5763,N_7443);
nor U9482 (N_9482,N_6178,N_4711);
nor U9483 (N_9483,N_7110,N_7371);
or U9484 (N_9484,N_5813,N_6560);
nor U9485 (N_9485,N_5737,N_7900);
or U9486 (N_9486,N_6492,N_4249);
nor U9487 (N_9487,N_4857,N_6590);
xor U9488 (N_9488,N_4090,N_6840);
and U9489 (N_9489,N_4820,N_6451);
and U9490 (N_9490,N_6536,N_5918);
nand U9491 (N_9491,N_6013,N_6132);
or U9492 (N_9492,N_6895,N_5436);
and U9493 (N_9493,N_4211,N_4624);
xor U9494 (N_9494,N_6079,N_7851);
or U9495 (N_9495,N_5222,N_4354);
xor U9496 (N_9496,N_4045,N_4136);
or U9497 (N_9497,N_6522,N_5183);
xnor U9498 (N_9498,N_6225,N_7390);
nand U9499 (N_9499,N_6345,N_7451);
nand U9500 (N_9500,N_6826,N_7082);
xor U9501 (N_9501,N_4049,N_5237);
nor U9502 (N_9502,N_7508,N_4629);
nand U9503 (N_9503,N_7919,N_6669);
xnor U9504 (N_9504,N_4770,N_7340);
and U9505 (N_9505,N_6558,N_7156);
nand U9506 (N_9506,N_6534,N_4151);
xor U9507 (N_9507,N_7088,N_7841);
and U9508 (N_9508,N_7802,N_6833);
nor U9509 (N_9509,N_4306,N_5193);
xor U9510 (N_9510,N_6863,N_6784);
and U9511 (N_9511,N_5724,N_6286);
xor U9512 (N_9512,N_5794,N_5400);
nand U9513 (N_9513,N_6510,N_7581);
nor U9514 (N_9514,N_6220,N_6599);
and U9515 (N_9515,N_7899,N_5799);
and U9516 (N_9516,N_5162,N_5531);
or U9517 (N_9517,N_7275,N_4417);
or U9518 (N_9518,N_5124,N_7141);
or U9519 (N_9519,N_7906,N_7936);
nand U9520 (N_9520,N_7165,N_7940);
xnor U9521 (N_9521,N_6901,N_7456);
nand U9522 (N_9522,N_7054,N_6796);
nor U9523 (N_9523,N_5880,N_5104);
nand U9524 (N_9524,N_7484,N_6391);
and U9525 (N_9525,N_5302,N_5523);
or U9526 (N_9526,N_7375,N_4251);
and U9527 (N_9527,N_7779,N_4981);
and U9528 (N_9528,N_6678,N_4398);
or U9529 (N_9529,N_7359,N_5197);
nand U9530 (N_9530,N_7933,N_5839);
nor U9531 (N_9531,N_7948,N_7116);
or U9532 (N_9532,N_4462,N_4554);
nor U9533 (N_9533,N_5675,N_7118);
and U9534 (N_9534,N_4285,N_6343);
nor U9535 (N_9535,N_6151,N_5313);
nand U9536 (N_9536,N_7235,N_5152);
and U9537 (N_9537,N_5992,N_4815);
nand U9538 (N_9538,N_6072,N_4416);
nand U9539 (N_9539,N_7237,N_7453);
and U9540 (N_9540,N_4252,N_5519);
nand U9541 (N_9541,N_7431,N_4656);
nand U9542 (N_9542,N_6742,N_4766);
and U9543 (N_9543,N_5804,N_5844);
or U9544 (N_9544,N_7719,N_7876);
xnor U9545 (N_9545,N_4463,N_6497);
xor U9546 (N_9546,N_6141,N_5471);
and U9547 (N_9547,N_6815,N_7301);
nand U9548 (N_9548,N_6875,N_5175);
and U9549 (N_9549,N_5857,N_7046);
nor U9550 (N_9550,N_5782,N_7692);
xnor U9551 (N_9551,N_7727,N_6668);
nand U9552 (N_9552,N_7840,N_5139);
or U9553 (N_9553,N_7960,N_5549);
nand U9554 (N_9554,N_5807,N_7680);
xnor U9555 (N_9555,N_7426,N_4860);
and U9556 (N_9556,N_4173,N_5626);
or U9557 (N_9557,N_4674,N_7467);
and U9558 (N_9558,N_4601,N_5333);
or U9559 (N_9559,N_5373,N_5833);
xnor U9560 (N_9560,N_4407,N_5871);
and U9561 (N_9561,N_6031,N_7526);
xnor U9562 (N_9562,N_4931,N_7089);
nor U9563 (N_9563,N_7389,N_4263);
xnor U9564 (N_9564,N_7812,N_6232);
and U9565 (N_9565,N_6803,N_5143);
nor U9566 (N_9566,N_6667,N_7717);
or U9567 (N_9567,N_4310,N_6647);
xnor U9568 (N_9568,N_7896,N_5187);
and U9569 (N_9569,N_4228,N_6591);
nand U9570 (N_9570,N_5274,N_5657);
xor U9571 (N_9571,N_7171,N_4142);
nand U9572 (N_9572,N_5272,N_5426);
and U9573 (N_9573,N_7664,N_7574);
and U9574 (N_9574,N_4568,N_7228);
nand U9575 (N_9575,N_5034,N_7133);
nor U9576 (N_9576,N_5157,N_7430);
or U9577 (N_9577,N_7870,N_6097);
xnor U9578 (N_9578,N_4278,N_6952);
xnor U9579 (N_9579,N_7720,N_6694);
nand U9580 (N_9580,N_5558,N_5595);
xor U9581 (N_9581,N_4939,N_6146);
xnor U9582 (N_9582,N_6682,N_4113);
nor U9583 (N_9583,N_5522,N_6463);
nor U9584 (N_9584,N_4364,N_6618);
and U9585 (N_9585,N_7051,N_4493);
nor U9586 (N_9586,N_7327,N_4794);
xor U9587 (N_9587,N_7927,N_4646);
xor U9588 (N_9588,N_5198,N_5751);
nor U9589 (N_9589,N_4682,N_5328);
and U9590 (N_9590,N_4681,N_5953);
nor U9591 (N_9591,N_4270,N_4728);
xnor U9592 (N_9592,N_7198,N_7395);
nand U9593 (N_9593,N_7942,N_7690);
or U9594 (N_9594,N_6581,N_5416);
xnor U9595 (N_9595,N_7829,N_4039);
and U9596 (N_9596,N_5854,N_5964);
nand U9597 (N_9597,N_5696,N_6740);
nor U9598 (N_9598,N_4376,N_4853);
xor U9599 (N_9599,N_7579,N_6670);
nand U9600 (N_9600,N_4399,N_5285);
xnor U9601 (N_9601,N_4772,N_5453);
xnor U9602 (N_9602,N_6302,N_6358);
xnor U9603 (N_9603,N_6513,N_5828);
nand U9604 (N_9604,N_5410,N_7593);
and U9605 (N_9605,N_6172,N_4916);
or U9606 (N_9606,N_5024,N_5010);
nand U9607 (N_9607,N_6487,N_6197);
nor U9608 (N_9608,N_5050,N_5064);
or U9609 (N_9609,N_7782,N_7473);
nand U9610 (N_9610,N_4230,N_6476);
or U9611 (N_9611,N_6637,N_4223);
xnor U9612 (N_9612,N_7465,N_5329);
xnor U9613 (N_9613,N_7396,N_7679);
nand U9614 (N_9614,N_5155,N_5905);
nor U9615 (N_9615,N_5046,N_4121);
and U9616 (N_9616,N_4483,N_4004);
xor U9617 (N_9617,N_6814,N_5508);
xnor U9618 (N_9618,N_7077,N_4679);
xor U9619 (N_9619,N_7611,N_5688);
nor U9620 (N_9620,N_7464,N_4509);
and U9621 (N_9621,N_7215,N_5520);
xor U9622 (N_9622,N_6690,N_4344);
xnor U9623 (N_9623,N_5478,N_4719);
nand U9624 (N_9624,N_4169,N_5575);
nand U9625 (N_9625,N_7529,N_7347);
nand U9626 (N_9626,N_7871,N_6212);
xnor U9627 (N_9627,N_7411,N_7482);
nand U9628 (N_9628,N_4533,N_7592);
nor U9629 (N_9629,N_5009,N_5552);
or U9630 (N_9630,N_5488,N_4375);
and U9631 (N_9631,N_6709,N_4480);
and U9632 (N_9632,N_4651,N_7277);
and U9633 (N_9633,N_7220,N_5787);
and U9634 (N_9634,N_6449,N_7219);
xor U9635 (N_9635,N_7490,N_5770);
xor U9636 (N_9636,N_4128,N_7283);
nand U9637 (N_9637,N_7654,N_6403);
nand U9638 (N_9638,N_5374,N_4775);
nor U9639 (N_9639,N_4801,N_7723);
and U9640 (N_9640,N_5331,N_7964);
nand U9641 (N_9641,N_6614,N_4290);
xor U9642 (N_9642,N_7494,N_4390);
and U9643 (N_9643,N_6862,N_7734);
nor U9644 (N_9644,N_5974,N_7807);
xnor U9645 (N_9645,N_4214,N_6267);
nor U9646 (N_9646,N_7628,N_4521);
xnor U9647 (N_9647,N_7015,N_7048);
xor U9648 (N_9648,N_6980,N_6794);
nand U9649 (N_9649,N_4535,N_7311);
xor U9650 (N_9650,N_6010,N_7878);
and U9651 (N_9651,N_5115,N_5732);
or U9652 (N_9652,N_4371,N_6696);
xor U9653 (N_9653,N_4064,N_4945);
or U9654 (N_9654,N_5585,N_5934);
and U9655 (N_9655,N_6938,N_7651);
nor U9656 (N_9656,N_4219,N_7058);
or U9657 (N_9657,N_4103,N_5425);
or U9658 (N_9658,N_5253,N_4437);
and U9659 (N_9659,N_4443,N_6047);
xnor U9660 (N_9660,N_4578,N_7555);
nand U9661 (N_9661,N_4152,N_6081);
nor U9662 (N_9662,N_7049,N_5120);
or U9663 (N_9663,N_5866,N_4171);
nand U9664 (N_9664,N_7621,N_7570);
nand U9665 (N_9665,N_4867,N_7553);
nand U9666 (N_9666,N_5135,N_4722);
nand U9667 (N_9667,N_7072,N_7912);
nand U9668 (N_9668,N_5908,N_5916);
nand U9669 (N_9669,N_5816,N_7238);
xnor U9670 (N_9670,N_7466,N_6357);
or U9671 (N_9671,N_6758,N_4827);
xnor U9672 (N_9672,N_5251,N_7505);
and U9673 (N_9673,N_4930,N_7120);
xnor U9674 (N_9674,N_5529,N_4224);
or U9675 (N_9675,N_4453,N_6717);
and U9676 (N_9676,N_6693,N_6779);
xor U9677 (N_9677,N_7630,N_7142);
nand U9678 (N_9678,N_7200,N_4704);
nand U9679 (N_9679,N_5930,N_4059);
and U9680 (N_9680,N_7668,N_4708);
nand U9681 (N_9681,N_5256,N_5057);
and U9682 (N_9682,N_4345,N_6240);
and U9683 (N_9683,N_4102,N_7794);
xor U9684 (N_9684,N_5105,N_5126);
and U9685 (N_9685,N_7636,N_7265);
or U9686 (N_9686,N_5068,N_7160);
xnor U9687 (N_9687,N_4415,N_6736);
and U9688 (N_9688,N_4623,N_5636);
nor U9689 (N_9689,N_5307,N_5168);
or U9690 (N_9690,N_7750,N_6261);
and U9691 (N_9691,N_7856,N_6477);
nand U9692 (N_9692,N_6730,N_7549);
and U9693 (N_9693,N_7042,N_7625);
nand U9694 (N_9694,N_7544,N_6632);
and U9695 (N_9695,N_4078,N_5849);
xor U9696 (N_9696,N_4072,N_7331);
or U9697 (N_9697,N_5039,N_4750);
or U9698 (N_9698,N_4611,N_6890);
nor U9699 (N_9699,N_4042,N_7619);
and U9700 (N_9700,N_4883,N_6530);
xor U9701 (N_9701,N_7528,N_5347);
and U9702 (N_9702,N_6037,N_6098);
or U9703 (N_9703,N_7706,N_4140);
nor U9704 (N_9704,N_5394,N_5788);
nand U9705 (N_9705,N_6504,N_6903);
xnor U9706 (N_9706,N_6278,N_5898);
nand U9707 (N_9707,N_6427,N_7677);
xnor U9708 (N_9708,N_6194,N_7286);
and U9709 (N_9709,N_4106,N_6633);
nand U9710 (N_9710,N_6745,N_5913);
xor U9711 (N_9711,N_7972,N_7749);
xor U9712 (N_9712,N_5759,N_7419);
nand U9713 (N_9713,N_4663,N_7150);
and U9714 (N_9714,N_6387,N_7185);
xnor U9715 (N_9715,N_4751,N_4791);
or U9716 (N_9716,N_7321,N_6209);
or U9717 (N_9717,N_7199,N_4370);
nand U9718 (N_9718,N_7554,N_5723);
and U9719 (N_9719,N_4793,N_4287);
and U9720 (N_9720,N_6781,N_6263);
or U9721 (N_9721,N_5640,N_7299);
xor U9722 (N_9722,N_6746,N_7316);
nor U9723 (N_9723,N_6900,N_4868);
nand U9724 (N_9724,N_6086,N_7254);
nand U9725 (N_9725,N_6725,N_5283);
and U9726 (N_9726,N_5092,N_4257);
xor U9727 (N_9727,N_4165,N_5784);
xor U9728 (N_9728,N_7511,N_4101);
nand U9729 (N_9729,N_7186,N_7685);
nor U9730 (N_9730,N_5070,N_7246);
and U9731 (N_9731,N_7368,N_7614);
nand U9732 (N_9732,N_5249,N_7769);
and U9733 (N_9733,N_5216,N_7129);
and U9734 (N_9734,N_4207,N_4964);
nor U9735 (N_9735,N_4243,N_4992);
and U9736 (N_9736,N_4175,N_6818);
nand U9737 (N_9737,N_5876,N_4665);
xnor U9738 (N_9738,N_6114,N_4458);
nor U9739 (N_9739,N_7161,N_6798);
nor U9740 (N_9740,N_5762,N_6651);
or U9741 (N_9741,N_7954,N_5548);
nor U9742 (N_9742,N_7610,N_5846);
nand U9743 (N_9743,N_5439,N_4281);
nand U9744 (N_9744,N_5468,N_5103);
nand U9745 (N_9745,N_5463,N_7414);
nor U9746 (N_9746,N_4147,N_4323);
xor U9747 (N_9747,N_4866,N_5205);
or U9748 (N_9748,N_6704,N_6911);
nand U9749 (N_9749,N_7064,N_7557);
nor U9750 (N_9750,N_4316,N_5924);
or U9751 (N_9751,N_7006,N_4020);
or U9752 (N_9752,N_6984,N_5567);
and U9753 (N_9753,N_7388,N_7166);
nor U9754 (N_9754,N_6057,N_6603);
or U9755 (N_9755,N_4471,N_5147);
xnor U9756 (N_9756,N_5848,N_5557);
nor U9757 (N_9757,N_4079,N_7694);
and U9758 (N_9758,N_4792,N_6969);
or U9759 (N_9759,N_7434,N_6104);
xnor U9760 (N_9760,N_4675,N_6356);
nand U9761 (N_9761,N_6501,N_5309);
nor U9762 (N_9762,N_5387,N_4998);
and U9763 (N_9763,N_6223,N_4439);
and U9764 (N_9764,N_7033,N_4977);
nor U9765 (N_9765,N_5709,N_6359);
xnor U9766 (N_9766,N_5005,N_6904);
or U9767 (N_9767,N_7469,N_4691);
and U9768 (N_9768,N_4718,N_7873);
and U9769 (N_9769,N_7248,N_7096);
nand U9770 (N_9770,N_5721,N_7291);
and U9771 (N_9771,N_4350,N_7493);
and U9772 (N_9772,N_6116,N_7792);
or U9773 (N_9773,N_5185,N_5798);
nand U9774 (N_9774,N_6089,N_4572);
nor U9775 (N_9775,N_4712,N_6366);
nand U9776 (N_9776,N_4494,N_6021);
or U9777 (N_9777,N_5096,N_6363);
or U9778 (N_9778,N_4225,N_4513);
or U9779 (N_9779,N_4446,N_7437);
and U9780 (N_9780,N_4032,N_6587);
or U9781 (N_9781,N_7346,N_7067);
and U9782 (N_9782,N_6738,N_6731);
and U9783 (N_9783,N_5078,N_5601);
nor U9784 (N_9784,N_6094,N_6421);
or U9785 (N_9785,N_5985,N_4724);
and U9786 (N_9786,N_4699,N_4381);
and U9787 (N_9787,N_7777,N_7194);
xnor U9788 (N_9788,N_6845,N_6695);
and U9789 (N_9789,N_7052,N_7123);
xor U9790 (N_9790,N_7424,N_6479);
xnor U9791 (N_9791,N_5995,N_6881);
nor U9792 (N_9792,N_6546,N_4468);
or U9793 (N_9793,N_5133,N_4019);
or U9794 (N_9794,N_4740,N_6200);
nor U9795 (N_9795,N_6077,N_7971);
nor U9796 (N_9796,N_7970,N_5278);
nand U9797 (N_9797,N_7422,N_5091);
nand U9798 (N_9798,N_4067,N_5170);
nor U9799 (N_9799,N_6296,N_6248);
nor U9800 (N_9800,N_7770,N_4960);
nand U9801 (N_9801,N_6101,N_5234);
nand U9802 (N_9802,N_5761,N_7626);
xnor U9803 (N_9803,N_4123,N_5850);
nor U9804 (N_9804,N_5428,N_7790);
nor U9805 (N_9805,N_7261,N_4332);
xnor U9806 (N_9806,N_5244,N_6490);
nor U9807 (N_9807,N_5513,N_7016);
or U9808 (N_9808,N_6210,N_4597);
or U9809 (N_9809,N_4638,N_7030);
xnor U9810 (N_9810,N_7378,N_5856);
and U9811 (N_9811,N_6108,N_5980);
or U9812 (N_9812,N_4200,N_6555);
or U9813 (N_9813,N_6411,N_4824);
nor U9814 (N_9814,N_4349,N_7716);
and U9815 (N_9815,N_6407,N_4063);
nand U9816 (N_9816,N_6878,N_4328);
xnor U9817 (N_9817,N_7921,N_4968);
or U9818 (N_9818,N_5089,N_4540);
nor U9819 (N_9819,N_4401,N_5227);
nor U9820 (N_9820,N_5184,N_7540);
nor U9821 (N_9821,N_7888,N_4216);
xor U9822 (N_9822,N_7725,N_7530);
nor U9823 (N_9823,N_6252,N_7392);
or U9824 (N_9824,N_7913,N_7348);
xor U9825 (N_9825,N_6657,N_4505);
and U9826 (N_9826,N_4482,N_5378);
and U9827 (N_9827,N_5705,N_7193);
or U9828 (N_9828,N_6467,N_4153);
nand U9829 (N_9829,N_7132,N_4484);
and U9830 (N_9830,N_4268,N_4680);
or U9831 (N_9831,N_6589,N_5395);
or U9832 (N_9832,N_7496,N_7344);
nor U9833 (N_9833,N_7005,N_4888);
or U9834 (N_9834,N_5907,N_5603);
and U9835 (N_9835,N_6175,N_5325);
nor U9836 (N_9836,N_5551,N_4098);
and U9837 (N_9837,N_5561,N_7673);
nor U9838 (N_9838,N_5577,N_5405);
nand U9839 (N_9839,N_5469,N_6519);
nor U9840 (N_9840,N_6706,N_6334);
nor U9841 (N_9841,N_7667,N_6585);
nor U9842 (N_9842,N_7406,N_7449);
and U9843 (N_9843,N_7559,N_4518);
and U9844 (N_9844,N_4124,N_5650);
nand U9845 (N_9845,N_7401,N_5053);
or U9846 (N_9846,N_5442,N_7604);
xor U9847 (N_9847,N_7515,N_5853);
xnor U9848 (N_9848,N_5774,N_4723);
nand U9849 (N_9849,N_4474,N_4733);
and U9850 (N_9850,N_6182,N_4758);
and U9851 (N_9851,N_7548,N_7122);
or U9852 (N_9852,N_4778,N_6478);
nand U9853 (N_9853,N_6595,N_7336);
nor U9854 (N_9854,N_4002,N_7189);
or U9855 (N_9855,N_5931,N_4847);
nor U9856 (N_9856,N_7584,N_4637);
nor U9857 (N_9857,N_4606,N_5191);
nand U9858 (N_9858,N_6640,N_7229);
xor U9859 (N_9859,N_6891,N_6643);
nor U9860 (N_9860,N_7304,N_4411);
or U9861 (N_9861,N_4570,N_4951);
and U9862 (N_9862,N_5945,N_6588);
nor U9863 (N_9863,N_6554,N_6544);
xor U9864 (N_9864,N_5447,N_7671);
nor U9865 (N_9865,N_6983,N_6070);
xor U9866 (N_9866,N_7887,N_4840);
nand U9867 (N_9867,N_7393,N_4950);
xor U9868 (N_9868,N_4383,N_6128);
xor U9869 (N_9869,N_7520,N_5268);
xor U9870 (N_9870,N_7034,N_5192);
xnor U9871 (N_9871,N_5286,N_6419);
nand U9872 (N_9872,N_5587,N_5800);
nor U9873 (N_9873,N_6568,N_7965);
and U9874 (N_9874,N_5411,N_5892);
nand U9875 (N_9875,N_5886,N_4621);
and U9876 (N_9876,N_5767,N_5223);
and U9877 (N_9877,N_6080,N_4561);
or U9878 (N_9878,N_4007,N_7184);
nor U9879 (N_9879,N_7711,N_7822);
and U9880 (N_9880,N_4051,N_5443);
or U9881 (N_9881,N_7147,N_6457);
nand U9882 (N_9882,N_4639,N_7480);
and U9883 (N_9883,N_6975,N_6383);
nor U9884 (N_9884,N_5811,N_7804);
xor U9885 (N_9885,N_5045,N_7944);
nor U9886 (N_9886,N_6936,N_6800);
and U9887 (N_9887,N_6771,N_6865);
or U9888 (N_9888,N_5579,N_6867);
and U9889 (N_9889,N_6033,N_4456);
xnor U9890 (N_9890,N_7751,N_7522);
xor U9891 (N_9891,N_4502,N_4172);
or U9892 (N_9892,N_4033,N_5697);
nor U9893 (N_9893,N_5327,N_4753);
xnor U9894 (N_9894,N_5785,N_5079);
nor U9895 (N_9895,N_7410,N_5766);
or U9896 (N_9896,N_5874,N_5749);
and U9897 (N_9897,N_7583,N_7973);
xor U9898 (N_9898,N_4030,N_6916);
or U9899 (N_9899,N_5852,N_5099);
and U9900 (N_9900,N_5209,N_5838);
or U9901 (N_9901,N_4489,N_6823);
or U9902 (N_9902,N_4897,N_4741);
nor U9903 (N_9903,N_5920,N_6170);
and U9904 (N_9904,N_4924,N_4445);
and U9905 (N_9905,N_4086,N_4726);
xor U9906 (N_9906,N_5140,N_4137);
and U9907 (N_9907,N_4120,N_7259);
nand U9908 (N_9908,N_5355,N_6475);
and U9909 (N_9909,N_6703,N_4209);
or U9910 (N_9910,N_4523,N_5894);
or U9911 (N_9911,N_5710,N_4941);
and U9912 (N_9912,N_7140,N_7732);
nand U9913 (N_9913,N_6914,N_7441);
xnor U9914 (N_9914,N_6584,N_7991);
and U9915 (N_9915,N_4186,N_5445);
nor U9916 (N_9916,N_4835,N_7645);
nand U9917 (N_9917,N_5484,N_6469);
nand U9918 (N_9918,N_5182,N_6937);
and U9919 (N_9919,N_4781,N_6472);
xnor U9920 (N_9920,N_5382,N_5706);
xor U9921 (N_9921,N_6685,N_7232);
nand U9922 (N_9922,N_5201,N_5474);
nand U9923 (N_9923,N_6331,N_4254);
xnor U9924 (N_9924,N_6619,N_6520);
xnor U9925 (N_9925,N_6650,N_4807);
nor U9926 (N_9926,N_5942,N_7500);
and U9927 (N_9927,N_6502,N_4393);
and U9928 (N_9928,N_5542,N_5858);
xnor U9929 (N_9929,N_7863,N_7495);
and U9930 (N_9930,N_7946,N_5910);
nor U9931 (N_9931,N_6095,N_7018);
nor U9932 (N_9932,N_4549,N_4832);
or U9933 (N_9933,N_7759,N_6466);
and U9934 (N_9934,N_5504,N_7687);
xor U9935 (N_9935,N_7952,N_6217);
or U9936 (N_9936,N_5019,N_5166);
and U9937 (N_9937,N_4813,N_5367);
nand U9938 (N_9938,N_6157,N_6935);
nand U9939 (N_9939,N_6245,N_4368);
nor U9940 (N_9940,N_4974,N_5052);
or U9941 (N_9941,N_4887,N_4006);
and U9942 (N_9942,N_6162,N_5363);
or U9943 (N_9943,N_6301,N_4745);
or U9944 (N_9944,N_6316,N_4319);
or U9945 (N_9945,N_6394,N_5406);
nand U9946 (N_9946,N_4066,N_7633);
xnor U9947 (N_9947,N_6734,N_7834);
nand U9948 (N_9948,N_4962,N_7601);
nor U9949 (N_9949,N_7622,N_5689);
nor U9950 (N_9950,N_7987,N_6483);
nand U9951 (N_9951,N_6060,N_4018);
or U9952 (N_9952,N_7305,N_6539);
and U9953 (N_9953,N_7582,N_4205);
xnor U9954 (N_9954,N_6844,N_6511);
nand U9955 (N_9955,N_6295,N_5284);
nand U9956 (N_9956,N_7455,N_4420);
or U9957 (N_9957,N_7231,N_6957);
or U9958 (N_9958,N_5923,N_7796);
nand U9959 (N_9959,N_5316,N_5013);
nand U9960 (N_9960,N_6462,N_6134);
and U9961 (N_9961,N_7489,N_7820);
nor U9962 (N_9962,N_6015,N_4017);
xnor U9963 (N_9963,N_4695,N_5506);
or U9964 (N_9964,N_5324,N_5340);
xor U9965 (N_9965,N_6557,N_7833);
xnor U9966 (N_9966,N_6338,N_4321);
and U9967 (N_9967,N_7920,N_5178);
and U9968 (N_9968,N_6986,N_4074);
nor U9969 (N_9969,N_6144,N_4394);
or U9970 (N_9970,N_7595,N_7826);
xor U9971 (N_9971,N_6954,N_7159);
nor U9972 (N_9972,N_4385,N_7427);
nor U9973 (N_9973,N_6029,N_7115);
and U9974 (N_9974,N_5792,N_5535);
and U9975 (N_9975,N_4947,N_7587);
and U9976 (N_9976,N_7950,N_5290);
and U9977 (N_9977,N_4581,N_5718);
nand U9978 (N_9978,N_4731,N_4598);
or U9979 (N_9979,N_4424,N_4929);
and U9980 (N_9980,N_5028,N_4573);
nor U9981 (N_9981,N_5392,N_4531);
nor U9982 (N_9982,N_5318,N_4655);
nand U9983 (N_9983,N_4642,N_7428);
and U9984 (N_9984,N_4911,N_5801);
nand U9985 (N_9985,N_6992,N_5298);
xnor U9986 (N_9986,N_4015,N_5860);
or U9987 (N_9987,N_4647,N_7468);
nor U9988 (N_9988,N_4284,N_6464);
nand U9989 (N_9989,N_5260,N_4732);
nand U9990 (N_9990,N_5783,N_5733);
nand U9991 (N_9991,N_6623,N_7041);
xnor U9992 (N_9992,N_4702,N_6188);
and U9993 (N_9993,N_7893,N_4182);
nand U9994 (N_9994,N_6894,N_6549);
nor U9995 (N_9995,N_4697,N_7011);
or U9996 (N_9996,N_4485,N_7318);
nand U9997 (N_9997,N_6600,N_6806);
or U9998 (N_9998,N_7861,N_5263);
and U9999 (N_9999,N_6726,N_4904);
nor U10000 (N_10000,N_4663,N_6454);
nand U10001 (N_10001,N_5577,N_6688);
nor U10002 (N_10002,N_6803,N_7702);
and U10003 (N_10003,N_5481,N_4526);
nand U10004 (N_10004,N_5283,N_6803);
nand U10005 (N_10005,N_7176,N_4714);
or U10006 (N_10006,N_7732,N_6496);
xor U10007 (N_10007,N_6296,N_6022);
xnor U10008 (N_10008,N_6595,N_4795);
or U10009 (N_10009,N_6692,N_7332);
or U10010 (N_10010,N_5392,N_6282);
and U10011 (N_10011,N_4974,N_5462);
xnor U10012 (N_10012,N_7481,N_6701);
nor U10013 (N_10013,N_6063,N_7164);
nor U10014 (N_10014,N_5233,N_6931);
nor U10015 (N_10015,N_4537,N_6620);
nor U10016 (N_10016,N_4426,N_4957);
nand U10017 (N_10017,N_5548,N_6144);
or U10018 (N_10018,N_4856,N_6186);
and U10019 (N_10019,N_5170,N_4436);
xor U10020 (N_10020,N_4853,N_4077);
nor U10021 (N_10021,N_7773,N_6661);
xnor U10022 (N_10022,N_7984,N_7956);
xor U10023 (N_10023,N_6435,N_7985);
nand U10024 (N_10024,N_4201,N_7577);
xnor U10025 (N_10025,N_7029,N_6089);
xor U10026 (N_10026,N_5630,N_7807);
or U10027 (N_10027,N_6646,N_6845);
nor U10028 (N_10028,N_5421,N_7319);
and U10029 (N_10029,N_5284,N_5330);
nor U10030 (N_10030,N_6572,N_6882);
and U10031 (N_10031,N_5366,N_6706);
nor U10032 (N_10032,N_5881,N_4883);
and U10033 (N_10033,N_5038,N_7013);
xor U10034 (N_10034,N_4934,N_5523);
nor U10035 (N_10035,N_6059,N_7475);
nor U10036 (N_10036,N_5339,N_6120);
and U10037 (N_10037,N_5448,N_7001);
nand U10038 (N_10038,N_7665,N_4957);
xor U10039 (N_10039,N_6908,N_5482);
nor U10040 (N_10040,N_7163,N_4893);
nand U10041 (N_10041,N_7964,N_6329);
xor U10042 (N_10042,N_7354,N_5523);
nor U10043 (N_10043,N_7056,N_5838);
or U10044 (N_10044,N_5813,N_7032);
nand U10045 (N_10045,N_7071,N_5508);
and U10046 (N_10046,N_7673,N_7215);
nand U10047 (N_10047,N_5751,N_4614);
and U10048 (N_10048,N_7889,N_4817);
or U10049 (N_10049,N_7925,N_4706);
xnor U10050 (N_10050,N_5350,N_5759);
and U10051 (N_10051,N_7234,N_7742);
xnor U10052 (N_10052,N_5652,N_7675);
xnor U10053 (N_10053,N_7609,N_6285);
or U10054 (N_10054,N_6600,N_5702);
and U10055 (N_10055,N_6197,N_5879);
or U10056 (N_10056,N_5620,N_6844);
nand U10057 (N_10057,N_6774,N_4958);
nand U10058 (N_10058,N_4907,N_6322);
nor U10059 (N_10059,N_4178,N_6035);
and U10060 (N_10060,N_7809,N_7506);
or U10061 (N_10061,N_6797,N_4498);
nand U10062 (N_10062,N_4548,N_5674);
nand U10063 (N_10063,N_4752,N_6247);
nor U10064 (N_10064,N_6969,N_4622);
and U10065 (N_10065,N_4216,N_6569);
or U10066 (N_10066,N_7394,N_6700);
and U10067 (N_10067,N_6352,N_6610);
nor U10068 (N_10068,N_7630,N_5826);
and U10069 (N_10069,N_6202,N_4261);
nor U10070 (N_10070,N_4344,N_5481);
nor U10071 (N_10071,N_6418,N_5638);
nand U10072 (N_10072,N_7435,N_4680);
xor U10073 (N_10073,N_4127,N_6999);
xnor U10074 (N_10074,N_7690,N_7704);
nand U10075 (N_10075,N_5268,N_4764);
nor U10076 (N_10076,N_5846,N_7530);
and U10077 (N_10077,N_7523,N_6142);
nand U10078 (N_10078,N_6128,N_5048);
nor U10079 (N_10079,N_6221,N_4659);
or U10080 (N_10080,N_5681,N_5068);
or U10081 (N_10081,N_4194,N_4896);
nand U10082 (N_10082,N_5425,N_6688);
and U10083 (N_10083,N_7128,N_5067);
nor U10084 (N_10084,N_4870,N_4303);
xnor U10085 (N_10085,N_5587,N_7378);
xnor U10086 (N_10086,N_7269,N_5352);
nor U10087 (N_10087,N_6527,N_5908);
xnor U10088 (N_10088,N_6528,N_5208);
and U10089 (N_10089,N_4598,N_4344);
nor U10090 (N_10090,N_7866,N_7607);
or U10091 (N_10091,N_5521,N_5465);
nor U10092 (N_10092,N_4267,N_5438);
nand U10093 (N_10093,N_7992,N_6680);
or U10094 (N_10094,N_6407,N_4881);
or U10095 (N_10095,N_4568,N_6510);
nor U10096 (N_10096,N_4767,N_6675);
nand U10097 (N_10097,N_6840,N_5540);
nor U10098 (N_10098,N_5157,N_4881);
and U10099 (N_10099,N_5819,N_7008);
or U10100 (N_10100,N_6893,N_6582);
and U10101 (N_10101,N_4056,N_7986);
nand U10102 (N_10102,N_4249,N_6185);
xnor U10103 (N_10103,N_6604,N_6435);
or U10104 (N_10104,N_7328,N_7409);
and U10105 (N_10105,N_6242,N_4784);
nor U10106 (N_10106,N_6973,N_4880);
nand U10107 (N_10107,N_6716,N_4783);
xnor U10108 (N_10108,N_7633,N_4405);
nor U10109 (N_10109,N_6727,N_5461);
nor U10110 (N_10110,N_7983,N_5106);
nand U10111 (N_10111,N_5929,N_5170);
and U10112 (N_10112,N_4515,N_4123);
nor U10113 (N_10113,N_6463,N_5605);
xor U10114 (N_10114,N_5872,N_6136);
or U10115 (N_10115,N_4165,N_6497);
nand U10116 (N_10116,N_5775,N_5718);
and U10117 (N_10117,N_6343,N_6004);
nor U10118 (N_10118,N_4357,N_5467);
nor U10119 (N_10119,N_6372,N_6694);
or U10120 (N_10120,N_6816,N_4242);
or U10121 (N_10121,N_7389,N_4305);
nor U10122 (N_10122,N_6548,N_7219);
nand U10123 (N_10123,N_7582,N_7512);
and U10124 (N_10124,N_7401,N_5707);
nor U10125 (N_10125,N_5477,N_4046);
or U10126 (N_10126,N_4723,N_4474);
nand U10127 (N_10127,N_5746,N_6460);
nor U10128 (N_10128,N_7570,N_5887);
and U10129 (N_10129,N_4951,N_5592);
and U10130 (N_10130,N_4560,N_4809);
xnor U10131 (N_10131,N_4287,N_6637);
xnor U10132 (N_10132,N_7072,N_7243);
xor U10133 (N_10133,N_5608,N_4619);
nor U10134 (N_10134,N_5179,N_6172);
nor U10135 (N_10135,N_4935,N_4210);
nand U10136 (N_10136,N_4948,N_6242);
nand U10137 (N_10137,N_5509,N_4439);
or U10138 (N_10138,N_7908,N_4424);
or U10139 (N_10139,N_5324,N_7607);
or U10140 (N_10140,N_5717,N_4581);
or U10141 (N_10141,N_6671,N_5228);
and U10142 (N_10142,N_7300,N_6231);
and U10143 (N_10143,N_7387,N_5048);
nand U10144 (N_10144,N_5634,N_7289);
xor U10145 (N_10145,N_5990,N_5348);
xnor U10146 (N_10146,N_5024,N_4032);
xnor U10147 (N_10147,N_6988,N_6416);
and U10148 (N_10148,N_4260,N_6680);
nand U10149 (N_10149,N_6372,N_7216);
xnor U10150 (N_10150,N_4041,N_6113);
or U10151 (N_10151,N_7546,N_5502);
and U10152 (N_10152,N_5330,N_6690);
nand U10153 (N_10153,N_6976,N_4923);
xnor U10154 (N_10154,N_7791,N_5021);
nand U10155 (N_10155,N_4070,N_7054);
nand U10156 (N_10156,N_4427,N_7001);
nor U10157 (N_10157,N_6627,N_6286);
xor U10158 (N_10158,N_6964,N_5045);
or U10159 (N_10159,N_6204,N_4028);
nor U10160 (N_10160,N_5218,N_6750);
nand U10161 (N_10161,N_4238,N_5469);
nor U10162 (N_10162,N_6248,N_7925);
and U10163 (N_10163,N_6909,N_4862);
and U10164 (N_10164,N_4949,N_5605);
nor U10165 (N_10165,N_7246,N_5611);
and U10166 (N_10166,N_4999,N_7528);
or U10167 (N_10167,N_7085,N_6902);
and U10168 (N_10168,N_5925,N_7321);
nand U10169 (N_10169,N_7305,N_4981);
and U10170 (N_10170,N_4091,N_6040);
nor U10171 (N_10171,N_7169,N_5347);
or U10172 (N_10172,N_4898,N_6742);
and U10173 (N_10173,N_7704,N_7184);
nand U10174 (N_10174,N_6646,N_4202);
or U10175 (N_10175,N_5044,N_4795);
or U10176 (N_10176,N_6430,N_4890);
nand U10177 (N_10177,N_5261,N_7686);
xnor U10178 (N_10178,N_7171,N_4667);
nor U10179 (N_10179,N_7194,N_7153);
xnor U10180 (N_10180,N_5152,N_7256);
xnor U10181 (N_10181,N_5153,N_5106);
and U10182 (N_10182,N_7036,N_6558);
nand U10183 (N_10183,N_4882,N_5763);
and U10184 (N_10184,N_5310,N_7428);
and U10185 (N_10185,N_6275,N_4380);
or U10186 (N_10186,N_4352,N_7123);
and U10187 (N_10187,N_6359,N_5901);
nor U10188 (N_10188,N_6946,N_5113);
and U10189 (N_10189,N_5191,N_7113);
or U10190 (N_10190,N_5168,N_6448);
xor U10191 (N_10191,N_4380,N_6719);
nor U10192 (N_10192,N_5061,N_5490);
xor U10193 (N_10193,N_6296,N_6758);
nor U10194 (N_10194,N_4337,N_6220);
and U10195 (N_10195,N_4491,N_6228);
or U10196 (N_10196,N_5946,N_6173);
nand U10197 (N_10197,N_6760,N_7998);
xor U10198 (N_10198,N_7429,N_5144);
or U10199 (N_10199,N_6004,N_6745);
or U10200 (N_10200,N_4911,N_4720);
nand U10201 (N_10201,N_5230,N_5299);
nor U10202 (N_10202,N_6594,N_7929);
and U10203 (N_10203,N_6375,N_6119);
nand U10204 (N_10204,N_7579,N_4020);
nor U10205 (N_10205,N_4616,N_5953);
xnor U10206 (N_10206,N_4782,N_5524);
nand U10207 (N_10207,N_4351,N_7789);
and U10208 (N_10208,N_7281,N_6987);
nand U10209 (N_10209,N_4634,N_7614);
or U10210 (N_10210,N_4621,N_5055);
and U10211 (N_10211,N_4872,N_6805);
xor U10212 (N_10212,N_6215,N_7856);
nor U10213 (N_10213,N_5378,N_4668);
nand U10214 (N_10214,N_7211,N_4970);
and U10215 (N_10215,N_6461,N_6261);
nor U10216 (N_10216,N_4614,N_4511);
xor U10217 (N_10217,N_7885,N_6968);
nand U10218 (N_10218,N_7916,N_5665);
xor U10219 (N_10219,N_7179,N_4674);
xnor U10220 (N_10220,N_7667,N_5123);
nand U10221 (N_10221,N_7673,N_6539);
nor U10222 (N_10222,N_4513,N_4885);
nand U10223 (N_10223,N_4750,N_4164);
xor U10224 (N_10224,N_7560,N_6217);
nand U10225 (N_10225,N_6536,N_7641);
nand U10226 (N_10226,N_5392,N_4107);
or U10227 (N_10227,N_4768,N_6636);
or U10228 (N_10228,N_6112,N_7576);
and U10229 (N_10229,N_4945,N_5356);
or U10230 (N_10230,N_5771,N_5876);
or U10231 (N_10231,N_4908,N_5917);
and U10232 (N_10232,N_6680,N_7143);
nor U10233 (N_10233,N_7011,N_7443);
and U10234 (N_10234,N_4173,N_6037);
and U10235 (N_10235,N_7057,N_5775);
and U10236 (N_10236,N_5343,N_7638);
nor U10237 (N_10237,N_6464,N_7292);
nor U10238 (N_10238,N_4013,N_7754);
and U10239 (N_10239,N_7550,N_5635);
nor U10240 (N_10240,N_7459,N_7709);
nor U10241 (N_10241,N_6083,N_6205);
or U10242 (N_10242,N_5026,N_6545);
nor U10243 (N_10243,N_7182,N_7491);
nand U10244 (N_10244,N_5330,N_6560);
xnor U10245 (N_10245,N_6553,N_4174);
nand U10246 (N_10246,N_6151,N_6330);
nand U10247 (N_10247,N_4708,N_4438);
or U10248 (N_10248,N_4570,N_5337);
nor U10249 (N_10249,N_7132,N_6028);
or U10250 (N_10250,N_6635,N_4181);
and U10251 (N_10251,N_6015,N_6028);
or U10252 (N_10252,N_5305,N_7980);
or U10253 (N_10253,N_5662,N_4291);
and U10254 (N_10254,N_6496,N_5731);
and U10255 (N_10255,N_7063,N_7556);
nand U10256 (N_10256,N_4560,N_7786);
or U10257 (N_10257,N_7067,N_7509);
xor U10258 (N_10258,N_7649,N_4567);
xor U10259 (N_10259,N_7950,N_7373);
nand U10260 (N_10260,N_5847,N_5964);
or U10261 (N_10261,N_4446,N_5649);
xnor U10262 (N_10262,N_5470,N_5241);
or U10263 (N_10263,N_6411,N_7421);
or U10264 (N_10264,N_6470,N_4436);
nand U10265 (N_10265,N_6826,N_7666);
xnor U10266 (N_10266,N_6611,N_7332);
xor U10267 (N_10267,N_5682,N_6115);
xnor U10268 (N_10268,N_5548,N_5479);
xor U10269 (N_10269,N_6426,N_6654);
xor U10270 (N_10270,N_5736,N_6745);
nand U10271 (N_10271,N_4924,N_5136);
nor U10272 (N_10272,N_4618,N_4171);
nor U10273 (N_10273,N_6399,N_6950);
nand U10274 (N_10274,N_6306,N_4822);
xor U10275 (N_10275,N_6435,N_6858);
and U10276 (N_10276,N_6837,N_5562);
nand U10277 (N_10277,N_4802,N_4235);
nor U10278 (N_10278,N_5871,N_7026);
xnor U10279 (N_10279,N_7815,N_7128);
or U10280 (N_10280,N_4939,N_6654);
and U10281 (N_10281,N_6454,N_4816);
or U10282 (N_10282,N_7008,N_5864);
nor U10283 (N_10283,N_4547,N_5267);
nor U10284 (N_10284,N_7895,N_7763);
and U10285 (N_10285,N_7363,N_4195);
xor U10286 (N_10286,N_5866,N_5200);
and U10287 (N_10287,N_4542,N_6653);
xor U10288 (N_10288,N_4134,N_6952);
xor U10289 (N_10289,N_5995,N_5310);
nor U10290 (N_10290,N_7868,N_4016);
xor U10291 (N_10291,N_5281,N_6571);
and U10292 (N_10292,N_5302,N_7222);
xnor U10293 (N_10293,N_7061,N_5532);
nand U10294 (N_10294,N_6836,N_4363);
nor U10295 (N_10295,N_7990,N_5055);
nor U10296 (N_10296,N_5872,N_5726);
nand U10297 (N_10297,N_7698,N_5526);
nor U10298 (N_10298,N_7960,N_7581);
nor U10299 (N_10299,N_4254,N_4931);
xnor U10300 (N_10300,N_5631,N_6913);
xor U10301 (N_10301,N_7822,N_7850);
nor U10302 (N_10302,N_5703,N_7337);
nand U10303 (N_10303,N_5771,N_7208);
xnor U10304 (N_10304,N_6170,N_6307);
or U10305 (N_10305,N_5594,N_7283);
nor U10306 (N_10306,N_4959,N_5774);
xnor U10307 (N_10307,N_6962,N_5144);
or U10308 (N_10308,N_7020,N_5349);
nand U10309 (N_10309,N_7817,N_6404);
nor U10310 (N_10310,N_6891,N_5024);
nor U10311 (N_10311,N_4517,N_6315);
nor U10312 (N_10312,N_5600,N_4296);
nor U10313 (N_10313,N_5827,N_7156);
xor U10314 (N_10314,N_7052,N_5958);
xor U10315 (N_10315,N_7733,N_7565);
nor U10316 (N_10316,N_7550,N_6258);
or U10317 (N_10317,N_5052,N_4242);
nor U10318 (N_10318,N_6954,N_6726);
and U10319 (N_10319,N_6607,N_6201);
xnor U10320 (N_10320,N_6013,N_7726);
nand U10321 (N_10321,N_5346,N_6273);
nor U10322 (N_10322,N_4182,N_5286);
nor U10323 (N_10323,N_7899,N_4584);
or U10324 (N_10324,N_5489,N_5455);
nor U10325 (N_10325,N_7139,N_4311);
nand U10326 (N_10326,N_4994,N_6021);
or U10327 (N_10327,N_6105,N_7041);
xor U10328 (N_10328,N_5485,N_5659);
nand U10329 (N_10329,N_6507,N_7760);
nor U10330 (N_10330,N_4569,N_7500);
nor U10331 (N_10331,N_7398,N_7002);
nor U10332 (N_10332,N_6276,N_7736);
or U10333 (N_10333,N_6231,N_5048);
and U10334 (N_10334,N_4133,N_7150);
or U10335 (N_10335,N_5795,N_6487);
xor U10336 (N_10336,N_4178,N_5924);
and U10337 (N_10337,N_6388,N_6198);
and U10338 (N_10338,N_4217,N_7942);
and U10339 (N_10339,N_4151,N_6302);
or U10340 (N_10340,N_5920,N_5405);
xor U10341 (N_10341,N_6041,N_6087);
xnor U10342 (N_10342,N_5530,N_6888);
and U10343 (N_10343,N_5044,N_6488);
and U10344 (N_10344,N_6033,N_7852);
nor U10345 (N_10345,N_4516,N_4609);
nor U10346 (N_10346,N_5364,N_5075);
xnor U10347 (N_10347,N_5244,N_5596);
xnor U10348 (N_10348,N_5245,N_4393);
or U10349 (N_10349,N_4124,N_7218);
nor U10350 (N_10350,N_6586,N_4743);
and U10351 (N_10351,N_5621,N_6236);
and U10352 (N_10352,N_7810,N_5719);
xnor U10353 (N_10353,N_5842,N_5412);
xor U10354 (N_10354,N_4123,N_5489);
nand U10355 (N_10355,N_6601,N_4171);
and U10356 (N_10356,N_4779,N_5189);
nand U10357 (N_10357,N_6264,N_5904);
and U10358 (N_10358,N_6185,N_4383);
xor U10359 (N_10359,N_5169,N_7146);
nand U10360 (N_10360,N_6079,N_5772);
and U10361 (N_10361,N_6725,N_6237);
nand U10362 (N_10362,N_4809,N_5631);
xor U10363 (N_10363,N_6490,N_4299);
xor U10364 (N_10364,N_7306,N_7179);
xor U10365 (N_10365,N_7926,N_7287);
and U10366 (N_10366,N_4067,N_7846);
or U10367 (N_10367,N_5831,N_4046);
nor U10368 (N_10368,N_6598,N_5280);
xor U10369 (N_10369,N_5965,N_6240);
xnor U10370 (N_10370,N_7689,N_5320);
and U10371 (N_10371,N_4027,N_5244);
or U10372 (N_10372,N_7530,N_5790);
nor U10373 (N_10373,N_7579,N_6068);
and U10374 (N_10374,N_6975,N_5971);
and U10375 (N_10375,N_5320,N_4812);
nand U10376 (N_10376,N_6752,N_5427);
xor U10377 (N_10377,N_7785,N_4112);
xor U10378 (N_10378,N_7706,N_6162);
nand U10379 (N_10379,N_6244,N_4931);
or U10380 (N_10380,N_7660,N_7997);
nand U10381 (N_10381,N_5185,N_6928);
xnor U10382 (N_10382,N_5646,N_4039);
and U10383 (N_10383,N_4461,N_6514);
or U10384 (N_10384,N_7563,N_7122);
or U10385 (N_10385,N_6946,N_6777);
xor U10386 (N_10386,N_6565,N_5160);
nand U10387 (N_10387,N_4854,N_4787);
or U10388 (N_10388,N_7853,N_4392);
nand U10389 (N_10389,N_7775,N_6868);
xnor U10390 (N_10390,N_5651,N_6668);
and U10391 (N_10391,N_7847,N_5303);
and U10392 (N_10392,N_7288,N_4491);
and U10393 (N_10393,N_5305,N_5652);
xor U10394 (N_10394,N_7514,N_7128);
xnor U10395 (N_10395,N_5539,N_7116);
or U10396 (N_10396,N_6667,N_5818);
or U10397 (N_10397,N_4762,N_7280);
nor U10398 (N_10398,N_7126,N_4434);
nor U10399 (N_10399,N_4650,N_7582);
or U10400 (N_10400,N_7324,N_6651);
or U10401 (N_10401,N_4822,N_6856);
nor U10402 (N_10402,N_5166,N_5379);
xnor U10403 (N_10403,N_7538,N_6705);
nand U10404 (N_10404,N_4953,N_5372);
nor U10405 (N_10405,N_5358,N_5549);
xor U10406 (N_10406,N_7251,N_5076);
xor U10407 (N_10407,N_6856,N_7207);
nor U10408 (N_10408,N_5806,N_5740);
or U10409 (N_10409,N_4423,N_5860);
nor U10410 (N_10410,N_4537,N_7950);
or U10411 (N_10411,N_4924,N_6992);
or U10412 (N_10412,N_4830,N_5605);
and U10413 (N_10413,N_4697,N_5089);
nand U10414 (N_10414,N_6750,N_4454);
or U10415 (N_10415,N_6213,N_6247);
nand U10416 (N_10416,N_4134,N_4570);
nand U10417 (N_10417,N_5471,N_7325);
nand U10418 (N_10418,N_7899,N_4531);
or U10419 (N_10419,N_6552,N_4600);
xnor U10420 (N_10420,N_5327,N_4087);
xnor U10421 (N_10421,N_6429,N_7058);
and U10422 (N_10422,N_4584,N_5402);
nor U10423 (N_10423,N_4396,N_4935);
nor U10424 (N_10424,N_6801,N_7308);
nand U10425 (N_10425,N_7266,N_5925);
and U10426 (N_10426,N_5709,N_7220);
xor U10427 (N_10427,N_4953,N_5680);
nor U10428 (N_10428,N_4846,N_4202);
nand U10429 (N_10429,N_4253,N_5218);
or U10430 (N_10430,N_7047,N_5063);
and U10431 (N_10431,N_5679,N_6843);
and U10432 (N_10432,N_5633,N_5557);
or U10433 (N_10433,N_4467,N_6212);
nor U10434 (N_10434,N_6591,N_4315);
and U10435 (N_10435,N_6972,N_7591);
and U10436 (N_10436,N_7475,N_7807);
xor U10437 (N_10437,N_7999,N_7368);
or U10438 (N_10438,N_4048,N_6653);
and U10439 (N_10439,N_5170,N_6500);
nor U10440 (N_10440,N_4236,N_7459);
xnor U10441 (N_10441,N_7684,N_5948);
nor U10442 (N_10442,N_5811,N_6091);
xor U10443 (N_10443,N_4938,N_6087);
xnor U10444 (N_10444,N_4297,N_4151);
xor U10445 (N_10445,N_7286,N_4125);
nor U10446 (N_10446,N_4182,N_4615);
or U10447 (N_10447,N_4330,N_5830);
and U10448 (N_10448,N_6415,N_4587);
or U10449 (N_10449,N_4722,N_4035);
nand U10450 (N_10450,N_6847,N_5357);
and U10451 (N_10451,N_6225,N_7369);
and U10452 (N_10452,N_5962,N_7600);
xor U10453 (N_10453,N_5412,N_4002);
and U10454 (N_10454,N_5142,N_4279);
or U10455 (N_10455,N_7479,N_4927);
nand U10456 (N_10456,N_7419,N_5403);
nor U10457 (N_10457,N_6863,N_7212);
nand U10458 (N_10458,N_6423,N_6146);
nor U10459 (N_10459,N_4846,N_7188);
nand U10460 (N_10460,N_6709,N_7831);
nand U10461 (N_10461,N_7301,N_5727);
nand U10462 (N_10462,N_4201,N_7999);
and U10463 (N_10463,N_7180,N_4386);
and U10464 (N_10464,N_4004,N_4013);
or U10465 (N_10465,N_6734,N_6308);
nand U10466 (N_10466,N_4780,N_5225);
nor U10467 (N_10467,N_4531,N_6905);
xnor U10468 (N_10468,N_4934,N_5407);
xnor U10469 (N_10469,N_4936,N_7675);
xnor U10470 (N_10470,N_6848,N_7553);
and U10471 (N_10471,N_4557,N_6060);
and U10472 (N_10472,N_6419,N_7015);
and U10473 (N_10473,N_6787,N_5901);
or U10474 (N_10474,N_6515,N_6118);
nor U10475 (N_10475,N_5275,N_7918);
nor U10476 (N_10476,N_5704,N_7536);
or U10477 (N_10477,N_4431,N_4000);
xor U10478 (N_10478,N_6514,N_7674);
nor U10479 (N_10479,N_5642,N_4029);
nand U10480 (N_10480,N_4878,N_6786);
and U10481 (N_10481,N_5790,N_6238);
xnor U10482 (N_10482,N_5997,N_4985);
xor U10483 (N_10483,N_4586,N_7077);
nor U10484 (N_10484,N_4771,N_4005);
nor U10485 (N_10485,N_6269,N_5070);
and U10486 (N_10486,N_5444,N_6242);
nand U10487 (N_10487,N_5056,N_6479);
and U10488 (N_10488,N_4446,N_5331);
xnor U10489 (N_10489,N_7453,N_7368);
xnor U10490 (N_10490,N_7523,N_6098);
nand U10491 (N_10491,N_7109,N_4074);
nor U10492 (N_10492,N_6347,N_7198);
or U10493 (N_10493,N_7465,N_5336);
nand U10494 (N_10494,N_6800,N_4327);
xor U10495 (N_10495,N_7793,N_7951);
and U10496 (N_10496,N_4119,N_5818);
nand U10497 (N_10497,N_6135,N_5583);
nor U10498 (N_10498,N_5192,N_4613);
xnor U10499 (N_10499,N_7088,N_6385);
nand U10500 (N_10500,N_5589,N_6112);
nor U10501 (N_10501,N_4210,N_7547);
and U10502 (N_10502,N_4476,N_6403);
nor U10503 (N_10503,N_5746,N_4328);
or U10504 (N_10504,N_4502,N_5523);
nor U10505 (N_10505,N_4831,N_5118);
and U10506 (N_10506,N_6908,N_4133);
nand U10507 (N_10507,N_7693,N_5563);
xor U10508 (N_10508,N_4402,N_6312);
and U10509 (N_10509,N_7540,N_7029);
nand U10510 (N_10510,N_7479,N_7369);
and U10511 (N_10511,N_4316,N_4466);
xnor U10512 (N_10512,N_7009,N_4656);
nor U10513 (N_10513,N_4152,N_7528);
or U10514 (N_10514,N_4711,N_5621);
nand U10515 (N_10515,N_4510,N_5647);
nor U10516 (N_10516,N_5238,N_4220);
xnor U10517 (N_10517,N_5722,N_6456);
nor U10518 (N_10518,N_7805,N_5853);
and U10519 (N_10519,N_4862,N_6534);
or U10520 (N_10520,N_6441,N_6885);
and U10521 (N_10521,N_4907,N_6489);
xor U10522 (N_10522,N_4195,N_4110);
nor U10523 (N_10523,N_5010,N_6771);
nor U10524 (N_10524,N_5975,N_5349);
or U10525 (N_10525,N_6743,N_7279);
nand U10526 (N_10526,N_4452,N_4959);
nor U10527 (N_10527,N_6294,N_4408);
or U10528 (N_10528,N_7476,N_5168);
nand U10529 (N_10529,N_4443,N_7526);
xnor U10530 (N_10530,N_5027,N_7546);
or U10531 (N_10531,N_4616,N_7446);
nand U10532 (N_10532,N_7512,N_7897);
or U10533 (N_10533,N_7677,N_5247);
xor U10534 (N_10534,N_7188,N_7666);
nand U10535 (N_10535,N_5286,N_4656);
and U10536 (N_10536,N_7884,N_4714);
nor U10537 (N_10537,N_5974,N_5151);
and U10538 (N_10538,N_7910,N_5835);
xnor U10539 (N_10539,N_5211,N_7544);
and U10540 (N_10540,N_7213,N_6777);
or U10541 (N_10541,N_7837,N_7052);
and U10542 (N_10542,N_4541,N_7012);
xor U10543 (N_10543,N_7741,N_7544);
nor U10544 (N_10544,N_5874,N_5882);
nor U10545 (N_10545,N_4920,N_5845);
nand U10546 (N_10546,N_7066,N_4345);
xnor U10547 (N_10547,N_6713,N_4276);
and U10548 (N_10548,N_4399,N_4978);
xor U10549 (N_10549,N_6130,N_6710);
nand U10550 (N_10550,N_7985,N_5394);
and U10551 (N_10551,N_4392,N_5333);
nor U10552 (N_10552,N_6687,N_7062);
xor U10553 (N_10553,N_7439,N_6516);
nor U10554 (N_10554,N_6276,N_6492);
xor U10555 (N_10555,N_4412,N_5738);
nand U10556 (N_10556,N_5220,N_6041);
or U10557 (N_10557,N_4436,N_7222);
nor U10558 (N_10558,N_4167,N_6741);
or U10559 (N_10559,N_5676,N_5860);
or U10560 (N_10560,N_4989,N_4407);
nand U10561 (N_10561,N_4086,N_5379);
and U10562 (N_10562,N_6232,N_4743);
xnor U10563 (N_10563,N_6731,N_6994);
and U10564 (N_10564,N_7101,N_5777);
nand U10565 (N_10565,N_7079,N_7636);
nand U10566 (N_10566,N_6516,N_6232);
nor U10567 (N_10567,N_4388,N_5656);
or U10568 (N_10568,N_7021,N_6510);
nor U10569 (N_10569,N_4469,N_7346);
nor U10570 (N_10570,N_7457,N_7348);
nand U10571 (N_10571,N_4033,N_4579);
and U10572 (N_10572,N_4260,N_4926);
nand U10573 (N_10573,N_5938,N_4013);
or U10574 (N_10574,N_4855,N_6497);
or U10575 (N_10575,N_4171,N_4910);
and U10576 (N_10576,N_5576,N_7461);
nand U10577 (N_10577,N_6312,N_5733);
or U10578 (N_10578,N_6496,N_4801);
nand U10579 (N_10579,N_5961,N_6887);
or U10580 (N_10580,N_6409,N_5701);
nand U10581 (N_10581,N_5067,N_6109);
nand U10582 (N_10582,N_7069,N_5735);
nand U10583 (N_10583,N_6779,N_6839);
and U10584 (N_10584,N_7768,N_5918);
and U10585 (N_10585,N_4387,N_5018);
nor U10586 (N_10586,N_6872,N_5066);
xor U10587 (N_10587,N_7271,N_4669);
or U10588 (N_10588,N_4202,N_4006);
nor U10589 (N_10589,N_4945,N_4765);
or U10590 (N_10590,N_5205,N_4275);
xnor U10591 (N_10591,N_6867,N_5058);
nand U10592 (N_10592,N_4952,N_5460);
xnor U10593 (N_10593,N_7994,N_6175);
nand U10594 (N_10594,N_5410,N_7076);
and U10595 (N_10595,N_7825,N_7307);
and U10596 (N_10596,N_7041,N_5059);
nand U10597 (N_10597,N_5447,N_7520);
nand U10598 (N_10598,N_5323,N_4544);
or U10599 (N_10599,N_7040,N_6759);
nand U10600 (N_10600,N_7123,N_7194);
or U10601 (N_10601,N_7234,N_4073);
nor U10602 (N_10602,N_4899,N_6693);
or U10603 (N_10603,N_4850,N_7996);
nor U10604 (N_10604,N_4379,N_6245);
or U10605 (N_10605,N_7809,N_6051);
and U10606 (N_10606,N_7858,N_4279);
nand U10607 (N_10607,N_6818,N_7262);
and U10608 (N_10608,N_7759,N_4122);
and U10609 (N_10609,N_5706,N_5190);
xnor U10610 (N_10610,N_7105,N_7141);
nor U10611 (N_10611,N_4483,N_7222);
nor U10612 (N_10612,N_7457,N_6204);
nand U10613 (N_10613,N_6473,N_6850);
nand U10614 (N_10614,N_6551,N_6698);
or U10615 (N_10615,N_6210,N_7623);
and U10616 (N_10616,N_5808,N_4281);
or U10617 (N_10617,N_7047,N_7632);
or U10618 (N_10618,N_7847,N_5665);
nand U10619 (N_10619,N_5064,N_6616);
nand U10620 (N_10620,N_7904,N_6313);
nor U10621 (N_10621,N_7916,N_6524);
xnor U10622 (N_10622,N_5272,N_5287);
nand U10623 (N_10623,N_5763,N_5898);
nor U10624 (N_10624,N_5091,N_6009);
and U10625 (N_10625,N_5247,N_5294);
or U10626 (N_10626,N_4831,N_4451);
xnor U10627 (N_10627,N_4451,N_5951);
nor U10628 (N_10628,N_4049,N_4387);
nand U10629 (N_10629,N_4943,N_7441);
and U10630 (N_10630,N_7197,N_6391);
nand U10631 (N_10631,N_7242,N_5115);
or U10632 (N_10632,N_5608,N_5292);
nand U10633 (N_10633,N_7845,N_4479);
nand U10634 (N_10634,N_5923,N_7116);
nand U10635 (N_10635,N_5154,N_6030);
nor U10636 (N_10636,N_5618,N_6301);
nand U10637 (N_10637,N_4041,N_7052);
xor U10638 (N_10638,N_5152,N_4634);
nor U10639 (N_10639,N_6937,N_5439);
xor U10640 (N_10640,N_4584,N_4277);
nand U10641 (N_10641,N_4050,N_6440);
xnor U10642 (N_10642,N_5880,N_6112);
xor U10643 (N_10643,N_4527,N_5680);
nor U10644 (N_10644,N_4844,N_7769);
nand U10645 (N_10645,N_5899,N_7328);
xor U10646 (N_10646,N_5235,N_7245);
xor U10647 (N_10647,N_7504,N_7990);
xor U10648 (N_10648,N_6571,N_6784);
and U10649 (N_10649,N_7437,N_4689);
and U10650 (N_10650,N_4875,N_4529);
xnor U10651 (N_10651,N_5140,N_6933);
and U10652 (N_10652,N_7887,N_5528);
and U10653 (N_10653,N_7333,N_7478);
nor U10654 (N_10654,N_4251,N_6279);
nor U10655 (N_10655,N_4467,N_4155);
nand U10656 (N_10656,N_6106,N_6825);
nor U10657 (N_10657,N_6525,N_6325);
and U10658 (N_10658,N_6838,N_5277);
nor U10659 (N_10659,N_7325,N_4272);
or U10660 (N_10660,N_7487,N_4844);
xnor U10661 (N_10661,N_7156,N_6610);
and U10662 (N_10662,N_7669,N_5057);
nand U10663 (N_10663,N_6035,N_4795);
or U10664 (N_10664,N_6006,N_6263);
nor U10665 (N_10665,N_4943,N_6079);
nor U10666 (N_10666,N_4083,N_6568);
nor U10667 (N_10667,N_7032,N_6425);
and U10668 (N_10668,N_4416,N_4158);
nor U10669 (N_10669,N_7212,N_6945);
or U10670 (N_10670,N_7091,N_5490);
xor U10671 (N_10671,N_7299,N_6607);
or U10672 (N_10672,N_6251,N_6541);
nand U10673 (N_10673,N_5344,N_5802);
nand U10674 (N_10674,N_6977,N_6113);
xnor U10675 (N_10675,N_5638,N_4358);
nor U10676 (N_10676,N_5819,N_5920);
and U10677 (N_10677,N_6573,N_5631);
and U10678 (N_10678,N_7603,N_5849);
nand U10679 (N_10679,N_7958,N_6234);
or U10680 (N_10680,N_7498,N_5862);
or U10681 (N_10681,N_5898,N_5747);
or U10682 (N_10682,N_6635,N_4957);
nand U10683 (N_10683,N_6081,N_5250);
nand U10684 (N_10684,N_7930,N_6745);
nand U10685 (N_10685,N_5521,N_7804);
nand U10686 (N_10686,N_6058,N_6477);
and U10687 (N_10687,N_7588,N_6386);
nor U10688 (N_10688,N_6890,N_7145);
nor U10689 (N_10689,N_5747,N_4234);
or U10690 (N_10690,N_7270,N_7644);
or U10691 (N_10691,N_4959,N_6141);
nor U10692 (N_10692,N_5242,N_7544);
nor U10693 (N_10693,N_6745,N_5126);
and U10694 (N_10694,N_7988,N_6922);
and U10695 (N_10695,N_4499,N_5338);
nand U10696 (N_10696,N_5667,N_7961);
xnor U10697 (N_10697,N_7090,N_4215);
or U10698 (N_10698,N_4331,N_5180);
xnor U10699 (N_10699,N_5646,N_5415);
nor U10700 (N_10700,N_7884,N_6872);
nor U10701 (N_10701,N_6814,N_6205);
nand U10702 (N_10702,N_5951,N_4849);
or U10703 (N_10703,N_5931,N_5903);
and U10704 (N_10704,N_4172,N_7747);
nor U10705 (N_10705,N_5035,N_5556);
nor U10706 (N_10706,N_4667,N_7407);
nor U10707 (N_10707,N_7123,N_4418);
nor U10708 (N_10708,N_7509,N_5103);
xnor U10709 (N_10709,N_4994,N_6465);
nor U10710 (N_10710,N_5808,N_5547);
and U10711 (N_10711,N_5122,N_4248);
nand U10712 (N_10712,N_5265,N_4871);
nor U10713 (N_10713,N_4980,N_5613);
and U10714 (N_10714,N_6419,N_5852);
nor U10715 (N_10715,N_5634,N_7316);
xnor U10716 (N_10716,N_7883,N_7326);
and U10717 (N_10717,N_7522,N_7393);
or U10718 (N_10718,N_4917,N_7770);
nand U10719 (N_10719,N_6409,N_7701);
or U10720 (N_10720,N_5253,N_4960);
nand U10721 (N_10721,N_5083,N_7197);
nand U10722 (N_10722,N_5157,N_5152);
nand U10723 (N_10723,N_5219,N_6508);
and U10724 (N_10724,N_6481,N_5475);
or U10725 (N_10725,N_4332,N_5613);
or U10726 (N_10726,N_5284,N_7804);
nor U10727 (N_10727,N_4376,N_5473);
or U10728 (N_10728,N_5920,N_6236);
nor U10729 (N_10729,N_6399,N_7289);
and U10730 (N_10730,N_7269,N_6805);
and U10731 (N_10731,N_5401,N_7042);
and U10732 (N_10732,N_6745,N_5038);
and U10733 (N_10733,N_7083,N_5634);
and U10734 (N_10734,N_7438,N_7727);
and U10735 (N_10735,N_4018,N_7220);
nor U10736 (N_10736,N_5192,N_6250);
and U10737 (N_10737,N_5477,N_7955);
nand U10738 (N_10738,N_5193,N_4408);
or U10739 (N_10739,N_6514,N_7778);
xnor U10740 (N_10740,N_4001,N_5209);
or U10741 (N_10741,N_6301,N_5756);
nor U10742 (N_10742,N_5437,N_5172);
nand U10743 (N_10743,N_7318,N_6029);
nand U10744 (N_10744,N_4144,N_7330);
nand U10745 (N_10745,N_4497,N_7135);
nor U10746 (N_10746,N_5447,N_7724);
and U10747 (N_10747,N_4151,N_6261);
xnor U10748 (N_10748,N_6741,N_4399);
or U10749 (N_10749,N_7722,N_7741);
nand U10750 (N_10750,N_4616,N_6945);
nand U10751 (N_10751,N_6773,N_7278);
nand U10752 (N_10752,N_4571,N_7374);
and U10753 (N_10753,N_6430,N_6966);
nor U10754 (N_10754,N_5750,N_4125);
xnor U10755 (N_10755,N_4518,N_7602);
nand U10756 (N_10756,N_4542,N_5321);
or U10757 (N_10757,N_7819,N_5736);
nor U10758 (N_10758,N_6642,N_5624);
nor U10759 (N_10759,N_5906,N_4367);
nor U10760 (N_10760,N_5752,N_6112);
xnor U10761 (N_10761,N_6302,N_4001);
xnor U10762 (N_10762,N_5355,N_7327);
nand U10763 (N_10763,N_6565,N_4080);
xor U10764 (N_10764,N_7635,N_4191);
nand U10765 (N_10765,N_6574,N_6757);
or U10766 (N_10766,N_7839,N_6945);
xor U10767 (N_10767,N_7101,N_6587);
and U10768 (N_10768,N_6284,N_6294);
nor U10769 (N_10769,N_4493,N_7323);
xor U10770 (N_10770,N_5899,N_7738);
and U10771 (N_10771,N_6864,N_5268);
xor U10772 (N_10772,N_4555,N_7992);
and U10773 (N_10773,N_5664,N_4835);
or U10774 (N_10774,N_5901,N_4938);
nor U10775 (N_10775,N_7136,N_5929);
xor U10776 (N_10776,N_6636,N_5021);
nand U10777 (N_10777,N_4382,N_4148);
and U10778 (N_10778,N_4011,N_6605);
nand U10779 (N_10779,N_6090,N_7524);
and U10780 (N_10780,N_7050,N_7640);
nand U10781 (N_10781,N_7076,N_7310);
or U10782 (N_10782,N_6745,N_4686);
and U10783 (N_10783,N_5999,N_6344);
nor U10784 (N_10784,N_5296,N_6786);
nor U10785 (N_10785,N_5129,N_5842);
nand U10786 (N_10786,N_4283,N_6781);
xor U10787 (N_10787,N_7615,N_7969);
nor U10788 (N_10788,N_4044,N_7116);
nand U10789 (N_10789,N_7411,N_5061);
or U10790 (N_10790,N_5308,N_4863);
nand U10791 (N_10791,N_5540,N_4500);
or U10792 (N_10792,N_7217,N_6794);
and U10793 (N_10793,N_7327,N_6035);
xnor U10794 (N_10794,N_6913,N_6742);
nor U10795 (N_10795,N_6512,N_6413);
nor U10796 (N_10796,N_7874,N_7099);
nand U10797 (N_10797,N_6782,N_7469);
and U10798 (N_10798,N_6523,N_4261);
nand U10799 (N_10799,N_7865,N_4839);
or U10800 (N_10800,N_4014,N_6805);
and U10801 (N_10801,N_4171,N_6461);
nor U10802 (N_10802,N_7351,N_4220);
and U10803 (N_10803,N_4045,N_7643);
and U10804 (N_10804,N_6402,N_4480);
nand U10805 (N_10805,N_7659,N_7892);
nand U10806 (N_10806,N_4542,N_6475);
xnor U10807 (N_10807,N_4361,N_4379);
or U10808 (N_10808,N_5589,N_7183);
xor U10809 (N_10809,N_6761,N_4863);
or U10810 (N_10810,N_5214,N_4056);
or U10811 (N_10811,N_4028,N_5888);
xor U10812 (N_10812,N_6461,N_7619);
xor U10813 (N_10813,N_4048,N_4479);
and U10814 (N_10814,N_6217,N_6405);
or U10815 (N_10815,N_5625,N_6411);
and U10816 (N_10816,N_5692,N_5170);
or U10817 (N_10817,N_6862,N_7442);
nor U10818 (N_10818,N_5346,N_7072);
or U10819 (N_10819,N_7588,N_7382);
or U10820 (N_10820,N_6098,N_4505);
or U10821 (N_10821,N_6133,N_5335);
xor U10822 (N_10822,N_5890,N_6870);
and U10823 (N_10823,N_7169,N_5200);
nor U10824 (N_10824,N_6670,N_7658);
nor U10825 (N_10825,N_6737,N_6512);
nor U10826 (N_10826,N_7352,N_4001);
nor U10827 (N_10827,N_4596,N_6685);
and U10828 (N_10828,N_5334,N_5491);
nor U10829 (N_10829,N_5307,N_7315);
and U10830 (N_10830,N_4683,N_6990);
xor U10831 (N_10831,N_4987,N_4039);
nor U10832 (N_10832,N_6635,N_7175);
xor U10833 (N_10833,N_7524,N_6501);
nand U10834 (N_10834,N_5475,N_5736);
xor U10835 (N_10835,N_7102,N_4162);
or U10836 (N_10836,N_6072,N_5640);
and U10837 (N_10837,N_5665,N_4049);
nor U10838 (N_10838,N_4752,N_6747);
xor U10839 (N_10839,N_6616,N_5931);
or U10840 (N_10840,N_6631,N_6885);
and U10841 (N_10841,N_5152,N_7547);
or U10842 (N_10842,N_5040,N_7641);
and U10843 (N_10843,N_4890,N_5319);
nor U10844 (N_10844,N_5318,N_6249);
xor U10845 (N_10845,N_7824,N_4420);
or U10846 (N_10846,N_7771,N_5994);
nor U10847 (N_10847,N_5883,N_7492);
or U10848 (N_10848,N_5385,N_4742);
xor U10849 (N_10849,N_7017,N_7381);
nand U10850 (N_10850,N_6333,N_7926);
and U10851 (N_10851,N_5974,N_6899);
and U10852 (N_10852,N_5729,N_7046);
and U10853 (N_10853,N_5525,N_4678);
xor U10854 (N_10854,N_4219,N_6503);
nand U10855 (N_10855,N_4345,N_4590);
xnor U10856 (N_10856,N_6014,N_7871);
xnor U10857 (N_10857,N_7154,N_4937);
and U10858 (N_10858,N_6155,N_6267);
nor U10859 (N_10859,N_6060,N_6810);
and U10860 (N_10860,N_5451,N_5250);
nor U10861 (N_10861,N_6448,N_6990);
nand U10862 (N_10862,N_4057,N_4389);
nand U10863 (N_10863,N_7339,N_7445);
nor U10864 (N_10864,N_6816,N_4787);
nand U10865 (N_10865,N_6671,N_6714);
nand U10866 (N_10866,N_7166,N_4345);
nor U10867 (N_10867,N_7958,N_7405);
and U10868 (N_10868,N_6778,N_5031);
or U10869 (N_10869,N_4105,N_6863);
nor U10870 (N_10870,N_5277,N_7995);
nor U10871 (N_10871,N_6444,N_7938);
or U10872 (N_10872,N_4298,N_4259);
or U10873 (N_10873,N_4838,N_7843);
xnor U10874 (N_10874,N_6252,N_7580);
or U10875 (N_10875,N_4206,N_4071);
nor U10876 (N_10876,N_5756,N_7783);
xnor U10877 (N_10877,N_6162,N_4905);
xnor U10878 (N_10878,N_5121,N_7644);
nor U10879 (N_10879,N_6354,N_5496);
xor U10880 (N_10880,N_6999,N_5558);
xnor U10881 (N_10881,N_6044,N_5455);
and U10882 (N_10882,N_6833,N_6642);
nand U10883 (N_10883,N_5142,N_5961);
xnor U10884 (N_10884,N_7787,N_4241);
nor U10885 (N_10885,N_4551,N_7379);
nand U10886 (N_10886,N_6255,N_7510);
and U10887 (N_10887,N_4909,N_7267);
or U10888 (N_10888,N_5251,N_5982);
nand U10889 (N_10889,N_5051,N_6985);
or U10890 (N_10890,N_4547,N_5923);
nor U10891 (N_10891,N_4649,N_5333);
nor U10892 (N_10892,N_5304,N_7628);
nor U10893 (N_10893,N_4458,N_4463);
nor U10894 (N_10894,N_7804,N_6114);
nor U10895 (N_10895,N_7854,N_7517);
nor U10896 (N_10896,N_6762,N_6673);
nand U10897 (N_10897,N_4096,N_7376);
and U10898 (N_10898,N_5571,N_7461);
and U10899 (N_10899,N_7122,N_4752);
nor U10900 (N_10900,N_5563,N_5315);
or U10901 (N_10901,N_4864,N_4589);
nand U10902 (N_10902,N_4188,N_4315);
or U10903 (N_10903,N_4544,N_5438);
nor U10904 (N_10904,N_4597,N_6324);
nor U10905 (N_10905,N_7506,N_4087);
or U10906 (N_10906,N_4867,N_7240);
and U10907 (N_10907,N_6017,N_6074);
and U10908 (N_10908,N_4747,N_5035);
and U10909 (N_10909,N_4259,N_6866);
xor U10910 (N_10910,N_4330,N_7784);
nand U10911 (N_10911,N_7727,N_4996);
and U10912 (N_10912,N_5688,N_6537);
and U10913 (N_10913,N_7225,N_5017);
and U10914 (N_10914,N_5143,N_7074);
xor U10915 (N_10915,N_7231,N_7776);
nand U10916 (N_10916,N_7507,N_5179);
and U10917 (N_10917,N_7932,N_6027);
xnor U10918 (N_10918,N_5074,N_5883);
and U10919 (N_10919,N_6758,N_5964);
xnor U10920 (N_10920,N_4167,N_7629);
and U10921 (N_10921,N_6490,N_6415);
or U10922 (N_10922,N_5475,N_4239);
or U10923 (N_10923,N_7271,N_7694);
nor U10924 (N_10924,N_4840,N_5923);
xnor U10925 (N_10925,N_7072,N_4030);
or U10926 (N_10926,N_6086,N_6430);
or U10927 (N_10927,N_5574,N_6661);
nor U10928 (N_10928,N_4264,N_4434);
xnor U10929 (N_10929,N_7005,N_7927);
nand U10930 (N_10930,N_6697,N_7908);
nand U10931 (N_10931,N_4823,N_4820);
and U10932 (N_10932,N_5648,N_4300);
xnor U10933 (N_10933,N_5114,N_5964);
xnor U10934 (N_10934,N_5009,N_6894);
or U10935 (N_10935,N_4859,N_4456);
or U10936 (N_10936,N_5877,N_4755);
or U10937 (N_10937,N_4855,N_5681);
nand U10938 (N_10938,N_6680,N_6791);
nor U10939 (N_10939,N_7893,N_5973);
nor U10940 (N_10940,N_5605,N_4260);
xor U10941 (N_10941,N_7671,N_7563);
nand U10942 (N_10942,N_6148,N_5256);
nand U10943 (N_10943,N_6789,N_4046);
or U10944 (N_10944,N_6227,N_5195);
nand U10945 (N_10945,N_5584,N_5145);
and U10946 (N_10946,N_6058,N_6524);
xor U10947 (N_10947,N_5288,N_5111);
nand U10948 (N_10948,N_5595,N_4443);
nor U10949 (N_10949,N_6445,N_4719);
and U10950 (N_10950,N_4674,N_4246);
xor U10951 (N_10951,N_6187,N_7845);
nor U10952 (N_10952,N_6378,N_4194);
and U10953 (N_10953,N_7208,N_4551);
nor U10954 (N_10954,N_4907,N_6899);
nand U10955 (N_10955,N_6648,N_6436);
and U10956 (N_10956,N_5018,N_7358);
and U10957 (N_10957,N_4099,N_7029);
nand U10958 (N_10958,N_4289,N_6399);
and U10959 (N_10959,N_7323,N_4613);
and U10960 (N_10960,N_5487,N_7658);
and U10961 (N_10961,N_6128,N_6827);
or U10962 (N_10962,N_7896,N_5763);
and U10963 (N_10963,N_7352,N_5880);
or U10964 (N_10964,N_7183,N_4485);
or U10965 (N_10965,N_7199,N_7012);
and U10966 (N_10966,N_6368,N_4758);
nor U10967 (N_10967,N_4997,N_6427);
nor U10968 (N_10968,N_7030,N_7470);
xnor U10969 (N_10969,N_4527,N_5987);
and U10970 (N_10970,N_5732,N_4858);
nor U10971 (N_10971,N_7362,N_6594);
and U10972 (N_10972,N_4928,N_7910);
and U10973 (N_10973,N_5250,N_4750);
xnor U10974 (N_10974,N_6371,N_4930);
xor U10975 (N_10975,N_6411,N_6084);
nand U10976 (N_10976,N_4926,N_4865);
or U10977 (N_10977,N_4710,N_7000);
nand U10978 (N_10978,N_5227,N_4454);
nor U10979 (N_10979,N_4270,N_6940);
nor U10980 (N_10980,N_7817,N_7892);
nor U10981 (N_10981,N_5703,N_5824);
xnor U10982 (N_10982,N_7721,N_5070);
nor U10983 (N_10983,N_4100,N_4385);
xnor U10984 (N_10984,N_5490,N_7286);
and U10985 (N_10985,N_5201,N_6287);
or U10986 (N_10986,N_5872,N_7509);
and U10987 (N_10987,N_4568,N_6097);
nor U10988 (N_10988,N_7268,N_6660);
nor U10989 (N_10989,N_5635,N_7513);
or U10990 (N_10990,N_4286,N_4208);
xor U10991 (N_10991,N_4547,N_7729);
nand U10992 (N_10992,N_5591,N_5157);
or U10993 (N_10993,N_4940,N_6041);
nor U10994 (N_10994,N_6421,N_5073);
xnor U10995 (N_10995,N_5794,N_4475);
or U10996 (N_10996,N_4091,N_4725);
nand U10997 (N_10997,N_7214,N_5673);
xor U10998 (N_10998,N_4781,N_7659);
nor U10999 (N_10999,N_4639,N_4267);
xnor U11000 (N_11000,N_4840,N_4751);
and U11001 (N_11001,N_6887,N_7240);
nor U11002 (N_11002,N_4644,N_5746);
nor U11003 (N_11003,N_4115,N_5080);
or U11004 (N_11004,N_6972,N_7021);
xnor U11005 (N_11005,N_7309,N_5088);
nand U11006 (N_11006,N_4062,N_6452);
xnor U11007 (N_11007,N_7681,N_7948);
or U11008 (N_11008,N_5347,N_5864);
or U11009 (N_11009,N_7986,N_6373);
xnor U11010 (N_11010,N_5299,N_4765);
and U11011 (N_11011,N_7202,N_5149);
nor U11012 (N_11012,N_6212,N_5104);
or U11013 (N_11013,N_4911,N_4199);
and U11014 (N_11014,N_7237,N_5552);
and U11015 (N_11015,N_5267,N_5469);
xor U11016 (N_11016,N_4777,N_5079);
and U11017 (N_11017,N_7214,N_7678);
nor U11018 (N_11018,N_5287,N_6878);
or U11019 (N_11019,N_5817,N_6293);
nor U11020 (N_11020,N_6034,N_7333);
and U11021 (N_11021,N_5545,N_6711);
nor U11022 (N_11022,N_4818,N_6001);
nor U11023 (N_11023,N_5262,N_6605);
nor U11024 (N_11024,N_4131,N_7317);
nand U11025 (N_11025,N_7756,N_4971);
xnor U11026 (N_11026,N_7649,N_7987);
nor U11027 (N_11027,N_5160,N_6902);
or U11028 (N_11028,N_4423,N_5521);
nand U11029 (N_11029,N_7656,N_6032);
or U11030 (N_11030,N_5237,N_7883);
nor U11031 (N_11031,N_7087,N_5953);
xnor U11032 (N_11032,N_6940,N_5880);
or U11033 (N_11033,N_4845,N_7886);
and U11034 (N_11034,N_5825,N_6032);
and U11035 (N_11035,N_5625,N_5635);
nand U11036 (N_11036,N_4354,N_6843);
and U11037 (N_11037,N_6205,N_7020);
nor U11038 (N_11038,N_5613,N_5164);
nor U11039 (N_11039,N_6094,N_5831);
nor U11040 (N_11040,N_6351,N_7646);
or U11041 (N_11041,N_4289,N_4464);
nor U11042 (N_11042,N_5390,N_6050);
xor U11043 (N_11043,N_6768,N_6811);
nor U11044 (N_11044,N_5406,N_4564);
nand U11045 (N_11045,N_4882,N_5928);
xnor U11046 (N_11046,N_6892,N_4683);
and U11047 (N_11047,N_6357,N_7554);
nor U11048 (N_11048,N_7181,N_7035);
and U11049 (N_11049,N_5957,N_7654);
and U11050 (N_11050,N_5222,N_4386);
xor U11051 (N_11051,N_6902,N_5355);
or U11052 (N_11052,N_7282,N_5444);
xor U11053 (N_11053,N_4442,N_5494);
nand U11054 (N_11054,N_5002,N_4753);
nand U11055 (N_11055,N_4731,N_7438);
nand U11056 (N_11056,N_6679,N_6793);
nand U11057 (N_11057,N_5980,N_4068);
xor U11058 (N_11058,N_6781,N_7920);
or U11059 (N_11059,N_4183,N_6649);
xor U11060 (N_11060,N_6616,N_5250);
nand U11061 (N_11061,N_4883,N_6307);
or U11062 (N_11062,N_6783,N_6632);
or U11063 (N_11063,N_4562,N_4226);
and U11064 (N_11064,N_4855,N_5084);
xnor U11065 (N_11065,N_7241,N_7264);
and U11066 (N_11066,N_7692,N_6894);
or U11067 (N_11067,N_4182,N_7892);
nand U11068 (N_11068,N_4360,N_5742);
xnor U11069 (N_11069,N_4156,N_4310);
nand U11070 (N_11070,N_4898,N_6651);
and U11071 (N_11071,N_6304,N_7729);
xor U11072 (N_11072,N_6895,N_4851);
nand U11073 (N_11073,N_4538,N_7697);
or U11074 (N_11074,N_7152,N_4180);
or U11075 (N_11075,N_4488,N_6217);
and U11076 (N_11076,N_5701,N_4759);
or U11077 (N_11077,N_4060,N_6565);
or U11078 (N_11078,N_6075,N_5829);
or U11079 (N_11079,N_6164,N_6449);
nand U11080 (N_11080,N_5454,N_4616);
or U11081 (N_11081,N_7616,N_7587);
nor U11082 (N_11082,N_4720,N_5721);
xnor U11083 (N_11083,N_7465,N_6898);
and U11084 (N_11084,N_7445,N_4837);
nand U11085 (N_11085,N_4205,N_5808);
xor U11086 (N_11086,N_5763,N_5076);
nor U11087 (N_11087,N_5516,N_6769);
and U11088 (N_11088,N_4909,N_6052);
or U11089 (N_11089,N_6150,N_7784);
and U11090 (N_11090,N_4383,N_7771);
and U11091 (N_11091,N_6568,N_7207);
nand U11092 (N_11092,N_6327,N_4202);
or U11093 (N_11093,N_4780,N_5964);
nand U11094 (N_11094,N_4097,N_5214);
nand U11095 (N_11095,N_5661,N_4297);
or U11096 (N_11096,N_6478,N_5884);
nand U11097 (N_11097,N_4346,N_7374);
or U11098 (N_11098,N_4425,N_6739);
nand U11099 (N_11099,N_6066,N_6060);
nand U11100 (N_11100,N_5369,N_6744);
xor U11101 (N_11101,N_6823,N_5772);
and U11102 (N_11102,N_7483,N_7679);
and U11103 (N_11103,N_7336,N_7033);
nor U11104 (N_11104,N_5597,N_4555);
or U11105 (N_11105,N_7187,N_6002);
xor U11106 (N_11106,N_6351,N_7660);
nor U11107 (N_11107,N_7959,N_4038);
and U11108 (N_11108,N_6690,N_5572);
or U11109 (N_11109,N_5007,N_7307);
or U11110 (N_11110,N_6155,N_7788);
and U11111 (N_11111,N_7025,N_6795);
and U11112 (N_11112,N_6978,N_7924);
nor U11113 (N_11113,N_5038,N_6798);
xnor U11114 (N_11114,N_4902,N_5060);
or U11115 (N_11115,N_5580,N_5252);
nor U11116 (N_11116,N_4057,N_4072);
xor U11117 (N_11117,N_7007,N_6857);
or U11118 (N_11118,N_6545,N_4590);
and U11119 (N_11119,N_5710,N_6599);
or U11120 (N_11120,N_4733,N_4086);
or U11121 (N_11121,N_7931,N_4646);
or U11122 (N_11122,N_4034,N_5083);
nand U11123 (N_11123,N_4280,N_4925);
xor U11124 (N_11124,N_6949,N_5235);
and U11125 (N_11125,N_5078,N_6936);
and U11126 (N_11126,N_4662,N_6837);
or U11127 (N_11127,N_5207,N_7124);
nand U11128 (N_11128,N_7431,N_7052);
or U11129 (N_11129,N_7063,N_6250);
nor U11130 (N_11130,N_7011,N_4455);
nor U11131 (N_11131,N_7065,N_7016);
nand U11132 (N_11132,N_4141,N_6530);
or U11133 (N_11133,N_7445,N_5088);
nand U11134 (N_11134,N_6695,N_6302);
xnor U11135 (N_11135,N_5568,N_5239);
and U11136 (N_11136,N_5743,N_5326);
xnor U11137 (N_11137,N_5648,N_4174);
nand U11138 (N_11138,N_4292,N_6173);
nand U11139 (N_11139,N_4915,N_5207);
and U11140 (N_11140,N_4080,N_5947);
nor U11141 (N_11141,N_4421,N_4446);
or U11142 (N_11142,N_7661,N_5490);
nor U11143 (N_11143,N_5419,N_7543);
nor U11144 (N_11144,N_7067,N_4032);
nand U11145 (N_11145,N_5633,N_6979);
nand U11146 (N_11146,N_4992,N_4741);
or U11147 (N_11147,N_6772,N_6172);
and U11148 (N_11148,N_4157,N_4280);
or U11149 (N_11149,N_4882,N_4623);
xnor U11150 (N_11150,N_6234,N_4721);
nor U11151 (N_11151,N_7851,N_5069);
nor U11152 (N_11152,N_7683,N_5176);
xnor U11153 (N_11153,N_6430,N_4170);
nor U11154 (N_11154,N_7255,N_5628);
or U11155 (N_11155,N_5832,N_4067);
xor U11156 (N_11156,N_7272,N_6077);
nor U11157 (N_11157,N_4741,N_5514);
xnor U11158 (N_11158,N_5691,N_7265);
xor U11159 (N_11159,N_6072,N_6567);
nand U11160 (N_11160,N_7743,N_4919);
or U11161 (N_11161,N_5418,N_5641);
and U11162 (N_11162,N_5296,N_7842);
xor U11163 (N_11163,N_4426,N_4825);
xnor U11164 (N_11164,N_6165,N_5900);
and U11165 (N_11165,N_6882,N_7415);
and U11166 (N_11166,N_5009,N_7376);
or U11167 (N_11167,N_6732,N_6596);
and U11168 (N_11168,N_4321,N_7006);
and U11169 (N_11169,N_7915,N_4411);
and U11170 (N_11170,N_7683,N_4885);
xor U11171 (N_11171,N_7880,N_4628);
xor U11172 (N_11172,N_6865,N_4293);
or U11173 (N_11173,N_5856,N_5129);
or U11174 (N_11174,N_5718,N_6623);
nor U11175 (N_11175,N_7779,N_5885);
xor U11176 (N_11176,N_5714,N_5136);
nor U11177 (N_11177,N_4134,N_6321);
xnor U11178 (N_11178,N_7992,N_5180);
nor U11179 (N_11179,N_5443,N_5845);
xor U11180 (N_11180,N_5881,N_4914);
or U11181 (N_11181,N_4759,N_4583);
nand U11182 (N_11182,N_5255,N_7879);
nand U11183 (N_11183,N_4608,N_6218);
xnor U11184 (N_11184,N_4361,N_4171);
and U11185 (N_11185,N_7826,N_6287);
nand U11186 (N_11186,N_5175,N_5548);
or U11187 (N_11187,N_7363,N_6958);
nor U11188 (N_11188,N_7454,N_4077);
xnor U11189 (N_11189,N_6741,N_6283);
nor U11190 (N_11190,N_6318,N_5618);
nor U11191 (N_11191,N_6487,N_4376);
nand U11192 (N_11192,N_7848,N_7046);
xnor U11193 (N_11193,N_5794,N_4133);
and U11194 (N_11194,N_4229,N_6567);
and U11195 (N_11195,N_4499,N_4245);
or U11196 (N_11196,N_6957,N_5024);
and U11197 (N_11197,N_6114,N_4648);
or U11198 (N_11198,N_4822,N_7265);
nand U11199 (N_11199,N_7388,N_5410);
xnor U11200 (N_11200,N_4526,N_6042);
xor U11201 (N_11201,N_4590,N_5676);
or U11202 (N_11202,N_4501,N_5664);
xnor U11203 (N_11203,N_6564,N_6833);
or U11204 (N_11204,N_5796,N_4759);
xor U11205 (N_11205,N_5556,N_6309);
xnor U11206 (N_11206,N_4743,N_6311);
nand U11207 (N_11207,N_6005,N_6600);
or U11208 (N_11208,N_6279,N_5675);
nand U11209 (N_11209,N_5026,N_4670);
nand U11210 (N_11210,N_4202,N_5431);
xnor U11211 (N_11211,N_7523,N_6480);
or U11212 (N_11212,N_4915,N_5206);
nor U11213 (N_11213,N_6318,N_5244);
or U11214 (N_11214,N_7593,N_7598);
nand U11215 (N_11215,N_5634,N_7875);
nor U11216 (N_11216,N_7322,N_5461);
and U11217 (N_11217,N_4970,N_7439);
and U11218 (N_11218,N_7188,N_4012);
and U11219 (N_11219,N_6012,N_6077);
xnor U11220 (N_11220,N_6363,N_5644);
xor U11221 (N_11221,N_4563,N_7835);
and U11222 (N_11222,N_4759,N_7381);
nor U11223 (N_11223,N_7166,N_7956);
nor U11224 (N_11224,N_6297,N_5307);
or U11225 (N_11225,N_4043,N_5229);
nor U11226 (N_11226,N_7916,N_5353);
xor U11227 (N_11227,N_7106,N_7803);
nor U11228 (N_11228,N_6292,N_7935);
nand U11229 (N_11229,N_4312,N_4601);
nand U11230 (N_11230,N_5192,N_5388);
nand U11231 (N_11231,N_7860,N_7910);
and U11232 (N_11232,N_5301,N_4986);
xnor U11233 (N_11233,N_4344,N_4249);
nand U11234 (N_11234,N_5163,N_4998);
and U11235 (N_11235,N_4901,N_5702);
xor U11236 (N_11236,N_4177,N_6640);
nand U11237 (N_11237,N_5080,N_5289);
nand U11238 (N_11238,N_5573,N_5303);
xor U11239 (N_11239,N_7244,N_5791);
xnor U11240 (N_11240,N_5823,N_5783);
nand U11241 (N_11241,N_4264,N_5263);
xnor U11242 (N_11242,N_4812,N_7307);
xnor U11243 (N_11243,N_6347,N_6911);
or U11244 (N_11244,N_6492,N_5953);
or U11245 (N_11245,N_7370,N_5079);
and U11246 (N_11246,N_5291,N_7171);
and U11247 (N_11247,N_5263,N_5715);
and U11248 (N_11248,N_7022,N_4848);
and U11249 (N_11249,N_4579,N_7437);
xnor U11250 (N_11250,N_7802,N_4987);
or U11251 (N_11251,N_5919,N_6148);
and U11252 (N_11252,N_6182,N_7180);
nand U11253 (N_11253,N_4897,N_6840);
nand U11254 (N_11254,N_5113,N_7656);
nor U11255 (N_11255,N_7238,N_7130);
and U11256 (N_11256,N_5683,N_4709);
and U11257 (N_11257,N_7500,N_6062);
or U11258 (N_11258,N_4800,N_4035);
nor U11259 (N_11259,N_5808,N_6222);
xnor U11260 (N_11260,N_4289,N_5007);
or U11261 (N_11261,N_6816,N_4953);
or U11262 (N_11262,N_5419,N_5049);
nand U11263 (N_11263,N_6270,N_5202);
nor U11264 (N_11264,N_7474,N_7701);
and U11265 (N_11265,N_7968,N_7794);
nor U11266 (N_11266,N_6607,N_6767);
or U11267 (N_11267,N_6588,N_6681);
nand U11268 (N_11268,N_4516,N_6245);
or U11269 (N_11269,N_7902,N_5298);
and U11270 (N_11270,N_5492,N_5059);
nor U11271 (N_11271,N_4451,N_7119);
and U11272 (N_11272,N_4871,N_7210);
nand U11273 (N_11273,N_7120,N_7813);
and U11274 (N_11274,N_6096,N_7637);
xor U11275 (N_11275,N_6847,N_4069);
or U11276 (N_11276,N_6767,N_7151);
nand U11277 (N_11277,N_7467,N_6653);
nor U11278 (N_11278,N_5148,N_7292);
xor U11279 (N_11279,N_4665,N_5406);
nor U11280 (N_11280,N_6330,N_4823);
nand U11281 (N_11281,N_5672,N_5857);
and U11282 (N_11282,N_6547,N_4045);
nor U11283 (N_11283,N_4091,N_7680);
or U11284 (N_11284,N_6679,N_7902);
nor U11285 (N_11285,N_6420,N_7592);
and U11286 (N_11286,N_4759,N_7122);
or U11287 (N_11287,N_4699,N_7061);
xnor U11288 (N_11288,N_5479,N_7570);
nor U11289 (N_11289,N_5662,N_7232);
or U11290 (N_11290,N_4431,N_5271);
nand U11291 (N_11291,N_6367,N_6812);
nor U11292 (N_11292,N_5579,N_5974);
nand U11293 (N_11293,N_7584,N_4604);
or U11294 (N_11294,N_7349,N_7080);
or U11295 (N_11295,N_6482,N_4821);
xor U11296 (N_11296,N_4558,N_5427);
xnor U11297 (N_11297,N_5613,N_4091);
or U11298 (N_11298,N_6899,N_6481);
nor U11299 (N_11299,N_6633,N_6610);
nand U11300 (N_11300,N_6346,N_4348);
xor U11301 (N_11301,N_5052,N_6822);
and U11302 (N_11302,N_7054,N_6906);
nand U11303 (N_11303,N_5979,N_7091);
nand U11304 (N_11304,N_5091,N_4845);
and U11305 (N_11305,N_5456,N_7138);
nand U11306 (N_11306,N_5585,N_6305);
nand U11307 (N_11307,N_7178,N_4317);
nor U11308 (N_11308,N_6340,N_4171);
nand U11309 (N_11309,N_7177,N_6425);
xor U11310 (N_11310,N_5746,N_7621);
nand U11311 (N_11311,N_5479,N_5986);
nand U11312 (N_11312,N_7457,N_4324);
and U11313 (N_11313,N_7996,N_4214);
or U11314 (N_11314,N_4640,N_7734);
and U11315 (N_11315,N_5688,N_7823);
xnor U11316 (N_11316,N_5775,N_6358);
or U11317 (N_11317,N_7579,N_7048);
xnor U11318 (N_11318,N_5394,N_5456);
or U11319 (N_11319,N_5806,N_7019);
or U11320 (N_11320,N_4845,N_5167);
and U11321 (N_11321,N_5921,N_5426);
nand U11322 (N_11322,N_5649,N_6427);
and U11323 (N_11323,N_5326,N_6269);
nand U11324 (N_11324,N_7729,N_7864);
nor U11325 (N_11325,N_7676,N_5974);
xnor U11326 (N_11326,N_4190,N_6092);
and U11327 (N_11327,N_7387,N_6249);
nor U11328 (N_11328,N_6091,N_4144);
nor U11329 (N_11329,N_5559,N_6810);
nor U11330 (N_11330,N_7752,N_6760);
and U11331 (N_11331,N_7389,N_5049);
nor U11332 (N_11332,N_6169,N_7737);
nor U11333 (N_11333,N_5256,N_7082);
and U11334 (N_11334,N_4223,N_5047);
and U11335 (N_11335,N_7547,N_5381);
nand U11336 (N_11336,N_4145,N_6929);
nand U11337 (N_11337,N_5058,N_5112);
and U11338 (N_11338,N_5657,N_5386);
nand U11339 (N_11339,N_4059,N_5131);
nand U11340 (N_11340,N_6061,N_4319);
and U11341 (N_11341,N_4596,N_4602);
xor U11342 (N_11342,N_6608,N_4952);
xor U11343 (N_11343,N_4487,N_5433);
nor U11344 (N_11344,N_5424,N_5354);
nand U11345 (N_11345,N_6330,N_5281);
xnor U11346 (N_11346,N_5844,N_5122);
and U11347 (N_11347,N_5604,N_6058);
nand U11348 (N_11348,N_5719,N_7138);
nand U11349 (N_11349,N_4399,N_6152);
or U11350 (N_11350,N_6544,N_7206);
nand U11351 (N_11351,N_6872,N_4391);
nor U11352 (N_11352,N_4834,N_6961);
xor U11353 (N_11353,N_7630,N_6829);
nand U11354 (N_11354,N_6294,N_4838);
or U11355 (N_11355,N_5206,N_5504);
and U11356 (N_11356,N_7849,N_7810);
nand U11357 (N_11357,N_5833,N_5260);
xnor U11358 (N_11358,N_5221,N_5606);
xnor U11359 (N_11359,N_5461,N_5145);
and U11360 (N_11360,N_5110,N_6224);
and U11361 (N_11361,N_6960,N_4982);
nor U11362 (N_11362,N_5578,N_6378);
and U11363 (N_11363,N_6676,N_4509);
xor U11364 (N_11364,N_7960,N_7687);
or U11365 (N_11365,N_5911,N_5501);
xor U11366 (N_11366,N_6585,N_7854);
nand U11367 (N_11367,N_7291,N_7458);
and U11368 (N_11368,N_6616,N_5851);
xor U11369 (N_11369,N_4376,N_7498);
or U11370 (N_11370,N_5014,N_4926);
or U11371 (N_11371,N_4001,N_7728);
nor U11372 (N_11372,N_5336,N_4780);
and U11373 (N_11373,N_5558,N_4837);
xor U11374 (N_11374,N_5465,N_7824);
and U11375 (N_11375,N_6507,N_7924);
and U11376 (N_11376,N_6204,N_6092);
xnor U11377 (N_11377,N_4449,N_5406);
xnor U11378 (N_11378,N_5570,N_5332);
or U11379 (N_11379,N_4703,N_4241);
nand U11380 (N_11380,N_7425,N_6351);
nor U11381 (N_11381,N_5622,N_7095);
nand U11382 (N_11382,N_4887,N_5398);
or U11383 (N_11383,N_4892,N_7901);
and U11384 (N_11384,N_5996,N_7256);
nor U11385 (N_11385,N_4053,N_4381);
xor U11386 (N_11386,N_6132,N_5770);
nand U11387 (N_11387,N_6774,N_5273);
nor U11388 (N_11388,N_7466,N_5850);
nor U11389 (N_11389,N_4997,N_6714);
nor U11390 (N_11390,N_7823,N_7850);
nand U11391 (N_11391,N_7364,N_5659);
nand U11392 (N_11392,N_7568,N_6467);
xor U11393 (N_11393,N_7935,N_7307);
xor U11394 (N_11394,N_4700,N_6875);
nor U11395 (N_11395,N_4892,N_6387);
and U11396 (N_11396,N_6591,N_7941);
nand U11397 (N_11397,N_4956,N_5268);
or U11398 (N_11398,N_6191,N_7781);
nor U11399 (N_11399,N_5831,N_5993);
xor U11400 (N_11400,N_5611,N_6278);
nor U11401 (N_11401,N_5491,N_7461);
nor U11402 (N_11402,N_5028,N_6531);
nand U11403 (N_11403,N_5932,N_4051);
and U11404 (N_11404,N_7324,N_7971);
xnor U11405 (N_11405,N_4311,N_5006);
or U11406 (N_11406,N_4401,N_6141);
nor U11407 (N_11407,N_7752,N_5829);
and U11408 (N_11408,N_5408,N_4156);
xor U11409 (N_11409,N_7726,N_6757);
or U11410 (N_11410,N_5014,N_5183);
xnor U11411 (N_11411,N_7021,N_6832);
or U11412 (N_11412,N_4034,N_4298);
xnor U11413 (N_11413,N_7792,N_5344);
nor U11414 (N_11414,N_5968,N_7137);
nand U11415 (N_11415,N_6341,N_5602);
and U11416 (N_11416,N_7229,N_7744);
nand U11417 (N_11417,N_4811,N_7879);
or U11418 (N_11418,N_4071,N_4819);
or U11419 (N_11419,N_4806,N_6250);
xor U11420 (N_11420,N_7416,N_5975);
nor U11421 (N_11421,N_5278,N_4569);
xnor U11422 (N_11422,N_7347,N_6512);
or U11423 (N_11423,N_7242,N_5436);
nand U11424 (N_11424,N_4060,N_4409);
or U11425 (N_11425,N_5828,N_6966);
nor U11426 (N_11426,N_7151,N_4138);
nor U11427 (N_11427,N_5220,N_7725);
xor U11428 (N_11428,N_5433,N_6164);
nand U11429 (N_11429,N_5098,N_5303);
or U11430 (N_11430,N_5598,N_7797);
and U11431 (N_11431,N_5316,N_4826);
nor U11432 (N_11432,N_5225,N_6878);
or U11433 (N_11433,N_5437,N_4233);
or U11434 (N_11434,N_4458,N_6921);
and U11435 (N_11435,N_6882,N_6639);
nor U11436 (N_11436,N_6278,N_6070);
or U11437 (N_11437,N_7556,N_5299);
nor U11438 (N_11438,N_6679,N_4823);
nand U11439 (N_11439,N_6045,N_5300);
nand U11440 (N_11440,N_6020,N_5141);
xnor U11441 (N_11441,N_4865,N_5230);
nor U11442 (N_11442,N_6355,N_4980);
nand U11443 (N_11443,N_4219,N_6258);
xnor U11444 (N_11444,N_7766,N_6261);
nor U11445 (N_11445,N_6999,N_5490);
xor U11446 (N_11446,N_7776,N_6226);
nand U11447 (N_11447,N_4470,N_4545);
nand U11448 (N_11448,N_5132,N_6352);
xor U11449 (N_11449,N_5295,N_4971);
or U11450 (N_11450,N_7438,N_4315);
nor U11451 (N_11451,N_4227,N_5279);
or U11452 (N_11452,N_4327,N_7163);
nand U11453 (N_11453,N_7633,N_4925);
nand U11454 (N_11454,N_6329,N_5346);
and U11455 (N_11455,N_4318,N_5481);
nor U11456 (N_11456,N_7002,N_4149);
xnor U11457 (N_11457,N_4004,N_6224);
nand U11458 (N_11458,N_5556,N_6610);
and U11459 (N_11459,N_7050,N_7277);
xnor U11460 (N_11460,N_4870,N_7667);
xor U11461 (N_11461,N_7881,N_7095);
nor U11462 (N_11462,N_6808,N_5922);
and U11463 (N_11463,N_4302,N_4241);
or U11464 (N_11464,N_6429,N_4740);
nor U11465 (N_11465,N_6148,N_7844);
xnor U11466 (N_11466,N_5143,N_6463);
xnor U11467 (N_11467,N_6984,N_7524);
and U11468 (N_11468,N_5680,N_6010);
nand U11469 (N_11469,N_7030,N_4115);
or U11470 (N_11470,N_4665,N_7601);
nand U11471 (N_11471,N_5674,N_6910);
nand U11472 (N_11472,N_5541,N_5187);
xnor U11473 (N_11473,N_7545,N_6430);
nor U11474 (N_11474,N_6230,N_7106);
and U11475 (N_11475,N_5028,N_4262);
and U11476 (N_11476,N_4933,N_6020);
xor U11477 (N_11477,N_4146,N_4628);
xor U11478 (N_11478,N_4140,N_4819);
nor U11479 (N_11479,N_4673,N_7450);
or U11480 (N_11480,N_4908,N_7978);
xor U11481 (N_11481,N_7775,N_7022);
and U11482 (N_11482,N_7260,N_6542);
nand U11483 (N_11483,N_5712,N_6377);
and U11484 (N_11484,N_5194,N_6989);
nor U11485 (N_11485,N_5912,N_4656);
nand U11486 (N_11486,N_4152,N_6519);
xor U11487 (N_11487,N_4163,N_7984);
and U11488 (N_11488,N_5319,N_5300);
and U11489 (N_11489,N_6928,N_4862);
or U11490 (N_11490,N_6589,N_6926);
or U11491 (N_11491,N_4493,N_5988);
nor U11492 (N_11492,N_5242,N_7106);
nand U11493 (N_11493,N_5987,N_7768);
or U11494 (N_11494,N_4385,N_6830);
nor U11495 (N_11495,N_6948,N_4794);
nand U11496 (N_11496,N_5635,N_5813);
and U11497 (N_11497,N_6547,N_7416);
nor U11498 (N_11498,N_6342,N_7906);
xor U11499 (N_11499,N_7203,N_7995);
nand U11500 (N_11500,N_7577,N_5705);
nand U11501 (N_11501,N_4289,N_5455);
nor U11502 (N_11502,N_7528,N_5541);
nand U11503 (N_11503,N_7035,N_7247);
nand U11504 (N_11504,N_4756,N_7255);
and U11505 (N_11505,N_5983,N_4747);
nand U11506 (N_11506,N_6844,N_7387);
xor U11507 (N_11507,N_6916,N_5678);
or U11508 (N_11508,N_5725,N_6952);
and U11509 (N_11509,N_7903,N_5370);
nand U11510 (N_11510,N_5885,N_6623);
xnor U11511 (N_11511,N_5011,N_6304);
nand U11512 (N_11512,N_7285,N_5304);
nand U11513 (N_11513,N_4810,N_4794);
nand U11514 (N_11514,N_4172,N_7443);
xor U11515 (N_11515,N_5791,N_4880);
or U11516 (N_11516,N_7887,N_6057);
nor U11517 (N_11517,N_6584,N_5170);
nand U11518 (N_11518,N_5379,N_5427);
or U11519 (N_11519,N_5308,N_6316);
nor U11520 (N_11520,N_5795,N_4487);
nor U11521 (N_11521,N_4974,N_4545);
nand U11522 (N_11522,N_5604,N_6214);
nand U11523 (N_11523,N_6835,N_4105);
or U11524 (N_11524,N_7196,N_5566);
or U11525 (N_11525,N_6387,N_4652);
or U11526 (N_11526,N_5472,N_4369);
and U11527 (N_11527,N_4666,N_4941);
nor U11528 (N_11528,N_4032,N_4027);
or U11529 (N_11529,N_4098,N_7039);
or U11530 (N_11530,N_5095,N_7110);
nand U11531 (N_11531,N_6213,N_6725);
and U11532 (N_11532,N_4839,N_5540);
nand U11533 (N_11533,N_6365,N_6458);
xnor U11534 (N_11534,N_6682,N_5352);
nand U11535 (N_11535,N_5684,N_6056);
and U11536 (N_11536,N_4298,N_6003);
or U11537 (N_11537,N_7086,N_4752);
or U11538 (N_11538,N_7037,N_6773);
or U11539 (N_11539,N_7270,N_6295);
or U11540 (N_11540,N_5157,N_4631);
nor U11541 (N_11541,N_7162,N_7488);
or U11542 (N_11542,N_4459,N_7663);
xnor U11543 (N_11543,N_6054,N_7623);
nand U11544 (N_11544,N_7022,N_6838);
and U11545 (N_11545,N_4777,N_7466);
xnor U11546 (N_11546,N_7573,N_6493);
or U11547 (N_11547,N_4921,N_4385);
xor U11548 (N_11548,N_4273,N_7921);
xor U11549 (N_11549,N_6890,N_6723);
or U11550 (N_11550,N_4897,N_4889);
or U11551 (N_11551,N_4543,N_6299);
xor U11552 (N_11552,N_5242,N_6873);
and U11553 (N_11553,N_6449,N_6168);
and U11554 (N_11554,N_4023,N_4084);
xnor U11555 (N_11555,N_4025,N_6473);
and U11556 (N_11556,N_4392,N_7011);
xnor U11557 (N_11557,N_7940,N_7226);
nand U11558 (N_11558,N_4991,N_6415);
nor U11559 (N_11559,N_6590,N_5298);
xnor U11560 (N_11560,N_6452,N_4132);
and U11561 (N_11561,N_6011,N_4214);
nand U11562 (N_11562,N_4167,N_4704);
or U11563 (N_11563,N_4509,N_5667);
nand U11564 (N_11564,N_5964,N_4871);
or U11565 (N_11565,N_6549,N_6473);
xnor U11566 (N_11566,N_4441,N_5164);
xor U11567 (N_11567,N_4500,N_5092);
or U11568 (N_11568,N_4052,N_7319);
and U11569 (N_11569,N_5173,N_5578);
and U11570 (N_11570,N_4360,N_7363);
xor U11571 (N_11571,N_4058,N_7476);
xor U11572 (N_11572,N_5583,N_4556);
xnor U11573 (N_11573,N_7736,N_7713);
and U11574 (N_11574,N_4051,N_6496);
nand U11575 (N_11575,N_7269,N_6238);
and U11576 (N_11576,N_4130,N_7958);
nor U11577 (N_11577,N_5616,N_6358);
or U11578 (N_11578,N_5639,N_4430);
nand U11579 (N_11579,N_5042,N_5672);
or U11580 (N_11580,N_4052,N_6460);
xor U11581 (N_11581,N_7321,N_7941);
and U11582 (N_11582,N_6690,N_7284);
nor U11583 (N_11583,N_6402,N_5244);
xor U11584 (N_11584,N_4434,N_5479);
xor U11585 (N_11585,N_6202,N_4557);
nor U11586 (N_11586,N_5727,N_6076);
xor U11587 (N_11587,N_6374,N_6841);
nand U11588 (N_11588,N_7682,N_4888);
nand U11589 (N_11589,N_7387,N_5814);
or U11590 (N_11590,N_5378,N_6892);
nand U11591 (N_11591,N_5229,N_5326);
and U11592 (N_11592,N_4543,N_4445);
nor U11593 (N_11593,N_4654,N_6356);
nand U11594 (N_11594,N_4459,N_6054);
and U11595 (N_11595,N_7377,N_5316);
xnor U11596 (N_11596,N_4626,N_5697);
nor U11597 (N_11597,N_5067,N_5971);
and U11598 (N_11598,N_5659,N_5942);
or U11599 (N_11599,N_4538,N_6758);
nor U11600 (N_11600,N_7407,N_6753);
nor U11601 (N_11601,N_6188,N_6521);
or U11602 (N_11602,N_5748,N_7769);
nand U11603 (N_11603,N_4434,N_7322);
and U11604 (N_11604,N_5871,N_6666);
nor U11605 (N_11605,N_7471,N_7974);
and U11606 (N_11606,N_6296,N_6136);
nand U11607 (N_11607,N_5916,N_6154);
nor U11608 (N_11608,N_5141,N_6429);
or U11609 (N_11609,N_7845,N_4870);
and U11610 (N_11610,N_7339,N_5270);
nor U11611 (N_11611,N_7799,N_7904);
and U11612 (N_11612,N_6627,N_6124);
xor U11613 (N_11613,N_7585,N_4849);
nand U11614 (N_11614,N_7195,N_7438);
nand U11615 (N_11615,N_7851,N_7262);
nand U11616 (N_11616,N_6728,N_5789);
xnor U11617 (N_11617,N_6637,N_5964);
nor U11618 (N_11618,N_4309,N_5333);
xor U11619 (N_11619,N_7502,N_5336);
and U11620 (N_11620,N_5716,N_5853);
nand U11621 (N_11621,N_6306,N_5145);
nor U11622 (N_11622,N_7270,N_5006);
xor U11623 (N_11623,N_7188,N_7063);
nor U11624 (N_11624,N_6533,N_6890);
nand U11625 (N_11625,N_6730,N_4763);
or U11626 (N_11626,N_6691,N_7400);
xor U11627 (N_11627,N_6456,N_5134);
and U11628 (N_11628,N_5463,N_5383);
and U11629 (N_11629,N_5306,N_6821);
nor U11630 (N_11630,N_6437,N_5736);
xor U11631 (N_11631,N_5534,N_6299);
xor U11632 (N_11632,N_5741,N_5378);
nor U11633 (N_11633,N_4107,N_4108);
nor U11634 (N_11634,N_4752,N_6557);
nor U11635 (N_11635,N_5194,N_7901);
nand U11636 (N_11636,N_7329,N_6281);
and U11637 (N_11637,N_5693,N_7964);
nand U11638 (N_11638,N_4308,N_6161);
xor U11639 (N_11639,N_7975,N_7258);
xor U11640 (N_11640,N_7632,N_4897);
xor U11641 (N_11641,N_4093,N_5000);
nand U11642 (N_11642,N_6847,N_4066);
nor U11643 (N_11643,N_6824,N_6099);
and U11644 (N_11644,N_6964,N_7719);
nand U11645 (N_11645,N_5401,N_4848);
nand U11646 (N_11646,N_7398,N_4177);
nand U11647 (N_11647,N_6146,N_5971);
nor U11648 (N_11648,N_4317,N_7133);
nor U11649 (N_11649,N_5075,N_7341);
xnor U11650 (N_11650,N_6866,N_4854);
xor U11651 (N_11651,N_5188,N_5332);
and U11652 (N_11652,N_6834,N_5607);
nor U11653 (N_11653,N_4362,N_5074);
and U11654 (N_11654,N_4422,N_6650);
or U11655 (N_11655,N_6903,N_5932);
or U11656 (N_11656,N_6533,N_7093);
or U11657 (N_11657,N_6427,N_6695);
and U11658 (N_11658,N_4720,N_4631);
nor U11659 (N_11659,N_7222,N_7661);
nand U11660 (N_11660,N_6481,N_7630);
xnor U11661 (N_11661,N_4225,N_6661);
and U11662 (N_11662,N_7373,N_5708);
or U11663 (N_11663,N_4595,N_6006);
nand U11664 (N_11664,N_7803,N_5054);
nor U11665 (N_11665,N_4132,N_5803);
xnor U11666 (N_11666,N_4076,N_5507);
or U11667 (N_11667,N_5995,N_7165);
xor U11668 (N_11668,N_5343,N_5460);
and U11669 (N_11669,N_6706,N_5935);
nand U11670 (N_11670,N_6943,N_4378);
or U11671 (N_11671,N_6085,N_5863);
or U11672 (N_11672,N_7915,N_4635);
nor U11673 (N_11673,N_6733,N_4765);
and U11674 (N_11674,N_7949,N_4346);
nand U11675 (N_11675,N_4915,N_7578);
nand U11676 (N_11676,N_6988,N_5621);
or U11677 (N_11677,N_6081,N_4032);
nand U11678 (N_11678,N_4882,N_4266);
nor U11679 (N_11679,N_5104,N_5088);
nand U11680 (N_11680,N_5679,N_6237);
nor U11681 (N_11681,N_4619,N_4189);
nand U11682 (N_11682,N_4972,N_6824);
or U11683 (N_11683,N_7084,N_7491);
nor U11684 (N_11684,N_6911,N_4436);
and U11685 (N_11685,N_7017,N_4403);
nor U11686 (N_11686,N_7695,N_7506);
and U11687 (N_11687,N_7224,N_5415);
xor U11688 (N_11688,N_6385,N_7773);
nor U11689 (N_11689,N_6282,N_4467);
or U11690 (N_11690,N_4716,N_7084);
and U11691 (N_11691,N_4166,N_7932);
or U11692 (N_11692,N_4973,N_7982);
nor U11693 (N_11693,N_5428,N_5519);
nand U11694 (N_11694,N_4519,N_6836);
and U11695 (N_11695,N_4483,N_7869);
nand U11696 (N_11696,N_5711,N_6884);
nand U11697 (N_11697,N_5835,N_4548);
nor U11698 (N_11698,N_5230,N_4853);
or U11699 (N_11699,N_7407,N_7887);
nand U11700 (N_11700,N_6238,N_5285);
and U11701 (N_11701,N_7090,N_5090);
or U11702 (N_11702,N_5819,N_7197);
nand U11703 (N_11703,N_4193,N_6870);
and U11704 (N_11704,N_4669,N_6429);
and U11705 (N_11705,N_4706,N_6066);
or U11706 (N_11706,N_6722,N_6580);
nor U11707 (N_11707,N_6115,N_6130);
nor U11708 (N_11708,N_7284,N_5380);
nand U11709 (N_11709,N_4092,N_4313);
xnor U11710 (N_11710,N_6606,N_4939);
nor U11711 (N_11711,N_4560,N_4471);
nand U11712 (N_11712,N_5271,N_6383);
and U11713 (N_11713,N_5254,N_7342);
nand U11714 (N_11714,N_5299,N_4819);
xnor U11715 (N_11715,N_7611,N_6935);
and U11716 (N_11716,N_7194,N_7192);
nand U11717 (N_11717,N_6815,N_7896);
nor U11718 (N_11718,N_7428,N_7389);
or U11719 (N_11719,N_7210,N_4168);
nor U11720 (N_11720,N_5181,N_7527);
or U11721 (N_11721,N_6113,N_6204);
or U11722 (N_11722,N_4646,N_5704);
nand U11723 (N_11723,N_5736,N_6507);
and U11724 (N_11724,N_4213,N_5366);
or U11725 (N_11725,N_6829,N_6017);
xor U11726 (N_11726,N_7763,N_5649);
and U11727 (N_11727,N_7653,N_6631);
nand U11728 (N_11728,N_7434,N_4022);
nand U11729 (N_11729,N_5054,N_5538);
nor U11730 (N_11730,N_4261,N_6044);
nor U11731 (N_11731,N_5743,N_7756);
xnor U11732 (N_11732,N_4139,N_5822);
nand U11733 (N_11733,N_6213,N_6985);
or U11734 (N_11734,N_5384,N_4238);
xor U11735 (N_11735,N_5735,N_7487);
xnor U11736 (N_11736,N_7260,N_4452);
nand U11737 (N_11737,N_4167,N_4844);
nor U11738 (N_11738,N_7615,N_6329);
xnor U11739 (N_11739,N_4716,N_7435);
nor U11740 (N_11740,N_4405,N_7394);
xor U11741 (N_11741,N_4744,N_5439);
nor U11742 (N_11742,N_6157,N_4602);
nand U11743 (N_11743,N_4006,N_6978);
and U11744 (N_11744,N_4702,N_7532);
and U11745 (N_11745,N_5352,N_6431);
nor U11746 (N_11746,N_5729,N_7207);
and U11747 (N_11747,N_4415,N_5259);
or U11748 (N_11748,N_5992,N_5427);
xor U11749 (N_11749,N_6397,N_7188);
nand U11750 (N_11750,N_7875,N_4556);
or U11751 (N_11751,N_6928,N_7355);
xor U11752 (N_11752,N_6254,N_4399);
xor U11753 (N_11753,N_6080,N_4000);
and U11754 (N_11754,N_4889,N_6427);
nand U11755 (N_11755,N_6830,N_6416);
nand U11756 (N_11756,N_5483,N_4923);
and U11757 (N_11757,N_6982,N_5536);
nand U11758 (N_11758,N_6822,N_5475);
xor U11759 (N_11759,N_4046,N_7740);
nor U11760 (N_11760,N_4397,N_5074);
nor U11761 (N_11761,N_6136,N_4621);
and U11762 (N_11762,N_4804,N_5550);
xor U11763 (N_11763,N_7217,N_6158);
and U11764 (N_11764,N_7452,N_6808);
xnor U11765 (N_11765,N_6294,N_5437);
xor U11766 (N_11766,N_4822,N_7959);
and U11767 (N_11767,N_7781,N_7701);
nor U11768 (N_11768,N_4902,N_5925);
xnor U11769 (N_11769,N_4374,N_6930);
nand U11770 (N_11770,N_6510,N_5010);
xnor U11771 (N_11771,N_4561,N_7577);
or U11772 (N_11772,N_5115,N_7910);
nor U11773 (N_11773,N_5615,N_5585);
nor U11774 (N_11774,N_6220,N_5047);
and U11775 (N_11775,N_6861,N_4186);
nor U11776 (N_11776,N_7045,N_6140);
nor U11777 (N_11777,N_7161,N_5287);
xor U11778 (N_11778,N_7325,N_6688);
or U11779 (N_11779,N_4854,N_4104);
xor U11780 (N_11780,N_5155,N_6537);
and U11781 (N_11781,N_7244,N_7584);
and U11782 (N_11782,N_7796,N_4991);
and U11783 (N_11783,N_4390,N_6312);
nor U11784 (N_11784,N_4738,N_4811);
or U11785 (N_11785,N_7683,N_5954);
and U11786 (N_11786,N_6602,N_7314);
nand U11787 (N_11787,N_7688,N_4336);
or U11788 (N_11788,N_6166,N_6613);
nor U11789 (N_11789,N_7689,N_4738);
or U11790 (N_11790,N_5470,N_6706);
nor U11791 (N_11791,N_4565,N_5606);
nand U11792 (N_11792,N_6186,N_5381);
or U11793 (N_11793,N_7056,N_5923);
nand U11794 (N_11794,N_5575,N_4780);
xnor U11795 (N_11795,N_5618,N_6895);
nor U11796 (N_11796,N_4983,N_4857);
nand U11797 (N_11797,N_6968,N_7623);
nor U11798 (N_11798,N_7850,N_7142);
nand U11799 (N_11799,N_7795,N_6184);
nor U11800 (N_11800,N_7663,N_7730);
xnor U11801 (N_11801,N_4400,N_7718);
and U11802 (N_11802,N_5046,N_6927);
or U11803 (N_11803,N_5920,N_4112);
and U11804 (N_11804,N_7167,N_6229);
nand U11805 (N_11805,N_4309,N_4658);
xor U11806 (N_11806,N_5248,N_6781);
and U11807 (N_11807,N_5662,N_4479);
or U11808 (N_11808,N_5114,N_7453);
and U11809 (N_11809,N_6895,N_5188);
xnor U11810 (N_11810,N_6536,N_6577);
nor U11811 (N_11811,N_5171,N_7286);
and U11812 (N_11812,N_4818,N_4549);
or U11813 (N_11813,N_4592,N_5378);
or U11814 (N_11814,N_4309,N_6665);
xor U11815 (N_11815,N_5875,N_7076);
nor U11816 (N_11816,N_4216,N_6345);
and U11817 (N_11817,N_7731,N_4505);
nor U11818 (N_11818,N_6093,N_6424);
nor U11819 (N_11819,N_4520,N_4916);
and U11820 (N_11820,N_7162,N_7381);
nand U11821 (N_11821,N_5198,N_7051);
and U11822 (N_11822,N_4046,N_6133);
nand U11823 (N_11823,N_4110,N_6248);
xor U11824 (N_11824,N_7474,N_5859);
xnor U11825 (N_11825,N_7360,N_7234);
nor U11826 (N_11826,N_4274,N_7693);
xnor U11827 (N_11827,N_4509,N_7351);
xnor U11828 (N_11828,N_7077,N_4672);
nand U11829 (N_11829,N_7654,N_7860);
xnor U11830 (N_11830,N_7962,N_6819);
and U11831 (N_11831,N_6122,N_7873);
nand U11832 (N_11832,N_7045,N_5418);
nand U11833 (N_11833,N_7991,N_4343);
nor U11834 (N_11834,N_7285,N_7981);
nor U11835 (N_11835,N_6315,N_6705);
nor U11836 (N_11836,N_7982,N_4409);
xnor U11837 (N_11837,N_7762,N_7343);
and U11838 (N_11838,N_6141,N_5037);
nor U11839 (N_11839,N_4542,N_6363);
and U11840 (N_11840,N_7079,N_4119);
or U11841 (N_11841,N_4861,N_5659);
nand U11842 (N_11842,N_4959,N_6546);
or U11843 (N_11843,N_4410,N_5769);
or U11844 (N_11844,N_6504,N_7821);
xor U11845 (N_11845,N_7048,N_6598);
nor U11846 (N_11846,N_5541,N_5105);
nor U11847 (N_11847,N_5688,N_4016);
or U11848 (N_11848,N_4261,N_4074);
and U11849 (N_11849,N_4507,N_6073);
or U11850 (N_11850,N_6695,N_7340);
xnor U11851 (N_11851,N_5047,N_5448);
xor U11852 (N_11852,N_6614,N_5599);
nor U11853 (N_11853,N_5480,N_6045);
xor U11854 (N_11854,N_5901,N_7341);
xor U11855 (N_11855,N_5593,N_5072);
xor U11856 (N_11856,N_5534,N_6914);
xnor U11857 (N_11857,N_5454,N_5660);
or U11858 (N_11858,N_7347,N_6955);
nor U11859 (N_11859,N_6256,N_7483);
nor U11860 (N_11860,N_5199,N_6644);
xor U11861 (N_11861,N_6412,N_4001);
nor U11862 (N_11862,N_7061,N_4278);
and U11863 (N_11863,N_7226,N_6164);
and U11864 (N_11864,N_4194,N_7445);
nand U11865 (N_11865,N_5514,N_4593);
or U11866 (N_11866,N_4726,N_5121);
xnor U11867 (N_11867,N_6834,N_4788);
xnor U11868 (N_11868,N_4159,N_7944);
nor U11869 (N_11869,N_5815,N_4685);
nand U11870 (N_11870,N_6322,N_5654);
and U11871 (N_11871,N_5957,N_4122);
or U11872 (N_11872,N_5742,N_4525);
or U11873 (N_11873,N_6885,N_6380);
nor U11874 (N_11874,N_6951,N_6432);
nor U11875 (N_11875,N_7554,N_7931);
nand U11876 (N_11876,N_7989,N_7255);
nor U11877 (N_11877,N_7401,N_5504);
nand U11878 (N_11878,N_4109,N_5173);
and U11879 (N_11879,N_6267,N_6369);
and U11880 (N_11880,N_4816,N_5758);
nand U11881 (N_11881,N_6243,N_4899);
nand U11882 (N_11882,N_6948,N_7290);
and U11883 (N_11883,N_6496,N_4594);
and U11884 (N_11884,N_7908,N_7575);
nand U11885 (N_11885,N_7522,N_7710);
or U11886 (N_11886,N_5187,N_6880);
or U11887 (N_11887,N_7810,N_7339);
nand U11888 (N_11888,N_5400,N_4493);
nand U11889 (N_11889,N_4958,N_4832);
nor U11890 (N_11890,N_7507,N_5299);
nand U11891 (N_11891,N_7316,N_5402);
nand U11892 (N_11892,N_5360,N_7412);
nand U11893 (N_11893,N_7306,N_4356);
nand U11894 (N_11894,N_4580,N_6095);
nand U11895 (N_11895,N_6559,N_5410);
or U11896 (N_11896,N_4049,N_7233);
nor U11897 (N_11897,N_5882,N_6817);
or U11898 (N_11898,N_4096,N_4506);
nand U11899 (N_11899,N_4211,N_4786);
xnor U11900 (N_11900,N_4520,N_4446);
nand U11901 (N_11901,N_6172,N_4920);
and U11902 (N_11902,N_7280,N_5373);
nor U11903 (N_11903,N_5848,N_5884);
and U11904 (N_11904,N_5946,N_5952);
or U11905 (N_11905,N_4968,N_7562);
and U11906 (N_11906,N_5934,N_5537);
nor U11907 (N_11907,N_5838,N_7094);
and U11908 (N_11908,N_7966,N_6376);
nor U11909 (N_11909,N_4203,N_5500);
nand U11910 (N_11910,N_6376,N_7692);
nand U11911 (N_11911,N_5290,N_7477);
and U11912 (N_11912,N_6340,N_5456);
nand U11913 (N_11913,N_4846,N_6686);
nor U11914 (N_11914,N_4997,N_5970);
and U11915 (N_11915,N_6295,N_6171);
or U11916 (N_11916,N_6132,N_7551);
and U11917 (N_11917,N_6442,N_5336);
nand U11918 (N_11918,N_6797,N_5948);
and U11919 (N_11919,N_5600,N_6253);
xnor U11920 (N_11920,N_7472,N_4612);
nand U11921 (N_11921,N_7337,N_6672);
xnor U11922 (N_11922,N_6042,N_7494);
nor U11923 (N_11923,N_7667,N_7362);
and U11924 (N_11924,N_5859,N_7643);
and U11925 (N_11925,N_5692,N_4161);
nand U11926 (N_11926,N_5060,N_5915);
xor U11927 (N_11927,N_6259,N_6837);
nand U11928 (N_11928,N_4665,N_6895);
nand U11929 (N_11929,N_4135,N_7273);
nor U11930 (N_11930,N_5172,N_6154);
nand U11931 (N_11931,N_4345,N_7529);
or U11932 (N_11932,N_5600,N_5824);
and U11933 (N_11933,N_6068,N_5223);
nor U11934 (N_11934,N_6776,N_5960);
xor U11935 (N_11935,N_4499,N_6779);
nor U11936 (N_11936,N_5584,N_6652);
or U11937 (N_11937,N_7610,N_6270);
or U11938 (N_11938,N_4203,N_5892);
nor U11939 (N_11939,N_5286,N_4780);
xnor U11940 (N_11940,N_7677,N_6932);
nand U11941 (N_11941,N_6781,N_7018);
or U11942 (N_11942,N_4406,N_5706);
or U11943 (N_11943,N_5060,N_4713);
or U11944 (N_11944,N_4513,N_5768);
or U11945 (N_11945,N_4184,N_5696);
or U11946 (N_11946,N_4353,N_4696);
and U11947 (N_11947,N_6300,N_7798);
nand U11948 (N_11948,N_6821,N_5908);
nand U11949 (N_11949,N_4432,N_6427);
or U11950 (N_11950,N_6999,N_7312);
or U11951 (N_11951,N_5727,N_5424);
xnor U11952 (N_11952,N_5354,N_7569);
and U11953 (N_11953,N_6869,N_6803);
and U11954 (N_11954,N_6841,N_4654);
nand U11955 (N_11955,N_6512,N_5675);
xor U11956 (N_11956,N_5553,N_6932);
or U11957 (N_11957,N_5374,N_4919);
or U11958 (N_11958,N_4326,N_4238);
nand U11959 (N_11959,N_5549,N_4702);
or U11960 (N_11960,N_6144,N_7121);
and U11961 (N_11961,N_7632,N_7322);
xnor U11962 (N_11962,N_7438,N_6856);
or U11963 (N_11963,N_7293,N_6370);
or U11964 (N_11964,N_6488,N_4793);
and U11965 (N_11965,N_5663,N_7064);
xnor U11966 (N_11966,N_5096,N_7243);
or U11967 (N_11967,N_4426,N_5802);
or U11968 (N_11968,N_7370,N_6234);
nand U11969 (N_11969,N_4327,N_7945);
or U11970 (N_11970,N_5043,N_4663);
or U11971 (N_11971,N_7570,N_6079);
xor U11972 (N_11972,N_7643,N_6160);
xor U11973 (N_11973,N_6723,N_7830);
or U11974 (N_11974,N_6330,N_4647);
xnor U11975 (N_11975,N_7682,N_4464);
and U11976 (N_11976,N_6654,N_5436);
or U11977 (N_11977,N_7407,N_5394);
or U11978 (N_11978,N_4191,N_5273);
or U11979 (N_11979,N_6113,N_7315);
nor U11980 (N_11980,N_4271,N_4983);
nand U11981 (N_11981,N_4080,N_6602);
or U11982 (N_11982,N_4131,N_5461);
and U11983 (N_11983,N_6045,N_4263);
or U11984 (N_11984,N_7778,N_7708);
or U11985 (N_11985,N_5937,N_4621);
nand U11986 (N_11986,N_5766,N_4588);
and U11987 (N_11987,N_6930,N_5991);
or U11988 (N_11988,N_6897,N_7253);
and U11989 (N_11989,N_6601,N_6451);
and U11990 (N_11990,N_4324,N_6162);
nor U11991 (N_11991,N_4791,N_6714);
nor U11992 (N_11992,N_7478,N_4972);
nor U11993 (N_11993,N_4768,N_6943);
nand U11994 (N_11994,N_6116,N_5107);
or U11995 (N_11995,N_6358,N_5430);
xnor U11996 (N_11996,N_5015,N_6312);
or U11997 (N_11997,N_6056,N_5017);
or U11998 (N_11998,N_6886,N_5663);
nor U11999 (N_11999,N_7045,N_6288);
and U12000 (N_12000,N_11135,N_11793);
xnor U12001 (N_12001,N_10308,N_10973);
and U12002 (N_12002,N_10289,N_10613);
nand U12003 (N_12003,N_10057,N_11147);
nor U12004 (N_12004,N_10907,N_8573);
nand U12005 (N_12005,N_10048,N_10174);
nor U12006 (N_12006,N_9917,N_11228);
nor U12007 (N_12007,N_8304,N_9272);
and U12008 (N_12008,N_11309,N_8741);
or U12009 (N_12009,N_11959,N_10855);
xnor U12010 (N_12010,N_9297,N_8324);
or U12011 (N_12011,N_11672,N_8205);
nor U12012 (N_12012,N_9466,N_8361);
or U12013 (N_12013,N_11547,N_10757);
or U12014 (N_12014,N_11012,N_9645);
and U12015 (N_12015,N_8629,N_11981);
nand U12016 (N_12016,N_9559,N_9700);
xor U12017 (N_12017,N_11446,N_9432);
xor U12018 (N_12018,N_11124,N_9424);
or U12019 (N_12019,N_10187,N_8370);
nor U12020 (N_12020,N_9288,N_11082);
nor U12021 (N_12021,N_8932,N_11339);
nand U12022 (N_12022,N_11937,N_10246);
xnor U12023 (N_12023,N_11166,N_8624);
nand U12024 (N_12024,N_9984,N_11398);
xor U12025 (N_12025,N_8257,N_9654);
or U12026 (N_12026,N_11516,N_9100);
nor U12027 (N_12027,N_9501,N_11351);
xor U12028 (N_12028,N_9863,N_10803);
xor U12029 (N_12029,N_11250,N_8434);
or U12030 (N_12030,N_8405,N_11814);
or U12031 (N_12031,N_9427,N_10843);
nor U12032 (N_12032,N_10463,N_8162);
xor U12033 (N_12033,N_9511,N_8698);
nand U12034 (N_12034,N_10767,N_10596);
and U12035 (N_12035,N_10965,N_8882);
or U12036 (N_12036,N_10001,N_10674);
and U12037 (N_12037,N_8504,N_10677);
nand U12038 (N_12038,N_8589,N_11899);
or U12039 (N_12039,N_9412,N_11257);
or U12040 (N_12040,N_8853,N_8955);
nand U12041 (N_12041,N_10029,N_11103);
or U12042 (N_12042,N_10486,N_11700);
nor U12043 (N_12043,N_8369,N_10266);
xor U12044 (N_12044,N_8283,N_9337);
xor U12045 (N_12045,N_9877,N_8725);
nor U12046 (N_12046,N_8851,N_11966);
or U12047 (N_12047,N_8497,N_9019);
nor U12048 (N_12048,N_9776,N_9249);
nor U12049 (N_12049,N_10951,N_9247);
xor U12050 (N_12050,N_11983,N_8272);
nand U12051 (N_12051,N_8436,N_8458);
or U12052 (N_12052,N_9475,N_8872);
nor U12053 (N_12053,N_10357,N_11428);
nor U12054 (N_12054,N_9349,N_8287);
nand U12055 (N_12055,N_9429,N_10250);
nor U12056 (N_12056,N_8648,N_11225);
nor U12057 (N_12057,N_11022,N_9954);
nor U12058 (N_12058,N_8663,N_10832);
nand U12059 (N_12059,N_8731,N_10570);
xnor U12060 (N_12060,N_8294,N_10205);
or U12061 (N_12061,N_9291,N_9862);
or U12062 (N_12062,N_9836,N_10884);
and U12063 (N_12063,N_10561,N_10799);
nor U12064 (N_12064,N_11549,N_10637);
or U12065 (N_12065,N_10631,N_11171);
and U12066 (N_12066,N_10894,N_8610);
nor U12067 (N_12067,N_10095,N_8373);
nor U12068 (N_12068,N_9772,N_8295);
nand U12069 (N_12069,N_11553,N_11485);
and U12070 (N_12070,N_9608,N_9464);
and U12071 (N_12071,N_8695,N_8035);
xnor U12072 (N_12072,N_8875,N_10905);
nand U12073 (N_12073,N_11435,N_9906);
xnor U12074 (N_12074,N_8511,N_10963);
xnor U12075 (N_12075,N_8661,N_9001);
nand U12076 (N_12076,N_8406,N_10685);
or U12077 (N_12077,N_9449,N_8620);
and U12078 (N_12078,N_11178,N_10571);
nor U12079 (N_12079,N_11923,N_11402);
and U12080 (N_12080,N_10504,N_9543);
xnor U12081 (N_12081,N_9164,N_8856);
or U12082 (N_12082,N_8429,N_11714);
xor U12083 (N_12083,N_8761,N_11896);
xor U12084 (N_12084,N_9675,N_9790);
or U12085 (N_12085,N_9871,N_8175);
xnor U12086 (N_12086,N_9026,N_8012);
nand U12087 (N_12087,N_8281,N_10477);
nor U12088 (N_12088,N_8630,N_9067);
xnor U12089 (N_12089,N_9218,N_9583);
or U12090 (N_12090,N_9133,N_11821);
nor U12091 (N_12091,N_11955,N_11784);
and U12092 (N_12092,N_10279,N_11445);
nor U12093 (N_12093,N_9656,N_11552);
or U12094 (N_12094,N_11872,N_11775);
xnor U12095 (N_12095,N_11709,N_9965);
or U12096 (N_12096,N_9439,N_11484);
or U12097 (N_12097,N_10554,N_9661);
and U12098 (N_12098,N_9155,N_8084);
or U12099 (N_12099,N_8049,N_11583);
xor U12100 (N_12100,N_9936,N_9185);
nand U12101 (N_12101,N_9597,N_10788);
nand U12102 (N_12102,N_9004,N_11227);
nand U12103 (N_12103,N_10460,N_9014);
or U12104 (N_12104,N_10831,N_11919);
nor U12105 (N_12105,N_10207,N_10660);
and U12106 (N_12106,N_10744,N_9097);
nor U12107 (N_12107,N_9735,N_9916);
xnor U12108 (N_12108,N_9295,N_8263);
nor U12109 (N_12109,N_9408,N_9558);
nand U12110 (N_12110,N_10420,N_11209);
or U12111 (N_12111,N_10966,N_11433);
xor U12112 (N_12112,N_11527,N_11278);
nor U12113 (N_12113,N_8172,N_10847);
nor U12114 (N_12114,N_9343,N_11990);
or U12115 (N_12115,N_9018,N_9183);
and U12116 (N_12116,N_10306,N_10382);
xor U12117 (N_12117,N_11529,N_8918);
nor U12118 (N_12118,N_11689,N_10740);
nor U12119 (N_12119,N_11002,N_8834);
or U12120 (N_12120,N_10950,N_8940);
nor U12121 (N_12121,N_8082,N_10047);
nor U12122 (N_12122,N_11436,N_11600);
nor U12123 (N_12123,N_10166,N_10569);
or U12124 (N_12124,N_8242,N_10453);
xnor U12125 (N_12125,N_11676,N_9098);
nand U12126 (N_12126,N_8948,N_9778);
or U12127 (N_12127,N_8377,N_8712);
nor U12128 (N_12128,N_8706,N_11623);
xnor U12129 (N_12129,N_9033,N_11644);
nand U12130 (N_12130,N_11790,N_9730);
nor U12131 (N_12131,N_8491,N_9973);
and U12132 (N_12132,N_8769,N_11316);
nand U12133 (N_12133,N_11076,N_11258);
nand U12134 (N_12134,N_11753,N_10114);
and U12135 (N_12135,N_10309,N_9806);
nand U12136 (N_12136,N_10506,N_8837);
or U12137 (N_12137,N_8969,N_8721);
xor U12138 (N_12138,N_10588,N_9178);
nand U12139 (N_12139,N_11439,N_8579);
and U12140 (N_12140,N_9647,N_10559);
and U12141 (N_12141,N_8785,N_8410);
or U12142 (N_12142,N_10086,N_8757);
nand U12143 (N_12143,N_11862,N_9823);
xor U12144 (N_12144,N_11144,N_9939);
nor U12145 (N_12145,N_9179,N_10818);
and U12146 (N_12146,N_8767,N_8719);
nand U12147 (N_12147,N_10734,N_10626);
nor U12148 (N_12148,N_9234,N_11046);
nor U12149 (N_12149,N_11734,N_9091);
or U12150 (N_12150,N_11964,N_8933);
nand U12151 (N_12151,N_11740,N_8789);
xor U12152 (N_12152,N_9056,N_10708);
nor U12153 (N_12153,N_10198,N_8562);
nand U12154 (N_12154,N_8705,N_9808);
nor U12155 (N_12155,N_10286,N_11570);
nand U12156 (N_12156,N_9321,N_9396);
or U12157 (N_12157,N_9054,N_10622);
xnor U12158 (N_12158,N_8156,N_11665);
and U12159 (N_12159,N_10795,N_9822);
nand U12160 (N_12160,N_9372,N_11898);
nand U12161 (N_12161,N_11168,N_9769);
nand U12162 (N_12162,N_11655,N_8805);
xor U12163 (N_12163,N_10967,N_10562);
xor U12164 (N_12164,N_10448,N_11156);
nand U12165 (N_12165,N_10703,N_10512);
and U12166 (N_12166,N_11997,N_8793);
nand U12167 (N_12167,N_8167,N_10124);
nor U12168 (N_12168,N_11337,N_11235);
nand U12169 (N_12169,N_8462,N_10438);
xor U12170 (N_12170,N_9519,N_11765);
nand U12171 (N_12171,N_10876,N_9901);
or U12172 (N_12172,N_10082,N_11755);
and U12173 (N_12173,N_11928,N_8115);
or U12174 (N_12174,N_9517,N_8245);
and U12175 (N_12175,N_11289,N_11972);
nor U12176 (N_12176,N_10028,N_9851);
nor U12177 (N_12177,N_10499,N_8148);
and U12178 (N_12178,N_10239,N_11048);
or U12179 (N_12179,N_8964,N_10919);
nand U12180 (N_12180,N_11831,N_11177);
xnor U12181 (N_12181,N_9002,N_9477);
nand U12182 (N_12182,N_8925,N_11275);
nor U12183 (N_12183,N_8604,N_10627);
xnor U12184 (N_12184,N_9109,N_10811);
xnor U12185 (N_12185,N_9262,N_8988);
and U12186 (N_12186,N_8655,N_8397);
nand U12187 (N_12187,N_11890,N_9749);
nor U12188 (N_12188,N_9191,N_11954);
xor U12189 (N_12189,N_10177,N_9542);
xor U12190 (N_12190,N_9833,N_10405);
and U12191 (N_12191,N_10396,N_10623);
and U12192 (N_12192,N_8591,N_11362);
or U12193 (N_12193,N_10635,N_9667);
or U12194 (N_12194,N_10657,N_8681);
and U12195 (N_12195,N_9145,N_9380);
and U12196 (N_12196,N_10064,N_11461);
xor U12197 (N_12197,N_10389,N_8502);
xor U12198 (N_12198,N_9505,N_8615);
nand U12199 (N_12199,N_9073,N_9677);
nand U12200 (N_12200,N_10122,N_11370);
or U12201 (N_12201,N_11030,N_8966);
xor U12202 (N_12202,N_8439,N_11538);
nand U12203 (N_12203,N_10979,N_8345);
or U12204 (N_12204,N_8994,N_9881);
nor U12205 (N_12205,N_9289,N_9705);
nand U12206 (N_12206,N_10317,N_10691);
and U12207 (N_12207,N_10084,N_9312);
xor U12208 (N_12208,N_8510,N_10327);
nand U12209 (N_12209,N_10806,N_8682);
nand U12210 (N_12210,N_9979,N_11916);
and U12211 (N_12211,N_8549,N_8337);
or U12212 (N_12212,N_11650,N_11804);
nor U12213 (N_12213,N_11089,N_11459);
nor U12214 (N_12214,N_9919,N_11377);
nand U12215 (N_12215,N_11400,N_8551);
or U12216 (N_12216,N_8599,N_8042);
nor U12217 (N_12217,N_8456,N_11957);
xor U12218 (N_12218,N_10737,N_10672);
xor U12219 (N_12219,N_8700,N_10013);
and U12220 (N_12220,N_8559,N_11546);
and U12221 (N_12221,N_8592,N_8710);
xor U12222 (N_12222,N_10595,N_10140);
and U12223 (N_12223,N_8413,N_11750);
and U12224 (N_12224,N_11332,N_11013);
nor U12225 (N_12225,N_9899,N_10071);
xor U12226 (N_12226,N_9471,N_8733);
and U12227 (N_12227,N_9199,N_11498);
nor U12228 (N_12228,N_10755,N_9679);
xnor U12229 (N_12229,N_11647,N_10826);
xnor U12230 (N_12230,N_11078,N_10742);
and U12231 (N_12231,N_10698,N_9831);
or U12232 (N_12232,N_10273,N_10036);
xnor U12233 (N_12233,N_10083,N_10654);
and U12234 (N_12234,N_10186,N_9951);
and U12235 (N_12235,N_11020,N_9669);
nand U12236 (N_12236,N_11929,N_8484);
nand U12237 (N_12237,N_8239,N_10902);
and U12238 (N_12238,N_10157,N_10406);
nor U12239 (N_12239,N_10556,N_8625);
xor U12240 (N_12240,N_9491,N_11496);
and U12241 (N_12241,N_10728,N_8357);
xnor U12242 (N_12242,N_10641,N_9142);
and U12243 (N_12243,N_9574,N_10575);
or U12244 (N_12244,N_11728,N_8829);
xnor U12245 (N_12245,N_11246,N_8611);
nor U12246 (N_12246,N_10912,N_11198);
nor U12247 (N_12247,N_8612,N_10819);
and U12248 (N_12248,N_11480,N_9923);
nor U12249 (N_12249,N_10434,N_10859);
nand U12250 (N_12250,N_10765,N_9430);
and U12251 (N_12251,N_8379,N_11738);
xor U12252 (N_12252,N_10074,N_11114);
nand U12253 (N_12253,N_9031,N_9390);
nand U12254 (N_12254,N_11083,N_10662);
nor U12255 (N_12255,N_8367,N_10000);
nand U12256 (N_12256,N_11965,N_9557);
nor U12257 (N_12257,N_8946,N_8653);
nor U12258 (N_12258,N_10194,N_9551);
nand U12259 (N_12259,N_8293,N_11961);
xnor U12260 (N_12260,N_10839,N_9339);
or U12261 (N_12261,N_8564,N_8658);
xnor U12262 (N_12262,N_8426,N_10834);
or U12263 (N_12263,N_8366,N_11540);
xnor U12264 (N_12264,N_11490,N_9999);
nor U12265 (N_12265,N_11152,N_10577);
and U12266 (N_12266,N_8024,N_9509);
and U12267 (N_12267,N_11087,N_11963);
nor U12268 (N_12268,N_10835,N_8605);
or U12269 (N_12269,N_9461,N_10123);
and U12270 (N_12270,N_10105,N_8158);
nand U12271 (N_12271,N_10299,N_9599);
or U12272 (N_12272,N_11544,N_11724);
or U12273 (N_12273,N_9589,N_8540);
nand U12274 (N_12274,N_8074,N_9307);
or U12275 (N_12275,N_11090,N_8784);
and U12276 (N_12276,N_9755,N_8586);
and U12277 (N_12277,N_11973,N_9032);
nand U12278 (N_12278,N_9607,N_11842);
nor U12279 (N_12279,N_9506,N_8895);
nor U12280 (N_12280,N_10731,N_9969);
nand U12281 (N_12281,N_9314,N_11696);
or U12282 (N_12282,N_9726,N_9022);
nor U12283 (N_12283,N_8996,N_11819);
nand U12284 (N_12284,N_11533,N_10712);
nand U12285 (N_12285,N_10175,N_8886);
nand U12286 (N_12286,N_8244,N_8139);
and U12287 (N_12287,N_10178,N_11186);
nor U12288 (N_12288,N_9839,N_11846);
xor U12289 (N_12289,N_8073,N_11904);
or U12290 (N_12290,N_8711,N_9819);
or U12291 (N_12291,N_11018,N_11486);
nand U12292 (N_12292,N_11379,N_9446);
nor U12293 (N_12293,N_10200,N_8218);
or U12294 (N_12294,N_10880,N_10464);
xor U12295 (N_12295,N_10974,N_8548);
nand U12296 (N_12296,N_11207,N_8897);
nand U12297 (N_12297,N_10805,N_10754);
or U12298 (N_12298,N_11758,N_8446);
or U12299 (N_12299,N_10344,N_8116);
nand U12300 (N_12300,N_9898,N_11868);
nor U12301 (N_12301,N_9887,N_9311);
or U12302 (N_12302,N_10391,N_10033);
xor U12303 (N_12303,N_8425,N_8038);
or U12304 (N_12304,N_9995,N_11358);
or U12305 (N_12305,N_10196,N_8544);
and U12306 (N_12306,N_10352,N_10227);
nor U12307 (N_12307,N_8000,N_10235);
xnor U12308 (N_12308,N_9629,N_8301);
nand U12309 (N_12309,N_11779,N_8971);
and U12310 (N_12310,N_9742,N_10751);
nand U12311 (N_12311,N_9886,N_11268);
xor U12312 (N_12312,N_8207,N_8529);
nand U12313 (N_12313,N_11385,N_9752);
or U12314 (N_12314,N_10517,N_9723);
xor U12315 (N_12315,N_9843,N_11707);
xor U12316 (N_12316,N_11204,N_9770);
and U12317 (N_12317,N_10376,N_11190);
nand U12318 (N_12318,N_11026,N_11052);
nor U12319 (N_12319,N_9725,N_9701);
or U12320 (N_12320,N_9930,N_10314);
or U12321 (N_12321,N_8993,N_9853);
xor U12322 (N_12322,N_11747,N_9585);
and U12323 (N_12323,N_9156,N_9125);
xor U12324 (N_12324,N_9596,N_8056);
and U12325 (N_12325,N_10021,N_10675);
xor U12326 (N_12326,N_8336,N_8223);
xnor U12327 (N_12327,N_11481,N_9024);
nor U12328 (N_12328,N_9500,N_8786);
nand U12329 (N_12329,N_10222,N_10519);
and U12330 (N_12330,N_10128,N_8449);
or U12331 (N_12331,N_8563,N_8110);
and U12332 (N_12332,N_9670,N_9365);
xor U12333 (N_12333,N_9208,N_11815);
and U12334 (N_12334,N_9784,N_11906);
nor U12335 (N_12335,N_9909,N_9550);
or U12336 (N_12336,N_10229,N_9618);
xor U12337 (N_12337,N_8122,N_8979);
nand U12338 (N_12338,N_8689,N_8654);
nor U12339 (N_12339,N_11004,N_11374);
and U12340 (N_12340,N_11824,N_9445);
or U12341 (N_12341,N_9941,N_8291);
nor U12342 (N_12342,N_11094,N_9416);
xnor U12343 (N_12343,N_10909,N_9384);
or U12344 (N_12344,N_9381,N_8776);
and U12345 (N_12345,N_10645,N_8728);
and U12346 (N_12346,N_11580,N_9369);
xnor U12347 (N_12347,N_11656,N_8327);
nand U12348 (N_12348,N_9359,N_11265);
and U12349 (N_12349,N_11160,N_11605);
and U12350 (N_12350,N_11902,N_11313);
xor U12351 (N_12351,N_9094,N_8628);
or U12352 (N_12352,N_11948,N_11652);
or U12353 (N_12353,N_10814,N_9421);
xor U12354 (N_12354,N_11708,N_9659);
or U12355 (N_12355,N_9653,N_11262);
or U12356 (N_12356,N_10355,N_8646);
nand U12357 (N_12357,N_10232,N_8537);
nand U12358 (N_12358,N_11762,N_8849);
and U12359 (N_12359,N_11736,N_10496);
xnor U12360 (N_12360,N_8550,N_8602);
nor U12361 (N_12361,N_8002,N_9874);
or U12362 (N_12362,N_10523,N_8486);
and U12363 (N_12363,N_11497,N_9143);
nand U12364 (N_12364,N_9211,N_9482);
or U12365 (N_12365,N_9630,N_9454);
nand U12366 (N_12366,N_9110,N_8739);
or U12367 (N_12367,N_10614,N_11703);
or U12368 (N_12368,N_11796,N_9912);
and U12369 (N_12369,N_10268,N_9932);
and U12370 (N_12370,N_8103,N_9872);
or U12371 (N_12371,N_9498,N_8150);
xor U12372 (N_12372,N_8393,N_11430);
or U12373 (N_12373,N_11181,N_10270);
nand U12374 (N_12374,N_11303,N_9610);
nand U12375 (N_12375,N_11763,N_8973);
xnor U12376 (N_12376,N_8417,N_10253);
nor U12377 (N_12377,N_8552,N_10202);
nor U12378 (N_12378,N_8214,N_11305);
nand U12379 (N_12379,N_11526,N_8729);
xnor U12380 (N_12380,N_11811,N_9304);
nand U12381 (N_12381,N_9021,N_10295);
xor U12382 (N_12382,N_10211,N_11891);
or U12383 (N_12383,N_9417,N_8983);
and U12384 (N_12384,N_8560,N_8346);
xnor U12385 (N_12385,N_8310,N_8161);
or U12386 (N_12386,N_9483,N_11120);
nand U12387 (N_12387,N_8905,N_9214);
and U12388 (N_12388,N_9078,N_9609);
nand U12389 (N_12389,N_11189,N_8430);
and U12390 (N_12390,N_10025,N_9260);
nor U12391 (N_12391,N_9269,N_11182);
and U12392 (N_12392,N_9783,N_11011);
and U12393 (N_12393,N_11192,N_8606);
nand U12394 (N_12394,N_8799,N_9433);
or U12395 (N_12395,N_10470,N_11193);
xor U12396 (N_12396,N_10774,N_11106);
or U12397 (N_12397,N_9452,N_10126);
and U12398 (N_12398,N_11705,N_9248);
nor U12399 (N_12399,N_9813,N_9937);
xor U12400 (N_12400,N_8222,N_10115);
nand U12401 (N_12401,N_8957,N_10764);
nor U12402 (N_12402,N_8666,N_8542);
and U12403 (N_12403,N_10241,N_11638);
or U12404 (N_12404,N_10267,N_11506);
or U12405 (N_12405,N_8618,N_11179);
nand U12406 (N_12406,N_11534,N_9059);
xor U12407 (N_12407,N_10108,N_9413);
and U12408 (N_12408,N_9130,N_11340);
and U12409 (N_12409,N_11989,N_9870);
nand U12410 (N_12410,N_8431,N_10930);
xor U12411 (N_12411,N_9401,N_8107);
and U12412 (N_12412,N_10428,N_8553);
nor U12413 (N_12413,N_8817,N_9007);
and U12414 (N_12414,N_9913,N_11849);
nand U12415 (N_12415,N_10053,N_9463);
nand U12416 (N_12416,N_8527,N_11167);
or U12417 (N_12417,N_11474,N_11914);
nor U12418 (N_12418,N_8561,N_10466);
xnor U12419 (N_12419,N_8086,N_11558);
xor U12420 (N_12420,N_11184,N_8099);
xnor U12421 (N_12421,N_11501,N_11286);
xor U12422 (N_12422,N_9182,N_10838);
nand U12423 (N_12423,N_8112,N_8105);
xnor U12424 (N_12424,N_11752,N_11597);
or U12425 (N_12425,N_9035,N_11025);
or U12426 (N_12426,N_10644,N_8171);
and U12427 (N_12427,N_8735,N_11099);
nor U12428 (N_12428,N_10233,N_9503);
nor U12429 (N_12429,N_9821,N_9860);
or U12430 (N_12430,N_11417,N_9945);
or U12431 (N_12431,N_11630,N_10706);
nor U12432 (N_12432,N_8478,N_10257);
nand U12433 (N_12433,N_8006,N_8667);
nor U12434 (N_12434,N_8095,N_9451);
xor U12435 (N_12435,N_10502,N_10667);
or U12436 (N_12436,N_9621,N_9083);
or U12437 (N_12437,N_10059,N_8688);
nor U12438 (N_12438,N_11742,N_11062);
or U12439 (N_12439,N_9761,N_8234);
xnor U12440 (N_12440,N_8928,N_8471);
xnor U12441 (N_12441,N_9244,N_10386);
nor U12442 (N_12442,N_8727,N_8202);
xor U12443 (N_12443,N_11832,N_8213);
nand U12444 (N_12444,N_10668,N_8299);
and U12445 (N_12445,N_11129,N_10432);
xnor U12446 (N_12446,N_10329,N_10103);
xor U12447 (N_12447,N_11039,N_9678);
nor U12448 (N_12448,N_9764,N_11962);
xnor U12449 (N_12449,N_8643,N_8958);
xor U12450 (N_12450,N_11933,N_11499);
or U12451 (N_12451,N_10332,N_9407);
nand U12452 (N_12452,N_10447,N_9329);
or U12453 (N_12453,N_9347,N_11881);
or U12454 (N_12454,N_10604,N_8468);
and U12455 (N_12455,N_10359,N_9717);
nand U12456 (N_12456,N_8203,N_9189);
and U12457 (N_12457,N_10829,N_8671);
nor U12458 (N_12458,N_9760,N_8773);
and U12459 (N_12459,N_10942,N_10172);
or U12460 (N_12460,N_8742,N_9231);
or U12461 (N_12461,N_9532,N_8376);
xor U12462 (N_12462,N_10601,N_11704);
nor U12463 (N_12463,N_11852,N_11231);
and U12464 (N_12464,N_10098,N_9023);
or U12465 (N_12465,N_9775,N_9318);
nor U12466 (N_12466,N_8558,N_8746);
and U12467 (N_12467,N_11851,N_9306);
and U12468 (N_12468,N_8541,N_8965);
and U12469 (N_12469,N_8864,N_9946);
xnor U12470 (N_12470,N_11095,N_9277);
and U12471 (N_12471,N_9472,N_8193);
and U12472 (N_12472,N_9338,N_8696);
nand U12473 (N_12473,N_10429,N_10969);
or U12474 (N_12474,N_11800,N_11776);
nand U12475 (N_12475,N_8692,N_8315);
or U12476 (N_12476,N_10444,N_8062);
nor U12477 (N_12477,N_9731,N_8123);
nand U12478 (N_12478,N_8396,N_11612);
nor U12479 (N_12479,N_8910,N_8296);
nor U12480 (N_12480,N_11255,N_11722);
xnor U12481 (N_12481,N_10791,N_9081);
or U12482 (N_12482,N_8435,N_10521);
and U12483 (N_12483,N_9593,N_10692);
xor U12484 (N_12484,N_11838,N_9903);
nand U12485 (N_12485,N_10955,N_8233);
or U12486 (N_12486,N_9027,N_9605);
nand U12487 (N_12487,N_10503,N_9695);
xor U12488 (N_12488,N_11589,N_10711);
nor U12489 (N_12489,N_9779,N_10243);
or U12490 (N_12490,N_11908,N_9470);
nand U12491 (N_12491,N_8642,N_9876);
xnor U12492 (N_12492,N_8052,N_8512);
xor U12493 (N_12493,N_8794,N_10209);
nor U12494 (N_12494,N_11673,N_9219);
nor U12495 (N_12495,N_9137,N_9299);
nor U12496 (N_12496,N_11871,N_8943);
or U12497 (N_12497,N_10563,N_8815);
nand U12498 (N_12498,N_9331,N_9920);
or U12499 (N_12499,N_11621,N_8515);
nand U12500 (N_12500,N_10240,N_10546);
or U12501 (N_12501,N_10097,N_9342);
or U12502 (N_12502,N_8034,N_9628);
nor U12503 (N_12503,N_8232,N_8403);
nand U12504 (N_12504,N_11487,N_11335);
nor U12505 (N_12505,N_11348,N_9548);
and U12506 (N_12506,N_11907,N_9613);
nor U12507 (N_12507,N_9163,N_9926);
nand U12508 (N_12508,N_11191,N_11284);
or U12509 (N_12509,N_10398,N_9907);
nand U12510 (N_12510,N_10899,N_9266);
nor U12511 (N_12511,N_9395,N_11127);
xor U12512 (N_12512,N_9484,N_11449);
nand U12513 (N_12513,N_8394,N_11174);
and U12514 (N_12514,N_11333,N_10639);
and U12515 (N_12515,N_8340,N_9789);
xnor U12516 (N_12516,N_11787,N_11699);
xnor U12517 (N_12517,N_11384,N_10526);
or U12518 (N_12518,N_9619,N_11737);
or U12519 (N_12519,N_10807,N_9070);
or U12520 (N_12520,N_10533,N_9444);
xnor U12521 (N_12521,N_10844,N_8745);
and U12522 (N_12522,N_11098,N_10959);
nor U12523 (N_12523,N_11925,N_9457);
nand U12524 (N_12524,N_8917,N_11014);
nand U12525 (N_12525,N_10410,N_11028);
nor U12526 (N_12526,N_8173,N_9869);
or U12527 (N_12527,N_9538,N_10006);
and U12528 (N_12528,N_8543,N_10846);
nor U12529 (N_12529,N_11783,N_10724);
nor U12530 (N_12530,N_9345,N_11967);
xor U12531 (N_12531,N_9787,N_8247);
nor U12532 (N_12532,N_9696,N_11602);
xor U12533 (N_12533,N_8069,N_9268);
and U12534 (N_12534,N_10479,N_10370);
and U12535 (N_12535,N_11802,N_9479);
xnor U12536 (N_12536,N_8603,N_10776);
nand U12537 (N_12537,N_11403,N_9368);
or U12538 (N_12538,N_10664,N_8118);
and U12539 (N_12539,N_9280,N_8483);
or U12540 (N_12540,N_11173,N_9290);
nand U12541 (N_12541,N_10061,N_8187);
nor U12542 (N_12542,N_11277,N_10032);
nand U12543 (N_12543,N_11112,N_10547);
xor U12544 (N_12544,N_9458,N_11049);
nand U12545 (N_12545,N_8229,N_10125);
or U12546 (N_12546,N_9530,N_10101);
or U12547 (N_12547,N_9927,N_11512);
nor U12548 (N_12548,N_10182,N_9341);
or U12549 (N_12549,N_10366,N_9165);
nor U12550 (N_12550,N_8622,N_8408);
xor U12551 (N_12551,N_9111,N_8530);
or U12552 (N_12552,N_11285,N_10746);
or U12553 (N_12553,N_10582,N_10958);
nand U12554 (N_12554,N_10682,N_9526);
and U12555 (N_12555,N_10558,N_10031);
xnor U12556 (N_12556,N_10137,N_8092);
or U12557 (N_12557,N_10045,N_8679);
and U12558 (N_12558,N_9437,N_9990);
xnor U12559 (N_12559,N_11613,N_11071);
nand U12560 (N_12560,N_10686,N_8952);
and U12561 (N_12561,N_8911,N_9611);
nand U12562 (N_12562,N_8869,N_11315);
or U12563 (N_12563,N_10649,N_10372);
nor U12564 (N_12564,N_11134,N_8970);
xor U12565 (N_12565,N_11903,N_11860);
nand U12566 (N_12566,N_9649,N_10848);
nor U12567 (N_12567,N_10416,N_8674);
nand U12568 (N_12568,N_9711,N_8423);
nand U12569 (N_12569,N_11476,N_9215);
nor U12570 (N_12570,N_8489,N_11507);
nand U12571 (N_12571,N_9967,N_9239);
or U12572 (N_12572,N_9614,N_11456);
xor U12573 (N_12573,N_8723,N_9317);
nor U12574 (N_12574,N_8616,N_10983);
nand U12575 (N_12575,N_8717,N_11163);
or U12576 (N_12576,N_11640,N_8019);
nor U12577 (N_12577,N_9037,N_11259);
xnor U12578 (N_12578,N_11766,N_10648);
or U12579 (N_12579,N_9225,N_11619);
or U12580 (N_12580,N_8338,N_8386);
xnor U12581 (N_12581,N_8503,N_11695);
or U12582 (N_12582,N_11319,N_11097);
xnor U12583 (N_12583,N_8221,N_11931);
xor U12584 (N_12584,N_9175,N_8378);
nand U12585 (N_12585,N_8566,N_11354);
and U12586 (N_12586,N_10565,N_10008);
nor U12587 (N_12587,N_11945,N_11205);
and U12588 (N_12588,N_9847,N_11940);
or U12589 (N_12589,N_11746,N_11222);
or U12590 (N_12590,N_8807,N_8180);
xnor U12591 (N_12591,N_11467,N_10864);
xor U12592 (N_12592,N_8126,N_9842);
nand U12593 (N_12593,N_11223,N_9328);
xor U12594 (N_12594,N_11702,N_8475);
and U12595 (N_12595,N_11847,N_9355);
nor U12596 (N_12596,N_11625,N_8358);
or U12597 (N_12597,N_9626,N_9353);
or U12598 (N_12598,N_8165,N_11888);
xor U12599 (N_12599,N_10085,N_8157);
and U12600 (N_12600,N_11109,N_9238);
nand U12601 (N_12601,N_9738,N_11560);
or U12602 (N_12602,N_8927,N_11944);
xor U12603 (N_12603,N_10535,N_9411);
or U12604 (N_12604,N_8701,N_9161);
and U12605 (N_12605,N_10615,N_8350);
nand U12606 (N_12606,N_9579,N_10271);
nand U12607 (N_12607,N_10056,N_8915);
nor U12608 (N_12608,N_11357,N_10529);
and U12609 (N_12609,N_9080,N_8372);
xor U12610 (N_12610,N_10591,N_9207);
and U12611 (N_12611,N_10713,N_11697);
nor U12612 (N_12612,N_11419,N_10075);
or U12613 (N_12613,N_9005,N_8580);
nand U12614 (N_12614,N_8136,N_10228);
or U12615 (N_12615,N_10718,N_10820);
or U12616 (N_12616,N_10952,N_10251);
xnor U12617 (N_12617,N_9719,N_9845);
and U12618 (N_12618,N_9960,N_9721);
nor U12619 (N_12619,N_8215,N_8399);
and U12620 (N_12620,N_8395,N_10112);
nand U12621 (N_12621,N_11180,N_10161);
xnor U12622 (N_12622,N_11220,N_10073);
and U12623 (N_12623,N_8102,N_8380);
and U12624 (N_12624,N_9072,N_10236);
nor U12625 (N_12625,N_8001,N_11261);
nand U12626 (N_12626,N_11162,N_10378);
xor U12627 (N_12627,N_9051,N_11007);
or U12628 (N_12628,N_8217,N_9053);
or U12629 (N_12629,N_9245,N_8098);
and U12630 (N_12630,N_11388,N_10078);
or U12631 (N_12631,N_11643,N_9236);
or U12632 (N_12632,N_10617,N_9232);
xnor U12633 (N_12633,N_9866,N_9117);
or U12634 (N_12634,N_10334,N_9071);
and U12635 (N_12635,N_8867,N_10980);
or U12636 (N_12636,N_11524,N_9642);
nand U12637 (N_12637,N_11217,N_10252);
xor U12638 (N_12638,N_9264,N_10322);
and U12639 (N_12639,N_9223,N_10374);
or U12640 (N_12640,N_9516,N_11288);
nand U12641 (N_12641,N_11185,N_11100);
nand U12642 (N_12642,N_10732,N_11988);
and U12643 (N_12643,N_11780,N_10164);
nor U12644 (N_12644,N_9241,N_11939);
xor U12645 (N_12645,N_10485,N_8258);
xnor U12646 (N_12646,N_10018,N_9844);
xnor U12647 (N_12647,N_8535,N_8758);
nand U12648 (N_12648,N_10911,N_11067);
and U12649 (N_12649,N_10516,N_8026);
nand U12650 (N_12650,N_10929,N_10011);
nor U12651 (N_12651,N_10468,N_8938);
nor U12652 (N_12652,N_11778,N_10070);
nor U12653 (N_12653,N_10651,N_8039);
nand U12654 (N_12654,N_9703,N_10995);
xnor U12655 (N_12655,N_10149,N_9048);
nand U12656 (N_12656,N_11292,N_10431);
and U12657 (N_12657,N_9030,N_9374);
and U12658 (N_12658,N_9058,N_10385);
nand U12659 (N_12659,N_11648,N_9540);
nand U12660 (N_12660,N_9782,N_10500);
or U12661 (N_12661,N_11720,N_10134);
or U12662 (N_12662,N_8037,N_9330);
xor U12663 (N_12663,N_10600,N_9216);
or U12664 (N_12664,N_11416,N_9688);
xnor U12665 (N_12665,N_8262,N_10874);
nand U12666 (N_12666,N_9710,N_9015);
xnor U12667 (N_12667,N_9332,N_8487);
and U12668 (N_12668,N_11713,N_9573);
or U12669 (N_12669,N_9652,N_11057);
or U12670 (N_12670,N_9774,N_11483);
or U12671 (N_12671,N_11041,N_9780);
nor U12672 (N_12672,N_9816,N_8833);
or U12673 (N_12673,N_11617,N_11047);
or U12674 (N_12674,N_9298,N_9003);
nor U12675 (N_12675,N_11883,N_10508);
or U12676 (N_12676,N_9282,N_11215);
xor U12677 (N_12677,N_11024,N_11008);
nor U12678 (N_12678,N_11325,N_8320);
or U12679 (N_12679,N_9859,N_9807);
or U12680 (N_12680,N_9278,N_10399);
and U12681 (N_12681,N_9838,N_9508);
nand U12682 (N_12682,N_8931,N_9074);
or U12683 (N_12683,N_8188,N_8677);
nor U12684 (N_12684,N_11006,N_10851);
nor U12685 (N_12685,N_11146,N_11917);
nand U12686 (N_12686,N_11301,N_11300);
nand U12687 (N_12687,N_11457,N_10527);
nand U12688 (N_12688,N_10189,N_11987);
nand U12689 (N_12689,N_11397,N_8210);
nor U12690 (N_12690,N_10625,N_10816);
xnor U12691 (N_12691,N_10867,N_10403);
and U12692 (N_12692,N_11693,N_11263);
or U12693 (N_12693,N_11145,N_8220);
and U12694 (N_12694,N_9697,N_9256);
and U12695 (N_12695,N_11718,N_8241);
or U12696 (N_12696,N_11934,N_9617);
and U12697 (N_12697,N_9894,N_8754);
xor U12698 (N_12698,N_8960,N_8490);
and U12699 (N_12699,N_8694,N_10079);
and U12700 (N_12700,N_11971,N_10418);
or U12701 (N_12701,N_10763,N_8982);
nand U12702 (N_12702,N_10646,N_11375);
and U12703 (N_12703,N_8470,N_8619);
nand U12704 (N_12704,N_10199,N_9134);
nor U12705 (N_12705,N_9443,N_8120);
or U12706 (N_12706,N_11281,N_8195);
nand U12707 (N_12707,N_10735,N_10379);
xnor U12708 (N_12708,N_8067,N_8756);
or U12709 (N_12709,N_10495,N_9283);
or U12710 (N_12710,N_11170,N_9754);
and U12711 (N_12711,N_11827,N_11294);
or U12712 (N_12712,N_9420,N_11777);
nand U12713 (N_12713,N_9102,N_8797);
and U12714 (N_12714,N_10766,N_11603);
and U12715 (N_12715,N_9402,N_11998);
nor U12716 (N_12716,N_11218,N_10191);
nand U12717 (N_12717,N_8868,N_9017);
or U12718 (N_12718,N_11343,N_9360);
nor U12719 (N_12719,N_11835,N_9552);
xor U12720 (N_12720,N_9316,N_11611);
nor U12721 (N_12721,N_11251,N_8312);
and U12722 (N_12722,N_11606,N_9173);
xor U12723 (N_12723,N_10609,N_10551);
or U12724 (N_12724,N_10055,N_8028);
nor U12725 (N_12725,N_10462,N_9915);
and U12726 (N_12726,N_10594,N_10323);
nor U12727 (N_12727,N_9956,N_10046);
xor U12728 (N_12728,N_11770,N_10782);
and U12729 (N_12729,N_8230,N_10883);
and U12730 (N_12730,N_10738,N_8859);
nand U12731 (N_12731,N_11040,N_9386);
or U12732 (N_12732,N_9305,N_11684);
and U12733 (N_12733,N_11329,N_8228);
or U12734 (N_12734,N_9529,N_8879);
nor U12735 (N_12735,N_8224,N_8828);
nand U12736 (N_12736,N_10469,N_9057);
xnor U12737 (N_12737,N_8058,N_11615);
xor U12738 (N_12738,N_8494,N_8297);
nand U12739 (N_12739,N_10170,N_11420);
or U12740 (N_12740,N_9150,N_11202);
nand U12741 (N_12741,N_9485,N_11440);
nand U12742 (N_12742,N_11404,N_10093);
nor U12743 (N_12743,N_11216,N_8876);
nor U12744 (N_12744,N_10455,N_10193);
nor U12745 (N_12745,N_8212,N_9891);
nand U12746 (N_12746,N_11065,N_8862);
nor U12747 (N_12747,N_9837,N_11153);
or U12748 (N_12748,N_8990,N_11667);
or U12749 (N_12749,N_8806,N_9541);
or U12750 (N_12750,N_10714,N_9180);
or U12751 (N_12751,N_9709,N_8392);
or U12752 (N_12752,N_9497,N_9625);
or U12753 (N_12753,N_10278,N_8045);
nor U12754 (N_12754,N_8743,N_9534);
nor U12755 (N_12755,N_10262,N_10536);
and U12756 (N_12756,N_8730,N_8474);
nand U12757 (N_12757,N_8569,N_9113);
and U12758 (N_12758,N_11296,N_11401);
nand U12759 (N_12759,N_9040,N_10568);
or U12760 (N_12760,N_9085,N_11968);
and U12761 (N_12761,N_11282,N_8186);
xor U12762 (N_12762,N_8108,N_8921);
nand U12763 (N_12763,N_10301,N_11561);
or U12764 (N_12764,N_11308,N_9882);
nor U12765 (N_12765,N_10892,N_11594);
and U12766 (N_12766,N_8924,N_9972);
or U12767 (N_12767,N_9949,N_9467);
nand U12768 (N_12768,N_11579,N_10442);
and U12769 (N_12769,N_11108,N_11244);
xor U12770 (N_12770,N_10155,N_10590);
or U12771 (N_12771,N_11659,N_11576);
xnor U12772 (N_12772,N_11508,N_10217);
nand U12773 (N_12773,N_10597,N_8521);
nand U12774 (N_12774,N_11344,N_9205);
nand U12775 (N_12775,N_9884,N_11175);
xor U12776 (N_12776,N_11794,N_11877);
nor U12777 (N_12777,N_10143,N_8791);
nor U12778 (N_12778,N_8164,N_10050);
and U12779 (N_12779,N_11588,N_9692);
and U12780 (N_12780,N_10815,N_9865);
or U12781 (N_12781,N_11117,N_10077);
nand U12782 (N_12782,N_10548,N_10787);
nand U12783 (N_12783,N_10810,N_10783);
xor U12784 (N_12784,N_8319,N_8104);
and U12785 (N_12785,N_8804,N_11462);
xor U12786 (N_12786,N_8321,N_9680);
nand U12787 (N_12787,N_9181,N_10413);
nor U12788 (N_12788,N_8441,N_8017);
xor U12789 (N_12789,N_11023,N_10505);
nor U12790 (N_12790,N_11726,N_8722);
nor U12791 (N_12791,N_10671,N_10984);
and U12792 (N_12792,N_9193,N_9377);
nand U12793 (N_12793,N_10784,N_11882);
nand U12794 (N_12794,N_9885,N_9136);
or U12795 (N_12795,N_10210,N_8636);
nor U12796 (N_12796,N_8131,N_8457);
or U12797 (N_12797,N_9796,N_9442);
nand U12798 (N_12798,N_8125,N_9950);
or U12799 (N_12799,N_9904,N_11515);
and U12800 (N_12800,N_9803,N_11645);
or U12801 (N_12801,N_9632,N_8669);
and U12802 (N_12802,N_11169,N_11649);
or U12803 (N_12803,N_8114,N_8763);
nor U12804 (N_12804,N_10017,N_9962);
nor U12805 (N_12805,N_9810,N_10044);
nand U12806 (N_12806,N_8855,N_10132);
nand U12807 (N_12807,N_9580,N_8040);
or U12808 (N_12808,N_10213,N_9537);
or U12809 (N_12809,N_8060,N_10135);
nand U12810 (N_12810,N_9861,N_8194);
nor U12811 (N_12811,N_11247,N_10861);
nor U12812 (N_12812,N_10484,N_11031);
and U12813 (N_12813,N_10067,N_11042);
nand U12814 (N_12814,N_10009,N_9817);
or U12815 (N_12815,N_9555,N_9729);
xnor U12816 (N_12816,N_8285,N_9379);
or U12817 (N_12817,N_10515,N_9985);
or U12818 (N_12818,N_9747,N_10195);
or U12819 (N_12819,N_9116,N_11367);
and U12820 (N_12820,N_10350,N_9327);
nor U12821 (N_12821,N_9947,N_11230);
and U12822 (N_12822,N_8787,N_8400);
nor U12823 (N_12823,N_10375,N_9481);
or U12824 (N_12824,N_8963,N_9952);
or U12825 (N_12825,N_8335,N_9988);
or U12826 (N_12826,N_11312,N_10647);
nor U12827 (N_12827,N_10870,N_10305);
xnor U12828 (N_12828,N_11555,N_11608);
nand U12829 (N_12829,N_8387,N_11138);
nand U12830 (N_12830,N_9896,N_8499);
and U12831 (N_12831,N_8750,N_9131);
xor U12832 (N_12832,N_11347,N_11196);
xor U12833 (N_12833,N_8809,N_11328);
nand U12834 (N_12834,N_8704,N_8514);
nand U12835 (N_12835,N_11646,N_11927);
and U12836 (N_12836,N_11844,N_11635);
nand U12837 (N_12837,N_9567,N_9435);
nand U12838 (N_12838,N_11488,N_9624);
xor U12839 (N_12839,N_9814,N_10524);
nand U12840 (N_12840,N_11273,N_10878);
nor U12841 (N_12841,N_10828,N_11422);
nand U12842 (N_12842,N_11918,N_8974);
or U12843 (N_12843,N_11241,N_10566);
xnor U12844 (N_12844,N_8967,N_8351);
nand U12845 (N_12845,N_9476,N_9334);
and U12846 (N_12846,N_10842,N_8831);
nor U12847 (N_12847,N_11033,N_8277);
or U12848 (N_12848,N_8816,N_10336);
or U12849 (N_12849,N_11234,N_10208);
nand U12850 (N_12850,N_8440,N_10365);
nor U12851 (N_12851,N_10106,N_11164);
xnor U12852 (N_12852,N_10642,N_8571);
or U12853 (N_12853,N_8053,N_9734);
xor U12854 (N_12854,N_9044,N_10060);
and U12855 (N_12855,N_8626,N_8482);
and U12856 (N_12856,N_11390,N_9724);
nor U12857 (N_12857,N_10868,N_9897);
xnor U12858 (N_12858,N_9856,N_10401);
nand U12859 (N_12859,N_9079,N_10886);
and U12860 (N_12860,N_8326,N_10457);
or U12861 (N_12861,N_11016,N_9086);
or U12862 (N_12862,N_10092,N_11123);
or U12863 (N_12863,N_9197,N_10887);
or U12864 (N_12864,N_9096,N_11366);
or U12865 (N_12865,N_10761,N_8880);
nor U12866 (N_12866,N_11980,N_9924);
and U12867 (N_12867,N_8526,N_8149);
nand U12868 (N_12868,N_10522,N_9398);
and U12869 (N_12869,N_8830,N_9310);
or U12870 (N_12870,N_8072,N_9468);
nor U12871 (N_12871,N_11797,N_8684);
nor U12872 (N_12872,N_11566,N_11463);
or U12873 (N_12873,N_11637,N_11743);
xor U12874 (N_12874,N_11056,N_10404);
nor U12875 (N_12875,N_10397,N_10338);
nor U12876 (N_12876,N_10180,N_9363);
and U12877 (N_12877,N_9522,N_8556);
nor U12878 (N_12878,N_8708,N_9034);
and U12879 (N_12879,N_8896,N_10552);
nor U12880 (N_12880,N_10809,N_8237);
nand U12881 (N_12881,N_10578,N_8355);
nand U12882 (N_12882,N_8584,N_10415);
and U12883 (N_12883,N_10914,N_10653);
nor U12884 (N_12884,N_9228,N_10333);
xor U12885 (N_12885,N_11036,N_11856);
nor U12886 (N_12886,N_8812,N_10822);
and U12887 (N_12887,N_9883,N_8022);
and U12888 (N_12888,N_10096,N_8536);
xor U12889 (N_12889,N_10099,N_10245);
nor U12890 (N_12890,N_10272,N_8138);
or U12891 (N_12891,N_10659,N_8984);
and U12892 (N_12892,N_9184,N_8783);
and U12893 (N_12893,N_9644,N_10610);
or U12894 (N_12894,N_8328,N_8051);
and U12895 (N_12895,N_10091,N_10043);
xnor U12896 (N_12896,N_11686,N_11287);
nand U12897 (N_12897,N_11077,N_8518);
or U12898 (N_12898,N_8877,N_11050);
nand U12899 (N_12899,N_9459,N_9082);
nand U12900 (N_12900,N_8881,N_11341);
and U12901 (N_12901,N_10445,N_9828);
and U12902 (N_12902,N_9751,N_8079);
xnor U12903 (N_12903,N_11751,N_10749);
nor U12904 (N_12904,N_11817,N_8308);
nor U12905 (N_12905,N_10298,N_8904);
xor U12906 (N_12906,N_9604,N_11032);
or U12907 (N_12907,N_10040,N_8445);
nand U12908 (N_12908,N_10530,N_11053);
nor U12909 (N_12909,N_8479,N_10537);
nand U12910 (N_12910,N_8753,N_11475);
or U12911 (N_12911,N_9938,N_10845);
nand U12912 (N_12912,N_8209,N_10857);
and U12913 (N_12913,N_9170,N_10318);
or U12914 (N_12914,N_11363,N_9084);
nor U12915 (N_12915,N_10088,N_10291);
or U12916 (N_12916,N_8765,N_10019);
and U12917 (N_12917,N_8623,N_8339);
nand U12918 (N_12918,N_9975,N_10585);
and U12919 (N_12919,N_11666,N_10801);
xnor U12920 (N_12920,N_11116,N_10394);
nand U12921 (N_12921,N_9303,N_10821);
nand U12922 (N_12922,N_11710,N_11113);
nor U12923 (N_12923,N_8939,N_10118);
nor U12924 (N_12924,N_8307,N_10917);
or U12925 (N_12925,N_11833,N_11632);
or U12926 (N_12926,N_11590,N_11051);
xor U12927 (N_12927,N_8041,N_8892);
nand U12928 (N_12928,N_10107,N_8811);
xor U12929 (N_12929,N_8013,N_11574);
and U12930 (N_12930,N_8243,N_11346);
or U12931 (N_12931,N_11599,N_8135);
nand U12932 (N_12932,N_10743,N_8235);
nand U12933 (N_12933,N_9367,N_10534);
and U12934 (N_12934,N_8737,N_11805);
nor U12935 (N_12935,N_10999,N_10297);
nor U12936 (N_12936,N_11295,N_9875);
or U12937 (N_12937,N_8178,N_11447);
nor U12938 (N_12938,N_10068,N_8699);
and U12939 (N_12939,N_11843,N_9622);
and U12940 (N_12940,N_11314,N_10129);
or U12941 (N_12941,N_10921,N_10572);
nor U12942 (N_12942,N_11975,N_10242);
xor U12943 (N_12943,N_10699,N_11055);
xor U12944 (N_12944,N_11748,N_11809);
or U12945 (N_12945,N_9699,N_9301);
nand U12946 (N_12946,N_9281,N_10281);
nor U12947 (N_12947,N_11542,N_10435);
nor U12948 (N_12948,N_8063,N_10244);
nor U12949 (N_12949,N_11941,N_11756);
and U12950 (N_12950,N_10369,N_10422);
and U12951 (N_12951,N_11759,N_10472);
nor U12952 (N_12952,N_8702,N_10311);
nor U12953 (N_12953,N_10156,N_11248);
nand U12954 (N_12954,N_11812,N_11880);
or U12955 (N_12955,N_9714,N_11541);
nor U12956 (N_12956,N_8587,N_10335);
or U12957 (N_12957,N_9112,N_8375);
and U12958 (N_12958,N_8991,N_8402);
nor U12959 (N_12959,N_8300,N_10022);
xor U12960 (N_12960,N_8909,N_11233);
nand U12961 (N_12961,N_11505,N_8197);
xnor U12962 (N_12962,N_11360,N_8595);
xnor U12963 (N_12963,N_9404,N_11415);
nor U12964 (N_12964,N_11893,N_9315);
nor U12965 (N_12965,N_9740,N_10608);
and U12966 (N_12966,N_8500,N_8176);
and U12967 (N_12967,N_9050,N_9460);
xnor U12968 (N_12968,N_11003,N_9284);
nor U12969 (N_12969,N_9641,N_9544);
or U12970 (N_12970,N_9495,N_11674);
or U12971 (N_12971,N_9263,N_9233);
nand U12972 (N_12972,N_11905,N_11493);
nand U12973 (N_12973,N_8447,N_8352);
or U12974 (N_12974,N_8046,N_9673);
or U12975 (N_12975,N_11500,N_10932);
or U12976 (N_12976,N_10991,N_10491);
xor U12977 (N_12977,N_8748,N_10856);
or U12978 (N_12978,N_11291,N_10866);
xor U12979 (N_12979,N_9286,N_9977);
nand U12980 (N_12980,N_9132,N_9092);
nor U12981 (N_12981,N_11869,N_11545);
nor U12982 (N_12982,N_10058,N_10873);
nor U12983 (N_12983,N_10321,N_11556);
nand U12984 (N_12984,N_11212,N_10087);
and U12985 (N_12985,N_8182,N_10538);
xnor U12986 (N_12986,N_11735,N_8011);
or U12987 (N_12987,N_11070,N_10450);
nand U12988 (N_12988,N_9728,N_8574);
or U12989 (N_12989,N_9545,N_10993);
or U12990 (N_12990,N_11976,N_9594);
nand U12991 (N_12991,N_11376,N_9115);
xnor U12992 (N_12992,N_9657,N_11969);
and U12993 (N_12993,N_11425,N_9631);
nand U12994 (N_12994,N_8848,N_8885);
xor U12995 (N_12995,N_11086,N_9253);
xor U12996 (N_12996,N_11072,N_10023);
or U12997 (N_12997,N_8585,N_10439);
nand U12998 (N_12998,N_10237,N_8651);
and U12999 (N_12999,N_8023,N_10775);
xor U13000 (N_13000,N_11518,N_10249);
and U13001 (N_13001,N_11816,N_11468);
nand U13002 (N_13002,N_8065,N_10218);
and U13003 (N_13003,N_9640,N_10363);
and U13004 (N_13004,N_8808,N_8360);
or U13005 (N_13005,N_11788,N_8368);
or U13006 (N_13006,N_10039,N_10409);
or U13007 (N_13007,N_9646,N_9160);
and U13008 (N_13008,N_8048,N_10388);
and U13009 (N_13009,N_8121,N_11627);
xnor U13010 (N_13010,N_8168,N_9168);
or U13011 (N_13011,N_8937,N_8290);
xnor U13012 (N_13012,N_10408,N_9135);
nor U13013 (N_13013,N_10707,N_9296);
and U13014 (N_13014,N_11381,N_10316);
nor U13015 (N_13015,N_11651,N_9765);
xnor U13016 (N_13016,N_8090,N_11364);
or U13017 (N_13017,N_11960,N_9006);
or U13018 (N_13018,N_11523,N_9996);
and U13019 (N_13019,N_9419,N_10633);
xor U13020 (N_13020,N_8467,N_11478);
xor U13021 (N_13021,N_11310,N_8461);
and U13022 (N_13022,N_11211,N_11993);
and U13023 (N_13023,N_10915,N_9258);
nand U13024 (N_13024,N_9651,N_10015);
or U13025 (N_13025,N_10889,N_10300);
and U13026 (N_13026,N_9637,N_9490);
nor U13027 (N_13027,N_10072,N_10998);
and U13028 (N_13028,N_8520,N_9690);
nor U13029 (N_13029,N_11949,N_10931);
and U13030 (N_13030,N_9835,N_9455);
xor U13031 (N_13031,N_10904,N_9128);
nor U13032 (N_13032,N_8155,N_8691);
nor U13033 (N_13033,N_8889,N_8068);
nor U13034 (N_13034,N_9388,N_10414);
nor U13035 (N_13035,N_9438,N_8657);
xor U13036 (N_13036,N_10800,N_9715);
nor U13037 (N_13037,N_8513,N_11214);
xnor U13038 (N_13038,N_9944,N_11575);
nor U13039 (N_13039,N_10340,N_9400);
xnor U13040 (N_13040,N_11038,N_9713);
xnor U13041 (N_13041,N_10313,N_11183);
and U13042 (N_13042,N_9867,N_11064);
nor U13043 (N_13043,N_8317,N_9858);
and U13044 (N_13044,N_8976,N_11119);
nand U13045 (N_13045,N_10430,N_8260);
xor U13046 (N_13046,N_11359,N_9361);
nor U13047 (N_13047,N_8601,N_11682);
xnor U13048 (N_13048,N_10402,N_8813);
and U13049 (N_13049,N_10638,N_11706);
nand U13050 (N_13050,N_11154,N_10133);
nand U13051 (N_13051,N_11491,N_8534);
nand U13052 (N_13052,N_10081,N_8935);
nor U13053 (N_13053,N_10827,N_8274);
or U13054 (N_13054,N_8863,N_9987);
and U13055 (N_13055,N_8803,N_8033);
xor U13056 (N_13056,N_10049,N_8179);
or U13057 (N_13057,N_11471,N_11254);
and U13058 (N_13058,N_10665,N_8775);
nor U13059 (N_13059,N_9756,N_10947);
nand U13060 (N_13060,N_10897,N_10310);
xnor U13061 (N_13061,N_9202,N_10607);
nand U13062 (N_13062,N_8077,N_10852);
and U13063 (N_13063,N_11151,N_10616);
nand U13064 (N_13064,N_9294,N_9302);
and U13065 (N_13065,N_9595,N_8609);
nand U13066 (N_13066,N_10024,N_8588);
xnor U13067 (N_13067,N_9512,N_9982);
nor U13068 (N_13068,N_9576,N_8344);
nand U13069 (N_13069,N_9357,N_9042);
or U13070 (N_13070,N_10640,N_8465);
nor U13071 (N_13071,N_8050,N_10474);
and U13072 (N_13072,N_8818,N_8614);
xor U13073 (N_13073,N_11520,N_11530);
nor U13074 (N_13074,N_11598,N_11754);
or U13075 (N_13075,N_10197,N_8253);
xor U13076 (N_13076,N_10989,N_10910);
and U13077 (N_13077,N_10158,N_8772);
or U13078 (N_13078,N_8525,N_9203);
xnor U13079 (N_13079,N_8565,N_9169);
or U13080 (N_13080,N_10119,N_10769);
nor U13081 (N_13081,N_9694,N_11015);
or U13082 (N_13082,N_10307,N_9154);
or U13083 (N_13083,N_8343,N_11626);
nor U13084 (N_13084,N_10264,N_9061);
and U13085 (N_13085,N_8198,N_10282);
nor U13086 (N_13086,N_11395,N_11409);
nand U13087 (N_13087,N_11823,N_11884);
nand U13088 (N_13088,N_9394,N_11539);
or U13089 (N_13089,N_8433,N_10159);
or U13090 (N_13090,N_9118,N_10656);
xnor U13091 (N_13091,N_9959,N_10934);
or U13092 (N_13092,N_10320,N_9536);
nor U13093 (N_13093,N_10720,N_9144);
nand U13094 (N_13094,N_10263,N_9063);
and U13095 (N_13095,N_11317,N_10680);
or U13096 (N_13096,N_8225,N_10727);
or U13097 (N_13097,N_9553,N_9171);
and U13098 (N_13098,N_10550,N_11460);
and U13099 (N_13099,N_9423,N_11806);
xnor U13100 (N_13100,N_8495,N_10296);
nand U13101 (N_13101,N_11239,N_10666);
xor U13102 (N_13102,N_8267,N_9352);
xnor U13103 (N_13103,N_11822,N_11396);
or U13104 (N_13104,N_9706,N_11732);
or U13105 (N_13105,N_9201,N_11330);
xor U13106 (N_13106,N_9854,N_8524);
nand U13107 (N_13107,N_10789,N_11892);
xor U13108 (N_13108,N_11290,N_11874);
nand U13109 (N_13109,N_11494,N_10802);
xnor U13110 (N_13110,N_10697,N_9743);
and U13111 (N_13111,N_8720,N_11088);
and U13112 (N_13112,N_11280,N_8903);
nand U13113 (N_13113,N_8453,N_8823);
nand U13114 (N_13114,N_11010,N_10634);
nand U13115 (N_13115,N_11922,N_11636);
nor U13116 (N_13116,N_11930,N_8989);
xnor U13117 (N_13117,N_10507,N_9188);
nand U13118 (N_13118,N_10812,N_10762);
nand U13119 (N_13119,N_8633,N_11876);
and U13120 (N_13120,N_9088,N_8388);
xor U13121 (N_13121,N_10437,N_8054);
xor U13122 (N_13122,N_11875,N_9992);
nor U13123 (N_13123,N_10918,N_10598);
or U13124 (N_13124,N_11355,N_8557);
nand U13125 (N_13125,N_9745,N_11452);
or U13126 (N_13126,N_10138,N_10150);
or U13127 (N_13127,N_8418,N_11005);
and U13128 (N_13128,N_11604,N_10778);
nor U13129 (N_13129,N_9864,N_8259);
and U13130 (N_13130,N_11272,N_10722);
and U13131 (N_13131,N_11999,N_9744);
xnor U13132 (N_13132,N_9757,N_8266);
xor U13133 (N_13133,N_10162,N_10684);
nor U13134 (N_13134,N_8954,N_11311);
xnor U13135 (N_13135,N_11423,N_10154);
or U13136 (N_13136,N_11813,N_9221);
xnor U13137 (N_13137,N_10825,N_11454);
nand U13138 (N_13138,N_9428,N_10953);
and U13139 (N_13139,N_9655,N_9591);
or U13140 (N_13140,N_9792,N_11798);
xnor U13141 (N_13141,N_9643,N_8081);
nand U13142 (N_13142,N_8030,N_11698);
or U13143 (N_13143,N_9786,N_8822);
xor U13144 (N_13144,N_9791,N_10772);
nor U13145 (N_13145,N_9146,N_8738);
and U13146 (N_13146,N_8945,N_9958);
nor U13147 (N_13147,N_10509,N_8778);
nor U13148 (N_13148,N_10557,N_11532);
nor U13149 (N_13149,N_9616,N_8975);
xnor U13150 (N_13150,N_10939,N_8124);
xor U13151 (N_13151,N_9313,N_10717);
and U13152 (N_13152,N_9261,N_8608);
and U13153 (N_13153,N_10461,N_8036);
xor U13154 (N_13154,N_8929,N_10473);
or U13155 (N_13155,N_9612,N_10837);
and U13156 (N_13156,N_10804,N_9008);
xnor U13157 (N_13157,N_11986,N_11322);
and U13158 (N_13158,N_9344,N_10274);
and U13159 (N_13159,N_8238,N_10906);
or U13160 (N_13160,N_10497,N_8064);
or U13161 (N_13161,N_8009,N_9356);
or U13162 (N_13162,N_9525,N_8890);
and U13163 (N_13163,N_10721,N_11394);
and U13164 (N_13164,N_10110,N_11828);
nor U13165 (N_13165,N_10606,N_10510);
nor U13166 (N_13166,N_11091,N_8858);
nor U13167 (N_13167,N_9486,N_10144);
nand U13168 (N_13168,N_9980,N_8744);
nor U13169 (N_13169,N_8845,N_11996);
xnor U13170 (N_13170,N_9456,N_11642);
xnor U13171 (N_13171,N_10773,N_8726);
and U13172 (N_13172,N_9047,N_10900);
and U13173 (N_13173,N_10676,N_11910);
nand U13174 (N_13174,N_8652,N_11938);
nand U13175 (N_13175,N_10142,N_9415);
xor U13176 (N_13176,N_10035,N_11681);
and U13177 (N_13177,N_8174,N_10544);
nand U13178 (N_13178,N_8286,N_11378);
nand U13179 (N_13179,N_11567,N_10065);
nand U13180 (N_13180,N_9240,N_11932);
nand U13181 (N_13181,N_9900,N_9777);
nor U13182 (N_13182,N_8061,N_8101);
nand U13183 (N_13183,N_8531,N_8501);
nand U13184 (N_13184,N_9217,N_9737);
xnor U13185 (N_13185,N_10377,N_9592);
nor U13186 (N_13186,N_9166,N_9251);
or U13187 (N_13187,N_9409,N_11901);
nor U13188 (N_13188,N_8678,N_9246);
nand U13189 (N_13189,N_11723,N_8313);
and U13190 (N_13190,N_9830,N_9087);
and U13191 (N_13191,N_9931,N_8860);
nand U13192 (N_13192,N_10380,N_11950);
nor U13193 (N_13193,N_8878,N_10304);
or U13194 (N_13194,N_10619,N_11855);
nand U13195 (N_13195,N_8840,N_11021);
nor U13196 (N_13196,N_8752,N_10944);
or U13197 (N_13197,N_11392,N_8496);
nor U13198 (N_13198,N_11554,N_9974);
or U13199 (N_13199,N_10968,N_8498);
nor U13200 (N_13200,N_8365,N_11001);
nor U13201 (N_13201,N_9758,N_10339);
nor U13202 (N_13202,N_9362,N_10488);
xor U13203 (N_13203,N_11837,N_11240);
or U13204 (N_13204,N_8509,N_10171);
or U13205 (N_13205,N_9978,N_10454);
or U13206 (N_13206,N_10525,N_9448);
nand U13207 (N_13207,N_9741,N_10863);
and U13208 (N_13208,N_10337,N_9487);
and U13209 (N_13209,N_10183,N_11745);
nand U13210 (N_13210,N_11513,N_9148);
or U13211 (N_13211,N_11653,N_8389);
nand U13212 (N_13212,N_8507,N_8716);
nor U13213 (N_13213,N_8740,N_8874);
nand U13214 (N_13214,N_9060,N_8519);
xnor U13215 (N_13215,N_9935,N_11629);
xnor U13216 (N_13216,N_11412,N_8707);
and U13217 (N_13217,N_8555,N_10975);
nor U13218 (N_13218,N_9852,N_10518);
nor U13219 (N_13219,N_10997,N_11767);
nand U13220 (N_13220,N_11349,N_11825);
or U13221 (N_13221,N_11307,N_11455);
xnor U13222 (N_13222,N_11913,N_10113);
or U13223 (N_13223,N_11935,N_11194);
nand U13224 (N_13224,N_10690,N_10695);
or U13225 (N_13225,N_11841,N_11079);
or U13226 (N_13226,N_8407,N_10725);
nor U13227 (N_13227,N_11489,N_8883);
nand U13228 (N_13228,N_10964,N_10943);
nor U13229 (N_13229,N_9152,N_10937);
xnor U13230 (N_13230,N_11102,N_10986);
xnor U13231 (N_13231,N_8318,N_11610);
and U13232 (N_13232,N_10100,N_8177);
and U13233 (N_13233,N_10630,N_10130);
xnor U13234 (N_13234,N_8533,N_10520);
or U13235 (N_13235,N_8117,N_8032);
and U13236 (N_13236,N_9123,N_10632);
nand U13237 (N_13237,N_8777,N_9383);
nor U13238 (N_13238,N_8044,N_9910);
xnor U13239 (N_13239,N_8353,N_11537);
nand U13240 (N_13240,N_8788,N_8523);
nor U13241 (N_13241,N_8770,N_8656);
nand U13242 (N_13242,N_11658,N_9683);
or U13243 (N_13243,N_8759,N_8085);
or U13244 (N_13244,N_11719,N_8273);
nor U13245 (N_13245,N_9308,N_10970);
nor U13246 (N_13246,N_10465,N_9496);
nand U13247 (N_13247,N_9274,N_9375);
nor U13248 (N_13248,N_11717,N_8422);
nor U13249 (N_13249,N_10758,N_8912);
xor U13250 (N_13250,N_8027,N_11338);
nor U13251 (N_13251,N_10513,N_11878);
nand U13252 (N_13252,N_9000,N_11101);
and U13253 (N_13253,N_9566,N_11886);
nor U13254 (N_13254,N_8986,N_10862);
and U13255 (N_13255,N_10269,N_10841);
or U13256 (N_13256,N_9068,N_10926);
and U13257 (N_13257,N_9664,N_8169);
or U13258 (N_13258,N_11578,N_9981);
nand U13259 (N_13259,N_9797,N_11469);
nor U13260 (N_13260,N_9149,N_8448);
nor U13261 (N_13261,N_8668,N_11105);
xnor U13262 (N_13262,N_9562,N_10010);
nand U13263 (N_13263,N_10992,N_11894);
and U13264 (N_13264,N_8768,N_9198);
nand U13265 (N_13265,N_11879,N_11596);
xnor U13266 (N_13266,N_11839,N_11786);
xnor U13267 (N_13267,N_10996,N_10364);
nand U13268 (N_13268,N_10949,N_11618);
nor U13269 (N_13269,N_8021,N_9389);
xnor U13270 (N_13270,N_11979,N_10002);
or U13271 (N_13271,N_11080,N_9615);
or U13272 (N_13272,N_11458,N_11584);
xnor U13273 (N_13273,N_10345,N_11424);
or U13274 (N_13274,N_8211,N_8264);
or U13275 (N_13275,N_8189,N_11104);
and U13276 (N_13276,N_11620,N_11685);
and U13277 (N_13277,N_10165,N_8270);
and U13278 (N_13278,N_9520,N_10817);
nor U13279 (N_13279,N_9733,N_10120);
or U13280 (N_13280,N_11897,N_9209);
or U13281 (N_13281,N_10709,N_11715);
nor U13282 (N_13282,N_9122,N_9319);
or U13283 (N_13283,N_8452,N_11535);
or U13284 (N_13284,N_8631,N_11159);
or U13285 (N_13285,N_10121,N_8196);
nand U13286 (N_13286,N_11356,N_10896);
nand U13287 (N_13287,N_9986,N_10745);
nor U13288 (N_13288,N_11140,N_9970);
nor U13289 (N_13289,N_8613,N_9465);
xor U13290 (N_13290,N_9892,N_8617);
nand U13291 (N_13291,N_10348,N_9039);
nand U13292 (N_13292,N_11383,N_11350);
nor U13293 (N_13293,N_9805,N_8075);
nand U13294 (N_13294,N_9554,N_11768);
xnor U13295 (N_13295,N_11176,N_11592);
or U13296 (N_13296,N_11426,N_9336);
and U13297 (N_13297,N_9447,N_8362);
xnor U13298 (N_13298,N_8451,N_10872);
and U13299 (N_13299,N_9799,N_10895);
nand U13300 (N_13300,N_8581,N_9370);
and U13301 (N_13301,N_10733,N_9488);
and U13302 (N_13302,N_8926,N_10730);
nand U13303 (N_13303,N_10265,N_8003);
xnor U13304 (N_13304,N_11757,N_8127);
nor U13305 (N_13305,N_8949,N_11372);
and U13306 (N_13306,N_8240,N_10901);
or U13307 (N_13307,N_11895,N_8959);
xnor U13308 (N_13308,N_10860,N_9933);
nor U13309 (N_13309,N_9426,N_8080);
nand U13310 (N_13310,N_11437,N_8472);
or U13311 (N_13311,N_9815,N_10371);
and U13312 (N_13312,N_9602,N_8992);
nand U13313 (N_13313,N_9672,N_10661);
and U13314 (N_13314,N_8981,N_10360);
nand U13315 (N_13315,N_8311,N_8690);
and U13316 (N_13316,N_11565,N_11382);
nor U13317 (N_13317,N_9195,N_8460);
nand U13318 (N_13318,N_10768,N_9075);
and U13319 (N_13319,N_9346,N_10747);
or U13320 (N_13320,N_8004,N_11387);
and U13321 (N_13321,N_8401,N_9855);
nor U13322 (N_13322,N_10584,N_8147);
nand U13323 (N_13323,N_9681,N_9373);
and U13324 (N_13324,N_8014,N_10553);
nand U13325 (N_13325,N_11326,N_8249);
nand U13326 (N_13326,N_9873,N_9908);
nor U13327 (N_13327,N_8428,N_9222);
nor U13328 (N_13328,N_8200,N_9929);
nor U13329 (N_13329,N_9879,N_10760);
xnor U13330 (N_13330,N_8279,N_11985);
nand U13331 (N_13331,N_11654,N_10542);
or U13332 (N_13332,N_8133,N_11121);
or U13333 (N_13333,N_8780,N_10564);
or U13334 (N_13334,N_10080,N_10007);
or U13335 (N_13335,N_10054,N_11634);
xor U13336 (N_13336,N_10145,N_9890);
nand U13337 (N_13337,N_8268,N_8538);
or U13338 (N_13338,N_10136,N_9090);
and U13339 (N_13339,N_10349,N_10190);
and U13340 (N_13340,N_11587,N_9569);
nor U13341 (N_13341,N_9578,N_9099);
nor U13342 (N_13342,N_8819,N_9285);
and U13343 (N_13343,N_10532,N_9739);
or U13344 (N_13344,N_9691,N_8505);
xor U13345 (N_13345,N_9750,N_10603);
nand U13346 (N_13346,N_9918,N_9793);
and U13347 (N_13347,N_11657,N_8455);
nand U13348 (N_13348,N_10903,N_8962);
and U13349 (N_13349,N_11668,N_9376);
nand U13350 (N_13350,N_10117,N_8539);
nor U13351 (N_13351,N_9682,N_8936);
nor U13352 (N_13352,N_9140,N_9539);
or U13353 (N_13353,N_10226,N_11371);
xnor U13354 (N_13354,N_8088,N_8206);
or U13355 (N_13355,N_11731,N_9518);
nor U13356 (N_13356,N_11143,N_8111);
xor U13357 (N_13357,N_11270,N_11243);
nor U13358 (N_13358,N_9300,N_10592);
nor U13359 (N_13359,N_8109,N_8106);
xor U13360 (N_13360,N_10224,N_11126);
xor U13361 (N_13361,N_11444,N_8980);
or U13362 (N_13362,N_9889,N_8231);
or U13363 (N_13363,N_11870,N_10748);
and U13364 (N_13364,N_10459,N_11473);
nor U13365 (N_13365,N_10581,N_10916);
nor U13366 (N_13366,N_8632,N_9192);
and U13367 (N_13367,N_9633,N_8709);
nand U13368 (N_13368,N_9718,N_9046);
and U13369 (N_13369,N_11550,N_9043);
xor U13370 (N_13370,N_8781,N_10255);
xor U13371 (N_13371,N_9162,N_11405);
nand U13372 (N_13372,N_11060,N_11517);
nor U13373 (N_13373,N_9489,N_9393);
nor U13374 (N_13374,N_9736,N_9326);
and U13375 (N_13375,N_9494,N_10636);
and U13376 (N_13376,N_10605,N_9707);
nand U13377 (N_13377,N_10354,N_8870);
or U13378 (N_13378,N_11236,N_11953);
and U13379 (N_13379,N_8839,N_10599);
xor U13380 (N_13380,N_11601,N_9213);
xor U13381 (N_13381,N_11427,N_10888);
nor U13382 (N_13382,N_10052,N_9620);
or U13383 (N_13383,N_10849,N_11283);
xor U13384 (N_13384,N_9829,N_11818);
nand U13385 (N_13385,N_9174,N_9235);
and U13386 (N_13386,N_9020,N_8251);
nor U13387 (N_13387,N_9687,N_10173);
xor U13388 (N_13388,N_9527,N_9848);
nand U13389 (N_13389,N_11900,N_9983);
nor U13390 (N_13390,N_8159,N_8650);
nand U13391 (N_13391,N_11773,N_8985);
nor U13392 (N_13392,N_10153,N_9586);
nand U13393 (N_13393,N_9660,N_9371);
nand U13394 (N_13394,N_11092,N_8141);
and U13395 (N_13395,N_11641,N_8201);
nor U13396 (N_13396,N_8181,N_8374);
or U13397 (N_13397,N_10689,N_8578);
xnor U13398 (N_13398,N_9065,N_10179);
or U13399 (N_13399,N_8686,N_9510);
xor U13400 (N_13400,N_11063,N_11150);
nor U13401 (N_13401,N_8309,N_11536);
xor U13402 (N_13402,N_11810,N_11229);
nor U13403 (N_13403,N_11557,N_8398);
and U13404 (N_13404,N_9422,N_9242);
xnor U13405 (N_13405,N_9940,N_9127);
and U13406 (N_13406,N_10141,N_8732);
nor U13407 (N_13407,N_10549,N_11563);
or U13408 (N_13408,N_8128,N_11970);
xnor U13409 (N_13409,N_8094,N_8680);
nand U13410 (N_13410,N_10893,N_10368);
nor U13411 (N_13411,N_11729,N_11683);
nor U13412 (N_13412,N_10514,N_8826);
and U13413 (N_13413,N_9141,N_11242);
or U13414 (N_13414,N_8246,N_9513);
xnor U13415 (N_13415,N_8997,N_10490);
nand U13416 (N_13416,N_11920,N_11694);
nor U13417 (N_13417,N_11721,N_8887);
nand U13418 (N_13418,N_8621,N_9036);
and U13419 (N_13419,N_10446,N_10293);
xnor U13420 (N_13420,N_11543,N_8923);
xor U13421 (N_13421,N_9107,N_8861);
xnor U13422 (N_13422,N_9811,N_11161);
and U13423 (N_13423,N_8432,N_10411);
nor U13424 (N_13424,N_10066,N_10261);
and U13425 (N_13425,N_9588,N_11921);
nand U13426 (N_13426,N_10798,N_11111);
nand U13427 (N_13427,N_8836,N_10041);
nor U13428 (N_13428,N_11820,N_8083);
xnor U13429 (N_13429,N_11361,N_9584);
or U13430 (N_13430,N_11840,N_10611);
nand U13431 (N_13431,N_11264,N_9187);
xor U13432 (N_13432,N_10347,N_9546);
and U13433 (N_13433,N_10501,N_10168);
or U13434 (N_13434,N_8029,N_9824);
or U13435 (N_13435,N_10579,N_10185);
or U13436 (N_13436,N_11411,N_9139);
and U13437 (N_13437,N_11219,N_11274);
nand U13438 (N_13438,N_11450,N_11302);
xnor U13439 (N_13439,N_11393,N_11942);
nor U13440 (N_13440,N_8089,N_8968);
xor U13441 (N_13441,N_10423,N_9227);
nand U13442 (N_13442,N_8987,N_11741);
nand U13443 (N_13443,N_10574,N_10424);
and U13444 (N_13444,N_9802,N_8493);
xor U13445 (N_13445,N_9674,N_9712);
and U13446 (N_13446,N_10476,N_9126);
nand U13447 (N_13447,N_10587,N_10528);
nand U13448 (N_13448,N_8634,N_10785);
nand U13449 (N_13449,N_9292,N_10116);
xor U13450 (N_13450,N_10946,N_10176);
or U13451 (N_13451,N_11431,N_9868);
xnor U13452 (N_13452,N_8227,N_11043);
or U13453 (N_13453,N_11521,N_10030);
or U13454 (N_13454,N_11044,N_8532);
and U13455 (N_13455,N_10192,N_11386);
xor U13456 (N_13456,N_11389,N_9571);
or U13457 (N_13457,N_8331,N_8252);
or U13458 (N_13458,N_10922,N_10038);
nor U13459 (N_13459,N_9934,N_10037);
xnor U13460 (N_13460,N_10258,N_9335);
and U13461 (N_13461,N_8888,N_10658);
nand U13462 (N_13462,N_9634,N_8153);
xnor U13463 (N_13463,N_8025,N_8600);
nand U13464 (N_13464,N_9392,N_10865);
xor U13465 (N_13465,N_11991,N_11318);
and U13466 (N_13466,N_11107,N_11093);
nand U13467 (N_13467,N_9159,N_8687);
nand U13468 (N_13468,N_11353,N_9069);
xnor U13469 (N_13469,N_9762,N_9720);
or U13470 (N_13470,N_10384,N_11808);
and U13471 (N_13471,N_9089,N_10051);
nor U13472 (N_13472,N_10913,N_11149);
xor U13473 (N_13473,N_8570,N_10492);
and U13474 (N_13474,N_9818,N_9684);
xnor U13475 (N_13475,N_10618,N_8256);
nor U13476 (N_13476,N_9502,N_8900);
nor U13477 (N_13477,N_11352,N_8302);
nor U13478 (N_13478,N_8288,N_10628);
or U13479 (N_13479,N_9841,N_10679);
xnor U13480 (N_13480,N_8020,N_10840);
or U13481 (N_13481,N_8736,N_11165);
nor U13482 (N_13482,N_10890,N_9186);
nand U13483 (N_13483,N_11564,N_8950);
nand U13484 (N_13484,N_8607,N_8978);
and U13485 (N_13485,N_11502,N_11691);
nor U13486 (N_13486,N_11414,N_9138);
nand U13487 (N_13487,N_9025,N_8659);
nor U13488 (N_13488,N_10936,N_9478);
or U13489 (N_13489,N_8627,N_9151);
or U13490 (N_13490,N_10440,N_8412);
nand U13491 (N_13491,N_8798,N_9382);
nand U13492 (N_13492,N_10487,N_8015);
and U13493 (N_13493,N_10373,N_8907);
nor U13494 (N_13494,N_11252,N_8100);
nand U13495 (N_13495,N_11519,N_9275);
xnor U13496 (N_13496,N_10478,N_8637);
or U13497 (N_13497,N_8546,N_10700);
or U13498 (N_13498,N_9103,N_8269);
xnor U13499 (N_13499,N_8146,N_9515);
and U13500 (N_13500,N_9572,N_10650);
or U13501 (N_13501,N_10678,N_11562);
nand U13502 (N_13502,N_9888,N_9358);
or U13503 (N_13503,N_9265,N_8995);
and U13504 (N_13504,N_11548,N_11692);
nand U13505 (N_13505,N_8847,N_10940);
or U13506 (N_13506,N_10489,N_10231);
and U13507 (N_13507,N_9953,N_10441);
or U13508 (N_13508,N_11845,N_9826);
nand U13509 (N_13509,N_10181,N_8492);
or U13510 (N_13510,N_11711,N_8640);
or U13511 (N_13511,N_10696,N_10203);
and U13512 (N_13512,N_9350,N_8390);
and U13513 (N_13513,N_9955,N_8464);
xor U13514 (N_13514,N_8208,N_8639);
xnor U13515 (N_13515,N_8226,N_10988);
nor U13516 (N_13516,N_8488,N_10960);
or U13517 (N_13517,N_9436,N_11830);
or U13518 (N_13518,N_11133,N_9785);
nand U13519 (N_13519,N_11073,N_11951);
and U13520 (N_13520,N_11873,N_10624);
and U13521 (N_13521,N_11128,N_11203);
nand U13522 (N_13522,N_11581,N_10216);
nor U13523 (N_13523,N_8547,N_8334);
nand U13524 (N_13524,N_10481,N_10223);
nand U13525 (N_13525,N_10945,N_11136);
or U13526 (N_13526,N_8919,N_10302);
nor U13527 (N_13527,N_9220,N_11299);
and U13528 (N_13528,N_8947,N_10219);
and U13529 (N_13529,N_10004,N_10303);
xnor U13530 (N_13530,N_11276,N_9521);
nor U13531 (N_13531,N_9638,N_11084);
xnor U13532 (N_13532,N_11858,N_11836);
and U13533 (N_13533,N_8724,N_8481);
nand U13534 (N_13534,N_9255,N_9921);
nand U13535 (N_13535,N_11271,N_9533);
nor U13536 (N_13536,N_11155,N_10312);
and U13537 (N_13537,N_9686,N_9514);
nand U13538 (N_13538,N_9157,N_10482);
nand U13539 (N_13539,N_10756,N_11320);
nor U13540 (N_13540,N_8333,N_8575);
nor U13541 (N_13541,N_10277,N_10104);
nor U13542 (N_13542,N_8771,N_11238);
or U13543 (N_13543,N_11195,N_11947);
and U13544 (N_13544,N_11864,N_10089);
xnor U13545 (N_13545,N_9474,N_10294);
nor U13546 (N_13546,N_10102,N_11479);
xnor U13547 (N_13547,N_8664,N_10395);
xnor U13548 (N_13548,N_10687,N_9598);
nand U13549 (N_13549,N_10753,N_11974);
nand U13550 (N_13550,N_8810,N_11995);
nor U13551 (N_13551,N_10694,N_10412);
and U13552 (N_13552,N_10287,N_9029);
nor U13553 (N_13553,N_11853,N_10663);
xnor U13554 (N_13554,N_9425,N_9905);
nor U13555 (N_13555,N_10127,N_11118);
nor U13556 (N_13556,N_11675,N_11863);
or U13557 (N_13557,N_11224,N_10824);
nor U13558 (N_13558,N_9922,N_11232);
nand U13559 (N_13559,N_10688,N_10436);
nand U13560 (N_13560,N_9603,N_9041);
or U13561 (N_13561,N_10670,N_10620);
and U13562 (N_13562,N_11760,N_11045);
and U13563 (N_13563,N_10276,N_10367);
and U13564 (N_13564,N_8057,N_8898);
or U13565 (N_13565,N_11470,N_10256);
and U13566 (N_13566,N_8644,N_11421);
nor U13567 (N_13567,N_10456,N_8385);
and U13568 (N_13568,N_8824,N_9716);
and U13569 (N_13569,N_10400,N_8314);
nand U13570 (N_13570,N_11321,N_8292);
nand U13571 (N_13571,N_9434,N_11464);
xnor U13572 (N_13572,N_9271,N_11139);
and U13573 (N_13573,N_11019,N_9504);
xnor U13574 (N_13574,N_8043,N_9011);
xnor U13575 (N_13575,N_8649,N_11936);
or U13576 (N_13576,N_10204,N_11586);
or U13577 (N_13577,N_9230,N_8873);
nand U13578 (N_13578,N_8871,N_9351);
and U13579 (N_13579,N_8322,N_11069);
nand U13580 (N_13580,N_11085,N_11664);
and U13581 (N_13581,N_10621,N_11122);
or U13582 (N_13582,N_10003,N_9561);
nor U13583 (N_13583,N_11441,N_11407);
nand U13584 (N_13584,N_10109,N_11631);
or U13585 (N_13585,N_10994,N_11687);
nor U13586 (N_13586,N_10879,N_9348);
xor U13587 (N_13587,N_8576,N_8265);
nand U13588 (N_13588,N_9722,N_10288);
xor U13589 (N_13589,N_8865,N_8371);
nand U13590 (N_13590,N_8018,N_11453);
xor U13591 (N_13591,N_8404,N_8473);
xor U13592 (N_13592,N_8411,N_9440);
xor U13593 (N_13593,N_8517,N_11725);
and U13594 (N_13594,N_8134,N_10160);
nor U13595 (N_13595,N_11677,N_9385);
and U13596 (N_13596,N_10794,N_8204);
xor U13597 (N_13597,N_9771,N_11148);
nand U13598 (N_13598,N_10471,N_8341);
and U13599 (N_13599,N_11035,N_8572);
xnor U13600 (N_13600,N_10971,N_8316);
or U13601 (N_13601,N_10419,N_11130);
and U13602 (N_13602,N_11434,N_10877);
or U13603 (N_13603,N_8795,N_11448);
nor U13604 (N_13604,N_10586,N_8166);
nand U13605 (N_13605,N_9834,N_9387);
nor U13606 (N_13606,N_11188,N_10421);
xor U13607 (N_13607,N_9991,N_11834);
nor U13608 (N_13608,N_10026,N_11952);
nand U13609 (N_13609,N_10324,N_9662);
nor U13610 (N_13610,N_11369,N_11607);
nor U13611 (N_13611,N_11789,N_8254);
or U13612 (N_13612,N_8363,N_10433);
xor U13613 (N_13613,N_8902,N_9639);
xor U13614 (N_13614,N_9224,N_9976);
or U13615 (N_13615,N_8248,N_10230);
or U13616 (N_13616,N_11595,N_11688);
and U13617 (N_13617,N_10545,N_10982);
nor U13618 (N_13618,N_9049,N_11269);
nand U13619 (N_13619,N_10729,N_10260);
nor U13620 (N_13620,N_8660,N_9378);
nor U13621 (N_13621,N_8093,N_8132);
nand U13622 (N_13622,N_11795,N_8714);
nor U13623 (N_13623,N_8841,N_10771);
xor U13624 (N_13624,N_8364,N_10188);
nor U13625 (N_13625,N_10716,N_8920);
and U13626 (N_13626,N_8914,N_11803);
and U13627 (N_13627,N_9693,N_8409);
and U13628 (N_13628,N_11826,N_9399);
nand U13629 (N_13629,N_10315,N_10259);
xnor U13630 (N_13630,N_9095,N_8096);
nor U13631 (N_13631,N_11739,N_11799);
xor U13632 (N_13632,N_9666,N_9009);
or U13633 (N_13633,N_11249,N_8137);
xnor U13634 (N_13634,N_8152,N_9406);
and U13635 (N_13635,N_11081,N_9431);
or U13636 (N_13636,N_11115,N_8289);
and U13637 (N_13637,N_10254,N_8443);
nand U13638 (N_13638,N_8703,N_11391);
and U13639 (N_13639,N_10602,N_11551);
and U13640 (N_13640,N_8348,N_10808);
or U13641 (N_13641,N_10854,N_11782);
nand U13642 (N_13642,N_11764,N_8170);
and U13643 (N_13643,N_10836,N_8662);
nor U13644 (N_13644,N_10393,N_11206);
or U13645 (N_13645,N_8480,N_11438);
and U13646 (N_13646,N_11443,N_8673);
or U13647 (N_13647,N_9176,N_11525);
nor U13648 (N_13648,N_9450,N_8485);
and U13649 (N_13649,N_9989,N_9781);
xnor U13650 (N_13650,N_8154,N_11670);
or U13651 (N_13651,N_11887,N_10451);
and U13652 (N_13652,N_10351,N_10924);
xnor U13653 (N_13653,N_11571,N_8119);
xor U13654 (N_13654,N_11671,N_11924);
or U13655 (N_13655,N_10452,N_10319);
and U13656 (N_13656,N_9119,N_9333);
and U13657 (N_13657,N_11769,N_10511);
xor U13658 (N_13658,N_8444,N_10325);
or U13659 (N_13659,N_10131,N_9911);
and U13660 (N_13660,N_10063,N_9196);
nand U13661 (N_13661,N_8143,N_11037);
nor U13662 (N_13662,N_8070,N_11889);
xor U13663 (N_13663,N_10681,N_10813);
nand U13664 (N_13664,N_10786,N_10407);
xnor U13665 (N_13665,N_9259,N_9746);
or U13666 (N_13666,N_9492,N_9418);
nand U13667 (N_13667,N_10220,N_11511);
nor U13668 (N_13668,N_8330,N_11609);
or U13669 (N_13669,N_11158,N_11510);
nand U13670 (N_13670,N_8944,N_10034);
nor U13671 (N_13671,N_8951,N_11327);
nand U13672 (N_13672,N_9668,N_8956);
xnor U13673 (N_13673,N_8384,N_11850);
or U13674 (N_13674,N_11857,N_11324);
or U13675 (N_13675,N_8922,N_8843);
nor U13676 (N_13676,N_11977,N_8391);
and U13677 (N_13677,N_10247,N_10933);
nand U13678 (N_13678,N_11712,N_8675);
nand U13679 (N_13679,N_8594,N_8469);
nand U13680 (N_13680,N_10741,N_10062);
nor U13681 (N_13681,N_11141,N_8893);
xor U13682 (N_13682,N_8016,N_11926);
and U13683 (N_13683,N_11624,N_8846);
nand U13684 (N_13684,N_10780,N_8437);
and U13685 (N_13685,N_9206,N_10458);
nor U13686 (N_13686,N_10573,N_9964);
nand U13687 (N_13687,N_10425,N_9997);
and U13688 (N_13688,N_11915,N_9895);
xor U13689 (N_13689,N_8190,N_8894);
nand U13690 (N_13690,N_11771,N_10643);
nand U13691 (N_13691,N_10206,N_10541);
xor U13692 (N_13692,N_8764,N_8144);
xnor U13693 (N_13693,N_8463,N_11342);
xor U13694 (N_13694,N_8151,N_9121);
xnor U13695 (N_13695,N_10248,N_10467);
or U13696 (N_13696,N_8583,N_9902);
xnor U13697 (N_13697,N_8554,N_10985);
and U13698 (N_13698,N_10797,N_9759);
xor U13699 (N_13699,N_10498,N_8071);
xnor U13700 (N_13700,N_10283,N_8747);
nand U13701 (N_13701,N_10449,N_8476);
nand U13702 (N_13702,N_9971,N_8059);
nor U13703 (N_13703,N_10151,N_8332);
nand U13704 (N_13704,N_11365,N_11911);
and U13705 (N_13705,N_11027,N_9601);
xnor U13706 (N_13706,N_11807,N_8852);
nand U13707 (N_13707,N_9798,N_9702);
nor U13708 (N_13708,N_10589,N_9147);
and U13709 (N_13709,N_9857,N_8097);
and U13710 (N_13710,N_9648,N_11000);
nand U13711 (N_13711,N_8199,N_8163);
and U13712 (N_13712,N_11572,N_11221);
nand U13713 (N_13713,N_10925,N_10383);
nor U13714 (N_13714,N_9524,N_11559);
nor U13715 (N_13715,N_10543,N_10381);
or U13716 (N_13716,N_11663,N_11068);
and U13717 (N_13717,N_8007,N_11616);
nor U13718 (N_13718,N_9606,N_11017);
xor U13719 (N_13719,N_10005,N_11958);
and U13720 (N_13720,N_11591,N_9708);
nand U13721 (N_13721,N_8884,N_9698);
and U13722 (N_13722,N_8008,N_9038);
or U13723 (N_13723,N_11848,N_10356);
or U13724 (N_13724,N_9028,N_10443);
nand U13725 (N_13725,N_8854,N_11492);
xor U13726 (N_13726,N_10343,N_9825);
nor U13727 (N_13727,N_9237,N_10941);
nor U13728 (N_13728,N_10781,N_10146);
or U13729 (N_13729,N_11399,N_10284);
and U13730 (N_13730,N_10723,N_11678);
xnor U13731 (N_13731,N_10426,N_9575);
nand U13732 (N_13732,N_9767,N_9963);
and U13733 (N_13733,N_9568,N_11829);
xor U13734 (N_13734,N_11157,N_9650);
or U13735 (N_13735,N_11279,N_9340);
nor U13736 (N_13736,N_9462,N_10152);
or U13737 (N_13737,N_8383,N_8590);
nor U13738 (N_13738,N_8999,N_10292);
xnor U13739 (N_13739,N_10710,N_10823);
nand U13740 (N_13740,N_9106,N_11504);
or U13741 (N_13741,N_9577,N_11201);
or U13742 (N_13742,N_8382,N_8416);
nor U13743 (N_13743,N_9177,N_9665);
nand U13744 (N_13744,N_11885,N_8420);
nand U13745 (N_13745,N_10669,N_9354);
or U13746 (N_13746,N_11096,N_9243);
nand U13747 (N_13747,N_9565,N_8734);
xor U13748 (N_13748,N_11943,N_10094);
and U13749 (N_13749,N_11978,N_9493);
and U13750 (N_13750,N_8779,N_9849);
nor U13751 (N_13751,N_10920,N_8766);
and U13752 (N_13752,N_11210,N_9287);
xnor U13753 (N_13753,N_8913,N_11569);
nor U13754 (N_13754,N_10853,N_8466);
nand U13755 (N_13755,N_10027,N_10234);
nand U13756 (N_13756,N_11245,N_11058);
and U13757 (N_13757,N_9535,N_8827);
or U13758 (N_13758,N_9108,N_9727);
nor U13759 (N_13759,N_10972,N_8508);
or U13760 (N_13760,N_9627,N_10358);
xnor U13761 (N_13761,N_10770,N_8676);
nand U13762 (N_13762,N_9948,N_9226);
and U13763 (N_13763,N_11582,N_9064);
and U13764 (N_13764,N_11256,N_8354);
nand U13765 (N_13765,N_9364,N_8442);
and U13766 (N_13766,N_10938,N_8516);
xor U13767 (N_13767,N_9194,N_8454);
nor U13768 (N_13768,N_9804,N_10882);
nor U13769 (N_13769,N_9405,N_9010);
nor U13770 (N_13770,N_8087,N_11482);
or U13771 (N_13771,N_8528,N_9732);
xor U13772 (N_13772,N_9507,N_9101);
xnor U13773 (N_13773,N_11690,N_8715);
nor U13774 (N_13774,N_11373,N_11585);
or U13775 (N_13775,N_9397,N_9172);
nand U13776 (N_13776,N_11304,N_8838);
nand U13777 (N_13777,N_10923,N_10655);
or U13778 (N_13778,N_11199,N_11633);
and U13779 (N_13779,N_11132,N_9531);
nor U13780 (N_13780,N_10531,N_10214);
nor U13781 (N_13781,N_11761,N_10948);
nand U13782 (N_13782,N_10326,N_9414);
nand U13783 (N_13783,N_8749,N_10012);
or U13784 (N_13784,N_8280,N_9499);
and U13785 (N_13785,N_10961,N_8185);
nand U13786 (N_13786,N_9120,N_9993);
nand U13787 (N_13787,N_10290,N_8596);
xnor U13788 (N_13788,N_10793,N_11946);
or U13789 (N_13789,N_11679,N_10076);
and U13790 (N_13790,N_8323,N_8857);
and U13791 (N_13791,N_9523,N_11293);
nand U13792 (N_13792,N_9850,N_11568);
nor U13793 (N_13793,N_9794,N_8953);
nand U13794 (N_13794,N_10392,N_8145);
or U13795 (N_13795,N_8278,N_11131);
nor U13796 (N_13796,N_11260,N_11413);
and U13797 (N_13797,N_8961,N_8005);
and U13798 (N_13798,N_10891,N_11334);
or U13799 (N_13799,N_8250,N_8047);
nand U13800 (N_13800,N_11075,N_10957);
xor U13801 (N_13801,N_8800,N_11380);
or U13802 (N_13802,N_9636,N_9968);
nand U13803 (N_13803,N_9250,N_9473);
nor U13804 (N_13804,N_8801,N_11866);
nor U13805 (N_13805,N_8645,N_9055);
or U13806 (N_13806,N_11909,N_9212);
nor U13807 (N_13807,N_9077,N_10792);
xor U13808 (N_13808,N_9600,N_8821);
and U13809 (N_13809,N_9925,N_11226);
xor U13810 (N_13810,N_9076,N_10427);
and U13811 (N_13811,N_11661,N_11622);
and U13812 (N_13812,N_8638,N_9998);
xnor U13813 (N_13813,N_9322,N_8683);
nor U13814 (N_13814,N_10928,N_10612);
or U13815 (N_13815,N_8835,N_9105);
and U13816 (N_13816,N_10275,N_9773);
nor U13817 (N_13817,N_8598,N_11781);
or U13818 (N_13818,N_8814,N_8076);
and U13819 (N_13819,N_9403,N_11054);
xor U13820 (N_13820,N_9104,N_8697);
nor U13821 (N_13821,N_10715,N_9469);
or U13822 (N_13822,N_9820,N_10167);
and U13823 (N_13823,N_9325,N_9114);
xnor U13824 (N_13824,N_8647,N_10221);
or U13825 (N_13825,N_9994,N_10683);
and U13826 (N_13826,N_11408,N_9704);
nand U13827 (N_13827,N_8582,N_9809);
or U13828 (N_13828,N_8450,N_11197);
nand U13829 (N_13829,N_9391,N_11066);
nor U13830 (N_13830,N_11531,N_11466);
xor U13831 (N_13831,N_8790,N_10858);
or U13832 (N_13832,N_8972,N_11442);
nand U13833 (N_13833,N_8191,N_8381);
and U13834 (N_13834,N_8421,N_8275);
nor U13835 (N_13835,N_9581,N_9635);
or U13836 (N_13836,N_8760,N_8305);
nor U13837 (N_13837,N_9800,N_10555);
xor U13838 (N_13838,N_11514,N_11791);
or U13839 (N_13839,N_11331,N_9200);
xor U13840 (N_13840,N_10702,N_10201);
xnor U13841 (N_13841,N_10163,N_10390);
or U13842 (N_13842,N_8419,N_10212);
or U13843 (N_13843,N_11992,N_10736);
nand U13844 (N_13844,N_9293,N_8665);
xor U13845 (N_13845,N_10978,N_11701);
xor U13846 (N_13846,N_8160,N_11418);
xnor U13847 (N_13847,N_8427,N_8236);
xor U13848 (N_13848,N_10539,N_10850);
nand U13849 (N_13849,N_11172,N_8329);
or U13850 (N_13850,N_10475,N_10719);
or U13851 (N_13851,N_11792,N_10726);
xor U13852 (N_13852,N_11110,N_9549);
and U13853 (N_13853,N_8359,N_10962);
or U13854 (N_13854,N_11982,N_9254);
nor U13855 (N_13855,N_10987,N_10341);
and U13856 (N_13856,N_9257,N_8567);
or U13857 (N_13857,N_11503,N_9943);
and U13858 (N_13858,N_9453,N_8941);
nand U13859 (N_13859,N_11465,N_9045);
xor U13860 (N_13860,N_9893,N_11774);
and U13861 (N_13861,N_11200,N_10387);
xor U13862 (N_13862,N_9966,N_9812);
xor U13863 (N_13863,N_8842,N_9658);
nor U13864 (N_13864,N_9204,N_11336);
nand U13865 (N_13865,N_9623,N_11368);
xnor U13866 (N_13866,N_10759,N_9158);
nand U13867 (N_13867,N_8718,N_8113);
nand U13868 (N_13868,N_8298,N_10593);
or U13869 (N_13869,N_8577,N_9528);
or U13870 (N_13870,N_10280,N_8762);
and U13871 (N_13871,N_11865,N_10881);
xnor U13872 (N_13872,N_11495,N_11680);
nor U13873 (N_13873,N_9560,N_9153);
nand U13874 (N_13874,N_9878,N_9846);
nor U13875 (N_13875,N_8349,N_11912);
and U13876 (N_13876,N_9267,N_11266);
or U13877 (N_13877,N_9066,N_11509);
nor U13878 (N_13878,N_11345,N_11472);
and U13879 (N_13879,N_8140,N_8751);
nor U13880 (N_13880,N_9663,N_8276);
xnor U13881 (N_13881,N_8693,N_10069);
nand U13882 (N_13882,N_9570,N_8342);
nand U13883 (N_13883,N_10830,N_9840);
and U13884 (N_13884,N_11522,N_8782);
nand U13885 (N_13885,N_8977,N_10111);
nor U13886 (N_13886,N_10750,N_10147);
nand U13887 (N_13887,N_8774,N_8670);
or U13888 (N_13888,N_8755,N_10285);
nor U13889 (N_13889,N_10908,N_10777);
or U13890 (N_13890,N_10042,N_9309);
or U13891 (N_13891,N_10576,N_9129);
nor U13892 (N_13892,N_11074,N_10567);
and U13893 (N_13893,N_9564,N_11009);
xor U13894 (N_13894,N_9590,N_9942);
nor U13895 (N_13895,N_11660,N_11267);
nand U13896 (N_13896,N_11142,N_11406);
and U13897 (N_13897,N_9582,N_9229);
nand U13898 (N_13898,N_10184,N_8192);
and U13899 (N_13899,N_9013,N_10652);
nand U13900 (N_13900,N_11528,N_10990);
xnor U13901 (N_13901,N_11727,N_8635);
xnor U13902 (N_13902,N_10956,N_8010);
or U13903 (N_13903,N_10701,N_11639);
and U13904 (N_13904,N_9167,N_8844);
and U13905 (N_13905,N_8901,N_8216);
and U13906 (N_13906,N_8597,N_8271);
and U13907 (N_13907,N_10020,N_10977);
xnor U13908 (N_13908,N_8477,N_8284);
or U13909 (N_13909,N_9320,N_9928);
or U13910 (N_13910,N_8545,N_8306);
nor U13911 (N_13911,N_11432,N_10148);
nand U13912 (N_13912,N_8414,N_8908);
nand U13913 (N_13913,N_8593,N_9410);
xnor U13914 (N_13914,N_9832,N_10331);
nor U13915 (N_13915,N_8031,N_10704);
and U13916 (N_13916,N_11984,N_8261);
nand U13917 (N_13917,N_11059,N_11208);
or U13918 (N_13918,N_10885,N_10480);
xor U13919 (N_13919,N_11253,N_9827);
nand U13920 (N_13920,N_10739,N_9753);
nor U13921 (N_13921,N_9190,N_9801);
nor U13922 (N_13922,N_8850,N_11744);
xor U13923 (N_13923,N_10833,N_8303);
nor U13924 (N_13924,N_10328,N_11994);
xnor U13925 (N_13925,N_8998,N_10673);
xnor U13926 (N_13926,N_10238,N_10790);
nor U13927 (N_13927,N_10342,N_10629);
and U13928 (N_13928,N_9276,N_8672);
xor U13929 (N_13929,N_8891,N_9324);
xor U13930 (N_13930,N_8713,N_9914);
and U13931 (N_13931,N_9556,N_10225);
and U13932 (N_13932,N_9480,N_8415);
xnor U13933 (N_13933,N_11867,N_10796);
xnor U13934 (N_13934,N_11614,N_10705);
and U13935 (N_13935,N_11861,N_11859);
nor U13936 (N_13936,N_9685,N_8130);
and U13937 (N_13937,N_9252,N_8820);
xnor U13938 (N_13938,N_11956,N_11801);
nor U13939 (N_13939,N_9547,N_11477);
nor U13940 (N_13940,N_10494,N_10417);
nor U13941 (N_13941,N_9768,N_10361);
nor U13942 (N_13942,N_10869,N_8802);
and U13943 (N_13943,N_8078,N_8424);
and U13944 (N_13944,N_11749,N_8356);
nand U13945 (N_13945,N_8255,N_11573);
nand U13946 (N_13946,N_11187,N_8506);
nor U13947 (N_13947,N_10981,N_9093);
and U13948 (N_13948,N_8641,N_8930);
nand U13949 (N_13949,N_11669,N_8066);
and U13950 (N_13950,N_11125,N_8091);
and U13951 (N_13951,N_11662,N_9366);
or U13952 (N_13952,N_11237,N_11410);
nand U13953 (N_13953,N_11429,N_11213);
nor U13954 (N_13954,N_9676,N_9961);
and U13955 (N_13955,N_9273,N_9671);
xor U13956 (N_13956,N_10976,N_9210);
and U13957 (N_13957,N_8934,N_8942);
xor U13958 (N_13958,N_11733,N_11137);
nor U13959 (N_13959,N_10583,N_9052);
and U13960 (N_13960,N_11306,N_8916);
and U13961 (N_13961,N_11061,N_8282);
xnor U13962 (N_13962,N_10215,N_9788);
xor U13963 (N_13963,N_9689,N_9270);
and U13964 (N_13964,N_10330,N_9012);
xnor U13965 (N_13965,N_10016,N_8347);
nor U13966 (N_13966,N_8899,N_10954);
nand U13967 (N_13967,N_10483,N_10693);
nor U13968 (N_13968,N_8568,N_9766);
or U13969 (N_13969,N_10014,N_11628);
nand U13970 (N_13970,N_10935,N_10580);
and U13971 (N_13971,N_11297,N_10362);
or U13972 (N_13972,N_8219,N_11772);
xor U13973 (N_13973,N_10540,N_9795);
and U13974 (N_13974,N_9279,N_10090);
nor U13975 (N_13975,N_9016,N_11451);
nor U13976 (N_13976,N_8796,N_8438);
nor U13977 (N_13977,N_11029,N_10898);
or U13978 (N_13978,N_9563,N_10346);
xnor U13979 (N_13979,N_11593,N_10493);
nand U13980 (N_13980,N_8142,N_9062);
and U13981 (N_13981,N_10779,N_8866);
and U13982 (N_13982,N_11730,N_10752);
nor U13983 (N_13983,N_9880,N_11785);
xnor U13984 (N_13984,N_11034,N_8129);
nor U13985 (N_13985,N_10927,N_8459);
or U13986 (N_13986,N_9124,N_8685);
or U13987 (N_13987,N_9748,N_8906);
or U13988 (N_13988,N_10353,N_8792);
xor U13989 (N_13989,N_10169,N_8184);
nor U13990 (N_13990,N_8325,N_8055);
nand U13991 (N_13991,N_11577,N_9441);
or U13992 (N_13992,N_8183,N_11854);
nand U13993 (N_13993,N_10871,N_8522);
nor U13994 (N_13994,N_10560,N_10139);
and U13995 (N_13995,N_8825,N_9957);
nor U13996 (N_13996,N_9763,N_10875);
nand U13997 (N_13997,N_9587,N_11716);
or U13998 (N_13998,N_8832,N_11298);
and U13999 (N_13999,N_9323,N_11323);
or U14000 (N_14000,N_8872,N_9550);
xor U14001 (N_14001,N_10431,N_10220);
nand U14002 (N_14002,N_10925,N_11278);
or U14003 (N_14003,N_11785,N_8777);
nand U14004 (N_14004,N_8815,N_10847);
nor U14005 (N_14005,N_11596,N_10980);
and U14006 (N_14006,N_8701,N_10328);
or U14007 (N_14007,N_9473,N_10535);
and U14008 (N_14008,N_11754,N_8441);
or U14009 (N_14009,N_10480,N_9616);
nor U14010 (N_14010,N_10901,N_9569);
or U14011 (N_14011,N_9266,N_9922);
nor U14012 (N_14012,N_9974,N_8067);
and U14013 (N_14013,N_8033,N_11981);
nor U14014 (N_14014,N_11634,N_10831);
nor U14015 (N_14015,N_8691,N_10914);
and U14016 (N_14016,N_11152,N_11531);
nor U14017 (N_14017,N_8152,N_9511);
nor U14018 (N_14018,N_9987,N_10968);
xor U14019 (N_14019,N_8780,N_8680);
or U14020 (N_14020,N_11032,N_10974);
xnor U14021 (N_14021,N_9455,N_11784);
or U14022 (N_14022,N_8084,N_9128);
nor U14023 (N_14023,N_8946,N_11984);
and U14024 (N_14024,N_9216,N_10134);
and U14025 (N_14025,N_8649,N_11923);
nor U14026 (N_14026,N_11272,N_8968);
and U14027 (N_14027,N_9797,N_9134);
and U14028 (N_14028,N_11646,N_11186);
xnor U14029 (N_14029,N_8284,N_11274);
xor U14030 (N_14030,N_11119,N_9903);
nor U14031 (N_14031,N_10010,N_10937);
nand U14032 (N_14032,N_10588,N_11744);
nor U14033 (N_14033,N_10198,N_11127);
and U14034 (N_14034,N_9002,N_11797);
or U14035 (N_14035,N_10337,N_11712);
xnor U14036 (N_14036,N_10157,N_8195);
xor U14037 (N_14037,N_9115,N_10285);
nand U14038 (N_14038,N_9490,N_8952);
xor U14039 (N_14039,N_11166,N_8501);
xnor U14040 (N_14040,N_9635,N_9895);
and U14041 (N_14041,N_9416,N_10280);
nand U14042 (N_14042,N_8937,N_9684);
nor U14043 (N_14043,N_10852,N_10100);
nor U14044 (N_14044,N_11242,N_10415);
nand U14045 (N_14045,N_11616,N_9529);
nand U14046 (N_14046,N_8313,N_9081);
and U14047 (N_14047,N_8724,N_10353);
nor U14048 (N_14048,N_11001,N_9287);
nand U14049 (N_14049,N_8958,N_11877);
or U14050 (N_14050,N_10884,N_11031);
or U14051 (N_14051,N_11818,N_9458);
nor U14052 (N_14052,N_10784,N_9266);
nand U14053 (N_14053,N_9325,N_11512);
nor U14054 (N_14054,N_11466,N_9360);
and U14055 (N_14055,N_11069,N_11854);
or U14056 (N_14056,N_9932,N_10331);
nor U14057 (N_14057,N_10353,N_10332);
and U14058 (N_14058,N_10488,N_9462);
xnor U14059 (N_14059,N_10694,N_9535);
xor U14060 (N_14060,N_8616,N_11244);
and U14061 (N_14061,N_10006,N_10063);
xor U14062 (N_14062,N_10405,N_10446);
xnor U14063 (N_14063,N_10423,N_11617);
xor U14064 (N_14064,N_10022,N_9861);
nand U14065 (N_14065,N_9329,N_9817);
xnor U14066 (N_14066,N_8602,N_11756);
and U14067 (N_14067,N_8912,N_8371);
nand U14068 (N_14068,N_9001,N_11607);
or U14069 (N_14069,N_11059,N_9539);
or U14070 (N_14070,N_11276,N_9142);
xnor U14071 (N_14071,N_11188,N_11182);
nand U14072 (N_14072,N_8153,N_9552);
and U14073 (N_14073,N_8679,N_8546);
nand U14074 (N_14074,N_8801,N_11790);
and U14075 (N_14075,N_9099,N_10911);
and U14076 (N_14076,N_10582,N_8415);
or U14077 (N_14077,N_10373,N_9488);
and U14078 (N_14078,N_11938,N_8232);
xnor U14079 (N_14079,N_11036,N_8619);
nand U14080 (N_14080,N_8968,N_8291);
nand U14081 (N_14081,N_10900,N_11300);
nand U14082 (N_14082,N_9759,N_10338);
nand U14083 (N_14083,N_8830,N_11090);
and U14084 (N_14084,N_11765,N_11078);
or U14085 (N_14085,N_10859,N_9205);
xor U14086 (N_14086,N_8748,N_9303);
nor U14087 (N_14087,N_9883,N_10591);
xor U14088 (N_14088,N_10137,N_8949);
nor U14089 (N_14089,N_11066,N_9836);
nand U14090 (N_14090,N_11063,N_8824);
nand U14091 (N_14091,N_10031,N_8265);
nand U14092 (N_14092,N_10754,N_9358);
or U14093 (N_14093,N_8555,N_9082);
and U14094 (N_14094,N_10789,N_10739);
nor U14095 (N_14095,N_8430,N_10751);
nor U14096 (N_14096,N_8958,N_8292);
xnor U14097 (N_14097,N_9501,N_11547);
nor U14098 (N_14098,N_11352,N_11022);
nand U14099 (N_14099,N_11468,N_8324);
nand U14100 (N_14100,N_10376,N_9521);
nor U14101 (N_14101,N_8495,N_8163);
xor U14102 (N_14102,N_8953,N_10154);
nand U14103 (N_14103,N_10973,N_11481);
or U14104 (N_14104,N_10325,N_11705);
nand U14105 (N_14105,N_10928,N_8897);
xor U14106 (N_14106,N_9764,N_8842);
or U14107 (N_14107,N_10824,N_11738);
nand U14108 (N_14108,N_11293,N_11209);
xnor U14109 (N_14109,N_9520,N_11852);
nor U14110 (N_14110,N_9772,N_9842);
and U14111 (N_14111,N_10610,N_9094);
nor U14112 (N_14112,N_10423,N_8616);
xor U14113 (N_14113,N_11962,N_11134);
xor U14114 (N_14114,N_9896,N_11949);
nand U14115 (N_14115,N_9941,N_10318);
xnor U14116 (N_14116,N_8144,N_8208);
nand U14117 (N_14117,N_11915,N_10479);
nand U14118 (N_14118,N_10473,N_11805);
or U14119 (N_14119,N_8493,N_8919);
and U14120 (N_14120,N_9150,N_10740);
xor U14121 (N_14121,N_8063,N_11541);
xor U14122 (N_14122,N_11462,N_10130);
nand U14123 (N_14123,N_11123,N_9517);
nor U14124 (N_14124,N_9523,N_10607);
nor U14125 (N_14125,N_10358,N_9770);
nor U14126 (N_14126,N_9892,N_10767);
or U14127 (N_14127,N_11757,N_8400);
xor U14128 (N_14128,N_9785,N_8185);
nand U14129 (N_14129,N_8181,N_10791);
nand U14130 (N_14130,N_8054,N_9833);
nand U14131 (N_14131,N_8754,N_11923);
nor U14132 (N_14132,N_9893,N_11193);
or U14133 (N_14133,N_11212,N_11239);
nor U14134 (N_14134,N_9152,N_11113);
nor U14135 (N_14135,N_10813,N_11740);
and U14136 (N_14136,N_8623,N_9346);
nor U14137 (N_14137,N_10183,N_8196);
xnor U14138 (N_14138,N_9723,N_10719);
and U14139 (N_14139,N_11484,N_8002);
or U14140 (N_14140,N_8284,N_10980);
and U14141 (N_14141,N_11732,N_8079);
nand U14142 (N_14142,N_11247,N_11647);
nor U14143 (N_14143,N_11348,N_9267);
xor U14144 (N_14144,N_9382,N_9839);
nand U14145 (N_14145,N_10835,N_10394);
or U14146 (N_14146,N_11912,N_11840);
nor U14147 (N_14147,N_11105,N_11460);
and U14148 (N_14148,N_9156,N_9284);
and U14149 (N_14149,N_9926,N_10761);
nand U14150 (N_14150,N_11043,N_8387);
nor U14151 (N_14151,N_10311,N_9997);
or U14152 (N_14152,N_11621,N_8305);
nand U14153 (N_14153,N_9620,N_9324);
and U14154 (N_14154,N_9238,N_8280);
nand U14155 (N_14155,N_10984,N_8928);
and U14156 (N_14156,N_8703,N_9384);
or U14157 (N_14157,N_10501,N_9529);
nor U14158 (N_14158,N_11499,N_9436);
nand U14159 (N_14159,N_9156,N_11672);
nand U14160 (N_14160,N_8619,N_9422);
nand U14161 (N_14161,N_10442,N_9371);
xnor U14162 (N_14162,N_11570,N_9955);
and U14163 (N_14163,N_8119,N_8047);
nor U14164 (N_14164,N_8394,N_11973);
and U14165 (N_14165,N_10137,N_11768);
nand U14166 (N_14166,N_8784,N_11453);
xor U14167 (N_14167,N_9865,N_8041);
nand U14168 (N_14168,N_11037,N_11803);
or U14169 (N_14169,N_10088,N_10348);
nand U14170 (N_14170,N_10612,N_10594);
nor U14171 (N_14171,N_10532,N_11291);
nand U14172 (N_14172,N_11597,N_8960);
and U14173 (N_14173,N_11565,N_11856);
nand U14174 (N_14174,N_9924,N_11866);
and U14175 (N_14175,N_8966,N_10217);
nor U14176 (N_14176,N_10262,N_9063);
xor U14177 (N_14177,N_9514,N_9184);
nor U14178 (N_14178,N_11050,N_10468);
xor U14179 (N_14179,N_10442,N_10774);
xor U14180 (N_14180,N_9056,N_9881);
or U14181 (N_14181,N_10573,N_10306);
or U14182 (N_14182,N_10295,N_10075);
nand U14183 (N_14183,N_11586,N_10596);
xor U14184 (N_14184,N_9030,N_10293);
or U14185 (N_14185,N_8759,N_10067);
nand U14186 (N_14186,N_8306,N_10965);
nand U14187 (N_14187,N_9725,N_9599);
and U14188 (N_14188,N_10294,N_9567);
nand U14189 (N_14189,N_9058,N_11003);
nand U14190 (N_14190,N_8334,N_10620);
xnor U14191 (N_14191,N_9419,N_8010);
and U14192 (N_14192,N_11620,N_10810);
xnor U14193 (N_14193,N_8553,N_10111);
and U14194 (N_14194,N_9322,N_9548);
nand U14195 (N_14195,N_8483,N_11337);
xor U14196 (N_14196,N_11072,N_9936);
or U14197 (N_14197,N_9166,N_10723);
or U14198 (N_14198,N_11591,N_9762);
nand U14199 (N_14199,N_11586,N_11878);
xor U14200 (N_14200,N_9211,N_10129);
or U14201 (N_14201,N_8923,N_10719);
nor U14202 (N_14202,N_10792,N_9339);
xor U14203 (N_14203,N_9223,N_9709);
nand U14204 (N_14204,N_9203,N_11218);
nor U14205 (N_14205,N_9905,N_10982);
and U14206 (N_14206,N_11588,N_8470);
nand U14207 (N_14207,N_9899,N_10387);
nor U14208 (N_14208,N_11813,N_9017);
and U14209 (N_14209,N_11114,N_9189);
nor U14210 (N_14210,N_11025,N_11021);
or U14211 (N_14211,N_8732,N_10077);
and U14212 (N_14212,N_11751,N_11856);
xor U14213 (N_14213,N_9894,N_11949);
xor U14214 (N_14214,N_9077,N_9834);
and U14215 (N_14215,N_11083,N_9379);
nand U14216 (N_14216,N_8875,N_10221);
and U14217 (N_14217,N_10368,N_10846);
and U14218 (N_14218,N_10366,N_11478);
and U14219 (N_14219,N_8776,N_9424);
nand U14220 (N_14220,N_9821,N_8357);
xnor U14221 (N_14221,N_9761,N_10920);
and U14222 (N_14222,N_10402,N_8519);
or U14223 (N_14223,N_9941,N_10350);
nand U14224 (N_14224,N_11699,N_10993);
or U14225 (N_14225,N_10061,N_11126);
or U14226 (N_14226,N_8813,N_11907);
nand U14227 (N_14227,N_11863,N_10976);
and U14228 (N_14228,N_11819,N_9381);
nor U14229 (N_14229,N_11030,N_11264);
and U14230 (N_14230,N_11819,N_9369);
nand U14231 (N_14231,N_8874,N_11381);
xnor U14232 (N_14232,N_10419,N_8990);
nand U14233 (N_14233,N_11016,N_9402);
and U14234 (N_14234,N_8723,N_11091);
and U14235 (N_14235,N_10555,N_8474);
xor U14236 (N_14236,N_10297,N_10793);
or U14237 (N_14237,N_10524,N_10346);
nor U14238 (N_14238,N_10150,N_9895);
and U14239 (N_14239,N_8703,N_8839);
nand U14240 (N_14240,N_10311,N_9615);
xor U14241 (N_14241,N_9706,N_11374);
and U14242 (N_14242,N_10793,N_9326);
nor U14243 (N_14243,N_11666,N_10694);
or U14244 (N_14244,N_9980,N_9587);
and U14245 (N_14245,N_11203,N_8429);
nand U14246 (N_14246,N_9366,N_8886);
nand U14247 (N_14247,N_8805,N_10396);
xnor U14248 (N_14248,N_9523,N_8661);
nor U14249 (N_14249,N_9918,N_9763);
or U14250 (N_14250,N_9331,N_10770);
nand U14251 (N_14251,N_11943,N_8844);
or U14252 (N_14252,N_9346,N_10837);
or U14253 (N_14253,N_9081,N_11419);
or U14254 (N_14254,N_11527,N_9860);
or U14255 (N_14255,N_10632,N_11980);
or U14256 (N_14256,N_10274,N_10875);
nand U14257 (N_14257,N_11914,N_9628);
or U14258 (N_14258,N_9791,N_11906);
or U14259 (N_14259,N_11935,N_8556);
xnor U14260 (N_14260,N_11332,N_9054);
or U14261 (N_14261,N_8690,N_8829);
nand U14262 (N_14262,N_10095,N_9434);
or U14263 (N_14263,N_10323,N_10164);
nor U14264 (N_14264,N_8465,N_9340);
nor U14265 (N_14265,N_8286,N_11455);
nor U14266 (N_14266,N_8731,N_9814);
nor U14267 (N_14267,N_10821,N_8083);
and U14268 (N_14268,N_10065,N_9119);
xnor U14269 (N_14269,N_10711,N_11393);
nor U14270 (N_14270,N_8110,N_8303);
xnor U14271 (N_14271,N_11171,N_10076);
xnor U14272 (N_14272,N_11953,N_11541);
nor U14273 (N_14273,N_11573,N_11909);
nor U14274 (N_14274,N_8571,N_8977);
nand U14275 (N_14275,N_9105,N_10606);
nor U14276 (N_14276,N_8903,N_11498);
xnor U14277 (N_14277,N_11880,N_9162);
or U14278 (N_14278,N_11284,N_9586);
nor U14279 (N_14279,N_10796,N_8211);
xor U14280 (N_14280,N_8788,N_11198);
and U14281 (N_14281,N_9953,N_9496);
xnor U14282 (N_14282,N_11503,N_8586);
and U14283 (N_14283,N_11189,N_9397);
and U14284 (N_14284,N_9276,N_9742);
and U14285 (N_14285,N_9028,N_8797);
nand U14286 (N_14286,N_11799,N_10756);
or U14287 (N_14287,N_10228,N_8044);
and U14288 (N_14288,N_8800,N_9248);
or U14289 (N_14289,N_8395,N_8955);
or U14290 (N_14290,N_11458,N_10269);
and U14291 (N_14291,N_8737,N_9283);
nor U14292 (N_14292,N_10186,N_9840);
nor U14293 (N_14293,N_9132,N_10737);
nand U14294 (N_14294,N_9878,N_8350);
nand U14295 (N_14295,N_11923,N_9844);
nand U14296 (N_14296,N_11044,N_10397);
nor U14297 (N_14297,N_11828,N_9756);
nor U14298 (N_14298,N_10109,N_8452);
or U14299 (N_14299,N_9534,N_9872);
and U14300 (N_14300,N_8048,N_11602);
nand U14301 (N_14301,N_10551,N_8100);
and U14302 (N_14302,N_10191,N_8936);
nand U14303 (N_14303,N_8521,N_9927);
nor U14304 (N_14304,N_9694,N_10653);
nor U14305 (N_14305,N_8306,N_10518);
xor U14306 (N_14306,N_8273,N_8099);
or U14307 (N_14307,N_8853,N_9540);
xnor U14308 (N_14308,N_8346,N_11320);
nand U14309 (N_14309,N_9428,N_11520);
or U14310 (N_14310,N_10536,N_10673);
or U14311 (N_14311,N_8002,N_9122);
or U14312 (N_14312,N_9989,N_8327);
or U14313 (N_14313,N_10649,N_10216);
or U14314 (N_14314,N_8176,N_10320);
or U14315 (N_14315,N_10905,N_11080);
and U14316 (N_14316,N_11549,N_8123);
nand U14317 (N_14317,N_11572,N_11312);
nand U14318 (N_14318,N_11037,N_8971);
nand U14319 (N_14319,N_11988,N_9853);
and U14320 (N_14320,N_10350,N_10363);
xor U14321 (N_14321,N_8332,N_8977);
nor U14322 (N_14322,N_10064,N_9201);
xor U14323 (N_14323,N_10182,N_11591);
xnor U14324 (N_14324,N_10091,N_9754);
or U14325 (N_14325,N_9413,N_10952);
nand U14326 (N_14326,N_9919,N_8080);
or U14327 (N_14327,N_10742,N_9635);
and U14328 (N_14328,N_11369,N_9932);
and U14329 (N_14329,N_10704,N_10309);
xor U14330 (N_14330,N_11967,N_10102);
xor U14331 (N_14331,N_10949,N_10534);
and U14332 (N_14332,N_11714,N_10067);
or U14333 (N_14333,N_11515,N_8967);
nand U14334 (N_14334,N_9000,N_9216);
xor U14335 (N_14335,N_9415,N_8579);
nand U14336 (N_14336,N_8740,N_11148);
nand U14337 (N_14337,N_9734,N_8317);
nor U14338 (N_14338,N_11874,N_9342);
and U14339 (N_14339,N_8986,N_11226);
or U14340 (N_14340,N_11749,N_9771);
xnor U14341 (N_14341,N_11843,N_8998);
or U14342 (N_14342,N_11724,N_11489);
and U14343 (N_14343,N_8848,N_8647);
or U14344 (N_14344,N_10202,N_10982);
xnor U14345 (N_14345,N_10202,N_11797);
xor U14346 (N_14346,N_8515,N_11771);
and U14347 (N_14347,N_11499,N_9234);
nor U14348 (N_14348,N_8393,N_8983);
nand U14349 (N_14349,N_9944,N_9310);
nand U14350 (N_14350,N_10269,N_10616);
xnor U14351 (N_14351,N_10707,N_10694);
nor U14352 (N_14352,N_8635,N_10769);
xor U14353 (N_14353,N_8693,N_8151);
and U14354 (N_14354,N_11653,N_11067);
xor U14355 (N_14355,N_11313,N_8966);
xnor U14356 (N_14356,N_9729,N_9211);
and U14357 (N_14357,N_9829,N_8294);
and U14358 (N_14358,N_10335,N_8490);
or U14359 (N_14359,N_9666,N_11451);
and U14360 (N_14360,N_11517,N_11492);
nand U14361 (N_14361,N_8321,N_10449);
nand U14362 (N_14362,N_11165,N_9167);
or U14363 (N_14363,N_10121,N_11047);
xnor U14364 (N_14364,N_11461,N_8970);
xor U14365 (N_14365,N_11629,N_11510);
nand U14366 (N_14366,N_11517,N_9330);
xor U14367 (N_14367,N_10154,N_11228);
xor U14368 (N_14368,N_11762,N_10068);
nor U14369 (N_14369,N_9161,N_10060);
xnor U14370 (N_14370,N_11625,N_11646);
nor U14371 (N_14371,N_10715,N_8940);
xor U14372 (N_14372,N_10837,N_9877);
or U14373 (N_14373,N_8928,N_10799);
nand U14374 (N_14374,N_10582,N_8985);
nand U14375 (N_14375,N_9304,N_11023);
xor U14376 (N_14376,N_9675,N_9246);
or U14377 (N_14377,N_10950,N_9056);
or U14378 (N_14378,N_9274,N_10445);
nand U14379 (N_14379,N_10875,N_8067);
xnor U14380 (N_14380,N_8565,N_8013);
xnor U14381 (N_14381,N_11104,N_9519);
and U14382 (N_14382,N_11695,N_9393);
nor U14383 (N_14383,N_9047,N_11440);
or U14384 (N_14384,N_11643,N_8264);
nor U14385 (N_14385,N_11110,N_8267);
xor U14386 (N_14386,N_10646,N_11574);
nor U14387 (N_14387,N_10085,N_11556);
and U14388 (N_14388,N_10631,N_9465);
and U14389 (N_14389,N_10328,N_11006);
and U14390 (N_14390,N_8044,N_10358);
nand U14391 (N_14391,N_11375,N_9348);
and U14392 (N_14392,N_9338,N_9680);
nor U14393 (N_14393,N_11156,N_10421);
and U14394 (N_14394,N_10235,N_10240);
nor U14395 (N_14395,N_11306,N_10345);
or U14396 (N_14396,N_11867,N_9164);
nor U14397 (N_14397,N_9709,N_8172);
nand U14398 (N_14398,N_11188,N_11930);
nor U14399 (N_14399,N_8133,N_10102);
nor U14400 (N_14400,N_11339,N_8693);
nand U14401 (N_14401,N_8876,N_10351);
nand U14402 (N_14402,N_10014,N_8057);
or U14403 (N_14403,N_9523,N_10691);
xor U14404 (N_14404,N_10028,N_9847);
xor U14405 (N_14405,N_11082,N_10551);
nor U14406 (N_14406,N_10851,N_10135);
and U14407 (N_14407,N_8933,N_10319);
nor U14408 (N_14408,N_11580,N_9134);
xor U14409 (N_14409,N_11910,N_11036);
and U14410 (N_14410,N_11683,N_10017);
or U14411 (N_14411,N_11442,N_10409);
xnor U14412 (N_14412,N_8924,N_9453);
or U14413 (N_14413,N_9565,N_10697);
and U14414 (N_14414,N_11531,N_9350);
and U14415 (N_14415,N_11532,N_8546);
nand U14416 (N_14416,N_11081,N_10593);
nor U14417 (N_14417,N_9536,N_10283);
xnor U14418 (N_14418,N_11229,N_9863);
nand U14419 (N_14419,N_8468,N_8651);
nand U14420 (N_14420,N_8495,N_9825);
nand U14421 (N_14421,N_11277,N_11314);
nand U14422 (N_14422,N_10100,N_10842);
xor U14423 (N_14423,N_10334,N_8552);
xnor U14424 (N_14424,N_10945,N_11853);
and U14425 (N_14425,N_9766,N_9555);
nand U14426 (N_14426,N_10924,N_11895);
nor U14427 (N_14427,N_8518,N_10074);
nor U14428 (N_14428,N_8734,N_8712);
nor U14429 (N_14429,N_9332,N_11830);
or U14430 (N_14430,N_11394,N_9281);
or U14431 (N_14431,N_10269,N_10629);
nand U14432 (N_14432,N_10924,N_8821);
and U14433 (N_14433,N_9864,N_11685);
and U14434 (N_14434,N_11395,N_10067);
xnor U14435 (N_14435,N_9061,N_10880);
nand U14436 (N_14436,N_11871,N_8871);
xnor U14437 (N_14437,N_10088,N_9311);
and U14438 (N_14438,N_10833,N_11426);
nand U14439 (N_14439,N_11098,N_9767);
xnor U14440 (N_14440,N_10313,N_10774);
nand U14441 (N_14441,N_10578,N_9720);
xor U14442 (N_14442,N_10999,N_10476);
xor U14443 (N_14443,N_10877,N_10124);
nor U14444 (N_14444,N_11738,N_9325);
nand U14445 (N_14445,N_10840,N_8173);
or U14446 (N_14446,N_11954,N_11639);
nor U14447 (N_14447,N_9611,N_11905);
and U14448 (N_14448,N_10537,N_8187);
nand U14449 (N_14449,N_8265,N_10266);
and U14450 (N_14450,N_8051,N_9969);
nor U14451 (N_14451,N_11056,N_9727);
nand U14452 (N_14452,N_10162,N_10013);
or U14453 (N_14453,N_10286,N_8588);
xnor U14454 (N_14454,N_8486,N_8633);
or U14455 (N_14455,N_8595,N_9105);
and U14456 (N_14456,N_9223,N_9126);
xnor U14457 (N_14457,N_11380,N_9625);
or U14458 (N_14458,N_10559,N_10630);
or U14459 (N_14459,N_9310,N_9309);
xor U14460 (N_14460,N_11901,N_8850);
nor U14461 (N_14461,N_10295,N_10937);
xnor U14462 (N_14462,N_11807,N_10363);
xor U14463 (N_14463,N_9992,N_11637);
nor U14464 (N_14464,N_10438,N_9631);
nand U14465 (N_14465,N_9043,N_8830);
xor U14466 (N_14466,N_10479,N_9295);
or U14467 (N_14467,N_11189,N_8619);
or U14468 (N_14468,N_10591,N_8044);
xnor U14469 (N_14469,N_9247,N_10468);
xor U14470 (N_14470,N_8594,N_8086);
xor U14471 (N_14471,N_11155,N_10615);
or U14472 (N_14472,N_10318,N_11453);
xor U14473 (N_14473,N_11776,N_10701);
or U14474 (N_14474,N_10812,N_10970);
nor U14475 (N_14475,N_8520,N_8429);
nor U14476 (N_14476,N_11411,N_11871);
xnor U14477 (N_14477,N_8447,N_9576);
nor U14478 (N_14478,N_8268,N_9109);
and U14479 (N_14479,N_8988,N_8518);
nand U14480 (N_14480,N_11117,N_8711);
xnor U14481 (N_14481,N_11171,N_11131);
and U14482 (N_14482,N_10651,N_10674);
and U14483 (N_14483,N_9719,N_9075);
and U14484 (N_14484,N_10182,N_10669);
nand U14485 (N_14485,N_10714,N_11603);
nor U14486 (N_14486,N_8495,N_8068);
nand U14487 (N_14487,N_10435,N_8909);
and U14488 (N_14488,N_11726,N_9142);
nand U14489 (N_14489,N_10423,N_9749);
and U14490 (N_14490,N_11920,N_9448);
nand U14491 (N_14491,N_8550,N_8680);
nor U14492 (N_14492,N_8015,N_8429);
and U14493 (N_14493,N_8853,N_8433);
nor U14494 (N_14494,N_8639,N_10194);
nor U14495 (N_14495,N_8856,N_8624);
and U14496 (N_14496,N_10622,N_8085);
and U14497 (N_14497,N_8823,N_11135);
nand U14498 (N_14498,N_9223,N_8697);
and U14499 (N_14499,N_8327,N_9476);
xor U14500 (N_14500,N_8311,N_9036);
or U14501 (N_14501,N_10499,N_11317);
and U14502 (N_14502,N_8600,N_11572);
and U14503 (N_14503,N_10664,N_10189);
nor U14504 (N_14504,N_11059,N_9895);
nor U14505 (N_14505,N_8038,N_9175);
nand U14506 (N_14506,N_9762,N_10713);
nor U14507 (N_14507,N_9643,N_8478);
nand U14508 (N_14508,N_8947,N_9881);
or U14509 (N_14509,N_9904,N_9668);
or U14510 (N_14510,N_11817,N_10919);
nor U14511 (N_14511,N_9698,N_9420);
xor U14512 (N_14512,N_9819,N_11484);
or U14513 (N_14513,N_11097,N_8671);
xnor U14514 (N_14514,N_9060,N_10012);
and U14515 (N_14515,N_9330,N_11315);
and U14516 (N_14516,N_10270,N_10219);
nand U14517 (N_14517,N_9245,N_8798);
nand U14518 (N_14518,N_11544,N_11488);
or U14519 (N_14519,N_11361,N_9445);
nand U14520 (N_14520,N_9183,N_8573);
or U14521 (N_14521,N_8232,N_11008);
and U14522 (N_14522,N_8800,N_8473);
and U14523 (N_14523,N_9382,N_11206);
xor U14524 (N_14524,N_8630,N_8216);
nor U14525 (N_14525,N_11486,N_11387);
xor U14526 (N_14526,N_9512,N_11605);
and U14527 (N_14527,N_10712,N_10599);
xor U14528 (N_14528,N_11536,N_10718);
or U14529 (N_14529,N_11960,N_9211);
nand U14530 (N_14530,N_10885,N_11191);
and U14531 (N_14531,N_10043,N_8584);
xor U14532 (N_14532,N_11059,N_9522);
xor U14533 (N_14533,N_8488,N_8919);
nand U14534 (N_14534,N_8871,N_10984);
and U14535 (N_14535,N_11643,N_9484);
and U14536 (N_14536,N_10023,N_10006);
and U14537 (N_14537,N_8923,N_10910);
or U14538 (N_14538,N_9058,N_11358);
and U14539 (N_14539,N_8706,N_9257);
xnor U14540 (N_14540,N_8418,N_11143);
nand U14541 (N_14541,N_8967,N_9121);
xor U14542 (N_14542,N_9456,N_11440);
and U14543 (N_14543,N_11391,N_11131);
nor U14544 (N_14544,N_8118,N_10571);
and U14545 (N_14545,N_11450,N_11708);
nor U14546 (N_14546,N_10529,N_9874);
and U14547 (N_14547,N_9570,N_11995);
and U14548 (N_14548,N_10680,N_8550);
nor U14549 (N_14549,N_9088,N_8821);
xor U14550 (N_14550,N_11282,N_9735);
nand U14551 (N_14551,N_10149,N_8612);
nand U14552 (N_14552,N_11283,N_10182);
nand U14553 (N_14553,N_10028,N_10445);
xor U14554 (N_14554,N_11420,N_10188);
and U14555 (N_14555,N_11613,N_9981);
or U14556 (N_14556,N_8471,N_10488);
nand U14557 (N_14557,N_9209,N_11076);
nor U14558 (N_14558,N_9832,N_11250);
xor U14559 (N_14559,N_11805,N_8552);
nor U14560 (N_14560,N_8402,N_9477);
nor U14561 (N_14561,N_11789,N_8541);
and U14562 (N_14562,N_11843,N_8634);
nor U14563 (N_14563,N_9335,N_8775);
nor U14564 (N_14564,N_11450,N_9083);
and U14565 (N_14565,N_8577,N_8221);
xor U14566 (N_14566,N_9066,N_8249);
and U14567 (N_14567,N_9841,N_11414);
xnor U14568 (N_14568,N_9401,N_11671);
nor U14569 (N_14569,N_10174,N_11156);
nor U14570 (N_14570,N_8279,N_8485);
and U14571 (N_14571,N_8739,N_10322);
xnor U14572 (N_14572,N_9173,N_9006);
and U14573 (N_14573,N_9849,N_8667);
and U14574 (N_14574,N_11278,N_8671);
nor U14575 (N_14575,N_9725,N_11208);
nand U14576 (N_14576,N_10016,N_10317);
nor U14577 (N_14577,N_10330,N_11155);
xnor U14578 (N_14578,N_11308,N_11660);
nand U14579 (N_14579,N_9031,N_8083);
or U14580 (N_14580,N_10267,N_9273);
nand U14581 (N_14581,N_10956,N_10872);
nand U14582 (N_14582,N_9291,N_9050);
nand U14583 (N_14583,N_10004,N_9885);
and U14584 (N_14584,N_11690,N_11038);
nor U14585 (N_14585,N_11315,N_8895);
xor U14586 (N_14586,N_8130,N_8246);
or U14587 (N_14587,N_11678,N_11260);
xnor U14588 (N_14588,N_11124,N_11166);
xnor U14589 (N_14589,N_8279,N_9222);
nor U14590 (N_14590,N_10026,N_9752);
xor U14591 (N_14591,N_10187,N_8691);
and U14592 (N_14592,N_10283,N_8448);
xor U14593 (N_14593,N_11617,N_8855);
nor U14594 (N_14594,N_10680,N_10231);
nor U14595 (N_14595,N_8024,N_9308);
nor U14596 (N_14596,N_8687,N_8938);
nand U14597 (N_14597,N_9133,N_9364);
nor U14598 (N_14598,N_11129,N_11340);
and U14599 (N_14599,N_9522,N_10676);
and U14600 (N_14600,N_10092,N_11657);
nor U14601 (N_14601,N_8965,N_8474);
nor U14602 (N_14602,N_10732,N_8606);
nand U14603 (N_14603,N_8457,N_8159);
and U14604 (N_14604,N_10271,N_10748);
xnor U14605 (N_14605,N_11733,N_10543);
nor U14606 (N_14606,N_10382,N_9136);
and U14607 (N_14607,N_9973,N_8174);
xor U14608 (N_14608,N_10762,N_9004);
nand U14609 (N_14609,N_8733,N_8514);
nand U14610 (N_14610,N_10457,N_10925);
and U14611 (N_14611,N_10822,N_11006);
and U14612 (N_14612,N_11326,N_10157);
and U14613 (N_14613,N_11501,N_8983);
or U14614 (N_14614,N_11745,N_11862);
or U14615 (N_14615,N_9055,N_8732);
xor U14616 (N_14616,N_8645,N_9529);
nand U14617 (N_14617,N_11220,N_9966);
or U14618 (N_14618,N_10731,N_11937);
xor U14619 (N_14619,N_11670,N_8721);
xor U14620 (N_14620,N_11483,N_10880);
and U14621 (N_14621,N_8290,N_9752);
or U14622 (N_14622,N_10667,N_11860);
xnor U14623 (N_14623,N_8687,N_9215);
or U14624 (N_14624,N_11346,N_10307);
xnor U14625 (N_14625,N_10833,N_10689);
xnor U14626 (N_14626,N_9047,N_8879);
and U14627 (N_14627,N_9289,N_8369);
nand U14628 (N_14628,N_9490,N_11591);
xor U14629 (N_14629,N_8352,N_10582);
and U14630 (N_14630,N_9049,N_9618);
or U14631 (N_14631,N_11009,N_11731);
and U14632 (N_14632,N_8072,N_11885);
xnor U14633 (N_14633,N_10668,N_10974);
and U14634 (N_14634,N_10274,N_10796);
nand U14635 (N_14635,N_10566,N_9544);
xnor U14636 (N_14636,N_9507,N_9984);
and U14637 (N_14637,N_8386,N_11451);
nor U14638 (N_14638,N_9774,N_9200);
nor U14639 (N_14639,N_9829,N_8382);
or U14640 (N_14640,N_9985,N_10633);
nand U14641 (N_14641,N_10158,N_11382);
or U14642 (N_14642,N_11414,N_10303);
xnor U14643 (N_14643,N_11697,N_9857);
xor U14644 (N_14644,N_8443,N_10296);
and U14645 (N_14645,N_8095,N_8972);
nand U14646 (N_14646,N_8498,N_11998);
and U14647 (N_14647,N_9018,N_11918);
nor U14648 (N_14648,N_8356,N_11241);
or U14649 (N_14649,N_10757,N_9959);
and U14650 (N_14650,N_8388,N_8136);
nand U14651 (N_14651,N_11289,N_11656);
xor U14652 (N_14652,N_11914,N_8205);
xor U14653 (N_14653,N_9626,N_10493);
xnor U14654 (N_14654,N_10919,N_10964);
nand U14655 (N_14655,N_9653,N_9765);
nand U14656 (N_14656,N_10549,N_9982);
and U14657 (N_14657,N_8429,N_11805);
nand U14658 (N_14658,N_8612,N_8785);
or U14659 (N_14659,N_10566,N_8881);
or U14660 (N_14660,N_8508,N_10855);
nand U14661 (N_14661,N_8850,N_9820);
xor U14662 (N_14662,N_11683,N_8649);
and U14663 (N_14663,N_8650,N_10352);
and U14664 (N_14664,N_9634,N_11143);
xor U14665 (N_14665,N_8534,N_11656);
and U14666 (N_14666,N_9058,N_10492);
and U14667 (N_14667,N_9937,N_9291);
and U14668 (N_14668,N_10937,N_10236);
xor U14669 (N_14669,N_9065,N_11039);
nor U14670 (N_14670,N_8691,N_9758);
and U14671 (N_14671,N_10224,N_10786);
nand U14672 (N_14672,N_9198,N_8826);
nand U14673 (N_14673,N_9891,N_8939);
xnor U14674 (N_14674,N_9166,N_11006);
nor U14675 (N_14675,N_9208,N_10120);
xor U14676 (N_14676,N_11744,N_10216);
xnor U14677 (N_14677,N_11691,N_10147);
and U14678 (N_14678,N_8885,N_10947);
and U14679 (N_14679,N_8322,N_11506);
and U14680 (N_14680,N_8778,N_11798);
or U14681 (N_14681,N_8929,N_8524);
nand U14682 (N_14682,N_11555,N_8983);
nor U14683 (N_14683,N_9897,N_8569);
or U14684 (N_14684,N_9514,N_10540);
xor U14685 (N_14685,N_9203,N_10331);
nor U14686 (N_14686,N_11731,N_10307);
or U14687 (N_14687,N_8167,N_11202);
nand U14688 (N_14688,N_11212,N_10603);
or U14689 (N_14689,N_9332,N_8421);
xor U14690 (N_14690,N_9804,N_8356);
and U14691 (N_14691,N_8299,N_11881);
or U14692 (N_14692,N_8881,N_8053);
or U14693 (N_14693,N_8437,N_9540);
xor U14694 (N_14694,N_9813,N_8989);
xor U14695 (N_14695,N_10333,N_9501);
nor U14696 (N_14696,N_9632,N_10487);
or U14697 (N_14697,N_11636,N_8150);
nand U14698 (N_14698,N_8272,N_10540);
nand U14699 (N_14699,N_10163,N_9086);
and U14700 (N_14700,N_11488,N_10039);
xnor U14701 (N_14701,N_11925,N_8202);
and U14702 (N_14702,N_9290,N_10882);
nor U14703 (N_14703,N_8522,N_11974);
or U14704 (N_14704,N_9062,N_10195);
and U14705 (N_14705,N_9038,N_11019);
xnor U14706 (N_14706,N_10313,N_11179);
nand U14707 (N_14707,N_9627,N_10445);
xnor U14708 (N_14708,N_10326,N_8574);
or U14709 (N_14709,N_9833,N_11136);
nor U14710 (N_14710,N_11115,N_11957);
or U14711 (N_14711,N_11175,N_11434);
or U14712 (N_14712,N_9463,N_10839);
and U14713 (N_14713,N_10217,N_10527);
or U14714 (N_14714,N_11027,N_10787);
nand U14715 (N_14715,N_9207,N_10695);
nand U14716 (N_14716,N_8204,N_9054);
or U14717 (N_14717,N_10491,N_9749);
xnor U14718 (N_14718,N_11678,N_10670);
nand U14719 (N_14719,N_9076,N_11412);
or U14720 (N_14720,N_10397,N_11012);
nand U14721 (N_14721,N_8585,N_10869);
or U14722 (N_14722,N_8345,N_8663);
xor U14723 (N_14723,N_8073,N_8103);
xnor U14724 (N_14724,N_10027,N_10939);
nand U14725 (N_14725,N_11516,N_8887);
xor U14726 (N_14726,N_11161,N_10864);
xor U14727 (N_14727,N_11060,N_8569);
and U14728 (N_14728,N_11558,N_8677);
and U14729 (N_14729,N_10315,N_9654);
xor U14730 (N_14730,N_10319,N_10533);
nor U14731 (N_14731,N_11914,N_11721);
xnor U14732 (N_14732,N_10697,N_11900);
nand U14733 (N_14733,N_10395,N_9622);
nand U14734 (N_14734,N_11934,N_11135);
or U14735 (N_14735,N_11108,N_11558);
or U14736 (N_14736,N_11398,N_8012);
and U14737 (N_14737,N_9484,N_8278);
xnor U14738 (N_14738,N_9064,N_9917);
nor U14739 (N_14739,N_8879,N_9308);
xor U14740 (N_14740,N_10859,N_8779);
xor U14741 (N_14741,N_11664,N_10828);
nand U14742 (N_14742,N_9152,N_10785);
or U14743 (N_14743,N_11069,N_8552);
or U14744 (N_14744,N_8731,N_10078);
or U14745 (N_14745,N_11378,N_11698);
and U14746 (N_14746,N_8176,N_9290);
nor U14747 (N_14747,N_9634,N_10685);
nor U14748 (N_14748,N_9231,N_8494);
and U14749 (N_14749,N_10090,N_11541);
and U14750 (N_14750,N_10542,N_9784);
or U14751 (N_14751,N_10077,N_9639);
xnor U14752 (N_14752,N_10939,N_10726);
nand U14753 (N_14753,N_8009,N_11317);
nand U14754 (N_14754,N_8606,N_8904);
or U14755 (N_14755,N_10363,N_8543);
and U14756 (N_14756,N_10001,N_8333);
nand U14757 (N_14757,N_11361,N_10494);
nor U14758 (N_14758,N_10651,N_11973);
and U14759 (N_14759,N_8794,N_10620);
nor U14760 (N_14760,N_10498,N_8686);
nand U14761 (N_14761,N_8762,N_10890);
or U14762 (N_14762,N_11506,N_10218);
or U14763 (N_14763,N_8452,N_10228);
xor U14764 (N_14764,N_10065,N_8076);
nor U14765 (N_14765,N_10471,N_9364);
or U14766 (N_14766,N_11880,N_9046);
or U14767 (N_14767,N_8109,N_11488);
xnor U14768 (N_14768,N_10584,N_10686);
nor U14769 (N_14769,N_10977,N_8143);
xnor U14770 (N_14770,N_9404,N_10995);
nor U14771 (N_14771,N_9393,N_11028);
or U14772 (N_14772,N_11581,N_8307);
or U14773 (N_14773,N_10764,N_11190);
nand U14774 (N_14774,N_8897,N_9796);
and U14775 (N_14775,N_9349,N_8462);
and U14776 (N_14776,N_8035,N_10843);
xor U14777 (N_14777,N_11428,N_9329);
nor U14778 (N_14778,N_10458,N_11730);
nor U14779 (N_14779,N_9378,N_8323);
xor U14780 (N_14780,N_9260,N_8211);
or U14781 (N_14781,N_11192,N_9930);
xor U14782 (N_14782,N_11778,N_9473);
nand U14783 (N_14783,N_8890,N_11346);
or U14784 (N_14784,N_11354,N_9465);
or U14785 (N_14785,N_8632,N_11618);
nand U14786 (N_14786,N_10451,N_8149);
and U14787 (N_14787,N_10584,N_8748);
nor U14788 (N_14788,N_9511,N_11342);
and U14789 (N_14789,N_10241,N_9864);
xor U14790 (N_14790,N_11470,N_11253);
nand U14791 (N_14791,N_9035,N_11146);
nand U14792 (N_14792,N_8020,N_11865);
nand U14793 (N_14793,N_10857,N_10248);
and U14794 (N_14794,N_8749,N_11543);
and U14795 (N_14795,N_10516,N_9255);
nand U14796 (N_14796,N_11112,N_9698);
nand U14797 (N_14797,N_8144,N_9330);
and U14798 (N_14798,N_9918,N_11554);
xnor U14799 (N_14799,N_10423,N_9751);
nor U14800 (N_14800,N_8405,N_11530);
xor U14801 (N_14801,N_11916,N_10687);
or U14802 (N_14802,N_11152,N_8703);
and U14803 (N_14803,N_10488,N_9429);
and U14804 (N_14804,N_9166,N_9480);
xor U14805 (N_14805,N_10117,N_11097);
or U14806 (N_14806,N_10402,N_8141);
nor U14807 (N_14807,N_9363,N_9075);
xnor U14808 (N_14808,N_11222,N_8318);
xor U14809 (N_14809,N_9544,N_10849);
or U14810 (N_14810,N_9874,N_10013);
nand U14811 (N_14811,N_8568,N_10722);
or U14812 (N_14812,N_8486,N_11045);
nor U14813 (N_14813,N_9083,N_11449);
nand U14814 (N_14814,N_8602,N_10099);
xnor U14815 (N_14815,N_10840,N_11325);
or U14816 (N_14816,N_10383,N_8652);
nand U14817 (N_14817,N_10941,N_11104);
nand U14818 (N_14818,N_11375,N_8386);
nor U14819 (N_14819,N_9191,N_9185);
or U14820 (N_14820,N_11531,N_11595);
xnor U14821 (N_14821,N_9669,N_10408);
xnor U14822 (N_14822,N_10231,N_9559);
xor U14823 (N_14823,N_11719,N_9614);
and U14824 (N_14824,N_10806,N_8197);
nand U14825 (N_14825,N_8626,N_9798);
and U14826 (N_14826,N_11229,N_11190);
nand U14827 (N_14827,N_9838,N_10212);
nor U14828 (N_14828,N_10698,N_10127);
or U14829 (N_14829,N_8923,N_9835);
xnor U14830 (N_14830,N_9754,N_8942);
and U14831 (N_14831,N_9611,N_10668);
xor U14832 (N_14832,N_8626,N_11078);
and U14833 (N_14833,N_10872,N_9139);
or U14834 (N_14834,N_8173,N_11156);
and U14835 (N_14835,N_10631,N_10504);
nand U14836 (N_14836,N_8592,N_10327);
or U14837 (N_14837,N_9502,N_9174);
nor U14838 (N_14838,N_10188,N_8544);
nor U14839 (N_14839,N_9825,N_11392);
nand U14840 (N_14840,N_9666,N_10762);
and U14841 (N_14841,N_10632,N_9866);
and U14842 (N_14842,N_8769,N_10747);
nor U14843 (N_14843,N_8704,N_11324);
or U14844 (N_14844,N_9956,N_9629);
xor U14845 (N_14845,N_11272,N_8138);
or U14846 (N_14846,N_9686,N_10287);
or U14847 (N_14847,N_10662,N_10150);
nor U14848 (N_14848,N_10120,N_11553);
or U14849 (N_14849,N_9171,N_11514);
and U14850 (N_14850,N_10161,N_10311);
nor U14851 (N_14851,N_11091,N_8919);
nor U14852 (N_14852,N_11123,N_10690);
xor U14853 (N_14853,N_8833,N_11257);
or U14854 (N_14854,N_8349,N_10660);
nor U14855 (N_14855,N_11912,N_11079);
or U14856 (N_14856,N_10977,N_11364);
or U14857 (N_14857,N_8618,N_10635);
or U14858 (N_14858,N_9497,N_8226);
or U14859 (N_14859,N_10782,N_11840);
or U14860 (N_14860,N_11718,N_11628);
and U14861 (N_14861,N_11033,N_10752);
and U14862 (N_14862,N_11171,N_8385);
nor U14863 (N_14863,N_9666,N_10709);
or U14864 (N_14864,N_8811,N_8837);
nor U14865 (N_14865,N_10998,N_9528);
or U14866 (N_14866,N_10737,N_11724);
and U14867 (N_14867,N_11972,N_10938);
and U14868 (N_14868,N_10332,N_8003);
nor U14869 (N_14869,N_9194,N_10641);
xnor U14870 (N_14870,N_11849,N_11507);
nor U14871 (N_14871,N_9758,N_8400);
nand U14872 (N_14872,N_10728,N_10529);
nor U14873 (N_14873,N_11230,N_11456);
xor U14874 (N_14874,N_10697,N_8550);
nand U14875 (N_14875,N_10736,N_8932);
xnor U14876 (N_14876,N_8754,N_8116);
and U14877 (N_14877,N_10644,N_11998);
nand U14878 (N_14878,N_10956,N_10107);
and U14879 (N_14879,N_8235,N_10429);
xor U14880 (N_14880,N_9533,N_11403);
xor U14881 (N_14881,N_9814,N_8886);
nand U14882 (N_14882,N_10420,N_11104);
xnor U14883 (N_14883,N_8930,N_8978);
nor U14884 (N_14884,N_9575,N_8866);
nor U14885 (N_14885,N_11176,N_8236);
xnor U14886 (N_14886,N_8967,N_11340);
xor U14887 (N_14887,N_9426,N_11639);
or U14888 (N_14888,N_11965,N_9287);
or U14889 (N_14889,N_10502,N_10929);
nor U14890 (N_14890,N_8952,N_10573);
xnor U14891 (N_14891,N_11245,N_11074);
nor U14892 (N_14892,N_10768,N_9478);
nand U14893 (N_14893,N_8354,N_11234);
xnor U14894 (N_14894,N_8935,N_10357);
nand U14895 (N_14895,N_9476,N_11813);
nand U14896 (N_14896,N_8251,N_8205);
nand U14897 (N_14897,N_11041,N_8506);
nand U14898 (N_14898,N_9622,N_10005);
nor U14899 (N_14899,N_11763,N_10141);
nand U14900 (N_14900,N_10037,N_9148);
and U14901 (N_14901,N_11916,N_11761);
or U14902 (N_14902,N_11124,N_8826);
xor U14903 (N_14903,N_8499,N_8291);
xnor U14904 (N_14904,N_11293,N_10633);
nor U14905 (N_14905,N_11809,N_9280);
or U14906 (N_14906,N_8078,N_8688);
xor U14907 (N_14907,N_10405,N_9640);
xnor U14908 (N_14908,N_9197,N_10784);
nand U14909 (N_14909,N_9786,N_10548);
nand U14910 (N_14910,N_8493,N_10935);
or U14911 (N_14911,N_9091,N_10827);
xnor U14912 (N_14912,N_10603,N_8302);
nor U14913 (N_14913,N_8040,N_11766);
or U14914 (N_14914,N_9540,N_10565);
and U14915 (N_14915,N_9668,N_10775);
xor U14916 (N_14916,N_11210,N_11092);
and U14917 (N_14917,N_9024,N_9980);
and U14918 (N_14918,N_11969,N_10263);
or U14919 (N_14919,N_8436,N_11674);
or U14920 (N_14920,N_8140,N_8534);
nor U14921 (N_14921,N_11212,N_9283);
xor U14922 (N_14922,N_9697,N_10909);
and U14923 (N_14923,N_8792,N_11556);
nor U14924 (N_14924,N_11492,N_11925);
xnor U14925 (N_14925,N_9114,N_10227);
and U14926 (N_14926,N_10310,N_10072);
xor U14927 (N_14927,N_11047,N_9928);
and U14928 (N_14928,N_11231,N_8982);
nor U14929 (N_14929,N_10619,N_9139);
and U14930 (N_14930,N_9037,N_11058);
nor U14931 (N_14931,N_9715,N_11757);
nand U14932 (N_14932,N_10168,N_8332);
nand U14933 (N_14933,N_11142,N_8631);
nand U14934 (N_14934,N_8648,N_8263);
xnor U14935 (N_14935,N_11111,N_8751);
nand U14936 (N_14936,N_8021,N_9982);
and U14937 (N_14937,N_10277,N_8896);
and U14938 (N_14938,N_9069,N_9946);
and U14939 (N_14939,N_9259,N_10774);
nand U14940 (N_14940,N_9818,N_8204);
nand U14941 (N_14941,N_11188,N_9249);
nor U14942 (N_14942,N_9644,N_11642);
nand U14943 (N_14943,N_11616,N_10561);
xnor U14944 (N_14944,N_9770,N_10477);
nand U14945 (N_14945,N_11615,N_8685);
and U14946 (N_14946,N_8936,N_11855);
and U14947 (N_14947,N_11754,N_8117);
or U14948 (N_14948,N_10462,N_8386);
xnor U14949 (N_14949,N_10635,N_8651);
and U14950 (N_14950,N_9709,N_9063);
nand U14951 (N_14951,N_10505,N_9120);
and U14952 (N_14952,N_10983,N_11257);
or U14953 (N_14953,N_9620,N_8396);
nand U14954 (N_14954,N_9512,N_9054);
and U14955 (N_14955,N_11582,N_10949);
nand U14956 (N_14956,N_9877,N_9560);
nor U14957 (N_14957,N_9704,N_10494);
nand U14958 (N_14958,N_11245,N_8264);
xor U14959 (N_14959,N_11273,N_11864);
nand U14960 (N_14960,N_9694,N_8557);
nor U14961 (N_14961,N_9510,N_9701);
or U14962 (N_14962,N_11514,N_9771);
nor U14963 (N_14963,N_8317,N_11662);
xnor U14964 (N_14964,N_8963,N_11382);
nand U14965 (N_14965,N_9499,N_9170);
nand U14966 (N_14966,N_11760,N_10518);
xor U14967 (N_14967,N_9728,N_10257);
and U14968 (N_14968,N_10763,N_11960);
and U14969 (N_14969,N_10857,N_8338);
nor U14970 (N_14970,N_10829,N_11255);
and U14971 (N_14971,N_8400,N_9261);
nand U14972 (N_14972,N_10208,N_10652);
nand U14973 (N_14973,N_8364,N_10965);
or U14974 (N_14974,N_11408,N_9826);
and U14975 (N_14975,N_11399,N_10151);
nand U14976 (N_14976,N_10317,N_8132);
nand U14977 (N_14977,N_9167,N_8509);
nor U14978 (N_14978,N_10441,N_9578);
and U14979 (N_14979,N_11558,N_11146);
xnor U14980 (N_14980,N_8706,N_9736);
nand U14981 (N_14981,N_9990,N_8851);
nand U14982 (N_14982,N_9735,N_9897);
nand U14983 (N_14983,N_10860,N_10862);
xnor U14984 (N_14984,N_8020,N_9426);
or U14985 (N_14985,N_10860,N_10478);
xor U14986 (N_14986,N_9376,N_11996);
and U14987 (N_14987,N_9065,N_9264);
xor U14988 (N_14988,N_11485,N_11345);
xnor U14989 (N_14989,N_9674,N_9799);
nor U14990 (N_14990,N_10415,N_8512);
xnor U14991 (N_14991,N_10037,N_8530);
nand U14992 (N_14992,N_8006,N_9726);
xnor U14993 (N_14993,N_10580,N_9127);
and U14994 (N_14994,N_10849,N_10391);
and U14995 (N_14995,N_10197,N_10787);
xnor U14996 (N_14996,N_9577,N_9868);
or U14997 (N_14997,N_8139,N_11013);
nor U14998 (N_14998,N_10700,N_9863);
or U14999 (N_14999,N_10624,N_10310);
xnor U15000 (N_15000,N_11017,N_10969);
or U15001 (N_15001,N_8277,N_9500);
or U15002 (N_15002,N_9504,N_9834);
nor U15003 (N_15003,N_11117,N_9892);
xnor U15004 (N_15004,N_8969,N_11208);
xnor U15005 (N_15005,N_8967,N_11217);
nand U15006 (N_15006,N_8268,N_11370);
and U15007 (N_15007,N_11716,N_9342);
and U15008 (N_15008,N_10262,N_9113);
and U15009 (N_15009,N_11293,N_11116);
or U15010 (N_15010,N_11799,N_9344);
xnor U15011 (N_15011,N_10063,N_11135);
and U15012 (N_15012,N_9223,N_10353);
nor U15013 (N_15013,N_9831,N_10626);
nand U15014 (N_15014,N_11429,N_8533);
xnor U15015 (N_15015,N_8059,N_10757);
xor U15016 (N_15016,N_9648,N_10291);
and U15017 (N_15017,N_10200,N_8595);
nor U15018 (N_15018,N_8221,N_9883);
nand U15019 (N_15019,N_11278,N_9956);
and U15020 (N_15020,N_8131,N_10357);
nor U15021 (N_15021,N_10318,N_10862);
nor U15022 (N_15022,N_8369,N_10746);
nor U15023 (N_15023,N_9242,N_9256);
or U15024 (N_15024,N_10559,N_9907);
nand U15025 (N_15025,N_10485,N_10701);
nor U15026 (N_15026,N_11128,N_11099);
nand U15027 (N_15027,N_10553,N_9197);
nor U15028 (N_15028,N_10784,N_11103);
or U15029 (N_15029,N_11027,N_11217);
and U15030 (N_15030,N_9851,N_11245);
xor U15031 (N_15031,N_9420,N_10799);
nand U15032 (N_15032,N_8991,N_8879);
nand U15033 (N_15033,N_9324,N_10957);
or U15034 (N_15034,N_10406,N_11219);
nand U15035 (N_15035,N_9474,N_8715);
xnor U15036 (N_15036,N_9978,N_11167);
xnor U15037 (N_15037,N_11410,N_9162);
and U15038 (N_15038,N_9636,N_8825);
xor U15039 (N_15039,N_8397,N_11707);
and U15040 (N_15040,N_9192,N_10238);
and U15041 (N_15041,N_9490,N_8997);
nand U15042 (N_15042,N_10308,N_10505);
and U15043 (N_15043,N_10366,N_11599);
xnor U15044 (N_15044,N_8967,N_10054);
and U15045 (N_15045,N_11819,N_8686);
and U15046 (N_15046,N_11023,N_11905);
and U15047 (N_15047,N_11797,N_10353);
and U15048 (N_15048,N_9668,N_11831);
or U15049 (N_15049,N_11161,N_8764);
nor U15050 (N_15050,N_9671,N_9526);
nor U15051 (N_15051,N_8048,N_9632);
or U15052 (N_15052,N_10324,N_11051);
and U15053 (N_15053,N_8415,N_8192);
xnor U15054 (N_15054,N_11234,N_9711);
xnor U15055 (N_15055,N_8341,N_9684);
nand U15056 (N_15056,N_11553,N_9385);
nand U15057 (N_15057,N_11815,N_10125);
nand U15058 (N_15058,N_9540,N_10709);
nand U15059 (N_15059,N_8390,N_9695);
nor U15060 (N_15060,N_10706,N_8665);
nand U15061 (N_15061,N_8499,N_10692);
nand U15062 (N_15062,N_11527,N_10849);
xor U15063 (N_15063,N_9731,N_9113);
nand U15064 (N_15064,N_11432,N_8698);
nor U15065 (N_15065,N_10872,N_9035);
xor U15066 (N_15066,N_9069,N_9412);
and U15067 (N_15067,N_8798,N_11220);
or U15068 (N_15068,N_11117,N_9065);
nor U15069 (N_15069,N_11720,N_9935);
and U15070 (N_15070,N_10528,N_11999);
or U15071 (N_15071,N_10318,N_11541);
nor U15072 (N_15072,N_11529,N_8890);
xor U15073 (N_15073,N_10021,N_11361);
xnor U15074 (N_15074,N_11245,N_10905);
nand U15075 (N_15075,N_8932,N_8167);
and U15076 (N_15076,N_10571,N_11232);
nor U15077 (N_15077,N_8662,N_11878);
nand U15078 (N_15078,N_8008,N_10452);
or U15079 (N_15079,N_9097,N_11204);
or U15080 (N_15080,N_11833,N_10580);
nor U15081 (N_15081,N_10484,N_11163);
nor U15082 (N_15082,N_8356,N_9281);
and U15083 (N_15083,N_11603,N_9497);
nor U15084 (N_15084,N_9585,N_11678);
and U15085 (N_15085,N_9505,N_9199);
nand U15086 (N_15086,N_11254,N_9515);
or U15087 (N_15087,N_9030,N_9812);
or U15088 (N_15088,N_9751,N_8295);
and U15089 (N_15089,N_9614,N_8550);
and U15090 (N_15090,N_10024,N_8469);
or U15091 (N_15091,N_9542,N_9021);
nand U15092 (N_15092,N_8981,N_8137);
xnor U15093 (N_15093,N_10637,N_11579);
nand U15094 (N_15094,N_11897,N_9901);
nor U15095 (N_15095,N_8368,N_9461);
or U15096 (N_15096,N_9277,N_11006);
nand U15097 (N_15097,N_10974,N_8549);
nand U15098 (N_15098,N_10916,N_8413);
xor U15099 (N_15099,N_9942,N_10778);
xor U15100 (N_15100,N_11784,N_8512);
and U15101 (N_15101,N_8648,N_10471);
nor U15102 (N_15102,N_10590,N_11021);
nor U15103 (N_15103,N_11634,N_10372);
nor U15104 (N_15104,N_10587,N_8116);
nor U15105 (N_15105,N_9857,N_10461);
nor U15106 (N_15106,N_10905,N_11741);
xnor U15107 (N_15107,N_9897,N_11186);
xor U15108 (N_15108,N_11202,N_10685);
xnor U15109 (N_15109,N_8378,N_9764);
xnor U15110 (N_15110,N_10287,N_9124);
and U15111 (N_15111,N_11305,N_9216);
or U15112 (N_15112,N_9160,N_10980);
nor U15113 (N_15113,N_8799,N_10351);
nor U15114 (N_15114,N_9356,N_8687);
nand U15115 (N_15115,N_10960,N_11905);
nand U15116 (N_15116,N_11760,N_10860);
xnor U15117 (N_15117,N_10851,N_10887);
nor U15118 (N_15118,N_8946,N_11701);
and U15119 (N_15119,N_9663,N_10501);
nor U15120 (N_15120,N_9504,N_9799);
and U15121 (N_15121,N_11579,N_9238);
nand U15122 (N_15122,N_10436,N_11003);
nand U15123 (N_15123,N_8754,N_10055);
or U15124 (N_15124,N_9376,N_9214);
or U15125 (N_15125,N_9095,N_10696);
xor U15126 (N_15126,N_8760,N_11907);
xor U15127 (N_15127,N_11093,N_10154);
nand U15128 (N_15128,N_9323,N_8666);
xnor U15129 (N_15129,N_11886,N_11985);
nor U15130 (N_15130,N_8201,N_9848);
nand U15131 (N_15131,N_9880,N_11266);
and U15132 (N_15132,N_8547,N_9315);
nand U15133 (N_15133,N_11360,N_8443);
nand U15134 (N_15134,N_11325,N_11405);
nand U15135 (N_15135,N_8000,N_10374);
or U15136 (N_15136,N_10971,N_9665);
or U15137 (N_15137,N_10032,N_10261);
or U15138 (N_15138,N_9382,N_11583);
nor U15139 (N_15139,N_10086,N_9323);
nor U15140 (N_15140,N_10044,N_11195);
xnor U15141 (N_15141,N_11675,N_9167);
xnor U15142 (N_15142,N_8275,N_9088);
nor U15143 (N_15143,N_9259,N_9777);
or U15144 (N_15144,N_10594,N_10642);
nand U15145 (N_15145,N_11046,N_8083);
or U15146 (N_15146,N_9893,N_11744);
nor U15147 (N_15147,N_8876,N_11812);
xnor U15148 (N_15148,N_11235,N_8272);
and U15149 (N_15149,N_10110,N_11294);
nand U15150 (N_15150,N_11323,N_9223);
and U15151 (N_15151,N_11993,N_8469);
and U15152 (N_15152,N_9799,N_9053);
or U15153 (N_15153,N_9042,N_9808);
xor U15154 (N_15154,N_9417,N_9952);
xor U15155 (N_15155,N_9468,N_11834);
or U15156 (N_15156,N_8326,N_10823);
or U15157 (N_15157,N_8397,N_9804);
or U15158 (N_15158,N_11117,N_9738);
and U15159 (N_15159,N_11655,N_8388);
and U15160 (N_15160,N_8902,N_10200);
nor U15161 (N_15161,N_8422,N_10835);
or U15162 (N_15162,N_8337,N_9201);
nor U15163 (N_15163,N_8492,N_10572);
nand U15164 (N_15164,N_10476,N_11311);
xor U15165 (N_15165,N_8734,N_9812);
or U15166 (N_15166,N_11879,N_9260);
nor U15167 (N_15167,N_9237,N_8546);
nor U15168 (N_15168,N_9637,N_9039);
xnor U15169 (N_15169,N_9708,N_8605);
and U15170 (N_15170,N_10741,N_10051);
and U15171 (N_15171,N_11517,N_8526);
xnor U15172 (N_15172,N_11735,N_10178);
and U15173 (N_15173,N_8049,N_11931);
or U15174 (N_15174,N_9983,N_11986);
xnor U15175 (N_15175,N_10745,N_11834);
or U15176 (N_15176,N_9040,N_10872);
xor U15177 (N_15177,N_11518,N_11205);
or U15178 (N_15178,N_10076,N_11791);
and U15179 (N_15179,N_10375,N_11846);
nand U15180 (N_15180,N_10505,N_9876);
or U15181 (N_15181,N_9685,N_10149);
nor U15182 (N_15182,N_10381,N_8665);
nor U15183 (N_15183,N_10027,N_11423);
xnor U15184 (N_15184,N_9486,N_10511);
nand U15185 (N_15185,N_10747,N_10359);
nand U15186 (N_15186,N_10137,N_11599);
and U15187 (N_15187,N_9074,N_10948);
nand U15188 (N_15188,N_9432,N_9296);
xnor U15189 (N_15189,N_10474,N_11587);
or U15190 (N_15190,N_8333,N_11604);
and U15191 (N_15191,N_8493,N_8337);
and U15192 (N_15192,N_8962,N_8407);
and U15193 (N_15193,N_9731,N_11003);
or U15194 (N_15194,N_10444,N_10872);
or U15195 (N_15195,N_10046,N_8805);
nor U15196 (N_15196,N_8137,N_11239);
nor U15197 (N_15197,N_9589,N_9750);
or U15198 (N_15198,N_8108,N_8419);
nor U15199 (N_15199,N_8002,N_11465);
nor U15200 (N_15200,N_11881,N_9828);
or U15201 (N_15201,N_9429,N_8265);
nor U15202 (N_15202,N_10057,N_11141);
nand U15203 (N_15203,N_8935,N_10752);
nand U15204 (N_15204,N_8345,N_11998);
or U15205 (N_15205,N_8872,N_9273);
or U15206 (N_15206,N_9822,N_9398);
xnor U15207 (N_15207,N_11904,N_10153);
nor U15208 (N_15208,N_8943,N_8540);
xor U15209 (N_15209,N_10741,N_8131);
xor U15210 (N_15210,N_8813,N_10026);
nand U15211 (N_15211,N_9727,N_11404);
nand U15212 (N_15212,N_11186,N_11803);
nor U15213 (N_15213,N_10814,N_8859);
and U15214 (N_15214,N_8691,N_10859);
or U15215 (N_15215,N_9240,N_11195);
or U15216 (N_15216,N_10710,N_8198);
nand U15217 (N_15217,N_8888,N_10999);
xor U15218 (N_15218,N_8580,N_8030);
xnor U15219 (N_15219,N_9440,N_8294);
and U15220 (N_15220,N_8963,N_10684);
nor U15221 (N_15221,N_11216,N_10604);
nor U15222 (N_15222,N_10935,N_8233);
or U15223 (N_15223,N_8893,N_9012);
nand U15224 (N_15224,N_8893,N_10573);
or U15225 (N_15225,N_10696,N_10655);
nand U15226 (N_15226,N_8625,N_9528);
and U15227 (N_15227,N_11075,N_10078);
or U15228 (N_15228,N_10766,N_11027);
xor U15229 (N_15229,N_10910,N_10721);
nor U15230 (N_15230,N_11144,N_11432);
nand U15231 (N_15231,N_11847,N_9932);
nand U15232 (N_15232,N_8376,N_8287);
and U15233 (N_15233,N_11015,N_9518);
nor U15234 (N_15234,N_8103,N_8842);
and U15235 (N_15235,N_11854,N_8279);
xor U15236 (N_15236,N_9538,N_11338);
nand U15237 (N_15237,N_11638,N_8113);
nor U15238 (N_15238,N_9586,N_11272);
and U15239 (N_15239,N_10945,N_10854);
and U15240 (N_15240,N_10870,N_10559);
xor U15241 (N_15241,N_9718,N_8156);
and U15242 (N_15242,N_11418,N_11687);
nor U15243 (N_15243,N_11394,N_10824);
or U15244 (N_15244,N_9908,N_11945);
nor U15245 (N_15245,N_10200,N_9719);
nand U15246 (N_15246,N_8499,N_9714);
nor U15247 (N_15247,N_11467,N_11202);
or U15248 (N_15248,N_10916,N_11326);
or U15249 (N_15249,N_10272,N_9099);
or U15250 (N_15250,N_9573,N_8077);
or U15251 (N_15251,N_11093,N_11756);
or U15252 (N_15252,N_11383,N_9752);
nor U15253 (N_15253,N_9428,N_8731);
or U15254 (N_15254,N_8988,N_8821);
nand U15255 (N_15255,N_8986,N_9339);
nor U15256 (N_15256,N_10813,N_9794);
xor U15257 (N_15257,N_10922,N_9648);
xnor U15258 (N_15258,N_10589,N_11004);
or U15259 (N_15259,N_9583,N_10888);
nand U15260 (N_15260,N_8760,N_9473);
and U15261 (N_15261,N_8527,N_8478);
and U15262 (N_15262,N_9767,N_10407);
nand U15263 (N_15263,N_10342,N_9696);
nor U15264 (N_15264,N_9421,N_11224);
or U15265 (N_15265,N_9281,N_11375);
or U15266 (N_15266,N_9103,N_8770);
nor U15267 (N_15267,N_11593,N_9840);
and U15268 (N_15268,N_11462,N_9009);
and U15269 (N_15269,N_8065,N_10241);
xor U15270 (N_15270,N_10490,N_11021);
and U15271 (N_15271,N_10025,N_11607);
or U15272 (N_15272,N_9002,N_11092);
nor U15273 (N_15273,N_11216,N_11964);
xnor U15274 (N_15274,N_8608,N_11843);
or U15275 (N_15275,N_11350,N_11185);
xnor U15276 (N_15276,N_11482,N_9894);
nand U15277 (N_15277,N_11738,N_8475);
and U15278 (N_15278,N_11321,N_10787);
or U15279 (N_15279,N_8608,N_9787);
nand U15280 (N_15280,N_8485,N_9210);
nand U15281 (N_15281,N_8557,N_8492);
nor U15282 (N_15282,N_10143,N_9206);
nor U15283 (N_15283,N_9539,N_9409);
xnor U15284 (N_15284,N_11300,N_11553);
or U15285 (N_15285,N_8986,N_11235);
and U15286 (N_15286,N_9845,N_10669);
nor U15287 (N_15287,N_11134,N_10576);
nor U15288 (N_15288,N_11134,N_8508);
nand U15289 (N_15289,N_8398,N_11116);
or U15290 (N_15290,N_9310,N_11441);
xor U15291 (N_15291,N_10402,N_8831);
nor U15292 (N_15292,N_8606,N_10873);
or U15293 (N_15293,N_9837,N_9462);
xnor U15294 (N_15294,N_10164,N_11072);
nand U15295 (N_15295,N_10320,N_9372);
nor U15296 (N_15296,N_9779,N_10213);
nand U15297 (N_15297,N_10623,N_10207);
and U15298 (N_15298,N_10706,N_9710);
nand U15299 (N_15299,N_9708,N_10467);
nor U15300 (N_15300,N_9261,N_9785);
or U15301 (N_15301,N_8499,N_9954);
xor U15302 (N_15302,N_9761,N_11246);
xnor U15303 (N_15303,N_10186,N_9844);
or U15304 (N_15304,N_8027,N_9735);
nor U15305 (N_15305,N_11648,N_8757);
and U15306 (N_15306,N_9474,N_11359);
xnor U15307 (N_15307,N_8336,N_10618);
nor U15308 (N_15308,N_10769,N_9360);
and U15309 (N_15309,N_8229,N_8499);
and U15310 (N_15310,N_9802,N_9364);
xnor U15311 (N_15311,N_8008,N_10855);
and U15312 (N_15312,N_11390,N_10462);
or U15313 (N_15313,N_8623,N_9609);
xor U15314 (N_15314,N_8678,N_8834);
or U15315 (N_15315,N_10922,N_8643);
or U15316 (N_15316,N_10401,N_11055);
nor U15317 (N_15317,N_11580,N_10303);
nor U15318 (N_15318,N_10254,N_11758);
nor U15319 (N_15319,N_8978,N_10183);
and U15320 (N_15320,N_8918,N_8991);
nor U15321 (N_15321,N_9539,N_8486);
or U15322 (N_15322,N_11127,N_9973);
and U15323 (N_15323,N_8331,N_10082);
nor U15324 (N_15324,N_8304,N_10459);
or U15325 (N_15325,N_9295,N_10214);
and U15326 (N_15326,N_9158,N_11334);
xor U15327 (N_15327,N_10708,N_10985);
and U15328 (N_15328,N_10018,N_9162);
xor U15329 (N_15329,N_10590,N_11421);
xor U15330 (N_15330,N_10127,N_9155);
or U15331 (N_15331,N_11186,N_9029);
nor U15332 (N_15332,N_11906,N_8169);
and U15333 (N_15333,N_11468,N_9036);
xnor U15334 (N_15334,N_9381,N_11880);
xnor U15335 (N_15335,N_9523,N_10991);
or U15336 (N_15336,N_10327,N_11646);
and U15337 (N_15337,N_10553,N_10818);
or U15338 (N_15338,N_8655,N_10279);
and U15339 (N_15339,N_9419,N_11839);
or U15340 (N_15340,N_9839,N_11625);
or U15341 (N_15341,N_10502,N_11990);
xor U15342 (N_15342,N_11229,N_10679);
or U15343 (N_15343,N_11272,N_8714);
nand U15344 (N_15344,N_8515,N_11530);
nor U15345 (N_15345,N_8823,N_10117);
or U15346 (N_15346,N_9025,N_11995);
nand U15347 (N_15347,N_11805,N_8386);
xnor U15348 (N_15348,N_8993,N_8064);
xor U15349 (N_15349,N_10406,N_11337);
and U15350 (N_15350,N_8922,N_9781);
and U15351 (N_15351,N_10379,N_10483);
or U15352 (N_15352,N_8937,N_11993);
nor U15353 (N_15353,N_8889,N_8412);
and U15354 (N_15354,N_10521,N_8020);
and U15355 (N_15355,N_8399,N_10611);
or U15356 (N_15356,N_9873,N_10180);
nand U15357 (N_15357,N_9172,N_10898);
and U15358 (N_15358,N_10399,N_11349);
xor U15359 (N_15359,N_9133,N_9503);
or U15360 (N_15360,N_8701,N_11791);
xor U15361 (N_15361,N_10028,N_10427);
and U15362 (N_15362,N_10343,N_10212);
xor U15363 (N_15363,N_11549,N_9300);
nor U15364 (N_15364,N_9538,N_11979);
xnor U15365 (N_15365,N_9897,N_9983);
nand U15366 (N_15366,N_9022,N_8849);
and U15367 (N_15367,N_9459,N_10556);
nor U15368 (N_15368,N_8014,N_11613);
and U15369 (N_15369,N_10136,N_8418);
or U15370 (N_15370,N_8934,N_10693);
nand U15371 (N_15371,N_9720,N_11138);
nand U15372 (N_15372,N_11581,N_8599);
and U15373 (N_15373,N_11031,N_8258);
nand U15374 (N_15374,N_9045,N_9916);
nand U15375 (N_15375,N_9772,N_8979);
xor U15376 (N_15376,N_11969,N_11489);
or U15377 (N_15377,N_8760,N_10379);
or U15378 (N_15378,N_8985,N_9256);
and U15379 (N_15379,N_11439,N_9233);
and U15380 (N_15380,N_8781,N_10962);
or U15381 (N_15381,N_9256,N_10539);
xor U15382 (N_15382,N_10931,N_8855);
and U15383 (N_15383,N_11389,N_9175);
and U15384 (N_15384,N_9076,N_8965);
xnor U15385 (N_15385,N_8194,N_10865);
or U15386 (N_15386,N_8541,N_8745);
nand U15387 (N_15387,N_10196,N_11785);
xnor U15388 (N_15388,N_10960,N_10202);
or U15389 (N_15389,N_9395,N_9513);
or U15390 (N_15390,N_10349,N_9638);
nand U15391 (N_15391,N_8889,N_11832);
nor U15392 (N_15392,N_10064,N_8093);
nand U15393 (N_15393,N_8145,N_11685);
or U15394 (N_15394,N_9372,N_8874);
and U15395 (N_15395,N_8687,N_8652);
nand U15396 (N_15396,N_9769,N_8391);
and U15397 (N_15397,N_11153,N_9170);
xnor U15398 (N_15398,N_10372,N_9514);
nand U15399 (N_15399,N_10833,N_8265);
xor U15400 (N_15400,N_10630,N_9842);
and U15401 (N_15401,N_10443,N_11831);
nor U15402 (N_15402,N_11415,N_9944);
xor U15403 (N_15403,N_10498,N_10416);
nor U15404 (N_15404,N_11898,N_8818);
nor U15405 (N_15405,N_8407,N_9557);
or U15406 (N_15406,N_9156,N_10044);
xnor U15407 (N_15407,N_8614,N_10682);
and U15408 (N_15408,N_9341,N_8692);
nand U15409 (N_15409,N_9282,N_11399);
nand U15410 (N_15410,N_10581,N_8447);
nand U15411 (N_15411,N_11404,N_8762);
nor U15412 (N_15412,N_8572,N_9040);
nor U15413 (N_15413,N_10831,N_9020);
nor U15414 (N_15414,N_9395,N_11461);
nand U15415 (N_15415,N_11995,N_11647);
nor U15416 (N_15416,N_10932,N_9815);
xnor U15417 (N_15417,N_8148,N_10185);
or U15418 (N_15418,N_10921,N_9787);
or U15419 (N_15419,N_11926,N_9360);
nor U15420 (N_15420,N_9012,N_8929);
and U15421 (N_15421,N_11604,N_8036);
nor U15422 (N_15422,N_8151,N_8204);
and U15423 (N_15423,N_8478,N_10396);
nor U15424 (N_15424,N_11701,N_9808);
or U15425 (N_15425,N_10088,N_10649);
and U15426 (N_15426,N_10163,N_8689);
or U15427 (N_15427,N_10038,N_9506);
xnor U15428 (N_15428,N_9524,N_10346);
or U15429 (N_15429,N_8221,N_11478);
xor U15430 (N_15430,N_10663,N_8544);
nand U15431 (N_15431,N_8043,N_9681);
xor U15432 (N_15432,N_9806,N_9988);
nor U15433 (N_15433,N_8507,N_9693);
and U15434 (N_15434,N_9700,N_10676);
nand U15435 (N_15435,N_9125,N_8375);
xor U15436 (N_15436,N_10018,N_10463);
nor U15437 (N_15437,N_8315,N_9218);
and U15438 (N_15438,N_9690,N_8851);
nor U15439 (N_15439,N_8072,N_8928);
xor U15440 (N_15440,N_10525,N_10347);
nand U15441 (N_15441,N_11970,N_11031);
and U15442 (N_15442,N_9144,N_9207);
nand U15443 (N_15443,N_8439,N_10391);
or U15444 (N_15444,N_8419,N_11063);
nor U15445 (N_15445,N_9942,N_8468);
and U15446 (N_15446,N_9533,N_11148);
and U15447 (N_15447,N_11782,N_8041);
nor U15448 (N_15448,N_9992,N_11262);
nand U15449 (N_15449,N_8733,N_11573);
xor U15450 (N_15450,N_9900,N_8462);
or U15451 (N_15451,N_9019,N_9113);
and U15452 (N_15452,N_10506,N_8798);
and U15453 (N_15453,N_11814,N_11600);
xor U15454 (N_15454,N_10145,N_9413);
or U15455 (N_15455,N_11954,N_8881);
and U15456 (N_15456,N_11047,N_11923);
nand U15457 (N_15457,N_9661,N_8488);
and U15458 (N_15458,N_8439,N_8507);
nand U15459 (N_15459,N_10644,N_10487);
and U15460 (N_15460,N_11685,N_11922);
or U15461 (N_15461,N_10534,N_11070);
nor U15462 (N_15462,N_10424,N_10490);
and U15463 (N_15463,N_11044,N_9594);
nand U15464 (N_15464,N_8304,N_9723);
nand U15465 (N_15465,N_11205,N_11382);
or U15466 (N_15466,N_10594,N_8420);
nand U15467 (N_15467,N_8359,N_10107);
xor U15468 (N_15468,N_9165,N_8049);
xor U15469 (N_15469,N_8127,N_10534);
or U15470 (N_15470,N_8622,N_10212);
and U15471 (N_15471,N_10359,N_10813);
and U15472 (N_15472,N_8911,N_10188);
nand U15473 (N_15473,N_11305,N_9618);
nand U15474 (N_15474,N_11911,N_10243);
and U15475 (N_15475,N_11971,N_11319);
and U15476 (N_15476,N_9760,N_11601);
or U15477 (N_15477,N_11834,N_11801);
nor U15478 (N_15478,N_11929,N_9995);
xor U15479 (N_15479,N_8235,N_9781);
or U15480 (N_15480,N_9826,N_11728);
nor U15481 (N_15481,N_9219,N_8704);
nand U15482 (N_15482,N_11797,N_10485);
xor U15483 (N_15483,N_11117,N_9298);
nand U15484 (N_15484,N_10145,N_10349);
nand U15485 (N_15485,N_9277,N_9041);
xor U15486 (N_15486,N_8249,N_8916);
nor U15487 (N_15487,N_9780,N_9571);
or U15488 (N_15488,N_10002,N_11909);
nor U15489 (N_15489,N_9348,N_9007);
nand U15490 (N_15490,N_11802,N_8002);
nand U15491 (N_15491,N_11394,N_9044);
xnor U15492 (N_15492,N_11284,N_8991);
xnor U15493 (N_15493,N_10099,N_8205);
nand U15494 (N_15494,N_11279,N_11568);
nand U15495 (N_15495,N_10076,N_11322);
nand U15496 (N_15496,N_11001,N_9472);
xnor U15497 (N_15497,N_8256,N_9696);
or U15498 (N_15498,N_9049,N_8460);
nor U15499 (N_15499,N_11597,N_11804);
nand U15500 (N_15500,N_8557,N_8635);
nand U15501 (N_15501,N_9827,N_8855);
nand U15502 (N_15502,N_10921,N_8435);
nand U15503 (N_15503,N_9061,N_10940);
xor U15504 (N_15504,N_9390,N_9623);
nor U15505 (N_15505,N_10966,N_9019);
or U15506 (N_15506,N_10031,N_8881);
xnor U15507 (N_15507,N_11253,N_8318);
nor U15508 (N_15508,N_10923,N_9759);
or U15509 (N_15509,N_10010,N_8821);
nor U15510 (N_15510,N_11639,N_11569);
xor U15511 (N_15511,N_8954,N_10811);
xor U15512 (N_15512,N_8460,N_8262);
or U15513 (N_15513,N_11211,N_10351);
nand U15514 (N_15514,N_8034,N_10530);
xnor U15515 (N_15515,N_10078,N_9007);
nand U15516 (N_15516,N_10094,N_8247);
nor U15517 (N_15517,N_9883,N_10001);
or U15518 (N_15518,N_11218,N_9804);
and U15519 (N_15519,N_10439,N_11922);
xnor U15520 (N_15520,N_10865,N_9480);
nor U15521 (N_15521,N_9353,N_9527);
or U15522 (N_15522,N_11909,N_8349);
xnor U15523 (N_15523,N_10625,N_11374);
nor U15524 (N_15524,N_11386,N_11589);
and U15525 (N_15525,N_11496,N_11293);
nor U15526 (N_15526,N_11960,N_9519);
nand U15527 (N_15527,N_9784,N_8797);
and U15528 (N_15528,N_9715,N_9309);
nand U15529 (N_15529,N_8009,N_8997);
and U15530 (N_15530,N_11146,N_10216);
nand U15531 (N_15531,N_9007,N_10839);
and U15532 (N_15532,N_11325,N_9643);
nor U15533 (N_15533,N_9534,N_11255);
nor U15534 (N_15534,N_9615,N_9601);
or U15535 (N_15535,N_9994,N_9212);
xor U15536 (N_15536,N_11133,N_9073);
or U15537 (N_15537,N_9594,N_9194);
and U15538 (N_15538,N_9890,N_8236);
and U15539 (N_15539,N_9835,N_9997);
xor U15540 (N_15540,N_9945,N_11090);
and U15541 (N_15541,N_10192,N_8899);
and U15542 (N_15542,N_9600,N_11842);
nor U15543 (N_15543,N_10754,N_10705);
xnor U15544 (N_15544,N_11217,N_10133);
or U15545 (N_15545,N_9566,N_11816);
xnor U15546 (N_15546,N_11425,N_10497);
xnor U15547 (N_15547,N_8414,N_9804);
nand U15548 (N_15548,N_9269,N_10853);
nand U15549 (N_15549,N_8154,N_11203);
nor U15550 (N_15550,N_8795,N_8215);
or U15551 (N_15551,N_10891,N_10093);
nor U15552 (N_15552,N_10705,N_11779);
nor U15553 (N_15553,N_10319,N_11646);
nor U15554 (N_15554,N_11972,N_9814);
nand U15555 (N_15555,N_10607,N_9849);
or U15556 (N_15556,N_10305,N_11492);
nor U15557 (N_15557,N_8646,N_11037);
xor U15558 (N_15558,N_9547,N_8885);
nor U15559 (N_15559,N_8186,N_10902);
or U15560 (N_15560,N_10337,N_11325);
nor U15561 (N_15561,N_11230,N_11929);
nand U15562 (N_15562,N_10870,N_8990);
nor U15563 (N_15563,N_10828,N_11617);
and U15564 (N_15564,N_10632,N_11887);
nand U15565 (N_15565,N_9318,N_9438);
nor U15566 (N_15566,N_10225,N_10932);
xnor U15567 (N_15567,N_11013,N_9197);
nand U15568 (N_15568,N_10716,N_11129);
and U15569 (N_15569,N_11045,N_10206);
xnor U15570 (N_15570,N_9466,N_10399);
or U15571 (N_15571,N_10326,N_11237);
nand U15572 (N_15572,N_9428,N_9559);
nor U15573 (N_15573,N_10766,N_10971);
xor U15574 (N_15574,N_9248,N_8028);
nand U15575 (N_15575,N_8049,N_9665);
nand U15576 (N_15576,N_8278,N_9100);
and U15577 (N_15577,N_10597,N_9095);
nand U15578 (N_15578,N_10628,N_10019);
or U15579 (N_15579,N_11119,N_8927);
and U15580 (N_15580,N_10274,N_9730);
nand U15581 (N_15581,N_8070,N_11063);
and U15582 (N_15582,N_11565,N_8314);
and U15583 (N_15583,N_9170,N_10345);
nor U15584 (N_15584,N_10092,N_10706);
or U15585 (N_15585,N_11129,N_10953);
and U15586 (N_15586,N_11723,N_10607);
nor U15587 (N_15587,N_10538,N_9113);
nand U15588 (N_15588,N_10861,N_8758);
nor U15589 (N_15589,N_10492,N_10760);
nor U15590 (N_15590,N_11512,N_8485);
or U15591 (N_15591,N_9740,N_11425);
xor U15592 (N_15592,N_9204,N_9042);
nor U15593 (N_15593,N_11297,N_9479);
xor U15594 (N_15594,N_8334,N_10345);
nand U15595 (N_15595,N_9008,N_11130);
xor U15596 (N_15596,N_11384,N_10788);
nor U15597 (N_15597,N_11825,N_11419);
and U15598 (N_15598,N_8685,N_10729);
and U15599 (N_15599,N_10244,N_11763);
nand U15600 (N_15600,N_8820,N_11606);
xor U15601 (N_15601,N_8616,N_11200);
and U15602 (N_15602,N_9185,N_8377);
nor U15603 (N_15603,N_11513,N_10276);
xor U15604 (N_15604,N_11152,N_11393);
nand U15605 (N_15605,N_10455,N_8203);
xor U15606 (N_15606,N_9747,N_10582);
nor U15607 (N_15607,N_10909,N_9275);
or U15608 (N_15608,N_8341,N_8255);
nand U15609 (N_15609,N_10706,N_11500);
or U15610 (N_15610,N_9885,N_9341);
and U15611 (N_15611,N_9068,N_10876);
or U15612 (N_15612,N_9263,N_11207);
or U15613 (N_15613,N_10027,N_9628);
nor U15614 (N_15614,N_10100,N_11120);
xnor U15615 (N_15615,N_9177,N_8650);
or U15616 (N_15616,N_10690,N_8911);
and U15617 (N_15617,N_11589,N_8505);
nor U15618 (N_15618,N_10750,N_10446);
nor U15619 (N_15619,N_8323,N_11744);
nand U15620 (N_15620,N_11564,N_8029);
or U15621 (N_15621,N_8407,N_11520);
nor U15622 (N_15622,N_9232,N_9463);
nor U15623 (N_15623,N_11623,N_10703);
nor U15624 (N_15624,N_9137,N_8073);
or U15625 (N_15625,N_11668,N_10118);
xnor U15626 (N_15626,N_10919,N_11677);
xor U15627 (N_15627,N_11283,N_10966);
and U15628 (N_15628,N_8249,N_10595);
and U15629 (N_15629,N_11635,N_11496);
nor U15630 (N_15630,N_9379,N_11055);
or U15631 (N_15631,N_11966,N_11207);
nor U15632 (N_15632,N_11114,N_11069);
and U15633 (N_15633,N_8974,N_9966);
nand U15634 (N_15634,N_11665,N_9286);
and U15635 (N_15635,N_9804,N_8640);
or U15636 (N_15636,N_8947,N_11831);
nor U15637 (N_15637,N_9276,N_11054);
xnor U15638 (N_15638,N_9358,N_10687);
xor U15639 (N_15639,N_8819,N_10956);
nand U15640 (N_15640,N_9786,N_11603);
nor U15641 (N_15641,N_10041,N_8040);
or U15642 (N_15642,N_11265,N_11207);
or U15643 (N_15643,N_11987,N_11656);
nor U15644 (N_15644,N_11358,N_9803);
xor U15645 (N_15645,N_9266,N_11485);
nand U15646 (N_15646,N_10066,N_8529);
nor U15647 (N_15647,N_10600,N_9195);
xor U15648 (N_15648,N_9378,N_11504);
or U15649 (N_15649,N_8817,N_8367);
or U15650 (N_15650,N_8495,N_11140);
nor U15651 (N_15651,N_8011,N_9674);
nor U15652 (N_15652,N_11834,N_9850);
or U15653 (N_15653,N_11855,N_8193);
nand U15654 (N_15654,N_8241,N_8469);
or U15655 (N_15655,N_8921,N_11058);
nor U15656 (N_15656,N_9707,N_11523);
or U15657 (N_15657,N_8599,N_8094);
and U15658 (N_15658,N_8359,N_9905);
nand U15659 (N_15659,N_11462,N_8695);
xnor U15660 (N_15660,N_10854,N_9180);
xor U15661 (N_15661,N_11286,N_10980);
nor U15662 (N_15662,N_9851,N_11509);
nand U15663 (N_15663,N_9420,N_9096);
and U15664 (N_15664,N_11577,N_8694);
nand U15665 (N_15665,N_10835,N_11814);
and U15666 (N_15666,N_11536,N_8034);
nor U15667 (N_15667,N_9356,N_9429);
nor U15668 (N_15668,N_9471,N_9597);
and U15669 (N_15669,N_10120,N_9835);
nand U15670 (N_15670,N_8609,N_9880);
and U15671 (N_15671,N_10007,N_10181);
or U15672 (N_15672,N_8131,N_10763);
and U15673 (N_15673,N_10265,N_11852);
nand U15674 (N_15674,N_11790,N_9240);
and U15675 (N_15675,N_11657,N_10910);
nor U15676 (N_15676,N_9573,N_11531);
and U15677 (N_15677,N_10115,N_8814);
or U15678 (N_15678,N_9513,N_8187);
xnor U15679 (N_15679,N_11118,N_11242);
nor U15680 (N_15680,N_8187,N_9087);
xor U15681 (N_15681,N_11415,N_10371);
xnor U15682 (N_15682,N_8501,N_9807);
nor U15683 (N_15683,N_11068,N_8895);
nand U15684 (N_15684,N_10799,N_10682);
xor U15685 (N_15685,N_10805,N_9907);
or U15686 (N_15686,N_9044,N_8571);
and U15687 (N_15687,N_8532,N_10330);
nand U15688 (N_15688,N_11351,N_8547);
nor U15689 (N_15689,N_8983,N_10252);
xnor U15690 (N_15690,N_10403,N_11727);
nor U15691 (N_15691,N_9870,N_8394);
xor U15692 (N_15692,N_11040,N_11848);
or U15693 (N_15693,N_10583,N_8343);
xnor U15694 (N_15694,N_8156,N_10641);
nand U15695 (N_15695,N_10598,N_11216);
nor U15696 (N_15696,N_11747,N_11135);
nand U15697 (N_15697,N_9598,N_11120);
and U15698 (N_15698,N_8411,N_10201);
and U15699 (N_15699,N_9415,N_9213);
and U15700 (N_15700,N_10592,N_8331);
nor U15701 (N_15701,N_11778,N_8215);
nand U15702 (N_15702,N_11534,N_10638);
nor U15703 (N_15703,N_8662,N_9155);
and U15704 (N_15704,N_11309,N_11195);
nand U15705 (N_15705,N_9223,N_10970);
and U15706 (N_15706,N_9247,N_10112);
nor U15707 (N_15707,N_10527,N_11104);
nor U15708 (N_15708,N_9004,N_11070);
xnor U15709 (N_15709,N_11406,N_10272);
or U15710 (N_15710,N_10680,N_9134);
nor U15711 (N_15711,N_8039,N_11822);
or U15712 (N_15712,N_11775,N_9377);
nor U15713 (N_15713,N_8725,N_10365);
or U15714 (N_15714,N_10646,N_8936);
or U15715 (N_15715,N_10707,N_9316);
nand U15716 (N_15716,N_8671,N_8177);
or U15717 (N_15717,N_9765,N_11016);
nor U15718 (N_15718,N_8191,N_10283);
nor U15719 (N_15719,N_11264,N_9535);
nor U15720 (N_15720,N_10736,N_11954);
nor U15721 (N_15721,N_8509,N_8737);
or U15722 (N_15722,N_10707,N_11365);
or U15723 (N_15723,N_11567,N_10057);
nor U15724 (N_15724,N_10771,N_10767);
and U15725 (N_15725,N_9437,N_11242);
xor U15726 (N_15726,N_11874,N_8227);
and U15727 (N_15727,N_8365,N_8498);
nor U15728 (N_15728,N_11988,N_8213);
nand U15729 (N_15729,N_11226,N_9172);
nor U15730 (N_15730,N_11902,N_11710);
or U15731 (N_15731,N_10684,N_9272);
nand U15732 (N_15732,N_9533,N_10364);
and U15733 (N_15733,N_11542,N_10730);
xnor U15734 (N_15734,N_11288,N_9141);
or U15735 (N_15735,N_8057,N_8491);
xor U15736 (N_15736,N_10900,N_10694);
nand U15737 (N_15737,N_11640,N_8584);
or U15738 (N_15738,N_11792,N_11232);
and U15739 (N_15739,N_8103,N_9874);
or U15740 (N_15740,N_8799,N_11664);
nand U15741 (N_15741,N_9581,N_8872);
or U15742 (N_15742,N_10905,N_9397);
xor U15743 (N_15743,N_10334,N_9193);
and U15744 (N_15744,N_11690,N_8270);
nor U15745 (N_15745,N_9752,N_10420);
nand U15746 (N_15746,N_8055,N_10676);
nand U15747 (N_15747,N_11727,N_8864);
and U15748 (N_15748,N_9996,N_11932);
nor U15749 (N_15749,N_8291,N_8694);
nor U15750 (N_15750,N_9061,N_8160);
nand U15751 (N_15751,N_11313,N_10632);
and U15752 (N_15752,N_9984,N_9039);
nand U15753 (N_15753,N_9989,N_10175);
or U15754 (N_15754,N_9338,N_11400);
and U15755 (N_15755,N_9662,N_8754);
nor U15756 (N_15756,N_8146,N_8168);
xor U15757 (N_15757,N_8039,N_8886);
and U15758 (N_15758,N_9902,N_11944);
nor U15759 (N_15759,N_8611,N_10480);
nor U15760 (N_15760,N_10903,N_8668);
nor U15761 (N_15761,N_8360,N_11664);
nor U15762 (N_15762,N_10220,N_8418);
or U15763 (N_15763,N_8928,N_8506);
or U15764 (N_15764,N_9290,N_11524);
and U15765 (N_15765,N_9405,N_11430);
and U15766 (N_15766,N_10002,N_11415);
nand U15767 (N_15767,N_11772,N_10430);
or U15768 (N_15768,N_10762,N_9600);
and U15769 (N_15769,N_9156,N_10170);
or U15770 (N_15770,N_11202,N_11955);
and U15771 (N_15771,N_11900,N_9691);
xor U15772 (N_15772,N_10033,N_8952);
or U15773 (N_15773,N_9341,N_9415);
xor U15774 (N_15774,N_8573,N_11951);
nand U15775 (N_15775,N_11416,N_11654);
or U15776 (N_15776,N_10039,N_8091);
and U15777 (N_15777,N_8615,N_9113);
nor U15778 (N_15778,N_9882,N_11432);
or U15779 (N_15779,N_10067,N_8865);
xnor U15780 (N_15780,N_10063,N_11460);
or U15781 (N_15781,N_11332,N_9250);
nand U15782 (N_15782,N_8083,N_8927);
and U15783 (N_15783,N_8526,N_9046);
nand U15784 (N_15784,N_11458,N_11567);
xnor U15785 (N_15785,N_11292,N_10768);
xor U15786 (N_15786,N_10025,N_10518);
or U15787 (N_15787,N_8506,N_9925);
xnor U15788 (N_15788,N_9472,N_10162);
and U15789 (N_15789,N_11446,N_11541);
xnor U15790 (N_15790,N_8652,N_10820);
nor U15791 (N_15791,N_10277,N_11442);
nand U15792 (N_15792,N_10368,N_11133);
xor U15793 (N_15793,N_10057,N_9367);
xor U15794 (N_15794,N_10751,N_11927);
or U15795 (N_15795,N_8254,N_8642);
nor U15796 (N_15796,N_8052,N_8111);
nand U15797 (N_15797,N_11246,N_10167);
nand U15798 (N_15798,N_8093,N_10870);
xor U15799 (N_15799,N_10183,N_9469);
and U15800 (N_15800,N_10417,N_11489);
nand U15801 (N_15801,N_11099,N_8110);
nand U15802 (N_15802,N_11167,N_10989);
nor U15803 (N_15803,N_9619,N_8409);
or U15804 (N_15804,N_9261,N_10890);
or U15805 (N_15805,N_11459,N_11631);
xor U15806 (N_15806,N_9243,N_10827);
nor U15807 (N_15807,N_11474,N_10197);
nor U15808 (N_15808,N_9033,N_9161);
or U15809 (N_15809,N_9928,N_9495);
and U15810 (N_15810,N_8044,N_9296);
and U15811 (N_15811,N_8834,N_11330);
or U15812 (N_15812,N_11845,N_8955);
nor U15813 (N_15813,N_10417,N_11445);
or U15814 (N_15814,N_10786,N_9209);
nand U15815 (N_15815,N_10514,N_9232);
xor U15816 (N_15816,N_10145,N_9055);
and U15817 (N_15817,N_8749,N_8468);
xor U15818 (N_15818,N_9448,N_9721);
nor U15819 (N_15819,N_10543,N_10981);
or U15820 (N_15820,N_11243,N_8098);
nand U15821 (N_15821,N_9130,N_10084);
xnor U15822 (N_15822,N_8341,N_11850);
nor U15823 (N_15823,N_11677,N_9004);
and U15824 (N_15824,N_11522,N_9432);
nand U15825 (N_15825,N_8158,N_11262);
nor U15826 (N_15826,N_11092,N_8155);
or U15827 (N_15827,N_11787,N_11986);
xnor U15828 (N_15828,N_10134,N_9610);
xnor U15829 (N_15829,N_8294,N_9182);
nor U15830 (N_15830,N_8042,N_9605);
nand U15831 (N_15831,N_11619,N_8717);
and U15832 (N_15832,N_8649,N_9675);
or U15833 (N_15833,N_9104,N_11214);
nor U15834 (N_15834,N_8173,N_10359);
nor U15835 (N_15835,N_11339,N_10946);
xor U15836 (N_15836,N_8608,N_9366);
nor U15837 (N_15837,N_9134,N_9524);
nor U15838 (N_15838,N_11423,N_9094);
and U15839 (N_15839,N_11137,N_10531);
or U15840 (N_15840,N_8456,N_9196);
and U15841 (N_15841,N_8706,N_8628);
xor U15842 (N_15842,N_9400,N_8053);
nand U15843 (N_15843,N_8793,N_9467);
nand U15844 (N_15844,N_9692,N_11734);
xnor U15845 (N_15845,N_10878,N_11991);
nand U15846 (N_15846,N_11571,N_11051);
and U15847 (N_15847,N_11582,N_10732);
nor U15848 (N_15848,N_10341,N_11060);
xor U15849 (N_15849,N_11227,N_9978);
and U15850 (N_15850,N_8396,N_11726);
nor U15851 (N_15851,N_10300,N_8466);
nor U15852 (N_15852,N_8617,N_8988);
or U15853 (N_15853,N_9094,N_8372);
or U15854 (N_15854,N_9840,N_11359);
xor U15855 (N_15855,N_8980,N_9187);
or U15856 (N_15856,N_9735,N_10940);
or U15857 (N_15857,N_9374,N_11207);
and U15858 (N_15858,N_10386,N_10466);
nor U15859 (N_15859,N_10892,N_8506);
xor U15860 (N_15860,N_10014,N_11995);
xnor U15861 (N_15861,N_11649,N_11964);
nand U15862 (N_15862,N_9067,N_10811);
nand U15863 (N_15863,N_10747,N_8988);
xor U15864 (N_15864,N_11199,N_10125);
xnor U15865 (N_15865,N_8963,N_8018);
and U15866 (N_15866,N_10794,N_8478);
or U15867 (N_15867,N_8671,N_10382);
and U15868 (N_15868,N_11954,N_10909);
and U15869 (N_15869,N_9567,N_11532);
nand U15870 (N_15870,N_9514,N_11915);
nand U15871 (N_15871,N_9794,N_9947);
nand U15872 (N_15872,N_9289,N_8044);
and U15873 (N_15873,N_10653,N_10918);
nor U15874 (N_15874,N_9269,N_10494);
nand U15875 (N_15875,N_9942,N_11907);
xnor U15876 (N_15876,N_11037,N_8652);
or U15877 (N_15877,N_9289,N_10026);
or U15878 (N_15878,N_11990,N_8888);
nand U15879 (N_15879,N_11487,N_11331);
or U15880 (N_15880,N_10929,N_10369);
or U15881 (N_15881,N_8402,N_10852);
and U15882 (N_15882,N_9174,N_11233);
nand U15883 (N_15883,N_10656,N_11546);
xor U15884 (N_15884,N_8393,N_11903);
and U15885 (N_15885,N_8480,N_9605);
nor U15886 (N_15886,N_10277,N_10065);
xor U15887 (N_15887,N_8016,N_8953);
nor U15888 (N_15888,N_10868,N_10933);
and U15889 (N_15889,N_11571,N_10768);
nor U15890 (N_15890,N_8118,N_11254);
nor U15891 (N_15891,N_8251,N_9440);
or U15892 (N_15892,N_9045,N_8657);
nand U15893 (N_15893,N_11041,N_9757);
or U15894 (N_15894,N_10942,N_11211);
nor U15895 (N_15895,N_11397,N_9426);
or U15896 (N_15896,N_10020,N_9959);
nor U15897 (N_15897,N_11983,N_9275);
nor U15898 (N_15898,N_9535,N_11935);
nand U15899 (N_15899,N_8999,N_8107);
xor U15900 (N_15900,N_10346,N_9247);
nand U15901 (N_15901,N_11581,N_8066);
and U15902 (N_15902,N_10810,N_11505);
nand U15903 (N_15903,N_8050,N_8080);
or U15904 (N_15904,N_11477,N_10668);
nor U15905 (N_15905,N_10926,N_8256);
nand U15906 (N_15906,N_8990,N_9452);
nor U15907 (N_15907,N_9154,N_11557);
xnor U15908 (N_15908,N_11564,N_9898);
or U15909 (N_15909,N_9987,N_10014);
xor U15910 (N_15910,N_10741,N_11158);
xor U15911 (N_15911,N_8075,N_10289);
or U15912 (N_15912,N_9161,N_11749);
or U15913 (N_15913,N_10267,N_10023);
and U15914 (N_15914,N_10865,N_10642);
nand U15915 (N_15915,N_9172,N_8504);
nand U15916 (N_15916,N_9978,N_8100);
and U15917 (N_15917,N_10982,N_8221);
and U15918 (N_15918,N_9390,N_10747);
nor U15919 (N_15919,N_11114,N_11231);
xnor U15920 (N_15920,N_10340,N_10920);
nor U15921 (N_15921,N_10047,N_9859);
nor U15922 (N_15922,N_10678,N_10052);
or U15923 (N_15923,N_10268,N_8136);
or U15924 (N_15924,N_10785,N_9522);
nand U15925 (N_15925,N_8969,N_8317);
and U15926 (N_15926,N_11606,N_10830);
or U15927 (N_15927,N_9059,N_10090);
nor U15928 (N_15928,N_8212,N_11449);
xor U15929 (N_15929,N_9958,N_11396);
xor U15930 (N_15930,N_8816,N_10540);
or U15931 (N_15931,N_11364,N_9371);
nand U15932 (N_15932,N_8876,N_11365);
nand U15933 (N_15933,N_11235,N_10022);
or U15934 (N_15934,N_8097,N_8129);
and U15935 (N_15935,N_11610,N_10723);
and U15936 (N_15936,N_11210,N_10267);
nor U15937 (N_15937,N_9137,N_10116);
nor U15938 (N_15938,N_10597,N_10466);
nand U15939 (N_15939,N_11684,N_9721);
or U15940 (N_15940,N_11564,N_8488);
or U15941 (N_15941,N_8994,N_8344);
or U15942 (N_15942,N_11041,N_11928);
nand U15943 (N_15943,N_10844,N_9784);
or U15944 (N_15944,N_8524,N_8320);
nand U15945 (N_15945,N_10115,N_11218);
and U15946 (N_15946,N_9231,N_10877);
and U15947 (N_15947,N_11342,N_8990);
xor U15948 (N_15948,N_10780,N_9414);
or U15949 (N_15949,N_8775,N_11945);
and U15950 (N_15950,N_9787,N_11930);
nor U15951 (N_15951,N_11213,N_9970);
nand U15952 (N_15952,N_8812,N_8095);
and U15953 (N_15953,N_9613,N_11635);
and U15954 (N_15954,N_11129,N_11127);
or U15955 (N_15955,N_8509,N_9123);
xnor U15956 (N_15956,N_8377,N_9839);
xor U15957 (N_15957,N_10444,N_10624);
xnor U15958 (N_15958,N_9340,N_8980);
xor U15959 (N_15959,N_10252,N_9624);
and U15960 (N_15960,N_10866,N_10555);
and U15961 (N_15961,N_11683,N_10862);
and U15962 (N_15962,N_11473,N_9831);
nand U15963 (N_15963,N_11023,N_11212);
and U15964 (N_15964,N_8037,N_8509);
nand U15965 (N_15965,N_10774,N_8528);
xor U15966 (N_15966,N_9737,N_8012);
nand U15967 (N_15967,N_11267,N_10852);
or U15968 (N_15968,N_10115,N_9019);
and U15969 (N_15969,N_8614,N_9151);
nor U15970 (N_15970,N_10768,N_10377);
nor U15971 (N_15971,N_9690,N_11805);
xnor U15972 (N_15972,N_8988,N_8712);
nor U15973 (N_15973,N_9546,N_8208);
nand U15974 (N_15974,N_11971,N_11882);
nand U15975 (N_15975,N_9336,N_9273);
nand U15976 (N_15976,N_11561,N_10843);
or U15977 (N_15977,N_8428,N_8982);
or U15978 (N_15978,N_11948,N_8518);
or U15979 (N_15979,N_8621,N_9305);
nor U15980 (N_15980,N_8018,N_11827);
and U15981 (N_15981,N_8022,N_8058);
nand U15982 (N_15982,N_8178,N_9673);
xor U15983 (N_15983,N_10279,N_9193);
or U15984 (N_15984,N_11630,N_8825);
and U15985 (N_15985,N_9610,N_11032);
nor U15986 (N_15986,N_11378,N_10913);
or U15987 (N_15987,N_10457,N_9132);
nand U15988 (N_15988,N_9527,N_11352);
nor U15989 (N_15989,N_10039,N_8528);
or U15990 (N_15990,N_10811,N_8885);
nor U15991 (N_15991,N_11791,N_8812);
and U15992 (N_15992,N_11337,N_10578);
xnor U15993 (N_15993,N_10172,N_10108);
and U15994 (N_15994,N_9438,N_8763);
or U15995 (N_15995,N_10537,N_10690);
xnor U15996 (N_15996,N_10919,N_11583);
and U15997 (N_15997,N_10788,N_10202);
xnor U15998 (N_15998,N_11430,N_10815);
or U15999 (N_15999,N_11893,N_8029);
or U16000 (N_16000,N_15930,N_13934);
nand U16001 (N_16001,N_12012,N_15753);
nand U16002 (N_16002,N_13646,N_15658);
nor U16003 (N_16003,N_12521,N_12390);
xor U16004 (N_16004,N_14259,N_12410);
nand U16005 (N_16005,N_14364,N_14699);
nor U16006 (N_16006,N_14762,N_15585);
nand U16007 (N_16007,N_14168,N_12797);
nor U16008 (N_16008,N_15641,N_12080);
nand U16009 (N_16009,N_15375,N_14972);
nand U16010 (N_16010,N_12174,N_15098);
and U16011 (N_16011,N_13165,N_14841);
xor U16012 (N_16012,N_14155,N_12468);
nor U16013 (N_16013,N_14409,N_14653);
xor U16014 (N_16014,N_12846,N_14974);
and U16015 (N_16015,N_15061,N_14264);
xnor U16016 (N_16016,N_12767,N_12498);
or U16017 (N_16017,N_14115,N_15947);
nor U16018 (N_16018,N_13027,N_12708);
nand U16019 (N_16019,N_14060,N_13502);
xnor U16020 (N_16020,N_12199,N_14515);
and U16021 (N_16021,N_14290,N_15144);
nand U16022 (N_16022,N_12799,N_15737);
xor U16023 (N_16023,N_12462,N_13058);
xnor U16024 (N_16024,N_12447,N_13788);
or U16025 (N_16025,N_13952,N_14840);
or U16026 (N_16026,N_14575,N_13471);
or U16027 (N_16027,N_14059,N_15519);
and U16028 (N_16028,N_12133,N_12152);
or U16029 (N_16029,N_13946,N_15323);
xnor U16030 (N_16030,N_12860,N_14689);
nand U16031 (N_16031,N_13481,N_12650);
or U16032 (N_16032,N_15435,N_12611);
xnor U16033 (N_16033,N_13314,N_15655);
and U16034 (N_16034,N_15589,N_12440);
and U16035 (N_16035,N_14873,N_13324);
nand U16036 (N_16036,N_12814,N_14539);
nand U16037 (N_16037,N_12908,N_13746);
nor U16038 (N_16038,N_14952,N_12657);
xnor U16039 (N_16039,N_12584,N_14506);
or U16040 (N_16040,N_14799,N_12942);
nor U16041 (N_16041,N_12121,N_15887);
or U16042 (N_16042,N_12671,N_15332);
nand U16043 (N_16043,N_14696,N_13288);
nor U16044 (N_16044,N_13115,N_14651);
or U16045 (N_16045,N_15401,N_15719);
nor U16046 (N_16046,N_12522,N_13967);
nor U16047 (N_16047,N_13672,N_12388);
nand U16048 (N_16048,N_13511,N_12513);
nand U16049 (N_16049,N_13100,N_14742);
nor U16050 (N_16050,N_13979,N_14177);
nor U16051 (N_16051,N_15409,N_12361);
xnor U16052 (N_16052,N_13220,N_15911);
nor U16053 (N_16053,N_13197,N_12758);
nand U16054 (N_16054,N_13602,N_13120);
nor U16055 (N_16055,N_14455,N_14489);
xor U16056 (N_16056,N_13011,N_13173);
xnor U16057 (N_16057,N_14353,N_15682);
or U16058 (N_16058,N_12682,N_13548);
nand U16059 (N_16059,N_13902,N_12897);
or U16060 (N_16060,N_14606,N_14114);
nand U16061 (N_16061,N_14293,N_15021);
xnor U16062 (N_16062,N_15559,N_13087);
xnor U16063 (N_16063,N_14861,N_12138);
nand U16064 (N_16064,N_14138,N_12986);
and U16065 (N_16065,N_13241,N_12808);
nand U16066 (N_16066,N_13963,N_14054);
and U16067 (N_16067,N_14932,N_13924);
and U16068 (N_16068,N_15917,N_15527);
and U16069 (N_16069,N_13785,N_12620);
xnor U16070 (N_16070,N_15076,N_12204);
nor U16071 (N_16071,N_15613,N_13650);
xnor U16072 (N_16072,N_15333,N_12379);
or U16073 (N_16073,N_14969,N_14746);
or U16074 (N_16074,N_13641,N_15366);
or U16075 (N_16075,N_13154,N_13781);
nand U16076 (N_16076,N_14786,N_13413);
nor U16077 (N_16077,N_15568,N_12987);
nand U16078 (N_16078,N_15827,N_15405);
and U16079 (N_16079,N_12068,N_12932);
nand U16080 (N_16080,N_13257,N_12725);
nand U16081 (N_16081,N_13069,N_13316);
and U16082 (N_16082,N_12069,N_13072);
nor U16083 (N_16083,N_13245,N_14686);
and U16084 (N_16084,N_15634,N_13224);
nand U16085 (N_16085,N_12426,N_14899);
and U16086 (N_16086,N_14436,N_13732);
and U16087 (N_16087,N_12718,N_15311);
nand U16088 (N_16088,N_13276,N_14169);
nand U16089 (N_16089,N_14101,N_15006);
xor U16090 (N_16090,N_12348,N_14791);
or U16091 (N_16091,N_15876,N_13848);
nand U16092 (N_16092,N_12867,N_15270);
xnor U16093 (N_16093,N_12691,N_14732);
and U16094 (N_16094,N_15805,N_13039);
xor U16095 (N_16095,N_13983,N_15328);
or U16096 (N_16096,N_14819,N_12640);
nand U16097 (N_16097,N_12639,N_14850);
nand U16098 (N_16098,N_15550,N_14597);
or U16099 (N_16099,N_12531,N_15709);
nor U16100 (N_16100,N_12707,N_15581);
nor U16101 (N_16101,N_12997,N_15046);
nand U16102 (N_16102,N_13139,N_15319);
nor U16103 (N_16103,N_13681,N_15960);
xnor U16104 (N_16104,N_13201,N_13737);
or U16105 (N_16105,N_12283,N_13371);
and U16106 (N_16106,N_12917,N_15592);
or U16107 (N_16107,N_15135,N_15163);
xnor U16108 (N_16108,N_14621,N_15958);
and U16109 (N_16109,N_12876,N_14598);
xor U16110 (N_16110,N_13459,N_12234);
nand U16111 (N_16111,N_14967,N_15809);
nor U16112 (N_16112,N_15793,N_13195);
and U16113 (N_16113,N_15150,N_14628);
nand U16114 (N_16114,N_15434,N_13327);
nand U16115 (N_16115,N_13700,N_13190);
or U16116 (N_16116,N_12652,N_15016);
or U16117 (N_16117,N_14717,N_12926);
xnor U16118 (N_16118,N_13347,N_12212);
nor U16119 (N_16119,N_14381,N_12399);
or U16120 (N_16120,N_12466,N_14073);
nand U16121 (N_16121,N_14363,N_14831);
nor U16122 (N_16122,N_15729,N_15885);
nor U16123 (N_16123,N_15059,N_12765);
nand U16124 (N_16124,N_12084,N_14801);
nand U16125 (N_16125,N_13889,N_15868);
and U16126 (N_16126,N_13845,N_12428);
or U16127 (N_16127,N_13596,N_12327);
nor U16128 (N_16128,N_14408,N_12480);
nand U16129 (N_16129,N_14476,N_12627);
and U16130 (N_16130,N_15367,N_13622);
nand U16131 (N_16131,N_12795,N_13517);
or U16132 (N_16132,N_15525,N_12649);
nand U16133 (N_16133,N_13364,N_13956);
nor U16134 (N_16134,N_14550,N_14412);
or U16135 (N_16135,N_15465,N_14512);
and U16136 (N_16136,N_12526,N_14958);
nor U16137 (N_16137,N_12565,N_15668);
nand U16138 (N_16138,N_12473,N_14357);
nand U16139 (N_16139,N_14084,N_13107);
or U16140 (N_16140,N_14808,N_14965);
nor U16141 (N_16141,N_15631,N_15777);
nor U16142 (N_16142,N_14745,N_12392);
or U16143 (N_16143,N_15529,N_12719);
nand U16144 (N_16144,N_15770,N_12634);
nand U16145 (N_16145,N_13576,N_13961);
nand U16146 (N_16146,N_13117,N_15358);
nor U16147 (N_16147,N_13996,N_12001);
or U16148 (N_16148,N_14713,N_12720);
xor U16149 (N_16149,N_15583,N_13805);
nand U16150 (N_16150,N_13321,N_15971);
xnor U16151 (N_16151,N_13608,N_13621);
and U16152 (N_16152,N_14174,N_12610);
and U16153 (N_16153,N_14453,N_12991);
or U16154 (N_16154,N_13759,N_14020);
nand U16155 (N_16155,N_12506,N_15292);
nor U16156 (N_16156,N_14505,N_14150);
nor U16157 (N_16157,N_15647,N_13658);
xor U16158 (N_16158,N_12203,N_15212);
xor U16159 (N_16159,N_12296,N_13232);
nand U16160 (N_16160,N_13794,N_13424);
nand U16161 (N_16161,N_15698,N_13496);
xnor U16162 (N_16162,N_14509,N_12044);
or U16163 (N_16163,N_14359,N_15850);
or U16164 (N_16164,N_14836,N_12684);
xor U16165 (N_16165,N_14592,N_13393);
nor U16166 (N_16166,N_15745,N_14750);
xor U16167 (N_16167,N_15051,N_15235);
or U16168 (N_16168,N_13643,N_14219);
or U16169 (N_16169,N_15446,N_12092);
or U16170 (N_16170,N_14761,N_14171);
nor U16171 (N_16171,N_14182,N_15466);
nand U16172 (N_16172,N_14739,N_15813);
nor U16173 (N_16173,N_15591,N_12857);
or U16174 (N_16174,N_15569,N_13551);
and U16175 (N_16175,N_12581,N_15158);
and U16176 (N_16176,N_12100,N_12651);
nand U16177 (N_16177,N_13624,N_13397);
xnor U16178 (N_16178,N_15293,N_14844);
xor U16179 (N_16179,N_12052,N_14806);
nand U16180 (N_16180,N_15686,N_15990);
or U16181 (N_16181,N_12231,N_15633);
nand U16182 (N_16182,N_13782,N_13251);
nand U16183 (N_16183,N_12501,N_15437);
and U16184 (N_16184,N_15732,N_12322);
nor U16185 (N_16185,N_12794,N_14532);
nand U16186 (N_16186,N_15062,N_13279);
xor U16187 (N_16187,N_13077,N_13707);
nor U16188 (N_16188,N_13368,N_14925);
and U16189 (N_16189,N_13935,N_15095);
xor U16190 (N_16190,N_15821,N_12006);
nor U16191 (N_16191,N_14501,N_13811);
nand U16192 (N_16192,N_14826,N_14682);
or U16193 (N_16193,N_15503,N_15417);
xor U16194 (N_16194,N_15862,N_14687);
or U16195 (N_16195,N_14767,N_12966);
nor U16196 (N_16196,N_13929,N_14782);
and U16197 (N_16197,N_14272,N_15210);
and U16198 (N_16198,N_15134,N_15878);
nand U16199 (N_16199,N_14567,N_12811);
and U16200 (N_16200,N_15981,N_12605);
nor U16201 (N_16201,N_13429,N_13547);
or U16202 (N_16202,N_15458,N_15567);
or U16203 (N_16203,N_14670,N_15067);
nor U16204 (N_16204,N_15861,N_12883);
or U16205 (N_16205,N_14581,N_12735);
and U16206 (N_16206,N_12820,N_14446);
and U16207 (N_16207,N_13891,N_14244);
nand U16208 (N_16208,N_13736,N_15101);
nand U16209 (N_16209,N_15251,N_15683);
nand U16210 (N_16210,N_14802,N_12191);
nor U16211 (N_16211,N_15110,N_13254);
nor U16212 (N_16212,N_13537,N_14153);
nand U16213 (N_16213,N_13567,N_13270);
nor U16214 (N_16214,N_13773,N_14946);
and U16215 (N_16215,N_12686,N_12353);
nand U16216 (N_16216,N_14633,N_15176);
xor U16217 (N_16217,N_15064,N_14499);
nor U16218 (N_16218,N_12551,N_13861);
and U16219 (N_16219,N_13724,N_12164);
nand U16220 (N_16220,N_12517,N_15873);
nand U16221 (N_16221,N_13696,N_12469);
nand U16222 (N_16222,N_15890,N_12437);
xnor U16223 (N_16223,N_13735,N_14005);
and U16224 (N_16224,N_12085,N_15301);
or U16225 (N_16225,N_12628,N_15548);
nand U16226 (N_16226,N_13063,N_15000);
nand U16227 (N_16227,N_15705,N_14339);
or U16228 (N_16228,N_13495,N_15931);
or U16229 (N_16229,N_13394,N_15702);
or U16230 (N_16230,N_13158,N_12586);
and U16231 (N_16231,N_15782,N_15028);
or U16232 (N_16232,N_13871,N_13940);
and U16233 (N_16233,N_13592,N_13671);
nand U16234 (N_16234,N_15999,N_12075);
and U16235 (N_16235,N_13632,N_14889);
or U16236 (N_16236,N_14076,N_12391);
and U16237 (N_16237,N_15822,N_15309);
xnor U16238 (N_16238,N_15199,N_12763);
or U16239 (N_16239,N_15280,N_12995);
nand U16240 (N_16240,N_15419,N_12726);
and U16241 (N_16241,N_14358,N_12463);
xor U16242 (N_16242,N_15125,N_14534);
xor U16243 (N_16243,N_15427,N_15320);
or U16244 (N_16244,N_14252,N_15893);
and U16245 (N_16245,N_14303,N_12738);
nor U16246 (N_16246,N_12877,N_14047);
xnor U16247 (N_16247,N_13354,N_12077);
and U16248 (N_16248,N_14878,N_14350);
nand U16249 (N_16249,N_14999,N_12434);
nand U16250 (N_16250,N_13231,N_14977);
xnor U16251 (N_16251,N_14292,N_14471);
or U16252 (N_16252,N_14203,N_12895);
xor U16253 (N_16253,N_14367,N_15528);
and U16254 (N_16254,N_12559,N_14647);
nor U16255 (N_16255,N_13470,N_14331);
or U16256 (N_16256,N_14964,N_15560);
xnor U16257 (N_16257,N_14305,N_14551);
or U16258 (N_16258,N_13262,N_12344);
nor U16259 (N_16259,N_12381,N_14148);
nand U16260 (N_16260,N_15362,N_15365);
nor U16261 (N_16261,N_15867,N_14388);
xor U16262 (N_16262,N_15943,N_12243);
and U16263 (N_16263,N_15757,N_15792);
or U16264 (N_16264,N_15264,N_12818);
nor U16265 (N_16265,N_14234,N_13006);
and U16266 (N_16266,N_13488,N_15070);
nand U16267 (N_16267,N_12177,N_13357);
xnor U16268 (N_16268,N_12073,N_13539);
xnor U16269 (N_16269,N_13026,N_15453);
or U16270 (N_16270,N_12982,N_14795);
nor U16271 (N_16271,N_15849,N_12484);
or U16272 (N_16272,N_15747,N_15115);
xnor U16273 (N_16273,N_13278,N_15407);
nor U16274 (N_16274,N_15149,N_13776);
and U16275 (N_16275,N_15495,N_12453);
or U16276 (N_16276,N_15678,N_15198);
and U16277 (N_16277,N_13148,N_12643);
or U16278 (N_16278,N_15207,N_14646);
nand U16279 (N_16279,N_12869,N_12830);
nand U16280 (N_16280,N_15584,N_13726);
nor U16281 (N_16281,N_12714,N_14865);
or U16282 (N_16282,N_15374,N_12490);
nor U16283 (N_16283,N_15639,N_12642);
or U16284 (N_16284,N_15985,N_15068);
xnor U16285 (N_16285,N_14362,N_12633);
nand U16286 (N_16286,N_15995,N_12339);
xor U16287 (N_16287,N_12335,N_15566);
or U16288 (N_16288,N_12448,N_12647);
xnor U16289 (N_16289,N_15392,N_15913);
nor U16290 (N_16290,N_13175,N_14924);
nor U16291 (N_16291,N_13466,N_15013);
xor U16292 (N_16292,N_13654,N_12163);
nor U16293 (N_16293,N_15720,N_14611);
nand U16294 (N_16294,N_13499,N_15588);
nand U16295 (N_16295,N_13119,N_12992);
or U16296 (N_16296,N_13128,N_15537);
nor U16297 (N_16297,N_13870,N_14624);
nand U16298 (N_16298,N_13949,N_15074);
or U16299 (N_16299,N_15368,N_15791);
nand U16300 (N_16300,N_13142,N_15448);
nand U16301 (N_16301,N_13688,N_13993);
nand U16302 (N_16302,N_13106,N_13941);
nor U16303 (N_16303,N_15806,N_13103);
nand U16304 (N_16304,N_15034,N_14010);
or U16305 (N_16305,N_12552,N_12578);
or U16306 (N_16306,N_14323,N_14268);
nor U16307 (N_16307,N_14052,N_15037);
xnor U16308 (N_16308,N_15287,N_15491);
xnor U16309 (N_16309,N_15182,N_12017);
and U16310 (N_16310,N_13887,N_15336);
nand U16311 (N_16311,N_12374,N_15089);
nand U16312 (N_16312,N_12248,N_12823);
nand U16313 (N_16313,N_13536,N_15425);
xnor U16314 (N_16314,N_15107,N_12492);
xnor U16315 (N_16315,N_14995,N_12919);
nand U16316 (N_16316,N_13644,N_12907);
and U16317 (N_16317,N_14495,N_13844);
xnor U16318 (N_16318,N_12508,N_15643);
xnor U16319 (N_16319,N_15146,N_12251);
or U16320 (N_16320,N_12931,N_13827);
and U16321 (N_16321,N_14594,N_14734);
nor U16322 (N_16322,N_14577,N_14049);
xor U16323 (N_16323,N_15096,N_15042);
nand U16324 (N_16324,N_12754,N_14810);
nand U16325 (N_16325,N_14674,N_12664);
or U16326 (N_16326,N_13711,N_13477);
and U16327 (N_16327,N_14116,N_13642);
and U16328 (N_16328,N_15079,N_15342);
xor U16329 (N_16329,N_14537,N_12699);
or U16330 (N_16330,N_12141,N_12479);
nand U16331 (N_16331,N_12158,N_13534);
xor U16332 (N_16332,N_12518,N_15549);
nor U16333 (N_16333,N_14492,N_15933);
or U16334 (N_16334,N_14097,N_14527);
or U16335 (N_16335,N_12904,N_13484);
or U16336 (N_16336,N_14652,N_15565);
xnor U16337 (N_16337,N_12020,N_12896);
or U16338 (N_16338,N_14212,N_13897);
nand U16339 (N_16339,N_12165,N_15728);
and U16340 (N_16340,N_14774,N_13412);
nor U16341 (N_16341,N_15353,N_14737);
nor U16342 (N_16342,N_13913,N_12749);
nor U16343 (N_16343,N_12299,N_12027);
and U16344 (N_16344,N_14036,N_13516);
and U16345 (N_16345,N_15291,N_14064);
nand U16346 (N_16346,N_15823,N_15273);
or U16347 (N_16347,N_12637,N_13603);
xnor U16348 (N_16348,N_13984,N_14137);
xor U16349 (N_16349,N_15189,N_12969);
or U16350 (N_16350,N_14159,N_13552);
xor U16351 (N_16351,N_15621,N_12487);
nand U16352 (N_16352,N_13761,N_12342);
and U16353 (N_16353,N_14275,N_12450);
or U16354 (N_16354,N_15384,N_15456);
and U16355 (N_16355,N_15611,N_14708);
or U16356 (N_16356,N_12264,N_14663);
nand U16357 (N_16357,N_15063,N_12695);
xnor U16358 (N_16358,N_15920,N_14333);
and U16359 (N_16359,N_15919,N_14752);
and U16360 (N_16360,N_12112,N_14405);
xnor U16361 (N_16361,N_12449,N_13853);
nand U16362 (N_16362,N_12829,N_12429);
xor U16363 (N_16363,N_13663,N_14927);
nand U16364 (N_16364,N_15496,N_14957);
xnor U16365 (N_16365,N_12800,N_13834);
xor U16366 (N_16366,N_12046,N_13689);
nand U16367 (N_16367,N_13525,N_13388);
nand U16368 (N_16368,N_15289,N_13655);
nand U16369 (N_16369,N_15632,N_12693);
xnor U16370 (N_16370,N_13016,N_13212);
nand U16371 (N_16371,N_13985,N_14441);
and U16372 (N_16372,N_13885,N_14636);
nand U16373 (N_16373,N_12089,N_13292);
nor U16374 (N_16374,N_12815,N_14540);
nor U16375 (N_16375,N_15471,N_13030);
nor U16376 (N_16376,N_14763,N_14871);
xor U16377 (N_16377,N_12476,N_14352);
and U16378 (N_16378,N_14199,N_14028);
xor U16379 (N_16379,N_13563,N_15617);
xor U16380 (N_16380,N_13291,N_13531);
nand U16381 (N_16381,N_12710,N_12841);
or U16382 (N_16382,N_15056,N_15928);
nand U16383 (N_16383,N_14538,N_13486);
nand U16384 (N_16384,N_15075,N_12345);
xnor U16385 (N_16385,N_13734,N_13256);
nand U16386 (N_16386,N_13923,N_15932);
and U16387 (N_16387,N_13937,N_14803);
or U16388 (N_16388,N_12178,N_13769);
nand U16389 (N_16389,N_12021,N_13793);
xnor U16390 (N_16390,N_13908,N_14288);
nor U16391 (N_16391,N_12802,N_15258);
nand U16392 (N_16392,N_13187,N_14574);
and U16393 (N_16393,N_12626,N_14984);
nand U16394 (N_16394,N_12537,N_14775);
or U16395 (N_16395,N_12337,N_13229);
and U16396 (N_16396,N_14705,N_13228);
or U16397 (N_16397,N_14562,N_12755);
and U16398 (N_16398,N_13783,N_13432);
nand U16399 (N_16399,N_14879,N_13819);
nand U16400 (N_16400,N_13543,N_13522);
or U16401 (N_16401,N_13804,N_15780);
nor U16402 (N_16402,N_12025,N_13982);
or U16403 (N_16403,N_12454,N_14829);
nand U16404 (N_16404,N_13741,N_12297);
and U16405 (N_16405,N_15508,N_13444);
nor U16406 (N_16406,N_12058,N_15662);
and U16407 (N_16407,N_12838,N_13064);
nand U16408 (N_16408,N_12849,N_13204);
or U16409 (N_16409,N_15015,N_14034);
nor U16410 (N_16410,N_13304,N_14792);
or U16411 (N_16411,N_14903,N_12423);
nor U16412 (N_16412,N_12901,N_15903);
and U16413 (N_16413,N_13753,N_15255);
nor U16414 (N_16414,N_14406,N_12443);
nand U16415 (N_16415,N_12854,N_13174);
nand U16416 (N_16416,N_15180,N_12419);
xnor U16417 (N_16417,N_15159,N_13922);
nand U16418 (N_16418,N_12090,N_14213);
or U16419 (N_16419,N_13750,N_13521);
or U16420 (N_16420,N_14085,N_15299);
and U16421 (N_16421,N_15359,N_12842);
or U16422 (N_16422,N_12858,N_12805);
and U16423 (N_16423,N_12056,N_12674);
nand U16424 (N_16424,N_14665,N_12134);
nor U16425 (N_16425,N_15058,N_13669);
and U16426 (N_16426,N_13931,N_12663);
nor U16427 (N_16427,N_12728,N_14250);
xnor U16428 (N_16428,N_14197,N_12798);
or U16429 (N_16429,N_15229,N_15530);
or U16430 (N_16430,N_15156,N_12185);
nand U16431 (N_16431,N_15544,N_12893);
xor U16432 (N_16432,N_15382,N_13075);
nor U16433 (N_16433,N_13057,N_15518);
nor U16434 (N_16434,N_15687,N_12539);
nor U16435 (N_16435,N_15173,N_14389);
xnor U16436 (N_16436,N_13150,N_13950);
xnor U16437 (N_16437,N_14493,N_13401);
and U16438 (N_16438,N_13789,N_15946);
nand U16439 (N_16439,N_14691,N_12403);
nor U16440 (N_16440,N_12589,N_14143);
or U16441 (N_16441,N_14165,N_14768);
xnor U16442 (N_16442,N_14172,N_14922);
nor U16443 (N_16443,N_13743,N_15276);
and U16444 (N_16444,N_12696,N_14864);
and U16445 (N_16445,N_14278,N_13065);
nor U16446 (N_16446,N_13351,N_14081);
or U16447 (N_16447,N_15211,N_15060);
and U16448 (N_16448,N_15536,N_13370);
or U16449 (N_16449,N_15915,N_15213);
nor U16450 (N_16450,N_15175,N_13515);
xnor U16451 (N_16451,N_12507,N_12129);
nand U16452 (N_16452,N_15347,N_15902);
or U16453 (N_16453,N_15924,N_15422);
nand U16454 (N_16454,N_12971,N_12421);
and U16455 (N_16455,N_14434,N_15670);
and U16456 (N_16456,N_12465,N_14091);
or U16457 (N_16457,N_12495,N_12687);
and U16458 (N_16458,N_15534,N_12511);
and U16459 (N_16459,N_13489,N_15084);
xnor U16460 (N_16460,N_13986,N_15140);
xor U16461 (N_16461,N_13857,N_15082);
nand U16462 (N_16462,N_15412,N_12538);
or U16463 (N_16463,N_13009,N_14196);
nand U16464 (N_16464,N_13374,N_14973);
and U16465 (N_16465,N_13493,N_15644);
nand U16466 (N_16466,N_13272,N_15024);
xor U16467 (N_16467,N_12839,N_15169);
xnor U16468 (N_16468,N_12870,N_15026);
and U16469 (N_16469,N_14511,N_15987);
nand U16470 (N_16470,N_15477,N_15974);
nand U16471 (N_16471,N_15214,N_14835);
or U16472 (N_16472,N_13705,N_14192);
xnor U16473 (N_16473,N_13659,N_12880);
and U16474 (N_16474,N_14279,N_13988);
nand U16475 (N_16475,N_15969,N_15267);
xor U16476 (N_16476,N_14832,N_13441);
or U16477 (N_16477,N_15463,N_14112);
nand U16478 (N_16478,N_13849,N_12645);
xor U16479 (N_16479,N_15455,N_12007);
or U16480 (N_16480,N_13972,N_14719);
xnor U16481 (N_16481,N_14778,N_13410);
and U16482 (N_16482,N_14113,N_15657);
nor U16483 (N_16483,N_13708,N_15234);
nand U16484 (N_16484,N_15845,N_12128);
xor U16485 (N_16485,N_13572,N_15616);
and U16486 (N_16486,N_13926,N_13300);
and U16487 (N_16487,N_14915,N_12051);
nand U16488 (N_16488,N_15892,N_14553);
or U16489 (N_16489,N_12279,N_14458);
and U16490 (N_16490,N_14510,N_12885);
and U16491 (N_16491,N_12301,N_12597);
xor U16492 (N_16492,N_15073,N_12183);
xnor U16493 (N_16493,N_12034,N_12146);
xnor U16494 (N_16494,N_14411,N_14890);
nor U16495 (N_16495,N_12142,N_14672);
or U16496 (N_16496,N_12115,N_13615);
nor U16497 (N_16497,N_14393,N_14867);
xnor U16498 (N_16498,N_12071,N_15798);
and U16499 (N_16499,N_12205,N_12737);
xnor U16500 (N_16500,N_12619,N_12488);
nor U16501 (N_16501,N_15078,N_13365);
or U16502 (N_16502,N_14484,N_13886);
or U16503 (N_16503,N_13498,N_14680);
xor U16504 (N_16504,N_13352,N_13312);
nand U16505 (N_16505,N_13605,N_15355);
xnor U16506 (N_16506,N_14726,N_12930);
and U16507 (N_16507,N_15030,N_15120);
nand U16508 (N_16508,N_13122,N_12011);
nand U16509 (N_16509,N_13638,N_13094);
and U16510 (N_16510,N_14083,N_12781);
xnor U16511 (N_16511,N_12851,N_13699);
xnor U16512 (N_16512,N_15010,N_12743);
xor U16513 (N_16513,N_13839,N_13830);
and U16514 (N_16514,N_15711,N_13969);
xnor U16515 (N_16515,N_13970,N_14781);
xor U16516 (N_16516,N_14843,N_13055);
nor U16517 (N_16517,N_12746,N_13146);
nand U16518 (N_16518,N_12984,N_12646);
xor U16519 (N_16519,N_14884,N_15283);
nor U16520 (N_16520,N_14257,N_12475);
and U16521 (N_16521,N_15041,N_15092);
and U16522 (N_16522,N_14923,N_14727);
nand U16523 (N_16523,N_14947,N_14356);
nand U16524 (N_16524,N_12612,N_12455);
nand U16525 (N_16525,N_14723,N_15499);
nand U16526 (N_16526,N_14160,N_14289);
nor U16527 (N_16527,N_12033,N_14721);
and U16528 (N_16528,N_13955,N_15261);
or U16529 (N_16529,N_13874,N_14514);
nor U16530 (N_16530,N_13007,N_14063);
and U16531 (N_16531,N_13180,N_15185);
xnor U16532 (N_16532,N_14729,N_15927);
xnor U16533 (N_16533,N_15093,N_14962);
xnor U16534 (N_16534,N_13465,N_13513);
xnor U16535 (N_16535,N_14710,N_15326);
xor U16536 (N_16536,N_15265,N_13701);
and U16537 (N_16537,N_14035,N_15117);
or U16538 (N_16538,N_12528,N_15807);
xor U16539 (N_16539,N_13530,N_15740);
nand U16540 (N_16540,N_15779,N_15145);
nor U16541 (N_16541,N_14233,N_13509);
and U16542 (N_16542,N_12601,N_15363);
nor U16543 (N_16543,N_12848,N_13482);
nor U16544 (N_16544,N_15500,N_14460);
xnor U16545 (N_16545,N_13652,N_14980);
xor U16546 (N_16546,N_13402,N_12861);
xnor U16547 (N_16547,N_15824,N_14907);
nand U16548 (N_16548,N_12996,N_13593);
or U16549 (N_16549,N_12644,N_15839);
xnor U16550 (N_16550,N_12218,N_15842);
xnor U16551 (N_16551,N_12785,N_15604);
or U16552 (N_16552,N_14119,N_15921);
xor U16553 (N_16553,N_15636,N_13613);
and U16554 (N_16554,N_14424,N_13085);
xor U16555 (N_16555,N_15579,N_13626);
and U16556 (N_16556,N_15464,N_13999);
and U16557 (N_16557,N_14731,N_13943);
or U16558 (N_16558,N_15590,N_14372);
nor U16559 (N_16559,N_14184,N_15840);
or U16560 (N_16560,N_14859,N_13125);
and U16561 (N_16561,N_13359,N_14796);
xor U16562 (N_16562,N_14759,N_15411);
and U16563 (N_16563,N_12274,N_15308);
nor U16564 (N_16564,N_13907,N_13556);
nor U16565 (N_16565,N_13812,N_12102);
and U16566 (N_16566,N_12585,N_12716);
xnor U16567 (N_16567,N_14866,N_14435);
or U16568 (N_16568,N_14198,N_13722);
or U16569 (N_16569,N_14173,N_14585);
and U16570 (N_16570,N_15083,N_13250);
nor U16571 (N_16571,N_13092,N_14329);
and U16572 (N_16572,N_13403,N_15143);
xnor U16573 (N_16573,N_14245,N_15296);
and U16574 (N_16574,N_14571,N_14144);
xnor U16575 (N_16575,N_12285,N_12500);
and U16576 (N_16576,N_12515,N_14224);
nand U16577 (N_16577,N_12157,N_15155);
or U16578 (N_16578,N_15672,N_15751);
or U16579 (N_16579,N_15936,N_12376);
nand U16580 (N_16580,N_15369,N_12807);
or U16581 (N_16581,N_12801,N_13311);
xor U16582 (N_16582,N_15897,N_15277);
nor U16583 (N_16583,N_13309,N_15443);
nor U16584 (N_16584,N_13442,N_13053);
xor U16585 (N_16585,N_13901,N_14325);
or U16586 (N_16586,N_14677,N_14287);
or U16587 (N_16587,N_14660,N_12575);
nor U16588 (N_16588,N_14026,N_12561);
nor U16589 (N_16589,N_13927,N_13062);
and U16590 (N_16590,N_12491,N_15618);
nand U16591 (N_16591,N_15970,N_13218);
xnor U16592 (N_16592,N_15023,N_12855);
xor U16593 (N_16593,N_14580,N_14022);
and U16594 (N_16594,N_14348,N_13267);
nor U16595 (N_16595,N_14678,N_15696);
nor U16596 (N_16596,N_12658,N_14040);
nor U16597 (N_16597,N_14648,N_12341);
and U16598 (N_16598,N_15874,N_12916);
and U16599 (N_16599,N_12072,N_13932);
xnor U16600 (N_16600,N_13587,N_14164);
nor U16601 (N_16601,N_13137,N_14454);
nand U16602 (N_16602,N_12588,N_13341);
nor U16603 (N_16603,N_15723,N_13758);
nor U16604 (N_16604,N_13091,N_12217);
xnor U16605 (N_16605,N_14985,N_13905);
or U16606 (N_16606,N_15557,N_14094);
nand U16607 (N_16607,N_15132,N_14074);
or U16608 (N_16608,N_15673,N_14230);
nand U16609 (N_16609,N_15473,N_13111);
xnor U16610 (N_16610,N_15350,N_12604);
nand U16611 (N_16611,N_13405,N_14218);
and U16612 (N_16612,N_15303,N_14161);
and U16613 (N_16613,N_14018,N_13953);
or U16614 (N_16614,N_14061,N_15721);
nor U16615 (N_16615,N_13431,N_15399);
and U16616 (N_16616,N_12208,N_14301);
nor U16617 (N_16617,N_15393,N_12557);
or U16618 (N_16618,N_15864,N_14365);
and U16619 (N_16619,N_13867,N_12990);
nor U16620 (N_16620,N_14024,N_12591);
and U16621 (N_16621,N_12734,N_12404);
nor U16622 (N_16622,N_13109,N_14311);
nand U16623 (N_16623,N_15324,N_12471);
nand U16624 (N_16624,N_15853,N_12312);
nand U16625 (N_16625,N_14645,N_12195);
xor U16626 (N_16626,N_15497,N_15577);
xor U16627 (N_16627,N_13396,N_15761);
or U16628 (N_16628,N_15978,N_12678);
or U16629 (N_16629,N_14324,N_13472);
and U16630 (N_16630,N_14563,N_13540);
or U16631 (N_16631,N_13991,N_12214);
or U16632 (N_16632,N_15020,N_13206);
nor U16633 (N_16633,N_14131,N_14322);
and U16634 (N_16634,N_14988,N_14658);
nand U16635 (N_16635,N_15300,N_13162);
and U16636 (N_16636,N_12951,N_12918);
or U16637 (N_16637,N_12370,N_13668);
or U16638 (N_16638,N_14519,N_14593);
nand U16639 (N_16639,N_13093,N_13575);
nor U16640 (N_16640,N_12512,N_12008);
and U16641 (N_16641,N_14068,N_15624);
and U16642 (N_16642,N_12401,N_15522);
nand U16643 (N_16643,N_12078,N_15253);
nor U16644 (N_16644,N_15398,N_15054);
nand U16645 (N_16645,N_13791,N_15097);
nand U16646 (N_16646,N_15288,N_13675);
nor U16647 (N_16647,N_14270,N_12669);
or U16648 (N_16648,N_15341,N_15638);
nor U16649 (N_16649,N_12689,N_13733);
and U16650 (N_16650,N_15451,N_15119);
nand U16651 (N_16651,N_14828,N_15241);
xnor U16652 (N_16652,N_14452,N_15240);
xnor U16653 (N_16653,N_14390,N_14355);
or U16654 (N_16654,N_14055,N_14217);
nor U16655 (N_16655,N_15997,N_14003);
nor U16656 (N_16656,N_15114,N_13921);
nand U16657 (N_16657,N_12950,N_13813);
nor U16658 (N_16658,N_14508,N_15959);
nand U16659 (N_16659,N_12256,N_14105);
nor U16660 (N_16660,N_14838,N_14560);
xor U16661 (N_16661,N_15428,N_12782);
and U16662 (N_16662,N_13807,N_14953);
and U16663 (N_16663,N_13727,N_15099);
and U16664 (N_16664,N_14078,N_14531);
xnor U16665 (N_16665,N_14715,N_12472);
or U16666 (N_16666,N_14856,N_15934);
nor U16667 (N_16667,N_15219,N_13906);
nand U16668 (N_16668,N_12953,N_14254);
and U16669 (N_16669,N_12970,N_14535);
nor U16670 (N_16670,N_15700,N_14163);
and U16671 (N_16671,N_13129,N_14370);
xor U16672 (N_16672,N_13473,N_12048);
xor U16673 (N_16673,N_13990,N_13061);
xor U16674 (N_16674,N_13558,N_14135);
nand U16675 (N_16675,N_15057,N_12127);
xor U16676 (N_16676,N_15756,N_14391);
nor U16677 (N_16677,N_12752,N_15268);
nor U16678 (N_16678,N_15168,N_14749);
nor U16679 (N_16679,N_14448,N_14426);
nor U16680 (N_16680,N_13760,N_13550);
and U16681 (N_16681,N_14983,N_13656);
and U16682 (N_16682,N_12617,N_15914);
nand U16683 (N_16683,N_13673,N_12067);
nor U16684 (N_16684,N_15713,N_12103);
nand U16685 (N_16685,N_15735,N_14996);
or U16686 (N_16686,N_12412,N_14766);
and U16687 (N_16687,N_13002,N_13285);
nand U16688 (N_16688,N_15812,N_14176);
nor U16689 (N_16689,N_12036,N_13600);
nor U16690 (N_16690,N_14524,N_13890);
xor U16691 (N_16691,N_15578,N_13266);
and U16692 (N_16692,N_13549,N_15200);
nand U16693 (N_16693,N_15582,N_13557);
and U16694 (N_16694,N_13647,N_15442);
and U16695 (N_16695,N_12360,N_15546);
nor U16696 (N_16696,N_12436,N_14392);
xnor U16697 (N_16697,N_14895,N_13698);
or U16698 (N_16698,N_15343,N_14189);
or U16699 (N_16699,N_14447,N_12233);
xor U16700 (N_16700,N_15139,N_13014);
nor U16701 (N_16701,N_13520,N_12375);
xnor U16702 (N_16702,N_14518,N_13980);
nand U16703 (N_16703,N_15554,N_12593);
xnor U16704 (N_16704,N_12010,N_13523);
and U16705 (N_16705,N_12690,N_12168);
nor U16706 (N_16706,N_13903,N_14554);
xnor U16707 (N_16707,N_13825,N_12150);
nand U16708 (N_16708,N_14753,N_15138);
xor U16709 (N_16709,N_13918,N_15808);
xor U16710 (N_16710,N_13144,N_15547);
nand U16711 (N_16711,N_13780,N_14477);
and U16712 (N_16712,N_13633,N_14893);
nor U16713 (N_16713,N_15224,N_14787);
nor U16714 (N_16714,N_13205,N_15502);
nor U16715 (N_16715,N_12744,N_14146);
nor U16716 (N_16716,N_12277,N_13056);
xnor U16717 (N_16717,N_15290,N_12606);
xnor U16718 (N_16718,N_15305,N_14006);
nor U16719 (N_16719,N_14188,N_12043);
nor U16720 (N_16720,N_13958,N_15193);
xor U16721 (N_16721,N_13102,N_14722);
or U16722 (N_16722,N_15916,N_14862);
xor U16723 (N_16723,N_15421,N_13260);
nand U16724 (N_16724,N_14222,N_15800);
or U16725 (N_16725,N_14202,N_12095);
or U16726 (N_16726,N_15423,N_15961);
xnor U16727 (N_16727,N_14949,N_13423);
or U16728 (N_16728,N_13084,N_14709);
or U16729 (N_16729,N_15710,N_15014);
xor U16730 (N_16730,N_12207,N_14586);
nand U16731 (N_16731,N_13744,N_13965);
nor U16732 (N_16732,N_14166,N_13518);
or U16733 (N_16733,N_13545,N_15833);
nor U16734 (N_16734,N_12457,N_12732);
xnor U16735 (N_16735,N_15033,N_15556);
xnor U16736 (N_16736,N_13639,N_15513);
nand U16737 (N_16737,N_12595,N_14811);
or U16738 (N_16738,N_12929,N_15859);
nor U16739 (N_16739,N_15484,N_14075);
xor U16740 (N_16740,N_12772,N_12653);
nand U16741 (N_16741,N_12055,N_13836);
and U16742 (N_16742,N_15220,N_15126);
xnor U16743 (N_16743,N_14248,N_14427);
and U16744 (N_16744,N_12656,N_12179);
xnor U16745 (N_16745,N_12002,N_13184);
nand U16746 (N_16746,N_15625,N_14281);
nand U16747 (N_16747,N_13096,N_14475);
nand U16748 (N_16748,N_13519,N_12405);
nor U16749 (N_16749,N_14384,N_13199);
xnor U16750 (N_16750,N_13771,N_15416);
and U16751 (N_16751,N_12332,N_14294);
and U16752 (N_16752,N_14332,N_15538);
nor U16753 (N_16753,N_13284,N_15734);
nand U16754 (N_16754,N_13553,N_14051);
or U16755 (N_16755,N_13446,N_14407);
nor U16756 (N_16756,N_14423,N_12520);
and U16757 (N_16757,N_13261,N_13510);
xor U16758 (N_16758,N_13389,N_15898);
nor U16759 (N_16759,N_15553,N_14221);
or U16760 (N_16760,N_15380,N_15712);
xnor U16761 (N_16761,N_14046,N_14588);
or U16762 (N_16762,N_14765,N_15619);
xnor U16763 (N_16763,N_14033,N_12965);
or U16764 (N_16764,N_15944,N_14888);
and U16765 (N_16765,N_13691,N_13089);
nor U16766 (N_16766,N_14297,N_15225);
nand U16767 (N_16767,N_13264,N_12294);
xor U16768 (N_16768,N_12709,N_15272);
xor U16769 (N_16769,N_12542,N_13379);
and U16770 (N_16770,N_15571,N_13020);
nand U16771 (N_16771,N_15480,N_12832);
nand U16772 (N_16772,N_15231,N_13840);
or U16773 (N_16773,N_13247,N_15739);
or U16774 (N_16774,N_15410,N_13747);
nand U16775 (N_16775,N_14383,N_12013);
xnor U16776 (N_16776,N_15708,N_13657);
nand U16777 (N_16777,N_13458,N_13099);
or U16778 (N_16778,N_15912,N_14271);
and U16779 (N_16779,N_14503,N_15237);
nor U16780 (N_16780,N_12349,N_14265);
or U16781 (N_16781,N_14100,N_13512);
and U16782 (N_16782,N_15019,N_12936);
and U16783 (N_16783,N_14309,N_13375);
nor U16784 (N_16784,N_14814,N_13436);
and U16785 (N_16785,N_13957,N_12303);
nor U16786 (N_16786,N_12865,N_12562);
nor U16787 (N_16787,N_15476,N_15482);
and U16788 (N_16788,N_12623,N_15982);
xor U16789 (N_16789,N_12884,N_12435);
and U16790 (N_16790,N_14185,N_12502);
or U16791 (N_16791,N_13238,N_12770);
nand U16792 (N_16792,N_13898,N_15085);
xor U16793 (N_16793,N_12560,N_12910);
nor U16794 (N_16794,N_12717,N_14368);
or U16795 (N_16795,N_13634,N_12638);
and U16796 (N_16796,N_13310,N_13457);
xor U16797 (N_16797,N_13203,N_12041);
xor U16798 (N_16798,N_12306,N_12053);
xor U16799 (N_16799,N_12227,N_14917);
xor U16800 (N_16800,N_13686,N_12567);
and U16801 (N_16801,N_13800,N_14487);
or U16802 (N_16802,N_13387,N_12514);
nand U16803 (N_16803,N_12603,N_14327);
and U16804 (N_16804,N_14186,N_15891);
xor U16805 (N_16805,N_15203,N_15949);
and U16806 (N_16806,N_12430,N_14127);
or U16807 (N_16807,N_13742,N_12268);
xor U16808 (N_16808,N_15017,N_13363);
nand U16809 (N_16809,N_13739,N_13059);
and U16810 (N_16810,N_12868,N_14870);
and U16811 (N_16811,N_14012,N_15284);
nand U16812 (N_16812,N_14754,N_12050);
nand U16813 (N_16813,N_13468,N_14283);
or U16814 (N_16814,N_12804,N_12887);
nor U16815 (N_16815,N_14247,N_12532);
nor U16816 (N_16816,N_14706,N_12505);
nand U16817 (N_16817,N_14625,N_12276);
nor U16818 (N_16818,N_14422,N_13784);
nand U16819 (N_16819,N_14472,N_12175);
nand U16820 (N_16820,N_15830,N_14183);
nand U16821 (N_16821,N_13038,N_13438);
and U16822 (N_16822,N_12176,N_12190);
nand U16823 (N_16823,N_14312,N_14504);
or U16824 (N_16824,N_12422,N_15778);
xnor U16825 (N_16825,N_14926,N_13582);
and U16826 (N_16826,N_14930,N_12170);
nand U16827 (N_16827,N_12534,N_14959);
and U16828 (N_16828,N_13070,N_12949);
and U16829 (N_16829,N_15656,N_12631);
and U16830 (N_16830,N_13487,N_15524);
nor U16831 (N_16831,N_13001,N_15361);
xnor U16832 (N_16832,N_13339,N_12250);
nor U16833 (N_16833,N_13872,N_15956);
and U16834 (N_16834,N_15627,N_13964);
xor U16835 (N_16835,N_12398,N_13338);
and U16836 (N_16836,N_14496,N_15860);
nor U16837 (N_16837,N_14366,N_15413);
and U16838 (N_16838,N_15642,N_15765);
nor U16839 (N_16839,N_12169,N_13360);
nand U16840 (N_16840,N_15029,N_12049);
and U16841 (N_16841,N_12026,N_13398);
or U16842 (N_16842,N_15783,N_15819);
and U16843 (N_16843,N_12130,N_14622);
nand U16844 (N_16844,N_13882,N_12676);
or U16845 (N_16845,N_15043,N_15103);
nand U16846 (N_16846,N_14943,N_12989);
or U16847 (N_16847,N_15346,N_15313);
xor U16848 (N_16848,N_14338,N_12239);
nor U16849 (N_16849,N_15854,N_14526);
nand U16850 (N_16850,N_13942,N_15131);
or U16851 (N_16851,N_13213,N_12762);
and U16852 (N_16852,N_14992,N_12523);
and U16853 (N_16853,N_13565,N_14698);
nor U16854 (N_16854,N_13851,N_13435);
nor U16855 (N_16855,N_12666,N_15420);
nor U16856 (N_16856,N_13259,N_12958);
nor U16857 (N_16857,N_15161,N_14124);
or U16858 (N_16858,N_12273,N_13674);
nand U16859 (N_16859,N_13217,N_13846);
and U16860 (N_16860,N_15205,N_12963);
nor U16861 (N_16861,N_15113,N_13323);
and U16862 (N_16862,N_12723,N_12715);
nand U16863 (N_16863,N_13445,N_14354);
or U16864 (N_16864,N_12618,N_12225);
and U16865 (N_16865,N_12145,N_14225);
xor U16866 (N_16866,N_14151,N_13879);
or U16867 (N_16867,N_14053,N_14800);
nand U16868 (N_16868,N_12812,N_14468);
and U16869 (N_16869,N_13127,N_13302);
nor U16870 (N_16870,N_15244,N_12365);
xor U16871 (N_16871,N_14707,N_13555);
or U16872 (N_16872,N_13200,N_12776);
xor U16873 (N_16873,N_14610,N_15615);
nor U16874 (N_16874,N_12788,N_13777);
nor U16875 (N_16875,N_13629,N_13386);
xnor U16876 (N_16876,N_13916,N_12625);
and U16877 (N_16877,N_14122,N_14690);
and U16878 (N_16878,N_12123,N_12040);
or U16879 (N_16879,N_15390,N_12324);
nand U16880 (N_16880,N_15693,N_15468);
nor U16881 (N_16881,N_13607,N_14688);
and U16882 (N_16882,N_12333,N_14481);
and U16883 (N_16883,N_13611,N_14549);
or U16884 (N_16884,N_15262,N_13198);
and U16885 (N_16885,N_12747,N_12483);
nand U16886 (N_16886,N_13149,N_13367);
xor U16887 (N_16887,N_13451,N_13223);
and U16888 (N_16888,N_12615,N_15196);
nor U16889 (N_16889,N_12793,N_15447);
and U16890 (N_16890,N_14464,N_14780);
nor U16891 (N_16891,N_12459,N_14086);
or U16892 (N_16892,N_14881,N_15462);
nand U16893 (N_16893,N_12395,N_14876);
xnor U16894 (N_16894,N_15882,N_14011);
and U16895 (N_16895,N_12113,N_15376);
nand U16896 (N_16896,N_13685,N_13366);
or U16897 (N_16897,N_15217,N_14004);
nor U16898 (N_16898,N_12915,N_15789);
nand U16899 (N_16899,N_14669,N_14897);
nand U16900 (N_16900,N_15165,N_13207);
nor U16901 (N_16901,N_13406,N_12621);
nor U16902 (N_16902,N_12149,N_13415);
xnor U16903 (N_16903,N_15232,N_15190);
or U16904 (N_16904,N_12673,N_14998);
or U16905 (N_16905,N_13809,N_13480);
xor U16906 (N_16906,N_13322,N_12367);
or U16907 (N_16907,N_12257,N_14874);
and U16908 (N_16908,N_13873,N_14241);
xor U16909 (N_16909,N_15153,N_15230);
nor U16910 (N_16910,N_12076,N_15724);
and U16911 (N_16911,N_15055,N_15857);
or U16912 (N_16912,N_15908,N_12057);
nand U16913 (N_16913,N_14525,N_12117);
nor U16914 (N_16914,N_15866,N_15081);
nand U16915 (N_16915,N_13706,N_13717);
nor U16916 (N_16916,N_12890,N_14382);
nor U16917 (N_16917,N_12874,N_14891);
xnor U16918 (N_16918,N_15252,N_12143);
xor U16919 (N_16919,N_15744,N_12497);
nor U16920 (N_16920,N_14756,N_12105);
xnor U16921 (N_16921,N_15450,N_14128);
and U16922 (N_16922,N_14568,N_13619);
and U16923 (N_16923,N_13306,N_13900);
and U16924 (N_16924,N_13185,N_14007);
nor U16925 (N_16925,N_13583,N_14318);
nand U16926 (N_16926,N_12654,N_15992);
xnor U16927 (N_16927,N_15470,N_15136);
xor U16928 (N_16928,N_14251,N_15895);
xnor U16929 (N_16929,N_15018,N_14711);
nor U16930 (N_16930,N_15976,N_12159);
xor U16931 (N_16931,N_12254,N_12439);
nor U16932 (N_16932,N_13133,N_13876);
or U16933 (N_16933,N_13335,N_14002);
or U16934 (N_16934,N_12221,N_14738);
or U16935 (N_16935,N_12184,N_14223);
nor U16936 (N_16936,N_13289,N_12244);
or U16937 (N_16937,N_13275,N_14321);
xnor U16938 (N_16938,N_15460,N_13485);
nand U16939 (N_16939,N_15439,N_13349);
xor U16940 (N_16940,N_15966,N_13731);
nor U16941 (N_16941,N_15814,N_14615);
or U16942 (N_16942,N_12192,N_14770);
xnor U16943 (N_16943,N_15228,N_12813);
nor U16944 (N_16944,N_15935,N_13108);
nand U16945 (N_16945,N_12357,N_15208);
or U16946 (N_16946,N_13821,N_13720);
xor U16947 (N_16947,N_14417,N_12023);
nor U16948 (N_16948,N_14757,N_14343);
nor U16949 (N_16949,N_13797,N_14675);
and U16950 (N_16950,N_15216,N_13529);
nor U16951 (N_16951,N_15483,N_13046);
or U16952 (N_16952,N_13326,N_12891);
nor U16953 (N_16953,N_12558,N_14483);
xnor U16954 (N_16954,N_13474,N_13013);
nand U16955 (N_16955,N_15005,N_13822);
or U16956 (N_16956,N_14008,N_14015);
and U16957 (N_16957,N_12819,N_12543);
xor U16958 (N_16958,N_15221,N_15105);
nor U16959 (N_16959,N_13277,N_15494);
nand U16960 (N_16960,N_14121,N_14486);
or U16961 (N_16961,N_13936,N_14944);
or U16962 (N_16962,N_15545,N_12099);
nand U16963 (N_16963,N_14149,N_13974);
nand U16964 (N_16964,N_14302,N_15889);
nand U16965 (N_16965,N_12994,N_14451);
nand U16966 (N_16966,N_14201,N_15766);
or U16967 (N_16967,N_12131,N_12570);
or U16968 (N_16968,N_14627,N_15371);
and U16969 (N_16969,N_14702,N_13350);
xor U16970 (N_16970,N_15172,N_15781);
nand U16971 (N_16971,N_15004,N_14442);
nor U16972 (N_16972,N_15162,N_14291);
xnor U16973 (N_16973,N_12999,N_15886);
nor U16974 (N_16974,N_13043,N_15315);
nor U16975 (N_16975,N_12680,N_13778);
nand U16976 (N_16976,N_15087,N_12675);
nand U16977 (N_16977,N_14162,N_13749);
nand U16978 (N_16978,N_15106,N_15142);
xnor U16979 (N_16979,N_15171,N_15730);
nand U16980 (N_16980,N_15152,N_14516);
nand U16981 (N_16981,N_15957,N_12414);
nor U16982 (N_16982,N_14616,N_12579);
nor U16983 (N_16983,N_15426,N_12156);
or U16984 (N_16984,N_13179,N_12330);
xor U16985 (N_16985,N_13697,N_15257);
and U16986 (N_16986,N_15454,N_13815);
or U16987 (N_16987,N_12668,N_14639);
nand U16988 (N_16988,N_13265,N_14102);
nand U16989 (N_16989,N_13023,N_13541);
xor U16990 (N_16990,N_14032,N_14269);
xnor U16991 (N_16991,N_15665,N_14583);
and U16992 (N_16992,N_13334,N_15178);
nand U16993 (N_16993,N_12569,N_14655);
nand U16994 (N_16994,N_14410,N_12331);
xor U16995 (N_16995,N_12242,N_13086);
xnor U16996 (N_16996,N_12305,N_15279);
nor U16997 (N_16997,N_15689,N_14530);
nand U16998 (N_16998,N_14425,N_14736);
nor U16999 (N_16999,N_12171,N_15758);
xnor U17000 (N_17000,N_14769,N_15441);
xor U17001 (N_17001,N_12122,N_15767);
and U17002 (N_17002,N_13152,N_12478);
xor U17003 (N_17003,N_15100,N_12028);
nand U17004 (N_17004,N_15661,N_12833);
xnor U17005 (N_17005,N_15429,N_12764);
nand U17006 (N_17006,N_12914,N_13712);
and U17007 (N_17007,N_14523,N_14894);
xor U17008 (N_17008,N_14883,N_12137);
nor U17009 (N_17009,N_14784,N_12927);
nor U17010 (N_17010,N_14142,N_15746);
or U17011 (N_17011,N_12037,N_15404);
or U17012 (N_17012,N_15659,N_15338);
nand U17013 (N_17013,N_13833,N_12154);
and U17014 (N_17014,N_14528,N_14236);
or U17015 (N_17015,N_12955,N_15040);
and U17016 (N_17016,N_14016,N_15151);
nand U17017 (N_17017,N_12742,N_15246);
nand U17018 (N_17018,N_14098,N_12816);
and U17019 (N_17019,N_15157,N_12736);
and U17020 (N_17020,N_14045,N_13772);
or U17021 (N_17021,N_13132,N_14533);
nand U17022 (N_17022,N_12240,N_12235);
or U17023 (N_17023,N_15869,N_12706);
and U17024 (N_17024,N_13947,N_14349);
or U17025 (N_17025,N_13283,N_15810);
nand U17026 (N_17026,N_15983,N_14319);
and U17027 (N_17027,N_13170,N_15909);
and U17028 (N_17028,N_13018,N_13035);
nor U17029 (N_17029,N_14596,N_15403);
and U17030 (N_17030,N_12139,N_14462);
and U17031 (N_17031,N_15788,N_12705);
nor U17032 (N_17032,N_15979,N_13380);
nand U17033 (N_17033,N_13191,N_14619);
and U17034 (N_17034,N_13571,N_13121);
nor U17035 (N_17035,N_12186,N_12864);
nor U17036 (N_17036,N_12946,N_14243);
xor U17037 (N_17037,N_14258,N_15964);
nand U17038 (N_17038,N_14057,N_14975);
nor U17039 (N_17039,N_15848,N_13467);
nand U17040 (N_17040,N_15671,N_12853);
xor U17041 (N_17041,N_15608,N_13928);
or U17042 (N_17042,N_13637,N_12739);
nand U17043 (N_17043,N_15794,N_13532);
nor U17044 (N_17044,N_12938,N_14330);
nor U17045 (N_17045,N_12160,N_15626);
nor U17046 (N_17046,N_13303,N_15490);
or U17047 (N_17047,N_13025,N_14232);
and U17048 (N_17048,N_13959,N_13880);
and U17049 (N_17049,N_14208,N_12094);
xnor U17050 (N_17050,N_14880,N_15856);
nand U17051 (N_17051,N_12826,N_13803);
nor U17052 (N_17052,N_13383,N_14679);
xnor U17053 (N_17053,N_13101,N_13421);
or U17054 (N_17054,N_14377,N_13210);
nor U17055 (N_17055,N_15851,N_15998);
xnor U17056 (N_17056,N_12271,N_13138);
nand U17057 (N_17057,N_12863,N_14603);
nor U17058 (N_17058,N_13987,N_15681);
nor U17059 (N_17059,N_13194,N_13838);
nor U17060 (N_17060,N_15009,N_15038);
nand U17061 (N_17061,N_13130,N_15938);
xor U17062 (N_17062,N_14041,N_15486);
nor U17063 (N_17063,N_13858,N_12960);
or U17064 (N_17064,N_15953,N_15197);
and U17065 (N_17065,N_15879,N_12408);
nand U17066 (N_17066,N_13329,N_13221);
xor U17067 (N_17067,N_12093,N_14887);
xor U17068 (N_17068,N_14755,N_12757);
or U17069 (N_17069,N_13635,N_15281);
and U17070 (N_17070,N_14714,N_12356);
nor U17071 (N_17071,N_14450,N_14179);
xnor U17072 (N_17072,N_15540,N_13045);
or U17073 (N_17073,N_13770,N_15731);
nand U17074 (N_17074,N_14228,N_12703);
and U17075 (N_17075,N_12821,N_15433);
or U17076 (N_17076,N_12302,N_13342);
or U17077 (N_17077,N_15762,N_14846);
and U17078 (N_17078,N_12882,N_14733);
or U17079 (N_17079,N_12648,N_14474);
nand U17080 (N_17080,N_14043,N_12576);
or U17081 (N_17081,N_14152,N_14431);
nor U17082 (N_17082,N_14079,N_12546);
nor U17083 (N_17083,N_14654,N_15736);
nor U17084 (N_17084,N_15801,N_14261);
or U17085 (N_17085,N_12151,N_15707);
or U17086 (N_17086,N_13418,N_14490);
and U17087 (N_17087,N_14299,N_13171);
or U17088 (N_17088,N_13343,N_13012);
xor U17089 (N_17089,N_12729,N_14058);
nor U17090 (N_17090,N_12313,N_13609);
or U17091 (N_17091,N_13449,N_12533);
and U17092 (N_17092,N_15950,N_14395);
xor U17093 (N_17093,N_13230,N_14335);
xnor U17094 (N_17094,N_12415,N_15387);
nand U17095 (N_17095,N_12661,N_13088);
nor U17096 (N_17096,N_13078,N_15706);
xnor U17097 (N_17097,N_12909,N_13762);
xor U17098 (N_17098,N_14274,N_13286);
nor U17099 (N_17099,N_14019,N_15877);
and U17100 (N_17100,N_14273,N_15835);
and U17101 (N_17101,N_15883,N_14868);
and U17102 (N_17102,N_12766,N_12935);
nand U17103 (N_17103,N_15052,N_14242);
nor U17104 (N_17104,N_12106,N_14704);
or U17105 (N_17105,N_14813,N_15785);
or U17106 (N_17106,N_14783,N_15716);
xnor U17107 (N_17107,N_13439,N_12384);
xnor U17108 (N_17108,N_15449,N_15984);
and U17109 (N_17109,N_13995,N_14657);
or U17110 (N_17110,N_15838,N_13440);
and U17111 (N_17111,N_14607,N_14429);
xor U17112 (N_17112,N_12249,N_12210);
and U17113 (N_17113,N_13390,N_15551);
nand U17114 (N_17114,N_14966,N_14089);
or U17115 (N_17115,N_15523,N_14582);
nand U17116 (N_17116,N_14809,N_12630);
and U17117 (N_17117,N_14397,N_13268);
xnor U17118 (N_17118,N_12596,N_12230);
nand U17119 (N_17119,N_15250,N_12481);
xor U17120 (N_17120,N_12265,N_13044);
nand U17121 (N_17121,N_13892,N_15090);
or U17122 (N_17122,N_15170,N_15102);
and U17123 (N_17123,N_15773,N_13837);
and U17124 (N_17124,N_15580,N_15939);
nor U17125 (N_17125,N_15675,N_12980);
and U17126 (N_17126,N_14906,N_15340);
nand U17127 (N_17127,N_14548,N_12116);
or U17128 (N_17128,N_14578,N_15357);
or U17129 (N_17129,N_12060,N_14419);
xor U17130 (N_17130,N_14123,N_15945);
nand U17131 (N_17131,N_14432,N_15727);
and U17132 (N_17132,N_14211,N_14991);
or U17133 (N_17133,N_13933,N_13294);
nand U17134 (N_17134,N_15510,N_12624);
nand U17135 (N_17135,N_14090,N_15167);
or U17136 (N_17136,N_12541,N_12967);
or U17137 (N_17137,N_13437,N_14193);
and U17138 (N_17138,N_13249,N_12494);
xnor U17139 (N_17139,N_14751,N_15594);
xnor U17140 (N_17140,N_15133,N_15329);
or U17141 (N_17141,N_13362,N_14145);
and U17142 (N_17142,N_13202,N_15316);
or U17143 (N_17143,N_13031,N_15243);
xor U17144 (N_17144,N_15485,N_14605);
xnor U17145 (N_17145,N_15431,N_15846);
nand U17146 (N_17146,N_12499,N_13597);
or U17147 (N_17147,N_13640,N_13019);
or U17148 (N_17148,N_15768,N_12878);
or U17149 (N_17149,N_12934,N_14989);
nand U17150 (N_17150,N_12263,N_13434);
or U17151 (N_17151,N_13948,N_12779);
xor U17152 (N_17152,N_14170,N_14215);
nor U17153 (N_17153,N_15684,N_12600);
or U17154 (N_17154,N_12336,N_12347);
or U17155 (N_17155,N_15461,N_13475);
nor U17156 (N_17156,N_14631,N_14282);
nor U17157 (N_17157,N_13036,N_15195);
xor U17158 (N_17158,N_15072,N_13246);
nand U17159 (N_17159,N_12252,N_15622);
and U17160 (N_17160,N_12672,N_13738);
and U17161 (N_17161,N_12196,N_14747);
nor U17162 (N_17162,N_12461,N_14158);
nand U17163 (N_17163,N_13966,N_12467);
or U17164 (N_17164,N_13730,N_14070);
nand U17165 (N_17165,N_15504,N_15259);
or U17166 (N_17166,N_14313,N_13155);
xor U17167 (N_17167,N_12503,N_12314);
and U17168 (N_17168,N_12629,N_12018);
xor U17169 (N_17169,N_15295,N_12803);
xor U17170 (N_17170,N_14916,N_15907);
xnor U17171 (N_17171,N_13960,N_12247);
and U17172 (N_17172,N_15888,N_13577);
xnor U17173 (N_17173,N_12211,N_15249);
or U17174 (N_17174,N_13628,N_15602);
or U17175 (N_17175,N_15088,N_13862);
nor U17176 (N_17176,N_15345,N_14807);
xor U17177 (N_17177,N_13135,N_12167);
and U17178 (N_17178,N_14986,N_15512);
nor U17179 (N_17179,N_12326,N_15501);
nor U17180 (N_17180,N_14937,N_14286);
xor U17181 (N_17181,N_12574,N_14681);
or U17182 (N_17182,N_14788,N_13768);
nand U17183 (N_17183,N_15963,N_13709);
or U17184 (N_17184,N_15795,N_13258);
xnor U17185 (N_17185,N_15065,N_15988);
and U17186 (N_17186,N_14214,N_13293);
nor U17187 (N_17187,N_14589,N_13899);
xor U17188 (N_17188,N_13914,N_12988);
and U17189 (N_17189,N_12545,N_13828);
xor U17190 (N_17190,N_13852,N_15539);
and U17191 (N_17191,N_15266,N_14227);
nor U17192 (N_17192,N_12275,N_13131);
xor U17193 (N_17193,N_13767,N_14181);
nand U17194 (N_17194,N_14764,N_15047);
or U17195 (N_17195,N_13649,N_12219);
or U17196 (N_17196,N_14304,N_15609);
nand U17197 (N_17197,N_14626,N_15192);
nand U17198 (N_17198,N_12825,N_12694);
or U17199 (N_17199,N_14692,N_12912);
and U17200 (N_17200,N_12284,N_15505);
nand U17201 (N_17201,N_14449,N_12834);
nor U17202 (N_17202,N_13598,N_13454);
nor U17203 (N_17203,N_14141,N_14566);
xnor U17204 (N_17204,N_14379,N_13041);
nand U17205 (N_17205,N_15614,N_13868);
and U17206 (N_17206,N_12328,N_15186);
nor U17207 (N_17207,N_13336,N_14667);
xor U17208 (N_17208,N_14239,N_14877);
and U17209 (N_17209,N_13196,N_14129);
xnor U17210 (N_17210,N_14640,N_15715);
and U17211 (N_17211,N_14773,N_12844);
and U17212 (N_17212,N_12964,N_13141);
and U17213 (N_17213,N_14623,N_14703);
nand U17214 (N_17214,N_13526,N_12385);
or U17215 (N_17215,N_12086,N_14498);
nor U17216 (N_17216,N_15370,N_14602);
and U17217 (N_17217,N_12679,N_13427);
nand U17218 (N_17218,N_13332,N_12281);
nor U17219 (N_17219,N_15492,N_15049);
and U17220 (N_17220,N_14336,N_15725);
and U17221 (N_17221,N_12940,N_15438);
nand U17222 (N_17222,N_15755,N_13305);
and U17223 (N_17223,N_12806,N_13620);
nand U17224 (N_17224,N_13456,N_14031);
xnor U17225 (N_17225,N_12109,N_14557);
xor U17226 (N_17226,N_12862,N_15077);
or U17227 (N_17227,N_12510,N_13409);
nand U17228 (N_17228,N_12761,N_13295);
and U17229 (N_17229,N_15726,N_13461);
nand U17230 (N_17230,N_13863,N_12504);
xor U17231 (N_17231,N_14875,N_14080);
xnor U17232 (N_17232,N_13648,N_15285);
or U17233 (N_17233,N_15587,N_15679);
xnor U17234 (N_17234,N_14009,N_15989);
or U17235 (N_17235,N_14608,N_15645);
and U17236 (N_17236,N_13183,N_13866);
nand U17237 (N_17237,N_13802,N_14632);
nor U17238 (N_17238,N_14463,N_15986);
nor U17239 (N_17239,N_15799,N_15881);
nand U17240 (N_17240,N_13680,N_13255);
and U17241 (N_17241,N_14649,N_12659);
xnor U17242 (N_17242,N_15335,N_13683);
nand U17243 (N_17243,N_14110,N_12189);
or U17244 (N_17244,N_15247,N_14376);
nor U17245 (N_17245,N_14825,N_12900);
or U17246 (N_17246,N_12899,N_12135);
nor U17247 (N_17247,N_12155,N_15129);
xnor U17248 (N_17248,N_12452,N_13372);
or U17249 (N_17249,N_12740,N_12607);
or U17250 (N_17250,N_12107,N_13407);
xor U17251 (N_17251,N_14882,N_13774);
xnor U17252 (N_17252,N_14823,N_15481);
nand U17253 (N_17253,N_13859,N_13714);
nand U17254 (N_17254,N_14369,N_13422);
and U17255 (N_17255,N_14120,N_15314);
or U17256 (N_17256,N_15601,N_14456);
nor U17257 (N_17257,N_14822,N_12300);
and U17258 (N_17258,N_13693,N_14671);
xnor U17259 (N_17259,N_13050,N_15109);
and U17260 (N_17260,N_12933,N_12925);
and U17261 (N_17261,N_14205,N_15666);
or U17262 (N_17262,N_12587,N_15804);
nor U17263 (N_17263,N_12905,N_12635);
xor U17264 (N_17264,N_15526,N_14697);
xor U17265 (N_17265,N_14386,N_15222);
nor U17266 (N_17266,N_14371,N_12704);
or U17267 (N_17267,N_15177,N_14351);
nand U17268 (N_17268,N_12074,N_14918);
nor U17269 (N_17269,N_13740,N_15298);
nand U17270 (N_17270,N_12236,N_12386);
nor U17271 (N_17271,N_14855,N_12255);
or U17272 (N_17272,N_12947,N_12082);
and U17273 (N_17273,N_13544,N_12822);
xor U17274 (N_17274,N_15256,N_15124);
nand U17275 (N_17275,N_15344,N_14157);
or U17276 (N_17276,N_14014,N_12363);
and U17277 (N_17277,N_12456,N_12432);
and U17278 (N_17278,N_14087,N_14987);
and U17279 (N_17279,N_15852,N_13561);
nor U17280 (N_17280,N_13679,N_12172);
and U17281 (N_17281,N_13353,N_13032);
xor U17282 (N_17282,N_15302,N_13573);
nor U17283 (N_17283,N_12898,N_15474);
and U17284 (N_17284,N_14797,N_12061);
and U17285 (N_17285,N_12228,N_13182);
and U17286 (N_17286,N_15066,N_12411);
nand U17287 (N_17287,N_13033,N_14347);
nand U17288 (N_17288,N_14295,N_13136);
xnor U17289 (N_17289,N_13578,N_14545);
nor U17290 (N_17290,N_15002,N_15011);
nor U17291 (N_17291,N_13816,N_12000);
xnor U17292 (N_17292,N_15942,N_15254);
or U17293 (N_17293,N_15894,N_12406);
or U17294 (N_17294,N_15748,N_13145);
nor U17295 (N_17295,N_13610,N_15201);
nand U17296 (N_17296,N_12118,N_14482);
nand U17297 (N_17297,N_13501,N_13297);
or U17298 (N_17298,N_14839,N_13453);
xnor U17299 (N_17299,N_12906,N_15629);
nor U17300 (N_17300,N_14569,N_14175);
and U17301 (N_17301,N_12098,N_15003);
nor U17302 (N_17302,N_15337,N_12549);
xor U17303 (N_17303,N_12193,N_15400);
and U17304 (N_17304,N_13678,N_15875);
xor U17305 (N_17305,N_14139,N_13010);
or U17306 (N_17306,N_14794,N_15188);
xor U17307 (N_17307,N_13159,N_15925);
nor U17308 (N_17308,N_12928,N_14724);
nor U17309 (N_17309,N_14913,N_15452);
and U17310 (N_17310,N_13225,N_14240);
nand U17311 (N_17311,N_12147,N_12554);
or U17312 (N_17312,N_15660,N_15118);
nor U17313 (N_17313,N_13463,N_13786);
xor U17314 (N_17314,N_13113,N_14478);
xnor U17315 (N_17315,N_12091,N_12261);
or U17316 (N_17316,N_13219,N_14316);
xnor U17317 (N_17317,N_14314,N_12241);
nand U17318 (N_17318,N_14334,N_15071);
nand U17319 (N_17319,N_14900,N_15586);
xnor U17320 (N_17320,N_15570,N_15685);
xnor U17321 (N_17321,N_13752,N_15900);
xor U17322 (N_17322,N_14818,N_14942);
or U17323 (N_17323,N_14617,N_15831);
xnor U17324 (N_17324,N_14934,N_13315);
xnor U17325 (N_17325,N_15763,N_14342);
or U17326 (N_17326,N_14438,N_14246);
nand U17327 (N_17327,N_14249,N_15191);
xnor U17328 (N_17328,N_13029,N_13348);
nand U17329 (N_17329,N_13826,N_12418);
xnor U17330 (N_17330,N_12859,N_12902);
nand U17331 (N_17331,N_13369,N_12201);
or U17332 (N_17332,N_14609,N_15871);
or U17333 (N_17333,N_14804,N_13723);
and U17334 (N_17334,N_15787,N_12030);
xor U17335 (N_17335,N_14167,N_12792);
nand U17336 (N_17336,N_14576,N_12272);
nor U17337 (N_17337,N_15148,N_14963);
xor U17338 (N_17338,N_14676,N_14284);
nand U17339 (N_17339,N_15948,N_13504);
nand U17340 (N_17340,N_13910,N_13992);
nor U17341 (N_17341,N_12525,N_12278);
nand U17342 (N_17342,N_12059,N_12120);
or U17343 (N_17343,N_12359,N_13865);
xnor U17344 (N_17344,N_14136,N_14025);
xnor U17345 (N_17345,N_14993,N_15855);
and U17346 (N_17346,N_15166,N_15032);
xnor U17347 (N_17347,N_13505,N_14095);
xor U17348 (N_17348,N_14673,N_15653);
and U17349 (N_17349,N_14945,N_14000);
and U17350 (N_17350,N_14457,N_14469);
or U17351 (N_17351,N_14816,N_14069);
nand U17352 (N_17352,N_13172,N_12751);
and U17353 (N_17353,N_14833,N_14178);
nand U17354 (N_17354,N_12843,N_14310);
or U17355 (N_17355,N_12580,N_13690);
and U17356 (N_17356,N_14470,N_13660);
or U17357 (N_17357,N_14976,N_13181);
xnor U17358 (N_17358,N_15226,N_14994);
nand U17359 (N_17359,N_12477,N_13263);
xor U17360 (N_17360,N_14741,N_13676);
and U17361 (N_17361,N_12712,N_13000);
nor U17362 (N_17362,N_13340,N_12956);
and U17363 (N_17363,N_13082,N_13665);
or U17364 (N_17364,N_12126,N_12974);
xor U17365 (N_17365,N_15776,N_12310);
nor U17366 (N_17366,N_12383,N_15847);
nor U17367 (N_17367,N_13400,N_15498);
and U17368 (N_17368,N_13824,N_15574);
nor U17369 (N_17369,N_13787,N_12973);
xnor U17370 (N_17370,N_14108,N_15688);
nor U17371 (N_17371,N_14910,N_12289);
nand U17372 (N_17372,N_13954,N_13331);
or U17373 (N_17373,N_13976,N_13694);
or U17374 (N_17374,N_12791,N_13274);
or U17375 (N_17375,N_13392,N_15307);
or U17376 (N_17376,N_13627,N_13978);
or U17377 (N_17377,N_13494,N_15383);
nor U17378 (N_17378,N_14187,N_13527);
xor U17379 (N_17379,N_13823,N_12670);
or U17380 (N_17380,N_13765,N_15334);
nor U17381 (N_17381,N_15784,N_12692);
and U17382 (N_17382,N_12209,N_13112);
xnor U17383 (N_17383,N_12258,N_12004);
xnor U17384 (N_17384,N_15160,N_15179);
or U17385 (N_17385,N_15511,N_14027);
nand U17386 (N_17386,N_14156,N_13796);
nor U17387 (N_17387,N_12713,N_13290);
or U17388 (N_17388,N_15994,N_12200);
or U17389 (N_17389,N_13584,N_15127);
or U17390 (N_17390,N_15108,N_14529);
or U17391 (N_17391,N_13968,N_14276);
xor U17392 (N_17392,N_14659,N_13391);
nand U17393 (N_17393,N_14830,N_13244);
nor U17394 (N_17394,N_14613,N_13599);
nor U17395 (N_17395,N_14445,N_12270);
nor U17396 (N_17396,N_15596,N_15242);
xnor U17397 (N_17397,N_15612,N_12564);
nand U17398 (N_17398,N_12943,N_13719);
nor U17399 (N_17399,N_14701,N_13616);
xnor U17400 (N_17400,N_14385,N_13930);
xnor U17401 (N_17401,N_12722,N_12568);
xor U17402 (N_17402,N_14190,N_14573);
nand U17403 (N_17403,N_13568,N_12444);
or U17404 (N_17404,N_15116,N_15121);
nand U17405 (N_17405,N_14912,N_14684);
xor U17406 (N_17406,N_12315,N_15825);
nand U17407 (N_17407,N_14191,N_13896);
xor U17408 (N_17408,N_12096,N_12759);
and U17409 (N_17409,N_14718,N_15395);
nor U17410 (N_17410,N_13188,N_12614);
xnor U17411 (N_17411,N_15086,N_15025);
or U17412 (N_17412,N_12777,N_15772);
or U17413 (N_17413,N_12976,N_15884);
nor U17414 (N_17414,N_13177,N_13507);
and U17415 (N_17415,N_12968,N_15968);
nand U17416 (N_17416,N_12320,N_15598);
nand U17417 (N_17417,N_12125,N_14326);
or U17418 (N_17418,N_12215,N_13022);
nor U17419 (N_17419,N_14106,N_13755);
and U17420 (N_17420,N_13817,N_12835);
or U17421 (N_17421,N_15573,N_12309);
and U17422 (N_17422,N_12259,N_12409);
nor U17423 (N_17423,N_15194,N_12413);
or U17424 (N_17424,N_15841,N_12188);
nor U17425 (N_17425,N_12355,N_12054);
nor U17426 (N_17426,N_14543,N_13066);
nand U17427 (N_17427,N_12769,N_12009);
xnor U17428 (N_17428,N_13308,N_13595);
or U17429 (N_17429,N_13042,N_14668);
xnor U17430 (N_17430,N_15652,N_14140);
and U17431 (N_17431,N_14195,N_14360);
nor U17432 (N_17432,N_15980,N_15506);
and U17433 (N_17433,N_15402,N_15394);
nand U17434 (N_17434,N_13097,N_14099);
and U17435 (N_17435,N_13835,N_12260);
nand U17436 (N_17436,N_14637,N_12380);
and U17437 (N_17437,N_13147,N_12937);
and U17438 (N_17438,N_15771,N_15954);
and U17439 (N_17439,N_15459,N_12003);
nor U17440 (N_17440,N_13452,N_15069);
nor U17441 (N_17441,N_13500,N_13925);
nand U17442 (N_17442,N_13166,N_14720);
and U17443 (N_17443,N_13430,N_15646);
nor U17444 (N_17444,N_12005,N_15951);
nand U17445 (N_17445,N_12886,N_14082);
nor U17446 (N_17446,N_14558,N_15215);
nor U17447 (N_17447,N_13361,N_15837);
nand U17448 (N_17448,N_15802,N_15863);
nor U17449 (N_17449,N_13433,N_14544);
or U17450 (N_17450,N_13559,N_12911);
nand U17451 (N_17451,N_13651,N_13623);
nand U17452 (N_17452,N_15738,N_12293);
and U17453 (N_17453,N_14997,N_13317);
and U17454 (N_17454,N_15187,N_12784);
or U17455 (N_17455,N_13282,N_15563);
xnor U17456 (N_17456,N_12194,N_13795);
xnor U17457 (N_17457,N_15991,N_12280);
or U17458 (N_17458,N_15348,N_15541);
xor U17459 (N_17459,N_14093,N_15123);
or U17460 (N_17460,N_14317,N_12097);
nand U17461 (N_17461,N_15360,N_13630);
nand U17462 (N_17462,N_13843,N_14337);
or U17463 (N_17463,N_13766,N_14590);
nand U17464 (N_17464,N_15364,N_13090);
and U17465 (N_17465,N_13248,N_15022);
or U17466 (N_17466,N_12417,N_12972);
xnor U17467 (N_17467,N_12441,N_15053);
and U17468 (N_17468,N_13617,N_13895);
nand U17469 (N_17469,N_12486,N_14017);
xor U17470 (N_17470,N_14013,N_15517);
nand U17471 (N_17471,N_13243,N_13328);
xor U17472 (N_17472,N_14200,N_15472);
or U17473 (N_17473,N_13015,N_12493);
xnor U17474 (N_17474,N_13856,N_12216);
nand U17475 (N_17475,N_12536,N_12400);
nor U17476 (N_17476,N_15600,N_12425);
and U17477 (N_17477,N_13799,N_14776);
nand U17478 (N_17478,N_14541,N_13313);
nor U17479 (N_17479,N_14928,N_13116);
or U17480 (N_17480,N_12451,N_13037);
nand U17481 (N_17481,N_12856,N_15415);
nor U17482 (N_17482,N_13820,N_12431);
or U17483 (N_17483,N_13841,N_15722);
xor U17484 (N_17484,N_14852,N_12232);
nand U17485 (N_17485,N_13564,N_15112);
nor U17486 (N_17486,N_14740,N_15209);
and U17487 (N_17487,N_14107,N_12066);
and U17488 (N_17488,N_13068,N_15607);
nand U17489 (N_17489,N_14117,N_12879);
or U17490 (N_17490,N_14982,N_12852);
and U17491 (N_17491,N_12286,N_15331);
xnor U17492 (N_17492,N_13614,N_14898);
xnor U17493 (N_17493,N_14307,N_15322);
or U17494 (N_17494,N_12110,N_14939);
nor U17495 (N_17495,N_13977,N_15487);
nand U17496 (N_17496,N_13625,N_15817);
nor U17497 (N_17497,N_12458,N_12571);
xor U17498 (N_17498,N_14023,N_12153);
or U17499 (N_17499,N_14088,N_14345);
nor U17500 (N_17500,N_15576,N_12688);
nor U17501 (N_17501,N_14266,N_14919);
nand U17502 (N_17502,N_13377,N_14072);
xor U17503 (N_17503,N_15542,N_14306);
or U17504 (N_17504,N_14748,N_14630);
nand U17505 (N_17505,N_14857,N_15475);
or U17506 (N_17506,N_13408,N_12181);
or U17507 (N_17507,N_13989,N_14824);
xor U17508 (N_17508,N_14860,N_13569);
and U17509 (N_17509,N_14904,N_12881);
xnor U17510 (N_17510,N_15648,N_15922);
or U17511 (N_17511,N_15965,N_13239);
or U17512 (N_17512,N_14629,N_13156);
nand U17513 (N_17513,N_15906,N_15640);
and U17514 (N_17514,N_14821,N_12817);
and U17515 (N_17515,N_12433,N_13233);
nor U17516 (N_17516,N_14542,N_12556);
nor U17517 (N_17517,N_12702,N_15274);
or U17518 (N_17518,N_12042,N_12609);
nor U17519 (N_17519,N_14415,N_12985);
xnor U17520 (N_17520,N_14620,N_12298);
nand U17521 (N_17521,N_14546,N_12366);
nand U17522 (N_17522,N_12962,N_12373);
nor U17523 (N_17523,N_15741,N_13745);
or U17524 (N_17524,N_13981,N_14929);
and U17525 (N_17525,N_12622,N_13506);
or U17526 (N_17526,N_13904,N_12894);
nor U17527 (N_17527,N_13385,N_15760);
nor U17528 (N_17528,N_13801,N_15227);
nor U17529 (N_17529,N_14403,N_15378);
xnor U17530 (N_17530,N_12489,N_15836);
xor U17531 (N_17531,N_14416,N_13376);
or U17532 (N_17532,N_13071,N_13860);
or U17533 (N_17533,N_14037,N_12346);
and U17534 (N_17534,N_15418,N_14414);
and U17535 (N_17535,N_12338,N_15045);
or U17536 (N_17536,N_13653,N_14579);
and U17537 (N_17537,N_15440,N_15509);
and U17538 (N_17538,N_12775,N_12582);
or U17539 (N_17539,N_15202,N_13395);
xnor U17540 (N_17540,N_12323,N_13296);
and U17541 (N_17541,N_13945,N_15717);
nor U17542 (N_17542,N_14820,N_15330);
and U17543 (N_17543,N_13917,N_14111);
nand U17544 (N_17544,N_12750,N_13601);
nand U17545 (N_17545,N_15044,N_14842);
xnor U17546 (N_17546,N_15901,N_12382);
nand U17547 (N_17547,N_12427,N_13728);
xnor U17548 (N_17548,N_13715,N_14413);
or U17549 (N_17549,N_12871,N_12977);
nor U17550 (N_17550,N_14280,N_12022);
nand U17551 (N_17551,N_14638,N_13612);
nand U17552 (N_17552,N_14226,N_13798);
xnor U17553 (N_17553,N_13271,N_15271);
and U17554 (N_17554,N_13855,N_12368);
nand U17555 (N_17555,N_13725,N_14695);
nor U17556 (N_17556,N_15239,N_12065);
or U17557 (N_17557,N_13176,N_15697);
nand U17558 (N_17558,N_12632,N_15445);
and U17559 (N_17559,N_12677,N_12774);
nand U17560 (N_17560,N_13562,N_12697);
and U17561 (N_17561,N_14990,N_13636);
xnor U17562 (N_17562,N_13808,N_13546);
nor U17563 (N_17563,N_12222,N_14960);
nand U17564 (N_17564,N_13479,N_13631);
or U17565 (N_17565,N_14921,N_12760);
xor U17566 (N_17566,N_14612,N_12866);
or U17567 (N_17567,N_13358,N_14591);
nor U17568 (N_17568,N_15742,N_12470);
and U17569 (N_17569,N_14030,N_13792);
nand U17570 (N_17570,N_14853,N_15815);
and U17571 (N_17571,N_15764,N_12246);
nand U17572 (N_17572,N_15385,N_14443);
nand U17573 (N_17573,N_14556,N_13151);
nor U17574 (N_17574,N_15844,N_13939);
and U17575 (N_17575,N_13514,N_15605);
and U17576 (N_17576,N_14614,N_14520);
xnor U17577 (N_17577,N_12524,N_13416);
nor U17578 (N_17578,N_12062,N_12269);
xor U17579 (N_17579,N_14479,N_15829);
or U17580 (N_17580,N_12741,N_13227);
and U17581 (N_17581,N_12087,N_12837);
or U17582 (N_17582,N_12206,N_15444);
and U17583 (N_17583,N_15993,N_12378);
nand U17584 (N_17584,N_14380,N_14154);
nand U17585 (N_17585,N_15294,N_12213);
and U17586 (N_17586,N_14256,N_14220);
nand U17587 (N_17587,N_12828,N_15750);
xnor U17588 (N_17588,N_14812,N_14968);
and U17589 (N_17589,N_14378,N_14237);
nor U17590 (N_17590,N_15356,N_13664);
xnor U17591 (N_17591,N_14599,N_13818);
and U17592 (N_17592,N_15543,N_15562);
nor U17593 (N_17593,N_12655,N_13938);
and U17594 (N_17594,N_14728,N_12544);
nor U17595 (N_17595,N_15694,N_12563);
xor U17596 (N_17596,N_15396,N_14936);
nor U17597 (N_17597,N_13017,N_12660);
or U17598 (N_17598,N_12237,N_14298);
and U17599 (N_17599,N_15406,N_14437);
nor U17600 (N_17600,N_13163,N_12875);
or U17601 (N_17601,N_13832,N_15973);
or U17602 (N_17602,N_13417,N_14118);
and U17603 (N_17603,N_12291,N_13345);
xnor U17604 (N_17604,N_15467,N_12783);
xor U17605 (N_17605,N_14536,N_12727);
and U17606 (N_17606,N_13713,N_15637);
and U17607 (N_17607,N_13164,N_14029);
nor U17608 (N_17608,N_12598,N_12924);
nor U17609 (N_17609,N_15275,N_14216);
and U17610 (N_17610,N_14001,N_12229);
and U17611 (N_17611,N_14404,N_15743);
or U17612 (N_17612,N_13186,N_13909);
or U17613 (N_17613,N_13211,N_13161);
or U17614 (N_17614,N_12731,N_14398);
nor U17615 (N_17615,N_14760,N_13443);
nor U17616 (N_17616,N_15870,N_12641);
nand U17617 (N_17617,N_13216,N_14635);
xnor U17618 (N_17618,N_14905,N_14077);
xor U17619 (N_17619,N_15535,N_14253);
nand U17620 (N_17620,N_14207,N_12014);
xor U17621 (N_17621,N_15391,N_14444);
xor U17622 (N_17622,N_12132,N_15962);
nand U17623 (N_17623,N_12407,N_12394);
nor U17624 (N_17624,N_14772,N_12304);
xor U17625 (N_17625,N_14849,N_15552);
xnor U17626 (N_17626,N_15774,N_15236);
and U17627 (N_17627,N_12921,N_12771);
or U17628 (N_17628,N_14320,N_12983);
nor U17629 (N_17629,N_12948,N_14869);
or U17630 (N_17630,N_15094,N_12667);
and U17631 (N_17631,N_13883,N_15351);
nand U17632 (N_17632,N_14743,N_13810);
nor U17633 (N_17633,N_14909,N_15651);
nor U17634 (N_17634,N_13528,N_13854);
or U17635 (N_17635,N_12789,N_13126);
or U17636 (N_17636,N_14735,N_15941);
or U17637 (N_17637,N_15828,N_15955);
nor U17638 (N_17638,N_14308,N_12321);
xor U17639 (N_17639,N_15233,N_13842);
or U17640 (N_17640,N_12681,N_15923);
nand U17641 (N_17641,N_13594,N_14938);
and U17642 (N_17642,N_13123,N_14595);
or U17643 (N_17643,N_13775,N_15327);
nand U17644 (N_17644,N_15352,N_15692);
nor U17645 (N_17645,N_13492,N_14914);
or U17646 (N_17646,N_15310,N_13178);
nor U17647 (N_17647,N_12352,N_15164);
nand U17648 (N_17648,N_15695,N_14285);
and U17649 (N_17649,N_13951,N_15749);
nand U17650 (N_17650,N_15031,N_15561);
nor U17651 (N_17651,N_15718,N_12047);
xor U17652 (N_17652,N_12509,N_12485);
and U17653 (N_17653,N_12845,N_14480);
nand U17654 (N_17654,N_15379,N_13580);
nand U17655 (N_17655,N_14555,N_14050);
nand U17656 (N_17656,N_15386,N_13005);
nor U17657 (N_17657,N_14328,N_13428);
xor U17658 (N_17658,N_13337,N_14650);
xnor U17659 (N_17659,N_12555,N_14656);
and U17660 (N_17660,N_12711,N_13104);
xnor U17661 (N_17661,N_14522,N_13318);
xnor U17662 (N_17662,N_12114,N_13414);
xor U17663 (N_17663,N_14488,N_12104);
or U17664 (N_17664,N_12350,N_12187);
nand U17665 (N_17665,N_12442,N_14570);
nor U17666 (N_17666,N_13048,N_15339);
xor U17667 (N_17667,N_12665,N_14461);
nand U17668 (N_17668,N_13535,N_12220);
xor U17669 (N_17669,N_13167,N_12290);
and U17670 (N_17670,N_14056,N_13667);
or U17671 (N_17671,N_12599,N_13208);
nor U17672 (N_17672,N_15669,N_15797);
xnor U17673 (N_17673,N_14229,N_12831);
nor U17674 (N_17674,N_14439,N_12847);
or U17675 (N_17675,N_14255,N_14716);
nor U17676 (N_17676,N_15493,N_13143);
nand U17677 (N_17677,N_14235,N_12202);
or U17678 (N_17678,N_13606,N_15654);
and U17679 (N_17679,N_13153,N_13024);
xor U17680 (N_17680,N_13281,N_13994);
and U17681 (N_17681,N_12311,N_13081);
xnor U17682 (N_17682,N_14935,N_13971);
and U17683 (N_17683,N_13047,N_12064);
nor U17684 (N_17684,N_13252,N_13462);
nand U17685 (N_17685,N_15457,N_12616);
nand U17686 (N_17686,N_14858,N_14744);
nand U17687 (N_17687,N_13662,N_15926);
nor U17688 (N_17688,N_14194,N_12371);
xor U17689 (N_17689,N_15572,N_13447);
nor U17690 (N_17690,N_12888,N_12548);
nand U17691 (N_17691,N_14730,N_15872);
and U17692 (N_17692,N_12786,N_13756);
nor U17693 (N_17693,N_12144,N_12724);
nand U17694 (N_17694,N_13687,N_13404);
nand U17695 (N_17695,N_13469,N_15122);
xor U17696 (N_17696,N_15206,N_14428);
xnor U17697 (N_17697,N_15260,N_13067);
or U17698 (N_17698,N_15752,N_12827);
or U17699 (N_17699,N_15269,N_15610);
or U17700 (N_17700,N_15940,N_14092);
and U17701 (N_17701,N_15865,N_15759);
xor U17702 (N_17702,N_13581,N_14430);
and U17703 (N_17703,N_15515,N_12945);
xnor U17704 (N_17704,N_13060,N_15479);
nor U17705 (N_17705,N_13912,N_13847);
nand U17706 (N_17706,N_14180,N_12836);
nor U17707 (N_17707,N_13585,N_14387);
nand U17708 (N_17708,N_15091,N_12372);
xnor U17709 (N_17709,N_15904,N_13320);
nand U17710 (N_17710,N_14132,N_14467);
or U17711 (N_17711,N_12402,N_15137);
and U17712 (N_17712,N_15373,N_13661);
and U17713 (N_17713,N_15325,N_12070);
xnor U17714 (N_17714,N_12318,N_15516);
or U17715 (N_17715,N_13021,N_14206);
nor U17716 (N_17716,N_15321,N_12892);
nand U17717 (N_17717,N_12590,N_14494);
xor U17718 (N_17718,N_13695,N_12245);
xnor U17719 (N_17719,N_12780,N_13764);
nand U17720 (N_17720,N_15514,N_13330);
xor U17721 (N_17721,N_15278,N_14661);
nand U17722 (N_17722,N_13124,N_13878);
nor U17723 (N_17723,N_13888,N_15424);
xor U17724 (N_17724,N_15436,N_13215);
nand U17725 (N_17725,N_12161,N_14847);
or U17726 (N_17726,N_15701,N_14433);
and U17727 (N_17727,N_14694,N_15703);
and U17728 (N_17728,N_14401,N_14420);
or U17729 (N_17729,N_15354,N_15035);
xnor U17730 (N_17730,N_12941,N_12913);
nand U17731 (N_17731,N_15130,N_14600);
or U17732 (N_17732,N_12529,N_14497);
and U17733 (N_17733,N_13645,N_12397);
xor U17734 (N_17734,N_14507,N_13590);
xnor U17735 (N_17735,N_14777,N_14970);
nand U17736 (N_17736,N_15414,N_12016);
nor U17737 (N_17737,N_15039,N_14210);
xor U17738 (N_17738,N_13114,N_12957);
or U17739 (N_17739,N_12464,N_14374);
and U17740 (N_17740,N_14130,N_15628);
nor U17741 (N_17741,N_15001,N_13079);
or U17742 (N_17742,N_12954,N_13591);
nand U17743 (N_17743,N_14361,N_15174);
xnor U17744 (N_17744,N_12081,N_15282);
or U17745 (N_17745,N_12790,N_13997);
and U17746 (N_17746,N_12768,N_13476);
or U17747 (N_17747,N_12438,N_12527);
nor U17748 (N_17748,N_15834,N_13319);
nand U17749 (N_17749,N_13169,N_12959);
nand U17750 (N_17750,N_12039,N_12809);
nor U17751 (N_17751,N_15204,N_13919);
nor U17752 (N_17752,N_14572,N_15397);
xor U17753 (N_17753,N_13560,N_15147);
nand U17754 (N_17754,N_15664,N_13975);
and U17755 (N_17755,N_12362,N_12393);
nand U17756 (N_17756,N_14961,N_14827);
nor U17757 (N_17757,N_13692,N_15818);
or U17758 (N_17758,N_13483,N_14396);
xor U17759 (N_17759,N_14948,N_14039);
and U17760 (N_17760,N_14931,N_12796);
xnor U17761 (N_17761,N_13790,N_13478);
and U17762 (N_17762,N_12340,N_14048);
or U17763 (N_17763,N_14851,N_15820);
xnor U17764 (N_17764,N_12334,N_14517);
xnor U17765 (N_17765,N_14854,N_15488);
or U17766 (N_17766,N_14758,N_14400);
nand U17767 (N_17767,N_15775,N_12101);
nor U17768 (N_17768,N_14067,N_13748);
and U17769 (N_17769,N_12961,N_13869);
nor U17770 (N_17770,N_13533,N_15555);
nand U17771 (N_17771,N_14038,N_14971);
xor U17772 (N_17772,N_14817,N_15996);
xor U17773 (N_17773,N_14231,N_15620);
or U17774 (N_17774,N_13325,N_15811);
nor U17775 (N_17775,N_12088,N_15796);
or U17776 (N_17776,N_13831,N_13864);
nor U17777 (N_17777,N_12369,N_15558);
nand U17778 (N_17778,N_12420,N_13915);
and U17779 (N_17779,N_14785,N_13618);
or U17780 (N_17780,N_13222,N_15910);
and U17781 (N_17781,N_14066,N_13333);
xnor U17782 (N_17782,N_12993,N_14834);
xnor U17783 (N_17783,N_14981,N_13721);
and U17784 (N_17784,N_12015,N_15183);
and U17785 (N_17785,N_13356,N_12474);
nand U17786 (N_17786,N_15238,N_12197);
or U17787 (N_17787,N_15677,N_13134);
nand U17788 (N_17788,N_14521,N_14941);
or U17789 (N_17789,N_13497,N_12662);
and U17790 (N_17790,N_15372,N_14238);
nand U17791 (N_17791,N_15680,N_12577);
and U17792 (N_17792,N_13875,N_15312);
nor U17793 (N_17793,N_14125,N_12516);
nand U17794 (N_17794,N_12292,N_13157);
nor U17795 (N_17795,N_14790,N_14373);
nand U17796 (N_17796,N_12329,N_12756);
xor U17797 (N_17797,N_15050,N_14837);
nor U17798 (N_17798,N_13524,N_12035);
nor U17799 (N_17799,N_15603,N_15754);
xnor U17800 (N_17800,N_13538,N_13508);
xnor U17801 (N_17801,N_14346,N_12287);
nand U17802 (N_17802,N_14886,N_13420);
nand U17803 (N_17803,N_12111,N_15389);
nand U17804 (N_17804,N_12063,N_13460);
and U17805 (N_17805,N_14465,N_13448);
nand U17806 (N_17806,N_13455,N_14641);
xor U17807 (N_17807,N_13382,N_12140);
and U17808 (N_17808,N_13298,N_12700);
nand U17809 (N_17809,N_14466,N_14126);
and U17810 (N_17810,N_12547,N_13280);
and U17811 (N_17811,N_12730,N_13682);
nand U17812 (N_17812,N_13579,N_13589);
or U17813 (N_17813,N_12903,N_13028);
and U17814 (N_17814,N_15832,N_12701);
or U17815 (N_17815,N_13729,N_12282);
nor U17816 (N_17816,N_15507,N_14262);
nor U17817 (N_17817,N_12920,N_12288);
or U17818 (N_17818,N_14344,N_13004);
or U17819 (N_17819,N_15595,N_15263);
nor U17820 (N_17820,N_14147,N_15218);
and U17821 (N_17821,N_14402,N_14700);
nand U17822 (N_17822,N_14815,N_14885);
and U17823 (N_17823,N_12307,N_14642);
or U17824 (N_17824,N_15858,N_12540);
nor U17825 (N_17825,N_13378,N_13301);
and U17826 (N_17826,N_15843,N_15790);
or U17827 (N_17827,N_13710,N_14260);
or U17828 (N_17828,N_12083,N_15027);
nor U17829 (N_17829,N_14940,N_14375);
nor U17830 (N_17830,N_15650,N_13008);
nor U17831 (N_17831,N_12566,N_12721);
xor U17832 (N_17832,N_12325,N_13209);
nor U17833 (N_17833,N_15223,N_14951);
or U17834 (N_17834,N_13684,N_15977);
nor U17835 (N_17835,N_15012,N_12872);
and U17836 (N_17836,N_14863,N_15432);
nor U17837 (N_17837,N_14561,N_12592);
or U17838 (N_17838,N_12173,N_12496);
and U17839 (N_17839,N_12180,N_13105);
xor U17840 (N_17840,N_13426,N_15532);
nor U17841 (N_17841,N_12317,N_15533);
xnor U17842 (N_17842,N_15769,N_14559);
nand U17843 (N_17843,N_15905,N_13381);
or U17844 (N_17844,N_15349,N_13893);
xor U17845 (N_17845,N_13080,N_14950);
and U17846 (N_17846,N_13073,N_14911);
xnor U17847 (N_17847,N_14634,N_15036);
or U17848 (N_17848,N_13192,N_14955);
nand U17849 (N_17849,N_15674,N_15690);
xor U17850 (N_17850,N_12182,N_14954);
xnor U17851 (N_17851,N_12594,N_12787);
xor U17852 (N_17852,N_15128,N_13003);
xnor U17853 (N_17853,N_12445,N_15245);
nor U17854 (N_17854,N_13160,N_13806);
nand U17855 (N_17855,N_15575,N_12602);
and U17856 (N_17856,N_13425,N_12396);
and U17857 (N_17857,N_15381,N_14340);
nand U17858 (N_17858,N_15714,N_12226);
xor U17859 (N_17859,N_13399,N_14296);
nor U17860 (N_17860,N_14896,N_14459);
and U17861 (N_17861,N_13236,N_13604);
or U17862 (N_17862,N_15676,N_12460);
nand U17863 (N_17863,N_12238,N_12944);
or U17864 (N_17864,N_13779,N_15154);
or U17865 (N_17865,N_13588,N_12308);
nor U17866 (N_17866,N_15184,N_12319);
xnor U17867 (N_17867,N_14513,N_13287);
or U17868 (N_17868,N_12745,N_13269);
nor U17869 (N_17869,N_12166,N_14491);
and U17870 (N_17870,N_14315,N_15297);
and U17871 (N_17871,N_13240,N_14712);
and U17872 (N_17872,N_14892,N_14666);
xor U17873 (N_17873,N_15286,N_12889);
nand U17874 (N_17874,N_15623,N_14664);
nor U17875 (N_17875,N_13110,N_14683);
nor U17876 (N_17876,N_14872,N_15007);
and U17877 (N_17877,N_14440,N_12998);
xnor U17878 (N_17878,N_12550,N_13877);
and U17879 (N_17879,N_12038,N_15111);
nand U17880 (N_17880,N_15593,N_12530);
nor U17881 (N_17881,N_14502,N_14473);
and U17882 (N_17882,N_15704,N_15635);
xor U17883 (N_17883,N_15816,N_13704);
and U17884 (N_17884,N_14071,N_12981);
nor U17885 (N_17885,N_12351,N_15248);
or U17886 (N_17886,N_12778,N_12573);
or U17887 (N_17887,N_14044,N_15377);
and U17888 (N_17888,N_15430,N_13850);
nand U17889 (N_17889,N_15952,N_15521);
nor U17890 (N_17890,N_13702,N_15388);
or U17891 (N_17891,N_12733,N_13373);
nand U17892 (N_17892,N_14956,N_14920);
or U17893 (N_17893,N_13829,N_12224);
nand U17894 (N_17894,N_15896,N_13049);
and U17895 (N_17895,N_12683,N_14418);
or U17896 (N_17896,N_14978,N_12266);
xnor U17897 (N_17897,N_15649,N_14601);
nor U17898 (N_17898,N_12748,N_13237);
xor U17899 (N_17899,N_14587,N_14394);
and U17900 (N_17900,N_15733,N_12519);
nand U17901 (N_17901,N_13881,N_13503);
or U17902 (N_17902,N_13299,N_12810);
or U17903 (N_17903,N_15008,N_12045);
xnor U17904 (N_17904,N_13040,N_13464);
and U17905 (N_17905,N_14277,N_12223);
and U17906 (N_17906,N_14399,N_13450);
xnor U17907 (N_17907,N_15929,N_14693);
nor U17908 (N_17908,N_13214,N_13574);
or U17909 (N_17909,N_15489,N_14263);
nor U17910 (N_17910,N_12316,N_14096);
nor U17911 (N_17911,N_12923,N_15899);
nand U17912 (N_17912,N_12136,N_14643);
nor U17913 (N_17913,N_15104,N_13307);
nand U17914 (N_17914,N_13542,N_13242);
nor U17915 (N_17915,N_14771,N_15663);
xnor U17916 (N_17916,N_15967,N_12267);
nor U17917 (N_17917,N_14798,N_12124);
or U17918 (N_17918,N_13716,N_14204);
nor U17919 (N_17919,N_12572,N_14104);
nor U17920 (N_17920,N_14662,N_15803);
or U17921 (N_17921,N_13419,N_13193);
xor U17922 (N_17922,N_15918,N_13666);
nor U17923 (N_17923,N_12416,N_13670);
and U17924 (N_17924,N_15667,N_13189);
and U17925 (N_17925,N_13998,N_13814);
nor U17926 (N_17926,N_13911,N_14908);
and U17927 (N_17927,N_15520,N_15937);
nand U17928 (N_17928,N_13677,N_13140);
nor U17929 (N_17929,N_12032,N_13051);
nand U17930 (N_17930,N_12019,N_15606);
xor U17931 (N_17931,N_12354,N_13083);
and U17932 (N_17932,N_15048,N_14584);
nor U17933 (N_17933,N_12029,N_13751);
or U17934 (N_17934,N_13973,N_12343);
or U17935 (N_17935,N_12446,N_12262);
and U17936 (N_17936,N_14618,N_13586);
xor U17937 (N_17937,N_14065,N_13034);
xor U17938 (N_17938,N_12253,N_12608);
and U17939 (N_17939,N_14103,N_13168);
nor U17940 (N_17940,N_14933,N_15141);
nand U17941 (N_17941,N_13234,N_12698);
nor U17942 (N_17942,N_14565,N_13052);
xor U17943 (N_17943,N_14793,N_12119);
xor U17944 (N_17944,N_14725,N_13273);
nor U17945 (N_17945,N_12079,N_12389);
and U17946 (N_17946,N_13074,N_15080);
xnor U17947 (N_17947,N_15972,N_14134);
xor U17948 (N_17948,N_14901,N_12031);
or U17949 (N_17949,N_12148,N_12535);
or U17950 (N_17950,N_15478,N_14209);
xnor U17951 (N_17951,N_13962,N_12840);
xor U17952 (N_17952,N_12024,N_12978);
or U17953 (N_17953,N_12613,N_13490);
nand U17954 (N_17954,N_14685,N_13566);
nand U17955 (N_17955,N_12685,N_13095);
and U17956 (N_17956,N_14564,N_14300);
or U17957 (N_17957,N_14979,N_14552);
nor U17958 (N_17958,N_15306,N_12198);
nand U17959 (N_17959,N_15975,N_14133);
and U17960 (N_17960,N_15880,N_13754);
nor U17961 (N_17961,N_15691,N_13570);
xor U17962 (N_17962,N_13763,N_13054);
or U17963 (N_17963,N_13226,N_15630);
nor U17964 (N_17964,N_15181,N_13098);
nand U17965 (N_17965,N_12482,N_12979);
and U17966 (N_17966,N_13944,N_15786);
xnor U17967 (N_17967,N_12377,N_12873);
or U17968 (N_17968,N_12939,N_15304);
nand U17969 (N_17969,N_13894,N_13253);
xor U17970 (N_17970,N_12753,N_15469);
xnor U17971 (N_17971,N_13491,N_12583);
nor U17972 (N_17972,N_13884,N_12850);
and U17973 (N_17973,N_14109,N_14779);
nor U17974 (N_17974,N_14267,N_12922);
and U17975 (N_17975,N_15597,N_13118);
nand U17976 (N_17976,N_12773,N_13554);
and U17977 (N_17977,N_14062,N_14902);
or U17978 (N_17978,N_15599,N_14644);
and U17979 (N_17979,N_14341,N_15564);
nor U17980 (N_17980,N_13920,N_15699);
nand U17981 (N_17981,N_13703,N_12952);
nand U17982 (N_17982,N_12636,N_14845);
nand U17983 (N_17983,N_14421,N_12824);
nand U17984 (N_17984,N_13076,N_15317);
nor U17985 (N_17985,N_14789,N_14604);
xnor U17986 (N_17986,N_12424,N_14042);
and U17987 (N_17987,N_12108,N_13355);
and U17988 (N_17988,N_14848,N_12162);
and U17989 (N_17989,N_12295,N_13757);
xor U17990 (N_17990,N_13235,N_14547);
nand U17991 (N_17991,N_15531,N_14485);
or U17992 (N_17992,N_12364,N_14500);
nand U17993 (N_17993,N_12553,N_15826);
nand U17994 (N_17994,N_12358,N_12387);
or U17995 (N_17995,N_14805,N_13346);
or U17996 (N_17996,N_13384,N_12975);
or U17997 (N_17997,N_15408,N_13718);
or U17998 (N_17998,N_13344,N_13411);
and U17999 (N_17999,N_15318,N_14021);
nand U18000 (N_18000,N_15196,N_12875);
and U18001 (N_18001,N_15819,N_15524);
and U18002 (N_18002,N_15283,N_13069);
nor U18003 (N_18003,N_13553,N_13808);
or U18004 (N_18004,N_15989,N_13673);
nor U18005 (N_18005,N_14428,N_13977);
and U18006 (N_18006,N_12771,N_12742);
nand U18007 (N_18007,N_13770,N_12885);
xor U18008 (N_18008,N_13657,N_14475);
xnor U18009 (N_18009,N_14779,N_14032);
and U18010 (N_18010,N_15986,N_13501);
and U18011 (N_18011,N_12115,N_14972);
nand U18012 (N_18012,N_15082,N_14383);
or U18013 (N_18013,N_14929,N_12368);
xnor U18014 (N_18014,N_15298,N_13946);
xnor U18015 (N_18015,N_13704,N_14757);
xnor U18016 (N_18016,N_13202,N_13794);
or U18017 (N_18017,N_13971,N_14981);
or U18018 (N_18018,N_13601,N_12552);
nor U18019 (N_18019,N_13818,N_14831);
xor U18020 (N_18020,N_12646,N_15605);
and U18021 (N_18021,N_15657,N_12884);
and U18022 (N_18022,N_14512,N_13012);
nor U18023 (N_18023,N_14410,N_14993);
or U18024 (N_18024,N_12521,N_12253);
nor U18025 (N_18025,N_13607,N_12735);
and U18026 (N_18026,N_14049,N_15735);
and U18027 (N_18027,N_15981,N_15621);
or U18028 (N_18028,N_13576,N_12699);
and U18029 (N_18029,N_13727,N_15361);
or U18030 (N_18030,N_14557,N_14339);
nor U18031 (N_18031,N_15463,N_14015);
nor U18032 (N_18032,N_14384,N_15140);
nand U18033 (N_18033,N_13342,N_14641);
and U18034 (N_18034,N_15711,N_12981);
nor U18035 (N_18035,N_13555,N_14325);
xor U18036 (N_18036,N_15559,N_12255);
nand U18037 (N_18037,N_12531,N_15375);
nor U18038 (N_18038,N_13444,N_13736);
nor U18039 (N_18039,N_13013,N_13858);
xor U18040 (N_18040,N_15912,N_13284);
nor U18041 (N_18041,N_13471,N_15223);
or U18042 (N_18042,N_14371,N_12677);
nor U18043 (N_18043,N_14697,N_12677);
nand U18044 (N_18044,N_13506,N_15144);
nand U18045 (N_18045,N_15479,N_15227);
nand U18046 (N_18046,N_14074,N_13551);
nand U18047 (N_18047,N_13311,N_12109);
xnor U18048 (N_18048,N_14749,N_12410);
xor U18049 (N_18049,N_14354,N_13966);
or U18050 (N_18050,N_12829,N_14005);
xnor U18051 (N_18051,N_12996,N_14488);
xor U18052 (N_18052,N_12871,N_15324);
or U18053 (N_18053,N_15864,N_12919);
xnor U18054 (N_18054,N_15732,N_13027);
and U18055 (N_18055,N_12766,N_14980);
or U18056 (N_18056,N_12623,N_12910);
nor U18057 (N_18057,N_13741,N_13228);
xor U18058 (N_18058,N_14514,N_14765);
or U18059 (N_18059,N_13089,N_15207);
nand U18060 (N_18060,N_15837,N_14608);
nor U18061 (N_18061,N_13119,N_13468);
xnor U18062 (N_18062,N_12979,N_13259);
or U18063 (N_18063,N_12558,N_14087);
or U18064 (N_18064,N_12756,N_12238);
and U18065 (N_18065,N_13466,N_12834);
or U18066 (N_18066,N_14323,N_14280);
nor U18067 (N_18067,N_15259,N_14406);
xor U18068 (N_18068,N_13848,N_12659);
nor U18069 (N_18069,N_13612,N_14035);
nand U18070 (N_18070,N_13678,N_14759);
xor U18071 (N_18071,N_12494,N_13210);
xnor U18072 (N_18072,N_12980,N_15001);
xnor U18073 (N_18073,N_12539,N_15535);
and U18074 (N_18074,N_14432,N_13824);
nor U18075 (N_18075,N_13865,N_13986);
xor U18076 (N_18076,N_12437,N_15067);
xor U18077 (N_18077,N_15688,N_13178);
nand U18078 (N_18078,N_12183,N_15687);
or U18079 (N_18079,N_14417,N_14756);
nand U18080 (N_18080,N_12070,N_14182);
and U18081 (N_18081,N_13092,N_12847);
nand U18082 (N_18082,N_13197,N_15425);
or U18083 (N_18083,N_14813,N_14153);
xor U18084 (N_18084,N_12559,N_15903);
and U18085 (N_18085,N_13049,N_12573);
or U18086 (N_18086,N_15654,N_12435);
xnor U18087 (N_18087,N_15499,N_12422);
nand U18088 (N_18088,N_13027,N_13647);
and U18089 (N_18089,N_13451,N_12406);
nor U18090 (N_18090,N_14912,N_13694);
or U18091 (N_18091,N_15583,N_15508);
xnor U18092 (N_18092,N_12850,N_13135);
and U18093 (N_18093,N_12456,N_12272);
nand U18094 (N_18094,N_13292,N_13035);
nand U18095 (N_18095,N_13694,N_15262);
nand U18096 (N_18096,N_13672,N_14351);
nand U18097 (N_18097,N_13969,N_15537);
nand U18098 (N_18098,N_12062,N_13022);
xor U18099 (N_18099,N_12327,N_13904);
and U18100 (N_18100,N_12101,N_14628);
and U18101 (N_18101,N_12734,N_13951);
or U18102 (N_18102,N_14595,N_15502);
xor U18103 (N_18103,N_13291,N_13116);
or U18104 (N_18104,N_15022,N_15450);
or U18105 (N_18105,N_13809,N_15041);
nand U18106 (N_18106,N_14949,N_14817);
and U18107 (N_18107,N_13882,N_15783);
nand U18108 (N_18108,N_13972,N_13536);
and U18109 (N_18109,N_12334,N_15154);
nor U18110 (N_18110,N_15999,N_13972);
and U18111 (N_18111,N_13696,N_12757);
xnor U18112 (N_18112,N_13842,N_14898);
and U18113 (N_18113,N_14296,N_15346);
or U18114 (N_18114,N_13957,N_13400);
or U18115 (N_18115,N_15966,N_12615);
nor U18116 (N_18116,N_15946,N_12667);
or U18117 (N_18117,N_12722,N_14480);
nand U18118 (N_18118,N_15242,N_14080);
xor U18119 (N_18119,N_15696,N_13689);
nand U18120 (N_18120,N_12519,N_15887);
nand U18121 (N_18121,N_12664,N_15304);
xor U18122 (N_18122,N_15130,N_13115);
nand U18123 (N_18123,N_15947,N_15899);
xor U18124 (N_18124,N_12292,N_12225);
xor U18125 (N_18125,N_14854,N_15905);
nand U18126 (N_18126,N_15332,N_12393);
nand U18127 (N_18127,N_13524,N_14277);
nor U18128 (N_18128,N_13627,N_14283);
nand U18129 (N_18129,N_14358,N_15504);
and U18130 (N_18130,N_12301,N_14928);
nand U18131 (N_18131,N_15144,N_12273);
xnor U18132 (N_18132,N_15231,N_15836);
or U18133 (N_18133,N_12806,N_15752);
or U18134 (N_18134,N_13988,N_12481);
nor U18135 (N_18135,N_15850,N_12529);
nand U18136 (N_18136,N_13022,N_12126);
xor U18137 (N_18137,N_12342,N_12848);
nor U18138 (N_18138,N_14553,N_14658);
and U18139 (N_18139,N_14114,N_15197);
xor U18140 (N_18140,N_14429,N_14170);
nor U18141 (N_18141,N_13045,N_15029);
or U18142 (N_18142,N_12997,N_14279);
xor U18143 (N_18143,N_13954,N_15763);
nand U18144 (N_18144,N_14869,N_13553);
nor U18145 (N_18145,N_14974,N_14744);
and U18146 (N_18146,N_13628,N_13771);
and U18147 (N_18147,N_15031,N_14814);
xor U18148 (N_18148,N_12666,N_14151);
xnor U18149 (N_18149,N_15077,N_14323);
or U18150 (N_18150,N_12786,N_12848);
nor U18151 (N_18151,N_12996,N_15437);
nor U18152 (N_18152,N_13474,N_13140);
nand U18153 (N_18153,N_12067,N_14280);
nor U18154 (N_18154,N_14656,N_15378);
or U18155 (N_18155,N_13688,N_14203);
nor U18156 (N_18156,N_12761,N_15842);
xor U18157 (N_18157,N_14277,N_14647);
or U18158 (N_18158,N_15298,N_14999);
xor U18159 (N_18159,N_13740,N_14052);
and U18160 (N_18160,N_12583,N_14296);
or U18161 (N_18161,N_14843,N_12707);
xnor U18162 (N_18162,N_15785,N_12361);
xnor U18163 (N_18163,N_14786,N_12286);
nor U18164 (N_18164,N_14537,N_15098);
or U18165 (N_18165,N_13505,N_13929);
or U18166 (N_18166,N_12182,N_12157);
nand U18167 (N_18167,N_12856,N_15684);
or U18168 (N_18168,N_12140,N_13067);
xor U18169 (N_18169,N_13903,N_15612);
nor U18170 (N_18170,N_14049,N_14671);
nor U18171 (N_18171,N_14226,N_14695);
nor U18172 (N_18172,N_12419,N_15321);
or U18173 (N_18173,N_13553,N_12232);
xor U18174 (N_18174,N_14606,N_13098);
nor U18175 (N_18175,N_13977,N_13078);
and U18176 (N_18176,N_15191,N_14533);
or U18177 (N_18177,N_15839,N_12177);
nor U18178 (N_18178,N_13497,N_14717);
or U18179 (N_18179,N_15896,N_15345);
nor U18180 (N_18180,N_15055,N_13296);
and U18181 (N_18181,N_13500,N_14000);
and U18182 (N_18182,N_15639,N_12706);
and U18183 (N_18183,N_15820,N_12199);
and U18184 (N_18184,N_14362,N_14036);
nor U18185 (N_18185,N_12996,N_14396);
or U18186 (N_18186,N_12692,N_12376);
xor U18187 (N_18187,N_15970,N_14948);
and U18188 (N_18188,N_14638,N_13798);
or U18189 (N_18189,N_12337,N_15635);
nor U18190 (N_18190,N_14732,N_14359);
nor U18191 (N_18191,N_14966,N_15778);
and U18192 (N_18192,N_15057,N_15609);
nor U18193 (N_18193,N_15550,N_13084);
xor U18194 (N_18194,N_14084,N_12801);
or U18195 (N_18195,N_13072,N_12646);
and U18196 (N_18196,N_13381,N_15034);
or U18197 (N_18197,N_13994,N_13614);
xnor U18198 (N_18198,N_15054,N_13174);
nand U18199 (N_18199,N_12462,N_14465);
nand U18200 (N_18200,N_12510,N_14992);
xor U18201 (N_18201,N_15581,N_12941);
and U18202 (N_18202,N_15969,N_12668);
nor U18203 (N_18203,N_13043,N_15577);
and U18204 (N_18204,N_15053,N_14814);
nor U18205 (N_18205,N_12772,N_12425);
or U18206 (N_18206,N_12887,N_15629);
nand U18207 (N_18207,N_15325,N_15004);
nand U18208 (N_18208,N_12828,N_12776);
nor U18209 (N_18209,N_14035,N_13424);
or U18210 (N_18210,N_14357,N_15157);
nor U18211 (N_18211,N_12442,N_15757);
and U18212 (N_18212,N_13199,N_15362);
nand U18213 (N_18213,N_13403,N_14572);
or U18214 (N_18214,N_12811,N_13669);
xnor U18215 (N_18215,N_14807,N_12940);
or U18216 (N_18216,N_13143,N_12374);
xnor U18217 (N_18217,N_12418,N_14053);
nand U18218 (N_18218,N_12757,N_12500);
xor U18219 (N_18219,N_12932,N_15303);
or U18220 (N_18220,N_14833,N_15729);
nand U18221 (N_18221,N_12358,N_13022);
nand U18222 (N_18222,N_14020,N_14882);
nor U18223 (N_18223,N_14924,N_14446);
nand U18224 (N_18224,N_13717,N_13337);
and U18225 (N_18225,N_14308,N_14495);
xor U18226 (N_18226,N_15551,N_14902);
and U18227 (N_18227,N_14792,N_15608);
nand U18228 (N_18228,N_12902,N_12277);
and U18229 (N_18229,N_14188,N_13771);
or U18230 (N_18230,N_13655,N_14538);
nor U18231 (N_18231,N_13955,N_14680);
nor U18232 (N_18232,N_13436,N_13129);
nand U18233 (N_18233,N_15981,N_15852);
and U18234 (N_18234,N_12679,N_14791);
or U18235 (N_18235,N_13731,N_14615);
xnor U18236 (N_18236,N_15307,N_15380);
and U18237 (N_18237,N_15271,N_12767);
nand U18238 (N_18238,N_14456,N_13211);
nor U18239 (N_18239,N_13208,N_15278);
xnor U18240 (N_18240,N_13118,N_12298);
nor U18241 (N_18241,N_13354,N_15104);
nand U18242 (N_18242,N_15360,N_13586);
and U18243 (N_18243,N_12128,N_15158);
or U18244 (N_18244,N_15978,N_12052);
and U18245 (N_18245,N_15316,N_12862);
nor U18246 (N_18246,N_12075,N_15493);
or U18247 (N_18247,N_15593,N_12331);
or U18248 (N_18248,N_14279,N_13254);
nand U18249 (N_18249,N_14511,N_12671);
or U18250 (N_18250,N_15749,N_13086);
nand U18251 (N_18251,N_13321,N_14436);
nor U18252 (N_18252,N_12881,N_13280);
or U18253 (N_18253,N_14637,N_13292);
and U18254 (N_18254,N_13911,N_12331);
and U18255 (N_18255,N_12616,N_14983);
or U18256 (N_18256,N_12270,N_13613);
nor U18257 (N_18257,N_13782,N_12270);
xor U18258 (N_18258,N_14793,N_15926);
nand U18259 (N_18259,N_12807,N_12754);
nor U18260 (N_18260,N_13163,N_13907);
and U18261 (N_18261,N_14359,N_15120);
or U18262 (N_18262,N_14336,N_12046);
nand U18263 (N_18263,N_14411,N_12178);
nor U18264 (N_18264,N_14766,N_12676);
xor U18265 (N_18265,N_15079,N_14765);
or U18266 (N_18266,N_13568,N_15844);
xnor U18267 (N_18267,N_12070,N_14495);
or U18268 (N_18268,N_12672,N_13330);
nor U18269 (N_18269,N_13925,N_15568);
or U18270 (N_18270,N_13885,N_12090);
nor U18271 (N_18271,N_13476,N_13979);
or U18272 (N_18272,N_14500,N_12911);
or U18273 (N_18273,N_13046,N_15629);
and U18274 (N_18274,N_15476,N_15575);
and U18275 (N_18275,N_14026,N_13761);
nor U18276 (N_18276,N_14570,N_15160);
nor U18277 (N_18277,N_12321,N_13221);
xnor U18278 (N_18278,N_13229,N_13531);
or U18279 (N_18279,N_12179,N_12526);
or U18280 (N_18280,N_12556,N_15601);
xor U18281 (N_18281,N_14282,N_12863);
xor U18282 (N_18282,N_12345,N_15579);
or U18283 (N_18283,N_12342,N_15801);
and U18284 (N_18284,N_13405,N_13389);
or U18285 (N_18285,N_12380,N_12575);
or U18286 (N_18286,N_15519,N_14356);
nor U18287 (N_18287,N_14135,N_14560);
or U18288 (N_18288,N_14690,N_13675);
nand U18289 (N_18289,N_13551,N_15221);
and U18290 (N_18290,N_14902,N_15754);
nand U18291 (N_18291,N_13827,N_14472);
and U18292 (N_18292,N_12905,N_15849);
nand U18293 (N_18293,N_12525,N_14440);
nor U18294 (N_18294,N_15441,N_15551);
nor U18295 (N_18295,N_13729,N_12275);
and U18296 (N_18296,N_12277,N_13846);
nor U18297 (N_18297,N_15013,N_15809);
xor U18298 (N_18298,N_13088,N_12690);
xor U18299 (N_18299,N_15834,N_12820);
and U18300 (N_18300,N_12115,N_12055);
or U18301 (N_18301,N_14659,N_15463);
or U18302 (N_18302,N_15459,N_14296);
xnor U18303 (N_18303,N_14953,N_13303);
and U18304 (N_18304,N_15077,N_15978);
or U18305 (N_18305,N_13202,N_13102);
or U18306 (N_18306,N_15046,N_15388);
or U18307 (N_18307,N_15596,N_13718);
or U18308 (N_18308,N_15125,N_14813);
and U18309 (N_18309,N_15113,N_12807);
or U18310 (N_18310,N_14214,N_14513);
and U18311 (N_18311,N_15413,N_12199);
xor U18312 (N_18312,N_15950,N_12612);
nand U18313 (N_18313,N_14845,N_13268);
xnor U18314 (N_18314,N_14527,N_12527);
or U18315 (N_18315,N_15067,N_13063);
nor U18316 (N_18316,N_15984,N_15670);
or U18317 (N_18317,N_13312,N_13531);
nand U18318 (N_18318,N_12015,N_15359);
nand U18319 (N_18319,N_13192,N_13318);
nand U18320 (N_18320,N_12502,N_14337);
and U18321 (N_18321,N_12191,N_14778);
and U18322 (N_18322,N_12307,N_14882);
xnor U18323 (N_18323,N_15200,N_14122);
xnor U18324 (N_18324,N_13746,N_13575);
and U18325 (N_18325,N_12974,N_12657);
xor U18326 (N_18326,N_15323,N_12972);
or U18327 (N_18327,N_14486,N_14439);
and U18328 (N_18328,N_13611,N_15476);
nand U18329 (N_18329,N_12737,N_14611);
xor U18330 (N_18330,N_12715,N_15698);
nand U18331 (N_18331,N_15631,N_12525);
or U18332 (N_18332,N_14507,N_13533);
xnor U18333 (N_18333,N_14880,N_14570);
nand U18334 (N_18334,N_13459,N_14332);
or U18335 (N_18335,N_14612,N_14805);
xnor U18336 (N_18336,N_14512,N_14447);
or U18337 (N_18337,N_12269,N_13227);
nor U18338 (N_18338,N_14913,N_15162);
nand U18339 (N_18339,N_15566,N_15569);
nor U18340 (N_18340,N_12684,N_12366);
xor U18341 (N_18341,N_14794,N_14877);
or U18342 (N_18342,N_14289,N_13692);
and U18343 (N_18343,N_14736,N_12003);
or U18344 (N_18344,N_13305,N_13427);
nor U18345 (N_18345,N_12531,N_14522);
xnor U18346 (N_18346,N_14663,N_13919);
or U18347 (N_18347,N_14899,N_13976);
nor U18348 (N_18348,N_14502,N_15218);
and U18349 (N_18349,N_12464,N_12873);
and U18350 (N_18350,N_12248,N_13298);
nor U18351 (N_18351,N_13729,N_15350);
and U18352 (N_18352,N_13889,N_14516);
nand U18353 (N_18353,N_12247,N_13680);
and U18354 (N_18354,N_12485,N_13375);
nor U18355 (N_18355,N_12132,N_14089);
and U18356 (N_18356,N_14309,N_15129);
xnor U18357 (N_18357,N_14924,N_14744);
xnor U18358 (N_18358,N_13433,N_12732);
or U18359 (N_18359,N_13223,N_13638);
and U18360 (N_18360,N_12099,N_13279);
xor U18361 (N_18361,N_15637,N_15085);
xor U18362 (N_18362,N_14811,N_13946);
nor U18363 (N_18363,N_13870,N_15392);
or U18364 (N_18364,N_12211,N_15115);
nand U18365 (N_18365,N_14386,N_15878);
xor U18366 (N_18366,N_13731,N_15491);
xor U18367 (N_18367,N_12378,N_13965);
nor U18368 (N_18368,N_12763,N_12846);
xor U18369 (N_18369,N_12546,N_15643);
and U18370 (N_18370,N_15633,N_13684);
xor U18371 (N_18371,N_14949,N_12840);
nor U18372 (N_18372,N_12197,N_15484);
xor U18373 (N_18373,N_12235,N_14016);
xor U18374 (N_18374,N_14468,N_15521);
xnor U18375 (N_18375,N_15795,N_12316);
and U18376 (N_18376,N_15922,N_15820);
xnor U18377 (N_18377,N_12488,N_12429);
xor U18378 (N_18378,N_12375,N_13413);
or U18379 (N_18379,N_13850,N_12768);
nor U18380 (N_18380,N_13968,N_15687);
nand U18381 (N_18381,N_13879,N_14233);
nand U18382 (N_18382,N_12793,N_14593);
xor U18383 (N_18383,N_14979,N_12099);
nor U18384 (N_18384,N_14695,N_14405);
nand U18385 (N_18385,N_15736,N_12875);
or U18386 (N_18386,N_13389,N_12756);
and U18387 (N_18387,N_14442,N_14362);
xnor U18388 (N_18388,N_15788,N_15756);
nand U18389 (N_18389,N_13726,N_13931);
xor U18390 (N_18390,N_14138,N_14400);
nand U18391 (N_18391,N_14779,N_15820);
nand U18392 (N_18392,N_12451,N_15974);
xnor U18393 (N_18393,N_12608,N_13423);
or U18394 (N_18394,N_13553,N_13162);
and U18395 (N_18395,N_15356,N_13179);
and U18396 (N_18396,N_12033,N_12052);
and U18397 (N_18397,N_15218,N_13030);
and U18398 (N_18398,N_14040,N_14802);
nand U18399 (N_18399,N_12275,N_12492);
and U18400 (N_18400,N_13114,N_15128);
xor U18401 (N_18401,N_15545,N_13277);
nor U18402 (N_18402,N_15845,N_12110);
nor U18403 (N_18403,N_14963,N_13610);
or U18404 (N_18404,N_12328,N_13821);
or U18405 (N_18405,N_14675,N_14624);
xnor U18406 (N_18406,N_13202,N_15184);
xnor U18407 (N_18407,N_13934,N_15440);
nand U18408 (N_18408,N_12467,N_14853);
xnor U18409 (N_18409,N_15967,N_15105);
nand U18410 (N_18410,N_13116,N_14644);
xnor U18411 (N_18411,N_13041,N_12420);
nor U18412 (N_18412,N_12057,N_14219);
or U18413 (N_18413,N_13071,N_12656);
and U18414 (N_18414,N_13607,N_13940);
xnor U18415 (N_18415,N_13166,N_15993);
or U18416 (N_18416,N_14785,N_14184);
and U18417 (N_18417,N_13381,N_12510);
nand U18418 (N_18418,N_15615,N_15246);
or U18419 (N_18419,N_14184,N_14424);
nand U18420 (N_18420,N_14191,N_15939);
nand U18421 (N_18421,N_14424,N_12549);
or U18422 (N_18422,N_13104,N_15404);
or U18423 (N_18423,N_13908,N_14036);
nor U18424 (N_18424,N_14116,N_13672);
nand U18425 (N_18425,N_12017,N_14942);
nor U18426 (N_18426,N_14395,N_15624);
or U18427 (N_18427,N_15853,N_15288);
xor U18428 (N_18428,N_13554,N_14182);
nand U18429 (N_18429,N_13974,N_12787);
or U18430 (N_18430,N_15915,N_15038);
nand U18431 (N_18431,N_14260,N_14041);
nand U18432 (N_18432,N_15300,N_14544);
and U18433 (N_18433,N_14452,N_14390);
nor U18434 (N_18434,N_13514,N_15943);
or U18435 (N_18435,N_14999,N_15759);
and U18436 (N_18436,N_13902,N_12915);
or U18437 (N_18437,N_14668,N_15367);
or U18438 (N_18438,N_13192,N_15364);
nand U18439 (N_18439,N_14625,N_13135);
or U18440 (N_18440,N_12479,N_14247);
xnor U18441 (N_18441,N_14120,N_14461);
nand U18442 (N_18442,N_12504,N_14121);
or U18443 (N_18443,N_14676,N_12423);
or U18444 (N_18444,N_14662,N_12940);
nor U18445 (N_18445,N_12210,N_13698);
and U18446 (N_18446,N_12555,N_15911);
nor U18447 (N_18447,N_14210,N_14351);
nor U18448 (N_18448,N_14253,N_14276);
and U18449 (N_18449,N_13001,N_15960);
nand U18450 (N_18450,N_15349,N_15820);
and U18451 (N_18451,N_14414,N_13096);
nor U18452 (N_18452,N_13449,N_14572);
or U18453 (N_18453,N_14923,N_14232);
or U18454 (N_18454,N_13478,N_12247);
xor U18455 (N_18455,N_14454,N_12117);
xnor U18456 (N_18456,N_13257,N_14562);
and U18457 (N_18457,N_14968,N_13440);
or U18458 (N_18458,N_14546,N_13945);
nor U18459 (N_18459,N_14649,N_12227);
xnor U18460 (N_18460,N_12144,N_15503);
xnor U18461 (N_18461,N_15934,N_13473);
nand U18462 (N_18462,N_15667,N_15503);
nand U18463 (N_18463,N_14318,N_14470);
nand U18464 (N_18464,N_12738,N_15119);
xor U18465 (N_18465,N_15426,N_13132);
and U18466 (N_18466,N_15424,N_12622);
nor U18467 (N_18467,N_15334,N_15437);
or U18468 (N_18468,N_12111,N_12014);
and U18469 (N_18469,N_12493,N_12180);
or U18470 (N_18470,N_12545,N_15545);
or U18471 (N_18471,N_15856,N_15123);
nand U18472 (N_18472,N_13063,N_12048);
nand U18473 (N_18473,N_13109,N_13106);
xnor U18474 (N_18474,N_14598,N_13441);
xor U18475 (N_18475,N_15778,N_12724);
or U18476 (N_18476,N_14323,N_13369);
nand U18477 (N_18477,N_14650,N_13088);
and U18478 (N_18478,N_13501,N_14008);
and U18479 (N_18479,N_15987,N_15091);
nand U18480 (N_18480,N_15922,N_12250);
or U18481 (N_18481,N_13163,N_14191);
xor U18482 (N_18482,N_13288,N_14656);
or U18483 (N_18483,N_12762,N_12180);
or U18484 (N_18484,N_14853,N_14500);
or U18485 (N_18485,N_15967,N_12373);
xor U18486 (N_18486,N_14011,N_14854);
nand U18487 (N_18487,N_12260,N_14825);
or U18488 (N_18488,N_13101,N_12933);
nor U18489 (N_18489,N_15072,N_14265);
nor U18490 (N_18490,N_12945,N_15289);
nor U18491 (N_18491,N_13325,N_13857);
nand U18492 (N_18492,N_15273,N_14098);
or U18493 (N_18493,N_14491,N_12347);
or U18494 (N_18494,N_13686,N_15955);
or U18495 (N_18495,N_15164,N_13331);
nor U18496 (N_18496,N_13429,N_14457);
nand U18497 (N_18497,N_14534,N_14698);
or U18498 (N_18498,N_14610,N_12408);
nor U18499 (N_18499,N_15265,N_12501);
nor U18500 (N_18500,N_14973,N_14211);
nand U18501 (N_18501,N_13251,N_14596);
and U18502 (N_18502,N_14651,N_12679);
or U18503 (N_18503,N_12924,N_12945);
or U18504 (N_18504,N_14874,N_14201);
or U18505 (N_18505,N_13192,N_15759);
nor U18506 (N_18506,N_13559,N_15416);
nand U18507 (N_18507,N_14989,N_13248);
or U18508 (N_18508,N_15778,N_14969);
or U18509 (N_18509,N_14188,N_14530);
xor U18510 (N_18510,N_14293,N_12189);
and U18511 (N_18511,N_14863,N_12987);
xnor U18512 (N_18512,N_14907,N_15443);
xnor U18513 (N_18513,N_14911,N_13976);
and U18514 (N_18514,N_13083,N_14149);
nand U18515 (N_18515,N_12250,N_14493);
or U18516 (N_18516,N_12480,N_15403);
nand U18517 (N_18517,N_13744,N_12927);
and U18518 (N_18518,N_12054,N_13716);
or U18519 (N_18519,N_14301,N_13730);
nand U18520 (N_18520,N_13802,N_15631);
nor U18521 (N_18521,N_13572,N_13345);
and U18522 (N_18522,N_12324,N_14309);
nor U18523 (N_18523,N_13109,N_13304);
nor U18524 (N_18524,N_15645,N_14658);
nand U18525 (N_18525,N_13288,N_14080);
and U18526 (N_18526,N_12061,N_14513);
or U18527 (N_18527,N_15913,N_12973);
nor U18528 (N_18528,N_12365,N_14668);
and U18529 (N_18529,N_12988,N_12845);
xnor U18530 (N_18530,N_13606,N_12977);
nand U18531 (N_18531,N_13463,N_14396);
and U18532 (N_18532,N_14465,N_14484);
and U18533 (N_18533,N_14169,N_15030);
nor U18534 (N_18534,N_14242,N_14976);
nand U18535 (N_18535,N_14669,N_14470);
and U18536 (N_18536,N_14997,N_13044);
or U18537 (N_18537,N_15988,N_12103);
xnor U18538 (N_18538,N_12251,N_12807);
nand U18539 (N_18539,N_14738,N_14710);
nor U18540 (N_18540,N_15807,N_14632);
nor U18541 (N_18541,N_15915,N_12005);
xnor U18542 (N_18542,N_15379,N_15015);
and U18543 (N_18543,N_13752,N_12389);
or U18544 (N_18544,N_14619,N_14496);
or U18545 (N_18545,N_13627,N_15705);
and U18546 (N_18546,N_13154,N_14523);
xnor U18547 (N_18547,N_15028,N_14584);
nand U18548 (N_18548,N_14040,N_13747);
or U18549 (N_18549,N_14444,N_15548);
and U18550 (N_18550,N_15844,N_14695);
xnor U18551 (N_18551,N_13720,N_13255);
and U18552 (N_18552,N_14776,N_12807);
xor U18553 (N_18553,N_14257,N_12023);
nor U18554 (N_18554,N_14658,N_13199);
nand U18555 (N_18555,N_12317,N_12765);
nor U18556 (N_18556,N_14962,N_13776);
xnor U18557 (N_18557,N_13511,N_13470);
xnor U18558 (N_18558,N_12967,N_15087);
nand U18559 (N_18559,N_13882,N_14557);
nor U18560 (N_18560,N_14245,N_13001);
and U18561 (N_18561,N_14955,N_13012);
nor U18562 (N_18562,N_13472,N_12641);
and U18563 (N_18563,N_12533,N_15665);
or U18564 (N_18564,N_14425,N_13722);
nand U18565 (N_18565,N_13002,N_13201);
xnor U18566 (N_18566,N_15976,N_15257);
nor U18567 (N_18567,N_13191,N_12172);
nand U18568 (N_18568,N_15933,N_12812);
nand U18569 (N_18569,N_15462,N_14234);
and U18570 (N_18570,N_13120,N_12575);
xnor U18571 (N_18571,N_13272,N_12717);
or U18572 (N_18572,N_13229,N_15893);
nand U18573 (N_18573,N_12074,N_12385);
xnor U18574 (N_18574,N_14189,N_15248);
nand U18575 (N_18575,N_14305,N_15272);
xnor U18576 (N_18576,N_15599,N_14098);
or U18577 (N_18577,N_13095,N_15594);
xnor U18578 (N_18578,N_15349,N_13181);
nand U18579 (N_18579,N_13891,N_13049);
nor U18580 (N_18580,N_13822,N_12307);
and U18581 (N_18581,N_14635,N_15625);
nand U18582 (N_18582,N_14051,N_12169);
or U18583 (N_18583,N_14687,N_13597);
and U18584 (N_18584,N_13072,N_13728);
nor U18585 (N_18585,N_14292,N_12229);
xor U18586 (N_18586,N_13527,N_15964);
nor U18587 (N_18587,N_15343,N_12131);
xor U18588 (N_18588,N_14788,N_15487);
nand U18589 (N_18589,N_15178,N_13401);
nor U18590 (N_18590,N_15144,N_13229);
xnor U18591 (N_18591,N_13581,N_13766);
or U18592 (N_18592,N_15891,N_12964);
and U18593 (N_18593,N_12809,N_12685);
or U18594 (N_18594,N_14403,N_13981);
nor U18595 (N_18595,N_15596,N_15050);
nand U18596 (N_18596,N_13906,N_12718);
and U18597 (N_18597,N_12926,N_13368);
or U18598 (N_18598,N_12915,N_12305);
xnor U18599 (N_18599,N_14398,N_15235);
xor U18600 (N_18600,N_13703,N_15067);
nand U18601 (N_18601,N_12082,N_13859);
nor U18602 (N_18602,N_14137,N_15223);
nand U18603 (N_18603,N_14922,N_14297);
or U18604 (N_18604,N_13951,N_15631);
xnor U18605 (N_18605,N_15378,N_14402);
nand U18606 (N_18606,N_15660,N_14310);
or U18607 (N_18607,N_13286,N_13548);
xnor U18608 (N_18608,N_13667,N_13112);
xnor U18609 (N_18609,N_15469,N_13144);
and U18610 (N_18610,N_13962,N_14253);
or U18611 (N_18611,N_15560,N_13023);
nand U18612 (N_18612,N_13204,N_12303);
nor U18613 (N_18613,N_14021,N_12941);
nand U18614 (N_18614,N_12942,N_15956);
nand U18615 (N_18615,N_15078,N_14545);
or U18616 (N_18616,N_12806,N_13085);
and U18617 (N_18617,N_14030,N_12075);
or U18618 (N_18618,N_15761,N_13571);
nand U18619 (N_18619,N_14862,N_13367);
nor U18620 (N_18620,N_13671,N_14018);
xor U18621 (N_18621,N_12272,N_15588);
or U18622 (N_18622,N_13893,N_14697);
or U18623 (N_18623,N_15405,N_15104);
nor U18624 (N_18624,N_13480,N_13196);
xor U18625 (N_18625,N_15987,N_13802);
xor U18626 (N_18626,N_15567,N_14328);
or U18627 (N_18627,N_12515,N_14452);
and U18628 (N_18628,N_15259,N_15832);
nand U18629 (N_18629,N_12969,N_13272);
or U18630 (N_18630,N_13849,N_15732);
or U18631 (N_18631,N_15046,N_13576);
nor U18632 (N_18632,N_14905,N_12963);
or U18633 (N_18633,N_15713,N_12918);
and U18634 (N_18634,N_12110,N_14950);
or U18635 (N_18635,N_14684,N_14652);
xor U18636 (N_18636,N_13496,N_12391);
nand U18637 (N_18637,N_13406,N_14995);
xor U18638 (N_18638,N_15493,N_14768);
xnor U18639 (N_18639,N_15423,N_12118);
nor U18640 (N_18640,N_13259,N_14298);
and U18641 (N_18641,N_13575,N_12339);
or U18642 (N_18642,N_13553,N_14720);
xnor U18643 (N_18643,N_15737,N_15849);
nor U18644 (N_18644,N_13592,N_15258);
or U18645 (N_18645,N_12362,N_15459);
and U18646 (N_18646,N_12794,N_14800);
and U18647 (N_18647,N_14019,N_13580);
or U18648 (N_18648,N_15163,N_12815);
and U18649 (N_18649,N_15461,N_15392);
xor U18650 (N_18650,N_12569,N_12610);
xnor U18651 (N_18651,N_15005,N_12724);
nand U18652 (N_18652,N_12576,N_13979);
or U18653 (N_18653,N_12030,N_13706);
and U18654 (N_18654,N_15664,N_13709);
and U18655 (N_18655,N_15756,N_14081);
or U18656 (N_18656,N_12076,N_13885);
nand U18657 (N_18657,N_12234,N_13230);
nor U18658 (N_18658,N_14874,N_13856);
xnor U18659 (N_18659,N_13708,N_12315);
and U18660 (N_18660,N_13974,N_14274);
nand U18661 (N_18661,N_15786,N_14127);
nor U18662 (N_18662,N_14557,N_15541);
nand U18663 (N_18663,N_13575,N_12864);
nor U18664 (N_18664,N_12584,N_14539);
nor U18665 (N_18665,N_14495,N_13207);
xnor U18666 (N_18666,N_15552,N_15624);
or U18667 (N_18667,N_13517,N_12391);
nand U18668 (N_18668,N_14399,N_13508);
and U18669 (N_18669,N_15241,N_13371);
or U18670 (N_18670,N_12215,N_13709);
xnor U18671 (N_18671,N_13274,N_13930);
nand U18672 (N_18672,N_14726,N_15209);
xor U18673 (N_18673,N_15144,N_14810);
or U18674 (N_18674,N_14952,N_14847);
nand U18675 (N_18675,N_14260,N_15459);
or U18676 (N_18676,N_14796,N_15243);
nor U18677 (N_18677,N_13270,N_14881);
nand U18678 (N_18678,N_14765,N_15661);
nand U18679 (N_18679,N_14035,N_15401);
xor U18680 (N_18680,N_15126,N_15776);
xor U18681 (N_18681,N_13550,N_13462);
or U18682 (N_18682,N_13144,N_13532);
xnor U18683 (N_18683,N_13188,N_13146);
xnor U18684 (N_18684,N_15912,N_12519);
or U18685 (N_18685,N_15810,N_15121);
and U18686 (N_18686,N_13471,N_15715);
nor U18687 (N_18687,N_14323,N_12982);
xor U18688 (N_18688,N_12923,N_13068);
nor U18689 (N_18689,N_14265,N_14030);
or U18690 (N_18690,N_13185,N_14951);
or U18691 (N_18691,N_14025,N_15745);
nand U18692 (N_18692,N_13899,N_15856);
xnor U18693 (N_18693,N_12130,N_12708);
nand U18694 (N_18694,N_12198,N_13138);
or U18695 (N_18695,N_15240,N_14114);
or U18696 (N_18696,N_14789,N_15374);
nand U18697 (N_18697,N_12531,N_15525);
xnor U18698 (N_18698,N_13789,N_12300);
and U18699 (N_18699,N_13600,N_13017);
and U18700 (N_18700,N_15036,N_14541);
or U18701 (N_18701,N_13389,N_15265);
or U18702 (N_18702,N_13896,N_15639);
or U18703 (N_18703,N_15619,N_13359);
nand U18704 (N_18704,N_15115,N_13913);
nor U18705 (N_18705,N_14725,N_13117);
or U18706 (N_18706,N_13621,N_15887);
nor U18707 (N_18707,N_14914,N_15201);
and U18708 (N_18708,N_15554,N_15609);
nor U18709 (N_18709,N_14377,N_13139);
nand U18710 (N_18710,N_14883,N_14760);
or U18711 (N_18711,N_13152,N_13846);
nor U18712 (N_18712,N_14871,N_15398);
nand U18713 (N_18713,N_14182,N_14002);
nor U18714 (N_18714,N_15289,N_12374);
nand U18715 (N_18715,N_14101,N_15323);
xnor U18716 (N_18716,N_14047,N_14643);
nor U18717 (N_18717,N_12524,N_12886);
nor U18718 (N_18718,N_14814,N_14067);
nor U18719 (N_18719,N_14230,N_13526);
xnor U18720 (N_18720,N_12596,N_14752);
and U18721 (N_18721,N_14158,N_13350);
and U18722 (N_18722,N_12332,N_13121);
nand U18723 (N_18723,N_12309,N_15196);
nor U18724 (N_18724,N_14339,N_15310);
or U18725 (N_18725,N_15104,N_15298);
or U18726 (N_18726,N_13371,N_15678);
and U18727 (N_18727,N_13025,N_13946);
or U18728 (N_18728,N_13409,N_14391);
or U18729 (N_18729,N_14674,N_12187);
nand U18730 (N_18730,N_12083,N_13176);
and U18731 (N_18731,N_14480,N_14081);
nor U18732 (N_18732,N_14065,N_12458);
or U18733 (N_18733,N_12170,N_15074);
or U18734 (N_18734,N_13630,N_15117);
or U18735 (N_18735,N_12678,N_13353);
or U18736 (N_18736,N_15700,N_12917);
or U18737 (N_18737,N_15810,N_13942);
and U18738 (N_18738,N_15826,N_12774);
and U18739 (N_18739,N_13461,N_12625);
or U18740 (N_18740,N_13456,N_13491);
or U18741 (N_18741,N_14183,N_13106);
and U18742 (N_18742,N_14720,N_15870);
xor U18743 (N_18743,N_12069,N_15626);
or U18744 (N_18744,N_14733,N_15607);
and U18745 (N_18745,N_14287,N_14864);
nand U18746 (N_18746,N_15277,N_15256);
or U18747 (N_18747,N_15185,N_14071);
and U18748 (N_18748,N_12377,N_13106);
nor U18749 (N_18749,N_12834,N_13091);
or U18750 (N_18750,N_14992,N_12184);
nor U18751 (N_18751,N_14301,N_15198);
nor U18752 (N_18752,N_15283,N_15146);
nand U18753 (N_18753,N_14609,N_12857);
nor U18754 (N_18754,N_13037,N_13671);
nor U18755 (N_18755,N_12559,N_13121);
or U18756 (N_18756,N_13224,N_13790);
or U18757 (N_18757,N_13244,N_15479);
nor U18758 (N_18758,N_14699,N_15711);
and U18759 (N_18759,N_14507,N_12098);
xor U18760 (N_18760,N_15627,N_14115);
and U18761 (N_18761,N_15466,N_13982);
nor U18762 (N_18762,N_15510,N_13900);
xnor U18763 (N_18763,N_13706,N_12730);
nor U18764 (N_18764,N_15840,N_12405);
nor U18765 (N_18765,N_13091,N_13193);
nand U18766 (N_18766,N_14932,N_13435);
nor U18767 (N_18767,N_13956,N_15059);
xnor U18768 (N_18768,N_13165,N_13467);
or U18769 (N_18769,N_12823,N_13723);
nor U18770 (N_18770,N_14828,N_14949);
xor U18771 (N_18771,N_12011,N_14474);
or U18772 (N_18772,N_13981,N_15697);
or U18773 (N_18773,N_14351,N_14797);
xor U18774 (N_18774,N_14500,N_12153);
and U18775 (N_18775,N_14585,N_13612);
nand U18776 (N_18776,N_15823,N_12587);
nor U18777 (N_18777,N_12806,N_12449);
nand U18778 (N_18778,N_12108,N_13479);
nor U18779 (N_18779,N_14362,N_12587);
or U18780 (N_18780,N_14515,N_14618);
xnor U18781 (N_18781,N_15260,N_15014);
xor U18782 (N_18782,N_12253,N_12725);
nor U18783 (N_18783,N_14580,N_12937);
or U18784 (N_18784,N_15307,N_14467);
nand U18785 (N_18785,N_13100,N_14971);
nand U18786 (N_18786,N_14443,N_13636);
nand U18787 (N_18787,N_15567,N_15508);
nor U18788 (N_18788,N_14420,N_14853);
nand U18789 (N_18789,N_14141,N_12113);
nand U18790 (N_18790,N_14896,N_13365);
and U18791 (N_18791,N_14221,N_14650);
or U18792 (N_18792,N_14669,N_15319);
nand U18793 (N_18793,N_15838,N_15508);
xnor U18794 (N_18794,N_12688,N_12953);
xor U18795 (N_18795,N_13956,N_12643);
or U18796 (N_18796,N_14289,N_14075);
nand U18797 (N_18797,N_14725,N_12503);
nor U18798 (N_18798,N_13479,N_14992);
nand U18799 (N_18799,N_12042,N_15369);
nand U18800 (N_18800,N_14431,N_14583);
and U18801 (N_18801,N_15198,N_15248);
and U18802 (N_18802,N_12629,N_12058);
nor U18803 (N_18803,N_12334,N_12848);
nor U18804 (N_18804,N_14433,N_13831);
or U18805 (N_18805,N_13152,N_15176);
xor U18806 (N_18806,N_12470,N_13173);
xor U18807 (N_18807,N_12019,N_14523);
nor U18808 (N_18808,N_14522,N_15144);
xor U18809 (N_18809,N_14025,N_12872);
or U18810 (N_18810,N_15624,N_15921);
and U18811 (N_18811,N_12163,N_14845);
nand U18812 (N_18812,N_14310,N_13265);
or U18813 (N_18813,N_13933,N_12098);
nor U18814 (N_18814,N_13553,N_13276);
and U18815 (N_18815,N_12503,N_12571);
xor U18816 (N_18816,N_12657,N_13380);
nor U18817 (N_18817,N_13310,N_15335);
nor U18818 (N_18818,N_12437,N_14888);
xor U18819 (N_18819,N_14309,N_14792);
nand U18820 (N_18820,N_15315,N_15284);
or U18821 (N_18821,N_15913,N_12795);
xor U18822 (N_18822,N_13041,N_15471);
or U18823 (N_18823,N_14433,N_15295);
and U18824 (N_18824,N_14526,N_15016);
nand U18825 (N_18825,N_12191,N_13656);
nand U18826 (N_18826,N_15189,N_14834);
nor U18827 (N_18827,N_14552,N_14728);
nand U18828 (N_18828,N_12705,N_14340);
nand U18829 (N_18829,N_12670,N_14196);
nand U18830 (N_18830,N_13300,N_13032);
nand U18831 (N_18831,N_15773,N_12714);
nor U18832 (N_18832,N_12764,N_12402);
nand U18833 (N_18833,N_13652,N_15093);
xor U18834 (N_18834,N_14191,N_12509);
or U18835 (N_18835,N_15291,N_14379);
nand U18836 (N_18836,N_15829,N_15674);
xor U18837 (N_18837,N_15568,N_14205);
nand U18838 (N_18838,N_14231,N_15867);
nor U18839 (N_18839,N_15450,N_14194);
nor U18840 (N_18840,N_15639,N_15703);
nand U18841 (N_18841,N_14634,N_12277);
nor U18842 (N_18842,N_15046,N_15044);
xnor U18843 (N_18843,N_14231,N_13080);
xor U18844 (N_18844,N_14432,N_12333);
and U18845 (N_18845,N_15948,N_12095);
xnor U18846 (N_18846,N_14398,N_14276);
nand U18847 (N_18847,N_15796,N_13652);
nor U18848 (N_18848,N_13622,N_12922);
and U18849 (N_18849,N_12967,N_15855);
nor U18850 (N_18850,N_15841,N_12486);
xor U18851 (N_18851,N_14930,N_13063);
nor U18852 (N_18852,N_13358,N_12113);
nand U18853 (N_18853,N_13526,N_13047);
and U18854 (N_18854,N_14447,N_14846);
xnor U18855 (N_18855,N_13592,N_15927);
xnor U18856 (N_18856,N_15017,N_13365);
nand U18857 (N_18857,N_14401,N_15828);
and U18858 (N_18858,N_14753,N_12943);
xnor U18859 (N_18859,N_13992,N_14478);
and U18860 (N_18860,N_15722,N_13130);
xor U18861 (N_18861,N_12810,N_12611);
xor U18862 (N_18862,N_13743,N_13953);
xnor U18863 (N_18863,N_14507,N_14900);
nand U18864 (N_18864,N_12296,N_15821);
nand U18865 (N_18865,N_13622,N_15270);
xnor U18866 (N_18866,N_12496,N_14067);
nor U18867 (N_18867,N_15389,N_13436);
and U18868 (N_18868,N_15065,N_15392);
nand U18869 (N_18869,N_14613,N_15718);
nand U18870 (N_18870,N_14802,N_13989);
and U18871 (N_18871,N_12285,N_14883);
and U18872 (N_18872,N_15536,N_15518);
or U18873 (N_18873,N_14801,N_13461);
or U18874 (N_18874,N_12439,N_12400);
and U18875 (N_18875,N_13599,N_15455);
and U18876 (N_18876,N_13980,N_14520);
nand U18877 (N_18877,N_13633,N_14214);
or U18878 (N_18878,N_13060,N_14879);
and U18879 (N_18879,N_13295,N_15757);
nand U18880 (N_18880,N_13153,N_15871);
nand U18881 (N_18881,N_12023,N_14828);
xor U18882 (N_18882,N_13315,N_14809);
xnor U18883 (N_18883,N_12603,N_15612);
xnor U18884 (N_18884,N_15403,N_15327);
or U18885 (N_18885,N_15672,N_12703);
or U18886 (N_18886,N_15726,N_14201);
xor U18887 (N_18887,N_14614,N_13813);
nor U18888 (N_18888,N_12088,N_14339);
xnor U18889 (N_18889,N_12344,N_13390);
and U18890 (N_18890,N_13065,N_12925);
nor U18891 (N_18891,N_12218,N_14392);
nor U18892 (N_18892,N_14269,N_12452);
xor U18893 (N_18893,N_14897,N_14881);
nand U18894 (N_18894,N_14038,N_14545);
nor U18895 (N_18895,N_14274,N_15740);
xor U18896 (N_18896,N_13294,N_12167);
or U18897 (N_18897,N_14273,N_12979);
xor U18898 (N_18898,N_13372,N_13344);
and U18899 (N_18899,N_15968,N_12287);
or U18900 (N_18900,N_14177,N_15344);
nor U18901 (N_18901,N_13785,N_12344);
and U18902 (N_18902,N_12192,N_14107);
nor U18903 (N_18903,N_12954,N_15616);
xor U18904 (N_18904,N_12298,N_14191);
or U18905 (N_18905,N_14984,N_13502);
xor U18906 (N_18906,N_13645,N_13337);
nor U18907 (N_18907,N_14814,N_15969);
nor U18908 (N_18908,N_14783,N_14804);
nand U18909 (N_18909,N_13969,N_12099);
and U18910 (N_18910,N_15946,N_14855);
xnor U18911 (N_18911,N_12306,N_13528);
nor U18912 (N_18912,N_12809,N_14657);
and U18913 (N_18913,N_15546,N_13405);
or U18914 (N_18914,N_15126,N_12505);
xor U18915 (N_18915,N_14812,N_13480);
xnor U18916 (N_18916,N_14146,N_15877);
and U18917 (N_18917,N_13802,N_15104);
xor U18918 (N_18918,N_15017,N_12527);
and U18919 (N_18919,N_13427,N_13286);
nand U18920 (N_18920,N_15115,N_14427);
or U18921 (N_18921,N_14138,N_12003);
xnor U18922 (N_18922,N_15167,N_12688);
nand U18923 (N_18923,N_15381,N_14274);
or U18924 (N_18924,N_14795,N_12679);
nor U18925 (N_18925,N_14090,N_13778);
nand U18926 (N_18926,N_15678,N_13876);
xor U18927 (N_18927,N_15973,N_12927);
or U18928 (N_18928,N_15540,N_12261);
xor U18929 (N_18929,N_14123,N_15691);
nor U18930 (N_18930,N_12790,N_15477);
and U18931 (N_18931,N_14883,N_13906);
and U18932 (N_18932,N_14755,N_14389);
and U18933 (N_18933,N_15192,N_14389);
xor U18934 (N_18934,N_12993,N_13543);
and U18935 (N_18935,N_15245,N_15043);
nand U18936 (N_18936,N_14576,N_15451);
or U18937 (N_18937,N_12908,N_14020);
xor U18938 (N_18938,N_12962,N_13485);
or U18939 (N_18939,N_13777,N_13677);
nor U18940 (N_18940,N_15231,N_14382);
or U18941 (N_18941,N_15090,N_12731);
xnor U18942 (N_18942,N_12847,N_12691);
xnor U18943 (N_18943,N_15892,N_14632);
xor U18944 (N_18944,N_13848,N_15080);
or U18945 (N_18945,N_12516,N_12403);
or U18946 (N_18946,N_14471,N_12499);
xnor U18947 (N_18947,N_14208,N_13092);
or U18948 (N_18948,N_13267,N_12147);
nor U18949 (N_18949,N_15056,N_12640);
nor U18950 (N_18950,N_15562,N_12241);
nand U18951 (N_18951,N_12368,N_13648);
or U18952 (N_18952,N_12837,N_13298);
or U18953 (N_18953,N_15285,N_15890);
xnor U18954 (N_18954,N_15433,N_15673);
or U18955 (N_18955,N_12846,N_12484);
nor U18956 (N_18956,N_15129,N_12937);
and U18957 (N_18957,N_13542,N_15828);
xor U18958 (N_18958,N_15099,N_12046);
or U18959 (N_18959,N_13955,N_12064);
nor U18960 (N_18960,N_14195,N_15184);
nor U18961 (N_18961,N_12218,N_12400);
and U18962 (N_18962,N_15508,N_14913);
xnor U18963 (N_18963,N_13488,N_13617);
nor U18964 (N_18964,N_13215,N_12057);
and U18965 (N_18965,N_14645,N_14207);
or U18966 (N_18966,N_12810,N_13041);
or U18967 (N_18967,N_15275,N_12849);
xor U18968 (N_18968,N_15246,N_15039);
or U18969 (N_18969,N_14660,N_13256);
nor U18970 (N_18970,N_14885,N_12963);
and U18971 (N_18971,N_15523,N_13553);
and U18972 (N_18972,N_14278,N_13109);
or U18973 (N_18973,N_14461,N_13793);
nand U18974 (N_18974,N_13904,N_15386);
xor U18975 (N_18975,N_13933,N_12824);
and U18976 (N_18976,N_15726,N_14694);
nand U18977 (N_18977,N_15303,N_13001);
xor U18978 (N_18978,N_12393,N_12349);
or U18979 (N_18979,N_13049,N_15348);
and U18980 (N_18980,N_14667,N_14831);
nor U18981 (N_18981,N_14968,N_13859);
nor U18982 (N_18982,N_13434,N_14899);
or U18983 (N_18983,N_14784,N_14552);
xnor U18984 (N_18984,N_15874,N_15809);
or U18985 (N_18985,N_15239,N_15487);
xnor U18986 (N_18986,N_14760,N_14275);
and U18987 (N_18987,N_13741,N_14857);
or U18988 (N_18988,N_15384,N_12058);
nor U18989 (N_18989,N_15698,N_12610);
or U18990 (N_18990,N_12892,N_14230);
nand U18991 (N_18991,N_14926,N_15708);
and U18992 (N_18992,N_15991,N_12083);
nor U18993 (N_18993,N_12766,N_15915);
nand U18994 (N_18994,N_13151,N_15874);
or U18995 (N_18995,N_12382,N_14276);
nand U18996 (N_18996,N_12332,N_12969);
xor U18997 (N_18997,N_14210,N_15602);
nor U18998 (N_18998,N_15382,N_14950);
xor U18999 (N_18999,N_13609,N_13491);
nor U19000 (N_19000,N_12660,N_13141);
and U19001 (N_19001,N_15685,N_13912);
xnor U19002 (N_19002,N_15675,N_13834);
xnor U19003 (N_19003,N_15891,N_13343);
nand U19004 (N_19004,N_13895,N_14727);
nor U19005 (N_19005,N_13141,N_15990);
nand U19006 (N_19006,N_13233,N_12907);
or U19007 (N_19007,N_13858,N_13172);
and U19008 (N_19008,N_14119,N_13384);
xnor U19009 (N_19009,N_14728,N_15185);
nand U19010 (N_19010,N_12157,N_15944);
xnor U19011 (N_19011,N_14628,N_14368);
nand U19012 (N_19012,N_13975,N_14233);
and U19013 (N_19013,N_14473,N_13211);
xor U19014 (N_19014,N_14800,N_12164);
xor U19015 (N_19015,N_15980,N_12677);
nand U19016 (N_19016,N_13345,N_14789);
and U19017 (N_19017,N_13881,N_14126);
and U19018 (N_19018,N_12966,N_13807);
or U19019 (N_19019,N_14051,N_15913);
or U19020 (N_19020,N_15556,N_13469);
and U19021 (N_19021,N_13405,N_12583);
or U19022 (N_19022,N_15403,N_15639);
nor U19023 (N_19023,N_13150,N_13049);
and U19024 (N_19024,N_14879,N_15359);
or U19025 (N_19025,N_13451,N_12709);
nand U19026 (N_19026,N_14990,N_12282);
xor U19027 (N_19027,N_14295,N_13835);
xor U19028 (N_19028,N_12464,N_13876);
nor U19029 (N_19029,N_14823,N_14844);
nand U19030 (N_19030,N_12196,N_15212);
or U19031 (N_19031,N_14286,N_14987);
xnor U19032 (N_19032,N_13852,N_14674);
xnor U19033 (N_19033,N_14633,N_13293);
or U19034 (N_19034,N_13322,N_12628);
nor U19035 (N_19035,N_12802,N_14232);
nand U19036 (N_19036,N_15740,N_14432);
and U19037 (N_19037,N_12739,N_14586);
or U19038 (N_19038,N_14757,N_13532);
nor U19039 (N_19039,N_12624,N_12727);
or U19040 (N_19040,N_12352,N_12566);
or U19041 (N_19041,N_15058,N_13792);
or U19042 (N_19042,N_13248,N_12958);
nor U19043 (N_19043,N_14227,N_13220);
xnor U19044 (N_19044,N_12194,N_13662);
or U19045 (N_19045,N_12786,N_15525);
nand U19046 (N_19046,N_12017,N_12756);
nor U19047 (N_19047,N_13888,N_15583);
or U19048 (N_19048,N_12493,N_13705);
nand U19049 (N_19049,N_15351,N_12957);
and U19050 (N_19050,N_15206,N_12198);
xnor U19051 (N_19051,N_15771,N_13069);
nand U19052 (N_19052,N_14015,N_13621);
or U19053 (N_19053,N_13264,N_15681);
nand U19054 (N_19054,N_15717,N_13355);
nand U19055 (N_19055,N_12723,N_13314);
nor U19056 (N_19056,N_13936,N_13154);
nand U19057 (N_19057,N_13829,N_13163);
xor U19058 (N_19058,N_13999,N_12512);
nor U19059 (N_19059,N_12602,N_14220);
nand U19060 (N_19060,N_13456,N_14107);
nor U19061 (N_19061,N_12429,N_15735);
nor U19062 (N_19062,N_14204,N_12185);
nor U19063 (N_19063,N_15885,N_15664);
and U19064 (N_19064,N_12741,N_13275);
nand U19065 (N_19065,N_15858,N_12498);
or U19066 (N_19066,N_15576,N_13810);
nand U19067 (N_19067,N_15643,N_12809);
xnor U19068 (N_19068,N_15472,N_15184);
or U19069 (N_19069,N_13409,N_12429);
and U19070 (N_19070,N_13618,N_15797);
or U19071 (N_19071,N_14010,N_12104);
nor U19072 (N_19072,N_14090,N_12872);
nor U19073 (N_19073,N_12330,N_13836);
and U19074 (N_19074,N_12760,N_13900);
nor U19075 (N_19075,N_15057,N_12885);
nor U19076 (N_19076,N_13788,N_15251);
nand U19077 (N_19077,N_13499,N_12498);
nor U19078 (N_19078,N_14309,N_14005);
xor U19079 (N_19079,N_13676,N_13672);
or U19080 (N_19080,N_15466,N_13509);
and U19081 (N_19081,N_12478,N_14623);
xnor U19082 (N_19082,N_13001,N_15117);
nor U19083 (N_19083,N_12902,N_14523);
or U19084 (N_19084,N_13441,N_14484);
nor U19085 (N_19085,N_12168,N_15571);
nand U19086 (N_19086,N_15492,N_14452);
or U19087 (N_19087,N_13581,N_12921);
xnor U19088 (N_19088,N_14199,N_12848);
nor U19089 (N_19089,N_15386,N_12136);
xnor U19090 (N_19090,N_13748,N_12983);
xor U19091 (N_19091,N_14316,N_15648);
nand U19092 (N_19092,N_14580,N_14381);
xnor U19093 (N_19093,N_13316,N_14148);
nand U19094 (N_19094,N_15962,N_15542);
nor U19095 (N_19095,N_13167,N_14961);
xor U19096 (N_19096,N_15003,N_14936);
or U19097 (N_19097,N_15070,N_14368);
nor U19098 (N_19098,N_14368,N_12809);
nor U19099 (N_19099,N_12404,N_14521);
and U19100 (N_19100,N_15256,N_15891);
nand U19101 (N_19101,N_15605,N_15105);
nand U19102 (N_19102,N_14379,N_14919);
or U19103 (N_19103,N_13142,N_12118);
and U19104 (N_19104,N_15908,N_13952);
xor U19105 (N_19105,N_12649,N_13434);
nor U19106 (N_19106,N_12293,N_13109);
xnor U19107 (N_19107,N_13538,N_12732);
xnor U19108 (N_19108,N_15005,N_13587);
xor U19109 (N_19109,N_15740,N_14725);
nor U19110 (N_19110,N_13488,N_13747);
nand U19111 (N_19111,N_14613,N_15516);
nand U19112 (N_19112,N_15126,N_15241);
nor U19113 (N_19113,N_12728,N_13346);
nor U19114 (N_19114,N_12359,N_12224);
or U19115 (N_19115,N_14078,N_13636);
xnor U19116 (N_19116,N_14439,N_12168);
xnor U19117 (N_19117,N_14573,N_14596);
nand U19118 (N_19118,N_12974,N_12889);
nor U19119 (N_19119,N_14718,N_14077);
nand U19120 (N_19120,N_14151,N_15625);
xor U19121 (N_19121,N_14010,N_14399);
and U19122 (N_19122,N_15023,N_12706);
nand U19123 (N_19123,N_12995,N_12566);
xnor U19124 (N_19124,N_14950,N_13827);
and U19125 (N_19125,N_12331,N_12397);
nor U19126 (N_19126,N_15893,N_12219);
and U19127 (N_19127,N_14012,N_14763);
nand U19128 (N_19128,N_15922,N_14052);
or U19129 (N_19129,N_13922,N_14902);
nor U19130 (N_19130,N_13822,N_14622);
and U19131 (N_19131,N_13556,N_14511);
or U19132 (N_19132,N_13402,N_15509);
xnor U19133 (N_19133,N_15182,N_13681);
xnor U19134 (N_19134,N_13506,N_14332);
nand U19135 (N_19135,N_12440,N_13733);
and U19136 (N_19136,N_13658,N_15500);
nor U19137 (N_19137,N_12820,N_15983);
or U19138 (N_19138,N_14722,N_15545);
nand U19139 (N_19139,N_15043,N_12481);
and U19140 (N_19140,N_14005,N_13796);
xor U19141 (N_19141,N_14694,N_12512);
nand U19142 (N_19142,N_12279,N_14437);
xor U19143 (N_19143,N_15973,N_13598);
and U19144 (N_19144,N_12342,N_15431);
nor U19145 (N_19145,N_14227,N_13800);
xnor U19146 (N_19146,N_15227,N_12095);
and U19147 (N_19147,N_12363,N_15030);
and U19148 (N_19148,N_12941,N_12322);
nor U19149 (N_19149,N_15766,N_15015);
nand U19150 (N_19150,N_15594,N_14931);
and U19151 (N_19151,N_14397,N_14989);
nand U19152 (N_19152,N_12146,N_15753);
or U19153 (N_19153,N_13018,N_13104);
nand U19154 (N_19154,N_12728,N_15756);
nand U19155 (N_19155,N_13341,N_12742);
nor U19156 (N_19156,N_12682,N_12573);
or U19157 (N_19157,N_13355,N_14237);
nand U19158 (N_19158,N_12585,N_14373);
or U19159 (N_19159,N_14003,N_12150);
or U19160 (N_19160,N_12364,N_14428);
nand U19161 (N_19161,N_14840,N_15464);
nor U19162 (N_19162,N_14616,N_15552);
nor U19163 (N_19163,N_15058,N_15091);
nand U19164 (N_19164,N_13255,N_12043);
and U19165 (N_19165,N_15521,N_13942);
nand U19166 (N_19166,N_12233,N_15721);
nand U19167 (N_19167,N_14312,N_12071);
and U19168 (N_19168,N_12642,N_13975);
nand U19169 (N_19169,N_12293,N_13387);
nand U19170 (N_19170,N_12450,N_14329);
xnor U19171 (N_19171,N_12789,N_12434);
xor U19172 (N_19172,N_14906,N_13527);
xor U19173 (N_19173,N_13534,N_12148);
or U19174 (N_19174,N_15617,N_14507);
nor U19175 (N_19175,N_15586,N_12360);
xnor U19176 (N_19176,N_12308,N_12899);
nand U19177 (N_19177,N_13776,N_14698);
nand U19178 (N_19178,N_12551,N_12600);
xor U19179 (N_19179,N_13081,N_15909);
and U19180 (N_19180,N_13257,N_12939);
nor U19181 (N_19181,N_12594,N_14184);
or U19182 (N_19182,N_13950,N_12115);
nor U19183 (N_19183,N_15620,N_14153);
or U19184 (N_19184,N_14339,N_12213);
or U19185 (N_19185,N_15826,N_15071);
xor U19186 (N_19186,N_13833,N_15278);
or U19187 (N_19187,N_15759,N_14559);
nand U19188 (N_19188,N_14081,N_15113);
and U19189 (N_19189,N_15263,N_12884);
or U19190 (N_19190,N_15694,N_12548);
and U19191 (N_19191,N_13811,N_15815);
nor U19192 (N_19192,N_13900,N_13509);
and U19193 (N_19193,N_13435,N_12033);
xor U19194 (N_19194,N_12672,N_14340);
and U19195 (N_19195,N_12260,N_12699);
nor U19196 (N_19196,N_12585,N_13526);
nand U19197 (N_19197,N_13324,N_15440);
and U19198 (N_19198,N_15718,N_13429);
xor U19199 (N_19199,N_12100,N_12392);
nand U19200 (N_19200,N_15105,N_15540);
or U19201 (N_19201,N_15877,N_14162);
nand U19202 (N_19202,N_13124,N_13152);
or U19203 (N_19203,N_15161,N_13666);
xor U19204 (N_19204,N_14840,N_14011);
nor U19205 (N_19205,N_12019,N_14750);
or U19206 (N_19206,N_15824,N_14074);
or U19207 (N_19207,N_13631,N_14919);
nand U19208 (N_19208,N_12602,N_15940);
and U19209 (N_19209,N_13363,N_14352);
and U19210 (N_19210,N_12015,N_12023);
xor U19211 (N_19211,N_12318,N_15833);
and U19212 (N_19212,N_13370,N_14408);
and U19213 (N_19213,N_13059,N_14859);
and U19214 (N_19214,N_12593,N_13319);
nor U19215 (N_19215,N_15659,N_14586);
nand U19216 (N_19216,N_15429,N_13979);
or U19217 (N_19217,N_14688,N_12263);
nor U19218 (N_19218,N_12647,N_12352);
nand U19219 (N_19219,N_12347,N_15559);
xnor U19220 (N_19220,N_15987,N_14295);
nand U19221 (N_19221,N_14135,N_14716);
or U19222 (N_19222,N_15653,N_12898);
nor U19223 (N_19223,N_12172,N_12149);
xnor U19224 (N_19224,N_14920,N_15682);
nor U19225 (N_19225,N_13806,N_12909);
or U19226 (N_19226,N_13679,N_15063);
or U19227 (N_19227,N_15539,N_14366);
xor U19228 (N_19228,N_14273,N_14099);
and U19229 (N_19229,N_12336,N_15253);
nor U19230 (N_19230,N_13189,N_14370);
xor U19231 (N_19231,N_14774,N_14404);
xor U19232 (N_19232,N_12276,N_13809);
nor U19233 (N_19233,N_15687,N_13880);
xnor U19234 (N_19234,N_14481,N_14405);
nand U19235 (N_19235,N_15687,N_13227);
or U19236 (N_19236,N_14092,N_13754);
nand U19237 (N_19237,N_12201,N_12924);
and U19238 (N_19238,N_12006,N_15099);
and U19239 (N_19239,N_14782,N_13849);
and U19240 (N_19240,N_14172,N_12314);
or U19241 (N_19241,N_13213,N_13609);
or U19242 (N_19242,N_14353,N_12348);
and U19243 (N_19243,N_13165,N_12098);
xnor U19244 (N_19244,N_15221,N_13459);
nor U19245 (N_19245,N_12553,N_15882);
nor U19246 (N_19246,N_13012,N_14042);
xor U19247 (N_19247,N_12350,N_12740);
or U19248 (N_19248,N_15471,N_14059);
and U19249 (N_19249,N_15933,N_13064);
and U19250 (N_19250,N_13634,N_12943);
xnor U19251 (N_19251,N_12191,N_14909);
nand U19252 (N_19252,N_13853,N_13817);
and U19253 (N_19253,N_15770,N_15161);
nor U19254 (N_19254,N_14263,N_12804);
or U19255 (N_19255,N_15235,N_15423);
and U19256 (N_19256,N_13388,N_15937);
or U19257 (N_19257,N_14313,N_14342);
xor U19258 (N_19258,N_14710,N_15563);
and U19259 (N_19259,N_12037,N_15876);
or U19260 (N_19260,N_12370,N_15266);
xor U19261 (N_19261,N_12905,N_13668);
or U19262 (N_19262,N_14326,N_12535);
nand U19263 (N_19263,N_12818,N_15339);
nor U19264 (N_19264,N_12899,N_14033);
or U19265 (N_19265,N_14296,N_14203);
nand U19266 (N_19266,N_14470,N_14903);
xor U19267 (N_19267,N_15732,N_15031);
or U19268 (N_19268,N_13660,N_14883);
nand U19269 (N_19269,N_14828,N_13194);
nor U19270 (N_19270,N_13523,N_15371);
and U19271 (N_19271,N_15612,N_14755);
nand U19272 (N_19272,N_12220,N_12808);
or U19273 (N_19273,N_12778,N_14094);
nor U19274 (N_19274,N_12804,N_14760);
and U19275 (N_19275,N_14693,N_12183);
nand U19276 (N_19276,N_13503,N_15116);
xnor U19277 (N_19277,N_12920,N_12679);
or U19278 (N_19278,N_12519,N_15185);
nor U19279 (N_19279,N_15757,N_15532);
and U19280 (N_19280,N_14296,N_14121);
nor U19281 (N_19281,N_15829,N_12366);
nor U19282 (N_19282,N_13014,N_15772);
and U19283 (N_19283,N_12177,N_12427);
and U19284 (N_19284,N_14632,N_13585);
and U19285 (N_19285,N_14609,N_13907);
nand U19286 (N_19286,N_14679,N_14008);
xnor U19287 (N_19287,N_15019,N_12839);
xor U19288 (N_19288,N_14499,N_15914);
nand U19289 (N_19289,N_15543,N_12860);
nand U19290 (N_19290,N_14737,N_13167);
or U19291 (N_19291,N_14481,N_13947);
xor U19292 (N_19292,N_15741,N_13307);
or U19293 (N_19293,N_14949,N_12707);
nor U19294 (N_19294,N_14735,N_12671);
xor U19295 (N_19295,N_12873,N_13367);
xor U19296 (N_19296,N_13948,N_13331);
xnor U19297 (N_19297,N_12667,N_15535);
and U19298 (N_19298,N_13886,N_12822);
and U19299 (N_19299,N_13263,N_14967);
or U19300 (N_19300,N_13683,N_15402);
or U19301 (N_19301,N_12240,N_13109);
and U19302 (N_19302,N_15260,N_14464);
xnor U19303 (N_19303,N_12203,N_13329);
nor U19304 (N_19304,N_14741,N_14591);
nor U19305 (N_19305,N_15758,N_13204);
nand U19306 (N_19306,N_13000,N_13014);
nand U19307 (N_19307,N_15476,N_13029);
and U19308 (N_19308,N_12857,N_13418);
and U19309 (N_19309,N_14915,N_14228);
nand U19310 (N_19310,N_12615,N_15410);
or U19311 (N_19311,N_15612,N_13859);
or U19312 (N_19312,N_15944,N_15824);
and U19313 (N_19313,N_12352,N_14379);
and U19314 (N_19314,N_14908,N_12646);
nand U19315 (N_19315,N_14922,N_14152);
nand U19316 (N_19316,N_14664,N_15925);
or U19317 (N_19317,N_15537,N_15749);
xor U19318 (N_19318,N_14117,N_12386);
xor U19319 (N_19319,N_13017,N_14571);
xor U19320 (N_19320,N_13882,N_14714);
nand U19321 (N_19321,N_12214,N_12906);
or U19322 (N_19322,N_15757,N_13329);
nand U19323 (N_19323,N_14665,N_14939);
and U19324 (N_19324,N_15803,N_12480);
and U19325 (N_19325,N_13356,N_12027);
or U19326 (N_19326,N_15055,N_12310);
and U19327 (N_19327,N_12486,N_12937);
xor U19328 (N_19328,N_12721,N_15481);
nand U19329 (N_19329,N_12121,N_13274);
or U19330 (N_19330,N_15088,N_15068);
or U19331 (N_19331,N_14225,N_12478);
xnor U19332 (N_19332,N_15101,N_14665);
nor U19333 (N_19333,N_12638,N_15429);
nor U19334 (N_19334,N_12445,N_12969);
and U19335 (N_19335,N_13657,N_15100);
and U19336 (N_19336,N_13159,N_13396);
nand U19337 (N_19337,N_12023,N_14102);
xor U19338 (N_19338,N_12916,N_15782);
xor U19339 (N_19339,N_14017,N_15354);
and U19340 (N_19340,N_15733,N_14941);
nor U19341 (N_19341,N_14041,N_12066);
and U19342 (N_19342,N_12556,N_15302);
nand U19343 (N_19343,N_14850,N_14953);
nand U19344 (N_19344,N_13771,N_12609);
nor U19345 (N_19345,N_14373,N_12060);
xnor U19346 (N_19346,N_13665,N_15962);
or U19347 (N_19347,N_12252,N_15776);
nor U19348 (N_19348,N_13874,N_15148);
nor U19349 (N_19349,N_15125,N_15884);
nand U19350 (N_19350,N_15461,N_12094);
or U19351 (N_19351,N_12420,N_13092);
and U19352 (N_19352,N_14214,N_13301);
xnor U19353 (N_19353,N_15423,N_12036);
and U19354 (N_19354,N_13722,N_13215);
nor U19355 (N_19355,N_15402,N_15717);
and U19356 (N_19356,N_14965,N_12451);
nand U19357 (N_19357,N_14835,N_15536);
xnor U19358 (N_19358,N_12769,N_15698);
or U19359 (N_19359,N_13412,N_13274);
nand U19360 (N_19360,N_13334,N_14128);
nand U19361 (N_19361,N_15903,N_14178);
nor U19362 (N_19362,N_12401,N_14513);
and U19363 (N_19363,N_14413,N_14927);
and U19364 (N_19364,N_15783,N_13065);
nand U19365 (N_19365,N_12042,N_14601);
or U19366 (N_19366,N_13212,N_13706);
nand U19367 (N_19367,N_15233,N_12837);
xor U19368 (N_19368,N_12602,N_13126);
xor U19369 (N_19369,N_13583,N_13521);
nor U19370 (N_19370,N_13351,N_12505);
xor U19371 (N_19371,N_15915,N_12597);
nor U19372 (N_19372,N_12603,N_14359);
nor U19373 (N_19373,N_14953,N_15045);
xor U19374 (N_19374,N_13848,N_12518);
nor U19375 (N_19375,N_14515,N_15517);
xnor U19376 (N_19376,N_12952,N_15595);
and U19377 (N_19377,N_12248,N_12783);
or U19378 (N_19378,N_15598,N_14260);
xnor U19379 (N_19379,N_13116,N_13489);
nor U19380 (N_19380,N_15958,N_12586);
or U19381 (N_19381,N_12388,N_12140);
or U19382 (N_19382,N_14731,N_13012);
nor U19383 (N_19383,N_14549,N_15384);
and U19384 (N_19384,N_14603,N_15046);
and U19385 (N_19385,N_15000,N_12284);
nand U19386 (N_19386,N_12134,N_12472);
and U19387 (N_19387,N_15562,N_15406);
nand U19388 (N_19388,N_14968,N_14465);
or U19389 (N_19389,N_14101,N_12155);
and U19390 (N_19390,N_15458,N_13969);
nand U19391 (N_19391,N_13953,N_13727);
nor U19392 (N_19392,N_12732,N_14014);
and U19393 (N_19393,N_14727,N_12513);
nand U19394 (N_19394,N_13363,N_12632);
xor U19395 (N_19395,N_14978,N_12427);
nor U19396 (N_19396,N_15636,N_12754);
xnor U19397 (N_19397,N_12986,N_12132);
and U19398 (N_19398,N_12799,N_15847);
or U19399 (N_19399,N_15501,N_13198);
and U19400 (N_19400,N_14816,N_13502);
and U19401 (N_19401,N_14300,N_12290);
or U19402 (N_19402,N_12312,N_14741);
and U19403 (N_19403,N_13249,N_14739);
and U19404 (N_19404,N_14939,N_15202);
nand U19405 (N_19405,N_12676,N_12608);
nor U19406 (N_19406,N_12174,N_13990);
xnor U19407 (N_19407,N_12180,N_15670);
nor U19408 (N_19408,N_13207,N_13181);
or U19409 (N_19409,N_14330,N_15527);
or U19410 (N_19410,N_12598,N_15750);
and U19411 (N_19411,N_14989,N_12020);
and U19412 (N_19412,N_15431,N_15081);
or U19413 (N_19413,N_15372,N_14056);
nor U19414 (N_19414,N_14340,N_14822);
or U19415 (N_19415,N_15006,N_15827);
xor U19416 (N_19416,N_15379,N_14708);
nand U19417 (N_19417,N_14606,N_12359);
or U19418 (N_19418,N_14618,N_13866);
nand U19419 (N_19419,N_15870,N_14604);
or U19420 (N_19420,N_13618,N_14573);
nand U19421 (N_19421,N_12426,N_15248);
or U19422 (N_19422,N_14595,N_12670);
xor U19423 (N_19423,N_13871,N_13531);
xor U19424 (N_19424,N_12430,N_12418);
or U19425 (N_19425,N_15178,N_14307);
nand U19426 (N_19426,N_12573,N_12994);
or U19427 (N_19427,N_14743,N_13716);
nand U19428 (N_19428,N_13234,N_12487);
and U19429 (N_19429,N_12459,N_15144);
xor U19430 (N_19430,N_14108,N_14974);
nand U19431 (N_19431,N_12944,N_12531);
xor U19432 (N_19432,N_14189,N_14921);
and U19433 (N_19433,N_14095,N_14134);
nand U19434 (N_19434,N_13385,N_13469);
xnor U19435 (N_19435,N_15720,N_12852);
or U19436 (N_19436,N_15710,N_12417);
or U19437 (N_19437,N_15814,N_14916);
nand U19438 (N_19438,N_12064,N_12686);
nand U19439 (N_19439,N_13827,N_14370);
nor U19440 (N_19440,N_14369,N_15596);
xor U19441 (N_19441,N_14014,N_15940);
xor U19442 (N_19442,N_12308,N_15472);
nand U19443 (N_19443,N_13206,N_13467);
or U19444 (N_19444,N_12197,N_12837);
xor U19445 (N_19445,N_13989,N_12691);
xnor U19446 (N_19446,N_14510,N_13419);
xor U19447 (N_19447,N_12597,N_13130);
and U19448 (N_19448,N_14425,N_15337);
or U19449 (N_19449,N_14454,N_15157);
nand U19450 (N_19450,N_12907,N_12072);
and U19451 (N_19451,N_14245,N_15963);
nor U19452 (N_19452,N_12337,N_13860);
or U19453 (N_19453,N_13566,N_13438);
nor U19454 (N_19454,N_15691,N_15112);
nand U19455 (N_19455,N_12786,N_15496);
nand U19456 (N_19456,N_13439,N_12680);
xnor U19457 (N_19457,N_12781,N_13469);
or U19458 (N_19458,N_15979,N_15218);
xnor U19459 (N_19459,N_14608,N_15387);
xnor U19460 (N_19460,N_14688,N_13251);
or U19461 (N_19461,N_12918,N_12252);
or U19462 (N_19462,N_12877,N_14567);
nor U19463 (N_19463,N_15198,N_12689);
nor U19464 (N_19464,N_15837,N_15013);
nand U19465 (N_19465,N_15417,N_15537);
nor U19466 (N_19466,N_15568,N_15655);
or U19467 (N_19467,N_13233,N_13035);
nor U19468 (N_19468,N_13227,N_15590);
nor U19469 (N_19469,N_14429,N_14448);
or U19470 (N_19470,N_14971,N_12164);
nand U19471 (N_19471,N_13557,N_12472);
xor U19472 (N_19472,N_13921,N_15041);
nor U19473 (N_19473,N_13789,N_15975);
xnor U19474 (N_19474,N_13866,N_14263);
nand U19475 (N_19475,N_13674,N_15671);
and U19476 (N_19476,N_13981,N_13069);
nand U19477 (N_19477,N_12564,N_14254);
nand U19478 (N_19478,N_14742,N_15374);
or U19479 (N_19479,N_12368,N_13156);
xnor U19480 (N_19480,N_15709,N_14070);
nor U19481 (N_19481,N_14702,N_13518);
nor U19482 (N_19482,N_14068,N_14405);
and U19483 (N_19483,N_13263,N_13194);
or U19484 (N_19484,N_15609,N_13634);
and U19485 (N_19485,N_13338,N_15305);
xnor U19486 (N_19486,N_15962,N_15594);
xor U19487 (N_19487,N_14108,N_13397);
and U19488 (N_19488,N_13070,N_12257);
and U19489 (N_19489,N_14281,N_15614);
nand U19490 (N_19490,N_13410,N_14025);
or U19491 (N_19491,N_13717,N_12846);
nand U19492 (N_19492,N_15101,N_12368);
nand U19493 (N_19493,N_15941,N_14016);
or U19494 (N_19494,N_13365,N_13287);
nor U19495 (N_19495,N_12130,N_15792);
and U19496 (N_19496,N_14921,N_14728);
nor U19497 (N_19497,N_14940,N_14812);
and U19498 (N_19498,N_14926,N_12650);
xnor U19499 (N_19499,N_15582,N_12415);
xnor U19500 (N_19500,N_14469,N_15002);
or U19501 (N_19501,N_14824,N_12352);
and U19502 (N_19502,N_14361,N_15688);
and U19503 (N_19503,N_14350,N_12395);
nor U19504 (N_19504,N_12348,N_14866);
nor U19505 (N_19505,N_14407,N_15249);
nor U19506 (N_19506,N_13528,N_12969);
nand U19507 (N_19507,N_14576,N_15337);
nand U19508 (N_19508,N_13757,N_14599);
nand U19509 (N_19509,N_14098,N_13133);
xnor U19510 (N_19510,N_15187,N_15175);
xor U19511 (N_19511,N_15000,N_15376);
and U19512 (N_19512,N_13363,N_14870);
or U19513 (N_19513,N_15319,N_15538);
xor U19514 (N_19514,N_14735,N_12524);
and U19515 (N_19515,N_13018,N_15451);
nand U19516 (N_19516,N_13539,N_12031);
or U19517 (N_19517,N_14734,N_13794);
xnor U19518 (N_19518,N_14064,N_15931);
xnor U19519 (N_19519,N_14330,N_15997);
xor U19520 (N_19520,N_13639,N_13605);
nor U19521 (N_19521,N_14219,N_15872);
xnor U19522 (N_19522,N_14676,N_13352);
or U19523 (N_19523,N_12836,N_15818);
and U19524 (N_19524,N_13289,N_12998);
nand U19525 (N_19525,N_12671,N_14412);
and U19526 (N_19526,N_12757,N_14634);
or U19527 (N_19527,N_13336,N_14543);
and U19528 (N_19528,N_13295,N_13614);
or U19529 (N_19529,N_13945,N_15495);
nor U19530 (N_19530,N_14578,N_14959);
and U19531 (N_19531,N_13583,N_14277);
or U19532 (N_19532,N_14405,N_15534);
nand U19533 (N_19533,N_14383,N_14610);
or U19534 (N_19534,N_12567,N_15339);
nand U19535 (N_19535,N_13061,N_12503);
nand U19536 (N_19536,N_14467,N_13316);
and U19537 (N_19537,N_14643,N_13687);
nor U19538 (N_19538,N_15920,N_12605);
or U19539 (N_19539,N_13241,N_12986);
nor U19540 (N_19540,N_14451,N_14002);
nor U19541 (N_19541,N_12517,N_13396);
nand U19542 (N_19542,N_14845,N_15867);
nor U19543 (N_19543,N_13799,N_14271);
or U19544 (N_19544,N_13245,N_15916);
or U19545 (N_19545,N_13990,N_15133);
nor U19546 (N_19546,N_13985,N_14573);
xnor U19547 (N_19547,N_13524,N_15459);
nand U19548 (N_19548,N_13149,N_15810);
or U19549 (N_19549,N_13885,N_15119);
xnor U19550 (N_19550,N_14245,N_15868);
nor U19551 (N_19551,N_14576,N_12728);
nor U19552 (N_19552,N_14835,N_12383);
nor U19553 (N_19553,N_12628,N_12233);
nand U19554 (N_19554,N_14105,N_15245);
nor U19555 (N_19555,N_15060,N_15571);
xor U19556 (N_19556,N_13057,N_12768);
or U19557 (N_19557,N_15907,N_14595);
or U19558 (N_19558,N_15341,N_12074);
or U19559 (N_19559,N_15801,N_14850);
or U19560 (N_19560,N_15677,N_14722);
xnor U19561 (N_19561,N_12543,N_15959);
nor U19562 (N_19562,N_13306,N_12340);
and U19563 (N_19563,N_12919,N_15170);
nor U19564 (N_19564,N_15274,N_14221);
nand U19565 (N_19565,N_15091,N_12157);
nand U19566 (N_19566,N_14774,N_14330);
xor U19567 (N_19567,N_15287,N_13166);
xnor U19568 (N_19568,N_13031,N_15081);
and U19569 (N_19569,N_15254,N_15512);
and U19570 (N_19570,N_15339,N_12586);
nor U19571 (N_19571,N_14309,N_13220);
and U19572 (N_19572,N_12899,N_15832);
and U19573 (N_19573,N_13393,N_15948);
nor U19574 (N_19574,N_13882,N_14399);
and U19575 (N_19575,N_13395,N_13617);
xnor U19576 (N_19576,N_14765,N_12033);
xnor U19577 (N_19577,N_13959,N_15294);
nor U19578 (N_19578,N_13598,N_14620);
or U19579 (N_19579,N_13045,N_12601);
nand U19580 (N_19580,N_13248,N_13067);
nor U19581 (N_19581,N_12411,N_13858);
or U19582 (N_19582,N_14415,N_12993);
or U19583 (N_19583,N_15218,N_13150);
or U19584 (N_19584,N_14586,N_13031);
nor U19585 (N_19585,N_14640,N_12606);
nand U19586 (N_19586,N_15809,N_15678);
and U19587 (N_19587,N_12408,N_13178);
xor U19588 (N_19588,N_15948,N_14193);
nand U19589 (N_19589,N_13255,N_14758);
nand U19590 (N_19590,N_15870,N_14845);
xor U19591 (N_19591,N_12804,N_12474);
nand U19592 (N_19592,N_13854,N_12993);
nor U19593 (N_19593,N_12436,N_12490);
xor U19594 (N_19594,N_15618,N_12196);
and U19595 (N_19595,N_15819,N_13629);
nand U19596 (N_19596,N_13887,N_15271);
nor U19597 (N_19597,N_13300,N_14633);
or U19598 (N_19598,N_15874,N_15382);
and U19599 (N_19599,N_14923,N_15428);
and U19600 (N_19600,N_15604,N_15266);
or U19601 (N_19601,N_14984,N_15957);
xor U19602 (N_19602,N_13115,N_14991);
nand U19603 (N_19603,N_12845,N_12823);
xor U19604 (N_19604,N_13227,N_14696);
or U19605 (N_19605,N_15275,N_14132);
or U19606 (N_19606,N_13285,N_14669);
nor U19607 (N_19607,N_14638,N_15260);
or U19608 (N_19608,N_15437,N_13494);
nand U19609 (N_19609,N_13088,N_15575);
nand U19610 (N_19610,N_14050,N_14766);
or U19611 (N_19611,N_12248,N_13997);
xor U19612 (N_19612,N_13555,N_12878);
and U19613 (N_19613,N_13785,N_14358);
nor U19614 (N_19614,N_12206,N_14731);
nand U19615 (N_19615,N_15131,N_15977);
nand U19616 (N_19616,N_15221,N_15491);
or U19617 (N_19617,N_12236,N_12476);
and U19618 (N_19618,N_15429,N_14520);
and U19619 (N_19619,N_13091,N_12147);
nand U19620 (N_19620,N_13645,N_13922);
nor U19621 (N_19621,N_14374,N_12669);
or U19622 (N_19622,N_15738,N_12928);
or U19623 (N_19623,N_13859,N_12710);
or U19624 (N_19624,N_14082,N_14390);
xnor U19625 (N_19625,N_13057,N_13060);
and U19626 (N_19626,N_13568,N_13421);
and U19627 (N_19627,N_13594,N_15069);
nand U19628 (N_19628,N_15072,N_13085);
or U19629 (N_19629,N_14642,N_15165);
or U19630 (N_19630,N_12270,N_12991);
or U19631 (N_19631,N_15919,N_13095);
nand U19632 (N_19632,N_14205,N_13733);
and U19633 (N_19633,N_13253,N_14711);
or U19634 (N_19634,N_14893,N_14223);
nor U19635 (N_19635,N_15923,N_13967);
or U19636 (N_19636,N_15789,N_14655);
and U19637 (N_19637,N_14324,N_14148);
xor U19638 (N_19638,N_12036,N_12237);
and U19639 (N_19639,N_13929,N_15380);
nor U19640 (N_19640,N_13271,N_15688);
nand U19641 (N_19641,N_14730,N_14995);
nand U19642 (N_19642,N_14463,N_12362);
or U19643 (N_19643,N_15842,N_14493);
and U19644 (N_19644,N_12770,N_15736);
and U19645 (N_19645,N_12245,N_14691);
nor U19646 (N_19646,N_12566,N_14192);
xnor U19647 (N_19647,N_14604,N_15584);
or U19648 (N_19648,N_12010,N_14868);
or U19649 (N_19649,N_13116,N_13366);
xnor U19650 (N_19650,N_13185,N_13796);
nor U19651 (N_19651,N_13892,N_12035);
xnor U19652 (N_19652,N_15544,N_14049);
nor U19653 (N_19653,N_13034,N_15488);
nor U19654 (N_19654,N_15605,N_14213);
nand U19655 (N_19655,N_15476,N_12241);
xnor U19656 (N_19656,N_12119,N_12460);
nand U19657 (N_19657,N_12120,N_12331);
and U19658 (N_19658,N_15995,N_14773);
nor U19659 (N_19659,N_15308,N_14489);
and U19660 (N_19660,N_12680,N_14679);
nand U19661 (N_19661,N_15345,N_15651);
or U19662 (N_19662,N_12167,N_14170);
nand U19663 (N_19663,N_12696,N_15340);
or U19664 (N_19664,N_13802,N_13513);
xnor U19665 (N_19665,N_15314,N_15495);
xnor U19666 (N_19666,N_14307,N_15403);
and U19667 (N_19667,N_12803,N_15265);
nor U19668 (N_19668,N_12258,N_13425);
nand U19669 (N_19669,N_14624,N_15436);
and U19670 (N_19670,N_15502,N_12919);
nand U19671 (N_19671,N_12990,N_14963);
and U19672 (N_19672,N_14995,N_15618);
xor U19673 (N_19673,N_12018,N_12663);
and U19674 (N_19674,N_14400,N_12176);
nor U19675 (N_19675,N_13119,N_14928);
or U19676 (N_19676,N_12724,N_12989);
or U19677 (N_19677,N_15353,N_14831);
or U19678 (N_19678,N_15467,N_13780);
and U19679 (N_19679,N_15886,N_13750);
or U19680 (N_19680,N_12805,N_13402);
and U19681 (N_19681,N_13202,N_12828);
nor U19682 (N_19682,N_14027,N_14272);
and U19683 (N_19683,N_14741,N_15647);
nor U19684 (N_19684,N_14371,N_12215);
xnor U19685 (N_19685,N_15986,N_14390);
or U19686 (N_19686,N_15595,N_13414);
xnor U19687 (N_19687,N_15507,N_15071);
xor U19688 (N_19688,N_13150,N_13113);
and U19689 (N_19689,N_12644,N_13661);
nand U19690 (N_19690,N_15472,N_14627);
nand U19691 (N_19691,N_14823,N_15432);
nand U19692 (N_19692,N_15035,N_13113);
xor U19693 (N_19693,N_15753,N_14139);
and U19694 (N_19694,N_14120,N_13054);
or U19695 (N_19695,N_12036,N_13191);
or U19696 (N_19696,N_14230,N_14418);
nand U19697 (N_19697,N_15660,N_14041);
xor U19698 (N_19698,N_13204,N_13505);
nand U19699 (N_19699,N_13597,N_13340);
xor U19700 (N_19700,N_14794,N_15075);
and U19701 (N_19701,N_14248,N_14570);
xor U19702 (N_19702,N_12780,N_12825);
nor U19703 (N_19703,N_12239,N_15888);
xor U19704 (N_19704,N_12444,N_14026);
and U19705 (N_19705,N_13799,N_14019);
nand U19706 (N_19706,N_13719,N_15590);
xnor U19707 (N_19707,N_13721,N_12774);
xor U19708 (N_19708,N_13101,N_13929);
and U19709 (N_19709,N_15862,N_13727);
and U19710 (N_19710,N_15135,N_14939);
and U19711 (N_19711,N_14061,N_13678);
xor U19712 (N_19712,N_13810,N_15161);
nand U19713 (N_19713,N_13687,N_15085);
nor U19714 (N_19714,N_12387,N_12660);
xnor U19715 (N_19715,N_15543,N_14199);
xnor U19716 (N_19716,N_15130,N_14197);
xnor U19717 (N_19717,N_15107,N_13555);
nand U19718 (N_19718,N_12337,N_14852);
and U19719 (N_19719,N_13616,N_12183);
or U19720 (N_19720,N_14626,N_15335);
nor U19721 (N_19721,N_13594,N_14915);
or U19722 (N_19722,N_14892,N_13723);
and U19723 (N_19723,N_14666,N_13047);
nor U19724 (N_19724,N_13212,N_12849);
xnor U19725 (N_19725,N_14122,N_12127);
nor U19726 (N_19726,N_13395,N_12525);
nand U19727 (N_19727,N_13129,N_12424);
and U19728 (N_19728,N_14047,N_13979);
xor U19729 (N_19729,N_13840,N_15307);
nor U19730 (N_19730,N_13662,N_13423);
nor U19731 (N_19731,N_14546,N_13795);
or U19732 (N_19732,N_14990,N_14481);
or U19733 (N_19733,N_15960,N_13430);
nor U19734 (N_19734,N_15754,N_15344);
or U19735 (N_19735,N_15477,N_12045);
nor U19736 (N_19736,N_12368,N_14876);
nand U19737 (N_19737,N_13716,N_12994);
or U19738 (N_19738,N_12263,N_14707);
xor U19739 (N_19739,N_13394,N_15347);
nand U19740 (N_19740,N_14302,N_15796);
and U19741 (N_19741,N_13916,N_13264);
and U19742 (N_19742,N_12006,N_15930);
xnor U19743 (N_19743,N_14616,N_12363);
nor U19744 (N_19744,N_13739,N_13516);
nand U19745 (N_19745,N_13856,N_12512);
xnor U19746 (N_19746,N_12289,N_14181);
and U19747 (N_19747,N_12429,N_15794);
nand U19748 (N_19748,N_13354,N_12188);
xnor U19749 (N_19749,N_15834,N_15901);
nand U19750 (N_19750,N_14927,N_13979);
xor U19751 (N_19751,N_15287,N_12296);
or U19752 (N_19752,N_12290,N_12278);
nand U19753 (N_19753,N_13800,N_15864);
nand U19754 (N_19754,N_12349,N_15824);
xor U19755 (N_19755,N_15448,N_13839);
nand U19756 (N_19756,N_15421,N_13621);
and U19757 (N_19757,N_13174,N_14170);
and U19758 (N_19758,N_15193,N_14967);
and U19759 (N_19759,N_15563,N_13714);
nand U19760 (N_19760,N_15270,N_15787);
and U19761 (N_19761,N_12747,N_13245);
nand U19762 (N_19762,N_15015,N_12949);
nand U19763 (N_19763,N_12247,N_15510);
nor U19764 (N_19764,N_14909,N_15340);
and U19765 (N_19765,N_12611,N_14768);
xnor U19766 (N_19766,N_15661,N_12893);
and U19767 (N_19767,N_12098,N_12613);
and U19768 (N_19768,N_13131,N_14996);
nor U19769 (N_19769,N_13438,N_13807);
nor U19770 (N_19770,N_15486,N_13628);
nand U19771 (N_19771,N_13274,N_13542);
nand U19772 (N_19772,N_14906,N_12139);
nor U19773 (N_19773,N_13102,N_13397);
and U19774 (N_19774,N_15209,N_14576);
nor U19775 (N_19775,N_12304,N_15498);
nand U19776 (N_19776,N_15263,N_12452);
nor U19777 (N_19777,N_15132,N_12106);
nor U19778 (N_19778,N_14709,N_13036);
and U19779 (N_19779,N_15801,N_14679);
or U19780 (N_19780,N_13048,N_15050);
or U19781 (N_19781,N_12607,N_13608);
xnor U19782 (N_19782,N_15702,N_14899);
nand U19783 (N_19783,N_15172,N_13414);
nor U19784 (N_19784,N_12468,N_13153);
xor U19785 (N_19785,N_15963,N_13980);
and U19786 (N_19786,N_12345,N_12331);
nor U19787 (N_19787,N_14026,N_15763);
nand U19788 (N_19788,N_12913,N_14980);
nand U19789 (N_19789,N_14092,N_12829);
or U19790 (N_19790,N_12634,N_15131);
xor U19791 (N_19791,N_15166,N_14109);
and U19792 (N_19792,N_13129,N_15641);
nor U19793 (N_19793,N_12274,N_14212);
nor U19794 (N_19794,N_12856,N_14033);
nor U19795 (N_19795,N_13832,N_15872);
nor U19796 (N_19796,N_12338,N_15497);
nor U19797 (N_19797,N_12677,N_12486);
and U19798 (N_19798,N_12000,N_15801);
or U19799 (N_19799,N_14348,N_14032);
and U19800 (N_19800,N_14644,N_13294);
xor U19801 (N_19801,N_13250,N_15883);
and U19802 (N_19802,N_15925,N_12661);
or U19803 (N_19803,N_14342,N_12854);
nor U19804 (N_19804,N_15666,N_14159);
and U19805 (N_19805,N_15294,N_12397);
xnor U19806 (N_19806,N_14931,N_12595);
or U19807 (N_19807,N_15719,N_13456);
nand U19808 (N_19808,N_14972,N_13269);
xor U19809 (N_19809,N_15724,N_14461);
nand U19810 (N_19810,N_14636,N_13395);
or U19811 (N_19811,N_14567,N_13422);
and U19812 (N_19812,N_15699,N_15308);
nor U19813 (N_19813,N_13993,N_15408);
or U19814 (N_19814,N_15560,N_15123);
and U19815 (N_19815,N_14382,N_13277);
nand U19816 (N_19816,N_15542,N_15950);
nor U19817 (N_19817,N_14834,N_14916);
nor U19818 (N_19818,N_15447,N_15583);
or U19819 (N_19819,N_15079,N_12197);
nand U19820 (N_19820,N_13050,N_14904);
nor U19821 (N_19821,N_14619,N_12332);
xor U19822 (N_19822,N_15359,N_12127);
xnor U19823 (N_19823,N_13671,N_13358);
or U19824 (N_19824,N_15458,N_15406);
nor U19825 (N_19825,N_14515,N_12859);
or U19826 (N_19826,N_15575,N_14738);
xnor U19827 (N_19827,N_13219,N_15111);
xor U19828 (N_19828,N_14965,N_15519);
nand U19829 (N_19829,N_12910,N_12004);
and U19830 (N_19830,N_13956,N_13495);
xor U19831 (N_19831,N_12809,N_12725);
or U19832 (N_19832,N_14700,N_15227);
nor U19833 (N_19833,N_14333,N_14279);
xor U19834 (N_19834,N_15385,N_13796);
and U19835 (N_19835,N_14430,N_14226);
or U19836 (N_19836,N_12923,N_13880);
or U19837 (N_19837,N_15396,N_12806);
and U19838 (N_19838,N_14295,N_13227);
xor U19839 (N_19839,N_15968,N_13920);
nand U19840 (N_19840,N_12203,N_15375);
nor U19841 (N_19841,N_14031,N_12663);
nand U19842 (N_19842,N_13142,N_15535);
nor U19843 (N_19843,N_14007,N_14561);
nor U19844 (N_19844,N_13335,N_13426);
nand U19845 (N_19845,N_13061,N_15150);
and U19846 (N_19846,N_14008,N_13523);
nand U19847 (N_19847,N_14574,N_13094);
nor U19848 (N_19848,N_13791,N_14686);
xor U19849 (N_19849,N_14246,N_12527);
and U19850 (N_19850,N_12633,N_15353);
xnor U19851 (N_19851,N_12596,N_15281);
and U19852 (N_19852,N_15782,N_15935);
and U19853 (N_19853,N_15888,N_12067);
and U19854 (N_19854,N_15856,N_15298);
xor U19855 (N_19855,N_12984,N_12897);
xnor U19856 (N_19856,N_12968,N_13861);
or U19857 (N_19857,N_12137,N_15320);
nor U19858 (N_19858,N_14029,N_12799);
or U19859 (N_19859,N_13620,N_15747);
or U19860 (N_19860,N_14951,N_14672);
xor U19861 (N_19861,N_13410,N_14103);
and U19862 (N_19862,N_14187,N_14231);
nor U19863 (N_19863,N_13620,N_15552);
xor U19864 (N_19864,N_15617,N_13184);
nand U19865 (N_19865,N_14856,N_14740);
nand U19866 (N_19866,N_12784,N_15229);
and U19867 (N_19867,N_13457,N_15361);
xor U19868 (N_19868,N_14646,N_14657);
xor U19869 (N_19869,N_12535,N_13470);
xor U19870 (N_19870,N_13518,N_12818);
and U19871 (N_19871,N_12989,N_15087);
xor U19872 (N_19872,N_14199,N_12932);
and U19873 (N_19873,N_13070,N_13854);
nor U19874 (N_19874,N_15114,N_13465);
nor U19875 (N_19875,N_15100,N_14851);
xnor U19876 (N_19876,N_15363,N_13049);
nand U19877 (N_19877,N_12487,N_12862);
xor U19878 (N_19878,N_15265,N_12648);
or U19879 (N_19879,N_13500,N_13878);
or U19880 (N_19880,N_13438,N_15971);
and U19881 (N_19881,N_12172,N_12296);
nor U19882 (N_19882,N_14902,N_14914);
nand U19883 (N_19883,N_13688,N_15370);
xnor U19884 (N_19884,N_14989,N_15650);
or U19885 (N_19885,N_15283,N_12842);
and U19886 (N_19886,N_15253,N_13024);
nand U19887 (N_19887,N_12027,N_12621);
xor U19888 (N_19888,N_14710,N_15974);
nor U19889 (N_19889,N_13360,N_15580);
nand U19890 (N_19890,N_13370,N_13172);
or U19891 (N_19891,N_15336,N_12404);
or U19892 (N_19892,N_14571,N_12560);
and U19893 (N_19893,N_12691,N_12636);
nand U19894 (N_19894,N_14850,N_12410);
and U19895 (N_19895,N_13335,N_13774);
nor U19896 (N_19896,N_15941,N_13907);
nor U19897 (N_19897,N_15166,N_15395);
nand U19898 (N_19898,N_13030,N_14266);
or U19899 (N_19899,N_12391,N_13562);
nand U19900 (N_19900,N_15101,N_12705);
and U19901 (N_19901,N_12849,N_13613);
and U19902 (N_19902,N_13770,N_13845);
xor U19903 (N_19903,N_13317,N_13444);
nand U19904 (N_19904,N_14748,N_12940);
nor U19905 (N_19905,N_13416,N_13189);
or U19906 (N_19906,N_13263,N_15794);
or U19907 (N_19907,N_13062,N_12786);
or U19908 (N_19908,N_15072,N_15337);
or U19909 (N_19909,N_13076,N_14960);
nand U19910 (N_19910,N_15378,N_15639);
nand U19911 (N_19911,N_13769,N_14332);
nand U19912 (N_19912,N_15913,N_14704);
nand U19913 (N_19913,N_12692,N_14434);
xnor U19914 (N_19914,N_12111,N_13040);
and U19915 (N_19915,N_12495,N_15950);
or U19916 (N_19916,N_15434,N_12676);
or U19917 (N_19917,N_13769,N_14974);
nor U19918 (N_19918,N_15612,N_12502);
or U19919 (N_19919,N_14053,N_14441);
xnor U19920 (N_19920,N_14597,N_12449);
nand U19921 (N_19921,N_12895,N_13818);
or U19922 (N_19922,N_13563,N_15848);
and U19923 (N_19923,N_14752,N_15798);
and U19924 (N_19924,N_12496,N_14348);
and U19925 (N_19925,N_14388,N_12724);
xnor U19926 (N_19926,N_14949,N_14905);
and U19927 (N_19927,N_13890,N_13830);
nor U19928 (N_19928,N_13814,N_14243);
nand U19929 (N_19929,N_15239,N_15255);
nand U19930 (N_19930,N_13511,N_14726);
and U19931 (N_19931,N_14491,N_12338);
or U19932 (N_19932,N_15611,N_13579);
and U19933 (N_19933,N_14644,N_13466);
or U19934 (N_19934,N_15348,N_15808);
xor U19935 (N_19935,N_12733,N_12681);
nor U19936 (N_19936,N_13098,N_12140);
and U19937 (N_19937,N_15585,N_15372);
or U19938 (N_19938,N_13926,N_14552);
nand U19939 (N_19939,N_13270,N_15304);
or U19940 (N_19940,N_14897,N_15743);
and U19941 (N_19941,N_12113,N_14549);
xnor U19942 (N_19942,N_14651,N_15967);
and U19943 (N_19943,N_15232,N_12571);
and U19944 (N_19944,N_13831,N_15911);
nor U19945 (N_19945,N_13585,N_14446);
or U19946 (N_19946,N_13265,N_13767);
xor U19947 (N_19947,N_15749,N_15000);
nor U19948 (N_19948,N_15388,N_13414);
nand U19949 (N_19949,N_14669,N_12497);
or U19950 (N_19950,N_15281,N_13796);
nand U19951 (N_19951,N_13620,N_13878);
nor U19952 (N_19952,N_12992,N_12200);
nor U19953 (N_19953,N_13147,N_13680);
or U19954 (N_19954,N_13624,N_15959);
nand U19955 (N_19955,N_13478,N_12411);
nor U19956 (N_19956,N_14713,N_14069);
and U19957 (N_19957,N_15159,N_15710);
xor U19958 (N_19958,N_14938,N_14747);
or U19959 (N_19959,N_13945,N_15302);
or U19960 (N_19960,N_12156,N_15025);
nor U19961 (N_19961,N_15439,N_15367);
and U19962 (N_19962,N_12122,N_12584);
and U19963 (N_19963,N_13487,N_12399);
nand U19964 (N_19964,N_12450,N_14391);
nor U19965 (N_19965,N_14372,N_14008);
nor U19966 (N_19966,N_14694,N_12867);
and U19967 (N_19967,N_13131,N_14259);
nand U19968 (N_19968,N_14558,N_13476);
nor U19969 (N_19969,N_12037,N_13618);
nand U19970 (N_19970,N_14114,N_12958);
or U19971 (N_19971,N_12221,N_14615);
and U19972 (N_19972,N_13537,N_14614);
and U19973 (N_19973,N_15583,N_15191);
or U19974 (N_19974,N_12255,N_15258);
and U19975 (N_19975,N_14104,N_14496);
xnor U19976 (N_19976,N_15726,N_12127);
nand U19977 (N_19977,N_13228,N_15611);
xnor U19978 (N_19978,N_13333,N_12647);
nand U19979 (N_19979,N_12866,N_14292);
and U19980 (N_19980,N_14414,N_13741);
or U19981 (N_19981,N_12174,N_13795);
and U19982 (N_19982,N_15339,N_13305);
and U19983 (N_19983,N_15941,N_15623);
or U19984 (N_19984,N_15971,N_15136);
nand U19985 (N_19985,N_12895,N_15508);
nor U19986 (N_19986,N_15458,N_12218);
xnor U19987 (N_19987,N_13681,N_14432);
and U19988 (N_19988,N_15741,N_14960);
nor U19989 (N_19989,N_15519,N_14325);
nand U19990 (N_19990,N_12921,N_15554);
or U19991 (N_19991,N_14723,N_12238);
nor U19992 (N_19992,N_14193,N_12376);
or U19993 (N_19993,N_12482,N_13005);
nor U19994 (N_19994,N_13809,N_12904);
or U19995 (N_19995,N_14028,N_12262);
or U19996 (N_19996,N_14005,N_14203);
nor U19997 (N_19997,N_14540,N_14200);
or U19998 (N_19998,N_15244,N_14799);
xor U19999 (N_19999,N_13119,N_13725);
nand UO_0 (O_0,N_17977,N_16110);
xor UO_1 (O_1,N_18993,N_16208);
and UO_2 (O_2,N_18347,N_18917);
nor UO_3 (O_3,N_19230,N_19374);
xnor UO_4 (O_4,N_19639,N_17703);
nand UO_5 (O_5,N_16486,N_18493);
or UO_6 (O_6,N_16659,N_19547);
nand UO_7 (O_7,N_18742,N_17646);
or UO_8 (O_8,N_18218,N_16268);
and UO_9 (O_9,N_19443,N_16962);
and UO_10 (O_10,N_16970,N_19316);
xnor UO_11 (O_11,N_19127,N_18362);
and UO_12 (O_12,N_17267,N_19404);
or UO_13 (O_13,N_18422,N_16055);
nand UO_14 (O_14,N_16401,N_17483);
xnor UO_15 (O_15,N_18022,N_18268);
or UO_16 (O_16,N_19099,N_19063);
nand UO_17 (O_17,N_19478,N_17757);
xor UO_18 (O_18,N_18160,N_18952);
nor UO_19 (O_19,N_16884,N_17366);
and UO_20 (O_20,N_17799,N_16163);
and UO_21 (O_21,N_19419,N_19197);
and UO_22 (O_22,N_18156,N_19831);
xor UO_23 (O_23,N_18924,N_18570);
and UO_24 (O_24,N_19482,N_18152);
and UO_25 (O_25,N_16390,N_17756);
nand UO_26 (O_26,N_16722,N_17443);
nand UO_27 (O_27,N_17017,N_19264);
nand UO_28 (O_28,N_19435,N_17473);
xnor UO_29 (O_29,N_16681,N_17255);
xor UO_30 (O_30,N_17834,N_19181);
and UO_31 (O_31,N_16651,N_19651);
nand UO_32 (O_32,N_19778,N_19371);
nand UO_33 (O_33,N_19534,N_17418);
nand UO_34 (O_34,N_17359,N_17328);
xnor UO_35 (O_35,N_19323,N_18516);
or UO_36 (O_36,N_17556,N_17074);
xor UO_37 (O_37,N_17452,N_19471);
or UO_38 (O_38,N_19647,N_19454);
nor UO_39 (O_39,N_16744,N_16222);
nand UO_40 (O_40,N_16778,N_19248);
and UO_41 (O_41,N_16426,N_19751);
and UO_42 (O_42,N_16934,N_19580);
xor UO_43 (O_43,N_17915,N_19554);
nor UO_44 (O_44,N_16142,N_19598);
xnor UO_45 (O_45,N_18401,N_16555);
nor UO_46 (O_46,N_19839,N_18800);
or UO_47 (O_47,N_19406,N_18717);
and UO_48 (O_48,N_17315,N_18146);
and UO_49 (O_49,N_17490,N_19948);
and UO_50 (O_50,N_18994,N_17529);
nor UO_51 (O_51,N_18096,N_16481);
xnor UO_52 (O_52,N_18874,N_19335);
and UO_53 (O_53,N_19157,N_16973);
nand UO_54 (O_54,N_19207,N_19000);
and UO_55 (O_55,N_17187,N_19758);
and UO_56 (O_56,N_17582,N_18382);
xor UO_57 (O_57,N_18468,N_17080);
and UO_58 (O_58,N_16507,N_16251);
nand UO_59 (O_59,N_18689,N_16636);
nor UO_60 (O_60,N_18655,N_16836);
xnor UO_61 (O_61,N_19211,N_16726);
nand UO_62 (O_62,N_17073,N_17912);
xor UO_63 (O_63,N_19975,N_19479);
or UO_64 (O_64,N_17895,N_17369);
nor UO_65 (O_65,N_17622,N_19887);
and UO_66 (O_66,N_17218,N_17934);
and UO_67 (O_67,N_19326,N_19518);
or UO_68 (O_68,N_18028,N_16427);
xor UO_69 (O_69,N_16605,N_18195);
and UO_70 (O_70,N_17543,N_16617);
nand UO_71 (O_71,N_17827,N_19017);
nor UO_72 (O_72,N_19811,N_19333);
nor UO_73 (O_73,N_18885,N_16322);
or UO_74 (O_74,N_16686,N_16933);
and UO_75 (O_75,N_17431,N_17486);
nor UO_76 (O_76,N_17678,N_19511);
nor UO_77 (O_77,N_16148,N_16914);
nand UO_78 (O_78,N_17435,N_16409);
and UO_79 (O_79,N_18436,N_18001);
nor UO_80 (O_80,N_16948,N_19638);
or UO_81 (O_81,N_19633,N_19744);
nand UO_82 (O_82,N_19086,N_19603);
nand UO_83 (O_83,N_18880,N_17110);
nor UO_84 (O_84,N_19210,N_19779);
xor UO_85 (O_85,N_18292,N_19311);
xor UO_86 (O_86,N_18899,N_16536);
nor UO_87 (O_87,N_16618,N_18479);
xor UO_88 (O_88,N_18421,N_18442);
nor UO_89 (O_89,N_19716,N_18872);
or UO_90 (O_90,N_16224,N_16628);
nor UO_91 (O_91,N_17152,N_16485);
nor UO_92 (O_92,N_16865,N_18098);
xnor UO_93 (O_93,N_16739,N_16186);
or UO_94 (O_94,N_19971,N_18371);
or UO_95 (O_95,N_19769,N_19919);
or UO_96 (O_96,N_19338,N_16429);
and UO_97 (O_97,N_19882,N_17013);
and UO_98 (O_98,N_16423,N_17956);
or UO_99 (O_99,N_18563,N_19420);
and UO_100 (O_100,N_18884,N_19946);
and UO_101 (O_101,N_16718,N_17441);
and UO_102 (O_102,N_16491,N_16683);
and UO_103 (O_103,N_17609,N_17989);
nand UO_104 (O_104,N_18741,N_16967);
xnor UO_105 (O_105,N_18558,N_19244);
xor UO_106 (O_106,N_18951,N_16078);
xor UO_107 (O_107,N_19134,N_16438);
nor UO_108 (O_108,N_19485,N_18728);
nand UO_109 (O_109,N_16408,N_19559);
xor UO_110 (O_110,N_19530,N_16368);
and UO_111 (O_111,N_18157,N_18178);
nor UO_112 (O_112,N_16277,N_18329);
nor UO_113 (O_113,N_18731,N_18345);
xor UO_114 (O_114,N_17580,N_19392);
nor UO_115 (O_115,N_17333,N_19569);
or UO_116 (O_116,N_18839,N_18982);
xor UO_117 (O_117,N_16985,N_19346);
nor UO_118 (O_118,N_18669,N_16587);
and UO_119 (O_119,N_17780,N_16315);
or UO_120 (O_120,N_18019,N_18848);
and UO_121 (O_121,N_18440,N_17843);
nor UO_122 (O_122,N_19465,N_16930);
xnor UO_123 (O_123,N_18696,N_17889);
nor UO_124 (O_124,N_17260,N_17925);
nand UO_125 (O_125,N_17548,N_19266);
and UO_126 (O_126,N_16370,N_16327);
xnor UO_127 (O_127,N_17997,N_17368);
xnor UO_128 (O_128,N_17511,N_17919);
and UO_129 (O_129,N_19848,N_19128);
and UO_130 (O_130,N_19049,N_17750);
nor UO_131 (O_131,N_17410,N_16477);
or UO_132 (O_132,N_17809,N_19468);
nand UO_133 (O_133,N_19423,N_19125);
xnor UO_134 (O_134,N_18437,N_19236);
nor UO_135 (O_135,N_16007,N_16273);
and UO_136 (O_136,N_18119,N_17286);
nor UO_137 (O_137,N_19683,N_18139);
and UO_138 (O_138,N_19376,N_18455);
and UO_139 (O_139,N_19330,N_16174);
xnor UO_140 (O_140,N_17037,N_16512);
nor UO_141 (O_141,N_16310,N_16927);
or UO_142 (O_142,N_19452,N_16118);
nand UO_143 (O_143,N_18398,N_18108);
nor UO_144 (O_144,N_19444,N_18283);
nand UO_145 (O_145,N_17371,N_18518);
xnor UO_146 (O_146,N_17349,N_17201);
nor UO_147 (O_147,N_18317,N_18460);
xnor UO_148 (O_148,N_18510,N_16124);
and UO_149 (O_149,N_19618,N_17726);
xnor UO_150 (O_150,N_17310,N_19274);
nand UO_151 (O_151,N_18652,N_17545);
xor UO_152 (O_152,N_18121,N_18344);
and UO_153 (O_153,N_16439,N_18122);
nand UO_154 (O_154,N_17098,N_17796);
or UO_155 (O_155,N_19901,N_17733);
or UO_156 (O_156,N_16283,N_19934);
nor UO_157 (O_157,N_16354,N_18990);
nor UO_158 (O_158,N_19498,N_18340);
and UO_159 (O_159,N_19621,N_18410);
nand UO_160 (O_160,N_19077,N_18960);
nand UO_161 (O_161,N_16036,N_16122);
and UO_162 (O_162,N_19808,N_17920);
or UO_163 (O_163,N_19868,N_18496);
xor UO_164 (O_164,N_19148,N_16334);
or UO_165 (O_165,N_16777,N_16538);
and UO_166 (O_166,N_18045,N_18651);
nand UO_167 (O_167,N_16756,N_18415);
and UO_168 (O_168,N_17148,N_16372);
nand UO_169 (O_169,N_18972,N_17983);
and UO_170 (O_170,N_18454,N_16420);
xnor UO_171 (O_171,N_17227,N_16434);
nor UO_172 (O_172,N_19929,N_18445);
or UO_173 (O_173,N_19825,N_18576);
nand UO_174 (O_174,N_16242,N_18920);
nand UO_175 (O_175,N_19881,N_16475);
nand UO_176 (O_176,N_18908,N_18766);
or UO_177 (O_177,N_18200,N_17439);
nor UO_178 (O_178,N_16500,N_18759);
or UO_179 (O_179,N_19456,N_16798);
nand UO_180 (O_180,N_17065,N_16254);
or UO_181 (O_181,N_18368,N_17601);
nand UO_182 (O_182,N_19736,N_17623);
xor UO_183 (O_183,N_17472,N_16623);
and UO_184 (O_184,N_19555,N_16936);
nand UO_185 (O_185,N_17096,N_16905);
and UO_186 (O_186,N_18678,N_19958);
nor UO_187 (O_187,N_19538,N_17566);
nor UO_188 (O_188,N_18303,N_19380);
or UO_189 (O_189,N_19467,N_19360);
xnor UO_190 (O_190,N_19166,N_19317);
and UO_191 (O_191,N_18099,N_17633);
xnor UO_192 (O_192,N_16346,N_19842);
nand UO_193 (O_193,N_16953,N_17021);
or UO_194 (O_194,N_16245,N_17588);
nand UO_195 (O_195,N_16518,N_17658);
or UO_196 (O_196,N_19009,N_18027);
or UO_197 (O_197,N_18458,N_16762);
nand UO_198 (O_198,N_19747,N_16307);
nor UO_199 (O_199,N_18177,N_16484);
and UO_200 (O_200,N_16127,N_19821);
nand UO_201 (O_201,N_17520,N_18086);
and UO_202 (O_202,N_19663,N_19358);
nor UO_203 (O_203,N_17466,N_16490);
xnor UO_204 (O_204,N_19413,N_16793);
xor UO_205 (O_205,N_18379,N_18720);
xnor UO_206 (O_206,N_19182,N_18589);
nand UO_207 (O_207,N_16604,N_19854);
nor UO_208 (O_208,N_18544,N_19593);
or UO_209 (O_209,N_19944,N_17667);
and UO_210 (O_210,N_18774,N_16529);
or UO_211 (O_211,N_18414,N_19059);
and UO_212 (O_212,N_19476,N_18280);
or UO_213 (O_213,N_16264,N_19287);
xnor UO_214 (O_214,N_19004,N_18430);
or UO_215 (O_215,N_19441,N_16897);
nand UO_216 (O_216,N_16214,N_18789);
nor UO_217 (O_217,N_17052,N_17685);
xnor UO_218 (O_218,N_19268,N_17729);
or UO_219 (O_219,N_19272,N_16923);
and UO_220 (O_220,N_19373,N_16995);
nor UO_221 (O_221,N_17420,N_16724);
nand UO_222 (O_222,N_16407,N_19728);
and UO_223 (O_223,N_18143,N_17892);
or UO_224 (O_224,N_16391,N_16029);
or UO_225 (O_225,N_16018,N_17654);
xor UO_226 (O_226,N_17957,N_17952);
nor UO_227 (O_227,N_18818,N_18792);
nor UO_228 (O_228,N_18873,N_18512);
and UO_229 (O_229,N_19251,N_16431);
xor UO_230 (O_230,N_17561,N_19002);
or UO_231 (O_231,N_17415,N_19090);
and UO_232 (O_232,N_18816,N_17116);
and UO_233 (O_233,N_18695,N_16414);
xor UO_234 (O_234,N_19167,N_18622);
xnor UO_235 (O_235,N_18024,N_18933);
xnor UO_236 (O_236,N_18444,N_17170);
nand UO_237 (O_237,N_19937,N_19710);
and UO_238 (O_238,N_19327,N_17665);
nand UO_239 (O_239,N_19344,N_17718);
nand UO_240 (O_240,N_18048,N_16976);
and UO_241 (O_241,N_16573,N_19885);
nand UO_242 (O_242,N_16599,N_17049);
and UO_243 (O_243,N_19616,N_17849);
or UO_244 (O_244,N_19656,N_17874);
nand UO_245 (O_245,N_16316,N_16991);
nand UO_246 (O_246,N_18074,N_16794);
or UO_247 (O_247,N_17280,N_18758);
nand UO_248 (O_248,N_19252,N_17253);
xor UO_249 (O_249,N_16693,N_19249);
xor UO_250 (O_250,N_19290,N_16012);
or UO_251 (O_251,N_19965,N_17205);
and UO_252 (O_252,N_18914,N_18120);
and UO_253 (O_253,N_18854,N_17981);
nor UO_254 (O_254,N_16709,N_19657);
and UO_255 (O_255,N_18066,N_16228);
xor UO_256 (O_256,N_16941,N_16688);
nor UO_257 (O_257,N_17176,N_18783);
xor UO_258 (O_258,N_19552,N_16041);
or UO_259 (O_259,N_19817,N_17374);
or UO_260 (O_260,N_18999,N_18756);
xor UO_261 (O_261,N_16524,N_16281);
xor UO_262 (O_262,N_16400,N_19109);
or UO_263 (O_263,N_16037,N_17532);
xor UO_264 (O_264,N_16916,N_17653);
and UO_265 (O_265,N_16206,N_17671);
or UO_266 (O_266,N_18539,N_19730);
xor UO_267 (O_267,N_19601,N_18897);
nand UO_268 (O_268,N_19038,N_16821);
nor UO_269 (O_269,N_16382,N_18072);
nor UO_270 (O_270,N_19301,N_16158);
or UO_271 (O_271,N_18697,N_19117);
and UO_272 (O_272,N_16788,N_19265);
nand UO_273 (O_273,N_16571,N_19959);
nor UO_274 (O_274,N_17399,N_18294);
or UO_275 (O_275,N_17759,N_19658);
or UO_276 (O_276,N_16954,N_16337);
nand UO_277 (O_277,N_18969,N_19499);
nor UO_278 (O_278,N_16637,N_17583);
or UO_279 (O_279,N_18588,N_19217);
xor UO_280 (O_280,N_19133,N_19674);
nor UO_281 (O_281,N_16893,N_18017);
nor UO_282 (O_282,N_18672,N_19357);
and UO_283 (O_283,N_18419,N_17035);
nand UO_284 (O_284,N_18757,N_16111);
nor UO_285 (O_285,N_19520,N_19802);
nor UO_286 (O_286,N_19258,N_17230);
nor UO_287 (O_287,N_16664,N_17605);
nor UO_288 (O_288,N_16544,N_18888);
and UO_289 (O_289,N_17632,N_16393);
nand UO_290 (O_290,N_17515,N_17692);
nor UO_291 (O_291,N_18977,N_17041);
xnor UO_292 (O_292,N_16625,N_19036);
and UO_293 (O_293,N_16170,N_19073);
xor UO_294 (O_294,N_18612,N_16318);
nand UO_295 (O_295,N_16763,N_19472);
nand UO_296 (O_296,N_17030,N_16033);
or UO_297 (O_297,N_18610,N_19438);
nor UO_298 (O_298,N_17656,N_16115);
nand UO_299 (O_299,N_19081,N_18314);
or UO_300 (O_300,N_19149,N_18232);
xor UO_301 (O_301,N_16630,N_19584);
or UO_302 (O_302,N_19798,N_18606);
nor UO_303 (O_303,N_18834,N_16417);
and UO_304 (O_304,N_16364,N_17456);
nor UO_305 (O_305,N_18094,N_18217);
and UO_306 (O_306,N_17612,N_19171);
or UO_307 (O_307,N_16644,N_16458);
or UO_308 (O_308,N_18926,N_18192);
nor UO_309 (O_309,N_17265,N_19537);
nand UO_310 (O_310,N_16638,N_18583);
and UO_311 (O_311,N_19761,N_16211);
and UO_312 (O_312,N_18786,N_18716);
or UO_313 (O_313,N_16737,N_18003);
nand UO_314 (O_314,N_16175,N_19544);
nand UO_315 (O_315,N_16422,N_19313);
and UO_316 (O_316,N_17271,N_16169);
nand UO_317 (O_317,N_18274,N_16061);
nor UO_318 (O_318,N_18286,N_17506);
xnor UO_319 (O_319,N_17360,N_17115);
nand UO_320 (O_320,N_16509,N_16881);
and UO_321 (O_321,N_17361,N_18657);
nor UO_322 (O_322,N_17629,N_19019);
or UO_323 (O_323,N_19421,N_18199);
and UO_324 (O_324,N_18773,N_16576);
or UO_325 (O_325,N_17059,N_19056);
xnor UO_326 (O_326,N_19714,N_17537);
nand UO_327 (O_327,N_16549,N_19451);
and UO_328 (O_328,N_16546,N_19399);
and UO_329 (O_329,N_19813,N_18748);
nand UO_330 (O_330,N_16972,N_19737);
nor UO_331 (O_331,N_16325,N_16561);
xor UO_332 (O_332,N_17329,N_19754);
xor UO_333 (O_333,N_19349,N_16149);
nand UO_334 (O_334,N_16702,N_18549);
nor UO_335 (O_335,N_18784,N_16750);
nand UO_336 (O_336,N_19042,N_17903);
xnor UO_337 (O_337,N_18273,N_17502);
xnor UO_338 (O_338,N_19806,N_19648);
nand UO_339 (O_339,N_16047,N_19995);
nand UO_340 (O_340,N_17001,N_19993);
or UO_341 (O_341,N_19936,N_16270);
and UO_342 (O_342,N_16855,N_16106);
and UO_343 (O_343,N_16234,N_19561);
nand UO_344 (O_344,N_16802,N_16690);
xnor UO_345 (O_345,N_18184,N_17158);
nor UO_346 (O_346,N_17248,N_16129);
or UO_347 (O_347,N_19093,N_16910);
nand UO_348 (O_348,N_16454,N_18405);
xor UO_349 (O_349,N_17365,N_19440);
xor UO_350 (O_350,N_16023,N_18018);
xnor UO_351 (O_351,N_17774,N_16049);
xnor UO_352 (O_352,N_18447,N_18233);
and UO_353 (O_353,N_18406,N_16667);
and UO_354 (O_354,N_19989,N_18466);
and UO_355 (O_355,N_16979,N_18416);
and UO_356 (O_356,N_16772,N_19354);
and UO_357 (O_357,N_17002,N_16648);
nand UO_358 (O_358,N_16974,N_18381);
nand UO_359 (O_359,N_18722,N_19632);
and UO_360 (O_360,N_16929,N_16097);
and UO_361 (O_361,N_18310,N_16043);
xor UO_362 (O_362,N_18660,N_16789);
and UO_363 (O_363,N_16731,N_17914);
and UO_364 (O_364,N_18395,N_19097);
and UO_365 (O_365,N_16021,N_18685);
nor UO_366 (O_366,N_17129,N_19701);
and UO_367 (O_367,N_19228,N_17928);
nor UO_368 (O_368,N_19673,N_17558);
nand UO_369 (O_369,N_17500,N_18937);
nand UO_370 (O_370,N_19840,N_16809);
and UO_371 (O_371,N_19720,N_17705);
and UO_372 (O_372,N_17967,N_17741);
nand UO_373 (O_373,N_17800,N_17801);
nor UO_374 (O_374,N_17747,N_19484);
xnor UO_375 (O_375,N_18278,N_18863);
nor UO_376 (O_376,N_16001,N_19863);
xnor UO_377 (O_377,N_18250,N_18646);
nand UO_378 (O_378,N_16958,N_17467);
nor UO_379 (O_379,N_19562,N_16306);
nor UO_380 (O_380,N_18076,N_18114);
xnor UO_381 (O_381,N_19583,N_16369);
nor UO_382 (O_382,N_17006,N_18112);
nor UO_383 (O_383,N_18733,N_19974);
xor UO_384 (O_384,N_19068,N_19961);
nor UO_385 (O_385,N_17215,N_16569);
and UO_386 (O_386,N_16497,N_17536);
xnor UO_387 (O_387,N_17303,N_19634);
and UO_388 (O_388,N_17586,N_18891);
or UO_389 (O_389,N_17807,N_17931);
nand UO_390 (O_390,N_16566,N_19542);
and UO_391 (O_391,N_17666,N_16460);
nand UO_392 (O_392,N_17727,N_19763);
xor UO_393 (O_393,N_17239,N_16463);
nor UO_394 (O_394,N_16700,N_16220);
or UO_395 (O_395,N_16394,N_19305);
xor UO_396 (O_396,N_19455,N_19669);
nor UO_397 (O_397,N_16918,N_16633);
or UO_398 (O_398,N_17269,N_18882);
xnor UO_399 (O_399,N_17236,N_19426);
nor UO_400 (O_400,N_18936,N_16679);
nand UO_401 (O_401,N_19949,N_19764);
nor UO_402 (O_402,N_18149,N_16155);
nor UO_403 (O_403,N_16996,N_18843);
nand UO_404 (O_404,N_17820,N_18257);
xor UO_405 (O_405,N_19293,N_16792);
nor UO_406 (O_406,N_18536,N_16296);
nand UO_407 (O_407,N_18423,N_18615);
xor UO_408 (O_408,N_16374,N_16217);
or UO_409 (O_409,N_19853,N_17651);
nand UO_410 (O_410,N_17738,N_17854);
nand UO_411 (O_411,N_18145,N_18862);
nand UO_412 (O_412,N_17694,N_16988);
or UO_413 (O_413,N_19070,N_18433);
nor UO_414 (O_414,N_19113,N_17033);
xor UO_415 (O_415,N_16537,N_19759);
and UO_416 (O_416,N_19895,N_19486);
nor UO_417 (O_417,N_18743,N_16366);
or UO_418 (O_418,N_16917,N_16532);
xor UO_419 (O_419,N_19640,N_17770);
xor UO_420 (O_420,N_19935,N_18580);
nor UO_421 (O_421,N_16017,N_19026);
xor UO_422 (O_422,N_19890,N_19024);
and UO_423 (O_423,N_17714,N_17542);
and UO_424 (O_424,N_17089,N_19889);
and UO_425 (O_425,N_16938,N_19628);
xnor UO_426 (O_426,N_17314,N_17425);
nand UO_427 (O_427,N_18461,N_17283);
xnor UO_428 (O_428,N_18568,N_18954);
nor UO_429 (O_429,N_18054,N_16919);
nor UO_430 (O_430,N_19461,N_17963);
and UO_431 (O_431,N_18590,N_17434);
xnor UO_432 (O_432,N_18047,N_18738);
xor UO_433 (O_433,N_17828,N_16410);
nor UO_434 (O_434,N_19080,N_19790);
and UO_435 (O_435,N_19370,N_16707);
nor UO_436 (O_436,N_16942,N_16889);
xnor UO_437 (O_437,N_18829,N_18690);
nor UO_438 (O_438,N_17897,N_18380);
nand UO_439 (O_439,N_18103,N_18367);
nand UO_440 (O_440,N_16692,N_16553);
xor UO_441 (O_441,N_19163,N_16492);
xnor UO_442 (O_442,N_17861,N_18796);
nor UO_443 (O_443,N_18713,N_16223);
or UO_444 (O_444,N_17492,N_19200);
or UO_445 (O_445,N_17647,N_17784);
or UO_446 (O_446,N_17400,N_18605);
nand UO_447 (O_447,N_19220,N_16098);
xor UO_448 (O_448,N_17906,N_18886);
or UO_449 (O_449,N_16353,N_18025);
nor UO_450 (O_450,N_17890,N_17829);
and UO_451 (O_451,N_18744,N_19925);
xnor UO_452 (O_452,N_18730,N_19263);
or UO_453 (O_453,N_19767,N_16137);
or UO_454 (O_454,N_17185,N_19835);
and UO_455 (O_455,N_19687,N_19585);
nand UO_456 (O_456,N_16768,N_17916);
xor UO_457 (O_457,N_18674,N_19702);
nor UO_458 (O_458,N_18039,N_17385);
or UO_459 (O_459,N_18671,N_16854);
nor UO_460 (O_460,N_18942,N_18219);
or UO_461 (O_461,N_16769,N_16805);
nand UO_462 (O_462,N_16025,N_18353);
nand UO_463 (O_463,N_17512,N_19660);
nor UO_464 (O_464,N_19749,N_17938);
nor UO_465 (O_465,N_18375,N_19191);
nor UO_466 (O_466,N_19165,N_17358);
xor UO_467 (O_467,N_16237,N_19428);
or UO_468 (O_468,N_16808,N_17064);
and UO_469 (O_469,N_19797,N_16708);
xnor UO_470 (O_470,N_17830,N_19847);
xnor UO_471 (O_471,N_18469,N_19218);
nor UO_472 (O_472,N_19084,N_18515);
and UO_473 (O_473,N_17857,N_19654);
xnor UO_474 (O_474,N_16581,N_19150);
xor UO_475 (O_475,N_17879,N_18623);
xnor UO_476 (O_476,N_19475,N_19696);
nor UO_477 (O_477,N_16540,N_16986);
and UO_478 (O_478,N_19688,N_18667);
nand UO_479 (O_479,N_18182,N_18239);
and UO_480 (O_480,N_17522,N_19625);
or UO_481 (O_481,N_18855,N_18448);
and UO_482 (O_482,N_17554,N_16776);
nand UO_483 (O_483,N_18501,N_16767);
xnor UO_484 (O_484,N_18038,N_18259);
xor UO_485 (O_485,N_17572,N_19368);
xor UO_486 (O_486,N_17216,N_16870);
and UO_487 (O_487,N_18833,N_19159);
or UO_488 (O_488,N_16773,N_18255);
nor UO_489 (O_489,N_19908,N_17155);
or UO_490 (O_490,N_18916,N_18204);
or UO_491 (O_491,N_17390,N_19902);
nand UO_492 (O_492,N_17308,N_17824);
nand UO_493 (O_493,N_17372,N_19886);
xor UO_494 (O_494,N_18905,N_16344);
nand UO_495 (O_495,N_17050,N_18385);
nand UO_496 (O_496,N_17894,N_19715);
nand UO_497 (O_497,N_19557,N_18567);
or UO_498 (O_498,N_18209,N_18289);
or UO_499 (O_499,N_17232,N_17144);
xnor UO_500 (O_500,N_17575,N_19051);
nor UO_501 (O_501,N_19108,N_19904);
xor UO_502 (O_502,N_16363,N_18413);
nor UO_503 (O_503,N_16323,N_17146);
xnor UO_504 (O_504,N_17427,N_16760);
nor UO_505 (O_505,N_16874,N_16719);
xnor UO_506 (O_506,N_17223,N_19259);
nor UO_507 (O_507,N_16554,N_17433);
nand UO_508 (O_508,N_19067,N_19874);
or UO_509 (O_509,N_18797,N_16665);
and UO_510 (O_510,N_19234,N_17783);
nand UO_511 (O_511,N_16030,N_18011);
or UO_512 (O_512,N_19748,N_18231);
xor UO_513 (O_513,N_16607,N_19830);
nor UO_514 (O_514,N_18585,N_16657);
and UO_515 (O_515,N_17421,N_16287);
xnor UO_516 (O_516,N_16074,N_17095);
and UO_517 (O_517,N_16673,N_18935);
and UO_518 (O_518,N_17825,N_19962);
and UO_519 (O_519,N_16123,N_18223);
nor UO_520 (O_520,N_17362,N_19463);
nor UO_521 (O_521,N_18923,N_19943);
or UO_522 (O_522,N_16162,N_18547);
xor UO_523 (O_523,N_16894,N_16472);
and UO_524 (O_524,N_16164,N_19493);
and UO_525 (O_525,N_17102,N_17258);
xnor UO_526 (O_526,N_19300,N_17295);
nor UO_527 (O_527,N_17610,N_19334);
nor UO_528 (O_528,N_17765,N_17881);
nand UO_529 (O_529,N_19665,N_18625);
nor UO_530 (O_530,N_16255,N_16856);
nand UO_531 (O_531,N_17724,N_18193);
and UO_532 (O_532,N_16866,N_19771);
xor UO_533 (O_533,N_16184,N_18021);
or UO_534 (O_534,N_18694,N_17626);
nand UO_535 (O_535,N_18307,N_18364);
nand UO_536 (O_536,N_19981,N_19996);
nand UO_537 (O_537,N_17876,N_19222);
or UO_538 (O_538,N_16112,N_17010);
xor UO_539 (O_539,N_17699,N_17868);
nand UO_540 (O_540,N_19775,N_19470);
or UO_541 (O_541,N_19152,N_19030);
or UO_542 (O_542,N_18427,N_19563);
and UO_543 (O_543,N_18117,N_18485);
nor UO_544 (O_544,N_19415,N_19578);
nor UO_545 (O_545,N_16799,N_17590);
nand UO_546 (O_546,N_19143,N_16761);
xnor UO_547 (O_547,N_19203,N_16671);
xnor UO_548 (O_548,N_19653,N_17547);
nor UO_549 (O_549,N_18983,N_19064);
and UO_550 (O_550,N_17287,N_16820);
nor UO_551 (O_551,N_17761,N_17028);
or UO_552 (O_552,N_17551,N_18527);
nand UO_553 (O_553,N_17292,N_19102);
xnor UO_554 (O_554,N_16662,N_17736);
xnor UO_555 (O_555,N_18502,N_16196);
nand UO_556 (O_556,N_16591,N_16766);
xor UO_557 (O_557,N_17014,N_19667);
or UO_558 (O_558,N_19364,N_16333);
or UO_559 (O_559,N_17811,N_17092);
or UO_560 (O_560,N_16733,N_19697);
or UO_561 (O_561,N_19214,N_19689);
nand UO_562 (O_562,N_19564,N_19926);
nor UO_563 (O_563,N_19433,N_17126);
xor UO_564 (O_564,N_19187,N_18554);
or UO_565 (O_565,N_16785,N_17711);
xnor UO_566 (O_566,N_16295,N_17901);
nand UO_567 (O_567,N_18906,N_16499);
and UO_568 (O_568,N_19286,N_19940);
xor UO_569 (O_569,N_16703,N_18878);
xnor UO_570 (O_570,N_18276,N_16040);
or UO_571 (O_571,N_18754,N_16660);
or UO_572 (O_572,N_16822,N_17053);
xnor UO_573 (O_573,N_18127,N_16067);
nor UO_574 (O_574,N_19285,N_18343);
or UO_575 (O_575,N_19124,N_16867);
nand UO_576 (O_576,N_16015,N_18249);
nand UO_577 (O_577,N_19548,N_18109);
nand UO_578 (O_578,N_19977,N_17513);
nor UO_579 (O_579,N_19492,N_16404);
nor UO_580 (O_580,N_19599,N_17165);
and UO_581 (O_581,N_19731,N_18537);
and UO_582 (O_582,N_19308,N_19545);
nor UO_583 (O_583,N_17213,N_17987);
and UO_584 (O_584,N_18335,N_19328);
nand UO_585 (O_585,N_19727,N_16356);
or UO_586 (O_586,N_18850,N_19637);
or UO_587 (O_587,N_17198,N_17514);
and UO_588 (O_588,N_18523,N_18531);
and UO_589 (O_589,N_18070,N_17458);
xnor UO_590 (O_590,N_16610,N_19606);
nor UO_591 (O_591,N_19532,N_17079);
nor UO_592 (O_592,N_17636,N_19092);
or UO_593 (O_593,N_16852,N_18677);
nand UO_594 (O_594,N_16505,N_19850);
nor UO_595 (O_595,N_16728,N_16982);
xor UO_596 (O_596,N_18135,N_18302);
xnor UO_597 (O_597,N_17238,N_19312);
nor UO_598 (O_598,N_18319,N_16863);
or UO_599 (O_599,N_18726,N_19614);
or UO_600 (O_600,N_17051,N_16412);
nand UO_601 (O_601,N_18893,N_16157);
and UO_602 (O_602,N_17955,N_19867);
and UO_603 (O_603,N_16669,N_19690);
or UO_604 (O_604,N_18814,N_18288);
and UO_605 (O_605,N_18456,N_16717);
nand UO_606 (O_606,N_17744,N_17555);
nand UO_607 (O_607,N_17336,N_19039);
xnor UO_608 (O_608,N_17816,N_19597);
and UO_609 (O_609,N_17091,N_19533);
or UO_610 (O_610,N_19910,N_16311);
and UO_611 (O_611,N_17099,N_17237);
nor UO_612 (O_612,N_18418,N_19613);
nand UO_613 (O_613,N_16746,N_16790);
nand UO_614 (O_614,N_16453,N_19031);
and UO_615 (O_615,N_18712,N_17019);
nor UO_616 (O_616,N_16583,N_17494);
xnor UO_617 (O_617,N_17855,N_16457);
or UO_618 (O_618,N_18277,N_17182);
nor UO_619 (O_619,N_19581,N_18487);
nor UO_620 (O_620,N_18929,N_16138);
nand UO_621 (O_621,N_18470,N_17300);
or UO_622 (O_622,N_18533,N_16649);
xnor UO_623 (O_623,N_18497,N_17261);
nand UO_624 (O_624,N_17405,N_18804);
or UO_625 (O_625,N_19595,N_18927);
nand UO_626 (O_626,N_18597,N_17081);
xor UO_627 (O_627,N_17573,N_18737);
nand UO_628 (O_628,N_17918,N_16466);
nor UO_629 (O_629,N_16229,N_19131);
nand UO_630 (O_630,N_17553,N_16993);
nand UO_631 (O_631,N_16935,N_19786);
nand UO_632 (O_632,N_18543,N_16488);
or UO_633 (O_633,N_17011,N_18042);
xnor UO_634 (O_634,N_19695,N_17639);
or UO_635 (O_635,N_19104,N_19057);
and UO_636 (O_636,N_16612,N_16629);
or UO_637 (O_637,N_18002,N_19643);
nand UO_638 (O_638,N_19396,N_16876);
or UO_639 (O_639,N_16031,N_19713);
nand UO_640 (O_640,N_17994,N_18500);
nand UO_641 (O_641,N_18187,N_16687);
nor UO_642 (O_642,N_17364,N_17787);
or UO_643 (O_643,N_16543,N_17954);
or UO_644 (O_644,N_17461,N_16194);
nand UO_645 (O_645,N_19956,N_16847);
nand UO_646 (O_646,N_17873,N_17523);
or UO_647 (O_647,N_17839,N_16068);
and UO_648 (O_648,N_16946,N_19350);
xnor UO_649 (O_649,N_16959,N_17686);
or UO_650 (O_650,N_19592,N_17577);
nand UO_651 (O_651,N_17311,N_17103);
or UO_652 (O_652,N_17319,N_16470);
or UO_653 (O_653,N_19060,N_16464);
or UO_654 (O_654,N_17428,N_17980);
nand UO_655 (O_655,N_19400,N_16961);
xor UO_656 (O_656,N_19698,N_16205);
nand UO_657 (O_657,N_17939,N_18740);
and UO_658 (O_658,N_19602,N_17484);
or UO_659 (O_659,N_18552,N_17161);
and UO_660 (O_660,N_17025,N_19137);
nand UO_661 (O_661,N_16525,N_18691);
nor UO_662 (O_662,N_17644,N_17713);
nor UO_663 (O_663,N_19670,N_18428);
or UO_664 (O_664,N_18093,N_17382);
xnor UO_665 (O_665,N_18185,N_18535);
xor UO_666 (O_666,N_16203,N_18264);
and UO_667 (O_667,N_19983,N_17533);
nor UO_668 (O_668,N_16489,N_19815);
xnor UO_669 (O_669,N_18441,N_18858);
or UO_670 (O_670,N_19671,N_19164);
and UO_671 (O_671,N_18647,N_17259);
or UO_672 (O_672,N_18150,N_19094);
xnor UO_673 (O_673,N_17250,N_19620);
nand UO_674 (O_674,N_18180,N_17550);
or UO_675 (O_675,N_17085,N_18659);
nand UO_676 (O_676,N_19504,N_19072);
and UO_677 (O_677,N_19495,N_18306);
or UO_678 (O_678,N_16631,N_16070);
and UO_679 (O_679,N_16308,N_16782);
xnor UO_680 (O_680,N_18102,N_18198);
xor UO_681 (O_681,N_17072,N_17312);
nand UO_682 (O_682,N_18564,N_19947);
xnor UO_683 (O_683,N_19646,N_18938);
or UO_684 (O_684,N_19836,N_16928);
and UO_685 (O_685,N_19750,N_17923);
xor UO_686 (O_686,N_17114,N_19588);
nor UO_687 (O_687,N_17352,N_19635);
xor UO_688 (O_688,N_16380,N_19047);
nor UO_689 (O_689,N_17598,N_19278);
and UO_690 (O_690,N_18097,N_18519);
and UO_691 (O_691,N_17326,N_19384);
or UO_692 (O_692,N_19352,N_17683);
or UO_693 (O_693,N_19088,N_18890);
nor UO_694 (O_694,N_17403,N_16578);
xnor UO_695 (O_695,N_19844,N_18113);
and UO_696 (O_696,N_19123,N_19630);
and UO_697 (O_697,N_16841,N_19083);
or UO_698 (O_698,N_19389,N_16116);
xor UO_699 (O_699,N_16132,N_17438);
nor UO_700 (O_700,N_17357,N_18007);
nand UO_701 (O_701,N_18238,N_16300);
or UO_702 (O_702,N_17027,N_17663);
nand UO_703 (O_703,N_16901,N_18069);
xnor UO_704 (O_704,N_18036,N_16216);
or UO_705 (O_705,N_18688,N_17781);
and UO_706 (O_706,N_17937,N_17730);
and UO_707 (O_707,N_18988,N_18296);
nor UO_708 (O_708,N_16172,N_16720);
xor UO_709 (O_709,N_19718,N_18168);
nor UO_710 (O_710,N_18877,N_17976);
xor UO_711 (O_711,N_17207,N_18144);
and UO_712 (O_712,N_19679,N_16383);
and UO_713 (O_713,N_16840,N_19500);
or UO_714 (O_714,N_17453,N_16080);
nor UO_715 (O_715,N_16447,N_18321);
nand UO_716 (O_716,N_19196,N_18365);
or UO_717 (O_717,N_19921,N_19006);
nand UO_718 (O_718,N_16005,N_18251);
xor UO_719 (O_719,N_18524,N_17974);
and UO_720 (O_720,N_17270,N_16028);
and UO_721 (O_721,N_19923,N_17469);
nand UO_722 (O_722,N_17125,N_18265);
or UO_723 (O_723,N_16526,N_16279);
and UO_724 (O_724,N_16695,N_16461);
nor UO_725 (O_725,N_17631,N_18719);
or UO_726 (O_726,N_17022,N_19899);
or UO_727 (O_727,N_19240,N_16360);
nor UO_728 (O_728,N_18836,N_18492);
and UO_729 (O_729,N_18864,N_19642);
nor UO_730 (O_730,N_16878,N_16002);
nor UO_731 (O_731,N_16879,N_19551);
and UO_732 (O_732,N_19875,N_16541);
xnor UO_733 (O_733,N_16083,N_18525);
nor UO_734 (O_734,N_16386,N_18844);
nand UO_735 (O_735,N_18711,N_18148);
nand UO_736 (O_736,N_18867,N_16054);
nor UO_737 (O_737,N_17249,N_18782);
xnor UO_738 (O_738,N_19048,N_16011);
and UO_739 (O_739,N_19035,N_18142);
nor UO_740 (O_740,N_16069,N_19314);
nand UO_741 (O_741,N_19512,N_18981);
nand UO_742 (O_742,N_16140,N_17875);
nor UO_743 (O_743,N_18755,N_17169);
nand UO_744 (O_744,N_19777,N_16506);
and UO_745 (O_745,N_18932,N_18092);
xnor UO_746 (O_746,N_17641,N_17965);
and UO_747 (O_747,N_16655,N_16355);
and UO_748 (O_748,N_18556,N_18111);
and UO_749 (O_749,N_16796,N_16684);
and UO_750 (O_750,N_16248,N_18845);
and UO_751 (O_751,N_16063,N_16085);
nand UO_752 (O_752,N_17754,N_17669);
and UO_753 (O_753,N_16749,N_19973);
xor UO_754 (O_754,N_18817,N_18167);
nor UO_755 (O_755,N_17327,N_17627);
nand UO_756 (O_756,N_16861,N_16415);
nand UO_757 (O_757,N_16094,N_17131);
nor UO_758 (O_758,N_17739,N_17409);
xnor UO_759 (O_759,N_19391,N_17755);
or UO_760 (O_760,N_17764,N_17785);
xnor UO_761 (O_761,N_18263,N_17379);
and UO_762 (O_762,N_19877,N_19623);
nor UO_763 (O_763,N_17173,N_18129);
nor UO_764 (O_764,N_17521,N_16797);
nand UO_765 (O_765,N_17417,N_19820);
or UO_766 (O_766,N_19735,N_18012);
nand UO_767 (O_767,N_16039,N_18034);
nand UO_768 (O_768,N_17437,N_17167);
or UO_769 (O_769,N_17935,N_16902);
and UO_770 (O_770,N_19525,N_17214);
and UO_771 (O_771,N_18170,N_19310);
nand UO_772 (O_772,N_18057,N_19202);
xnor UO_773 (O_773,N_19477,N_19819);
and UO_774 (O_774,N_17959,N_18465);
nor UO_775 (O_775,N_16341,N_18621);
nor UO_776 (O_776,N_18224,N_17619);
nor UO_777 (O_777,N_18875,N_18643);
or UO_778 (O_778,N_19276,N_16285);
or UO_779 (O_779,N_19565,N_16831);
nand UO_780 (O_780,N_17406,N_19785);
xnor UO_781 (O_781,N_18339,N_17530);
nand UO_782 (O_782,N_18407,N_18734);
nand UO_783 (O_783,N_19412,N_17680);
or UO_784 (O_784,N_17040,N_18928);
nor UO_785 (O_785,N_17481,N_16759);
or UO_786 (O_786,N_17317,N_19076);
xor UO_787 (O_787,N_18010,N_18587);
and UO_788 (O_788,N_18649,N_18172);
nor UO_789 (O_789,N_18222,N_16912);
and UO_790 (O_790,N_18186,N_19353);
nor UO_791 (O_791,N_17111,N_18281);
nand UO_792 (O_792,N_16253,N_19238);
xnor UO_793 (O_793,N_16579,N_18979);
nand UO_794 (O_794,N_17637,N_18808);
xnor UO_795 (O_795,N_17604,N_16324);
xor UO_796 (O_796,N_16560,N_18628);
nor UO_797 (O_797,N_17332,N_16551);
and UO_798 (O_798,N_17226,N_17606);
xor UO_799 (O_799,N_16890,N_16613);
or UO_800 (O_800,N_19998,N_16738);
nand UO_801 (O_801,N_17274,N_19717);
nand UO_802 (O_802,N_17772,N_16089);
xor UO_803 (O_803,N_16994,N_19458);
xor UO_804 (O_804,N_17109,N_17008);
nor UO_805 (O_805,N_18334,N_16403);
nand UO_806 (O_806,N_18451,N_19507);
or UO_807 (O_807,N_16764,N_19876);
and UO_808 (O_808,N_18600,N_19664);
xor UO_809 (O_809,N_19058,N_18154);
and UO_810 (O_810,N_17324,N_19022);
and UO_811 (O_811,N_19362,N_16634);
and UO_812 (O_812,N_19257,N_16071);
and UO_813 (O_813,N_19608,N_17948);
nor UO_814 (O_814,N_18573,N_16900);
and UO_815 (O_815,N_19509,N_16392);
nor UO_816 (O_816,N_19743,N_19755);
nor UO_817 (O_817,N_17426,N_17331);
or UO_818 (O_818,N_19082,N_18384);
xor UO_819 (O_819,N_17408,N_17068);
nand UO_820 (O_820,N_17748,N_18707);
nand UO_821 (O_821,N_19462,N_18665);
or UO_822 (O_822,N_19267,N_19385);
xor UO_823 (O_823,N_17090,N_16236);
and UO_824 (O_824,N_19957,N_19237);
and UO_825 (O_825,N_18235,N_16685);
nand UO_826 (O_826,N_18077,N_18698);
or UO_827 (O_827,N_17595,N_18494);
xnor UO_828 (O_828,N_17517,N_16385);
and UO_829 (O_829,N_18909,N_17302);
nand UO_830 (O_830,N_18046,N_18090);
or UO_831 (O_831,N_17196,N_18000);
or UO_832 (O_832,N_17313,N_16042);
nand UO_833 (O_833,N_18328,N_19115);
xor UO_834 (O_834,N_19550,N_19153);
or UO_835 (O_835,N_19883,N_16860);
or UO_836 (O_836,N_18110,N_18491);
and UO_837 (O_837,N_19273,N_17156);
and UO_838 (O_838,N_17337,N_18629);
or UO_839 (O_839,N_19221,N_18747);
and UO_840 (O_840,N_18593,N_16668);
nand UO_841 (O_841,N_19930,N_17943);
nand UO_842 (O_842,N_18495,N_18624);
nand UO_843 (O_843,N_16812,N_18913);
nand UO_844 (O_844,N_19801,N_18349);
xor UO_845 (O_845,N_19052,N_18220);
and UO_846 (O_846,N_18577,N_16304);
or UO_847 (O_847,N_19911,N_19138);
xnor UO_848 (O_848,N_17546,N_16871);
nand UO_849 (O_849,N_18673,N_16260);
or UO_850 (O_850,N_17347,N_19295);
xor UO_851 (O_851,N_16173,N_16003);
and UO_852 (O_852,N_17584,N_17034);
nor UO_853 (O_853,N_16807,N_18974);
and UO_854 (O_854,N_16301,N_16202);
nand UO_855 (O_855,N_19007,N_17621);
xor UO_856 (O_856,N_16419,N_17272);
or UO_857 (O_857,N_17932,N_16949);
xor UO_858 (O_858,N_17964,N_17592);
nand UO_859 (O_859,N_17200,N_18687);
nor UO_860 (O_860,N_17802,N_18599);
or UO_861 (O_861,N_17465,N_18530);
xnor UO_862 (O_862,N_18091,N_18115);
and UO_863 (O_863,N_17661,N_17866);
nor UO_864 (O_864,N_17039,N_17460);
xor UO_865 (O_865,N_18846,N_16416);
xor UO_866 (O_866,N_17301,N_16666);
nor UO_867 (O_867,N_17618,N_19909);
nor UO_868 (O_868,N_19106,N_16875);
and UO_869 (O_869,N_19922,N_18258);
xnor UO_870 (O_870,N_17565,N_19074);
or UO_871 (O_871,N_16256,N_17518);
and UO_872 (O_872,N_19609,N_18134);
nand UO_873 (O_873,N_17803,N_17607);
xor UO_874 (O_874,N_18798,N_18883);
and UO_875 (O_875,N_19279,N_16534);
and UO_876 (O_876,N_17808,N_19570);
nand UO_877 (O_877,N_17602,N_19756);
and UO_878 (O_878,N_17717,N_18498);
xnor UO_879 (O_879,N_19587,N_19960);
nand UO_880 (O_880,N_18431,N_19624);
xnor UO_881 (O_881,N_18820,N_16450);
nor UO_882 (O_882,N_16735,N_16027);
nand UO_883 (O_883,N_16519,N_17070);
nand UO_884 (O_884,N_19768,N_16969);
xor UO_885 (O_885,N_17166,N_19447);
nand UO_886 (O_886,N_18813,N_16844);
nand UO_887 (O_887,N_18636,N_16858);
or UO_888 (O_888,N_16827,N_19087);
or UO_889 (O_889,N_16670,N_18333);
xor UO_890 (O_890,N_16517,N_18962);
nor UO_891 (O_891,N_19322,N_16804);
or UO_892 (O_892,N_17143,N_18842);
xnor UO_893 (O_893,N_19791,N_18291);
xnor UO_894 (O_894,N_16073,N_16082);
xor UO_895 (O_895,N_16181,N_19931);
or UO_896 (O_896,N_17288,N_17712);
and UO_897 (O_897,N_19254,N_18216);
xor UO_898 (O_898,N_19681,N_17579);
and UO_899 (O_899,N_17163,N_19540);
nor UO_900 (O_900,N_19568,N_19855);
nand UO_901 (O_901,N_17266,N_19990);
nand UO_902 (O_902,N_19866,N_16926);
nor UO_903 (O_903,N_17858,N_16743);
nor UO_904 (O_904,N_18100,N_18404);
nor UO_905 (O_905,N_16803,N_17505);
and UO_906 (O_906,N_17233,N_18718);
and UO_907 (O_907,N_17568,N_18082);
nor UO_908 (O_908,N_16786,N_16920);
nor UO_909 (O_909,N_16171,N_19436);
nand UO_910 (O_910,N_19536,N_17038);
nor UO_911 (O_911,N_19055,N_16734);
nand UO_912 (O_912,N_16757,N_19549);
and UO_913 (O_913,N_19069,N_16891);
or UO_914 (O_914,N_19037,N_19997);
nor UO_915 (O_915,N_19969,N_18489);
or UO_916 (O_916,N_17268,N_18138);
nor UO_917 (O_917,N_17128,N_19410);
nand UO_918 (O_918,N_17624,N_18912);
nor UO_919 (O_919,N_18206,N_18316);
and UO_920 (O_920,N_19980,N_17463);
or UO_921 (O_921,N_18008,N_16606);
nor UO_922 (O_922,N_17222,N_17544);
and UO_923 (O_923,N_19424,N_17284);
xor UO_924 (O_924,N_16515,N_18879);
and UO_925 (O_925,N_18627,N_16121);
nor UO_926 (O_926,N_18663,N_17078);
nand UO_927 (O_927,N_19920,N_16079);
or UO_928 (O_928,N_19849,N_17700);
xor UO_929 (O_929,N_19915,N_16187);
or UO_930 (O_930,N_18560,N_16653);
xor UO_931 (O_931,N_19315,N_17867);
nor UO_932 (O_932,N_18968,N_17510);
xnor UO_933 (O_933,N_17157,N_19986);
nand UO_934 (O_934,N_17171,N_16826);
and UO_935 (O_935,N_19071,N_17525);
and UO_936 (O_936,N_19116,N_18966);
and UO_937 (O_937,N_16406,N_16272);
nor UO_938 (O_938,N_16869,N_17650);
nand UO_939 (O_939,N_16833,N_17234);
or UO_940 (O_940,N_17350,N_17373);
and UO_941 (O_941,N_19757,N_17851);
and UO_942 (O_942,N_17067,N_17203);
nand UO_943 (O_943,N_17842,N_19363);
or UO_944 (O_944,N_17130,N_19025);
and UO_945 (O_945,N_18684,N_19193);
and UO_946 (O_946,N_18601,N_18188);
nor UO_947 (O_947,N_19034,N_19403);
nor UO_948 (O_948,N_17562,N_19898);
nor UO_949 (O_949,N_16977,N_17202);
nor UO_950 (O_950,N_19740,N_17732);
or UO_951 (O_951,N_16365,N_18870);
nor UO_952 (O_952,N_19079,N_16725);
xnor UO_953 (O_953,N_16008,N_19968);
nor UO_954 (O_954,N_19560,N_16159);
and UO_955 (O_955,N_17291,N_16195);
nor UO_956 (O_956,N_16645,N_19794);
or UO_957 (O_957,N_16964,N_19837);
xor UO_958 (O_958,N_19029,N_17767);
nand UO_959 (O_959,N_18559,N_16190);
nand UO_960 (O_960,N_17725,N_18984);
xnor UO_961 (O_961,N_19480,N_19226);
and UO_962 (O_962,N_19448,N_19824);
nand UO_963 (O_963,N_17384,N_16332);
or UO_964 (O_964,N_19297,N_16004);
or UO_965 (O_965,N_16226,N_16795);
nor UO_966 (O_966,N_16857,N_19397);
or UO_967 (O_967,N_17388,N_19589);
nand UO_968 (O_968,N_18898,N_18584);
xor UO_969 (O_969,N_19241,N_19140);
nor UO_970 (O_970,N_16883,N_19411);
xor UO_971 (O_971,N_18369,N_16824);
nor UO_972 (O_972,N_17933,N_16877);
and UO_973 (O_973,N_18400,N_19450);
xnor UO_974 (O_974,N_18534,N_16320);
and UO_975 (O_975,N_19573,N_17883);
and UO_976 (O_976,N_19043,N_18298);
and UO_977 (O_977,N_18023,N_18948);
and UO_978 (O_978,N_16741,N_16182);
and UO_979 (O_979,N_19188,N_18941);
nand UO_980 (O_980,N_17758,N_16705);
or UO_981 (O_981,N_17684,N_16204);
and UO_982 (O_982,N_16987,N_19590);
or UO_983 (O_983,N_16832,N_16432);
nor UO_984 (O_984,N_16661,N_18260);
nor UO_985 (O_985,N_17009,N_17191);
and UO_986 (O_986,N_18191,N_18793);
and UO_987 (O_987,N_18033,N_17751);
or UO_988 (O_988,N_18555,N_18040);
or UO_989 (O_989,N_17097,N_18607);
xnor UO_990 (O_990,N_19250,N_17869);
nand UO_991 (O_991,N_16405,N_16084);
xor UO_992 (O_992,N_18499,N_16539);
nor UO_993 (O_993,N_18208,N_19515);
or UO_994 (O_994,N_19114,N_19954);
nor UO_995 (O_995,N_18705,N_16595);
xor UO_996 (O_996,N_18822,N_19617);
and UO_997 (O_997,N_17018,N_17320);
nand UO_998 (O_998,N_16895,N_16014);
and UO_999 (O_999,N_19449,N_19827);
xnor UO_1000 (O_1000,N_17204,N_18272);
nor UO_1001 (O_1001,N_18080,N_19491);
nor UO_1002 (O_1002,N_18823,N_18958);
and UO_1003 (O_1003,N_19299,N_16952);
nor UO_1004 (O_1004,N_17762,N_18248);
nor UO_1005 (O_1005,N_19377,N_17262);
or UO_1006 (O_1006,N_17264,N_17742);
nor UO_1007 (O_1007,N_18881,N_17709);
xor UO_1008 (O_1008,N_16131,N_18571);
or UO_1009 (O_1009,N_17872,N_17930);
and UO_1010 (O_1010,N_16627,N_19126);
xnor UO_1011 (O_1011,N_16603,N_16710);
nand UO_1012 (O_1012,N_19607,N_18795);
and UO_1013 (O_1013,N_19232,N_18073);
nand UO_1014 (O_1014,N_19927,N_18124);
or UO_1015 (O_1015,N_19177,N_17206);
and UO_1016 (O_1016,N_17257,N_17478);
nand UO_1017 (O_1017,N_19970,N_16698);
nand UO_1018 (O_1018,N_19277,N_18778);
xnor UO_1019 (O_1019,N_16088,N_19804);
nand UO_1020 (O_1020,N_18921,N_16289);
xnor UO_1021 (O_1021,N_16915,N_18346);
xor UO_1022 (O_1022,N_17242,N_17710);
or UO_1023 (O_1023,N_16119,N_18639);
nor UO_1024 (O_1024,N_17477,N_17150);
xnor UO_1025 (O_1025,N_19343,N_19682);
and UO_1026 (O_1026,N_16528,N_16609);
or UO_1027 (O_1027,N_17723,N_18215);
nand UO_1028 (O_1028,N_17978,N_18162);
nand UO_1029 (O_1029,N_19355,N_18900);
xnor UO_1030 (O_1030,N_18569,N_19789);
or UO_1031 (O_1031,N_17988,N_19028);
or UO_1032 (O_1032,N_17355,N_17887);
and UO_1033 (O_1033,N_18267,N_17630);
or UO_1034 (O_1034,N_16828,N_18044);
and UO_1035 (O_1035,N_16247,N_19383);
and UO_1036 (O_1036,N_16911,N_18490);
nand UO_1037 (O_1037,N_16048,N_18126);
xnor UO_1038 (O_1038,N_16144,N_18383);
nor UO_1039 (O_1039,N_17042,N_19223);
nand UO_1040 (O_1040,N_18598,N_17354);
nor UO_1041 (O_1041,N_16034,N_17036);
or UO_1042 (O_1042,N_19553,N_16520);
xnor UO_1043 (O_1043,N_18477,N_19726);
xnor UO_1044 (O_1044,N_16819,N_18484);
nor UO_1045 (O_1045,N_19933,N_18965);
nor UO_1046 (O_1046,N_16153,N_17489);
nand UO_1047 (O_1047,N_19611,N_19430);
nand UO_1048 (O_1048,N_19008,N_17377);
nor UO_1049 (O_1049,N_18056,N_16455);
and UO_1050 (O_1050,N_19409,N_19641);
xnor UO_1051 (O_1051,N_18318,N_16035);
nor UO_1052 (O_1052,N_16150,N_18026);
nor UO_1053 (O_1053,N_17289,N_19179);
or UO_1054 (O_1054,N_17189,N_16680);
xnor UO_1055 (O_1055,N_18887,N_19490);
nand UO_1056 (O_1056,N_17596,N_19439);
or UO_1057 (O_1057,N_19422,N_16997);
or UO_1058 (O_1058,N_16087,N_19417);
nor UO_1059 (O_1059,N_18095,N_17782);
nand UO_1060 (O_1060,N_16238,N_17913);
nand UO_1061 (O_1061,N_18372,N_17127);
nor UO_1062 (O_1062,N_16747,N_19145);
xor UO_1063 (O_1063,N_19514,N_16752);
nor UO_1064 (O_1064,N_16943,N_16250);
nor UO_1065 (O_1065,N_16641,N_18290);
or UO_1066 (O_1066,N_19722,N_18031);
nand UO_1067 (O_1067,N_19100,N_17853);
nor UO_1068 (O_1068,N_19388,N_16899);
xor UO_1069 (O_1069,N_19275,N_17082);
nand UO_1070 (O_1070,N_18356,N_17471);
xor UO_1071 (O_1071,N_17845,N_18837);
or UO_1072 (O_1072,N_19018,N_19803);
and UO_1073 (O_1073,N_16387,N_19173);
or UO_1074 (O_1074,N_19280,N_19984);
nand UO_1075 (O_1075,N_18254,N_17459);
or UO_1076 (O_1076,N_18128,N_18866);
nor UO_1077 (O_1077,N_16299,N_19703);
nor UO_1078 (O_1078,N_17015,N_17275);
xor UO_1079 (O_1079,N_17407,N_18141);
nor UO_1080 (O_1080,N_19262,N_18775);
xor UO_1081 (O_1081,N_17031,N_18931);
or UO_1082 (O_1082,N_18325,N_17936);
xor UO_1083 (O_1083,N_16656,N_16176);
or UO_1084 (O_1084,N_18337,N_17674);
nor UO_1085 (O_1085,N_16376,N_16596);
or UO_1086 (O_1086,N_16151,N_19180);
or UO_1087 (O_1087,N_16358,N_18911);
or UO_1088 (O_1088,N_16261,N_19781);
or UO_1089 (O_1089,N_16714,N_16577);
xnor UO_1090 (O_1090,N_16559,N_18749);
nor UO_1091 (O_1091,N_16727,N_19320);
or UO_1092 (O_1092,N_19178,N_18550);
and UO_1093 (O_1093,N_18551,N_19046);
or UO_1094 (O_1094,N_19650,N_19707);
xor UO_1095 (O_1095,N_18043,N_16780);
and UO_1096 (O_1096,N_16501,N_18637);
or UO_1097 (O_1097,N_16288,N_17339);
or UO_1098 (O_1098,N_16924,N_17348);
and UO_1099 (O_1099,N_19382,N_18925);
and UO_1100 (O_1100,N_16221,N_16467);
and UO_1101 (O_1101,N_16388,N_18475);
nor UO_1102 (O_1102,N_16770,N_17084);
nor UO_1103 (O_1103,N_16677,N_16117);
and UO_1104 (O_1104,N_18805,N_17728);
and UO_1105 (O_1105,N_18953,N_19541);
or UO_1106 (O_1106,N_17707,N_17670);
nand UO_1107 (O_1107,N_17910,N_19395);
nand UO_1108 (O_1108,N_18631,N_17942);
and UO_1109 (O_1109,N_17975,N_18443);
and UO_1110 (O_1110,N_19020,N_16090);
or UO_1111 (O_1111,N_18940,N_18363);
xnor UO_1112 (O_1112,N_17541,N_17104);
or UO_1113 (O_1113,N_16135,N_17793);
nand UO_1114 (O_1114,N_19351,N_17318);
nor UO_1115 (O_1115,N_19506,N_18207);
or UO_1116 (O_1116,N_19833,N_17693);
xnor UO_1117 (O_1117,N_16514,N_17147);
xor UO_1118 (O_1118,N_19543,N_19023);
xor UO_1119 (O_1119,N_17507,N_19186);
xor UO_1120 (O_1120,N_19676,N_16567);
nand UO_1121 (O_1121,N_17946,N_19571);
or UO_1122 (O_1122,N_17133,N_17856);
xnor UO_1123 (O_1123,N_18075,N_18261);
and UO_1124 (O_1124,N_19011,N_19894);
and UO_1125 (O_1125,N_18323,N_19416);
nor UO_1126 (O_1126,N_19579,N_19119);
and UO_1127 (O_1127,N_16399,N_17482);
nand UO_1128 (O_1128,N_19787,N_17325);
or UO_1129 (O_1129,N_17297,N_18579);
xnor UO_1130 (O_1130,N_18950,N_19828);
and UO_1131 (O_1131,N_16160,N_18304);
nor UO_1132 (O_1132,N_18616,N_17643);
and UO_1133 (O_1133,N_16654,N_19414);
nand UO_1134 (O_1134,N_16535,N_18166);
nor UO_1135 (O_1135,N_17953,N_16053);
nor UO_1136 (O_1136,N_18201,N_17293);
and UO_1137 (O_1137,N_19845,N_19519);
nand UO_1138 (O_1138,N_16101,N_17991);
xnor UO_1139 (O_1139,N_19209,N_16314);
nand UO_1140 (O_1140,N_18163,N_19985);
xnor UO_1141 (O_1141,N_18970,N_16697);
or UO_1142 (O_1142,N_16593,N_16139);
nand UO_1143 (O_1143,N_16213,N_16179);
or UO_1144 (O_1144,N_18473,N_18654);
nor UO_1145 (O_1145,N_19800,N_19445);
nor UO_1146 (O_1146,N_18642,N_17720);
xor UO_1147 (O_1147,N_18322,N_16601);
and UO_1148 (O_1148,N_19098,N_17746);
and UO_1149 (O_1149,N_18706,N_16678);
or UO_1150 (O_1150,N_16589,N_17071);
and UO_1151 (O_1151,N_17792,N_18700);
nor UO_1152 (O_1152,N_16456,N_17278);
nor UO_1153 (O_1153,N_17900,N_18996);
or UO_1154 (O_1154,N_16436,N_19741);
xnor UO_1155 (O_1155,N_17491,N_19566);
xnor UO_1156 (O_1156,N_19225,N_16125);
nor UO_1157 (O_1157,N_16696,N_16830);
and UO_1158 (O_1158,N_18764,N_17649);
nand UO_1159 (O_1159,N_16062,N_19142);
nand UO_1160 (O_1160,N_17958,N_17119);
or UO_1161 (O_1161,N_18609,N_16806);
and UO_1162 (O_1162,N_16284,N_19870);
xnor UO_1163 (O_1163,N_17047,N_17380);
xor UO_1164 (O_1164,N_19497,N_19945);
and UO_1165 (O_1165,N_17316,N_16614);
or UO_1166 (O_1166,N_16189,N_18165);
and UO_1167 (O_1167,N_19891,N_18787);
or UO_1168 (O_1168,N_16413,N_18980);
and UO_1169 (O_1169,N_16508,N_17087);
or UO_1170 (O_1170,N_17123,N_18106);
nor UO_1171 (O_1171,N_19652,N_16582);
nor UO_1172 (O_1172,N_17689,N_17821);
xor UO_1173 (O_1173,N_19010,N_16845);
nor UO_1174 (O_1174,N_18645,N_18619);
or UO_1175 (O_1175,N_17281,N_16286);
xnor UO_1176 (O_1176,N_18425,N_17549);
or UO_1177 (O_1177,N_17679,N_16207);
and UO_1178 (O_1178,N_19302,N_17993);
nand UO_1179 (O_1179,N_19402,N_16791);
nor UO_1180 (O_1180,N_19605,N_16274);
and UO_1181 (O_1181,N_19873,N_16096);
xnor UO_1182 (O_1182,N_19631,N_19814);
and UO_1183 (O_1183,N_18392,N_16398);
nand UO_1184 (O_1184,N_18871,N_19600);
nor UO_1185 (O_1185,N_17599,N_17046);
or UO_1186 (O_1186,N_16944,N_18955);
nor UO_1187 (O_1187,N_16347,N_19528);
xor UO_1188 (O_1188,N_18378,N_18892);
and UO_1189 (O_1189,N_16058,N_16302);
nor UO_1190 (O_1190,N_16275,N_16736);
xnor UO_1191 (O_1191,N_17112,N_17831);
nand UO_1192 (O_1192,N_16842,N_19880);
nand UO_1193 (O_1193,N_19269,N_18373);
nand UO_1194 (O_1194,N_18930,N_18151);
and UO_1195 (O_1195,N_19672,N_16850);
xor UO_1196 (O_1196,N_16632,N_16829);
xnor UO_1197 (O_1197,N_18176,N_19649);
nor UO_1198 (O_1198,N_17924,N_18732);
xnor UO_1199 (O_1199,N_16584,N_16745);
xnor UO_1200 (O_1200,N_19752,N_17121);
and UO_1201 (O_1201,N_18729,N_19016);
xnor UO_1202 (O_1202,N_16955,N_18557);
xor UO_1203 (O_1203,N_16598,N_18553);
and UO_1204 (O_1204,N_16230,N_18449);
xnor UO_1205 (O_1205,N_17593,N_17862);
xor UO_1206 (O_1206,N_19526,N_17672);
and UO_1207 (O_1207,N_17395,N_18155);
nor UO_1208 (O_1208,N_19387,N_16572);
nand UO_1209 (O_1209,N_18826,N_19572);
xnor UO_1210 (O_1210,N_17891,N_18715);
nand UO_1211 (O_1211,N_19857,N_18675);
and UO_1212 (O_1212,N_16183,N_18803);
nand UO_1213 (O_1213,N_17229,N_17888);
or UO_1214 (O_1214,N_16292,N_16600);
nand UO_1215 (O_1215,N_16013,N_16921);
or UO_1216 (O_1216,N_16193,N_17118);
or UO_1217 (O_1217,N_19577,N_18902);
nor UO_1218 (O_1218,N_19916,N_17690);
and UO_1219 (O_1219,N_17835,N_18256);
nor UO_1220 (O_1220,N_17149,N_17905);
and UO_1221 (O_1221,N_17448,N_18446);
xor UO_1222 (O_1222,N_18770,N_17378);
and UO_1223 (O_1223,N_17423,N_16682);
nand UO_1224 (O_1224,N_16585,N_17341);
nand UO_1225 (O_1225,N_19398,N_17662);
nand UO_1226 (O_1226,N_16586,N_16556);
nand UO_1227 (O_1227,N_18617,N_17446);
or UO_1228 (O_1228,N_17841,N_19170);
nor UO_1229 (O_1229,N_17850,N_17470);
nor UO_1230 (O_1230,N_17922,N_17655);
nor UO_1231 (O_1231,N_16990,N_18078);
nor UO_1232 (O_1232,N_16635,N_19356);
xor UO_1233 (O_1233,N_18998,N_17251);
and UO_1234 (O_1234,N_17468,N_16496);
or UO_1235 (O_1235,N_19508,N_19139);
nor UO_1236 (O_1236,N_18632,N_19734);
nand UO_1237 (O_1237,N_18284,N_18225);
nor UO_1238 (O_1238,N_16487,N_16446);
and UO_1239 (O_1239,N_18301,N_16197);
or UO_1240 (O_1240,N_17197,N_18030);
nor UO_1241 (O_1241,N_19888,N_19517);
xnor UO_1242 (O_1242,N_16907,N_16338);
nand UO_1243 (O_1243,N_18471,N_17760);
nand UO_1244 (O_1244,N_16904,N_16433);
nand UO_1245 (O_1245,N_16147,N_19204);
xnor UO_1246 (O_1246,N_19711,N_19972);
or UO_1247 (O_1247,N_18735,N_17066);
nand UO_1248 (O_1248,N_17973,N_19136);
or UO_1249 (O_1249,N_16712,N_18653);
or UO_1250 (O_1250,N_18903,N_18197);
nor UO_1251 (O_1251,N_18635,N_18995);
and UO_1252 (O_1252,N_18608,N_19005);
nand UO_1253 (O_1253,N_19596,N_19619);
nor UO_1254 (O_1254,N_17306,N_17445);
nand UO_1255 (O_1255,N_18959,N_16588);
nand UO_1256 (O_1256,N_17620,N_17414);
and UO_1257 (O_1257,N_16448,N_18752);
nor UO_1258 (O_1258,N_18949,N_19705);
xor UO_1259 (O_1259,N_17159,N_19185);
nand UO_1260 (O_1260,N_17763,N_19078);
nand UO_1261 (O_1261,N_18548,N_16440);
xnor UO_1262 (O_1262,N_16885,N_18085);
xnor UO_1263 (O_1263,N_17926,N_16241);
xor UO_1264 (O_1264,N_17908,N_16838);
and UO_1265 (O_1265,N_19366,N_19992);
and UO_1266 (O_1266,N_16839,N_19982);
nand UO_1267 (O_1267,N_17966,N_17657);
nor UO_1268 (O_1268,N_19612,N_18083);
xor UO_1269 (O_1269,N_19816,N_16235);
and UO_1270 (O_1270,N_18241,N_16019);
nand UO_1271 (O_1271,N_17735,N_17026);
nand UO_1272 (O_1272,N_16691,N_19135);
xnor UO_1273 (O_1273,N_16742,N_16114);
and UO_1274 (O_1274,N_17597,N_19680);
and UO_1275 (O_1275,N_18602,N_16823);
nand UO_1276 (O_1276,N_16266,N_19032);
nand UO_1277 (O_1277,N_17069,N_16199);
xnor UO_1278 (O_1278,N_17810,N_18388);
xor UO_1279 (O_1279,N_19976,N_17172);
and UO_1280 (O_1280,N_16072,N_17704);
and UO_1281 (O_1281,N_19062,N_16978);
nand UO_1282 (O_1282,N_17154,N_18967);
and UO_1283 (O_1283,N_17241,N_17638);
or UO_1284 (O_1284,N_17398,N_16371);
or UO_1285 (O_1285,N_19838,N_19281);
and UO_1286 (O_1286,N_19245,N_17677);
or UO_1287 (O_1287,N_18591,N_17304);
nand UO_1288 (O_1288,N_19615,N_18101);
nor UO_1289 (O_1289,N_17882,N_19446);
nor UO_1290 (O_1290,N_17961,N_17921);
nor UO_1291 (O_1291,N_18029,N_16478);
nand UO_1292 (O_1292,N_17578,N_16896);
and UO_1293 (O_1293,N_18205,N_19199);
and UO_1294 (O_1294,N_18282,N_16957);
nor UO_1295 (O_1295,N_17951,N_19662);
nand UO_1296 (O_1296,N_18402,N_16378);
and UO_1297 (O_1297,N_17795,N_16362);
nand UO_1298 (O_1298,N_18279,N_17969);
and UO_1299 (O_1299,N_17945,N_19539);
xor UO_1300 (O_1300,N_17740,N_17645);
xor UO_1301 (O_1301,N_19318,N_17832);
or UO_1302 (O_1302,N_18153,N_18359);
or UO_1303 (O_1303,N_18595,N_17225);
nand UO_1304 (O_1304,N_16471,N_18847);
nand UO_1305 (O_1305,N_16624,N_16898);
xnor UO_1306 (O_1306,N_16326,N_18824);
or UO_1307 (O_1307,N_16892,N_19270);
or UO_1308 (O_1308,N_16026,N_18596);
xnor UO_1309 (O_1309,N_19809,N_17370);
or UO_1310 (O_1310,N_18634,N_19304);
and UO_1311 (O_1311,N_17475,N_19027);
xnor UO_1312 (O_1312,N_16305,N_18271);
nor UO_1313 (O_1313,N_19513,N_18309);
xnor UO_1314 (O_1314,N_19939,N_18409);
nor UO_1315 (O_1315,N_17668,N_18408);
and UO_1316 (O_1316,N_17044,N_16107);
nor UO_1317 (O_1317,N_19834,N_17826);
and UO_1318 (O_1318,N_19001,N_16402);
nand UO_1319 (O_1319,N_17282,N_18915);
and UO_1320 (O_1320,N_17608,N_19659);
xnor UO_1321 (O_1321,N_18393,N_19247);
or UO_1322 (O_1322,N_19189,N_18638);
nand UO_1323 (O_1323,N_18360,N_17083);
xor UO_1324 (O_1324,N_18270,N_18483);
nor UO_1325 (O_1325,N_16564,N_16523);
and UO_1326 (O_1326,N_17120,N_18840);
nand UO_1327 (O_1327,N_16361,N_19967);
xor UO_1328 (O_1328,N_16336,N_16779);
nand UO_1329 (O_1329,N_17885,N_18790);
or UO_1330 (O_1330,N_16351,N_17992);
xnor UO_1331 (O_1331,N_16825,N_19987);
xor UO_1332 (O_1332,N_19271,N_16459);
xor UO_1333 (O_1333,N_19739,N_16435);
and UO_1334 (O_1334,N_19003,N_18240);
or UO_1335 (O_1335,N_16329,N_16908);
nor UO_1336 (O_1336,N_18032,N_17749);
xnor UO_1337 (O_1337,N_16516,N_18352);
nand UO_1338 (O_1338,N_19709,N_18943);
nand UO_1339 (O_1339,N_18305,N_16818);
nor UO_1340 (O_1340,N_19879,N_17455);
and UO_1341 (O_1341,N_19381,N_17432);
xor UO_1342 (O_1342,N_17335,N_19401);
nand UO_1343 (O_1343,N_19795,N_16009);
nand UO_1344 (O_1344,N_18324,N_16282);
or UO_1345 (O_1345,N_17804,N_17054);
xnor UO_1346 (O_1346,N_18295,N_17886);
nand UO_1347 (O_1347,N_16263,N_19503);
or UO_1348 (O_1348,N_19852,N_19645);
or UO_1349 (O_1349,N_19129,N_16252);
nand UO_1350 (O_1350,N_16482,N_17745);
and UO_1351 (O_1351,N_17587,N_17058);
or UO_1352 (O_1352,N_17968,N_16445);
nand UO_1353 (O_1353,N_18417,N_19260);
or UO_1354 (O_1354,N_16348,N_19655);
nor UO_1355 (O_1355,N_17346,N_19208);
or UO_1356 (O_1356,N_16956,N_17178);
nor UO_1357 (O_1357,N_18650,N_16319);
xor UO_1358 (O_1358,N_16552,N_17340);
xnor UO_1359 (O_1359,N_16154,N_16590);
xor UO_1360 (O_1360,N_18701,N_16886);
nand UO_1361 (O_1361,N_19843,N_18084);
or UO_1362 (O_1362,N_17029,N_17768);
or UO_1363 (O_1363,N_18050,N_17701);
xnor UO_1364 (O_1364,N_18478,N_18693);
nor UO_1365 (O_1365,N_17356,N_17321);
nand UO_1366 (O_1366,N_16813,N_19516);
nand UO_1367 (O_1367,N_17188,N_19339);
nand UO_1368 (O_1368,N_17877,N_19132);
or UO_1369 (O_1369,N_17776,N_17817);
xnor UO_1370 (O_1370,N_17393,N_19175);
nand UO_1371 (O_1371,N_17508,N_18342);
or UO_1372 (O_1372,N_18538,N_18946);
nor UO_1373 (O_1373,N_16732,N_16783);
nor UO_1374 (O_1374,N_19953,N_18065);
xor UO_1375 (O_1375,N_17927,N_17193);
nand UO_1376 (O_1376,N_16511,N_16652);
and UO_1377 (O_1377,N_18079,N_16384);
nand UO_1378 (O_1378,N_19212,N_18604);
and UO_1379 (O_1379,N_18123,N_17375);
and UO_1380 (O_1380,N_16443,N_19331);
and UO_1381 (O_1381,N_16227,N_18247);
xor UO_1382 (O_1382,N_16239,N_19807);
nand UO_1383 (O_1383,N_19033,N_16650);
and UO_1384 (O_1384,N_16580,N_18771);
or UO_1385 (O_1385,N_17898,N_17531);
or UO_1386 (O_1386,N_16984,N_19215);
and UO_1387 (O_1387,N_17611,N_16562);
or UO_1388 (O_1388,N_16113,N_16533);
nand UO_1389 (O_1389,N_17086,N_19089);
or UO_1390 (O_1390,N_16639,N_18221);
nor UO_1391 (O_1391,N_16178,N_19708);
nand UO_1392 (O_1392,N_17252,N_17616);
and UO_1393 (O_1393,N_19229,N_18330);
nor UO_1394 (O_1394,N_19481,N_17285);
nand UO_1395 (O_1395,N_19337,N_19489);
or UO_1396 (O_1396,N_19742,N_19298);
or UO_1397 (O_1397,N_16608,N_17305);
xor UO_1398 (O_1398,N_17160,N_17024);
and UO_1399 (O_1399,N_19288,N_17457);
xnor UO_1400 (O_1400,N_17664,N_16126);
nor UO_1401 (O_1401,N_16643,N_18971);
or UO_1402 (O_1402,N_18680,N_18230);
nor UO_1403 (O_1403,N_17753,N_18603);
and UO_1404 (O_1404,N_18088,N_18174);
or UO_1405 (O_1405,N_18164,N_19859);
nor UO_1406 (O_1406,N_18227,N_16024);
nand UO_1407 (O_1407,N_18061,N_19586);
xor UO_1408 (O_1408,N_19195,N_17844);
or UO_1409 (O_1409,N_16851,N_18105);
xnor UO_1410 (O_1410,N_18781,N_16557);
nand UO_1411 (O_1411,N_19418,N_18811);
nand UO_1412 (O_1412,N_17422,N_19283);
nor UO_1413 (O_1413,N_19591,N_18068);
or UO_1414 (O_1414,N_19892,N_16367);
and UO_1415 (O_1415,N_16723,N_17812);
nand UO_1416 (O_1416,N_19044,N_18961);
and UO_1417 (O_1417,N_17982,N_17342);
xnor UO_1418 (O_1418,N_19522,N_16424);
xor UO_1419 (O_1419,N_16619,N_19156);
xor UO_1420 (O_1420,N_18354,N_18865);
and UO_1421 (O_1421,N_17635,N_16888);
xor UO_1422 (O_1422,N_18944,N_17904);
nor UO_1423 (O_1423,N_19459,N_18118);
xnor UO_1424 (O_1424,N_17219,N_18236);
nand UO_1425 (O_1425,N_18807,N_16060);
nor UO_1426 (O_1426,N_17263,N_16706);
and UO_1427 (O_1427,N_17105,N_17162);
xnor UO_1428 (O_1428,N_18821,N_17007);
or UO_1429 (O_1429,N_19851,N_17600);
xnor UO_1430 (O_1430,N_16120,N_16476);
and UO_1431 (O_1431,N_19190,N_16095);
and UO_1432 (O_1432,N_17837,N_18828);
nor UO_1433 (O_1433,N_16530,N_19487);
or UO_1434 (O_1434,N_19999,N_16330);
and UO_1435 (O_1435,N_18459,N_17822);
nor UO_1436 (O_1436,N_17673,N_16715);
nor UO_1437 (O_1437,N_18486,N_19721);
and UO_1438 (O_1438,N_19255,N_19979);
xor UO_1439 (O_1439,N_16513,N_18904);
nand UO_1440 (O_1440,N_17020,N_17322);
nor UO_1441 (O_1441,N_17045,N_16704);
nand UO_1442 (O_1442,N_16616,N_17353);
and UO_1443 (O_1443,N_18411,N_18020);
nand UO_1444 (O_1444,N_16729,N_17695);
or UO_1445 (O_1445,N_19122,N_16093);
nand UO_1446 (O_1446,N_17210,N_19644);
nand UO_1447 (O_1447,N_18312,N_16444);
xor UO_1448 (O_1448,N_16050,N_19829);
nand UO_1449 (O_1449,N_17389,N_19289);
nor UO_1450 (O_1450,N_19685,N_18809);
and UO_1451 (O_1451,N_18234,N_19699);
and UO_1452 (O_1452,N_19567,N_17387);
nor UO_1453 (O_1453,N_17323,N_17101);
xor UO_1454 (O_1454,N_18869,N_18396);
nand UO_1455 (O_1455,N_16473,N_19460);
and UO_1456 (O_1456,N_16143,N_18785);
xor UO_1457 (O_1457,N_16059,N_18387);
nor UO_1458 (O_1458,N_18299,N_19282);
or UO_1459 (O_1459,N_16495,N_18572);
and UO_1460 (O_1460,N_17057,N_18529);
and UO_1461 (O_1461,N_19144,N_16146);
nand UO_1462 (O_1462,N_17062,N_19812);
xnor UO_1463 (O_1463,N_18059,N_18386);
or UO_1464 (O_1464,N_18055,N_19120);
xor UO_1465 (O_1465,N_19494,N_16006);
and UO_1466 (O_1466,N_16294,N_19483);
xnor UO_1467 (O_1467,N_17524,N_16999);
xnor UO_1468 (O_1468,N_16814,N_18358);
xnor UO_1469 (O_1469,N_17814,N_16922);
or UO_1470 (O_1470,N_19745,N_16989);
nor UO_1471 (O_1471,N_17055,N_17496);
nor UO_1472 (O_1472,N_17211,N_19622);
nand UO_1473 (O_1473,N_16056,N_18147);
and UO_1474 (O_1474,N_19924,N_16931);
xor UO_1475 (O_1475,N_19021,N_16479);
or UO_1476 (O_1476,N_16721,N_19437);
nor UO_1477 (O_1477,N_19161,N_17338);
nand UO_1478 (O_1478,N_16504,N_18704);
nand UO_1479 (O_1479,N_18760,N_17528);
or UO_1480 (O_1480,N_18780,N_19732);
nand UO_1481 (O_1481,N_18035,N_19694);
nor UO_1482 (O_1482,N_18739,N_18452);
nor UO_1483 (O_1483,N_16177,N_18228);
xnor UO_1484 (O_1484,N_16602,N_18670);
or UO_1485 (O_1485,N_16425,N_19325);
nand UO_1486 (O_1486,N_16550,N_18041);
xor UO_1487 (O_1487,N_17023,N_17944);
xnor UO_1488 (O_1488,N_16395,N_16971);
nand UO_1489 (O_1489,N_18768,N_16968);
nor UO_1490 (O_1490,N_17209,N_16699);
or UO_1491 (O_1491,N_18708,N_16396);
or UO_1492 (O_1492,N_19955,N_18644);
nand UO_1493 (O_1493,N_16474,N_19158);
and UO_1494 (O_1494,N_18819,N_18750);
nor UO_1495 (O_1495,N_17563,N_19464);
nor UO_1496 (O_1496,N_18997,N_18130);
and UO_1497 (O_1497,N_16864,N_19390);
or UO_1498 (O_1498,N_16099,N_18956);
or UO_1499 (O_1499,N_16992,N_16859);
nand UO_1500 (O_1500,N_19151,N_19332);
nor UO_1501 (O_1501,N_16246,N_17625);
nand UO_1502 (O_1502,N_17212,N_16339);
xor UO_1503 (O_1503,N_18838,N_18327);
or UO_1504 (O_1504,N_16998,N_16198);
nor UO_1505 (O_1505,N_17094,N_19319);
nor UO_1506 (O_1506,N_19917,N_19050);
nand UO_1507 (O_1507,N_18266,N_17990);
and UO_1508 (O_1508,N_16834,N_16480);
or UO_1509 (O_1509,N_16032,N_19784);
nor UO_1510 (O_1510,N_19938,N_19799);
xor UO_1511 (O_1511,N_18801,N_17279);
xnor UO_1512 (O_1512,N_19348,N_19369);
or UO_1513 (O_1513,N_19832,N_16676);
or UO_1514 (O_1514,N_18434,N_17847);
and UO_1515 (O_1515,N_19780,N_18037);
nor UO_1516 (O_1516,N_16379,N_18158);
nor UO_1517 (O_1517,N_18761,N_19684);
nand UO_1518 (O_1518,N_16835,N_16317);
and UO_1519 (O_1519,N_16755,N_18753);
nand UO_1520 (O_1520,N_16209,N_17838);
xor UO_1521 (O_1521,N_17731,N_18472);
nor UO_1522 (O_1522,N_18210,N_17495);
xor UO_1523 (O_1523,N_17687,N_18081);
xor UO_1524 (O_1524,N_18661,N_19216);
xor UO_1525 (O_1525,N_17794,N_18676);
and UO_1526 (O_1526,N_17231,N_19626);
or UO_1527 (O_1527,N_16521,N_17790);
nand UO_1528 (O_1528,N_16020,N_19884);
nand UO_1529 (O_1529,N_18376,N_19375);
nand UO_1530 (O_1530,N_17594,N_19903);
and UO_1531 (O_1531,N_16418,N_18293);
and UO_1532 (O_1532,N_16937,N_19869);
nor UO_1533 (O_1533,N_18746,N_17949);
and UO_1534 (O_1534,N_19677,N_18181);
xor UO_1535 (O_1535,N_19704,N_19823);
or UO_1536 (O_1536,N_16951,N_17722);
and UO_1537 (O_1537,N_17779,N_17893);
nor UO_1538 (O_1538,N_17907,N_16303);
or UO_1539 (O_1539,N_17004,N_18989);
xnor UO_1540 (O_1540,N_16309,N_16134);
nand UO_1541 (O_1541,N_16775,N_16843);
xor UO_1542 (O_1542,N_17195,N_17108);
and UO_1543 (O_1543,N_19505,N_18252);
xnor UO_1544 (O_1544,N_16849,N_19501);
or UO_1545 (O_1545,N_18934,N_17436);
or UO_1546 (O_1546,N_16377,N_18918);
or UO_1547 (O_1547,N_16259,N_18964);
nor UO_1548 (O_1548,N_18767,N_17818);
and UO_1549 (O_1549,N_18620,N_18939);
nand UO_1550 (O_1550,N_17240,N_18586);
and UO_1551 (O_1551,N_16493,N_17474);
nor UO_1552 (O_1552,N_17444,N_17186);
or UO_1553 (O_1553,N_16647,N_19432);
xnor UO_1554 (O_1554,N_19183,N_16748);
xnor UO_1555 (O_1555,N_17394,N_17005);
nor UO_1556 (O_1556,N_16862,N_18975);
nor UO_1557 (O_1557,N_17823,N_18285);
nand UO_1558 (O_1558,N_18067,N_17451);
xnor UO_1559 (O_1559,N_16711,N_18852);
xnor UO_1560 (O_1560,N_16689,N_19627);
or UO_1561 (O_1561,N_17571,N_18910);
xnor UO_1562 (O_1562,N_19111,N_17124);
or UO_1563 (O_1563,N_19782,N_17552);
nor UO_1564 (O_1564,N_18849,N_18397);
nor UO_1565 (O_1565,N_18412,N_18107);
nor UO_1566 (O_1566,N_17276,N_16784);
or UO_1567 (O_1567,N_16674,N_19162);
xor UO_1568 (O_1568,N_16740,N_19110);
nor UO_1569 (O_1569,N_16574,N_16966);
and UO_1570 (O_1570,N_16716,N_19118);
nand UO_1571 (O_1571,N_19905,N_17970);
or UO_1572 (O_1572,N_18137,N_17852);
nand UO_1573 (O_1573,N_18682,N_17534);
nand UO_1574 (O_1574,N_17708,N_17343);
and UO_1575 (O_1575,N_17397,N_16233);
or UO_1576 (O_1576,N_18987,N_18269);
and UO_1577 (O_1577,N_16345,N_18692);
nor UO_1578 (O_1578,N_19425,N_17290);
or UO_1579 (O_1579,N_19546,N_17567);
and UO_1580 (O_1580,N_19253,N_17960);
nor UO_1581 (O_1581,N_17917,N_19174);
and UO_1582 (O_1582,N_16200,N_18196);
xnor UO_1583 (O_1583,N_19201,N_19893);
xnor UO_1584 (O_1584,N_19130,N_16801);
xor UO_1585 (O_1585,N_16373,N_18474);
or UO_1586 (O_1586,N_18005,N_18226);
or UO_1587 (O_1587,N_18169,N_17691);
or UO_1588 (O_1588,N_18063,N_16038);
and UO_1589 (O_1589,N_17396,N_17164);
xor UO_1590 (O_1590,N_19796,N_19991);
and UO_1591 (O_1591,N_18506,N_17244);
xor UO_1592 (O_1592,N_17256,N_17367);
xnor UO_1593 (O_1593,N_17499,N_18777);
nor UO_1594 (O_1594,N_16887,N_19733);
xnor UO_1595 (O_1595,N_19760,N_19810);
nand UO_1596 (O_1596,N_19574,N_16102);
nand UO_1597 (O_1597,N_17181,N_16502);
and UO_1598 (O_1598,N_16185,N_19386);
nand UO_1599 (O_1599,N_18399,N_17199);
and UO_1600 (O_1600,N_19978,N_17273);
nor UO_1601 (O_1601,N_16452,N_18374);
nor UO_1602 (O_1602,N_17032,N_19994);
or UO_1603 (O_1603,N_16640,N_18370);
and UO_1604 (O_1604,N_16950,N_17766);
nor UO_1605 (O_1605,N_16754,N_16077);
xor UO_1606 (O_1606,N_17648,N_16430);
nand UO_1607 (O_1607,N_16880,N_18481);
nand UO_1608 (O_1608,N_16091,N_16498);
xnor UO_1609 (O_1609,N_19474,N_18004);
nor UO_1610 (O_1610,N_18183,N_19594);
and UO_1611 (O_1611,N_18237,N_19527);
nand UO_1612 (O_1612,N_18013,N_17228);
xor UO_1613 (O_1613,N_16451,N_19746);
xor UO_1614 (O_1614,N_16321,N_19294);
and UO_1615 (O_1615,N_16774,N_19176);
or UO_1616 (O_1616,N_18366,N_16016);
nor UO_1617 (O_1617,N_16352,N_17797);
and UO_1618 (O_1618,N_17652,N_19261);
nor UO_1619 (O_1619,N_19896,N_17122);
nand UO_1620 (O_1620,N_17813,N_17682);
or UO_1621 (O_1621,N_18528,N_19095);
nor UO_1622 (O_1622,N_18681,N_18194);
nand UO_1623 (O_1623,N_19155,N_17716);
or UO_1624 (O_1624,N_19091,N_18992);
nand UO_1625 (O_1625,N_19012,N_17309);
nor UO_1626 (O_1626,N_18520,N_17247);
or UO_1627 (O_1627,N_16932,N_18140);
and UO_1628 (O_1628,N_18542,N_19379);
or UO_1629 (O_1629,N_16191,N_18453);
nand UO_1630 (O_1630,N_17719,N_19878);
nor UO_1631 (O_1631,N_17175,N_18957);
xor UO_1632 (O_1632,N_18211,N_16694);
and UO_1633 (O_1633,N_18361,N_17277);
and UO_1634 (O_1634,N_17413,N_17299);
or UO_1635 (O_1635,N_19066,N_18794);
nor UO_1636 (O_1636,N_18308,N_17076);
nand UO_1637 (O_1637,N_19766,N_18614);
xor UO_1638 (O_1638,N_17194,N_17334);
nor UO_1639 (O_1639,N_19719,N_16108);
nor UO_1640 (O_1640,N_17016,N_18633);
and UO_1641 (O_1641,N_19706,N_18546);
and UO_1642 (O_1642,N_17294,N_16225);
or UO_1643 (O_1643,N_18332,N_17246);
xnor UO_1644 (O_1644,N_18860,N_16269);
nand UO_1645 (O_1645,N_18763,N_18450);
nand UO_1646 (O_1646,N_19324,N_19488);
nor UO_1647 (O_1647,N_16811,N_18922);
xor UO_1648 (O_1648,N_19558,N_19224);
nand UO_1649 (O_1649,N_19861,N_19918);
or UO_1650 (O_1650,N_17134,N_16981);
and UO_1651 (O_1651,N_19184,N_17183);
xor UO_1652 (O_1652,N_18432,N_16342);
xnor UO_1653 (O_1653,N_19168,N_17777);
nand UO_1654 (O_1654,N_19793,N_19914);
nor UO_1655 (O_1655,N_19407,N_16945);
and UO_1656 (O_1656,N_16548,N_19303);
and UO_1657 (O_1657,N_17060,N_16597);
or UO_1658 (O_1658,N_19235,N_16621);
xor UO_1659 (O_1659,N_18132,N_19045);
nand UO_1660 (O_1660,N_16421,N_17488);
or UO_1661 (O_1661,N_18791,N_17145);
xor UO_1662 (O_1662,N_18015,N_19724);
or UO_1663 (O_1663,N_18429,N_18709);
nand UO_1664 (O_1664,N_17871,N_18575);
or UO_1665 (O_1665,N_17585,N_18727);
or UO_1666 (O_1666,N_17840,N_19686);
xnor UO_1667 (O_1667,N_17243,N_19466);
or UO_1668 (O_1668,N_18578,N_16575);
nor UO_1669 (O_1669,N_18131,N_19054);
or UO_1670 (O_1670,N_18161,N_18901);
nor UO_1671 (O_1671,N_17752,N_17962);
nand UO_1672 (O_1672,N_19668,N_19963);
nand UO_1673 (O_1673,N_17454,N_18978);
xor UO_1674 (O_1674,N_16340,N_18064);
nand UO_1675 (O_1675,N_18889,N_19966);
nand UO_1676 (O_1676,N_19160,N_16903);
nand UO_1677 (O_1677,N_19473,N_18053);
nor UO_1678 (O_1678,N_19342,N_19112);
nand UO_1679 (O_1679,N_19776,N_16765);
and UO_1680 (O_1680,N_17688,N_18116);
nor UO_1681 (O_1681,N_17911,N_16675);
xor UO_1682 (O_1682,N_18439,N_19367);
xor UO_1683 (O_1683,N_16167,N_19336);
nand UO_1684 (O_1684,N_16545,N_16565);
nor UO_1685 (O_1685,N_16156,N_18769);
nor UO_1686 (O_1686,N_19227,N_16570);
nor UO_1687 (O_1687,N_17848,N_16109);
xor UO_1688 (O_1688,N_19393,N_17526);
and UO_1689 (O_1689,N_19347,N_17141);
or UO_1690 (O_1690,N_19762,N_19951);
xor UO_1691 (O_1691,N_18592,N_17743);
and UO_1692 (O_1692,N_18357,N_18394);
or UO_1693 (O_1693,N_19860,N_18214);
or UO_1694 (O_1694,N_16663,N_16558);
or UO_1695 (O_1695,N_19906,N_18058);
nand UO_1696 (O_1696,N_18089,N_17979);
nor UO_1697 (O_1697,N_19610,N_19103);
xor UO_1698 (O_1698,N_17344,N_17048);
and UO_1699 (O_1699,N_18815,N_19361);
xor UO_1700 (O_1700,N_19556,N_18420);
or UO_1701 (O_1701,N_19146,N_18336);
nor UO_1702 (O_1702,N_17416,N_17298);
and UO_1703 (O_1703,N_18171,N_17192);
nor UO_1704 (O_1704,N_19510,N_18509);
xor UO_1705 (O_1705,N_19105,N_19405);
or UO_1706 (O_1706,N_16219,N_17805);
or UO_1707 (O_1707,N_17462,N_19531);
nor UO_1708 (O_1708,N_16939,N_16468);
nor UO_1709 (O_1709,N_16940,N_18658);
and UO_1710 (O_1710,N_16297,N_16271);
or UO_1711 (O_1711,N_18179,N_19826);
or UO_1712 (O_1712,N_16462,N_16848);
or UO_1713 (O_1713,N_18350,N_19678);
nand UO_1714 (O_1714,N_17697,N_18348);
xor UO_1715 (O_1715,N_16010,N_18762);
xnor UO_1716 (O_1716,N_16278,N_17788);
and UO_1717 (O_1717,N_18331,N_16469);
and UO_1718 (O_1718,N_18765,N_18522);
nor UO_1719 (O_1719,N_17789,N_17860);
nor UO_1720 (O_1720,N_16244,N_16052);
nand UO_1721 (O_1721,N_19666,N_17538);
nor UO_1722 (O_1722,N_18613,N_17775);
nor UO_1723 (O_1723,N_19738,N_18945);
nor UO_1724 (O_1724,N_19061,N_19529);
nand UO_1725 (O_1725,N_19172,N_16152);
nor UO_1726 (O_1726,N_19434,N_16965);
and UO_1727 (O_1727,N_16066,N_19865);
and UO_1728 (O_1728,N_19065,N_18831);
xnor UO_1729 (O_1729,N_18242,N_19629);
nor UO_1730 (O_1730,N_17870,N_19675);
nand UO_1731 (O_1731,N_18714,N_18985);
nor UO_1732 (O_1732,N_17603,N_16868);
nor UO_1733 (O_1733,N_18505,N_19408);
nand UO_1734 (O_1734,N_16980,N_18159);
and UO_1735 (O_1735,N_17527,N_19107);
nor UO_1736 (O_1736,N_17778,N_19774);
xnor UO_1737 (O_1737,N_16626,N_18724);
or UO_1738 (O_1738,N_18594,N_18806);
or UO_1739 (O_1739,N_18896,N_17180);
nor UO_1740 (O_1740,N_16265,N_17819);
or UO_1741 (O_1741,N_17786,N_19907);
and UO_1742 (O_1742,N_18351,N_18297);
xor UO_1743 (O_1743,N_19194,N_19928);
nor UO_1744 (O_1744,N_17675,N_16389);
or UO_1745 (O_1745,N_18574,N_19846);
nand UO_1746 (O_1746,N_17613,N_16081);
nor UO_1747 (O_1747,N_18582,N_19783);
and UO_1748 (O_1748,N_16104,N_19912);
nor UO_1749 (O_1749,N_19246,N_19243);
xor UO_1750 (O_1750,N_16441,N_19431);
nor UO_1751 (O_1751,N_18071,N_16168);
xnor UO_1752 (O_1752,N_16192,N_18703);
nor UO_1753 (O_1753,N_17100,N_18907);
and UO_1754 (O_1754,N_17769,N_16350);
nor UO_1755 (O_1755,N_17863,N_17971);
xor UO_1756 (O_1756,N_16751,N_18526);
nor UO_1757 (O_1757,N_16044,N_16622);
nand UO_1758 (O_1758,N_18341,N_18618);
and UO_1759 (O_1759,N_16810,N_17012);
nor UO_1760 (O_1760,N_18190,N_18861);
and UO_1761 (O_1761,N_17485,N_18435);
nand UO_1762 (O_1762,N_16161,N_17737);
and UO_1763 (O_1763,N_19691,N_19014);
xnor UO_1764 (O_1764,N_16442,N_16730);
and UO_1765 (O_1765,N_17878,N_18125);
xnor UO_1766 (O_1766,N_18963,N_17383);
and UO_1767 (O_1767,N_18052,N_16267);
and UO_1768 (O_1768,N_16672,N_16092);
xor UO_1769 (O_1769,N_19296,N_19013);
xor UO_1770 (O_1770,N_16243,N_17088);
and UO_1771 (O_1771,N_19788,N_18245);
nor UO_1772 (O_1772,N_17696,N_18287);
nand UO_1773 (O_1773,N_18229,N_17902);
nand UO_1774 (O_1774,N_18503,N_16963);
xnor UO_1775 (O_1775,N_16276,N_17464);
or UO_1776 (O_1776,N_19818,N_16909);
nand UO_1777 (O_1777,N_17504,N_16397);
and UO_1778 (O_1778,N_17424,N_18016);
and UO_1779 (O_1779,N_19427,N_18851);
or UO_1780 (O_1780,N_19378,N_18391);
xor UO_1781 (O_1781,N_18049,N_18841);
and UO_1782 (O_1782,N_18611,N_18779);
nor UO_1783 (O_1783,N_16503,N_17581);
xor UO_1784 (O_1784,N_19502,N_17640);
nand UO_1785 (O_1785,N_17509,N_18175);
nand UO_1786 (O_1786,N_19792,N_19521);
nand UO_1787 (O_1787,N_16359,N_19359);
or UO_1788 (O_1788,N_17986,N_17798);
nand UO_1789 (O_1789,N_17659,N_19700);
and UO_1790 (O_1790,N_17833,N_16882);
or UO_1791 (O_1791,N_19053,N_19075);
or UO_1792 (O_1792,N_16906,N_17896);
nand UO_1793 (O_1793,N_16837,N_18776);
nor UO_1794 (O_1794,N_17296,N_18702);
nor UO_1795 (O_1795,N_16076,N_16086);
and UO_1796 (O_1796,N_17000,N_17899);
xnor UO_1797 (O_1797,N_18213,N_16262);
xnor UO_1798 (O_1798,N_17487,N_16231);
nand UO_1799 (O_1799,N_18482,N_17056);
and UO_1800 (O_1800,N_17392,N_18723);
nor UO_1801 (O_1801,N_17617,N_17224);
or UO_1802 (O_1802,N_16257,N_19693);
and UO_1803 (O_1803,N_16658,N_16510);
xnor UO_1804 (O_1804,N_17235,N_17591);
nor UO_1805 (O_1805,N_18311,N_19206);
and UO_1806 (O_1806,N_18464,N_17429);
or UO_1807 (O_1807,N_17419,N_17698);
xnor UO_1808 (O_1808,N_16210,N_18664);
nand UO_1809 (O_1809,N_18189,N_18488);
nor UO_1810 (O_1810,N_19453,N_17061);
nand UO_1811 (O_1811,N_16437,N_16136);
and UO_1812 (O_1812,N_18476,N_18338);
nor UO_1813 (O_1813,N_16180,N_17412);
or UO_1814 (O_1814,N_16075,N_17307);
or UO_1815 (O_1815,N_18859,N_19321);
xnor UO_1816 (O_1816,N_16873,N_19575);
nand UO_1817 (O_1817,N_16522,N_18424);
nand UO_1818 (O_1818,N_18060,N_16531);
and UO_1819 (O_1819,N_17564,N_19219);
xnor UO_1820 (O_1820,N_19147,N_18390);
nor UO_1821 (O_1821,N_19988,N_16335);
nor UO_1822 (O_1822,N_18751,N_17479);
nor UO_1823 (O_1823,N_16960,N_16298);
and UO_1824 (O_1824,N_17569,N_17574);
nand UO_1825 (O_1825,N_18683,N_18246);
and UO_1826 (O_1826,N_17576,N_16331);
xnor UO_1827 (O_1827,N_18532,N_16913);
or UO_1828 (O_1828,N_18710,N_19307);
xnor UO_1829 (O_1829,N_18876,N_17615);
or UO_1830 (O_1830,N_17995,N_18104);
nor UO_1831 (O_1831,N_17442,N_18517);
or UO_1832 (O_1832,N_18630,N_18262);
nand UO_1833 (O_1833,N_16611,N_18062);
nand UO_1834 (O_1834,N_17539,N_19822);
nand UO_1835 (O_1835,N_17998,N_17734);
or UO_1836 (O_1836,N_17063,N_17940);
or UO_1837 (O_1837,N_19858,N_17135);
or UO_1838 (O_1838,N_16642,N_18788);
and UO_1839 (O_1839,N_17430,N_17136);
and UO_1840 (O_1840,N_17401,N_18825);
xor UO_1841 (O_1841,N_18802,N_16046);
nor UO_1842 (O_1842,N_16100,N_17865);
and UO_1843 (O_1843,N_18686,N_16594);
xor UO_1844 (O_1844,N_18521,N_16166);
and UO_1845 (O_1845,N_19856,N_17836);
nor UO_1846 (O_1846,N_16022,N_17351);
nor UO_1847 (O_1847,N_17503,N_17941);
nand UO_1848 (O_1848,N_16141,N_16465);
nor UO_1849 (O_1849,N_16343,N_18562);
nand UO_1850 (O_1850,N_17498,N_17168);
and UO_1851 (O_1851,N_17447,N_16568);
xnor UO_1852 (O_1852,N_17570,N_18566);
xnor UO_1853 (O_1853,N_19950,N_17540);
or UO_1854 (O_1854,N_17142,N_18640);
or UO_1855 (O_1855,N_19256,N_19604);
xor UO_1856 (O_1856,N_19770,N_17113);
and UO_1857 (O_1857,N_18009,N_17815);
and UO_1858 (O_1858,N_16713,N_17003);
nor UO_1859 (O_1859,N_19841,N_19964);
nor UO_1860 (O_1860,N_18508,N_17929);
nand UO_1861 (O_1861,N_19306,N_16065);
or UO_1862 (O_1862,N_19329,N_17497);
nor UO_1863 (O_1863,N_17381,N_16846);
nor UO_1864 (O_1864,N_17642,N_19900);
and UO_1865 (O_1865,N_18253,N_19753);
xnor UO_1866 (O_1866,N_19942,N_18507);
and UO_1867 (O_1867,N_19213,N_16188);
nor UO_1868 (O_1868,N_17589,N_19805);
xor UO_1869 (O_1869,N_19242,N_16771);
and UO_1870 (O_1870,N_19729,N_16201);
and UO_1871 (O_1871,N_18561,N_18212);
or UO_1872 (O_1872,N_16411,N_17516);
xor UO_1873 (O_1873,N_17628,N_19429);
xor UO_1874 (O_1874,N_17440,N_18203);
and UO_1875 (O_1875,N_19205,N_17480);
xor UO_1876 (O_1876,N_19932,N_18641);
nand UO_1877 (O_1877,N_19773,N_19372);
nand UO_1878 (O_1878,N_18244,N_18853);
and UO_1879 (O_1879,N_16547,N_18976);
and UO_1880 (O_1880,N_18894,N_18745);
xnor UO_1881 (O_1881,N_17771,N_16787);
xor UO_1882 (O_1882,N_18835,N_17614);
nor UO_1883 (O_1883,N_18014,N_17220);
xnor UO_1884 (O_1884,N_18377,N_19345);
and UO_1885 (O_1885,N_17972,N_19198);
nor UO_1886 (O_1886,N_17107,N_19169);
and UO_1887 (O_1887,N_18202,N_16947);
nor UO_1888 (O_1888,N_16753,N_16103);
xnor UO_1889 (O_1889,N_16349,N_16130);
or UO_1890 (O_1890,N_17996,N_16983);
or UO_1891 (O_1891,N_18947,N_18403);
or UO_1892 (O_1892,N_18462,N_19864);
and UO_1893 (O_1893,N_18504,N_19457);
and UO_1894 (O_1894,N_19015,N_18315);
nor UO_1895 (O_1895,N_16800,N_17449);
and UO_1896 (O_1896,N_18656,N_16975);
nor UO_1897 (O_1897,N_17139,N_17404);
nand UO_1898 (O_1898,N_17984,N_16758);
or UO_1899 (O_1899,N_16701,N_18668);
xor UO_1900 (O_1900,N_17179,N_16375);
xor UO_1901 (O_1901,N_17706,N_19394);
xnor UO_1902 (O_1902,N_17151,N_16542);
nor UO_1903 (O_1903,N_18173,N_18426);
nor UO_1904 (O_1904,N_19341,N_17043);
nor UO_1905 (O_1905,N_16449,N_17208);
nor UO_1906 (O_1906,N_17386,N_17773);
nand UO_1907 (O_1907,N_17153,N_16853);
nand UO_1908 (O_1908,N_16815,N_17660);
xnor UO_1909 (O_1909,N_17093,N_18300);
nor UO_1910 (O_1910,N_18919,N_16313);
nand UO_1911 (O_1911,N_19913,N_17846);
and UO_1912 (O_1912,N_18467,N_17245);
xor UO_1913 (O_1913,N_17950,N_17791);
xnor UO_1914 (O_1914,N_17184,N_17077);
nor UO_1915 (O_1915,N_19101,N_18320);
and UO_1916 (O_1916,N_19952,N_17880);
or UO_1917 (O_1917,N_17402,N_17117);
nor UO_1918 (O_1918,N_16280,N_19524);
or UO_1919 (O_1919,N_19661,N_16045);
nor UO_1920 (O_1920,N_17177,N_19284);
nor UO_1921 (O_1921,N_17132,N_18355);
and UO_1922 (O_1922,N_19862,N_19340);
nand UO_1923 (O_1923,N_17557,N_16290);
nand UO_1924 (O_1924,N_17254,N_16218);
nand UO_1925 (O_1925,N_19535,N_18581);
xnor UO_1926 (O_1926,N_16145,N_18565);
nor UO_1927 (O_1927,N_19872,N_16620);
nor UO_1928 (O_1928,N_18087,N_18856);
or UO_1929 (O_1929,N_19725,N_16563);
nand UO_1930 (O_1930,N_17174,N_17363);
and UO_1931 (O_1931,N_17411,N_18626);
nor UO_1932 (O_1932,N_17345,N_17493);
or UO_1933 (O_1933,N_18463,N_16817);
and UO_1934 (O_1934,N_17138,N_17476);
nor UO_1935 (O_1935,N_16215,N_18679);
or UO_1936 (O_1936,N_19041,N_19233);
nand UO_1937 (O_1937,N_16133,N_19772);
nor UO_1938 (O_1938,N_18868,N_17806);
nor UO_1939 (O_1939,N_19154,N_17075);
xor UO_1940 (O_1940,N_18736,N_16240);
nor UO_1941 (O_1941,N_18699,N_19040);
and UO_1942 (O_1942,N_18136,N_19096);
nand UO_1943 (O_1943,N_16357,N_16925);
nor UO_1944 (O_1944,N_17676,N_18827);
xnor UO_1945 (O_1945,N_18051,N_19085);
nand UO_1946 (O_1946,N_19712,N_18514);
and UO_1947 (O_1947,N_18313,N_19309);
and UO_1948 (O_1948,N_18991,N_17721);
xnor UO_1949 (O_1949,N_19365,N_18721);
nand UO_1950 (O_1950,N_17859,N_19141);
xor UO_1951 (O_1951,N_17376,N_18662);
or UO_1952 (O_1952,N_17137,N_18857);
nand UO_1953 (O_1953,N_18973,N_16592);
or UO_1954 (O_1954,N_17864,N_16328);
or UO_1955 (O_1955,N_18389,N_16646);
nor UO_1956 (O_1956,N_19723,N_17999);
nand UO_1957 (O_1957,N_17909,N_16258);
or UO_1958 (O_1958,N_19121,N_16615);
and UO_1959 (O_1959,N_16057,N_16249);
nor UO_1960 (O_1960,N_18832,N_17985);
or UO_1961 (O_1961,N_17190,N_17106);
and UO_1962 (O_1962,N_19192,N_16128);
nor UO_1963 (O_1963,N_18725,N_19469);
or UO_1964 (O_1964,N_19239,N_18480);
xor UO_1965 (O_1965,N_16064,N_18438);
or UO_1966 (O_1966,N_18133,N_16212);
xnor UO_1967 (O_1967,N_16105,N_16381);
or UO_1968 (O_1968,N_19231,N_16232);
nor UO_1969 (O_1969,N_19523,N_18006);
and UO_1970 (O_1970,N_19292,N_16051);
nand UO_1971 (O_1971,N_18666,N_17634);
and UO_1972 (O_1972,N_16293,N_19576);
or UO_1973 (O_1973,N_18799,N_17535);
nand UO_1974 (O_1974,N_18326,N_18545);
or UO_1975 (O_1975,N_17559,N_17702);
nand UO_1976 (O_1976,N_18830,N_17221);
or UO_1977 (O_1977,N_19765,N_18513);
xnor UO_1978 (O_1978,N_19496,N_16816);
xnor UO_1979 (O_1979,N_18540,N_18812);
or UO_1980 (O_1980,N_19636,N_17715);
xor UO_1981 (O_1981,N_18810,N_16781);
or UO_1982 (O_1982,N_16000,N_17450);
and UO_1983 (O_1983,N_18243,N_17560);
xnor UO_1984 (O_1984,N_16312,N_18511);
nand UO_1985 (O_1985,N_19442,N_17519);
nor UO_1986 (O_1986,N_16494,N_17947);
or UO_1987 (O_1987,N_19582,N_17140);
xnor UO_1988 (O_1988,N_18772,N_18986);
xor UO_1989 (O_1989,N_19871,N_19291);
xnor UO_1990 (O_1990,N_18275,N_16428);
nand UO_1991 (O_1991,N_19941,N_18895);
nor UO_1992 (O_1992,N_16165,N_17884);
or UO_1993 (O_1993,N_19692,N_18541);
nor UO_1994 (O_1994,N_18648,N_16483);
nor UO_1995 (O_1995,N_16872,N_19897);
xor UO_1996 (O_1996,N_17217,N_17681);
nor UO_1997 (O_1997,N_17501,N_17330);
or UO_1998 (O_1998,N_17391,N_16291);
nand UO_1999 (O_1999,N_18457,N_16527);
nand UO_2000 (O_2000,N_18635,N_18259);
or UO_2001 (O_2001,N_16960,N_19032);
xnor UO_2002 (O_2002,N_18016,N_16066);
nand UO_2003 (O_2003,N_16065,N_18899);
nand UO_2004 (O_2004,N_17737,N_16415);
xor UO_2005 (O_2005,N_16585,N_17247);
or UO_2006 (O_2006,N_18994,N_17423);
xor UO_2007 (O_2007,N_18923,N_17434);
and UO_2008 (O_2008,N_16576,N_17839);
xnor UO_2009 (O_2009,N_18667,N_19885);
nor UO_2010 (O_2010,N_17044,N_18268);
and UO_2011 (O_2011,N_16215,N_18489);
and UO_2012 (O_2012,N_17339,N_19030);
or UO_2013 (O_2013,N_19258,N_16500);
and UO_2014 (O_2014,N_19200,N_19008);
and UO_2015 (O_2015,N_19713,N_19681);
nand UO_2016 (O_2016,N_16262,N_19972);
nor UO_2017 (O_2017,N_16847,N_19769);
nor UO_2018 (O_2018,N_16788,N_18313);
or UO_2019 (O_2019,N_16196,N_17038);
nor UO_2020 (O_2020,N_18856,N_19298);
xor UO_2021 (O_2021,N_17810,N_19319);
or UO_2022 (O_2022,N_16336,N_18573);
nand UO_2023 (O_2023,N_18470,N_16419);
nor UO_2024 (O_2024,N_17427,N_19023);
nand UO_2025 (O_2025,N_17614,N_16435);
or UO_2026 (O_2026,N_18573,N_19947);
or UO_2027 (O_2027,N_16380,N_18112);
nor UO_2028 (O_2028,N_17090,N_16165);
xor UO_2029 (O_2029,N_18647,N_16223);
nor UO_2030 (O_2030,N_19292,N_17668);
nor UO_2031 (O_2031,N_17343,N_17863);
and UO_2032 (O_2032,N_16060,N_17179);
and UO_2033 (O_2033,N_18675,N_19466);
and UO_2034 (O_2034,N_19241,N_19078);
and UO_2035 (O_2035,N_17748,N_16955);
nand UO_2036 (O_2036,N_19650,N_18016);
and UO_2037 (O_2037,N_16898,N_16246);
nor UO_2038 (O_2038,N_17944,N_17426);
and UO_2039 (O_2039,N_18241,N_19053);
nor UO_2040 (O_2040,N_16304,N_16286);
and UO_2041 (O_2041,N_18036,N_18996);
nor UO_2042 (O_2042,N_18546,N_18651);
and UO_2043 (O_2043,N_17886,N_18462);
and UO_2044 (O_2044,N_17658,N_16441);
or UO_2045 (O_2045,N_16093,N_18153);
nor UO_2046 (O_2046,N_19656,N_18655);
nand UO_2047 (O_2047,N_17066,N_18559);
or UO_2048 (O_2048,N_17401,N_19737);
and UO_2049 (O_2049,N_17168,N_17345);
or UO_2050 (O_2050,N_16112,N_17115);
xor UO_2051 (O_2051,N_19389,N_19275);
and UO_2052 (O_2052,N_17635,N_17947);
xnor UO_2053 (O_2053,N_18911,N_18218);
nand UO_2054 (O_2054,N_18676,N_19919);
and UO_2055 (O_2055,N_16219,N_17609);
xor UO_2056 (O_2056,N_16432,N_17005);
nor UO_2057 (O_2057,N_17647,N_19717);
nand UO_2058 (O_2058,N_16945,N_16313);
xnor UO_2059 (O_2059,N_19182,N_19254);
xnor UO_2060 (O_2060,N_18559,N_18825);
and UO_2061 (O_2061,N_18111,N_19585);
nor UO_2062 (O_2062,N_17358,N_16181);
nor UO_2063 (O_2063,N_17756,N_18533);
and UO_2064 (O_2064,N_17299,N_16777);
xnor UO_2065 (O_2065,N_17480,N_18914);
nand UO_2066 (O_2066,N_19413,N_19906);
xor UO_2067 (O_2067,N_17711,N_17213);
and UO_2068 (O_2068,N_17352,N_17101);
nand UO_2069 (O_2069,N_18754,N_16311);
or UO_2070 (O_2070,N_16112,N_18728);
nor UO_2071 (O_2071,N_18901,N_18098);
and UO_2072 (O_2072,N_19981,N_16501);
nand UO_2073 (O_2073,N_16888,N_17578);
nor UO_2074 (O_2074,N_16480,N_19734);
nand UO_2075 (O_2075,N_17838,N_17224);
or UO_2076 (O_2076,N_18728,N_17084);
xor UO_2077 (O_2077,N_17727,N_16016);
or UO_2078 (O_2078,N_18849,N_19489);
nand UO_2079 (O_2079,N_19710,N_17834);
and UO_2080 (O_2080,N_18899,N_16609);
nand UO_2081 (O_2081,N_18438,N_17568);
xor UO_2082 (O_2082,N_19423,N_19295);
and UO_2083 (O_2083,N_17904,N_16038);
xor UO_2084 (O_2084,N_16494,N_19952);
nand UO_2085 (O_2085,N_17610,N_19368);
xor UO_2086 (O_2086,N_19340,N_16645);
and UO_2087 (O_2087,N_17281,N_16267);
nor UO_2088 (O_2088,N_18634,N_16247);
nor UO_2089 (O_2089,N_16120,N_18922);
nor UO_2090 (O_2090,N_18218,N_16226);
xnor UO_2091 (O_2091,N_18218,N_16021);
nand UO_2092 (O_2092,N_16071,N_17154);
xnor UO_2093 (O_2093,N_17183,N_19593);
and UO_2094 (O_2094,N_19769,N_18356);
or UO_2095 (O_2095,N_16855,N_16276);
and UO_2096 (O_2096,N_18707,N_19195);
nor UO_2097 (O_2097,N_18464,N_19890);
nand UO_2098 (O_2098,N_17331,N_16513);
or UO_2099 (O_2099,N_16217,N_19186);
xnor UO_2100 (O_2100,N_16389,N_16875);
nand UO_2101 (O_2101,N_18040,N_18202);
or UO_2102 (O_2102,N_19804,N_17238);
nand UO_2103 (O_2103,N_17695,N_16000);
nor UO_2104 (O_2104,N_18559,N_16639);
or UO_2105 (O_2105,N_16790,N_17280);
nor UO_2106 (O_2106,N_16515,N_18387);
nand UO_2107 (O_2107,N_17752,N_19665);
nor UO_2108 (O_2108,N_19794,N_16369);
or UO_2109 (O_2109,N_18921,N_17932);
or UO_2110 (O_2110,N_18846,N_18209);
or UO_2111 (O_2111,N_18492,N_16162);
and UO_2112 (O_2112,N_16895,N_18379);
nand UO_2113 (O_2113,N_19904,N_16807);
and UO_2114 (O_2114,N_18777,N_16056);
or UO_2115 (O_2115,N_17399,N_17806);
or UO_2116 (O_2116,N_19014,N_19350);
or UO_2117 (O_2117,N_17011,N_16517);
nand UO_2118 (O_2118,N_19073,N_18360);
or UO_2119 (O_2119,N_16605,N_16332);
or UO_2120 (O_2120,N_18641,N_19251);
nand UO_2121 (O_2121,N_16652,N_16557);
and UO_2122 (O_2122,N_18329,N_19704);
nand UO_2123 (O_2123,N_18018,N_16835);
nand UO_2124 (O_2124,N_19649,N_17251);
or UO_2125 (O_2125,N_16370,N_17231);
nor UO_2126 (O_2126,N_17496,N_19565);
or UO_2127 (O_2127,N_16812,N_19810);
nand UO_2128 (O_2128,N_17793,N_16600);
and UO_2129 (O_2129,N_18329,N_17355);
and UO_2130 (O_2130,N_17397,N_16996);
nor UO_2131 (O_2131,N_19996,N_19928);
and UO_2132 (O_2132,N_19158,N_16358);
and UO_2133 (O_2133,N_19083,N_17277);
nand UO_2134 (O_2134,N_18587,N_17972);
nand UO_2135 (O_2135,N_18177,N_17752);
or UO_2136 (O_2136,N_16444,N_18872);
nor UO_2137 (O_2137,N_19073,N_17926);
nor UO_2138 (O_2138,N_18350,N_18582);
or UO_2139 (O_2139,N_18699,N_16187);
or UO_2140 (O_2140,N_16384,N_18989);
xnor UO_2141 (O_2141,N_17897,N_19979);
and UO_2142 (O_2142,N_18669,N_19198);
xor UO_2143 (O_2143,N_16342,N_18290);
or UO_2144 (O_2144,N_18549,N_16287);
nand UO_2145 (O_2145,N_16482,N_19635);
nand UO_2146 (O_2146,N_16005,N_19760);
xor UO_2147 (O_2147,N_18885,N_18663);
nor UO_2148 (O_2148,N_17057,N_17863);
and UO_2149 (O_2149,N_16965,N_18715);
nor UO_2150 (O_2150,N_17726,N_16191);
and UO_2151 (O_2151,N_19522,N_16068);
nor UO_2152 (O_2152,N_19382,N_16661);
and UO_2153 (O_2153,N_17671,N_17447);
nand UO_2154 (O_2154,N_17813,N_16188);
xor UO_2155 (O_2155,N_19280,N_17603);
or UO_2156 (O_2156,N_17564,N_18714);
xnor UO_2157 (O_2157,N_18525,N_19314);
or UO_2158 (O_2158,N_18744,N_19379);
or UO_2159 (O_2159,N_16556,N_19694);
nor UO_2160 (O_2160,N_18288,N_16661);
xnor UO_2161 (O_2161,N_18702,N_18514);
nor UO_2162 (O_2162,N_19119,N_19688);
or UO_2163 (O_2163,N_19039,N_19404);
xor UO_2164 (O_2164,N_17505,N_16900);
xor UO_2165 (O_2165,N_18955,N_16046);
xor UO_2166 (O_2166,N_16203,N_19947);
or UO_2167 (O_2167,N_16690,N_16539);
nand UO_2168 (O_2168,N_18403,N_16073);
nor UO_2169 (O_2169,N_16956,N_16169);
xor UO_2170 (O_2170,N_19642,N_16391);
nand UO_2171 (O_2171,N_16883,N_18845);
and UO_2172 (O_2172,N_18179,N_18319);
xnor UO_2173 (O_2173,N_18070,N_18821);
nand UO_2174 (O_2174,N_16803,N_17714);
xor UO_2175 (O_2175,N_16103,N_17282);
xor UO_2176 (O_2176,N_19577,N_17862);
or UO_2177 (O_2177,N_16627,N_16024);
nor UO_2178 (O_2178,N_16851,N_18667);
and UO_2179 (O_2179,N_18473,N_17140);
nor UO_2180 (O_2180,N_17504,N_18686);
or UO_2181 (O_2181,N_16433,N_17701);
and UO_2182 (O_2182,N_17780,N_17265);
nor UO_2183 (O_2183,N_16634,N_17527);
or UO_2184 (O_2184,N_17276,N_19558);
and UO_2185 (O_2185,N_19242,N_17990);
xnor UO_2186 (O_2186,N_18169,N_17141);
nor UO_2187 (O_2187,N_18476,N_17492);
or UO_2188 (O_2188,N_16041,N_19478);
nor UO_2189 (O_2189,N_18980,N_18150);
nor UO_2190 (O_2190,N_16476,N_19790);
nor UO_2191 (O_2191,N_16367,N_19822);
xnor UO_2192 (O_2192,N_16497,N_16777);
xor UO_2193 (O_2193,N_18047,N_16683);
and UO_2194 (O_2194,N_18473,N_18124);
or UO_2195 (O_2195,N_16015,N_17787);
or UO_2196 (O_2196,N_16795,N_17076);
and UO_2197 (O_2197,N_16111,N_17558);
or UO_2198 (O_2198,N_19963,N_19574);
and UO_2199 (O_2199,N_17687,N_16762);
and UO_2200 (O_2200,N_17057,N_16346);
nand UO_2201 (O_2201,N_18163,N_18347);
and UO_2202 (O_2202,N_19639,N_18791);
or UO_2203 (O_2203,N_16083,N_19504);
nor UO_2204 (O_2204,N_17935,N_16924);
nand UO_2205 (O_2205,N_17460,N_17279);
xnor UO_2206 (O_2206,N_17000,N_16198);
xor UO_2207 (O_2207,N_17043,N_16542);
nor UO_2208 (O_2208,N_17814,N_17410);
and UO_2209 (O_2209,N_16442,N_19377);
nand UO_2210 (O_2210,N_19022,N_19668);
xnor UO_2211 (O_2211,N_16966,N_19991);
xor UO_2212 (O_2212,N_18333,N_16329);
or UO_2213 (O_2213,N_16152,N_19348);
nor UO_2214 (O_2214,N_19440,N_19509);
nand UO_2215 (O_2215,N_16527,N_17264);
nor UO_2216 (O_2216,N_19226,N_18613);
nand UO_2217 (O_2217,N_18591,N_19238);
and UO_2218 (O_2218,N_16647,N_17758);
xnor UO_2219 (O_2219,N_19060,N_19316);
xor UO_2220 (O_2220,N_19390,N_16968);
or UO_2221 (O_2221,N_19302,N_17804);
nand UO_2222 (O_2222,N_18801,N_16169);
nor UO_2223 (O_2223,N_17239,N_16362);
nor UO_2224 (O_2224,N_18981,N_16530);
nand UO_2225 (O_2225,N_18197,N_18452);
nor UO_2226 (O_2226,N_18507,N_17261);
xor UO_2227 (O_2227,N_18814,N_19500);
xor UO_2228 (O_2228,N_19303,N_18660);
nand UO_2229 (O_2229,N_18235,N_19776);
nand UO_2230 (O_2230,N_16256,N_18788);
xnor UO_2231 (O_2231,N_17145,N_17288);
or UO_2232 (O_2232,N_17289,N_17843);
xor UO_2233 (O_2233,N_19055,N_18135);
nor UO_2234 (O_2234,N_17709,N_18698);
nand UO_2235 (O_2235,N_19124,N_17732);
nand UO_2236 (O_2236,N_18099,N_18028);
and UO_2237 (O_2237,N_16255,N_19844);
nor UO_2238 (O_2238,N_17219,N_16009);
nor UO_2239 (O_2239,N_19059,N_17084);
and UO_2240 (O_2240,N_18965,N_16737);
or UO_2241 (O_2241,N_19559,N_18148);
and UO_2242 (O_2242,N_19712,N_18210);
and UO_2243 (O_2243,N_18648,N_16050);
nand UO_2244 (O_2244,N_16507,N_19211);
xor UO_2245 (O_2245,N_19013,N_16340);
nand UO_2246 (O_2246,N_17718,N_16089);
or UO_2247 (O_2247,N_17522,N_17851);
and UO_2248 (O_2248,N_16037,N_16797);
nor UO_2249 (O_2249,N_19857,N_16965);
nor UO_2250 (O_2250,N_17672,N_16552);
nor UO_2251 (O_2251,N_16328,N_18660);
nand UO_2252 (O_2252,N_16008,N_16348);
or UO_2253 (O_2253,N_18126,N_19085);
or UO_2254 (O_2254,N_18634,N_19065);
nor UO_2255 (O_2255,N_19171,N_17973);
xor UO_2256 (O_2256,N_16707,N_16426);
and UO_2257 (O_2257,N_19952,N_19043);
or UO_2258 (O_2258,N_19169,N_16041);
xor UO_2259 (O_2259,N_17377,N_19790);
nor UO_2260 (O_2260,N_16182,N_16807);
and UO_2261 (O_2261,N_18429,N_18805);
and UO_2262 (O_2262,N_18352,N_18680);
and UO_2263 (O_2263,N_17595,N_17707);
nand UO_2264 (O_2264,N_16838,N_19574);
nor UO_2265 (O_2265,N_18666,N_19506);
xor UO_2266 (O_2266,N_17030,N_19122);
xor UO_2267 (O_2267,N_19699,N_17582);
xor UO_2268 (O_2268,N_17167,N_18972);
nor UO_2269 (O_2269,N_19461,N_17253);
and UO_2270 (O_2270,N_18879,N_17349);
or UO_2271 (O_2271,N_19107,N_16086);
and UO_2272 (O_2272,N_16998,N_16959);
nand UO_2273 (O_2273,N_18957,N_18407);
and UO_2274 (O_2274,N_17053,N_16715);
or UO_2275 (O_2275,N_16277,N_17281);
nor UO_2276 (O_2276,N_16209,N_19939);
xor UO_2277 (O_2277,N_17479,N_17232);
or UO_2278 (O_2278,N_18779,N_17622);
nand UO_2279 (O_2279,N_16086,N_16631);
xnor UO_2280 (O_2280,N_18991,N_16306);
xor UO_2281 (O_2281,N_19842,N_18009);
or UO_2282 (O_2282,N_16120,N_17296);
and UO_2283 (O_2283,N_16421,N_18280);
nand UO_2284 (O_2284,N_16105,N_19619);
xnor UO_2285 (O_2285,N_16102,N_19421);
xnor UO_2286 (O_2286,N_17344,N_19750);
nand UO_2287 (O_2287,N_16502,N_17818);
nor UO_2288 (O_2288,N_17942,N_16913);
or UO_2289 (O_2289,N_17970,N_19931);
xnor UO_2290 (O_2290,N_16350,N_17361);
nor UO_2291 (O_2291,N_19759,N_16710);
nand UO_2292 (O_2292,N_16109,N_18794);
xnor UO_2293 (O_2293,N_19818,N_19302);
xor UO_2294 (O_2294,N_16625,N_16867);
and UO_2295 (O_2295,N_16555,N_18323);
nand UO_2296 (O_2296,N_16222,N_16373);
or UO_2297 (O_2297,N_16625,N_16140);
nand UO_2298 (O_2298,N_17748,N_16188);
and UO_2299 (O_2299,N_16197,N_17727);
xor UO_2300 (O_2300,N_16121,N_16716);
xor UO_2301 (O_2301,N_19663,N_19418);
xor UO_2302 (O_2302,N_19017,N_16710);
nand UO_2303 (O_2303,N_16054,N_18240);
xor UO_2304 (O_2304,N_19377,N_19429);
and UO_2305 (O_2305,N_16574,N_17090);
nand UO_2306 (O_2306,N_19470,N_17615);
or UO_2307 (O_2307,N_18604,N_19456);
nand UO_2308 (O_2308,N_18268,N_16725);
nand UO_2309 (O_2309,N_19581,N_19901);
nor UO_2310 (O_2310,N_19415,N_16711);
and UO_2311 (O_2311,N_16772,N_17696);
and UO_2312 (O_2312,N_16761,N_19744);
nand UO_2313 (O_2313,N_17619,N_17775);
or UO_2314 (O_2314,N_16942,N_17568);
xor UO_2315 (O_2315,N_18455,N_19481);
or UO_2316 (O_2316,N_16907,N_16975);
nand UO_2317 (O_2317,N_17578,N_19235);
or UO_2318 (O_2318,N_18662,N_16337);
nand UO_2319 (O_2319,N_16042,N_19265);
and UO_2320 (O_2320,N_19279,N_16103);
xnor UO_2321 (O_2321,N_17194,N_19116);
nand UO_2322 (O_2322,N_18587,N_16084);
or UO_2323 (O_2323,N_19188,N_16038);
nand UO_2324 (O_2324,N_17230,N_18643);
or UO_2325 (O_2325,N_19703,N_16984);
nor UO_2326 (O_2326,N_18767,N_18270);
xnor UO_2327 (O_2327,N_19624,N_17716);
xor UO_2328 (O_2328,N_18842,N_17895);
xnor UO_2329 (O_2329,N_19759,N_16590);
or UO_2330 (O_2330,N_16019,N_17192);
or UO_2331 (O_2331,N_16949,N_16276);
nor UO_2332 (O_2332,N_17876,N_18533);
nor UO_2333 (O_2333,N_16988,N_17533);
nand UO_2334 (O_2334,N_18971,N_17444);
and UO_2335 (O_2335,N_16784,N_18840);
nor UO_2336 (O_2336,N_18535,N_19264);
or UO_2337 (O_2337,N_18544,N_19130);
nand UO_2338 (O_2338,N_16101,N_19717);
or UO_2339 (O_2339,N_19850,N_18628);
xnor UO_2340 (O_2340,N_19583,N_17457);
or UO_2341 (O_2341,N_19258,N_16750);
nor UO_2342 (O_2342,N_16921,N_19466);
xnor UO_2343 (O_2343,N_17487,N_17569);
or UO_2344 (O_2344,N_17722,N_16779);
or UO_2345 (O_2345,N_17056,N_19828);
xor UO_2346 (O_2346,N_17959,N_19100);
nor UO_2347 (O_2347,N_16795,N_17283);
xor UO_2348 (O_2348,N_18377,N_16551);
xor UO_2349 (O_2349,N_18060,N_19658);
or UO_2350 (O_2350,N_17712,N_19605);
xor UO_2351 (O_2351,N_19446,N_16966);
or UO_2352 (O_2352,N_17290,N_18637);
nand UO_2353 (O_2353,N_16914,N_17286);
and UO_2354 (O_2354,N_17396,N_18572);
and UO_2355 (O_2355,N_16978,N_18515);
nor UO_2356 (O_2356,N_18830,N_17468);
nor UO_2357 (O_2357,N_18547,N_19547);
nand UO_2358 (O_2358,N_19658,N_18414);
and UO_2359 (O_2359,N_17743,N_16600);
nand UO_2360 (O_2360,N_18917,N_18938);
xnor UO_2361 (O_2361,N_17905,N_16930);
xnor UO_2362 (O_2362,N_19917,N_18556);
xor UO_2363 (O_2363,N_18093,N_18297);
xnor UO_2364 (O_2364,N_16796,N_19661);
xor UO_2365 (O_2365,N_16837,N_19443);
xnor UO_2366 (O_2366,N_17514,N_17768);
and UO_2367 (O_2367,N_19145,N_16932);
nand UO_2368 (O_2368,N_18063,N_19505);
nor UO_2369 (O_2369,N_16909,N_16468);
and UO_2370 (O_2370,N_19802,N_18295);
nor UO_2371 (O_2371,N_18970,N_17564);
nor UO_2372 (O_2372,N_18120,N_19681);
and UO_2373 (O_2373,N_18657,N_18106);
nor UO_2374 (O_2374,N_17263,N_16390);
and UO_2375 (O_2375,N_19224,N_17743);
nor UO_2376 (O_2376,N_18383,N_16745);
or UO_2377 (O_2377,N_16313,N_16339);
xnor UO_2378 (O_2378,N_17443,N_16669);
xor UO_2379 (O_2379,N_16992,N_19729);
nand UO_2380 (O_2380,N_17545,N_16650);
nor UO_2381 (O_2381,N_16206,N_17102);
and UO_2382 (O_2382,N_18713,N_17264);
nand UO_2383 (O_2383,N_19868,N_16970);
nor UO_2384 (O_2384,N_19332,N_18532);
nand UO_2385 (O_2385,N_16740,N_17968);
or UO_2386 (O_2386,N_19341,N_16641);
nor UO_2387 (O_2387,N_18119,N_18405);
xor UO_2388 (O_2388,N_16664,N_16014);
nor UO_2389 (O_2389,N_16785,N_18636);
nor UO_2390 (O_2390,N_18666,N_16965);
nand UO_2391 (O_2391,N_17501,N_16172);
xnor UO_2392 (O_2392,N_18058,N_18101);
or UO_2393 (O_2393,N_17896,N_18085);
or UO_2394 (O_2394,N_19858,N_18638);
nand UO_2395 (O_2395,N_19447,N_17599);
and UO_2396 (O_2396,N_16657,N_16660);
and UO_2397 (O_2397,N_17524,N_16929);
and UO_2398 (O_2398,N_16069,N_16529);
nor UO_2399 (O_2399,N_16907,N_18112);
nor UO_2400 (O_2400,N_18252,N_18317);
nor UO_2401 (O_2401,N_18718,N_18123);
nand UO_2402 (O_2402,N_16653,N_19285);
or UO_2403 (O_2403,N_18549,N_19071);
nand UO_2404 (O_2404,N_17375,N_18657);
nand UO_2405 (O_2405,N_19499,N_19817);
nor UO_2406 (O_2406,N_16101,N_17449);
and UO_2407 (O_2407,N_18585,N_16937);
and UO_2408 (O_2408,N_19479,N_19503);
nor UO_2409 (O_2409,N_16007,N_16872);
nand UO_2410 (O_2410,N_18804,N_19455);
and UO_2411 (O_2411,N_17557,N_17585);
nor UO_2412 (O_2412,N_19879,N_17536);
and UO_2413 (O_2413,N_19926,N_17629);
and UO_2414 (O_2414,N_17879,N_18744);
and UO_2415 (O_2415,N_19219,N_16444);
xnor UO_2416 (O_2416,N_16875,N_18609);
and UO_2417 (O_2417,N_19140,N_17294);
or UO_2418 (O_2418,N_18365,N_17465);
or UO_2419 (O_2419,N_19446,N_17523);
xor UO_2420 (O_2420,N_16913,N_18142);
nand UO_2421 (O_2421,N_19062,N_19161);
nor UO_2422 (O_2422,N_16969,N_17383);
and UO_2423 (O_2423,N_16136,N_17599);
nand UO_2424 (O_2424,N_19654,N_18817);
nand UO_2425 (O_2425,N_16833,N_17263);
or UO_2426 (O_2426,N_17455,N_17898);
nor UO_2427 (O_2427,N_19226,N_18516);
and UO_2428 (O_2428,N_16279,N_18683);
and UO_2429 (O_2429,N_19139,N_18456);
nand UO_2430 (O_2430,N_18088,N_19351);
xor UO_2431 (O_2431,N_19917,N_18683);
or UO_2432 (O_2432,N_17087,N_17480);
xnor UO_2433 (O_2433,N_17862,N_17559);
nand UO_2434 (O_2434,N_17444,N_19642);
and UO_2435 (O_2435,N_16198,N_17036);
and UO_2436 (O_2436,N_16512,N_18730);
xnor UO_2437 (O_2437,N_18416,N_16129);
nand UO_2438 (O_2438,N_19450,N_17495);
or UO_2439 (O_2439,N_17886,N_19617);
nor UO_2440 (O_2440,N_16269,N_17703);
xor UO_2441 (O_2441,N_16991,N_19415);
or UO_2442 (O_2442,N_16477,N_17773);
or UO_2443 (O_2443,N_17758,N_19390);
or UO_2444 (O_2444,N_19337,N_17947);
nor UO_2445 (O_2445,N_16601,N_17246);
and UO_2446 (O_2446,N_17402,N_19403);
xnor UO_2447 (O_2447,N_16248,N_18943);
nor UO_2448 (O_2448,N_17405,N_18955);
or UO_2449 (O_2449,N_16046,N_17508);
nor UO_2450 (O_2450,N_18545,N_19200);
nand UO_2451 (O_2451,N_18353,N_17517);
nor UO_2452 (O_2452,N_17795,N_19459);
xor UO_2453 (O_2453,N_16317,N_17637);
nand UO_2454 (O_2454,N_16248,N_19549);
and UO_2455 (O_2455,N_17200,N_17920);
and UO_2456 (O_2456,N_18363,N_19376);
and UO_2457 (O_2457,N_16384,N_18982);
xor UO_2458 (O_2458,N_17703,N_16748);
and UO_2459 (O_2459,N_19313,N_17025);
xnor UO_2460 (O_2460,N_18386,N_19851);
xor UO_2461 (O_2461,N_19860,N_18687);
xor UO_2462 (O_2462,N_19094,N_16708);
nor UO_2463 (O_2463,N_16627,N_19009);
and UO_2464 (O_2464,N_19468,N_19083);
nor UO_2465 (O_2465,N_16889,N_16275);
nand UO_2466 (O_2466,N_18919,N_17075);
and UO_2467 (O_2467,N_19159,N_19429);
or UO_2468 (O_2468,N_16103,N_19173);
xnor UO_2469 (O_2469,N_17768,N_18465);
nand UO_2470 (O_2470,N_16465,N_17253);
and UO_2471 (O_2471,N_18107,N_17566);
nand UO_2472 (O_2472,N_19943,N_19258);
or UO_2473 (O_2473,N_17425,N_17803);
xnor UO_2474 (O_2474,N_17695,N_19835);
nand UO_2475 (O_2475,N_17652,N_18244);
or UO_2476 (O_2476,N_18578,N_18754);
nand UO_2477 (O_2477,N_18617,N_19412);
and UO_2478 (O_2478,N_17473,N_19651);
xor UO_2479 (O_2479,N_16911,N_17646);
xor UO_2480 (O_2480,N_17704,N_17019);
nand UO_2481 (O_2481,N_17666,N_19486);
nor UO_2482 (O_2482,N_18423,N_16160);
and UO_2483 (O_2483,N_19422,N_16564);
nand UO_2484 (O_2484,N_16400,N_18287);
or UO_2485 (O_2485,N_19078,N_18000);
xor UO_2486 (O_2486,N_17387,N_19613);
or UO_2487 (O_2487,N_19646,N_17832);
nand UO_2488 (O_2488,N_18795,N_19756);
and UO_2489 (O_2489,N_17822,N_17962);
nand UO_2490 (O_2490,N_16903,N_19993);
nor UO_2491 (O_2491,N_18489,N_16880);
nor UO_2492 (O_2492,N_19796,N_19553);
or UO_2493 (O_2493,N_19307,N_18119);
nor UO_2494 (O_2494,N_16415,N_18870);
nor UO_2495 (O_2495,N_16781,N_17508);
xor UO_2496 (O_2496,N_17383,N_19001);
nor UO_2497 (O_2497,N_16612,N_16769);
xor UO_2498 (O_2498,N_18888,N_17003);
nor UO_2499 (O_2499,N_19528,N_16651);
endmodule