module basic_500_3000_500_6_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_284,In_322);
nor U1 (N_1,In_302,In_1);
nor U2 (N_2,In_312,In_62);
or U3 (N_3,In_324,In_48);
and U4 (N_4,In_201,In_78);
or U5 (N_5,In_289,In_105);
and U6 (N_6,In_444,In_80);
or U7 (N_7,In_304,In_433);
and U8 (N_8,In_151,In_251);
or U9 (N_9,In_461,In_336);
nor U10 (N_10,In_83,In_208);
nor U11 (N_11,In_497,In_197);
nand U12 (N_12,In_200,In_474);
and U13 (N_13,In_396,In_182);
and U14 (N_14,In_256,In_173);
nor U15 (N_15,In_193,In_495);
nor U16 (N_16,In_373,In_56);
nand U17 (N_17,In_181,In_153);
or U18 (N_18,In_491,In_332);
and U19 (N_19,In_8,In_81);
or U20 (N_20,In_142,In_326);
nand U21 (N_21,In_429,In_306);
or U22 (N_22,In_21,In_46);
or U23 (N_23,In_162,In_316);
or U24 (N_24,In_262,In_119);
or U25 (N_25,In_436,In_113);
or U26 (N_26,In_426,In_4);
nand U27 (N_27,In_93,In_406);
or U28 (N_28,In_325,In_219);
nor U29 (N_29,In_32,In_252);
or U30 (N_30,In_482,In_458);
and U31 (N_31,In_263,In_65);
nand U32 (N_32,In_176,In_104);
nand U33 (N_33,In_18,In_213);
nand U34 (N_34,In_390,In_337);
and U35 (N_35,In_179,In_156);
or U36 (N_36,In_449,In_67);
and U37 (N_37,In_191,In_260);
and U38 (N_38,In_146,In_335);
nor U39 (N_39,In_383,In_91);
xor U40 (N_40,In_116,In_237);
and U41 (N_41,In_283,In_69);
or U42 (N_42,In_408,In_211);
nand U43 (N_43,In_7,In_82);
and U44 (N_44,In_216,In_488);
nor U45 (N_45,In_374,In_245);
and U46 (N_46,In_346,In_441);
nand U47 (N_47,In_27,In_384);
and U48 (N_48,In_72,In_180);
nand U49 (N_49,In_25,In_432);
nand U50 (N_50,In_29,In_147);
or U51 (N_51,In_290,In_448);
nor U52 (N_52,In_218,In_363);
or U53 (N_53,In_455,In_440);
and U54 (N_54,In_372,In_349);
nor U55 (N_55,In_257,In_35);
nor U56 (N_56,In_207,In_102);
nand U57 (N_57,In_274,In_221);
and U58 (N_58,In_343,In_275);
or U59 (N_59,In_414,In_170);
nor U60 (N_60,In_97,In_84);
nor U61 (N_61,In_100,In_393);
nand U62 (N_62,In_189,In_413);
nand U63 (N_63,In_354,In_2);
nand U64 (N_64,In_468,In_492);
nor U65 (N_65,In_470,In_453);
and U66 (N_66,In_259,In_229);
and U67 (N_67,In_117,In_43);
and U68 (N_68,In_489,In_199);
nand U69 (N_69,In_339,In_136);
and U70 (N_70,In_300,In_63);
or U71 (N_71,In_228,In_165);
nor U72 (N_72,In_389,In_313);
and U73 (N_73,In_49,In_348);
nand U74 (N_74,In_244,In_490);
or U75 (N_75,In_369,In_410);
and U76 (N_76,In_96,In_273);
xor U77 (N_77,In_277,In_185);
and U78 (N_78,In_460,In_89);
nand U79 (N_79,In_291,In_194);
or U80 (N_80,In_301,In_479);
or U81 (N_81,In_196,In_51);
and U82 (N_82,In_452,In_439);
or U83 (N_83,In_230,In_403);
nand U84 (N_84,In_368,In_271);
and U85 (N_85,In_272,In_386);
nand U86 (N_86,In_344,In_109);
or U87 (N_87,In_26,In_99);
and U88 (N_88,In_480,In_421);
or U89 (N_89,In_74,In_225);
nand U90 (N_90,In_148,In_317);
xor U91 (N_91,In_129,In_445);
nand U92 (N_92,In_447,In_411);
nor U93 (N_93,In_477,In_39);
nor U94 (N_94,In_236,In_235);
and U95 (N_95,In_112,In_209);
nand U96 (N_96,In_295,In_347);
and U97 (N_97,In_476,In_184);
or U98 (N_98,In_38,In_164);
and U99 (N_99,In_50,In_15);
nand U100 (N_100,In_210,In_366);
nand U101 (N_101,In_419,In_159);
or U102 (N_102,In_94,In_279);
and U103 (N_103,In_76,In_438);
nor U104 (N_104,In_463,In_123);
nand U105 (N_105,In_103,In_364);
nand U106 (N_106,In_6,In_132);
and U107 (N_107,In_454,In_203);
and U108 (N_108,In_415,In_120);
nor U109 (N_109,In_68,In_37);
nor U110 (N_110,In_265,In_77);
or U111 (N_111,In_114,In_55);
nor U112 (N_112,In_376,In_267);
or U113 (N_113,In_446,In_166);
and U114 (N_114,In_484,In_172);
nor U115 (N_115,In_350,In_443);
or U116 (N_116,In_36,In_90);
nor U117 (N_117,In_282,In_266);
nor U118 (N_118,In_138,In_160);
or U119 (N_119,In_281,In_293);
nor U120 (N_120,In_107,In_308);
or U121 (N_121,In_155,In_286);
nor U122 (N_122,In_143,In_169);
or U123 (N_123,In_47,In_395);
and U124 (N_124,In_59,In_355);
and U125 (N_125,In_190,In_467);
and U126 (N_126,In_42,In_122);
nand U127 (N_127,In_417,In_303);
nor U128 (N_128,In_360,In_177);
nand U129 (N_129,In_405,In_334);
xnor U130 (N_130,In_398,In_288);
nand U131 (N_131,In_400,In_434);
or U132 (N_132,In_330,In_328);
and U133 (N_133,In_247,In_478);
or U134 (N_134,In_380,In_214);
or U135 (N_135,In_377,In_361);
nand U136 (N_136,In_168,In_111);
nand U137 (N_137,In_115,In_431);
nor U138 (N_138,In_250,In_135);
or U139 (N_139,In_345,In_154);
nor U140 (N_140,In_375,In_342);
or U141 (N_141,In_422,In_269);
nor U142 (N_142,In_285,In_456);
and U143 (N_143,In_9,In_58);
nand U144 (N_144,In_459,In_133);
or U145 (N_145,In_401,In_382);
or U146 (N_146,In_53,In_430);
and U147 (N_147,In_493,In_70);
nor U148 (N_148,In_409,In_23);
and U149 (N_149,In_246,In_110);
and U150 (N_150,In_486,In_305);
and U151 (N_151,In_424,In_223);
or U152 (N_152,In_367,In_362);
and U153 (N_153,In_243,In_121);
nor U154 (N_154,In_356,In_278);
or U155 (N_155,In_387,In_254);
nor U156 (N_156,In_397,In_158);
nor U157 (N_157,In_351,In_268);
and U158 (N_158,In_315,In_297);
or U159 (N_159,In_30,In_457);
nand U160 (N_160,In_473,In_124);
and U161 (N_161,In_204,In_388);
nand U162 (N_162,In_258,In_311);
or U163 (N_163,In_494,In_44);
nand U164 (N_164,In_139,In_248);
nand U165 (N_165,In_292,In_242);
and U166 (N_166,In_137,In_427);
nand U167 (N_167,In_41,In_496);
nand U168 (N_168,In_358,In_296);
nand U169 (N_169,In_323,In_222);
nor U170 (N_170,In_5,In_101);
nand U171 (N_171,In_391,In_60);
or U172 (N_172,In_270,In_378);
and U173 (N_173,In_294,In_309);
and U174 (N_174,In_195,In_220);
nor U175 (N_175,In_130,In_416);
or U176 (N_176,In_359,In_92);
or U177 (N_177,In_118,In_475);
or U178 (N_178,In_321,In_174);
or U179 (N_179,In_412,In_353);
nand U180 (N_180,In_498,In_319);
or U181 (N_181,In_287,In_171);
nand U182 (N_182,In_418,In_483);
and U183 (N_183,In_52,In_75);
and U184 (N_184,In_188,In_98);
and U185 (N_185,In_141,In_227);
nand U186 (N_186,In_144,In_34);
nor U187 (N_187,In_404,In_134);
nand U188 (N_188,In_333,In_442);
or U189 (N_189,In_87,In_365);
and U190 (N_190,In_66,In_239);
or U191 (N_191,In_464,In_255);
nand U192 (N_192,In_140,In_276);
and U193 (N_193,In_95,In_178);
nand U194 (N_194,In_61,In_234);
or U195 (N_195,In_340,In_40);
or U196 (N_196,In_17,In_423);
nor U197 (N_197,In_24,In_152);
and U198 (N_198,In_299,In_20);
and U199 (N_199,In_261,In_450);
or U200 (N_200,In_85,In_469);
nor U201 (N_201,In_217,In_79);
nand U202 (N_202,In_462,In_466);
or U203 (N_203,In_331,In_127);
nand U204 (N_204,In_370,In_86);
nor U205 (N_205,In_205,In_371);
or U206 (N_206,In_108,In_33);
nor U207 (N_207,In_232,In_88);
or U208 (N_208,In_149,In_341);
nor U209 (N_209,In_318,In_338);
nor U210 (N_210,In_145,In_314);
or U211 (N_211,In_379,In_13);
and U212 (N_212,In_249,In_264);
or U213 (N_213,In_215,In_16);
nor U214 (N_214,In_186,In_435);
nand U215 (N_215,In_106,In_150);
nor U216 (N_216,In_402,In_240);
or U217 (N_217,In_329,In_54);
and U218 (N_218,In_212,In_224);
nand U219 (N_219,In_472,In_22);
and U220 (N_220,In_11,In_451);
and U221 (N_221,In_357,In_28);
and U222 (N_222,In_485,In_428);
and U223 (N_223,In_226,In_128);
nand U224 (N_224,In_407,In_381);
and U225 (N_225,In_481,In_198);
or U226 (N_226,In_10,In_420);
or U227 (N_227,In_183,In_392);
nor U228 (N_228,In_399,In_167);
or U229 (N_229,In_231,In_64);
nand U230 (N_230,In_19,In_12);
and U231 (N_231,In_425,In_487);
nor U232 (N_232,In_0,In_73);
or U233 (N_233,In_163,In_280);
and U234 (N_234,In_202,In_192);
nor U235 (N_235,In_465,In_157);
nand U236 (N_236,In_57,In_125);
nand U237 (N_237,In_3,In_327);
nand U238 (N_238,In_307,In_126);
nor U239 (N_239,In_499,In_161);
or U240 (N_240,In_71,In_385);
or U241 (N_241,In_320,In_298);
and U242 (N_242,In_241,In_14);
and U243 (N_243,In_394,In_437);
and U244 (N_244,In_131,In_45);
or U245 (N_245,In_187,In_310);
and U246 (N_246,In_206,In_233);
and U247 (N_247,In_238,In_471);
and U248 (N_248,In_352,In_175);
nor U249 (N_249,In_253,In_31);
nor U250 (N_250,In_230,In_489);
nand U251 (N_251,In_383,In_32);
or U252 (N_252,In_429,In_296);
or U253 (N_253,In_5,In_15);
nand U254 (N_254,In_191,In_214);
and U255 (N_255,In_203,In_467);
nor U256 (N_256,In_450,In_158);
nor U257 (N_257,In_99,In_33);
and U258 (N_258,In_236,In_209);
nor U259 (N_259,In_195,In_129);
or U260 (N_260,In_197,In_464);
nor U261 (N_261,In_489,In_265);
or U262 (N_262,In_176,In_292);
nand U263 (N_263,In_238,In_245);
nand U264 (N_264,In_113,In_444);
xor U265 (N_265,In_91,In_9);
and U266 (N_266,In_99,In_455);
or U267 (N_267,In_198,In_86);
and U268 (N_268,In_340,In_287);
nand U269 (N_269,In_177,In_242);
or U270 (N_270,In_486,In_288);
nand U271 (N_271,In_334,In_218);
and U272 (N_272,In_115,In_355);
and U273 (N_273,In_113,In_36);
or U274 (N_274,In_321,In_453);
nand U275 (N_275,In_59,In_230);
or U276 (N_276,In_89,In_476);
nand U277 (N_277,In_492,In_267);
and U278 (N_278,In_8,In_144);
or U279 (N_279,In_140,In_128);
or U280 (N_280,In_134,In_33);
nand U281 (N_281,In_472,In_323);
and U282 (N_282,In_326,In_455);
or U283 (N_283,In_228,In_93);
nand U284 (N_284,In_422,In_322);
or U285 (N_285,In_188,In_145);
xnor U286 (N_286,In_297,In_461);
nand U287 (N_287,In_404,In_403);
nand U288 (N_288,In_4,In_375);
or U289 (N_289,In_6,In_172);
nor U290 (N_290,In_393,In_327);
nor U291 (N_291,In_59,In_199);
nand U292 (N_292,In_36,In_55);
nand U293 (N_293,In_245,In_265);
and U294 (N_294,In_40,In_347);
nor U295 (N_295,In_135,In_110);
nor U296 (N_296,In_160,In_265);
or U297 (N_297,In_33,In_468);
or U298 (N_298,In_251,In_17);
or U299 (N_299,In_350,In_1);
nor U300 (N_300,In_42,In_22);
nor U301 (N_301,In_167,In_321);
nor U302 (N_302,In_283,In_98);
nand U303 (N_303,In_199,In_383);
and U304 (N_304,In_268,In_110);
and U305 (N_305,In_357,In_20);
nor U306 (N_306,In_312,In_303);
nor U307 (N_307,In_301,In_359);
or U308 (N_308,In_475,In_364);
or U309 (N_309,In_353,In_452);
nor U310 (N_310,In_490,In_411);
and U311 (N_311,In_196,In_339);
nor U312 (N_312,In_230,In_211);
nand U313 (N_313,In_109,In_343);
nor U314 (N_314,In_132,In_287);
nor U315 (N_315,In_109,In_54);
nor U316 (N_316,In_440,In_83);
and U317 (N_317,In_301,In_173);
or U318 (N_318,In_180,In_349);
and U319 (N_319,In_74,In_354);
and U320 (N_320,In_72,In_253);
or U321 (N_321,In_131,In_333);
and U322 (N_322,In_366,In_478);
nand U323 (N_323,In_463,In_475);
nor U324 (N_324,In_278,In_466);
nor U325 (N_325,In_171,In_407);
xnor U326 (N_326,In_467,In_181);
nor U327 (N_327,In_427,In_389);
nand U328 (N_328,In_484,In_87);
or U329 (N_329,In_237,In_6);
nor U330 (N_330,In_434,In_6);
and U331 (N_331,In_248,In_311);
nor U332 (N_332,In_299,In_449);
and U333 (N_333,In_337,In_420);
nand U334 (N_334,In_129,In_96);
and U335 (N_335,In_168,In_374);
and U336 (N_336,In_212,In_257);
or U337 (N_337,In_26,In_426);
nand U338 (N_338,In_166,In_45);
nor U339 (N_339,In_100,In_200);
or U340 (N_340,In_33,In_0);
nor U341 (N_341,In_32,In_203);
nor U342 (N_342,In_432,In_413);
nand U343 (N_343,In_392,In_472);
nand U344 (N_344,In_33,In_314);
and U345 (N_345,In_223,In_267);
nand U346 (N_346,In_237,In_409);
nor U347 (N_347,In_479,In_135);
nor U348 (N_348,In_17,In_30);
nor U349 (N_349,In_135,In_326);
or U350 (N_350,In_56,In_463);
nand U351 (N_351,In_138,In_227);
nor U352 (N_352,In_471,In_159);
or U353 (N_353,In_183,In_486);
nand U354 (N_354,In_267,In_179);
and U355 (N_355,In_225,In_86);
or U356 (N_356,In_347,In_47);
nand U357 (N_357,In_88,In_473);
nor U358 (N_358,In_68,In_85);
nor U359 (N_359,In_206,In_404);
nand U360 (N_360,In_242,In_213);
nor U361 (N_361,In_322,In_15);
nand U362 (N_362,In_119,In_334);
or U363 (N_363,In_236,In_170);
nor U364 (N_364,In_435,In_441);
or U365 (N_365,In_449,In_446);
nor U366 (N_366,In_432,In_47);
xnor U367 (N_367,In_469,In_336);
and U368 (N_368,In_440,In_287);
nand U369 (N_369,In_493,In_18);
and U370 (N_370,In_234,In_490);
nand U371 (N_371,In_142,In_288);
or U372 (N_372,In_303,In_468);
xor U373 (N_373,In_159,In_413);
xnor U374 (N_374,In_67,In_140);
or U375 (N_375,In_90,In_389);
and U376 (N_376,In_443,In_160);
nand U377 (N_377,In_9,In_279);
and U378 (N_378,In_423,In_78);
or U379 (N_379,In_75,In_274);
nand U380 (N_380,In_446,In_383);
and U381 (N_381,In_368,In_334);
and U382 (N_382,In_92,In_440);
nor U383 (N_383,In_367,In_377);
and U384 (N_384,In_69,In_66);
or U385 (N_385,In_291,In_292);
nor U386 (N_386,In_322,In_153);
and U387 (N_387,In_373,In_191);
and U388 (N_388,In_210,In_190);
or U389 (N_389,In_69,In_250);
or U390 (N_390,In_350,In_447);
nor U391 (N_391,In_237,In_179);
xnor U392 (N_392,In_142,In_322);
nand U393 (N_393,In_266,In_482);
or U394 (N_394,In_75,In_293);
or U395 (N_395,In_118,In_380);
and U396 (N_396,In_91,In_12);
nand U397 (N_397,In_256,In_35);
and U398 (N_398,In_151,In_450);
nor U399 (N_399,In_257,In_113);
or U400 (N_400,In_367,In_190);
nand U401 (N_401,In_96,In_265);
or U402 (N_402,In_246,In_127);
nand U403 (N_403,In_111,In_335);
nor U404 (N_404,In_397,In_43);
and U405 (N_405,In_270,In_66);
and U406 (N_406,In_195,In_384);
or U407 (N_407,In_247,In_458);
nor U408 (N_408,In_3,In_356);
xor U409 (N_409,In_147,In_11);
nand U410 (N_410,In_252,In_381);
and U411 (N_411,In_396,In_244);
nor U412 (N_412,In_236,In_328);
nor U413 (N_413,In_51,In_82);
nand U414 (N_414,In_470,In_311);
and U415 (N_415,In_445,In_193);
and U416 (N_416,In_311,In_203);
or U417 (N_417,In_318,In_273);
nand U418 (N_418,In_236,In_26);
and U419 (N_419,In_429,In_240);
or U420 (N_420,In_390,In_449);
or U421 (N_421,In_413,In_214);
nor U422 (N_422,In_346,In_67);
nor U423 (N_423,In_17,In_405);
nor U424 (N_424,In_350,In_259);
nor U425 (N_425,In_1,In_98);
and U426 (N_426,In_489,In_469);
nand U427 (N_427,In_329,In_278);
or U428 (N_428,In_229,In_224);
and U429 (N_429,In_410,In_104);
or U430 (N_430,In_463,In_312);
nor U431 (N_431,In_108,In_134);
and U432 (N_432,In_469,In_196);
and U433 (N_433,In_333,In_499);
and U434 (N_434,In_31,In_9);
or U435 (N_435,In_237,In_23);
nor U436 (N_436,In_446,In_108);
and U437 (N_437,In_234,In_137);
and U438 (N_438,In_7,In_358);
nor U439 (N_439,In_159,In_395);
nor U440 (N_440,In_255,In_417);
or U441 (N_441,In_467,In_32);
or U442 (N_442,In_424,In_405);
nor U443 (N_443,In_212,In_474);
or U444 (N_444,In_94,In_73);
xor U445 (N_445,In_301,In_369);
and U446 (N_446,In_361,In_44);
nor U447 (N_447,In_392,In_84);
or U448 (N_448,In_214,In_5);
and U449 (N_449,In_42,In_332);
and U450 (N_450,In_43,In_300);
nor U451 (N_451,In_335,In_327);
and U452 (N_452,In_459,In_328);
or U453 (N_453,In_120,In_222);
nand U454 (N_454,In_196,In_55);
nand U455 (N_455,In_235,In_87);
and U456 (N_456,In_381,In_244);
or U457 (N_457,In_378,In_233);
and U458 (N_458,In_20,In_154);
or U459 (N_459,In_461,In_323);
or U460 (N_460,In_372,In_193);
or U461 (N_461,In_174,In_180);
nor U462 (N_462,In_243,In_447);
and U463 (N_463,In_383,In_46);
nand U464 (N_464,In_8,In_429);
nand U465 (N_465,In_250,In_454);
nor U466 (N_466,In_345,In_363);
nor U467 (N_467,In_215,In_170);
or U468 (N_468,In_91,In_59);
nand U469 (N_469,In_323,In_57);
nor U470 (N_470,In_61,In_481);
nor U471 (N_471,In_243,In_175);
nand U472 (N_472,In_153,In_257);
or U473 (N_473,In_450,In_123);
nor U474 (N_474,In_100,In_361);
nor U475 (N_475,In_391,In_170);
and U476 (N_476,In_360,In_141);
and U477 (N_477,In_182,In_282);
or U478 (N_478,In_443,In_138);
or U479 (N_479,In_130,In_442);
or U480 (N_480,In_31,In_137);
nand U481 (N_481,In_92,In_83);
nor U482 (N_482,In_210,In_108);
and U483 (N_483,In_390,In_190);
and U484 (N_484,In_245,In_0);
and U485 (N_485,In_263,In_89);
nand U486 (N_486,In_330,In_50);
nand U487 (N_487,In_277,In_19);
or U488 (N_488,In_48,In_208);
or U489 (N_489,In_59,In_362);
nor U490 (N_490,In_112,In_454);
or U491 (N_491,In_469,In_125);
and U492 (N_492,In_455,In_100);
or U493 (N_493,In_223,In_169);
or U494 (N_494,In_353,In_381);
nand U495 (N_495,In_200,In_377);
and U496 (N_496,In_207,In_275);
and U497 (N_497,In_268,In_109);
and U498 (N_498,In_170,In_73);
nand U499 (N_499,In_368,In_195);
and U500 (N_500,N_184,N_303);
nand U501 (N_501,N_387,N_337);
and U502 (N_502,N_438,N_401);
nor U503 (N_503,N_79,N_412);
and U504 (N_504,N_213,N_4);
nand U505 (N_505,N_437,N_279);
nor U506 (N_506,N_222,N_317);
nor U507 (N_507,N_174,N_59);
or U508 (N_508,N_262,N_381);
or U509 (N_509,N_442,N_443);
or U510 (N_510,N_81,N_444);
or U511 (N_511,N_390,N_340);
nor U512 (N_512,N_54,N_382);
or U513 (N_513,N_7,N_467);
and U514 (N_514,N_158,N_487);
or U515 (N_515,N_452,N_197);
and U516 (N_516,N_426,N_259);
nand U517 (N_517,N_394,N_298);
nor U518 (N_518,N_205,N_207);
and U519 (N_519,N_44,N_344);
nor U520 (N_520,N_245,N_406);
nor U521 (N_521,N_86,N_297);
xnor U522 (N_522,N_481,N_186);
or U523 (N_523,N_52,N_29);
nand U524 (N_524,N_399,N_459);
and U525 (N_525,N_348,N_370);
nor U526 (N_526,N_121,N_127);
nor U527 (N_527,N_314,N_351);
and U528 (N_528,N_172,N_322);
nand U529 (N_529,N_103,N_447);
nor U530 (N_530,N_239,N_100);
nor U531 (N_531,N_469,N_91);
nor U532 (N_532,N_28,N_154);
and U533 (N_533,N_66,N_236);
and U534 (N_534,N_138,N_369);
nor U535 (N_535,N_450,N_41);
nor U536 (N_536,N_34,N_335);
nand U537 (N_537,N_339,N_324);
or U538 (N_538,N_408,N_313);
nand U539 (N_539,N_157,N_198);
or U540 (N_540,N_88,N_456);
or U541 (N_541,N_376,N_55);
and U542 (N_542,N_393,N_130);
nor U543 (N_543,N_446,N_72);
and U544 (N_544,N_219,N_22);
or U545 (N_545,N_416,N_389);
nor U546 (N_546,N_73,N_92);
nand U547 (N_547,N_232,N_187);
or U548 (N_548,N_165,N_206);
and U549 (N_549,N_252,N_74);
nand U550 (N_550,N_167,N_392);
nand U551 (N_551,N_129,N_256);
and U552 (N_552,N_257,N_250);
and U553 (N_553,N_425,N_168);
or U554 (N_554,N_478,N_46);
and U555 (N_555,N_361,N_420);
or U556 (N_556,N_462,N_153);
or U557 (N_557,N_355,N_491);
nand U558 (N_558,N_273,N_366);
and U559 (N_559,N_359,N_451);
nand U560 (N_560,N_325,N_440);
and U561 (N_561,N_377,N_396);
nand U562 (N_562,N_276,N_435);
nor U563 (N_563,N_208,N_38);
and U564 (N_564,N_490,N_260);
or U565 (N_565,N_78,N_196);
and U566 (N_566,N_71,N_163);
nand U567 (N_567,N_221,N_357);
nor U568 (N_568,N_16,N_371);
or U569 (N_569,N_421,N_118);
nand U570 (N_570,N_114,N_286);
nand U571 (N_571,N_83,N_5);
xnor U572 (N_572,N_87,N_281);
and U573 (N_573,N_65,N_191);
or U574 (N_574,N_306,N_115);
nor U575 (N_575,N_363,N_234);
nor U576 (N_576,N_480,N_282);
or U577 (N_577,N_228,N_182);
and U578 (N_578,N_328,N_265);
nor U579 (N_579,N_270,N_296);
or U580 (N_580,N_316,N_64);
nor U581 (N_581,N_75,N_455);
nor U582 (N_582,N_27,N_101);
nor U583 (N_583,N_152,N_11);
nor U584 (N_584,N_51,N_58);
nand U585 (N_585,N_235,N_460);
nor U586 (N_586,N_274,N_39);
and U587 (N_587,N_224,N_20);
nand U588 (N_588,N_427,N_227);
and U589 (N_589,N_246,N_135);
and U590 (N_590,N_485,N_69);
or U591 (N_591,N_334,N_36);
nor U592 (N_592,N_181,N_431);
or U593 (N_593,N_284,N_60);
nand U594 (N_594,N_63,N_278);
or U595 (N_595,N_295,N_68);
or U596 (N_596,N_343,N_411);
nor U597 (N_597,N_386,N_137);
nand U598 (N_598,N_277,N_307);
nor U599 (N_599,N_145,N_470);
nor U600 (N_600,N_77,N_150);
nand U601 (N_601,N_151,N_179);
or U602 (N_602,N_241,N_433);
nand U603 (N_603,N_409,N_49);
or U604 (N_604,N_464,N_323);
and U605 (N_605,N_413,N_423);
nand U606 (N_606,N_410,N_358);
nor U607 (N_607,N_12,N_280);
nor U608 (N_608,N_251,N_458);
nand U609 (N_609,N_300,N_327);
nor U610 (N_610,N_0,N_243);
or U611 (N_611,N_275,N_312);
and U612 (N_612,N_217,N_18);
and U613 (N_613,N_108,N_321);
nor U614 (N_614,N_190,N_488);
nor U615 (N_615,N_90,N_407);
nor U616 (N_616,N_67,N_373);
nor U617 (N_617,N_98,N_10);
and U618 (N_618,N_449,N_202);
nand U619 (N_619,N_489,N_220);
nand U620 (N_620,N_117,N_47);
nand U621 (N_621,N_105,N_486);
nand U622 (N_622,N_112,N_258);
and U623 (N_623,N_175,N_80);
nor U624 (N_624,N_212,N_56);
nor U625 (N_625,N_99,N_237);
nand U626 (N_626,N_136,N_177);
or U627 (N_627,N_9,N_148);
nand U628 (N_628,N_21,N_388);
and U629 (N_629,N_364,N_139);
nand U630 (N_630,N_436,N_285);
nand U631 (N_631,N_31,N_82);
or U632 (N_632,N_331,N_292);
nor U633 (N_633,N_493,N_418);
nand U634 (N_634,N_497,N_261);
xor U635 (N_635,N_482,N_463);
nand U636 (N_636,N_404,N_301);
nor U637 (N_637,N_379,N_122);
nand U638 (N_638,N_330,N_125);
nor U639 (N_639,N_32,N_253);
or U640 (N_640,N_142,N_332);
and U641 (N_641,N_329,N_25);
nand U642 (N_642,N_374,N_162);
nor U643 (N_643,N_14,N_468);
and U644 (N_644,N_33,N_304);
nand U645 (N_645,N_144,N_395);
nand U646 (N_646,N_180,N_320);
or U647 (N_647,N_171,N_448);
nor U648 (N_648,N_155,N_305);
nor U649 (N_649,N_384,N_288);
or U650 (N_650,N_141,N_318);
nor U651 (N_651,N_495,N_203);
nor U652 (N_652,N_476,N_309);
and U653 (N_653,N_211,N_453);
and U654 (N_654,N_432,N_95);
nand U655 (N_655,N_445,N_417);
or U656 (N_656,N_209,N_93);
nand U657 (N_657,N_166,N_465);
or U658 (N_658,N_400,N_26);
or U659 (N_659,N_248,N_161);
and U660 (N_660,N_147,N_160);
or U661 (N_661,N_70,N_457);
nand U662 (N_662,N_189,N_113);
nor U663 (N_663,N_454,N_254);
and U664 (N_664,N_310,N_414);
nor U665 (N_665,N_383,N_53);
or U666 (N_666,N_378,N_146);
or U667 (N_667,N_474,N_345);
and U668 (N_668,N_424,N_120);
or U669 (N_669,N_173,N_192);
and U670 (N_670,N_104,N_471);
nand U671 (N_671,N_422,N_473);
nor U672 (N_672,N_164,N_45);
or U673 (N_673,N_218,N_362);
or U674 (N_674,N_178,N_268);
or U675 (N_675,N_472,N_42);
and U676 (N_676,N_240,N_35);
and U677 (N_677,N_6,N_143);
and U678 (N_678,N_415,N_183);
nand U679 (N_679,N_391,N_402);
or U680 (N_680,N_499,N_483);
nand U681 (N_681,N_293,N_365);
nor U682 (N_682,N_159,N_116);
and U683 (N_683,N_111,N_349);
and U684 (N_684,N_484,N_333);
nor U685 (N_685,N_124,N_57);
nor U686 (N_686,N_375,N_403);
or U687 (N_687,N_283,N_397);
or U688 (N_688,N_347,N_419);
nor U689 (N_689,N_350,N_62);
nor U690 (N_690,N_194,N_249);
or U691 (N_691,N_479,N_214);
or U692 (N_692,N_24,N_441);
nor U693 (N_693,N_199,N_244);
and U694 (N_694,N_15,N_185);
nor U695 (N_695,N_200,N_430);
nand U696 (N_696,N_40,N_354);
and U697 (N_697,N_193,N_494);
or U698 (N_698,N_43,N_215);
or U699 (N_699,N_128,N_315);
and U700 (N_700,N_216,N_231);
nand U701 (N_701,N_272,N_169);
and U702 (N_702,N_461,N_311);
nor U703 (N_703,N_294,N_356);
nand U704 (N_704,N_84,N_2);
nand U705 (N_705,N_308,N_102);
or U706 (N_706,N_291,N_367);
nand U707 (N_707,N_8,N_1);
or U708 (N_708,N_201,N_156);
nand U709 (N_709,N_110,N_97);
nand U710 (N_710,N_223,N_23);
nor U711 (N_711,N_229,N_385);
nor U712 (N_712,N_123,N_233);
nand U713 (N_713,N_204,N_346);
nand U714 (N_714,N_492,N_17);
nor U715 (N_715,N_50,N_299);
nand U716 (N_716,N_271,N_302);
or U717 (N_717,N_360,N_372);
nor U718 (N_718,N_13,N_368);
and U719 (N_719,N_405,N_30);
or U720 (N_720,N_149,N_319);
or U721 (N_721,N_255,N_131);
and U722 (N_722,N_225,N_267);
nor U723 (N_723,N_434,N_61);
nand U724 (N_724,N_76,N_429);
nand U725 (N_725,N_380,N_269);
nand U726 (N_726,N_287,N_85);
nor U727 (N_727,N_289,N_290);
or U728 (N_728,N_195,N_496);
and U729 (N_729,N_3,N_107);
nand U730 (N_730,N_230,N_352);
nand U731 (N_731,N_19,N_48);
and U732 (N_732,N_338,N_475);
and U733 (N_733,N_353,N_176);
nand U734 (N_734,N_226,N_188);
and U735 (N_735,N_133,N_498);
nor U736 (N_736,N_170,N_398);
nand U737 (N_737,N_238,N_106);
nor U738 (N_738,N_326,N_242);
nand U739 (N_739,N_264,N_263);
or U740 (N_740,N_342,N_134);
or U741 (N_741,N_94,N_266);
or U742 (N_742,N_37,N_466);
or U743 (N_743,N_247,N_140);
nand U744 (N_744,N_439,N_132);
or U745 (N_745,N_119,N_428);
nand U746 (N_746,N_89,N_96);
and U747 (N_747,N_477,N_126);
nor U748 (N_748,N_109,N_341);
and U749 (N_749,N_210,N_336);
nor U750 (N_750,N_65,N_50);
and U751 (N_751,N_123,N_193);
or U752 (N_752,N_46,N_174);
nor U753 (N_753,N_323,N_252);
or U754 (N_754,N_218,N_484);
nand U755 (N_755,N_22,N_322);
nor U756 (N_756,N_147,N_176);
nand U757 (N_757,N_455,N_405);
nor U758 (N_758,N_413,N_215);
and U759 (N_759,N_396,N_129);
and U760 (N_760,N_320,N_294);
or U761 (N_761,N_253,N_422);
nor U762 (N_762,N_25,N_176);
and U763 (N_763,N_160,N_300);
and U764 (N_764,N_44,N_478);
or U765 (N_765,N_333,N_144);
nor U766 (N_766,N_307,N_70);
and U767 (N_767,N_216,N_311);
or U768 (N_768,N_481,N_310);
and U769 (N_769,N_116,N_420);
nand U770 (N_770,N_371,N_144);
and U771 (N_771,N_72,N_113);
nand U772 (N_772,N_391,N_182);
or U773 (N_773,N_307,N_25);
nand U774 (N_774,N_213,N_41);
or U775 (N_775,N_230,N_390);
or U776 (N_776,N_307,N_49);
and U777 (N_777,N_382,N_292);
or U778 (N_778,N_338,N_3);
nor U779 (N_779,N_273,N_402);
nor U780 (N_780,N_412,N_473);
or U781 (N_781,N_237,N_102);
nand U782 (N_782,N_467,N_304);
or U783 (N_783,N_3,N_329);
nor U784 (N_784,N_188,N_259);
and U785 (N_785,N_161,N_317);
nand U786 (N_786,N_258,N_159);
xnor U787 (N_787,N_185,N_444);
nor U788 (N_788,N_475,N_17);
nand U789 (N_789,N_150,N_234);
and U790 (N_790,N_267,N_200);
and U791 (N_791,N_67,N_233);
nor U792 (N_792,N_432,N_67);
nor U793 (N_793,N_121,N_237);
and U794 (N_794,N_455,N_428);
and U795 (N_795,N_89,N_314);
or U796 (N_796,N_164,N_361);
or U797 (N_797,N_45,N_312);
or U798 (N_798,N_76,N_328);
or U799 (N_799,N_464,N_49);
or U800 (N_800,N_80,N_42);
and U801 (N_801,N_124,N_427);
or U802 (N_802,N_353,N_412);
nor U803 (N_803,N_194,N_153);
nand U804 (N_804,N_110,N_19);
and U805 (N_805,N_472,N_427);
or U806 (N_806,N_55,N_175);
or U807 (N_807,N_290,N_325);
or U808 (N_808,N_17,N_348);
or U809 (N_809,N_12,N_134);
nor U810 (N_810,N_129,N_451);
xor U811 (N_811,N_63,N_292);
nand U812 (N_812,N_18,N_210);
nand U813 (N_813,N_20,N_284);
or U814 (N_814,N_38,N_489);
nand U815 (N_815,N_230,N_233);
or U816 (N_816,N_446,N_226);
and U817 (N_817,N_242,N_132);
xor U818 (N_818,N_246,N_440);
xnor U819 (N_819,N_30,N_289);
or U820 (N_820,N_351,N_1);
and U821 (N_821,N_301,N_497);
nor U822 (N_822,N_27,N_453);
nand U823 (N_823,N_115,N_6);
nand U824 (N_824,N_449,N_290);
nor U825 (N_825,N_275,N_429);
nor U826 (N_826,N_197,N_158);
and U827 (N_827,N_297,N_212);
nor U828 (N_828,N_149,N_82);
and U829 (N_829,N_228,N_399);
and U830 (N_830,N_484,N_277);
and U831 (N_831,N_308,N_137);
nand U832 (N_832,N_481,N_456);
nor U833 (N_833,N_110,N_78);
nand U834 (N_834,N_326,N_475);
or U835 (N_835,N_91,N_383);
xnor U836 (N_836,N_89,N_193);
and U837 (N_837,N_334,N_303);
or U838 (N_838,N_45,N_176);
nor U839 (N_839,N_368,N_459);
nand U840 (N_840,N_13,N_149);
nand U841 (N_841,N_23,N_124);
xnor U842 (N_842,N_420,N_61);
and U843 (N_843,N_377,N_78);
or U844 (N_844,N_324,N_100);
nor U845 (N_845,N_275,N_359);
and U846 (N_846,N_223,N_55);
xor U847 (N_847,N_354,N_148);
or U848 (N_848,N_101,N_240);
nand U849 (N_849,N_394,N_117);
and U850 (N_850,N_401,N_183);
nand U851 (N_851,N_144,N_56);
or U852 (N_852,N_463,N_159);
nand U853 (N_853,N_111,N_73);
nor U854 (N_854,N_211,N_459);
and U855 (N_855,N_27,N_395);
nor U856 (N_856,N_370,N_158);
nand U857 (N_857,N_212,N_100);
or U858 (N_858,N_329,N_418);
and U859 (N_859,N_157,N_163);
or U860 (N_860,N_179,N_221);
and U861 (N_861,N_10,N_207);
nor U862 (N_862,N_257,N_144);
nor U863 (N_863,N_383,N_371);
and U864 (N_864,N_86,N_307);
nor U865 (N_865,N_497,N_169);
and U866 (N_866,N_499,N_328);
nand U867 (N_867,N_196,N_289);
nand U868 (N_868,N_478,N_139);
nor U869 (N_869,N_290,N_151);
nor U870 (N_870,N_279,N_460);
and U871 (N_871,N_415,N_434);
and U872 (N_872,N_68,N_27);
or U873 (N_873,N_262,N_131);
nor U874 (N_874,N_298,N_88);
or U875 (N_875,N_364,N_231);
nand U876 (N_876,N_464,N_2);
or U877 (N_877,N_218,N_465);
nor U878 (N_878,N_493,N_297);
or U879 (N_879,N_412,N_133);
and U880 (N_880,N_51,N_116);
or U881 (N_881,N_309,N_78);
or U882 (N_882,N_376,N_259);
nor U883 (N_883,N_125,N_395);
or U884 (N_884,N_309,N_163);
and U885 (N_885,N_331,N_169);
or U886 (N_886,N_408,N_255);
nor U887 (N_887,N_415,N_55);
and U888 (N_888,N_222,N_298);
or U889 (N_889,N_295,N_48);
and U890 (N_890,N_386,N_499);
nor U891 (N_891,N_438,N_395);
or U892 (N_892,N_337,N_406);
and U893 (N_893,N_206,N_37);
or U894 (N_894,N_418,N_52);
nor U895 (N_895,N_289,N_142);
nand U896 (N_896,N_102,N_202);
nand U897 (N_897,N_479,N_488);
or U898 (N_898,N_235,N_108);
or U899 (N_899,N_303,N_146);
nor U900 (N_900,N_398,N_100);
or U901 (N_901,N_65,N_199);
nor U902 (N_902,N_229,N_164);
nand U903 (N_903,N_11,N_238);
nand U904 (N_904,N_264,N_237);
or U905 (N_905,N_437,N_18);
nor U906 (N_906,N_196,N_473);
and U907 (N_907,N_56,N_127);
nor U908 (N_908,N_70,N_431);
nand U909 (N_909,N_464,N_218);
nand U910 (N_910,N_114,N_10);
and U911 (N_911,N_193,N_274);
nand U912 (N_912,N_91,N_395);
nand U913 (N_913,N_52,N_412);
nand U914 (N_914,N_167,N_261);
nor U915 (N_915,N_201,N_328);
nor U916 (N_916,N_361,N_458);
nor U917 (N_917,N_439,N_387);
or U918 (N_918,N_370,N_76);
nor U919 (N_919,N_403,N_349);
nand U920 (N_920,N_39,N_28);
or U921 (N_921,N_61,N_286);
nand U922 (N_922,N_303,N_450);
nor U923 (N_923,N_324,N_37);
and U924 (N_924,N_153,N_403);
nor U925 (N_925,N_273,N_26);
and U926 (N_926,N_115,N_453);
nand U927 (N_927,N_432,N_64);
or U928 (N_928,N_101,N_436);
xnor U929 (N_929,N_160,N_5);
nand U930 (N_930,N_419,N_257);
nand U931 (N_931,N_497,N_18);
nand U932 (N_932,N_55,N_156);
nor U933 (N_933,N_360,N_255);
nor U934 (N_934,N_495,N_323);
and U935 (N_935,N_239,N_219);
and U936 (N_936,N_293,N_407);
nand U937 (N_937,N_381,N_330);
or U938 (N_938,N_183,N_74);
nand U939 (N_939,N_29,N_46);
and U940 (N_940,N_445,N_77);
or U941 (N_941,N_455,N_226);
or U942 (N_942,N_268,N_491);
nand U943 (N_943,N_383,N_128);
nor U944 (N_944,N_38,N_307);
nand U945 (N_945,N_396,N_465);
nor U946 (N_946,N_376,N_295);
or U947 (N_947,N_227,N_310);
nor U948 (N_948,N_242,N_270);
or U949 (N_949,N_402,N_119);
nor U950 (N_950,N_235,N_52);
or U951 (N_951,N_269,N_370);
nor U952 (N_952,N_475,N_50);
nand U953 (N_953,N_114,N_485);
and U954 (N_954,N_197,N_201);
and U955 (N_955,N_363,N_435);
nor U956 (N_956,N_211,N_177);
nor U957 (N_957,N_412,N_51);
and U958 (N_958,N_354,N_284);
and U959 (N_959,N_34,N_338);
or U960 (N_960,N_134,N_159);
xor U961 (N_961,N_289,N_464);
nand U962 (N_962,N_393,N_59);
and U963 (N_963,N_404,N_392);
and U964 (N_964,N_256,N_474);
nand U965 (N_965,N_295,N_286);
or U966 (N_966,N_417,N_470);
and U967 (N_967,N_255,N_60);
nand U968 (N_968,N_430,N_7);
nand U969 (N_969,N_10,N_392);
and U970 (N_970,N_471,N_111);
nor U971 (N_971,N_449,N_193);
nand U972 (N_972,N_338,N_15);
or U973 (N_973,N_200,N_170);
nor U974 (N_974,N_428,N_338);
or U975 (N_975,N_37,N_451);
nor U976 (N_976,N_93,N_68);
and U977 (N_977,N_32,N_410);
or U978 (N_978,N_459,N_16);
xor U979 (N_979,N_334,N_234);
or U980 (N_980,N_38,N_211);
or U981 (N_981,N_473,N_149);
or U982 (N_982,N_109,N_130);
nand U983 (N_983,N_341,N_2);
nor U984 (N_984,N_41,N_472);
nand U985 (N_985,N_158,N_404);
or U986 (N_986,N_468,N_38);
nor U987 (N_987,N_56,N_345);
nand U988 (N_988,N_412,N_323);
nand U989 (N_989,N_421,N_223);
nor U990 (N_990,N_296,N_415);
nor U991 (N_991,N_187,N_450);
nor U992 (N_992,N_144,N_135);
nand U993 (N_993,N_423,N_191);
or U994 (N_994,N_68,N_493);
nand U995 (N_995,N_117,N_388);
and U996 (N_996,N_218,N_128);
nand U997 (N_997,N_157,N_161);
nand U998 (N_998,N_50,N_231);
nand U999 (N_999,N_337,N_175);
and U1000 (N_1000,N_770,N_715);
and U1001 (N_1001,N_868,N_917);
nand U1002 (N_1002,N_680,N_657);
or U1003 (N_1003,N_577,N_778);
or U1004 (N_1004,N_576,N_754);
or U1005 (N_1005,N_565,N_732);
or U1006 (N_1006,N_784,N_789);
nand U1007 (N_1007,N_767,N_834);
nand U1008 (N_1008,N_591,N_589);
and U1009 (N_1009,N_974,N_950);
and U1010 (N_1010,N_907,N_527);
xor U1011 (N_1011,N_551,N_507);
or U1012 (N_1012,N_859,N_983);
nand U1013 (N_1013,N_911,N_750);
nand U1014 (N_1014,N_888,N_587);
and U1015 (N_1015,N_891,N_547);
and U1016 (N_1016,N_634,N_906);
or U1017 (N_1017,N_875,N_599);
nor U1018 (N_1018,N_515,N_597);
and U1019 (N_1019,N_815,N_549);
nand U1020 (N_1020,N_632,N_532);
nand U1021 (N_1021,N_731,N_923);
nand U1022 (N_1022,N_668,N_658);
or U1023 (N_1023,N_713,N_830);
nor U1024 (N_1024,N_598,N_896);
nor U1025 (N_1025,N_762,N_782);
nor U1026 (N_1026,N_573,N_763);
nand U1027 (N_1027,N_989,N_707);
nor U1028 (N_1028,N_552,N_566);
nand U1029 (N_1029,N_776,N_948);
and U1030 (N_1030,N_753,N_991);
or U1031 (N_1031,N_909,N_742);
and U1032 (N_1032,N_662,N_640);
nor U1033 (N_1033,N_942,N_884);
nand U1034 (N_1034,N_864,N_572);
nand U1035 (N_1035,N_843,N_933);
nor U1036 (N_1036,N_929,N_590);
and U1037 (N_1037,N_535,N_669);
or U1038 (N_1038,N_853,N_897);
or U1039 (N_1039,N_749,N_813);
nor U1040 (N_1040,N_554,N_980);
nand U1041 (N_1041,N_930,N_705);
nor U1042 (N_1042,N_977,N_799);
or U1043 (N_1043,N_604,N_758);
nand U1044 (N_1044,N_663,N_880);
nand U1045 (N_1045,N_964,N_628);
nor U1046 (N_1046,N_956,N_938);
or U1047 (N_1047,N_722,N_866);
or U1048 (N_1048,N_733,N_684);
nand U1049 (N_1049,N_586,N_655);
or U1050 (N_1050,N_686,N_530);
or U1051 (N_1051,N_766,N_683);
nor U1052 (N_1052,N_903,N_534);
or U1053 (N_1053,N_809,N_806);
nand U1054 (N_1054,N_699,N_656);
and U1055 (N_1055,N_693,N_728);
or U1056 (N_1056,N_779,N_970);
and U1057 (N_1057,N_675,N_570);
nor U1058 (N_1058,N_642,N_837);
nor U1059 (N_1059,N_526,N_893);
nor U1060 (N_1060,N_624,N_678);
nor U1061 (N_1061,N_616,N_998);
or U1062 (N_1062,N_984,N_521);
nand U1063 (N_1063,N_506,N_646);
or U1064 (N_1064,N_730,N_787);
nand U1065 (N_1065,N_615,N_701);
nand U1066 (N_1066,N_503,N_921);
nand U1067 (N_1067,N_636,N_756);
or U1068 (N_1068,N_568,N_601);
nor U1069 (N_1069,N_714,N_982);
and U1070 (N_1070,N_919,N_945);
or U1071 (N_1071,N_772,N_935);
and U1072 (N_1072,N_988,N_650);
nand U1073 (N_1073,N_710,N_666);
nor U1074 (N_1074,N_553,N_500);
and U1075 (N_1075,N_606,N_882);
nor U1076 (N_1076,N_827,N_962);
and U1077 (N_1077,N_596,N_602);
nor U1078 (N_1078,N_621,N_873);
and U1079 (N_1079,N_865,N_785);
or U1080 (N_1080,N_965,N_517);
nand U1081 (N_1081,N_810,N_540);
nand U1082 (N_1082,N_892,N_777);
or U1083 (N_1083,N_968,N_605);
or U1084 (N_1084,N_885,N_995);
nor U1085 (N_1085,N_820,N_687);
and U1086 (N_1086,N_941,N_790);
nand U1087 (N_1087,N_940,N_773);
nand U1088 (N_1088,N_555,N_994);
nor U1089 (N_1089,N_594,N_505);
nor U1090 (N_1090,N_635,N_560);
and U1091 (N_1091,N_898,N_608);
nor U1092 (N_1092,N_775,N_856);
nand U1093 (N_1093,N_781,N_522);
and U1094 (N_1094,N_894,N_920);
nand U1095 (N_1095,N_845,N_957);
nand U1096 (N_1096,N_702,N_912);
nand U1097 (N_1097,N_824,N_890);
nor U1098 (N_1098,N_627,N_654);
or U1099 (N_1099,N_852,N_519);
and U1100 (N_1100,N_791,N_672);
and U1101 (N_1101,N_706,N_513);
and U1102 (N_1102,N_690,N_924);
and U1103 (N_1103,N_755,N_671);
nand U1104 (N_1104,N_703,N_708);
or U1105 (N_1105,N_895,N_871);
nand U1106 (N_1106,N_819,N_510);
and U1107 (N_1107,N_583,N_825);
nand U1108 (N_1108,N_881,N_694);
or U1109 (N_1109,N_518,N_828);
nor U1110 (N_1110,N_633,N_631);
or U1111 (N_1111,N_817,N_937);
or U1112 (N_1112,N_712,N_867);
nand U1113 (N_1113,N_639,N_508);
nand U1114 (N_1114,N_972,N_925);
nand U1115 (N_1115,N_794,N_764);
nor U1116 (N_1116,N_847,N_677);
and U1117 (N_1117,N_550,N_768);
nor U1118 (N_1118,N_936,N_543);
or U1119 (N_1119,N_927,N_786);
or U1120 (N_1120,N_709,N_716);
nand U1121 (N_1121,N_512,N_916);
nor U1122 (N_1122,N_674,N_575);
nor U1123 (N_1123,N_797,N_861);
or U1124 (N_1124,N_638,N_679);
or U1125 (N_1125,N_899,N_637);
nor U1126 (N_1126,N_878,N_665);
nand U1127 (N_1127,N_934,N_595);
or U1128 (N_1128,N_870,N_711);
nor U1129 (N_1129,N_939,N_879);
or U1130 (N_1130,N_719,N_826);
or U1131 (N_1131,N_533,N_973);
or U1132 (N_1132,N_954,N_793);
and U1133 (N_1133,N_664,N_643);
or U1134 (N_1134,N_805,N_823);
nor U1135 (N_1135,N_574,N_509);
or U1136 (N_1136,N_739,N_647);
nor U1137 (N_1137,N_821,N_800);
or U1138 (N_1138,N_831,N_996);
and U1139 (N_1139,N_611,N_959);
nand U1140 (N_1140,N_949,N_952);
or U1141 (N_1141,N_600,N_862);
and U1142 (N_1142,N_751,N_748);
and U1143 (N_1143,N_838,N_741);
or U1144 (N_1144,N_692,N_697);
nand U1145 (N_1145,N_963,N_734);
nand U1146 (N_1146,N_908,N_951);
and U1147 (N_1147,N_511,N_501);
nand U1148 (N_1148,N_557,N_607);
nor U1149 (N_1149,N_537,N_943);
nor U1150 (N_1150,N_584,N_807);
nand U1151 (N_1151,N_883,N_738);
nor U1152 (N_1152,N_997,N_849);
and U1153 (N_1153,N_999,N_617);
nor U1154 (N_1154,N_556,N_851);
and U1155 (N_1155,N_761,N_812);
nor U1156 (N_1156,N_542,N_516);
and U1157 (N_1157,N_649,N_618);
or U1158 (N_1158,N_946,N_659);
nand U1159 (N_1159,N_564,N_966);
nor U1160 (N_1160,N_769,N_569);
nor U1161 (N_1161,N_524,N_641);
nand U1162 (N_1162,N_613,N_676);
nand U1163 (N_1163,N_696,N_992);
nor U1164 (N_1164,N_774,N_840);
nand U1165 (N_1165,N_765,N_872);
nand U1166 (N_1166,N_900,N_736);
nand U1167 (N_1167,N_928,N_905);
and U1168 (N_1168,N_619,N_848);
nor U1169 (N_1169,N_660,N_829);
and U1170 (N_1170,N_609,N_889);
nand U1171 (N_1171,N_685,N_986);
nand U1172 (N_1172,N_653,N_582);
or U1173 (N_1173,N_559,N_585);
nor U1174 (N_1174,N_682,N_832);
nand U1175 (N_1175,N_796,N_610);
nand U1176 (N_1176,N_740,N_953);
or U1177 (N_1177,N_629,N_814);
nor U1178 (N_1178,N_944,N_546);
and U1179 (N_1179,N_688,N_645);
or U1180 (N_1180,N_743,N_985);
nor U1181 (N_1181,N_630,N_571);
and U1182 (N_1182,N_681,N_744);
nand U1183 (N_1183,N_700,N_661);
nor U1184 (N_1184,N_623,N_673);
or U1185 (N_1185,N_857,N_914);
nor U1186 (N_1186,N_579,N_548);
nor U1187 (N_1187,N_822,N_874);
and U1188 (N_1188,N_504,N_704);
or U1189 (N_1189,N_528,N_561);
and U1190 (N_1190,N_625,N_717);
and U1191 (N_1191,N_759,N_913);
and U1192 (N_1192,N_960,N_745);
nor U1193 (N_1193,N_648,N_538);
or U1194 (N_1194,N_808,N_816);
nand U1195 (N_1195,N_592,N_727);
and U1196 (N_1196,N_525,N_651);
nand U1197 (N_1197,N_918,N_798);
or U1198 (N_1198,N_863,N_689);
and U1199 (N_1199,N_698,N_969);
or U1200 (N_1200,N_620,N_588);
nand U1201 (N_1201,N_626,N_818);
and U1202 (N_1202,N_841,N_842);
and U1203 (N_1203,N_967,N_746);
and U1204 (N_1204,N_955,N_523);
and U1205 (N_1205,N_855,N_720);
or U1206 (N_1206,N_839,N_854);
and U1207 (N_1207,N_723,N_979);
and U1208 (N_1208,N_780,N_529);
and U1209 (N_1209,N_783,N_981);
or U1210 (N_1210,N_718,N_612);
xnor U1211 (N_1211,N_904,N_502);
or U1212 (N_1212,N_887,N_721);
and U1213 (N_1213,N_975,N_858);
or U1214 (N_1214,N_695,N_726);
and U1215 (N_1215,N_835,N_541);
or U1216 (N_1216,N_520,N_811);
and U1217 (N_1217,N_725,N_926);
nand U1218 (N_1218,N_987,N_978);
or U1219 (N_1219,N_578,N_536);
or U1220 (N_1220,N_846,N_729);
and U1221 (N_1221,N_932,N_788);
or U1222 (N_1222,N_910,N_947);
nand U1223 (N_1223,N_603,N_869);
and U1224 (N_1224,N_795,N_961);
or U1225 (N_1225,N_652,N_558);
or U1226 (N_1226,N_802,N_990);
nor U1227 (N_1227,N_563,N_792);
nand U1228 (N_1228,N_958,N_737);
and U1229 (N_1229,N_614,N_976);
nand U1230 (N_1230,N_735,N_545);
nand U1231 (N_1231,N_531,N_752);
or U1232 (N_1232,N_724,N_539);
and U1233 (N_1233,N_771,N_593);
nor U1234 (N_1234,N_670,N_747);
nor U1235 (N_1235,N_876,N_803);
nor U1236 (N_1236,N_562,N_902);
and U1237 (N_1237,N_544,N_931);
or U1238 (N_1238,N_757,N_836);
nand U1239 (N_1239,N_581,N_850);
or U1240 (N_1240,N_801,N_971);
nor U1241 (N_1241,N_760,N_804);
nand U1242 (N_1242,N_580,N_901);
or U1243 (N_1243,N_860,N_667);
nor U1244 (N_1244,N_567,N_877);
or U1245 (N_1245,N_886,N_993);
and U1246 (N_1246,N_514,N_844);
or U1247 (N_1247,N_833,N_915);
nor U1248 (N_1248,N_922,N_691);
or U1249 (N_1249,N_622,N_644);
and U1250 (N_1250,N_819,N_849);
and U1251 (N_1251,N_576,N_828);
and U1252 (N_1252,N_730,N_891);
nor U1253 (N_1253,N_712,N_718);
or U1254 (N_1254,N_787,N_988);
and U1255 (N_1255,N_505,N_651);
and U1256 (N_1256,N_669,N_572);
nand U1257 (N_1257,N_876,N_753);
nand U1258 (N_1258,N_995,N_726);
nand U1259 (N_1259,N_530,N_737);
nor U1260 (N_1260,N_661,N_757);
and U1261 (N_1261,N_666,N_949);
nand U1262 (N_1262,N_536,N_810);
and U1263 (N_1263,N_531,N_898);
nand U1264 (N_1264,N_905,N_577);
or U1265 (N_1265,N_950,N_805);
nor U1266 (N_1266,N_884,N_918);
and U1267 (N_1267,N_792,N_977);
or U1268 (N_1268,N_875,N_801);
xnor U1269 (N_1269,N_523,N_984);
and U1270 (N_1270,N_860,N_601);
or U1271 (N_1271,N_954,N_656);
or U1272 (N_1272,N_721,N_692);
nor U1273 (N_1273,N_946,N_838);
nor U1274 (N_1274,N_866,N_940);
nor U1275 (N_1275,N_603,N_620);
nand U1276 (N_1276,N_656,N_894);
and U1277 (N_1277,N_652,N_933);
nand U1278 (N_1278,N_519,N_622);
nor U1279 (N_1279,N_834,N_598);
nand U1280 (N_1280,N_887,N_634);
and U1281 (N_1281,N_595,N_570);
and U1282 (N_1282,N_748,N_505);
and U1283 (N_1283,N_882,N_869);
and U1284 (N_1284,N_866,N_529);
nor U1285 (N_1285,N_945,N_843);
nand U1286 (N_1286,N_636,N_710);
and U1287 (N_1287,N_910,N_797);
nand U1288 (N_1288,N_588,N_867);
nor U1289 (N_1289,N_598,N_574);
nand U1290 (N_1290,N_782,N_812);
and U1291 (N_1291,N_677,N_681);
or U1292 (N_1292,N_647,N_567);
nand U1293 (N_1293,N_636,N_964);
or U1294 (N_1294,N_707,N_547);
or U1295 (N_1295,N_510,N_589);
nand U1296 (N_1296,N_797,N_570);
nor U1297 (N_1297,N_990,N_993);
nor U1298 (N_1298,N_692,N_699);
nor U1299 (N_1299,N_926,N_601);
and U1300 (N_1300,N_736,N_905);
and U1301 (N_1301,N_785,N_925);
nand U1302 (N_1302,N_744,N_762);
and U1303 (N_1303,N_544,N_809);
or U1304 (N_1304,N_825,N_538);
and U1305 (N_1305,N_622,N_541);
and U1306 (N_1306,N_774,N_913);
nand U1307 (N_1307,N_851,N_852);
nor U1308 (N_1308,N_744,N_628);
nand U1309 (N_1309,N_676,N_624);
nor U1310 (N_1310,N_900,N_958);
and U1311 (N_1311,N_871,N_794);
nor U1312 (N_1312,N_618,N_619);
nor U1313 (N_1313,N_856,N_648);
or U1314 (N_1314,N_582,N_577);
nand U1315 (N_1315,N_877,N_668);
nand U1316 (N_1316,N_634,N_530);
and U1317 (N_1317,N_504,N_686);
nand U1318 (N_1318,N_575,N_547);
and U1319 (N_1319,N_968,N_610);
nor U1320 (N_1320,N_648,N_542);
or U1321 (N_1321,N_908,N_729);
nand U1322 (N_1322,N_694,N_800);
or U1323 (N_1323,N_893,N_895);
and U1324 (N_1324,N_544,N_798);
or U1325 (N_1325,N_700,N_906);
and U1326 (N_1326,N_513,N_917);
or U1327 (N_1327,N_752,N_796);
nand U1328 (N_1328,N_643,N_627);
nor U1329 (N_1329,N_650,N_763);
or U1330 (N_1330,N_614,N_879);
or U1331 (N_1331,N_606,N_593);
nand U1332 (N_1332,N_608,N_867);
or U1333 (N_1333,N_580,N_958);
or U1334 (N_1334,N_734,N_574);
nand U1335 (N_1335,N_730,N_651);
or U1336 (N_1336,N_954,N_533);
and U1337 (N_1337,N_759,N_820);
and U1338 (N_1338,N_888,N_925);
and U1339 (N_1339,N_745,N_883);
nor U1340 (N_1340,N_550,N_825);
nand U1341 (N_1341,N_879,N_785);
nand U1342 (N_1342,N_910,N_988);
or U1343 (N_1343,N_933,N_880);
or U1344 (N_1344,N_684,N_865);
and U1345 (N_1345,N_572,N_884);
nand U1346 (N_1346,N_791,N_675);
nor U1347 (N_1347,N_799,N_999);
nand U1348 (N_1348,N_838,N_994);
and U1349 (N_1349,N_876,N_730);
nand U1350 (N_1350,N_898,N_924);
nor U1351 (N_1351,N_570,N_694);
nand U1352 (N_1352,N_571,N_856);
or U1353 (N_1353,N_965,N_703);
nand U1354 (N_1354,N_985,N_937);
nand U1355 (N_1355,N_810,N_670);
and U1356 (N_1356,N_545,N_538);
nor U1357 (N_1357,N_786,N_944);
nand U1358 (N_1358,N_966,N_727);
nor U1359 (N_1359,N_722,N_852);
nand U1360 (N_1360,N_695,N_725);
or U1361 (N_1361,N_935,N_771);
and U1362 (N_1362,N_567,N_505);
or U1363 (N_1363,N_979,N_878);
nor U1364 (N_1364,N_785,N_923);
nor U1365 (N_1365,N_623,N_678);
nor U1366 (N_1366,N_722,N_511);
or U1367 (N_1367,N_997,N_951);
nor U1368 (N_1368,N_879,N_981);
or U1369 (N_1369,N_916,N_968);
and U1370 (N_1370,N_764,N_851);
nand U1371 (N_1371,N_608,N_848);
nand U1372 (N_1372,N_930,N_996);
nand U1373 (N_1373,N_503,N_612);
nand U1374 (N_1374,N_782,N_680);
or U1375 (N_1375,N_967,N_798);
nand U1376 (N_1376,N_767,N_807);
nor U1377 (N_1377,N_541,N_843);
nand U1378 (N_1378,N_607,N_757);
nor U1379 (N_1379,N_642,N_838);
nand U1380 (N_1380,N_659,N_746);
nor U1381 (N_1381,N_876,N_901);
or U1382 (N_1382,N_684,N_932);
and U1383 (N_1383,N_635,N_515);
nand U1384 (N_1384,N_786,N_995);
nor U1385 (N_1385,N_843,N_867);
nor U1386 (N_1386,N_940,N_507);
nand U1387 (N_1387,N_886,N_875);
nand U1388 (N_1388,N_655,N_973);
nand U1389 (N_1389,N_810,N_768);
or U1390 (N_1390,N_519,N_704);
and U1391 (N_1391,N_934,N_701);
and U1392 (N_1392,N_698,N_866);
nor U1393 (N_1393,N_821,N_600);
nor U1394 (N_1394,N_796,N_862);
nor U1395 (N_1395,N_584,N_937);
nand U1396 (N_1396,N_841,N_959);
nand U1397 (N_1397,N_650,N_814);
and U1398 (N_1398,N_508,N_790);
nor U1399 (N_1399,N_757,N_938);
nand U1400 (N_1400,N_806,N_546);
or U1401 (N_1401,N_534,N_966);
nor U1402 (N_1402,N_821,N_791);
xor U1403 (N_1403,N_663,N_614);
nor U1404 (N_1404,N_631,N_583);
nor U1405 (N_1405,N_831,N_851);
or U1406 (N_1406,N_962,N_594);
nand U1407 (N_1407,N_896,N_672);
and U1408 (N_1408,N_728,N_632);
and U1409 (N_1409,N_832,N_915);
nand U1410 (N_1410,N_870,N_856);
and U1411 (N_1411,N_722,N_624);
nor U1412 (N_1412,N_727,N_723);
nor U1413 (N_1413,N_582,N_891);
and U1414 (N_1414,N_563,N_528);
nand U1415 (N_1415,N_770,N_626);
nand U1416 (N_1416,N_864,N_682);
nand U1417 (N_1417,N_715,N_602);
and U1418 (N_1418,N_841,N_895);
or U1419 (N_1419,N_954,N_758);
or U1420 (N_1420,N_933,N_917);
nand U1421 (N_1421,N_629,N_682);
or U1422 (N_1422,N_914,N_509);
nor U1423 (N_1423,N_833,N_683);
or U1424 (N_1424,N_538,N_813);
or U1425 (N_1425,N_724,N_974);
and U1426 (N_1426,N_782,N_996);
nand U1427 (N_1427,N_558,N_949);
nand U1428 (N_1428,N_959,N_536);
nand U1429 (N_1429,N_811,N_696);
or U1430 (N_1430,N_715,N_653);
or U1431 (N_1431,N_562,N_720);
nand U1432 (N_1432,N_834,N_658);
nor U1433 (N_1433,N_815,N_825);
and U1434 (N_1434,N_726,N_851);
or U1435 (N_1435,N_554,N_811);
nor U1436 (N_1436,N_577,N_636);
nand U1437 (N_1437,N_894,N_881);
nand U1438 (N_1438,N_850,N_817);
or U1439 (N_1439,N_963,N_742);
or U1440 (N_1440,N_790,N_654);
nor U1441 (N_1441,N_823,N_591);
nor U1442 (N_1442,N_855,N_787);
and U1443 (N_1443,N_702,N_838);
xnor U1444 (N_1444,N_927,N_573);
or U1445 (N_1445,N_908,N_690);
nor U1446 (N_1446,N_667,N_976);
nor U1447 (N_1447,N_671,N_522);
nor U1448 (N_1448,N_674,N_733);
and U1449 (N_1449,N_858,N_781);
and U1450 (N_1450,N_503,N_764);
or U1451 (N_1451,N_668,N_786);
nor U1452 (N_1452,N_856,N_761);
nor U1453 (N_1453,N_632,N_667);
nor U1454 (N_1454,N_974,N_939);
nor U1455 (N_1455,N_607,N_953);
and U1456 (N_1456,N_892,N_548);
or U1457 (N_1457,N_748,N_853);
xor U1458 (N_1458,N_515,N_897);
nand U1459 (N_1459,N_733,N_964);
nor U1460 (N_1460,N_742,N_808);
nor U1461 (N_1461,N_739,N_511);
nand U1462 (N_1462,N_732,N_546);
or U1463 (N_1463,N_993,N_646);
nor U1464 (N_1464,N_853,N_912);
and U1465 (N_1465,N_914,N_931);
nor U1466 (N_1466,N_785,N_755);
nand U1467 (N_1467,N_513,N_976);
nor U1468 (N_1468,N_784,N_796);
or U1469 (N_1469,N_703,N_748);
or U1470 (N_1470,N_828,N_563);
or U1471 (N_1471,N_608,N_951);
nor U1472 (N_1472,N_659,N_660);
or U1473 (N_1473,N_581,N_825);
nor U1474 (N_1474,N_678,N_861);
nand U1475 (N_1475,N_600,N_788);
nor U1476 (N_1476,N_852,N_958);
or U1477 (N_1477,N_718,N_689);
nand U1478 (N_1478,N_938,N_583);
nor U1479 (N_1479,N_610,N_667);
nand U1480 (N_1480,N_778,N_688);
or U1481 (N_1481,N_967,N_869);
nand U1482 (N_1482,N_501,N_566);
or U1483 (N_1483,N_997,N_675);
or U1484 (N_1484,N_988,N_992);
xnor U1485 (N_1485,N_977,N_608);
nor U1486 (N_1486,N_577,N_509);
or U1487 (N_1487,N_624,N_877);
or U1488 (N_1488,N_818,N_504);
nand U1489 (N_1489,N_937,N_689);
nor U1490 (N_1490,N_556,N_695);
and U1491 (N_1491,N_684,N_690);
or U1492 (N_1492,N_982,N_685);
nand U1493 (N_1493,N_755,N_851);
and U1494 (N_1494,N_586,N_630);
and U1495 (N_1495,N_560,N_944);
or U1496 (N_1496,N_868,N_962);
and U1497 (N_1497,N_700,N_961);
or U1498 (N_1498,N_668,N_617);
and U1499 (N_1499,N_533,N_931);
nor U1500 (N_1500,N_1094,N_1486);
or U1501 (N_1501,N_1192,N_1251);
nor U1502 (N_1502,N_1349,N_1239);
nor U1503 (N_1503,N_1353,N_1404);
nor U1504 (N_1504,N_1198,N_1100);
nand U1505 (N_1505,N_1216,N_1218);
and U1506 (N_1506,N_1029,N_1378);
nor U1507 (N_1507,N_1053,N_1327);
or U1508 (N_1508,N_1169,N_1394);
or U1509 (N_1509,N_1446,N_1184);
and U1510 (N_1510,N_1114,N_1163);
nor U1511 (N_1511,N_1158,N_1146);
nor U1512 (N_1512,N_1337,N_1347);
or U1513 (N_1513,N_1051,N_1009);
and U1514 (N_1514,N_1076,N_1030);
or U1515 (N_1515,N_1139,N_1263);
nand U1516 (N_1516,N_1466,N_1361);
and U1517 (N_1517,N_1342,N_1215);
nor U1518 (N_1518,N_1127,N_1264);
nor U1519 (N_1519,N_1448,N_1429);
nor U1520 (N_1520,N_1091,N_1256);
xor U1521 (N_1521,N_1052,N_1095);
and U1522 (N_1522,N_1267,N_1444);
or U1523 (N_1523,N_1284,N_1418);
nand U1524 (N_1524,N_1307,N_1379);
and U1525 (N_1525,N_1490,N_1219);
nand U1526 (N_1526,N_1289,N_1322);
or U1527 (N_1527,N_1045,N_1299);
nand U1528 (N_1528,N_1381,N_1447);
or U1529 (N_1529,N_1089,N_1047);
nand U1530 (N_1530,N_1057,N_1334);
and U1531 (N_1531,N_1135,N_1093);
nor U1532 (N_1532,N_1373,N_1406);
nor U1533 (N_1533,N_1323,N_1084);
nor U1534 (N_1534,N_1385,N_1302);
nor U1535 (N_1535,N_1443,N_1066);
and U1536 (N_1536,N_1485,N_1255);
and U1537 (N_1537,N_1034,N_1123);
nand U1538 (N_1538,N_1027,N_1088);
nand U1539 (N_1539,N_1185,N_1132);
or U1540 (N_1540,N_1085,N_1395);
xnor U1541 (N_1541,N_1212,N_1413);
nand U1542 (N_1542,N_1268,N_1393);
or U1543 (N_1543,N_1261,N_1338);
nand U1544 (N_1544,N_1332,N_1205);
nand U1545 (N_1545,N_1040,N_1345);
and U1546 (N_1546,N_1285,N_1427);
and U1547 (N_1547,N_1401,N_1072);
nor U1548 (N_1548,N_1273,N_1229);
or U1549 (N_1549,N_1487,N_1206);
xor U1550 (N_1550,N_1309,N_1242);
and U1551 (N_1551,N_1455,N_1033);
nand U1552 (N_1552,N_1423,N_1121);
nor U1553 (N_1553,N_1343,N_1493);
or U1554 (N_1554,N_1318,N_1425);
nor U1555 (N_1555,N_1159,N_1037);
or U1556 (N_1556,N_1249,N_1228);
and U1557 (N_1557,N_1063,N_1010);
or U1558 (N_1558,N_1087,N_1186);
nor U1559 (N_1559,N_1213,N_1367);
and U1560 (N_1560,N_1305,N_1428);
nor U1561 (N_1561,N_1207,N_1131);
nand U1562 (N_1562,N_1036,N_1464);
or U1563 (N_1563,N_1293,N_1065);
or U1564 (N_1564,N_1150,N_1432);
nand U1565 (N_1565,N_1283,N_1203);
nor U1566 (N_1566,N_1227,N_1238);
nor U1567 (N_1567,N_1405,N_1271);
nand U1568 (N_1568,N_1116,N_1387);
and U1569 (N_1569,N_1001,N_1226);
nand U1570 (N_1570,N_1079,N_1004);
nand U1571 (N_1571,N_1300,N_1118);
nand U1572 (N_1572,N_1356,N_1411);
or U1573 (N_1573,N_1357,N_1348);
nand U1574 (N_1574,N_1438,N_1471);
nand U1575 (N_1575,N_1458,N_1380);
nor U1576 (N_1576,N_1086,N_1482);
nand U1577 (N_1577,N_1097,N_1152);
or U1578 (N_1578,N_1137,N_1360);
nand U1579 (N_1579,N_1117,N_1194);
and U1580 (N_1580,N_1246,N_1274);
nor U1581 (N_1581,N_1102,N_1195);
or U1582 (N_1582,N_1454,N_1382);
nand U1583 (N_1583,N_1422,N_1200);
or U1584 (N_1584,N_1377,N_1191);
or U1585 (N_1585,N_1145,N_1153);
or U1586 (N_1586,N_1155,N_1431);
nor U1587 (N_1587,N_1341,N_1176);
nor U1588 (N_1588,N_1397,N_1115);
or U1589 (N_1589,N_1151,N_1408);
or U1590 (N_1590,N_1005,N_1473);
and U1591 (N_1591,N_1099,N_1328);
nor U1592 (N_1592,N_1232,N_1056);
nor U1593 (N_1593,N_1237,N_1161);
nor U1594 (N_1594,N_1017,N_1269);
or U1595 (N_1595,N_1365,N_1409);
and U1596 (N_1596,N_1286,N_1080);
nand U1597 (N_1597,N_1225,N_1179);
nor U1598 (N_1598,N_1461,N_1495);
and U1599 (N_1599,N_1336,N_1164);
and U1600 (N_1600,N_1166,N_1025);
or U1601 (N_1601,N_1096,N_1190);
and U1602 (N_1602,N_1296,N_1217);
or U1603 (N_1603,N_1498,N_1193);
nand U1604 (N_1604,N_1488,N_1064);
nor U1605 (N_1605,N_1480,N_1149);
nor U1606 (N_1606,N_1110,N_1280);
and U1607 (N_1607,N_1074,N_1248);
and U1608 (N_1608,N_1259,N_1478);
and U1609 (N_1609,N_1143,N_1325);
or U1610 (N_1610,N_1371,N_1372);
and U1611 (N_1611,N_1124,N_1419);
and U1612 (N_1612,N_1060,N_1172);
nor U1613 (N_1613,N_1319,N_1039);
or U1614 (N_1614,N_1412,N_1188);
nor U1615 (N_1615,N_1333,N_1223);
or U1616 (N_1616,N_1407,N_1330);
and U1617 (N_1617,N_1295,N_1441);
nand U1618 (N_1618,N_1062,N_1258);
or U1619 (N_1619,N_1098,N_1277);
and U1620 (N_1620,N_1317,N_1230);
nor U1621 (N_1621,N_1463,N_1477);
nand U1622 (N_1622,N_1173,N_1003);
nor U1623 (N_1623,N_1414,N_1452);
nand U1624 (N_1624,N_1312,N_1031);
or U1625 (N_1625,N_1208,N_1311);
nor U1626 (N_1626,N_1374,N_1041);
nor U1627 (N_1627,N_1054,N_1292);
nand U1628 (N_1628,N_1134,N_1165);
and U1629 (N_1629,N_1083,N_1389);
or U1630 (N_1630,N_1388,N_1492);
nor U1631 (N_1631,N_1061,N_1266);
nand U1632 (N_1632,N_1018,N_1476);
and U1633 (N_1633,N_1043,N_1399);
and U1634 (N_1634,N_1433,N_1231);
xnor U1635 (N_1635,N_1294,N_1276);
nand U1636 (N_1636,N_1306,N_1346);
nand U1637 (N_1637,N_1424,N_1331);
or U1638 (N_1638,N_1032,N_1437);
and U1639 (N_1639,N_1368,N_1019);
and U1640 (N_1640,N_1105,N_1439);
nor U1641 (N_1641,N_1475,N_1253);
nand U1642 (N_1642,N_1339,N_1494);
nor U1643 (N_1643,N_1224,N_1314);
nor U1644 (N_1644,N_1375,N_1288);
and U1645 (N_1645,N_1055,N_1440);
nand U1646 (N_1646,N_1304,N_1035);
nor U1647 (N_1647,N_1484,N_1141);
and U1648 (N_1648,N_1369,N_1024);
and U1649 (N_1649,N_1092,N_1358);
nor U1650 (N_1650,N_1390,N_1026);
nand U1651 (N_1651,N_1257,N_1214);
and U1652 (N_1652,N_1170,N_1415);
nand U1653 (N_1653,N_1250,N_1303);
or U1654 (N_1654,N_1420,N_1351);
nand U1655 (N_1655,N_1221,N_1370);
and U1656 (N_1656,N_1016,N_1386);
nand U1657 (N_1657,N_1281,N_1260);
or U1658 (N_1658,N_1148,N_1142);
and U1659 (N_1659,N_1316,N_1359);
nand U1660 (N_1660,N_1081,N_1119);
or U1661 (N_1661,N_1362,N_1182);
nand U1662 (N_1662,N_1046,N_1183);
and U1663 (N_1663,N_1282,N_1021);
xnor U1664 (N_1664,N_1279,N_1136);
nor U1665 (N_1665,N_1298,N_1366);
nand U1666 (N_1666,N_1022,N_1403);
or U1667 (N_1667,N_1075,N_1210);
or U1668 (N_1668,N_1474,N_1107);
and U1669 (N_1669,N_1090,N_1197);
or U1670 (N_1670,N_1147,N_1180);
nor U1671 (N_1671,N_1236,N_1038);
and U1672 (N_1672,N_1398,N_1391);
nor U1673 (N_1673,N_1489,N_1290);
nand U1674 (N_1674,N_1417,N_1129);
or U1675 (N_1675,N_1340,N_1211);
and U1676 (N_1676,N_1326,N_1457);
or U1677 (N_1677,N_1077,N_1416);
nor U1678 (N_1678,N_1315,N_1156);
and U1679 (N_1679,N_1272,N_1450);
nor U1680 (N_1680,N_1234,N_1383);
or U1681 (N_1681,N_1042,N_1201);
or U1682 (N_1682,N_1265,N_1442);
nand U1683 (N_1683,N_1308,N_1449);
or U1684 (N_1684,N_1350,N_1059);
nor U1685 (N_1685,N_1128,N_1101);
nor U1686 (N_1686,N_1468,N_1291);
or U1687 (N_1687,N_1069,N_1011);
nand U1688 (N_1688,N_1483,N_1481);
nor U1689 (N_1689,N_1177,N_1028);
or U1690 (N_1690,N_1174,N_1111);
and U1691 (N_1691,N_1070,N_1058);
nor U1692 (N_1692,N_1122,N_1235);
and U1693 (N_1693,N_1199,N_1355);
or U1694 (N_1694,N_1469,N_1167);
and U1695 (N_1695,N_1071,N_1301);
and U1696 (N_1696,N_1049,N_1002);
or U1697 (N_1697,N_1426,N_1073);
and U1698 (N_1698,N_1445,N_1410);
and U1699 (N_1699,N_1321,N_1241);
nor U1700 (N_1700,N_1462,N_1364);
nor U1701 (N_1701,N_1310,N_1157);
nand U1702 (N_1702,N_1006,N_1344);
nand U1703 (N_1703,N_1275,N_1243);
and U1704 (N_1704,N_1352,N_1120);
nand U1705 (N_1705,N_1000,N_1392);
or U1706 (N_1706,N_1467,N_1082);
nand U1707 (N_1707,N_1112,N_1456);
nor U1708 (N_1708,N_1222,N_1181);
or U1709 (N_1709,N_1233,N_1220);
nor U1710 (N_1710,N_1068,N_1472);
or U1711 (N_1711,N_1434,N_1459);
nor U1712 (N_1712,N_1078,N_1106);
xnor U1713 (N_1713,N_1126,N_1320);
nand U1714 (N_1714,N_1144,N_1023);
nor U1715 (N_1715,N_1324,N_1244);
nor U1716 (N_1716,N_1154,N_1245);
or U1717 (N_1717,N_1113,N_1202);
or U1718 (N_1718,N_1050,N_1402);
and U1719 (N_1719,N_1460,N_1430);
nand U1720 (N_1720,N_1007,N_1189);
nand U1721 (N_1721,N_1162,N_1453);
and U1722 (N_1722,N_1209,N_1435);
or U1723 (N_1723,N_1178,N_1140);
nand U1724 (N_1724,N_1048,N_1013);
or U1725 (N_1725,N_1497,N_1020);
and U1726 (N_1726,N_1313,N_1204);
nor U1727 (N_1727,N_1109,N_1171);
or U1728 (N_1728,N_1384,N_1108);
nand U1729 (N_1729,N_1479,N_1499);
nand U1730 (N_1730,N_1125,N_1187);
nand U1731 (N_1731,N_1396,N_1067);
or U1732 (N_1732,N_1103,N_1354);
nand U1733 (N_1733,N_1044,N_1451);
and U1734 (N_1734,N_1014,N_1196);
nor U1735 (N_1735,N_1470,N_1104);
and U1736 (N_1736,N_1465,N_1363);
nor U1737 (N_1737,N_1240,N_1015);
and U1738 (N_1738,N_1130,N_1247);
or U1739 (N_1739,N_1491,N_1168);
nand U1740 (N_1740,N_1287,N_1436);
or U1741 (N_1741,N_1400,N_1160);
nor U1742 (N_1742,N_1254,N_1421);
xnor U1743 (N_1743,N_1376,N_1262);
and U1744 (N_1744,N_1012,N_1329);
xor U1745 (N_1745,N_1252,N_1278);
nand U1746 (N_1746,N_1297,N_1138);
nand U1747 (N_1747,N_1008,N_1335);
and U1748 (N_1748,N_1496,N_1133);
or U1749 (N_1749,N_1270,N_1175);
nor U1750 (N_1750,N_1369,N_1492);
nand U1751 (N_1751,N_1325,N_1323);
and U1752 (N_1752,N_1360,N_1098);
or U1753 (N_1753,N_1305,N_1209);
and U1754 (N_1754,N_1142,N_1247);
and U1755 (N_1755,N_1211,N_1259);
nor U1756 (N_1756,N_1284,N_1405);
and U1757 (N_1757,N_1174,N_1180);
nor U1758 (N_1758,N_1276,N_1259);
and U1759 (N_1759,N_1192,N_1244);
or U1760 (N_1760,N_1220,N_1276);
nand U1761 (N_1761,N_1304,N_1049);
nor U1762 (N_1762,N_1441,N_1168);
or U1763 (N_1763,N_1149,N_1453);
and U1764 (N_1764,N_1315,N_1105);
or U1765 (N_1765,N_1183,N_1304);
and U1766 (N_1766,N_1323,N_1466);
nand U1767 (N_1767,N_1271,N_1315);
and U1768 (N_1768,N_1375,N_1403);
or U1769 (N_1769,N_1370,N_1163);
or U1770 (N_1770,N_1083,N_1341);
nand U1771 (N_1771,N_1162,N_1038);
nand U1772 (N_1772,N_1478,N_1357);
nor U1773 (N_1773,N_1391,N_1034);
and U1774 (N_1774,N_1406,N_1042);
nor U1775 (N_1775,N_1192,N_1328);
nand U1776 (N_1776,N_1258,N_1197);
nor U1777 (N_1777,N_1247,N_1330);
nor U1778 (N_1778,N_1234,N_1470);
nand U1779 (N_1779,N_1234,N_1098);
and U1780 (N_1780,N_1033,N_1129);
and U1781 (N_1781,N_1256,N_1270);
or U1782 (N_1782,N_1419,N_1178);
nor U1783 (N_1783,N_1308,N_1336);
nand U1784 (N_1784,N_1422,N_1087);
nand U1785 (N_1785,N_1300,N_1469);
nor U1786 (N_1786,N_1319,N_1301);
nor U1787 (N_1787,N_1351,N_1116);
or U1788 (N_1788,N_1448,N_1484);
or U1789 (N_1789,N_1497,N_1243);
and U1790 (N_1790,N_1206,N_1365);
nand U1791 (N_1791,N_1098,N_1430);
or U1792 (N_1792,N_1055,N_1493);
nor U1793 (N_1793,N_1398,N_1043);
xor U1794 (N_1794,N_1498,N_1262);
or U1795 (N_1795,N_1270,N_1437);
or U1796 (N_1796,N_1377,N_1337);
or U1797 (N_1797,N_1290,N_1138);
or U1798 (N_1798,N_1194,N_1206);
and U1799 (N_1799,N_1371,N_1430);
and U1800 (N_1800,N_1443,N_1310);
nand U1801 (N_1801,N_1016,N_1294);
nor U1802 (N_1802,N_1490,N_1180);
and U1803 (N_1803,N_1128,N_1462);
nor U1804 (N_1804,N_1264,N_1474);
nor U1805 (N_1805,N_1417,N_1172);
and U1806 (N_1806,N_1268,N_1034);
or U1807 (N_1807,N_1461,N_1080);
and U1808 (N_1808,N_1470,N_1006);
nand U1809 (N_1809,N_1163,N_1368);
nor U1810 (N_1810,N_1181,N_1269);
or U1811 (N_1811,N_1477,N_1355);
and U1812 (N_1812,N_1054,N_1225);
nand U1813 (N_1813,N_1486,N_1050);
nand U1814 (N_1814,N_1303,N_1185);
and U1815 (N_1815,N_1318,N_1476);
or U1816 (N_1816,N_1345,N_1189);
nor U1817 (N_1817,N_1228,N_1159);
nand U1818 (N_1818,N_1303,N_1087);
nand U1819 (N_1819,N_1232,N_1405);
and U1820 (N_1820,N_1055,N_1060);
nor U1821 (N_1821,N_1283,N_1184);
nor U1822 (N_1822,N_1487,N_1448);
nor U1823 (N_1823,N_1248,N_1306);
or U1824 (N_1824,N_1014,N_1428);
and U1825 (N_1825,N_1119,N_1115);
nor U1826 (N_1826,N_1199,N_1175);
or U1827 (N_1827,N_1140,N_1462);
nor U1828 (N_1828,N_1083,N_1016);
nor U1829 (N_1829,N_1345,N_1457);
nand U1830 (N_1830,N_1052,N_1302);
nor U1831 (N_1831,N_1285,N_1288);
or U1832 (N_1832,N_1269,N_1455);
and U1833 (N_1833,N_1141,N_1235);
nand U1834 (N_1834,N_1218,N_1321);
or U1835 (N_1835,N_1419,N_1340);
nor U1836 (N_1836,N_1172,N_1307);
nor U1837 (N_1837,N_1194,N_1198);
nor U1838 (N_1838,N_1430,N_1448);
and U1839 (N_1839,N_1134,N_1078);
nor U1840 (N_1840,N_1002,N_1150);
and U1841 (N_1841,N_1250,N_1014);
or U1842 (N_1842,N_1496,N_1088);
nor U1843 (N_1843,N_1239,N_1232);
nor U1844 (N_1844,N_1037,N_1465);
or U1845 (N_1845,N_1293,N_1197);
nand U1846 (N_1846,N_1456,N_1211);
nor U1847 (N_1847,N_1289,N_1215);
nand U1848 (N_1848,N_1036,N_1092);
or U1849 (N_1849,N_1378,N_1413);
nand U1850 (N_1850,N_1377,N_1058);
nor U1851 (N_1851,N_1392,N_1299);
or U1852 (N_1852,N_1266,N_1445);
and U1853 (N_1853,N_1336,N_1317);
nand U1854 (N_1854,N_1264,N_1390);
nor U1855 (N_1855,N_1010,N_1380);
or U1856 (N_1856,N_1163,N_1451);
nand U1857 (N_1857,N_1223,N_1417);
or U1858 (N_1858,N_1145,N_1186);
xnor U1859 (N_1859,N_1465,N_1354);
nor U1860 (N_1860,N_1498,N_1367);
nor U1861 (N_1861,N_1358,N_1280);
and U1862 (N_1862,N_1240,N_1200);
nand U1863 (N_1863,N_1330,N_1273);
nand U1864 (N_1864,N_1344,N_1382);
and U1865 (N_1865,N_1366,N_1387);
and U1866 (N_1866,N_1412,N_1069);
nand U1867 (N_1867,N_1161,N_1063);
nor U1868 (N_1868,N_1151,N_1230);
and U1869 (N_1869,N_1144,N_1098);
and U1870 (N_1870,N_1389,N_1123);
nand U1871 (N_1871,N_1363,N_1091);
nand U1872 (N_1872,N_1306,N_1024);
nand U1873 (N_1873,N_1019,N_1202);
nor U1874 (N_1874,N_1411,N_1116);
nor U1875 (N_1875,N_1201,N_1158);
or U1876 (N_1876,N_1495,N_1036);
and U1877 (N_1877,N_1263,N_1191);
and U1878 (N_1878,N_1292,N_1216);
nand U1879 (N_1879,N_1492,N_1402);
and U1880 (N_1880,N_1456,N_1235);
and U1881 (N_1881,N_1487,N_1327);
and U1882 (N_1882,N_1333,N_1019);
and U1883 (N_1883,N_1116,N_1114);
and U1884 (N_1884,N_1377,N_1432);
nor U1885 (N_1885,N_1391,N_1010);
nor U1886 (N_1886,N_1103,N_1384);
or U1887 (N_1887,N_1322,N_1397);
and U1888 (N_1888,N_1498,N_1170);
or U1889 (N_1889,N_1391,N_1151);
xor U1890 (N_1890,N_1476,N_1280);
nand U1891 (N_1891,N_1361,N_1139);
nor U1892 (N_1892,N_1176,N_1021);
nor U1893 (N_1893,N_1043,N_1300);
and U1894 (N_1894,N_1056,N_1457);
nand U1895 (N_1895,N_1143,N_1221);
nor U1896 (N_1896,N_1371,N_1031);
nor U1897 (N_1897,N_1341,N_1042);
or U1898 (N_1898,N_1009,N_1210);
nor U1899 (N_1899,N_1074,N_1315);
or U1900 (N_1900,N_1385,N_1245);
or U1901 (N_1901,N_1266,N_1003);
nand U1902 (N_1902,N_1235,N_1461);
and U1903 (N_1903,N_1373,N_1433);
or U1904 (N_1904,N_1283,N_1207);
and U1905 (N_1905,N_1115,N_1450);
nor U1906 (N_1906,N_1340,N_1481);
nand U1907 (N_1907,N_1432,N_1367);
nor U1908 (N_1908,N_1209,N_1451);
or U1909 (N_1909,N_1377,N_1495);
or U1910 (N_1910,N_1140,N_1370);
xnor U1911 (N_1911,N_1327,N_1122);
and U1912 (N_1912,N_1046,N_1257);
nand U1913 (N_1913,N_1399,N_1167);
or U1914 (N_1914,N_1412,N_1313);
and U1915 (N_1915,N_1000,N_1236);
and U1916 (N_1916,N_1119,N_1421);
nor U1917 (N_1917,N_1330,N_1268);
nand U1918 (N_1918,N_1199,N_1281);
nor U1919 (N_1919,N_1126,N_1381);
nor U1920 (N_1920,N_1474,N_1425);
nand U1921 (N_1921,N_1353,N_1011);
nor U1922 (N_1922,N_1315,N_1259);
and U1923 (N_1923,N_1254,N_1424);
nand U1924 (N_1924,N_1275,N_1475);
nand U1925 (N_1925,N_1443,N_1469);
and U1926 (N_1926,N_1354,N_1331);
and U1927 (N_1927,N_1430,N_1148);
or U1928 (N_1928,N_1351,N_1020);
nand U1929 (N_1929,N_1190,N_1229);
and U1930 (N_1930,N_1197,N_1417);
nand U1931 (N_1931,N_1227,N_1308);
and U1932 (N_1932,N_1222,N_1365);
and U1933 (N_1933,N_1478,N_1121);
and U1934 (N_1934,N_1456,N_1024);
nand U1935 (N_1935,N_1195,N_1244);
nor U1936 (N_1936,N_1367,N_1010);
and U1937 (N_1937,N_1028,N_1475);
nand U1938 (N_1938,N_1454,N_1183);
or U1939 (N_1939,N_1495,N_1180);
or U1940 (N_1940,N_1284,N_1058);
or U1941 (N_1941,N_1200,N_1457);
and U1942 (N_1942,N_1094,N_1174);
or U1943 (N_1943,N_1344,N_1122);
or U1944 (N_1944,N_1413,N_1355);
and U1945 (N_1945,N_1402,N_1404);
and U1946 (N_1946,N_1197,N_1065);
nand U1947 (N_1947,N_1065,N_1499);
and U1948 (N_1948,N_1163,N_1037);
or U1949 (N_1949,N_1458,N_1146);
nand U1950 (N_1950,N_1143,N_1387);
nand U1951 (N_1951,N_1372,N_1035);
nor U1952 (N_1952,N_1329,N_1245);
or U1953 (N_1953,N_1137,N_1430);
nor U1954 (N_1954,N_1280,N_1064);
and U1955 (N_1955,N_1146,N_1497);
nand U1956 (N_1956,N_1390,N_1402);
and U1957 (N_1957,N_1386,N_1231);
nand U1958 (N_1958,N_1251,N_1132);
nand U1959 (N_1959,N_1102,N_1438);
or U1960 (N_1960,N_1369,N_1031);
nand U1961 (N_1961,N_1346,N_1426);
and U1962 (N_1962,N_1351,N_1384);
nand U1963 (N_1963,N_1222,N_1079);
nand U1964 (N_1964,N_1176,N_1490);
or U1965 (N_1965,N_1385,N_1050);
nor U1966 (N_1966,N_1388,N_1391);
nor U1967 (N_1967,N_1060,N_1352);
and U1968 (N_1968,N_1010,N_1048);
nand U1969 (N_1969,N_1318,N_1427);
or U1970 (N_1970,N_1218,N_1059);
and U1971 (N_1971,N_1192,N_1023);
or U1972 (N_1972,N_1485,N_1004);
or U1973 (N_1973,N_1046,N_1497);
nor U1974 (N_1974,N_1297,N_1159);
nand U1975 (N_1975,N_1277,N_1377);
and U1976 (N_1976,N_1268,N_1128);
nand U1977 (N_1977,N_1373,N_1325);
nand U1978 (N_1978,N_1247,N_1325);
and U1979 (N_1979,N_1078,N_1113);
nor U1980 (N_1980,N_1230,N_1069);
and U1981 (N_1981,N_1158,N_1150);
or U1982 (N_1982,N_1193,N_1220);
nor U1983 (N_1983,N_1318,N_1166);
nor U1984 (N_1984,N_1339,N_1065);
and U1985 (N_1985,N_1322,N_1027);
or U1986 (N_1986,N_1140,N_1471);
or U1987 (N_1987,N_1357,N_1427);
nand U1988 (N_1988,N_1473,N_1260);
or U1989 (N_1989,N_1003,N_1052);
nand U1990 (N_1990,N_1111,N_1361);
and U1991 (N_1991,N_1273,N_1366);
and U1992 (N_1992,N_1156,N_1035);
nor U1993 (N_1993,N_1297,N_1214);
and U1994 (N_1994,N_1076,N_1185);
and U1995 (N_1995,N_1443,N_1018);
nand U1996 (N_1996,N_1460,N_1126);
and U1997 (N_1997,N_1152,N_1413);
or U1998 (N_1998,N_1162,N_1084);
or U1999 (N_1999,N_1072,N_1033);
nand U2000 (N_2000,N_1622,N_1507);
or U2001 (N_2001,N_1550,N_1871);
or U2002 (N_2002,N_1561,N_1925);
nand U2003 (N_2003,N_1753,N_1944);
nand U2004 (N_2004,N_1694,N_1981);
nand U2005 (N_2005,N_1829,N_1835);
nor U2006 (N_2006,N_1548,N_1711);
or U2007 (N_2007,N_1921,N_1770);
nor U2008 (N_2008,N_1596,N_1978);
nor U2009 (N_2009,N_1927,N_1765);
nand U2010 (N_2010,N_1962,N_1710);
or U2011 (N_2011,N_1784,N_1931);
and U2012 (N_2012,N_1783,N_1680);
nor U2013 (N_2013,N_1964,N_1741);
xnor U2014 (N_2014,N_1778,N_1584);
nor U2015 (N_2015,N_1712,N_1594);
or U2016 (N_2016,N_1938,N_1716);
nor U2017 (N_2017,N_1677,N_1563);
and U2018 (N_2018,N_1565,N_1794);
nand U2019 (N_2019,N_1887,N_1847);
nor U2020 (N_2020,N_1913,N_1980);
nand U2021 (N_2021,N_1676,N_1575);
and U2022 (N_2022,N_1880,N_1874);
nand U2023 (N_2023,N_1841,N_1525);
nand U2024 (N_2024,N_1616,N_1828);
nand U2025 (N_2025,N_1678,N_1690);
or U2026 (N_2026,N_1912,N_1929);
nor U2027 (N_2027,N_1762,N_1823);
and U2028 (N_2028,N_1693,N_1569);
nor U2029 (N_2029,N_1918,N_1746);
and U2030 (N_2030,N_1990,N_1519);
and U2031 (N_2031,N_1708,N_1850);
or U2032 (N_2032,N_1568,N_1706);
nand U2033 (N_2033,N_1760,N_1956);
nor U2034 (N_2034,N_1599,N_1897);
or U2035 (N_2035,N_1904,N_1605);
or U2036 (N_2036,N_1894,N_1846);
nor U2037 (N_2037,N_1864,N_1876);
nand U2038 (N_2038,N_1902,N_1722);
or U2039 (N_2039,N_1739,N_1977);
and U2040 (N_2040,N_1907,N_1808);
nor U2041 (N_2041,N_1941,N_1609);
or U2042 (N_2042,N_1667,N_1911);
nand U2043 (N_2043,N_1951,N_1662);
nor U2044 (N_2044,N_1679,N_1703);
nor U2045 (N_2045,N_1836,N_1700);
nand U2046 (N_2046,N_1578,N_1500);
nor U2047 (N_2047,N_1772,N_1786);
nand U2048 (N_2048,N_1669,N_1810);
and U2049 (N_2049,N_1627,N_1825);
nand U2050 (N_2050,N_1534,N_1623);
nand U2051 (N_2051,N_1502,N_1571);
nand U2052 (N_2052,N_1636,N_1792);
or U2053 (N_2053,N_1645,N_1892);
and U2054 (N_2054,N_1940,N_1854);
nor U2055 (N_2055,N_1668,N_1558);
nand U2056 (N_2056,N_1625,N_1769);
or U2057 (N_2057,N_1849,N_1795);
nor U2058 (N_2058,N_1952,N_1691);
or U2059 (N_2059,N_1949,N_1654);
nor U2060 (N_2060,N_1814,N_1666);
or U2061 (N_2061,N_1920,N_1861);
nor U2062 (N_2062,N_1801,N_1501);
and U2063 (N_2063,N_1833,N_1603);
nor U2064 (N_2064,N_1615,N_1805);
or U2065 (N_2065,N_1663,N_1881);
nand U2066 (N_2066,N_1511,N_1560);
or U2067 (N_2067,N_1797,N_1540);
and U2068 (N_2068,N_1509,N_1858);
or U2069 (N_2069,N_1592,N_1909);
nor U2070 (N_2070,N_1877,N_1777);
and U2071 (N_2071,N_1544,N_1910);
or U2072 (N_2072,N_1838,N_1787);
and U2073 (N_2073,N_1837,N_1776);
nand U2074 (N_2074,N_1661,N_1974);
xnor U2075 (N_2075,N_1896,N_1705);
nand U2076 (N_2076,N_1597,N_1843);
and U2077 (N_2077,N_1779,N_1689);
nand U2078 (N_2078,N_1785,N_1757);
nand U2079 (N_2079,N_1885,N_1947);
nor U2080 (N_2080,N_1960,N_1923);
nand U2081 (N_2081,N_1901,N_1748);
or U2082 (N_2082,N_1724,N_1988);
nor U2083 (N_2083,N_1524,N_1655);
or U2084 (N_2084,N_1733,N_1798);
and U2085 (N_2085,N_1506,N_1844);
nand U2086 (N_2086,N_1728,N_1732);
nand U2087 (N_2087,N_1889,N_1867);
nand U2088 (N_2088,N_1868,N_1687);
nand U2089 (N_2089,N_1865,N_1851);
nand U2090 (N_2090,N_1698,N_1780);
nor U2091 (N_2091,N_1755,N_1989);
and U2092 (N_2092,N_1613,N_1933);
and U2093 (N_2093,N_1611,N_1945);
xor U2094 (N_2094,N_1857,N_1660);
nand U2095 (N_2095,N_1782,N_1827);
nand U2096 (N_2096,N_1866,N_1517);
nor U2097 (N_2097,N_1740,N_1715);
or U2098 (N_2098,N_1527,N_1656);
nor U2099 (N_2099,N_1598,N_1738);
nor U2100 (N_2100,N_1518,N_1766);
xnor U2101 (N_2101,N_1817,N_1872);
nor U2102 (N_2102,N_1917,N_1900);
nand U2103 (N_2103,N_1618,N_1950);
and U2104 (N_2104,N_1652,N_1556);
or U2105 (N_2105,N_1579,N_1580);
or U2106 (N_2106,N_1685,N_1873);
or U2107 (N_2107,N_1612,N_1670);
and U2108 (N_2108,N_1818,N_1649);
nand U2109 (N_2109,N_1862,N_1528);
nor U2110 (N_2110,N_1961,N_1747);
or U2111 (N_2111,N_1713,N_1538);
nor U2112 (N_2112,N_1939,N_1781);
or U2113 (N_2113,N_1632,N_1574);
nor U2114 (N_2114,N_1800,N_1984);
nand U2115 (N_2115,N_1750,N_1727);
nor U2116 (N_2116,N_1513,N_1635);
and U2117 (N_2117,N_1788,N_1566);
or U2118 (N_2118,N_1930,N_1811);
nor U2119 (N_2119,N_1614,N_1620);
nor U2120 (N_2120,N_1761,N_1503);
or U2121 (N_2121,N_1752,N_1600);
and U2122 (N_2122,N_1692,N_1659);
and U2123 (N_2123,N_1512,N_1729);
or U2124 (N_2124,N_1573,N_1948);
and U2125 (N_2125,N_1975,N_1546);
or U2126 (N_2126,N_1651,N_1553);
or U2127 (N_2127,N_1510,N_1842);
nor U2128 (N_2128,N_1957,N_1735);
nand U2129 (N_2129,N_1799,N_1943);
and U2130 (N_2130,N_1526,N_1533);
nor U2131 (N_2131,N_1815,N_1520);
and U2132 (N_2132,N_1775,N_1886);
or U2133 (N_2133,N_1767,N_1759);
nand U2134 (N_2134,N_1906,N_1914);
nor U2135 (N_2135,N_1522,N_1826);
nand U2136 (N_2136,N_1791,N_1768);
nor U2137 (N_2137,N_1664,N_1591);
nor U2138 (N_2138,N_1607,N_1514);
or U2139 (N_2139,N_1640,N_1999);
nor U2140 (N_2140,N_1884,N_1725);
nor U2141 (N_2141,N_1587,N_1505);
nand U2142 (N_2142,N_1545,N_1987);
and U2143 (N_2143,N_1971,N_1749);
or U2144 (N_2144,N_1863,N_1982);
and U2145 (N_2145,N_1848,N_1870);
or U2146 (N_2146,N_1802,N_1852);
or U2147 (N_2147,N_1672,N_1806);
nor U2148 (N_2148,N_1572,N_1602);
nand U2149 (N_2149,N_1995,N_1665);
and U2150 (N_2150,N_1972,N_1695);
and U2151 (N_2151,N_1963,N_1754);
xor U2152 (N_2152,N_1993,N_1644);
nand U2153 (N_2153,N_1577,N_1634);
nor U2154 (N_2154,N_1824,N_1744);
and U2155 (N_2155,N_1552,N_1922);
nand U2156 (N_2156,N_1629,N_1919);
nand U2157 (N_2157,N_1721,N_1576);
nor U2158 (N_2158,N_1883,N_1646);
or U2159 (N_2159,N_1719,N_1859);
nand U2160 (N_2160,N_1899,N_1832);
nor U2161 (N_2161,N_1586,N_1756);
nor U2162 (N_2162,N_1658,N_1955);
nand U2163 (N_2163,N_1953,N_1840);
nand U2164 (N_2164,N_1581,N_1585);
or U2165 (N_2165,N_1908,N_1699);
nand U2166 (N_2166,N_1819,N_1875);
nand U2167 (N_2167,N_1926,N_1869);
nand U2168 (N_2168,N_1954,N_1935);
or U2169 (N_2169,N_1589,N_1895);
and U2170 (N_2170,N_1773,N_1682);
and U2171 (N_2171,N_1970,N_1532);
xnor U2172 (N_2172,N_1630,N_1915);
or U2173 (N_2173,N_1504,N_1812);
or U2174 (N_2174,N_1834,N_1718);
and U2175 (N_2175,N_1822,N_1588);
and U2176 (N_2176,N_1643,N_1707);
nand U2177 (N_2177,N_1702,N_1709);
nand U2178 (N_2178,N_1638,N_1606);
nand U2179 (N_2179,N_1946,N_1958);
or U2180 (N_2180,N_1617,N_1582);
nand U2181 (N_2181,N_1839,N_1903);
nor U2182 (N_2182,N_1515,N_1924);
nor U2183 (N_2183,N_1973,N_1541);
or U2184 (N_2184,N_1555,N_1998);
nor U2185 (N_2185,N_1619,N_1816);
and U2186 (N_2186,N_1539,N_1845);
and U2187 (N_2187,N_1821,N_1804);
or U2188 (N_2188,N_1969,N_1564);
nand U2189 (N_2189,N_1893,N_1905);
nand U2190 (N_2190,N_1967,N_1976);
or U2191 (N_2191,N_1542,N_1774);
nand U2192 (N_2192,N_1628,N_1830);
or U2193 (N_2193,N_1763,N_1535);
and U2194 (N_2194,N_1531,N_1593);
and U2195 (N_2195,N_1683,N_1523);
nand U2196 (N_2196,N_1916,N_1701);
nand U2197 (N_2197,N_1626,N_1809);
xnor U2198 (N_2198,N_1608,N_1742);
or U2199 (N_2199,N_1521,N_1820);
and U2200 (N_2200,N_1991,N_1583);
and U2201 (N_2201,N_1994,N_1734);
nand U2202 (N_2202,N_1537,N_1888);
nor U2203 (N_2203,N_1595,N_1688);
nand U2204 (N_2204,N_1932,N_1726);
and U2205 (N_2205,N_1601,N_1997);
nand U2206 (N_2206,N_1547,N_1697);
or U2207 (N_2207,N_1717,N_1959);
nand U2208 (N_2208,N_1704,N_1807);
and U2209 (N_2209,N_1675,N_1508);
nand U2210 (N_2210,N_1657,N_1966);
or U2211 (N_2211,N_1559,N_1631);
nand U2212 (N_2212,N_1771,N_1639);
or U2213 (N_2213,N_1604,N_1879);
and U2214 (N_2214,N_1684,N_1673);
nor U2215 (N_2215,N_1793,N_1714);
and U2216 (N_2216,N_1890,N_1562);
nand U2217 (N_2217,N_1731,N_1557);
nand U2218 (N_2218,N_1554,N_1621);
nor U2219 (N_2219,N_1751,N_1551);
and U2220 (N_2220,N_1674,N_1648);
and U2221 (N_2221,N_1720,N_1567);
nand U2222 (N_2222,N_1745,N_1856);
or U2223 (N_2223,N_1996,N_1671);
and U2224 (N_2224,N_1965,N_1985);
or U2225 (N_2225,N_1516,N_1743);
nor U2226 (N_2226,N_1853,N_1813);
and U2227 (N_2227,N_1543,N_1878);
and U2228 (N_2228,N_1570,N_1653);
nor U2229 (N_2229,N_1928,N_1641);
and U2230 (N_2230,N_1992,N_1764);
nor U2231 (N_2231,N_1898,N_1530);
and U2232 (N_2232,N_1647,N_1855);
or U2233 (N_2233,N_1979,N_1937);
nand U2234 (N_2234,N_1803,N_1737);
or U2235 (N_2235,N_1624,N_1882);
or U2236 (N_2236,N_1681,N_1790);
nor U2237 (N_2237,N_1891,N_1736);
nor U2238 (N_2238,N_1936,N_1723);
or U2239 (N_2239,N_1529,N_1642);
nor U2240 (N_2240,N_1610,N_1789);
and U2241 (N_2241,N_1983,N_1686);
nand U2242 (N_2242,N_1536,N_1549);
nor U2243 (N_2243,N_1934,N_1637);
or U2244 (N_2244,N_1796,N_1831);
or U2245 (N_2245,N_1968,N_1986);
or U2246 (N_2246,N_1942,N_1590);
nand U2247 (N_2247,N_1758,N_1633);
or U2248 (N_2248,N_1730,N_1650);
nor U2249 (N_2249,N_1696,N_1860);
nor U2250 (N_2250,N_1958,N_1763);
or U2251 (N_2251,N_1713,N_1535);
or U2252 (N_2252,N_1748,N_1744);
nand U2253 (N_2253,N_1840,N_1875);
and U2254 (N_2254,N_1690,N_1739);
or U2255 (N_2255,N_1943,N_1571);
and U2256 (N_2256,N_1934,N_1775);
xnor U2257 (N_2257,N_1961,N_1950);
or U2258 (N_2258,N_1674,N_1805);
nand U2259 (N_2259,N_1993,N_1705);
and U2260 (N_2260,N_1678,N_1961);
and U2261 (N_2261,N_1632,N_1540);
nand U2262 (N_2262,N_1853,N_1577);
or U2263 (N_2263,N_1661,N_1822);
nor U2264 (N_2264,N_1839,N_1955);
nor U2265 (N_2265,N_1512,N_1882);
nand U2266 (N_2266,N_1590,N_1579);
and U2267 (N_2267,N_1642,N_1809);
or U2268 (N_2268,N_1643,N_1653);
or U2269 (N_2269,N_1937,N_1630);
or U2270 (N_2270,N_1885,N_1533);
or U2271 (N_2271,N_1715,N_1959);
and U2272 (N_2272,N_1593,N_1631);
nand U2273 (N_2273,N_1624,N_1781);
nor U2274 (N_2274,N_1721,N_1983);
or U2275 (N_2275,N_1523,N_1716);
or U2276 (N_2276,N_1516,N_1570);
or U2277 (N_2277,N_1850,N_1902);
nor U2278 (N_2278,N_1578,N_1590);
and U2279 (N_2279,N_1936,N_1536);
nand U2280 (N_2280,N_1844,N_1661);
and U2281 (N_2281,N_1769,N_1758);
nand U2282 (N_2282,N_1722,N_1623);
nand U2283 (N_2283,N_1572,N_1611);
nor U2284 (N_2284,N_1578,N_1589);
and U2285 (N_2285,N_1904,N_1527);
or U2286 (N_2286,N_1927,N_1869);
and U2287 (N_2287,N_1599,N_1669);
and U2288 (N_2288,N_1994,N_1995);
or U2289 (N_2289,N_1739,N_1553);
and U2290 (N_2290,N_1711,N_1872);
and U2291 (N_2291,N_1896,N_1654);
nand U2292 (N_2292,N_1842,N_1638);
and U2293 (N_2293,N_1990,N_1979);
nand U2294 (N_2294,N_1552,N_1570);
nand U2295 (N_2295,N_1897,N_1596);
and U2296 (N_2296,N_1590,N_1551);
and U2297 (N_2297,N_1537,N_1542);
and U2298 (N_2298,N_1850,N_1529);
or U2299 (N_2299,N_1949,N_1551);
and U2300 (N_2300,N_1517,N_1902);
nand U2301 (N_2301,N_1841,N_1811);
and U2302 (N_2302,N_1603,N_1952);
and U2303 (N_2303,N_1850,N_1797);
or U2304 (N_2304,N_1798,N_1537);
and U2305 (N_2305,N_1590,N_1705);
nand U2306 (N_2306,N_1737,N_1755);
nand U2307 (N_2307,N_1602,N_1779);
or U2308 (N_2308,N_1927,N_1779);
or U2309 (N_2309,N_1991,N_1978);
and U2310 (N_2310,N_1880,N_1798);
or U2311 (N_2311,N_1748,N_1730);
nand U2312 (N_2312,N_1570,N_1905);
and U2313 (N_2313,N_1682,N_1993);
and U2314 (N_2314,N_1941,N_1924);
nand U2315 (N_2315,N_1622,N_1571);
nor U2316 (N_2316,N_1550,N_1699);
and U2317 (N_2317,N_1785,N_1996);
or U2318 (N_2318,N_1816,N_1925);
nand U2319 (N_2319,N_1839,N_1878);
and U2320 (N_2320,N_1525,N_1924);
and U2321 (N_2321,N_1647,N_1754);
xnor U2322 (N_2322,N_1641,N_1806);
or U2323 (N_2323,N_1761,N_1573);
and U2324 (N_2324,N_1538,N_1595);
or U2325 (N_2325,N_1945,N_1985);
and U2326 (N_2326,N_1882,N_1671);
and U2327 (N_2327,N_1663,N_1791);
or U2328 (N_2328,N_1829,N_1689);
or U2329 (N_2329,N_1666,N_1703);
nand U2330 (N_2330,N_1819,N_1889);
and U2331 (N_2331,N_1738,N_1655);
nor U2332 (N_2332,N_1536,N_1542);
nand U2333 (N_2333,N_1571,N_1569);
nand U2334 (N_2334,N_1602,N_1901);
nor U2335 (N_2335,N_1622,N_1891);
nand U2336 (N_2336,N_1573,N_1688);
nor U2337 (N_2337,N_1516,N_1676);
or U2338 (N_2338,N_1673,N_1792);
nor U2339 (N_2339,N_1644,N_1805);
nand U2340 (N_2340,N_1730,N_1526);
or U2341 (N_2341,N_1619,N_1837);
nand U2342 (N_2342,N_1701,N_1802);
or U2343 (N_2343,N_1829,N_1603);
nor U2344 (N_2344,N_1805,N_1647);
or U2345 (N_2345,N_1830,N_1910);
and U2346 (N_2346,N_1668,N_1970);
and U2347 (N_2347,N_1503,N_1567);
or U2348 (N_2348,N_1808,N_1891);
nor U2349 (N_2349,N_1626,N_1786);
nand U2350 (N_2350,N_1994,N_1704);
or U2351 (N_2351,N_1707,N_1648);
nor U2352 (N_2352,N_1657,N_1836);
nand U2353 (N_2353,N_1546,N_1810);
or U2354 (N_2354,N_1926,N_1747);
and U2355 (N_2355,N_1741,N_1745);
and U2356 (N_2356,N_1870,N_1896);
or U2357 (N_2357,N_1986,N_1504);
or U2358 (N_2358,N_1721,N_1601);
or U2359 (N_2359,N_1727,N_1959);
nor U2360 (N_2360,N_1565,N_1608);
nor U2361 (N_2361,N_1546,N_1878);
nor U2362 (N_2362,N_1973,N_1873);
and U2363 (N_2363,N_1885,N_1943);
nor U2364 (N_2364,N_1634,N_1635);
and U2365 (N_2365,N_1561,N_1886);
nor U2366 (N_2366,N_1646,N_1825);
and U2367 (N_2367,N_1545,N_1801);
or U2368 (N_2368,N_1914,N_1939);
nand U2369 (N_2369,N_1882,N_1568);
nor U2370 (N_2370,N_1623,N_1870);
nand U2371 (N_2371,N_1877,N_1739);
nor U2372 (N_2372,N_1639,N_1978);
and U2373 (N_2373,N_1899,N_1517);
and U2374 (N_2374,N_1943,N_1993);
or U2375 (N_2375,N_1781,N_1944);
nor U2376 (N_2376,N_1966,N_1563);
and U2377 (N_2377,N_1574,N_1960);
and U2378 (N_2378,N_1735,N_1921);
nor U2379 (N_2379,N_1593,N_1976);
nand U2380 (N_2380,N_1521,N_1654);
nand U2381 (N_2381,N_1578,N_1942);
nand U2382 (N_2382,N_1907,N_1715);
nand U2383 (N_2383,N_1600,N_1857);
or U2384 (N_2384,N_1601,N_1671);
or U2385 (N_2385,N_1995,N_1979);
and U2386 (N_2386,N_1624,N_1594);
nor U2387 (N_2387,N_1859,N_1642);
nand U2388 (N_2388,N_1597,N_1815);
or U2389 (N_2389,N_1725,N_1890);
and U2390 (N_2390,N_1736,N_1905);
and U2391 (N_2391,N_1590,N_1980);
or U2392 (N_2392,N_1937,N_1637);
nor U2393 (N_2393,N_1802,N_1770);
nor U2394 (N_2394,N_1629,N_1941);
nand U2395 (N_2395,N_1784,N_1635);
and U2396 (N_2396,N_1596,N_1648);
nand U2397 (N_2397,N_1593,N_1916);
nor U2398 (N_2398,N_1522,N_1754);
nor U2399 (N_2399,N_1779,N_1957);
or U2400 (N_2400,N_1722,N_1921);
or U2401 (N_2401,N_1972,N_1532);
nor U2402 (N_2402,N_1716,N_1755);
and U2403 (N_2403,N_1676,N_1936);
nand U2404 (N_2404,N_1650,N_1978);
nand U2405 (N_2405,N_1935,N_1512);
or U2406 (N_2406,N_1740,N_1744);
and U2407 (N_2407,N_1674,N_1660);
nand U2408 (N_2408,N_1764,N_1530);
nor U2409 (N_2409,N_1737,N_1954);
or U2410 (N_2410,N_1918,N_1683);
or U2411 (N_2411,N_1826,N_1968);
nand U2412 (N_2412,N_1953,N_1698);
or U2413 (N_2413,N_1996,N_1570);
nor U2414 (N_2414,N_1646,N_1880);
and U2415 (N_2415,N_1595,N_1500);
nand U2416 (N_2416,N_1708,N_1800);
nand U2417 (N_2417,N_1875,N_1728);
nor U2418 (N_2418,N_1730,N_1963);
nor U2419 (N_2419,N_1658,N_1768);
or U2420 (N_2420,N_1542,N_1758);
nor U2421 (N_2421,N_1893,N_1522);
nor U2422 (N_2422,N_1532,N_1976);
xor U2423 (N_2423,N_1805,N_1940);
and U2424 (N_2424,N_1810,N_1803);
or U2425 (N_2425,N_1809,N_1904);
nand U2426 (N_2426,N_1755,N_1601);
nor U2427 (N_2427,N_1593,N_1984);
or U2428 (N_2428,N_1869,N_1726);
or U2429 (N_2429,N_1536,N_1965);
and U2430 (N_2430,N_1939,N_1548);
or U2431 (N_2431,N_1561,N_1879);
or U2432 (N_2432,N_1673,N_1765);
nand U2433 (N_2433,N_1775,N_1923);
and U2434 (N_2434,N_1521,N_1579);
xnor U2435 (N_2435,N_1802,N_1539);
or U2436 (N_2436,N_1981,N_1633);
nand U2437 (N_2437,N_1567,N_1713);
nor U2438 (N_2438,N_1655,N_1636);
and U2439 (N_2439,N_1511,N_1676);
and U2440 (N_2440,N_1551,N_1915);
or U2441 (N_2441,N_1757,N_1527);
and U2442 (N_2442,N_1935,N_1966);
and U2443 (N_2443,N_1844,N_1809);
nor U2444 (N_2444,N_1526,N_1797);
and U2445 (N_2445,N_1774,N_1595);
or U2446 (N_2446,N_1787,N_1526);
or U2447 (N_2447,N_1662,N_1800);
or U2448 (N_2448,N_1606,N_1817);
nor U2449 (N_2449,N_1945,N_1634);
or U2450 (N_2450,N_1647,N_1556);
or U2451 (N_2451,N_1685,N_1760);
and U2452 (N_2452,N_1544,N_1584);
and U2453 (N_2453,N_1567,N_1988);
nor U2454 (N_2454,N_1875,N_1791);
nor U2455 (N_2455,N_1797,N_1582);
or U2456 (N_2456,N_1695,N_1646);
or U2457 (N_2457,N_1955,N_1966);
nor U2458 (N_2458,N_1755,N_1731);
xnor U2459 (N_2459,N_1902,N_1893);
and U2460 (N_2460,N_1854,N_1881);
and U2461 (N_2461,N_1898,N_1949);
and U2462 (N_2462,N_1607,N_1652);
or U2463 (N_2463,N_1923,N_1902);
nor U2464 (N_2464,N_1910,N_1590);
or U2465 (N_2465,N_1600,N_1888);
nand U2466 (N_2466,N_1555,N_1780);
nor U2467 (N_2467,N_1766,N_1578);
nand U2468 (N_2468,N_1860,N_1790);
and U2469 (N_2469,N_1773,N_1563);
nand U2470 (N_2470,N_1826,N_1745);
nand U2471 (N_2471,N_1863,N_1742);
and U2472 (N_2472,N_1681,N_1920);
and U2473 (N_2473,N_1522,N_1911);
or U2474 (N_2474,N_1511,N_1526);
and U2475 (N_2475,N_1962,N_1849);
nand U2476 (N_2476,N_1691,N_1962);
nor U2477 (N_2477,N_1989,N_1829);
nor U2478 (N_2478,N_1540,N_1947);
and U2479 (N_2479,N_1793,N_1800);
nor U2480 (N_2480,N_1882,N_1844);
nand U2481 (N_2481,N_1694,N_1794);
and U2482 (N_2482,N_1722,N_1500);
and U2483 (N_2483,N_1683,N_1934);
or U2484 (N_2484,N_1774,N_1701);
nand U2485 (N_2485,N_1568,N_1825);
nand U2486 (N_2486,N_1681,N_1646);
or U2487 (N_2487,N_1736,N_1829);
nor U2488 (N_2488,N_1809,N_1643);
and U2489 (N_2489,N_1637,N_1796);
nand U2490 (N_2490,N_1980,N_1513);
nor U2491 (N_2491,N_1929,N_1635);
nand U2492 (N_2492,N_1967,N_1569);
or U2493 (N_2493,N_1876,N_1548);
nand U2494 (N_2494,N_1931,N_1776);
or U2495 (N_2495,N_1950,N_1620);
nor U2496 (N_2496,N_1724,N_1631);
and U2497 (N_2497,N_1756,N_1934);
nand U2498 (N_2498,N_1891,N_1892);
or U2499 (N_2499,N_1965,N_1812);
nor U2500 (N_2500,N_2111,N_2162);
and U2501 (N_2501,N_2453,N_2201);
nor U2502 (N_2502,N_2418,N_2362);
nand U2503 (N_2503,N_2285,N_2126);
or U2504 (N_2504,N_2323,N_2032);
and U2505 (N_2505,N_2460,N_2397);
nand U2506 (N_2506,N_2328,N_2202);
or U2507 (N_2507,N_2245,N_2449);
or U2508 (N_2508,N_2193,N_2273);
and U2509 (N_2509,N_2342,N_2015);
nor U2510 (N_2510,N_2174,N_2478);
or U2511 (N_2511,N_2334,N_2167);
or U2512 (N_2512,N_2425,N_2263);
nor U2513 (N_2513,N_2026,N_2219);
nor U2514 (N_2514,N_2114,N_2001);
and U2515 (N_2515,N_2420,N_2288);
or U2516 (N_2516,N_2214,N_2246);
nand U2517 (N_2517,N_2172,N_2042);
or U2518 (N_2518,N_2030,N_2311);
or U2519 (N_2519,N_2255,N_2447);
nor U2520 (N_2520,N_2081,N_2499);
and U2521 (N_2521,N_2356,N_2325);
or U2522 (N_2522,N_2095,N_2475);
and U2523 (N_2523,N_2127,N_2474);
or U2524 (N_2524,N_2261,N_2016);
nand U2525 (N_2525,N_2140,N_2266);
nor U2526 (N_2526,N_2437,N_2170);
nor U2527 (N_2527,N_2105,N_2180);
nand U2528 (N_2528,N_2443,N_2231);
or U2529 (N_2529,N_2380,N_2086);
nand U2530 (N_2530,N_2476,N_2317);
nor U2531 (N_2531,N_2054,N_2045);
or U2532 (N_2532,N_2074,N_2448);
and U2533 (N_2533,N_2454,N_2213);
nand U2534 (N_2534,N_2291,N_2358);
nand U2535 (N_2535,N_2403,N_2368);
and U2536 (N_2536,N_2239,N_2367);
nand U2537 (N_2537,N_2057,N_2484);
nand U2538 (N_2538,N_2135,N_2248);
nor U2539 (N_2539,N_2050,N_2413);
nand U2540 (N_2540,N_2154,N_2371);
and U2541 (N_2541,N_2190,N_2148);
and U2542 (N_2542,N_2345,N_2034);
or U2543 (N_2543,N_2068,N_2136);
or U2544 (N_2544,N_2428,N_2277);
or U2545 (N_2545,N_2299,N_2468);
and U2546 (N_2546,N_2477,N_2459);
nand U2547 (N_2547,N_2071,N_2028);
nand U2548 (N_2548,N_2194,N_2061);
xor U2549 (N_2549,N_2179,N_2287);
and U2550 (N_2550,N_2452,N_2008);
nor U2551 (N_2551,N_2142,N_2218);
nor U2552 (N_2552,N_2377,N_2432);
nand U2553 (N_2553,N_2365,N_2326);
and U2554 (N_2554,N_2318,N_2336);
and U2555 (N_2555,N_2217,N_2196);
nor U2556 (N_2556,N_2348,N_2346);
nor U2557 (N_2557,N_2364,N_2108);
nand U2558 (N_2558,N_2143,N_2150);
and U2559 (N_2559,N_2085,N_2049);
nor U2560 (N_2560,N_2441,N_2004);
nand U2561 (N_2561,N_2215,N_2024);
nor U2562 (N_2562,N_2269,N_2464);
or U2563 (N_2563,N_2315,N_2404);
nor U2564 (N_2564,N_2019,N_2455);
nand U2565 (N_2565,N_2394,N_2153);
nor U2566 (N_2566,N_2234,N_2000);
or U2567 (N_2567,N_2075,N_2379);
or U2568 (N_2568,N_2097,N_2298);
nor U2569 (N_2569,N_2438,N_2178);
or U2570 (N_2570,N_2304,N_2253);
nor U2571 (N_2571,N_2274,N_2184);
and U2572 (N_2572,N_2416,N_2144);
nor U2573 (N_2573,N_2243,N_2103);
nand U2574 (N_2574,N_2374,N_2470);
or U2575 (N_2575,N_2165,N_2372);
nor U2576 (N_2576,N_2055,N_2237);
and U2577 (N_2577,N_2440,N_2270);
or U2578 (N_2578,N_2417,N_2396);
nor U2579 (N_2579,N_2122,N_2225);
nand U2580 (N_2580,N_2017,N_2233);
nor U2581 (N_2581,N_2181,N_2493);
nor U2582 (N_2582,N_2436,N_2080);
or U2583 (N_2583,N_2496,N_2435);
nand U2584 (N_2584,N_2360,N_2433);
nand U2585 (N_2585,N_2350,N_2262);
nand U2586 (N_2586,N_2164,N_2079);
and U2587 (N_2587,N_2092,N_2301);
nor U2588 (N_2588,N_2244,N_2232);
nor U2589 (N_2589,N_2195,N_2398);
and U2590 (N_2590,N_2044,N_2223);
nor U2591 (N_2591,N_2241,N_2145);
and U2592 (N_2592,N_2098,N_2275);
or U2593 (N_2593,N_2087,N_2296);
and U2594 (N_2594,N_2006,N_2236);
nor U2595 (N_2595,N_2444,N_2387);
nand U2596 (N_2596,N_2056,N_2163);
or U2597 (N_2597,N_2469,N_2330);
or U2598 (N_2598,N_2324,N_2102);
nand U2599 (N_2599,N_2258,N_2012);
and U2600 (N_2600,N_2070,N_2113);
xor U2601 (N_2601,N_2267,N_2156);
nand U2602 (N_2602,N_2088,N_2109);
and U2603 (N_2603,N_2395,N_2300);
nor U2604 (N_2604,N_2216,N_2212);
or U2605 (N_2605,N_2322,N_2158);
and U2606 (N_2606,N_2106,N_2199);
or U2607 (N_2607,N_2307,N_2278);
nand U2608 (N_2608,N_2421,N_2058);
and U2609 (N_2609,N_2490,N_2497);
nor U2610 (N_2610,N_2466,N_2339);
nor U2611 (N_2611,N_2222,N_2128);
and U2612 (N_2612,N_2383,N_2405);
nand U2613 (N_2613,N_2036,N_2419);
nand U2614 (N_2614,N_2207,N_2110);
and U2615 (N_2615,N_2066,N_2283);
nor U2616 (N_2616,N_2333,N_2189);
nor U2617 (N_2617,N_2047,N_2238);
or U2618 (N_2618,N_2250,N_2009);
nor U2619 (N_2619,N_2020,N_2121);
or U2620 (N_2620,N_2227,N_2073);
nor U2621 (N_2621,N_2224,N_2046);
nand U2622 (N_2622,N_2359,N_2002);
nor U2623 (N_2623,N_2187,N_2228);
and U2624 (N_2624,N_2256,N_2293);
or U2625 (N_2625,N_2072,N_2198);
nor U2626 (N_2626,N_2200,N_2076);
or U2627 (N_2627,N_2221,N_2369);
nand U2628 (N_2628,N_2146,N_2445);
nand U2629 (N_2629,N_2063,N_2132);
and U2630 (N_2630,N_2041,N_2357);
and U2631 (N_2631,N_2492,N_2467);
nor U2632 (N_2632,N_2251,N_2343);
nand U2633 (N_2633,N_2119,N_2320);
or U2634 (N_2634,N_2118,N_2029);
xnor U2635 (N_2635,N_2259,N_2062);
nand U2636 (N_2636,N_2276,N_2309);
or U2637 (N_2637,N_2147,N_2295);
nor U2638 (N_2638,N_2176,N_2314);
or U2639 (N_2639,N_2099,N_2264);
and U2640 (N_2640,N_2023,N_2129);
nand U2641 (N_2641,N_2382,N_2053);
nor U2642 (N_2642,N_2352,N_2185);
or U2643 (N_2643,N_2037,N_2204);
nor U2644 (N_2644,N_2462,N_2117);
or U2645 (N_2645,N_2077,N_2282);
or U2646 (N_2646,N_2473,N_2465);
or U2647 (N_2647,N_2409,N_2060);
or U2648 (N_2648,N_2220,N_2388);
xnor U2649 (N_2649,N_2399,N_2093);
and U2650 (N_2650,N_2271,N_2089);
and U2651 (N_2651,N_2321,N_2337);
nand U2652 (N_2652,N_2386,N_2412);
nand U2653 (N_2653,N_2033,N_2434);
nor U2654 (N_2654,N_2123,N_2480);
nand U2655 (N_2655,N_2151,N_2485);
or U2656 (N_2656,N_2188,N_2354);
nand U2657 (N_2657,N_2229,N_2010);
nor U2658 (N_2658,N_2115,N_2400);
nor U2659 (N_2659,N_2373,N_2491);
nand U2660 (N_2660,N_2384,N_2082);
nand U2661 (N_2661,N_2391,N_2302);
or U2662 (N_2662,N_2206,N_2494);
nor U2663 (N_2663,N_2422,N_2192);
nand U2664 (N_2664,N_2442,N_2332);
nand U2665 (N_2665,N_2393,N_2280);
nand U2666 (N_2666,N_2303,N_2257);
or U2667 (N_2667,N_2451,N_2096);
nor U2668 (N_2668,N_2025,N_2402);
nor U2669 (N_2669,N_2335,N_2363);
nor U2670 (N_2670,N_2414,N_2240);
or U2671 (N_2671,N_2078,N_2160);
nor U2672 (N_2672,N_2308,N_2101);
nand U2673 (N_2673,N_2408,N_2039);
nand U2674 (N_2674,N_2249,N_2112);
or U2675 (N_2675,N_2166,N_2366);
and U2676 (N_2676,N_2120,N_2031);
or U2677 (N_2677,N_2430,N_2131);
nor U2678 (N_2678,N_2427,N_2272);
and U2679 (N_2679,N_2489,N_2247);
and U2680 (N_2680,N_2027,N_2313);
and U2681 (N_2681,N_2084,N_2035);
or U2682 (N_2682,N_2059,N_2392);
or U2683 (N_2683,N_2139,N_2171);
nor U2684 (N_2684,N_2268,N_2355);
and U2685 (N_2685,N_2439,N_2124);
and U2686 (N_2686,N_2498,N_2292);
and U2687 (N_2687,N_2390,N_2381);
nor U2688 (N_2688,N_2411,N_2310);
or U2689 (N_2689,N_2294,N_2137);
or U2690 (N_2690,N_2327,N_2107);
or U2691 (N_2691,N_2007,N_2173);
and U2692 (N_2692,N_2265,N_2378);
nor U2693 (N_2693,N_2094,N_2083);
nand U2694 (N_2694,N_2209,N_2457);
and U2695 (N_2695,N_2260,N_2479);
and U2696 (N_2696,N_2289,N_2340);
or U2697 (N_2697,N_2091,N_2067);
nor U2698 (N_2698,N_2021,N_2018);
or U2699 (N_2699,N_2252,N_2149);
nor U2700 (N_2700,N_2279,N_2487);
nand U2701 (N_2701,N_2203,N_2456);
nor U2702 (N_2702,N_2370,N_2306);
and U2703 (N_2703,N_2011,N_2483);
and U2704 (N_2704,N_2090,N_2461);
nor U2705 (N_2705,N_2116,N_2242);
nor U2706 (N_2706,N_2048,N_2152);
nor U2707 (N_2707,N_2161,N_2488);
and U2708 (N_2708,N_2022,N_2191);
nor U2709 (N_2709,N_2375,N_2472);
or U2710 (N_2710,N_2155,N_2312);
nor U2711 (N_2711,N_2186,N_2141);
nor U2712 (N_2712,N_2407,N_2481);
and U2713 (N_2713,N_2254,N_2401);
or U2714 (N_2714,N_2423,N_2351);
nand U2715 (N_2715,N_2065,N_2226);
or U2716 (N_2716,N_2347,N_2415);
nand U2717 (N_2717,N_2389,N_2424);
nor U2718 (N_2718,N_2344,N_2486);
nor U2719 (N_2719,N_2406,N_2329);
and U2720 (N_2720,N_2205,N_2175);
nor U2721 (N_2721,N_2177,N_2446);
and U2722 (N_2722,N_2211,N_2230);
nand U2723 (N_2723,N_2104,N_2331);
and U2724 (N_2724,N_2138,N_2431);
nand U2725 (N_2725,N_2130,N_2471);
and U2726 (N_2726,N_2005,N_2014);
and U2727 (N_2727,N_2003,N_2361);
nand U2728 (N_2728,N_2286,N_2183);
and U2729 (N_2729,N_2168,N_2182);
nand U2730 (N_2730,N_2341,N_2038);
or U2731 (N_2731,N_2210,N_2064);
and U2732 (N_2732,N_2235,N_2316);
and U2733 (N_2733,N_2134,N_2281);
nor U2734 (N_2734,N_2429,N_2169);
or U2735 (N_2735,N_2100,N_2450);
nand U2736 (N_2736,N_2013,N_2069);
or U2737 (N_2737,N_2208,N_2159);
and U2738 (N_2738,N_2284,N_2305);
and U2739 (N_2739,N_2482,N_2052);
nand U2740 (N_2740,N_2197,N_2157);
and U2741 (N_2741,N_2290,N_2043);
or U2742 (N_2742,N_2410,N_2426);
nand U2743 (N_2743,N_2463,N_2040);
nor U2744 (N_2744,N_2376,N_2349);
or U2745 (N_2745,N_2051,N_2385);
nand U2746 (N_2746,N_2338,N_2458);
and U2747 (N_2747,N_2125,N_2297);
or U2748 (N_2748,N_2353,N_2133);
nor U2749 (N_2749,N_2495,N_2319);
nor U2750 (N_2750,N_2102,N_2449);
and U2751 (N_2751,N_2087,N_2044);
nor U2752 (N_2752,N_2142,N_2293);
nor U2753 (N_2753,N_2353,N_2226);
and U2754 (N_2754,N_2245,N_2028);
and U2755 (N_2755,N_2323,N_2313);
nor U2756 (N_2756,N_2477,N_2264);
and U2757 (N_2757,N_2385,N_2090);
nor U2758 (N_2758,N_2279,N_2366);
or U2759 (N_2759,N_2324,N_2325);
nor U2760 (N_2760,N_2493,N_2444);
nor U2761 (N_2761,N_2427,N_2349);
and U2762 (N_2762,N_2119,N_2367);
nand U2763 (N_2763,N_2293,N_2344);
or U2764 (N_2764,N_2275,N_2040);
nor U2765 (N_2765,N_2012,N_2273);
and U2766 (N_2766,N_2064,N_2437);
or U2767 (N_2767,N_2132,N_2474);
and U2768 (N_2768,N_2457,N_2375);
and U2769 (N_2769,N_2108,N_2449);
nand U2770 (N_2770,N_2400,N_2287);
and U2771 (N_2771,N_2427,N_2133);
nor U2772 (N_2772,N_2025,N_2362);
and U2773 (N_2773,N_2040,N_2424);
nor U2774 (N_2774,N_2488,N_2119);
nor U2775 (N_2775,N_2411,N_2379);
or U2776 (N_2776,N_2110,N_2000);
nor U2777 (N_2777,N_2265,N_2122);
nand U2778 (N_2778,N_2288,N_2374);
and U2779 (N_2779,N_2356,N_2495);
nand U2780 (N_2780,N_2101,N_2473);
nand U2781 (N_2781,N_2239,N_2253);
and U2782 (N_2782,N_2431,N_2457);
nor U2783 (N_2783,N_2072,N_2335);
nand U2784 (N_2784,N_2162,N_2446);
nand U2785 (N_2785,N_2118,N_2379);
nor U2786 (N_2786,N_2204,N_2214);
xnor U2787 (N_2787,N_2177,N_2435);
nand U2788 (N_2788,N_2037,N_2472);
or U2789 (N_2789,N_2444,N_2447);
nor U2790 (N_2790,N_2204,N_2316);
nand U2791 (N_2791,N_2172,N_2461);
nand U2792 (N_2792,N_2392,N_2147);
and U2793 (N_2793,N_2353,N_2265);
or U2794 (N_2794,N_2429,N_2499);
nor U2795 (N_2795,N_2339,N_2048);
nand U2796 (N_2796,N_2462,N_2324);
nor U2797 (N_2797,N_2025,N_2404);
nor U2798 (N_2798,N_2227,N_2275);
nor U2799 (N_2799,N_2292,N_2019);
and U2800 (N_2800,N_2122,N_2066);
or U2801 (N_2801,N_2233,N_2164);
nand U2802 (N_2802,N_2419,N_2260);
and U2803 (N_2803,N_2153,N_2025);
or U2804 (N_2804,N_2454,N_2499);
nand U2805 (N_2805,N_2138,N_2238);
nand U2806 (N_2806,N_2026,N_2260);
or U2807 (N_2807,N_2332,N_2148);
nor U2808 (N_2808,N_2082,N_2070);
or U2809 (N_2809,N_2420,N_2188);
nor U2810 (N_2810,N_2403,N_2105);
nor U2811 (N_2811,N_2021,N_2301);
nand U2812 (N_2812,N_2019,N_2160);
nand U2813 (N_2813,N_2032,N_2322);
or U2814 (N_2814,N_2166,N_2104);
nor U2815 (N_2815,N_2168,N_2459);
and U2816 (N_2816,N_2313,N_2436);
nor U2817 (N_2817,N_2078,N_2124);
nor U2818 (N_2818,N_2006,N_2256);
or U2819 (N_2819,N_2361,N_2075);
and U2820 (N_2820,N_2041,N_2246);
or U2821 (N_2821,N_2063,N_2054);
or U2822 (N_2822,N_2389,N_2056);
and U2823 (N_2823,N_2399,N_2360);
and U2824 (N_2824,N_2171,N_2117);
nor U2825 (N_2825,N_2218,N_2253);
nand U2826 (N_2826,N_2137,N_2234);
or U2827 (N_2827,N_2183,N_2066);
nand U2828 (N_2828,N_2471,N_2040);
or U2829 (N_2829,N_2196,N_2094);
nand U2830 (N_2830,N_2451,N_2393);
xnor U2831 (N_2831,N_2124,N_2289);
or U2832 (N_2832,N_2422,N_2172);
and U2833 (N_2833,N_2113,N_2448);
or U2834 (N_2834,N_2283,N_2485);
nor U2835 (N_2835,N_2347,N_2362);
and U2836 (N_2836,N_2195,N_2415);
or U2837 (N_2837,N_2057,N_2046);
nand U2838 (N_2838,N_2413,N_2037);
and U2839 (N_2839,N_2185,N_2046);
nand U2840 (N_2840,N_2204,N_2104);
nand U2841 (N_2841,N_2408,N_2457);
nand U2842 (N_2842,N_2168,N_2209);
or U2843 (N_2843,N_2122,N_2291);
or U2844 (N_2844,N_2226,N_2258);
or U2845 (N_2845,N_2364,N_2467);
or U2846 (N_2846,N_2239,N_2046);
nor U2847 (N_2847,N_2043,N_2446);
or U2848 (N_2848,N_2494,N_2254);
nand U2849 (N_2849,N_2133,N_2364);
nor U2850 (N_2850,N_2058,N_2410);
nand U2851 (N_2851,N_2064,N_2306);
nor U2852 (N_2852,N_2392,N_2050);
nor U2853 (N_2853,N_2014,N_2242);
and U2854 (N_2854,N_2148,N_2418);
or U2855 (N_2855,N_2009,N_2476);
nor U2856 (N_2856,N_2271,N_2013);
or U2857 (N_2857,N_2219,N_2126);
or U2858 (N_2858,N_2020,N_2157);
nand U2859 (N_2859,N_2033,N_2374);
nand U2860 (N_2860,N_2495,N_2005);
and U2861 (N_2861,N_2040,N_2279);
and U2862 (N_2862,N_2172,N_2238);
and U2863 (N_2863,N_2091,N_2344);
nor U2864 (N_2864,N_2102,N_2117);
nand U2865 (N_2865,N_2218,N_2041);
nor U2866 (N_2866,N_2252,N_2230);
or U2867 (N_2867,N_2224,N_2097);
and U2868 (N_2868,N_2403,N_2494);
and U2869 (N_2869,N_2463,N_2331);
or U2870 (N_2870,N_2176,N_2306);
or U2871 (N_2871,N_2410,N_2049);
and U2872 (N_2872,N_2223,N_2302);
nand U2873 (N_2873,N_2081,N_2162);
nand U2874 (N_2874,N_2110,N_2229);
or U2875 (N_2875,N_2498,N_2181);
and U2876 (N_2876,N_2000,N_2089);
nand U2877 (N_2877,N_2377,N_2305);
nand U2878 (N_2878,N_2266,N_2399);
nand U2879 (N_2879,N_2045,N_2038);
or U2880 (N_2880,N_2027,N_2417);
xnor U2881 (N_2881,N_2210,N_2083);
nor U2882 (N_2882,N_2015,N_2205);
and U2883 (N_2883,N_2032,N_2414);
nand U2884 (N_2884,N_2368,N_2099);
nand U2885 (N_2885,N_2386,N_2200);
or U2886 (N_2886,N_2377,N_2453);
xor U2887 (N_2887,N_2380,N_2051);
and U2888 (N_2888,N_2312,N_2364);
nand U2889 (N_2889,N_2358,N_2287);
or U2890 (N_2890,N_2113,N_2383);
nand U2891 (N_2891,N_2402,N_2412);
nand U2892 (N_2892,N_2028,N_2145);
nor U2893 (N_2893,N_2354,N_2256);
nor U2894 (N_2894,N_2423,N_2137);
or U2895 (N_2895,N_2352,N_2126);
or U2896 (N_2896,N_2033,N_2342);
and U2897 (N_2897,N_2077,N_2095);
nor U2898 (N_2898,N_2483,N_2311);
or U2899 (N_2899,N_2406,N_2354);
and U2900 (N_2900,N_2405,N_2020);
nor U2901 (N_2901,N_2435,N_2323);
or U2902 (N_2902,N_2393,N_2299);
and U2903 (N_2903,N_2140,N_2118);
and U2904 (N_2904,N_2293,N_2023);
and U2905 (N_2905,N_2360,N_2081);
nor U2906 (N_2906,N_2357,N_2355);
and U2907 (N_2907,N_2150,N_2402);
nor U2908 (N_2908,N_2088,N_2235);
nand U2909 (N_2909,N_2295,N_2090);
and U2910 (N_2910,N_2310,N_2071);
or U2911 (N_2911,N_2210,N_2295);
nand U2912 (N_2912,N_2231,N_2361);
nor U2913 (N_2913,N_2484,N_2098);
and U2914 (N_2914,N_2323,N_2049);
and U2915 (N_2915,N_2009,N_2429);
nand U2916 (N_2916,N_2062,N_2068);
nor U2917 (N_2917,N_2396,N_2356);
and U2918 (N_2918,N_2251,N_2439);
or U2919 (N_2919,N_2215,N_2413);
or U2920 (N_2920,N_2358,N_2411);
nand U2921 (N_2921,N_2244,N_2251);
and U2922 (N_2922,N_2364,N_2470);
and U2923 (N_2923,N_2126,N_2308);
nand U2924 (N_2924,N_2386,N_2343);
nor U2925 (N_2925,N_2008,N_2283);
or U2926 (N_2926,N_2060,N_2145);
nand U2927 (N_2927,N_2114,N_2299);
and U2928 (N_2928,N_2015,N_2378);
and U2929 (N_2929,N_2420,N_2308);
and U2930 (N_2930,N_2478,N_2257);
or U2931 (N_2931,N_2237,N_2222);
nor U2932 (N_2932,N_2203,N_2472);
and U2933 (N_2933,N_2153,N_2077);
or U2934 (N_2934,N_2282,N_2062);
nor U2935 (N_2935,N_2022,N_2308);
and U2936 (N_2936,N_2430,N_2037);
and U2937 (N_2937,N_2041,N_2135);
nand U2938 (N_2938,N_2244,N_2473);
or U2939 (N_2939,N_2036,N_2174);
or U2940 (N_2940,N_2326,N_2080);
or U2941 (N_2941,N_2172,N_2406);
nand U2942 (N_2942,N_2297,N_2149);
nor U2943 (N_2943,N_2497,N_2347);
nand U2944 (N_2944,N_2242,N_2073);
or U2945 (N_2945,N_2251,N_2200);
or U2946 (N_2946,N_2036,N_2392);
nor U2947 (N_2947,N_2349,N_2227);
and U2948 (N_2948,N_2269,N_2372);
or U2949 (N_2949,N_2162,N_2379);
nand U2950 (N_2950,N_2210,N_2224);
nor U2951 (N_2951,N_2182,N_2443);
or U2952 (N_2952,N_2020,N_2453);
nor U2953 (N_2953,N_2266,N_2204);
and U2954 (N_2954,N_2387,N_2376);
and U2955 (N_2955,N_2480,N_2371);
or U2956 (N_2956,N_2372,N_2332);
nor U2957 (N_2957,N_2370,N_2221);
nor U2958 (N_2958,N_2181,N_2454);
nand U2959 (N_2959,N_2026,N_2044);
nand U2960 (N_2960,N_2448,N_2433);
or U2961 (N_2961,N_2322,N_2090);
nor U2962 (N_2962,N_2470,N_2315);
nor U2963 (N_2963,N_2366,N_2039);
nor U2964 (N_2964,N_2319,N_2493);
nand U2965 (N_2965,N_2233,N_2107);
nor U2966 (N_2966,N_2068,N_2381);
nor U2967 (N_2967,N_2277,N_2243);
and U2968 (N_2968,N_2263,N_2089);
nand U2969 (N_2969,N_2178,N_2333);
or U2970 (N_2970,N_2438,N_2289);
and U2971 (N_2971,N_2405,N_2485);
and U2972 (N_2972,N_2363,N_2320);
nand U2973 (N_2973,N_2111,N_2059);
nand U2974 (N_2974,N_2344,N_2345);
nor U2975 (N_2975,N_2208,N_2277);
and U2976 (N_2976,N_2308,N_2070);
nand U2977 (N_2977,N_2189,N_2476);
and U2978 (N_2978,N_2413,N_2174);
or U2979 (N_2979,N_2148,N_2059);
nand U2980 (N_2980,N_2172,N_2168);
nor U2981 (N_2981,N_2237,N_2009);
and U2982 (N_2982,N_2108,N_2075);
or U2983 (N_2983,N_2052,N_2298);
nand U2984 (N_2984,N_2209,N_2440);
or U2985 (N_2985,N_2157,N_2200);
and U2986 (N_2986,N_2065,N_2297);
nor U2987 (N_2987,N_2291,N_2130);
or U2988 (N_2988,N_2153,N_2285);
or U2989 (N_2989,N_2454,N_2251);
or U2990 (N_2990,N_2046,N_2012);
and U2991 (N_2991,N_2073,N_2205);
nand U2992 (N_2992,N_2197,N_2499);
nor U2993 (N_2993,N_2388,N_2298);
or U2994 (N_2994,N_2185,N_2005);
nand U2995 (N_2995,N_2344,N_2329);
nor U2996 (N_2996,N_2257,N_2234);
or U2997 (N_2997,N_2085,N_2115);
nand U2998 (N_2998,N_2082,N_2350);
or U2999 (N_2999,N_2175,N_2484);
or UO_0 (O_0,N_2746,N_2658);
xnor UO_1 (O_1,N_2888,N_2563);
nor UO_2 (O_2,N_2649,N_2812);
and UO_3 (O_3,N_2700,N_2808);
nor UO_4 (O_4,N_2854,N_2532);
xor UO_5 (O_5,N_2573,N_2687);
nand UO_6 (O_6,N_2823,N_2694);
and UO_7 (O_7,N_2980,N_2741);
nand UO_8 (O_8,N_2972,N_2776);
nand UO_9 (O_9,N_2765,N_2558);
or UO_10 (O_10,N_2851,N_2511);
nor UO_11 (O_11,N_2908,N_2653);
nor UO_12 (O_12,N_2946,N_2677);
nor UO_13 (O_13,N_2860,N_2736);
or UO_14 (O_14,N_2531,N_2766);
or UO_15 (O_15,N_2883,N_2685);
or UO_16 (O_16,N_2600,N_2764);
or UO_17 (O_17,N_2698,N_2757);
or UO_18 (O_18,N_2804,N_2767);
nand UO_19 (O_19,N_2996,N_2753);
nand UO_20 (O_20,N_2551,N_2556);
nand UO_21 (O_21,N_2831,N_2589);
nor UO_22 (O_22,N_2948,N_2936);
or UO_23 (O_23,N_2749,N_2599);
and UO_24 (O_24,N_2582,N_2706);
nand UO_25 (O_25,N_2622,N_2884);
nor UO_26 (O_26,N_2762,N_2528);
nand UO_27 (O_27,N_2782,N_2756);
nor UO_28 (O_28,N_2939,N_2518);
nand UO_29 (O_29,N_2843,N_2695);
and UO_30 (O_30,N_2905,N_2988);
nor UO_31 (O_31,N_2932,N_2772);
nor UO_32 (O_32,N_2886,N_2570);
nor UO_33 (O_33,N_2858,N_2543);
nand UO_34 (O_34,N_2937,N_2674);
and UO_35 (O_35,N_2805,N_2569);
nor UO_36 (O_36,N_2799,N_2775);
nor UO_37 (O_37,N_2639,N_2873);
nand UO_38 (O_38,N_2847,N_2990);
and UO_39 (O_39,N_2501,N_2703);
nand UO_40 (O_40,N_2657,N_2867);
nor UO_41 (O_41,N_2759,N_2929);
nor UO_42 (O_42,N_2548,N_2602);
or UO_43 (O_43,N_2593,N_2914);
and UO_44 (O_44,N_2739,N_2624);
nor UO_45 (O_45,N_2839,N_2862);
and UO_46 (O_46,N_2592,N_2950);
nand UO_47 (O_47,N_2568,N_2615);
nor UO_48 (O_48,N_2664,N_2953);
nor UO_49 (O_49,N_2834,N_2533);
nand UO_50 (O_50,N_2740,N_2966);
nor UO_51 (O_51,N_2688,N_2967);
or UO_52 (O_52,N_2801,N_2876);
nand UO_53 (O_53,N_2923,N_2607);
nor UO_54 (O_54,N_2806,N_2572);
and UO_55 (O_55,N_2842,N_2735);
nor UO_56 (O_56,N_2915,N_2802);
and UO_57 (O_57,N_2835,N_2961);
or UO_58 (O_58,N_2594,N_2763);
nand UO_59 (O_59,N_2933,N_2794);
nand UO_60 (O_60,N_2527,N_2822);
nand UO_61 (O_61,N_2612,N_2743);
and UO_62 (O_62,N_2913,N_2675);
and UO_63 (O_63,N_2715,N_2726);
nand UO_64 (O_64,N_2526,N_2561);
nor UO_65 (O_65,N_2720,N_2667);
nand UO_66 (O_66,N_2807,N_2796);
or UO_67 (O_67,N_2541,N_2712);
and UO_68 (O_68,N_2791,N_2960);
and UO_69 (O_69,N_2654,N_2951);
nand UO_70 (O_70,N_2676,N_2999);
nor UO_71 (O_71,N_2965,N_2985);
or UO_72 (O_72,N_2724,N_2959);
nor UO_73 (O_73,N_2719,N_2971);
nor UO_74 (O_74,N_2895,N_2663);
or UO_75 (O_75,N_2742,N_2727);
nand UO_76 (O_76,N_2689,N_2671);
nand UO_77 (O_77,N_2636,N_2737);
or UO_78 (O_78,N_2912,N_2969);
or UO_79 (O_79,N_2870,N_2829);
nand UO_80 (O_80,N_2538,N_2603);
or UO_81 (O_81,N_2513,N_2711);
or UO_82 (O_82,N_2683,N_2918);
nand UO_83 (O_83,N_2942,N_2516);
nor UO_84 (O_84,N_2717,N_2577);
nor UO_85 (O_85,N_2991,N_2745);
nor UO_86 (O_86,N_2670,N_2833);
or UO_87 (O_87,N_2872,N_2827);
nor UO_88 (O_88,N_2928,N_2809);
nor UO_89 (O_89,N_2718,N_2750);
nand UO_90 (O_90,N_2580,N_2944);
or UO_91 (O_91,N_2813,N_2557);
nand UO_92 (O_92,N_2574,N_2679);
nand UO_93 (O_93,N_2566,N_2824);
or UO_94 (O_94,N_2792,N_2828);
nor UO_95 (O_95,N_2877,N_2637);
nand UO_96 (O_96,N_2938,N_2641);
or UO_97 (O_97,N_2546,N_2856);
or UO_98 (O_98,N_2909,N_2708);
and UO_99 (O_99,N_2692,N_2705);
and UO_100 (O_100,N_2841,N_2904);
nor UO_101 (O_101,N_2869,N_2787);
nor UO_102 (O_102,N_2826,N_2690);
or UO_103 (O_103,N_2783,N_2986);
nand UO_104 (O_104,N_2571,N_2789);
or UO_105 (O_105,N_2837,N_2896);
or UO_106 (O_106,N_2553,N_2784);
nor UO_107 (O_107,N_2621,N_2963);
or UO_108 (O_108,N_2554,N_2875);
nand UO_109 (O_109,N_2924,N_2898);
nor UO_110 (O_110,N_2627,N_2604);
or UO_111 (O_111,N_2779,N_2505);
nor UO_112 (O_112,N_2633,N_2970);
and UO_113 (O_113,N_2900,N_2761);
xnor UO_114 (O_114,N_2975,N_2979);
or UO_115 (O_115,N_2581,N_2682);
nand UO_116 (O_116,N_2696,N_2669);
and UO_117 (O_117,N_2725,N_2539);
or UO_118 (O_118,N_2917,N_2544);
xnor UO_119 (O_119,N_2710,N_2906);
or UO_120 (O_120,N_2853,N_2650);
or UO_121 (O_121,N_2850,N_2512);
nor UO_122 (O_122,N_2586,N_2508);
nor UO_123 (O_123,N_2744,N_2704);
or UO_124 (O_124,N_2655,N_2800);
and UO_125 (O_125,N_2997,N_2626);
or UO_126 (O_126,N_2998,N_2956);
nor UO_127 (O_127,N_2585,N_2769);
or UO_128 (O_128,N_2709,N_2559);
nand UO_129 (O_129,N_2993,N_2754);
and UO_130 (O_130,N_2686,N_2830);
nor UO_131 (O_131,N_2878,N_2921);
nand UO_132 (O_132,N_2894,N_2760);
nor UO_133 (O_133,N_2729,N_2907);
nand UO_134 (O_134,N_2635,N_2803);
or UO_135 (O_135,N_2617,N_2608);
nand UO_136 (O_136,N_2549,N_2910);
or UO_137 (O_137,N_2885,N_2609);
nand UO_138 (O_138,N_2732,N_2651);
or UO_139 (O_139,N_2623,N_2611);
and UO_140 (O_140,N_2786,N_2631);
and UO_141 (O_141,N_2857,N_2530);
or UO_142 (O_142,N_2846,N_2935);
nand UO_143 (O_143,N_2673,N_2550);
or UO_144 (O_144,N_2903,N_2973);
and UO_145 (O_145,N_2911,N_2931);
and UO_146 (O_146,N_2596,N_2934);
or UO_147 (O_147,N_2722,N_2902);
and UO_148 (O_148,N_2701,N_2672);
and UO_149 (O_149,N_2645,N_2734);
nand UO_150 (O_150,N_2535,N_2811);
and UO_151 (O_151,N_2793,N_2660);
and UO_152 (O_152,N_2506,N_2922);
nor UO_153 (O_153,N_2537,N_2575);
and UO_154 (O_154,N_2994,N_2520);
or UO_155 (O_155,N_2534,N_2995);
nand UO_156 (O_156,N_2976,N_2542);
nand UO_157 (O_157,N_2893,N_2514);
nand UO_158 (O_158,N_2816,N_2866);
nor UO_159 (O_159,N_2652,N_2591);
or UO_160 (O_160,N_2616,N_2521);
nand UO_161 (O_161,N_2984,N_2983);
or UO_162 (O_162,N_2778,N_2500);
or UO_163 (O_163,N_2781,N_2955);
nor UO_164 (O_164,N_2714,N_2733);
nor UO_165 (O_165,N_2721,N_2524);
nand UO_166 (O_166,N_2693,N_2713);
nor UO_167 (O_167,N_2605,N_2868);
nand UO_168 (O_168,N_2941,N_2865);
or UO_169 (O_169,N_2871,N_2640);
nor UO_170 (O_170,N_2901,N_2987);
or UO_171 (O_171,N_2855,N_2659);
and UO_172 (O_172,N_2583,N_2891);
nor UO_173 (O_173,N_2819,N_2771);
or UO_174 (O_174,N_2785,N_2977);
or UO_175 (O_175,N_2889,N_2795);
xor UO_176 (O_176,N_2661,N_2780);
or UO_177 (O_177,N_2880,N_2864);
nand UO_178 (O_178,N_2588,N_2666);
or UO_179 (O_179,N_2519,N_2723);
and UO_180 (O_180,N_2920,N_2560);
and UO_181 (O_181,N_2684,N_2555);
or UO_182 (O_182,N_2978,N_2510);
nand UO_183 (O_183,N_2777,N_2668);
and UO_184 (O_184,N_2892,N_2992);
nor UO_185 (O_185,N_2529,N_2517);
and UO_186 (O_186,N_2874,N_2576);
and UO_187 (O_187,N_2678,N_2601);
nor UO_188 (O_188,N_2610,N_2848);
nand UO_189 (O_189,N_2788,N_2964);
nand UO_190 (O_190,N_2629,N_2613);
and UO_191 (O_191,N_2926,N_2861);
nand UO_192 (O_192,N_2989,N_2879);
nand UO_193 (O_193,N_2797,N_2584);
and UO_194 (O_194,N_2838,N_2536);
nand UO_195 (O_195,N_2863,N_2646);
or UO_196 (O_196,N_2817,N_2825);
or UO_197 (O_197,N_2628,N_2567);
nand UO_198 (O_198,N_2947,N_2598);
or UO_199 (O_199,N_2974,N_2821);
and UO_200 (O_200,N_2731,N_2925);
nand UO_201 (O_201,N_2547,N_2702);
and UO_202 (O_202,N_2844,N_2587);
and UO_203 (O_203,N_2832,N_2770);
or UO_204 (O_204,N_2509,N_2810);
xor UO_205 (O_205,N_2815,N_2728);
and UO_206 (O_206,N_2680,N_2755);
xnor UO_207 (O_207,N_2620,N_2504);
nand UO_208 (O_208,N_2916,N_2840);
nand UO_209 (O_209,N_2738,N_2940);
and UO_210 (O_210,N_2751,N_2927);
or UO_211 (O_211,N_2818,N_2730);
nor UO_212 (O_212,N_2502,N_2630);
or UO_213 (O_213,N_2647,N_2747);
nand UO_214 (O_214,N_2887,N_2656);
or UO_215 (O_215,N_2882,N_2618);
or UO_216 (O_216,N_2919,N_2614);
or UO_217 (O_217,N_2758,N_2597);
or UO_218 (O_218,N_2968,N_2820);
nand UO_219 (O_219,N_2849,N_2943);
nand UO_220 (O_220,N_2774,N_2503);
nor UO_221 (O_221,N_2899,N_2619);
or UO_222 (O_222,N_2897,N_2958);
or UO_223 (O_223,N_2681,N_2945);
and UO_224 (O_224,N_2634,N_2638);
nand UO_225 (O_225,N_2595,N_2949);
nor UO_226 (O_226,N_2564,N_2642);
and UO_227 (O_227,N_2836,N_2930);
nand UO_228 (O_228,N_2507,N_2881);
nand UO_229 (O_229,N_2814,N_2579);
nor UO_230 (O_230,N_2606,N_2697);
or UO_231 (O_231,N_2981,N_2515);
and UO_232 (O_232,N_2773,N_2790);
nor UO_233 (O_233,N_2845,N_2540);
nor UO_234 (O_234,N_2752,N_2982);
or UO_235 (O_235,N_2957,N_2691);
and UO_236 (O_236,N_2523,N_2562);
nand UO_237 (O_237,N_2578,N_2699);
nor UO_238 (O_238,N_2625,N_2632);
or UO_239 (O_239,N_2707,N_2643);
xnor UO_240 (O_240,N_2522,N_2590);
nor UO_241 (O_241,N_2665,N_2716);
and UO_242 (O_242,N_2859,N_2852);
nand UO_243 (O_243,N_2962,N_2748);
nand UO_244 (O_244,N_2662,N_2644);
nand UO_245 (O_245,N_2648,N_2952);
nand UO_246 (O_246,N_2565,N_2768);
and UO_247 (O_247,N_2954,N_2890);
nand UO_248 (O_248,N_2552,N_2798);
or UO_249 (O_249,N_2545,N_2525);
or UO_250 (O_250,N_2981,N_2713);
and UO_251 (O_251,N_2725,N_2736);
and UO_252 (O_252,N_2613,N_2835);
or UO_253 (O_253,N_2601,N_2745);
and UO_254 (O_254,N_2533,N_2644);
nand UO_255 (O_255,N_2780,N_2935);
and UO_256 (O_256,N_2736,N_2836);
or UO_257 (O_257,N_2811,N_2699);
nor UO_258 (O_258,N_2953,N_2792);
and UO_259 (O_259,N_2630,N_2548);
or UO_260 (O_260,N_2948,N_2860);
nand UO_261 (O_261,N_2822,N_2980);
or UO_262 (O_262,N_2731,N_2795);
and UO_263 (O_263,N_2790,N_2936);
nand UO_264 (O_264,N_2567,N_2622);
nor UO_265 (O_265,N_2654,N_2600);
nand UO_266 (O_266,N_2523,N_2752);
and UO_267 (O_267,N_2602,N_2582);
or UO_268 (O_268,N_2682,N_2780);
and UO_269 (O_269,N_2736,N_2992);
and UO_270 (O_270,N_2814,N_2803);
or UO_271 (O_271,N_2912,N_2551);
nand UO_272 (O_272,N_2693,N_2659);
nor UO_273 (O_273,N_2960,N_2517);
or UO_274 (O_274,N_2534,N_2910);
or UO_275 (O_275,N_2982,N_2706);
or UO_276 (O_276,N_2560,N_2677);
nand UO_277 (O_277,N_2987,N_2968);
nor UO_278 (O_278,N_2802,N_2762);
or UO_279 (O_279,N_2856,N_2697);
nand UO_280 (O_280,N_2566,N_2665);
and UO_281 (O_281,N_2686,N_2615);
or UO_282 (O_282,N_2654,N_2863);
xor UO_283 (O_283,N_2560,N_2791);
nand UO_284 (O_284,N_2933,N_2581);
nor UO_285 (O_285,N_2877,N_2608);
and UO_286 (O_286,N_2720,N_2941);
nand UO_287 (O_287,N_2876,N_2723);
nand UO_288 (O_288,N_2712,N_2591);
or UO_289 (O_289,N_2609,N_2593);
and UO_290 (O_290,N_2984,N_2752);
or UO_291 (O_291,N_2710,N_2525);
and UO_292 (O_292,N_2655,N_2650);
nor UO_293 (O_293,N_2960,N_2522);
nor UO_294 (O_294,N_2677,N_2731);
nand UO_295 (O_295,N_2969,N_2506);
nor UO_296 (O_296,N_2778,N_2848);
or UO_297 (O_297,N_2531,N_2749);
and UO_298 (O_298,N_2871,N_2683);
nand UO_299 (O_299,N_2500,N_2596);
or UO_300 (O_300,N_2712,N_2845);
or UO_301 (O_301,N_2802,N_2501);
nor UO_302 (O_302,N_2583,N_2952);
and UO_303 (O_303,N_2691,N_2715);
nand UO_304 (O_304,N_2902,N_2814);
and UO_305 (O_305,N_2933,N_2705);
and UO_306 (O_306,N_2574,N_2883);
nand UO_307 (O_307,N_2918,N_2739);
and UO_308 (O_308,N_2523,N_2820);
or UO_309 (O_309,N_2694,N_2566);
xor UO_310 (O_310,N_2645,N_2911);
and UO_311 (O_311,N_2691,N_2656);
and UO_312 (O_312,N_2781,N_2867);
or UO_313 (O_313,N_2686,N_2559);
and UO_314 (O_314,N_2530,N_2988);
nand UO_315 (O_315,N_2990,N_2984);
nand UO_316 (O_316,N_2707,N_2571);
nor UO_317 (O_317,N_2630,N_2692);
or UO_318 (O_318,N_2571,N_2726);
nor UO_319 (O_319,N_2889,N_2988);
or UO_320 (O_320,N_2747,N_2559);
and UO_321 (O_321,N_2787,N_2629);
nand UO_322 (O_322,N_2645,N_2905);
nand UO_323 (O_323,N_2816,N_2502);
nor UO_324 (O_324,N_2978,N_2635);
nand UO_325 (O_325,N_2930,N_2824);
and UO_326 (O_326,N_2748,N_2752);
nand UO_327 (O_327,N_2592,N_2781);
nand UO_328 (O_328,N_2899,N_2913);
nor UO_329 (O_329,N_2932,N_2568);
and UO_330 (O_330,N_2803,N_2780);
and UO_331 (O_331,N_2548,N_2735);
nand UO_332 (O_332,N_2571,N_2752);
and UO_333 (O_333,N_2859,N_2888);
or UO_334 (O_334,N_2756,N_2936);
nor UO_335 (O_335,N_2632,N_2510);
or UO_336 (O_336,N_2518,N_2711);
or UO_337 (O_337,N_2807,N_2980);
nand UO_338 (O_338,N_2755,N_2959);
nand UO_339 (O_339,N_2638,N_2566);
or UO_340 (O_340,N_2953,N_2814);
nor UO_341 (O_341,N_2977,N_2913);
and UO_342 (O_342,N_2739,N_2976);
or UO_343 (O_343,N_2912,N_2678);
nor UO_344 (O_344,N_2565,N_2719);
or UO_345 (O_345,N_2569,N_2615);
nand UO_346 (O_346,N_2886,N_2905);
and UO_347 (O_347,N_2976,N_2970);
nor UO_348 (O_348,N_2691,N_2778);
and UO_349 (O_349,N_2546,N_2600);
and UO_350 (O_350,N_2956,N_2841);
or UO_351 (O_351,N_2827,N_2823);
nand UO_352 (O_352,N_2986,N_2634);
and UO_353 (O_353,N_2994,N_2929);
and UO_354 (O_354,N_2552,N_2867);
nor UO_355 (O_355,N_2587,N_2566);
and UO_356 (O_356,N_2691,N_2566);
nor UO_357 (O_357,N_2802,N_2821);
nor UO_358 (O_358,N_2887,N_2969);
and UO_359 (O_359,N_2916,N_2556);
and UO_360 (O_360,N_2732,N_2594);
or UO_361 (O_361,N_2678,N_2719);
or UO_362 (O_362,N_2862,N_2889);
nand UO_363 (O_363,N_2589,N_2853);
or UO_364 (O_364,N_2737,N_2519);
nand UO_365 (O_365,N_2677,N_2898);
and UO_366 (O_366,N_2653,N_2695);
or UO_367 (O_367,N_2785,N_2850);
nor UO_368 (O_368,N_2603,N_2646);
nand UO_369 (O_369,N_2662,N_2546);
nand UO_370 (O_370,N_2708,N_2674);
or UO_371 (O_371,N_2882,N_2974);
nand UO_372 (O_372,N_2867,N_2715);
nand UO_373 (O_373,N_2525,N_2696);
nand UO_374 (O_374,N_2705,N_2641);
and UO_375 (O_375,N_2808,N_2506);
nor UO_376 (O_376,N_2861,N_2785);
nor UO_377 (O_377,N_2661,N_2774);
nand UO_378 (O_378,N_2770,N_2737);
nand UO_379 (O_379,N_2576,N_2554);
nor UO_380 (O_380,N_2724,N_2674);
and UO_381 (O_381,N_2711,N_2736);
or UO_382 (O_382,N_2864,N_2582);
and UO_383 (O_383,N_2606,N_2525);
or UO_384 (O_384,N_2785,N_2818);
or UO_385 (O_385,N_2856,N_2539);
and UO_386 (O_386,N_2732,N_2949);
nor UO_387 (O_387,N_2771,N_2518);
and UO_388 (O_388,N_2814,N_2504);
and UO_389 (O_389,N_2579,N_2699);
nor UO_390 (O_390,N_2875,N_2892);
and UO_391 (O_391,N_2744,N_2660);
nand UO_392 (O_392,N_2840,N_2773);
and UO_393 (O_393,N_2927,N_2737);
nand UO_394 (O_394,N_2799,N_2784);
or UO_395 (O_395,N_2781,N_2549);
and UO_396 (O_396,N_2567,N_2917);
nand UO_397 (O_397,N_2978,N_2566);
and UO_398 (O_398,N_2947,N_2656);
nand UO_399 (O_399,N_2599,N_2753);
or UO_400 (O_400,N_2907,N_2657);
nor UO_401 (O_401,N_2884,N_2820);
nor UO_402 (O_402,N_2897,N_2885);
nand UO_403 (O_403,N_2983,N_2864);
or UO_404 (O_404,N_2716,N_2805);
or UO_405 (O_405,N_2751,N_2951);
nor UO_406 (O_406,N_2822,N_2876);
nor UO_407 (O_407,N_2897,N_2506);
nor UO_408 (O_408,N_2851,N_2970);
nand UO_409 (O_409,N_2711,N_2919);
or UO_410 (O_410,N_2613,N_2900);
or UO_411 (O_411,N_2546,N_2850);
or UO_412 (O_412,N_2566,N_2922);
nand UO_413 (O_413,N_2910,N_2665);
nor UO_414 (O_414,N_2616,N_2592);
nor UO_415 (O_415,N_2657,N_2597);
nor UO_416 (O_416,N_2709,N_2676);
nand UO_417 (O_417,N_2966,N_2659);
nor UO_418 (O_418,N_2983,N_2508);
and UO_419 (O_419,N_2809,N_2580);
nand UO_420 (O_420,N_2947,N_2772);
and UO_421 (O_421,N_2582,N_2919);
nand UO_422 (O_422,N_2899,N_2788);
nor UO_423 (O_423,N_2787,N_2724);
or UO_424 (O_424,N_2869,N_2992);
nand UO_425 (O_425,N_2734,N_2552);
or UO_426 (O_426,N_2867,N_2669);
or UO_427 (O_427,N_2657,N_2826);
nand UO_428 (O_428,N_2798,N_2638);
and UO_429 (O_429,N_2513,N_2823);
and UO_430 (O_430,N_2959,N_2896);
or UO_431 (O_431,N_2530,N_2931);
nand UO_432 (O_432,N_2526,N_2874);
nand UO_433 (O_433,N_2911,N_2890);
or UO_434 (O_434,N_2712,N_2568);
nand UO_435 (O_435,N_2590,N_2573);
and UO_436 (O_436,N_2983,N_2854);
nor UO_437 (O_437,N_2700,N_2995);
and UO_438 (O_438,N_2568,N_2999);
or UO_439 (O_439,N_2547,N_2899);
nor UO_440 (O_440,N_2674,N_2968);
or UO_441 (O_441,N_2555,N_2656);
nor UO_442 (O_442,N_2937,N_2516);
or UO_443 (O_443,N_2875,N_2982);
nand UO_444 (O_444,N_2882,N_2866);
nor UO_445 (O_445,N_2784,N_2972);
nand UO_446 (O_446,N_2743,N_2791);
nand UO_447 (O_447,N_2932,N_2787);
or UO_448 (O_448,N_2936,N_2892);
nor UO_449 (O_449,N_2537,N_2740);
and UO_450 (O_450,N_2932,N_2559);
nor UO_451 (O_451,N_2972,N_2857);
or UO_452 (O_452,N_2530,N_2697);
nor UO_453 (O_453,N_2528,N_2777);
and UO_454 (O_454,N_2888,N_2913);
nor UO_455 (O_455,N_2589,N_2968);
and UO_456 (O_456,N_2938,N_2740);
and UO_457 (O_457,N_2614,N_2664);
and UO_458 (O_458,N_2858,N_2738);
and UO_459 (O_459,N_2810,N_2618);
nand UO_460 (O_460,N_2555,N_2594);
nand UO_461 (O_461,N_2689,N_2968);
or UO_462 (O_462,N_2540,N_2850);
or UO_463 (O_463,N_2923,N_2728);
nor UO_464 (O_464,N_2945,N_2791);
nand UO_465 (O_465,N_2754,N_2768);
nand UO_466 (O_466,N_2806,N_2817);
or UO_467 (O_467,N_2725,N_2938);
nor UO_468 (O_468,N_2793,N_2887);
and UO_469 (O_469,N_2536,N_2907);
or UO_470 (O_470,N_2991,N_2844);
nand UO_471 (O_471,N_2737,N_2500);
nor UO_472 (O_472,N_2793,N_2923);
or UO_473 (O_473,N_2713,N_2880);
nand UO_474 (O_474,N_2701,N_2584);
or UO_475 (O_475,N_2571,N_2731);
and UO_476 (O_476,N_2691,N_2744);
or UO_477 (O_477,N_2818,N_2857);
or UO_478 (O_478,N_2751,N_2921);
or UO_479 (O_479,N_2774,N_2626);
and UO_480 (O_480,N_2938,N_2966);
or UO_481 (O_481,N_2746,N_2990);
or UO_482 (O_482,N_2815,N_2777);
or UO_483 (O_483,N_2706,N_2883);
and UO_484 (O_484,N_2799,N_2546);
nor UO_485 (O_485,N_2692,N_2696);
nand UO_486 (O_486,N_2644,N_2864);
or UO_487 (O_487,N_2644,N_2873);
or UO_488 (O_488,N_2826,N_2957);
nor UO_489 (O_489,N_2601,N_2519);
nor UO_490 (O_490,N_2877,N_2879);
or UO_491 (O_491,N_2542,N_2731);
nand UO_492 (O_492,N_2912,N_2723);
nand UO_493 (O_493,N_2763,N_2715);
nor UO_494 (O_494,N_2986,N_2564);
and UO_495 (O_495,N_2701,N_2694);
or UO_496 (O_496,N_2811,N_2683);
and UO_497 (O_497,N_2653,N_2528);
nor UO_498 (O_498,N_2645,N_2828);
nor UO_499 (O_499,N_2931,N_2635);
endmodule