module basic_1000_10000_1500_4_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_834,In_860);
xnor U1 (N_1,In_399,In_342);
nor U2 (N_2,In_246,In_906);
or U3 (N_3,In_242,In_603);
and U4 (N_4,In_710,In_71);
and U5 (N_5,In_219,In_248);
and U6 (N_6,In_544,In_194);
xor U7 (N_7,In_718,In_138);
and U8 (N_8,In_769,In_363);
nand U9 (N_9,In_359,In_182);
nand U10 (N_10,In_193,In_371);
and U11 (N_11,In_421,In_628);
or U12 (N_12,In_930,In_383);
nand U13 (N_13,In_841,In_514);
xnor U14 (N_14,In_118,In_878);
and U15 (N_15,In_882,In_444);
and U16 (N_16,In_588,In_65);
nor U17 (N_17,In_941,In_216);
nor U18 (N_18,In_899,In_497);
nand U19 (N_19,In_129,In_637);
or U20 (N_20,In_554,In_477);
nand U21 (N_21,In_354,In_794);
nand U22 (N_22,In_706,In_20);
and U23 (N_23,In_453,In_745);
nor U24 (N_24,In_967,In_229);
nor U25 (N_25,In_534,In_387);
or U26 (N_26,In_867,In_367);
or U27 (N_27,In_462,In_110);
or U28 (N_28,In_600,In_936);
or U29 (N_29,In_950,In_673);
nand U30 (N_30,In_679,In_349);
nand U31 (N_31,In_379,In_774);
nand U32 (N_32,In_664,In_251);
xor U33 (N_33,In_776,In_59);
and U34 (N_34,In_144,In_921);
nor U35 (N_35,In_966,In_148);
nor U36 (N_36,In_202,In_322);
nand U37 (N_37,In_463,In_592);
and U38 (N_38,In_807,In_250);
and U39 (N_39,In_33,In_333);
nand U40 (N_40,In_137,In_700);
and U41 (N_41,In_605,In_760);
xor U42 (N_42,In_509,In_294);
xnor U43 (N_43,In_960,In_73);
nor U44 (N_44,In_908,In_666);
nor U45 (N_45,In_988,In_5);
xor U46 (N_46,In_397,In_441);
or U47 (N_47,In_757,In_39);
and U48 (N_48,In_364,In_729);
xnor U49 (N_49,In_844,In_842);
and U50 (N_50,In_264,In_321);
xor U51 (N_51,In_398,In_344);
and U52 (N_52,In_702,In_355);
nand U53 (N_53,In_647,In_295);
xnor U54 (N_54,In_775,In_366);
nand U55 (N_55,In_997,In_581);
xnor U56 (N_56,In_817,In_318);
nand U57 (N_57,In_106,In_580);
and U58 (N_58,In_429,In_991);
nand U59 (N_59,In_262,In_939);
nor U60 (N_60,In_88,In_586);
nand U61 (N_61,In_224,In_912);
nor U62 (N_62,In_886,In_206);
nor U63 (N_63,In_112,In_909);
and U64 (N_64,In_46,In_782);
xnor U65 (N_65,In_515,In_986);
nand U66 (N_66,In_963,In_542);
or U67 (N_67,In_707,In_495);
xnor U68 (N_68,In_676,In_286);
or U69 (N_69,In_197,In_597);
or U70 (N_70,In_492,In_215);
xor U71 (N_71,In_61,In_887);
or U72 (N_72,In_334,In_984);
nor U73 (N_73,In_907,In_640);
or U74 (N_74,In_473,In_155);
nor U75 (N_75,In_633,In_320);
or U76 (N_76,In_890,In_271);
and U77 (N_77,In_725,In_313);
and U78 (N_78,In_783,In_470);
and U79 (N_79,In_560,In_977);
and U80 (N_80,In_884,In_837);
xor U81 (N_81,In_516,In_96);
nand U82 (N_82,In_213,In_501);
xnor U83 (N_83,In_356,In_770);
and U84 (N_84,In_653,In_937);
nor U85 (N_85,In_563,In_763);
nand U86 (N_86,In_846,In_613);
nor U87 (N_87,In_170,In_734);
nor U88 (N_88,In_927,In_49);
nand U89 (N_89,In_51,In_21);
and U90 (N_90,In_704,In_975);
and U91 (N_91,In_851,In_690);
and U92 (N_92,In_722,In_925);
and U93 (N_93,In_768,In_481);
nor U94 (N_94,In_522,In_451);
nand U95 (N_95,In_715,In_735);
nor U96 (N_96,In_802,In_86);
and U97 (N_97,In_133,In_317);
nor U98 (N_98,In_864,In_716);
and U99 (N_99,In_773,In_787);
nor U100 (N_100,In_616,In_232);
nand U101 (N_101,In_839,In_486);
or U102 (N_102,In_430,In_684);
or U103 (N_103,In_460,In_401);
nor U104 (N_104,In_200,In_798);
or U105 (N_105,In_184,In_27);
or U106 (N_106,In_162,In_352);
nand U107 (N_107,In_693,In_845);
and U108 (N_108,In_237,In_924);
nand U109 (N_109,In_645,In_132);
and U110 (N_110,In_268,In_56);
or U111 (N_111,In_620,In_981);
and U112 (N_112,In_69,In_928);
or U113 (N_113,In_272,In_404);
nor U114 (N_114,In_256,In_524);
nand U115 (N_115,In_150,In_705);
and U116 (N_116,In_15,In_553);
xnor U117 (N_117,In_743,In_391);
or U118 (N_118,In_119,In_999);
or U119 (N_119,In_468,In_736);
nand U120 (N_120,In_141,In_573);
nor U121 (N_121,In_151,In_233);
nor U122 (N_122,In_708,In_897);
or U123 (N_123,In_260,In_900);
nor U124 (N_124,In_149,In_120);
nand U125 (N_125,In_183,In_953);
nand U126 (N_126,In_862,In_425);
nor U127 (N_127,In_888,In_538);
nor U128 (N_128,In_815,In_266);
xor U129 (N_129,In_961,In_191);
nor U130 (N_130,In_18,In_228);
or U131 (N_131,In_612,In_362);
nand U132 (N_132,In_423,In_916);
or U133 (N_133,In_668,In_669);
nand U134 (N_134,In_723,In_587);
and U135 (N_135,In_885,In_324);
nor U136 (N_136,In_315,In_856);
nor U137 (N_137,In_656,In_830);
or U138 (N_138,In_348,In_225);
nand U139 (N_139,In_488,In_91);
or U140 (N_140,In_732,In_582);
and U141 (N_141,In_572,In_389);
nor U142 (N_142,In_220,In_730);
nand U143 (N_143,In_208,In_617);
nor U144 (N_144,In_503,In_944);
xnor U145 (N_145,In_316,In_214);
and U146 (N_146,In_595,In_848);
nor U147 (N_147,In_697,In_124);
xor U148 (N_148,In_40,In_337);
nand U149 (N_149,In_667,In_147);
and U150 (N_150,In_373,In_518);
nor U151 (N_151,In_11,In_414);
or U152 (N_152,In_555,In_788);
and U153 (N_153,In_771,In_350);
or U154 (N_154,In_341,In_83);
and U155 (N_155,In_520,In_703);
and U156 (N_156,In_559,In_254);
nand U157 (N_157,In_499,In_335);
and U158 (N_158,In_995,In_166);
nor U159 (N_159,In_614,In_978);
or U160 (N_160,In_591,In_942);
nand U161 (N_161,In_824,In_467);
or U162 (N_162,In_100,In_458);
and U163 (N_163,In_820,In_370);
xor U164 (N_164,In_738,In_546);
and U165 (N_165,In_75,In_750);
or U166 (N_166,In_808,In_236);
nand U167 (N_167,In_935,In_479);
and U168 (N_168,In_828,In_279);
nand U169 (N_169,In_245,In_827);
or U170 (N_170,In_3,In_529);
and U171 (N_171,In_455,In_759);
xor U172 (N_172,In_934,In_374);
nor U173 (N_173,In_556,In_993);
or U174 (N_174,In_408,In_28);
nor U175 (N_175,In_861,In_478);
nor U176 (N_176,In_606,In_660);
or U177 (N_177,In_426,In_831);
nand U178 (N_178,In_583,In_390);
and U179 (N_179,In_179,In_611);
or U180 (N_180,In_417,In_375);
nor U181 (N_181,In_810,In_577);
xnor U182 (N_182,In_416,In_41);
and U183 (N_183,In_386,In_525);
and U184 (N_184,In_513,In_159);
nor U185 (N_185,In_276,In_169);
xnor U186 (N_186,In_24,In_466);
and U187 (N_187,In_552,In_594);
and U188 (N_188,In_376,In_168);
or U189 (N_189,In_8,In_319);
nand U190 (N_190,In_93,In_484);
and U191 (N_191,In_517,In_154);
nand U192 (N_192,In_331,In_1);
and U193 (N_193,In_671,In_608);
xnor U194 (N_194,In_982,In_528);
or U195 (N_195,In_532,In_480);
and U196 (N_196,In_267,In_34);
and U197 (N_197,In_461,In_662);
and U198 (N_198,In_285,In_923);
nor U199 (N_199,In_139,In_626);
nor U200 (N_200,In_502,In_911);
xor U201 (N_201,In_762,In_474);
nand U202 (N_202,In_792,In_761);
or U203 (N_203,In_403,In_955);
nand U204 (N_204,In_485,In_439);
nor U205 (N_205,In_167,In_510);
xor U206 (N_206,In_687,In_454);
and U207 (N_207,In_918,In_629);
or U208 (N_208,In_283,In_678);
nor U209 (N_209,In_415,In_48);
or U210 (N_210,In_239,In_959);
xor U211 (N_211,In_622,In_130);
nand U212 (N_212,In_692,In_646);
and U213 (N_213,In_186,In_914);
nor U214 (N_214,In_14,In_744);
xor U215 (N_215,In_63,In_109);
nor U216 (N_216,In_803,In_160);
and U217 (N_217,In_464,In_602);
nor U218 (N_218,In_411,In_819);
or U219 (N_219,In_128,In_537);
nor U220 (N_220,In_895,In_306);
and U221 (N_221,In_437,In_420);
and U222 (N_222,In_876,In_883);
nor U223 (N_223,In_192,In_288);
and U224 (N_224,In_952,In_541);
nor U225 (N_225,In_311,In_372);
nand U226 (N_226,In_994,In_593);
xnor U227 (N_227,In_325,In_70);
or U228 (N_228,In_104,In_619);
or U229 (N_229,In_789,In_241);
and U230 (N_230,In_983,In_257);
and U231 (N_231,In_47,In_507);
nand U232 (N_232,In_418,In_790);
nand U233 (N_233,In_6,In_125);
nor U234 (N_234,In_670,In_171);
nor U235 (N_235,In_134,In_742);
and U236 (N_236,In_490,In_599);
nand U237 (N_237,In_938,In_832);
and U238 (N_238,In_747,In_596);
nor U239 (N_239,In_658,In_701);
and U240 (N_240,In_623,In_469);
nor U241 (N_241,In_946,In_579);
nor U242 (N_242,In_339,In_615);
nor U243 (N_243,In_252,In_30);
and U244 (N_244,In_407,In_32);
nor U245 (N_245,In_235,In_330);
or U246 (N_246,In_209,In_145);
nor U247 (N_247,In_574,In_521);
nor U248 (N_248,In_287,In_400);
or U249 (N_249,In_432,In_643);
nor U250 (N_250,In_314,In_569);
nor U251 (N_251,In_299,In_44);
or U252 (N_252,In_627,In_199);
and U253 (N_253,In_865,In_858);
and U254 (N_254,In_135,In_530);
or U255 (N_255,In_326,In_227);
xor U256 (N_256,In_230,In_970);
nor U257 (N_257,In_452,In_487);
nor U258 (N_258,In_631,In_724);
nor U259 (N_259,In_836,In_175);
and U260 (N_260,In_31,In_739);
nand U261 (N_261,In_717,In_855);
nor U262 (N_262,In_238,In_728);
nor U263 (N_263,In_207,In_465);
nor U264 (N_264,In_825,In_859);
nand U265 (N_265,In_576,In_434);
and U266 (N_266,In_847,In_726);
or U267 (N_267,In_632,In_709);
or U268 (N_268,In_508,In_903);
nor U269 (N_269,In_327,In_741);
nand U270 (N_270,In_79,In_217);
nand U271 (N_271,In_796,In_877);
or U272 (N_272,In_377,In_29);
or U273 (N_273,In_598,In_351);
nand U274 (N_274,In_338,In_113);
and U275 (N_275,In_805,In_277);
nand U276 (N_276,In_68,In_97);
and U277 (N_277,In_570,In_53);
or U278 (N_278,In_987,In_410);
or U279 (N_279,In_731,In_292);
nand U280 (N_280,In_0,In_625);
nor U281 (N_281,In_663,In_764);
and U282 (N_282,In_752,In_800);
xor U283 (N_283,In_748,In_558);
and U284 (N_284,In_694,In_2);
and U285 (N_285,In_117,In_565);
nor U286 (N_286,In_969,In_38);
and U287 (N_287,In_797,In_644);
and U288 (N_288,In_826,In_945);
or U289 (N_289,In_940,In_161);
nor U290 (N_290,In_265,In_714);
nor U291 (N_291,In_852,In_17);
and U292 (N_292,In_7,In_875);
nand U293 (N_293,In_66,In_650);
xor U294 (N_294,In_164,In_240);
or U295 (N_295,In_234,In_504);
nor U296 (N_296,In_298,In_177);
and U297 (N_297,In_523,In_749);
or U298 (N_298,In_290,In_419);
xnor U299 (N_299,In_691,In_55);
or U300 (N_300,In_695,In_578);
xnor U301 (N_301,In_243,In_590);
and U302 (N_302,In_816,In_733);
or U303 (N_303,In_84,In_123);
nand U304 (N_304,In_158,In_87);
nor U305 (N_305,In_893,In_607);
nor U306 (N_306,In_998,In_740);
nand U307 (N_307,In_780,In_482);
or U308 (N_308,In_801,In_98);
nand U309 (N_309,In_822,In_108);
nor U310 (N_310,In_428,In_649);
nand U311 (N_311,In_360,In_833);
or U312 (N_312,In_77,In_853);
and U313 (N_313,In_89,In_345);
nor U314 (N_314,In_122,In_424);
xor U315 (N_315,In_665,In_329);
nand U316 (N_316,In_926,In_871);
nand U317 (N_317,In_943,In_821);
nand U318 (N_318,In_526,In_686);
nand U319 (N_319,In_835,In_874);
and U320 (N_320,In_94,In_57);
and U321 (N_321,In_101,In_621);
nor U322 (N_322,In_720,In_567);
and U323 (N_323,In_917,In_795);
and U324 (N_324,In_196,In_436);
nor U325 (N_325,In_639,In_571);
nor U326 (N_326,In_549,In_378);
or U327 (N_327,In_811,In_527);
or U328 (N_328,In_312,In_618);
nand U329 (N_329,In_442,In_261);
and U330 (N_330,In_712,In_231);
nand U331 (N_331,In_711,In_74);
xnor U332 (N_332,In_919,In_672);
nand U333 (N_333,In_965,In_449);
nor U334 (N_334,In_755,In_476);
and U335 (N_335,In_624,In_512);
or U336 (N_336,In_548,In_247);
and U337 (N_337,In_394,In_178);
nor U338 (N_338,In_443,In_433);
xor U339 (N_339,In_396,In_758);
nand U340 (N_340,In_221,In_323);
and U341 (N_341,In_369,In_872);
nand U342 (N_342,In_804,In_146);
nor U343 (N_343,In_547,In_651);
nand U344 (N_344,In_153,In_103);
or U345 (N_345,In_980,In_683);
or U346 (N_346,In_636,In_920);
nand U347 (N_347,In_869,In_222);
or U348 (N_348,In_968,In_358);
nor U349 (N_349,In_902,In_840);
and U350 (N_350,In_721,In_962);
nor U351 (N_351,In_772,In_385);
or U352 (N_352,In_630,In_737);
nor U353 (N_353,In_519,In_682);
nor U354 (N_354,In_812,In_450);
nand U355 (N_355,In_568,In_45);
nand U356 (N_356,In_881,In_187);
and U357 (N_357,In_12,In_785);
or U358 (N_358,In_402,In_849);
nor U359 (N_359,In_990,In_289);
and U360 (N_360,In_427,In_185);
or U361 (N_361,In_80,In_974);
or U362 (N_362,In_244,In_95);
nand U363 (N_363,In_301,In_648);
and U364 (N_364,In_483,In_889);
and U365 (N_365,In_674,In_566);
nand U366 (N_366,In_136,In_879);
nand U367 (N_367,In_72,In_604);
nor U368 (N_368,In_43,In_67);
nor U369 (N_369,In_652,In_438);
or U370 (N_370,In_395,In_412);
xnor U371 (N_371,In_309,In_85);
nor U372 (N_372,In_806,In_380);
nor U373 (N_373,In_947,In_10);
xor U374 (N_374,In_910,In_964);
nor U375 (N_375,In_357,In_23);
nand U376 (N_376,In_562,In_756);
nand U377 (N_377,In_866,In_156);
or U378 (N_378,In_76,In_259);
nor U379 (N_379,In_751,In_62);
nand U380 (N_380,In_300,In_188);
and U381 (N_381,In_440,In_829);
or U382 (N_382,In_37,In_972);
nand U383 (N_383,In_857,In_791);
nor U384 (N_384,In_445,In_223);
and U385 (N_385,In_269,In_302);
nand U386 (N_386,In_82,In_505);
or U387 (N_387,In_195,In_713);
or U388 (N_388,In_680,In_753);
or U389 (N_389,In_675,In_173);
and U390 (N_390,In_561,In_564);
nand U391 (N_391,In_343,In_746);
nand U392 (N_392,In_281,In_174);
and U393 (N_393,In_280,In_901);
and U394 (N_394,In_814,In_661);
nand U395 (N_395,In_448,In_635);
or U396 (N_396,In_19,In_340);
nand U397 (N_397,In_610,In_543);
nor U398 (N_398,In_754,In_533);
and U399 (N_399,In_152,In_36);
xnor U400 (N_400,In_293,In_111);
and U401 (N_401,In_446,In_413);
xor U402 (N_402,In_255,In_346);
or U403 (N_403,In_699,In_305);
or U404 (N_404,In_212,In_551);
nand U405 (N_405,In_843,In_368);
nand U406 (N_406,In_489,In_64);
nand U407 (N_407,In_81,In_353);
nand U408 (N_408,In_22,In_498);
nor U409 (N_409,In_540,In_54);
and U410 (N_410,In_838,In_303);
nor U411 (N_411,In_898,In_655);
and U412 (N_412,In_308,In_949);
nor U413 (N_413,In_634,In_52);
nand U414 (N_414,In_304,In_275);
nor U415 (N_415,In_765,In_896);
and U416 (N_416,In_818,In_107);
or U417 (N_417,In_201,In_979);
nor U418 (N_418,In_258,In_913);
nor U419 (N_419,In_105,In_190);
or U420 (N_420,In_163,In_584);
and U421 (N_421,In_471,In_870);
nor U422 (N_422,In_456,In_511);
nand U423 (N_423,In_689,In_850);
xor U424 (N_424,In_60,In_659);
and U425 (N_425,In_929,In_557);
and U426 (N_426,In_274,In_210);
or U427 (N_427,In_78,In_270);
and U428 (N_428,In_328,In_9);
and U429 (N_429,In_809,In_863);
or U430 (N_430,In_115,In_905);
nand U431 (N_431,In_172,In_472);
xnor U432 (N_432,In_971,In_204);
xnor U433 (N_433,In_140,In_50);
nand U434 (N_434,In_892,In_99);
nor U435 (N_435,In_297,In_102);
or U436 (N_436,In_786,In_126);
xnor U437 (N_437,In_696,In_127);
and U438 (N_438,In_585,In_657);
nand U439 (N_439,In_435,In_958);
nor U440 (N_440,In_915,In_575);
or U441 (N_441,In_58,In_422);
nand U442 (N_442,In_951,In_799);
nor U443 (N_443,In_431,In_116);
nand U444 (N_444,In_347,In_891);
nand U445 (N_445,In_406,In_957);
nand U446 (N_446,In_218,In_121);
nand U447 (N_447,In_550,In_189);
nand U448 (N_448,In_13,In_642);
xnor U449 (N_449,In_609,In_641);
nor U450 (N_450,In_654,In_205);
xor U451 (N_451,In_16,In_589);
nor U452 (N_452,In_545,In_296);
xor U453 (N_453,In_813,In_500);
nor U454 (N_454,In_181,In_948);
or U455 (N_455,In_365,In_392);
nor U456 (N_456,In_361,In_447);
nand U457 (N_457,In_211,In_601);
nor U458 (N_458,In_868,In_779);
or U459 (N_459,In_932,In_35);
nand U460 (N_460,In_719,In_698);
and U461 (N_461,In_685,In_535);
nand U462 (N_462,In_727,In_336);
and U463 (N_463,In_131,In_793);
nor U464 (N_464,In_291,In_203);
and U465 (N_465,In_781,In_976);
nand U466 (N_466,In_382,In_996);
nand U467 (N_467,In_491,In_496);
xor U468 (N_468,In_989,In_4);
nand U469 (N_469,In_854,In_494);
and U470 (N_470,In_677,In_198);
nor U471 (N_471,In_278,In_475);
nor U472 (N_472,In_273,In_284);
or U473 (N_473,In_310,In_536);
or U474 (N_474,In_142,In_457);
nand U475 (N_475,In_638,In_681);
nor U476 (N_476,In_539,In_384);
nor U477 (N_477,In_933,In_493);
nand U478 (N_478,In_506,In_531);
nor U479 (N_479,In_992,In_332);
and U480 (N_480,In_157,In_114);
nor U481 (N_481,In_25,In_778);
xnor U482 (N_482,In_409,In_904);
and U483 (N_483,In_226,In_307);
nor U484 (N_484,In_688,In_823);
or U485 (N_485,In_954,In_42);
nor U486 (N_486,In_931,In_894);
or U487 (N_487,In_176,In_393);
nor U488 (N_488,In_973,In_766);
nand U489 (N_489,In_767,In_459);
nand U490 (N_490,In_26,In_405);
and U491 (N_491,In_282,In_784);
and U492 (N_492,In_180,In_249);
and U493 (N_493,In_956,In_253);
or U494 (N_494,In_388,In_777);
xor U495 (N_495,In_165,In_263);
or U496 (N_496,In_143,In_873);
or U497 (N_497,In_880,In_985);
nor U498 (N_498,In_381,In_92);
and U499 (N_499,In_90,In_922);
nand U500 (N_500,In_958,In_887);
xnor U501 (N_501,In_138,In_36);
nor U502 (N_502,In_247,In_561);
nand U503 (N_503,In_703,In_707);
and U504 (N_504,In_891,In_838);
or U505 (N_505,In_249,In_692);
or U506 (N_506,In_718,In_311);
and U507 (N_507,In_163,In_280);
or U508 (N_508,In_743,In_666);
or U509 (N_509,In_19,In_590);
and U510 (N_510,In_381,In_637);
and U511 (N_511,In_794,In_357);
nand U512 (N_512,In_64,In_544);
nand U513 (N_513,In_516,In_859);
nand U514 (N_514,In_427,In_142);
and U515 (N_515,In_77,In_786);
or U516 (N_516,In_267,In_166);
and U517 (N_517,In_693,In_309);
nor U518 (N_518,In_150,In_408);
xnor U519 (N_519,In_586,In_9);
nand U520 (N_520,In_361,In_980);
nand U521 (N_521,In_297,In_415);
and U522 (N_522,In_44,In_422);
nor U523 (N_523,In_452,In_559);
xor U524 (N_524,In_877,In_405);
nand U525 (N_525,In_159,In_789);
nor U526 (N_526,In_74,In_750);
nand U527 (N_527,In_882,In_725);
xor U528 (N_528,In_918,In_756);
or U529 (N_529,In_880,In_657);
nor U530 (N_530,In_815,In_143);
and U531 (N_531,In_521,In_492);
nand U532 (N_532,In_869,In_311);
and U533 (N_533,In_580,In_504);
nand U534 (N_534,In_985,In_192);
and U535 (N_535,In_521,In_712);
nand U536 (N_536,In_743,In_815);
nor U537 (N_537,In_52,In_611);
nand U538 (N_538,In_923,In_762);
nand U539 (N_539,In_661,In_874);
and U540 (N_540,In_938,In_873);
nand U541 (N_541,In_823,In_242);
or U542 (N_542,In_128,In_323);
nand U543 (N_543,In_457,In_535);
or U544 (N_544,In_359,In_266);
and U545 (N_545,In_894,In_304);
and U546 (N_546,In_367,In_731);
nand U547 (N_547,In_424,In_912);
nand U548 (N_548,In_330,In_717);
nand U549 (N_549,In_332,In_741);
and U550 (N_550,In_154,In_729);
nor U551 (N_551,In_723,In_532);
and U552 (N_552,In_492,In_120);
or U553 (N_553,In_790,In_678);
nand U554 (N_554,In_221,In_977);
or U555 (N_555,In_274,In_183);
nand U556 (N_556,In_371,In_14);
and U557 (N_557,In_698,In_716);
nand U558 (N_558,In_468,In_134);
nor U559 (N_559,In_832,In_661);
nand U560 (N_560,In_169,In_983);
and U561 (N_561,In_930,In_921);
and U562 (N_562,In_704,In_147);
nand U563 (N_563,In_396,In_470);
xor U564 (N_564,In_713,In_841);
nor U565 (N_565,In_848,In_956);
nand U566 (N_566,In_364,In_498);
nand U567 (N_567,In_197,In_146);
or U568 (N_568,In_991,In_459);
xor U569 (N_569,In_626,In_890);
or U570 (N_570,In_80,In_411);
and U571 (N_571,In_319,In_393);
nand U572 (N_572,In_869,In_211);
and U573 (N_573,In_69,In_423);
nand U574 (N_574,In_451,In_906);
and U575 (N_575,In_655,In_912);
xnor U576 (N_576,In_547,In_754);
or U577 (N_577,In_981,In_899);
nor U578 (N_578,In_567,In_810);
xor U579 (N_579,In_549,In_713);
nor U580 (N_580,In_460,In_59);
or U581 (N_581,In_923,In_722);
xnor U582 (N_582,In_635,In_869);
nor U583 (N_583,In_809,In_739);
or U584 (N_584,In_567,In_504);
xnor U585 (N_585,In_124,In_805);
nor U586 (N_586,In_171,In_243);
and U587 (N_587,In_318,In_422);
or U588 (N_588,In_868,In_973);
nand U589 (N_589,In_660,In_205);
or U590 (N_590,In_623,In_446);
and U591 (N_591,In_615,In_996);
and U592 (N_592,In_816,In_585);
nor U593 (N_593,In_508,In_484);
and U594 (N_594,In_573,In_233);
nand U595 (N_595,In_627,In_808);
xor U596 (N_596,In_502,In_425);
nand U597 (N_597,In_550,In_865);
xor U598 (N_598,In_486,In_217);
and U599 (N_599,In_527,In_682);
or U600 (N_600,In_587,In_140);
and U601 (N_601,In_881,In_738);
nand U602 (N_602,In_371,In_703);
xor U603 (N_603,In_575,In_567);
and U604 (N_604,In_728,In_996);
and U605 (N_605,In_930,In_860);
and U606 (N_606,In_283,In_302);
or U607 (N_607,In_56,In_608);
nor U608 (N_608,In_124,In_666);
and U609 (N_609,In_374,In_186);
or U610 (N_610,In_295,In_472);
or U611 (N_611,In_240,In_942);
and U612 (N_612,In_382,In_230);
and U613 (N_613,In_545,In_647);
nor U614 (N_614,In_295,In_883);
or U615 (N_615,In_865,In_753);
or U616 (N_616,In_877,In_999);
nand U617 (N_617,In_849,In_1);
xor U618 (N_618,In_612,In_797);
nor U619 (N_619,In_429,In_809);
or U620 (N_620,In_559,In_632);
nand U621 (N_621,In_330,In_770);
xnor U622 (N_622,In_679,In_240);
or U623 (N_623,In_247,In_272);
nand U624 (N_624,In_24,In_768);
nor U625 (N_625,In_712,In_32);
or U626 (N_626,In_95,In_28);
nor U627 (N_627,In_369,In_435);
nor U628 (N_628,In_220,In_528);
nor U629 (N_629,In_482,In_976);
and U630 (N_630,In_794,In_403);
xor U631 (N_631,In_569,In_211);
and U632 (N_632,In_602,In_329);
or U633 (N_633,In_986,In_575);
xnor U634 (N_634,In_575,In_917);
nor U635 (N_635,In_578,In_783);
nand U636 (N_636,In_515,In_718);
or U637 (N_637,In_817,In_493);
nor U638 (N_638,In_823,In_789);
nor U639 (N_639,In_840,In_240);
nand U640 (N_640,In_967,In_594);
or U641 (N_641,In_591,In_151);
nand U642 (N_642,In_672,In_199);
xnor U643 (N_643,In_578,In_808);
nor U644 (N_644,In_810,In_963);
nor U645 (N_645,In_23,In_480);
or U646 (N_646,In_179,In_484);
and U647 (N_647,In_888,In_399);
or U648 (N_648,In_495,In_475);
nor U649 (N_649,In_141,In_560);
nand U650 (N_650,In_352,In_191);
nor U651 (N_651,In_42,In_875);
and U652 (N_652,In_481,In_763);
xnor U653 (N_653,In_866,In_21);
nand U654 (N_654,In_177,In_503);
and U655 (N_655,In_748,In_487);
nor U656 (N_656,In_571,In_332);
or U657 (N_657,In_482,In_270);
and U658 (N_658,In_690,In_127);
nand U659 (N_659,In_314,In_46);
and U660 (N_660,In_635,In_390);
nand U661 (N_661,In_289,In_399);
and U662 (N_662,In_831,In_32);
nor U663 (N_663,In_95,In_978);
nand U664 (N_664,In_591,In_165);
or U665 (N_665,In_132,In_379);
or U666 (N_666,In_210,In_614);
or U667 (N_667,In_27,In_639);
or U668 (N_668,In_9,In_677);
nor U669 (N_669,In_467,In_823);
and U670 (N_670,In_129,In_425);
xnor U671 (N_671,In_80,In_472);
nand U672 (N_672,In_830,In_944);
xnor U673 (N_673,In_752,In_256);
or U674 (N_674,In_218,In_232);
nor U675 (N_675,In_121,In_497);
xor U676 (N_676,In_884,In_559);
nor U677 (N_677,In_373,In_497);
nor U678 (N_678,In_58,In_168);
or U679 (N_679,In_949,In_863);
xnor U680 (N_680,In_501,In_592);
or U681 (N_681,In_829,In_84);
nand U682 (N_682,In_5,In_548);
nor U683 (N_683,In_719,In_187);
nor U684 (N_684,In_173,In_151);
nor U685 (N_685,In_195,In_785);
or U686 (N_686,In_536,In_499);
nand U687 (N_687,In_45,In_705);
nand U688 (N_688,In_928,In_472);
or U689 (N_689,In_257,In_818);
or U690 (N_690,In_60,In_389);
nand U691 (N_691,In_750,In_971);
nand U692 (N_692,In_978,In_32);
and U693 (N_693,In_315,In_951);
xor U694 (N_694,In_294,In_11);
nand U695 (N_695,In_348,In_360);
nand U696 (N_696,In_448,In_918);
nand U697 (N_697,In_335,In_966);
and U698 (N_698,In_236,In_712);
xnor U699 (N_699,In_327,In_313);
and U700 (N_700,In_127,In_314);
nor U701 (N_701,In_982,In_593);
nor U702 (N_702,In_17,In_726);
nand U703 (N_703,In_639,In_292);
nor U704 (N_704,In_528,In_859);
nand U705 (N_705,In_382,In_525);
and U706 (N_706,In_32,In_390);
nand U707 (N_707,In_785,In_521);
or U708 (N_708,In_270,In_234);
nand U709 (N_709,In_857,In_420);
xor U710 (N_710,In_304,In_303);
and U711 (N_711,In_236,In_958);
nand U712 (N_712,In_701,In_115);
nor U713 (N_713,In_282,In_956);
nand U714 (N_714,In_563,In_270);
nand U715 (N_715,In_92,In_703);
and U716 (N_716,In_542,In_329);
nand U717 (N_717,In_970,In_538);
and U718 (N_718,In_272,In_788);
and U719 (N_719,In_784,In_968);
nor U720 (N_720,In_266,In_551);
nor U721 (N_721,In_277,In_700);
nor U722 (N_722,In_120,In_678);
and U723 (N_723,In_246,In_439);
nor U724 (N_724,In_252,In_983);
and U725 (N_725,In_409,In_829);
nand U726 (N_726,In_941,In_652);
nor U727 (N_727,In_351,In_165);
nand U728 (N_728,In_581,In_944);
and U729 (N_729,In_409,In_28);
and U730 (N_730,In_866,In_638);
or U731 (N_731,In_522,In_911);
nand U732 (N_732,In_441,In_573);
nor U733 (N_733,In_393,In_375);
and U734 (N_734,In_290,In_930);
and U735 (N_735,In_581,In_964);
nand U736 (N_736,In_910,In_715);
nor U737 (N_737,In_655,In_608);
nor U738 (N_738,In_793,In_820);
xor U739 (N_739,In_18,In_247);
nor U740 (N_740,In_635,In_107);
nand U741 (N_741,In_883,In_917);
nand U742 (N_742,In_513,In_184);
and U743 (N_743,In_642,In_819);
and U744 (N_744,In_991,In_648);
nand U745 (N_745,In_303,In_724);
nand U746 (N_746,In_324,In_987);
and U747 (N_747,In_635,In_35);
xor U748 (N_748,In_60,In_692);
or U749 (N_749,In_595,In_169);
or U750 (N_750,In_177,In_5);
and U751 (N_751,In_522,In_17);
nand U752 (N_752,In_7,In_282);
or U753 (N_753,In_720,In_255);
xor U754 (N_754,In_352,In_354);
and U755 (N_755,In_133,In_515);
nand U756 (N_756,In_601,In_250);
and U757 (N_757,In_441,In_898);
nor U758 (N_758,In_860,In_656);
and U759 (N_759,In_405,In_346);
nand U760 (N_760,In_529,In_279);
or U761 (N_761,In_343,In_332);
and U762 (N_762,In_798,In_677);
nand U763 (N_763,In_997,In_513);
nand U764 (N_764,In_77,In_427);
and U765 (N_765,In_151,In_562);
nor U766 (N_766,In_809,In_205);
nand U767 (N_767,In_69,In_575);
nor U768 (N_768,In_897,In_416);
and U769 (N_769,In_163,In_348);
or U770 (N_770,In_975,In_677);
xor U771 (N_771,In_258,In_717);
xor U772 (N_772,In_878,In_180);
or U773 (N_773,In_277,In_701);
nor U774 (N_774,In_82,In_117);
xnor U775 (N_775,In_568,In_242);
nor U776 (N_776,In_702,In_585);
nand U777 (N_777,In_101,In_313);
xnor U778 (N_778,In_966,In_884);
nor U779 (N_779,In_86,In_245);
or U780 (N_780,In_336,In_212);
nand U781 (N_781,In_760,In_443);
nand U782 (N_782,In_512,In_684);
nor U783 (N_783,In_721,In_53);
or U784 (N_784,In_444,In_238);
nor U785 (N_785,In_741,In_165);
nor U786 (N_786,In_991,In_59);
or U787 (N_787,In_658,In_747);
and U788 (N_788,In_18,In_9);
xnor U789 (N_789,In_659,In_632);
or U790 (N_790,In_972,In_904);
nand U791 (N_791,In_755,In_575);
nor U792 (N_792,In_953,In_447);
or U793 (N_793,In_244,In_242);
nand U794 (N_794,In_306,In_618);
and U795 (N_795,In_271,In_460);
and U796 (N_796,In_430,In_402);
nand U797 (N_797,In_614,In_64);
and U798 (N_798,In_716,In_930);
xnor U799 (N_799,In_585,In_669);
nand U800 (N_800,In_665,In_78);
nand U801 (N_801,In_443,In_176);
xor U802 (N_802,In_718,In_637);
or U803 (N_803,In_536,In_503);
or U804 (N_804,In_159,In_793);
or U805 (N_805,In_664,In_556);
nor U806 (N_806,In_961,In_286);
nor U807 (N_807,In_399,In_531);
xor U808 (N_808,In_464,In_776);
nand U809 (N_809,In_14,In_399);
or U810 (N_810,In_914,In_588);
and U811 (N_811,In_661,In_666);
nand U812 (N_812,In_981,In_807);
nand U813 (N_813,In_581,In_857);
xor U814 (N_814,In_159,In_799);
nand U815 (N_815,In_903,In_826);
nor U816 (N_816,In_75,In_793);
nand U817 (N_817,In_814,In_63);
xnor U818 (N_818,In_782,In_602);
nand U819 (N_819,In_529,In_956);
nor U820 (N_820,In_678,In_785);
nor U821 (N_821,In_83,In_54);
and U822 (N_822,In_666,In_516);
xnor U823 (N_823,In_911,In_295);
or U824 (N_824,In_716,In_603);
or U825 (N_825,In_72,In_135);
nor U826 (N_826,In_117,In_956);
or U827 (N_827,In_234,In_505);
or U828 (N_828,In_57,In_672);
xor U829 (N_829,In_551,In_599);
and U830 (N_830,In_302,In_393);
and U831 (N_831,In_865,In_879);
nor U832 (N_832,In_151,In_763);
or U833 (N_833,In_653,In_230);
and U834 (N_834,In_993,In_278);
or U835 (N_835,In_638,In_806);
nor U836 (N_836,In_655,In_250);
or U837 (N_837,In_30,In_907);
xor U838 (N_838,In_376,In_324);
and U839 (N_839,In_140,In_502);
nor U840 (N_840,In_726,In_197);
xor U841 (N_841,In_631,In_93);
nor U842 (N_842,In_144,In_709);
xnor U843 (N_843,In_643,In_80);
nand U844 (N_844,In_904,In_393);
and U845 (N_845,In_669,In_655);
or U846 (N_846,In_203,In_637);
or U847 (N_847,In_170,In_252);
xnor U848 (N_848,In_825,In_670);
and U849 (N_849,In_51,In_574);
nand U850 (N_850,In_605,In_738);
or U851 (N_851,In_314,In_503);
nand U852 (N_852,In_135,In_295);
nand U853 (N_853,In_304,In_379);
nor U854 (N_854,In_120,In_327);
nor U855 (N_855,In_770,In_736);
or U856 (N_856,In_64,In_126);
and U857 (N_857,In_486,In_658);
nor U858 (N_858,In_842,In_687);
and U859 (N_859,In_678,In_532);
xnor U860 (N_860,In_23,In_364);
xnor U861 (N_861,In_575,In_568);
nor U862 (N_862,In_786,In_961);
or U863 (N_863,In_851,In_176);
xnor U864 (N_864,In_929,In_131);
and U865 (N_865,In_747,In_278);
or U866 (N_866,In_471,In_425);
and U867 (N_867,In_518,In_974);
nor U868 (N_868,In_630,In_147);
nor U869 (N_869,In_128,In_114);
or U870 (N_870,In_130,In_613);
nand U871 (N_871,In_619,In_78);
or U872 (N_872,In_58,In_51);
or U873 (N_873,In_995,In_745);
nand U874 (N_874,In_127,In_753);
nor U875 (N_875,In_451,In_329);
nor U876 (N_876,In_155,In_906);
or U877 (N_877,In_90,In_564);
and U878 (N_878,In_2,In_592);
or U879 (N_879,In_211,In_218);
nor U880 (N_880,In_118,In_670);
and U881 (N_881,In_880,In_285);
nor U882 (N_882,In_796,In_221);
nand U883 (N_883,In_229,In_89);
or U884 (N_884,In_255,In_966);
and U885 (N_885,In_776,In_524);
nand U886 (N_886,In_599,In_60);
nor U887 (N_887,In_823,In_552);
nand U888 (N_888,In_515,In_374);
and U889 (N_889,In_252,In_245);
nand U890 (N_890,In_741,In_385);
or U891 (N_891,In_943,In_49);
nor U892 (N_892,In_255,In_881);
xor U893 (N_893,In_836,In_797);
and U894 (N_894,In_89,In_594);
nand U895 (N_895,In_230,In_322);
or U896 (N_896,In_596,In_227);
nor U897 (N_897,In_749,In_516);
and U898 (N_898,In_238,In_824);
nand U899 (N_899,In_873,In_803);
nand U900 (N_900,In_998,In_235);
or U901 (N_901,In_137,In_490);
nor U902 (N_902,In_51,In_255);
or U903 (N_903,In_198,In_89);
nor U904 (N_904,In_122,In_607);
nor U905 (N_905,In_561,In_497);
or U906 (N_906,In_762,In_200);
or U907 (N_907,In_354,In_439);
nand U908 (N_908,In_823,In_8);
nor U909 (N_909,In_739,In_840);
xor U910 (N_910,In_703,In_713);
or U911 (N_911,In_463,In_583);
and U912 (N_912,In_167,In_927);
nor U913 (N_913,In_338,In_516);
nand U914 (N_914,In_922,In_277);
nor U915 (N_915,In_242,In_38);
and U916 (N_916,In_302,In_175);
and U917 (N_917,In_56,In_919);
nor U918 (N_918,In_454,In_406);
nand U919 (N_919,In_620,In_264);
and U920 (N_920,In_952,In_852);
nor U921 (N_921,In_449,In_82);
nor U922 (N_922,In_427,In_557);
or U923 (N_923,In_107,In_648);
and U924 (N_924,In_296,In_876);
nand U925 (N_925,In_929,In_518);
nor U926 (N_926,In_605,In_828);
or U927 (N_927,In_605,In_781);
nand U928 (N_928,In_227,In_934);
xor U929 (N_929,In_691,In_638);
nand U930 (N_930,In_857,In_865);
or U931 (N_931,In_301,In_12);
xnor U932 (N_932,In_642,In_523);
or U933 (N_933,In_742,In_704);
and U934 (N_934,In_714,In_334);
and U935 (N_935,In_301,In_320);
or U936 (N_936,In_740,In_86);
and U937 (N_937,In_873,In_729);
xor U938 (N_938,In_558,In_588);
and U939 (N_939,In_708,In_920);
xor U940 (N_940,In_29,In_512);
or U941 (N_941,In_240,In_235);
nor U942 (N_942,In_766,In_639);
or U943 (N_943,In_756,In_740);
nand U944 (N_944,In_22,In_358);
nand U945 (N_945,In_478,In_44);
xnor U946 (N_946,In_881,In_979);
nand U947 (N_947,In_623,In_953);
nand U948 (N_948,In_727,In_749);
nor U949 (N_949,In_222,In_702);
nor U950 (N_950,In_330,In_91);
nand U951 (N_951,In_374,In_200);
nor U952 (N_952,In_260,In_465);
or U953 (N_953,In_212,In_206);
xor U954 (N_954,In_981,In_340);
or U955 (N_955,In_162,In_78);
nor U956 (N_956,In_111,In_701);
or U957 (N_957,In_886,In_76);
nand U958 (N_958,In_953,In_717);
nor U959 (N_959,In_198,In_904);
or U960 (N_960,In_881,In_468);
or U961 (N_961,In_224,In_595);
nand U962 (N_962,In_378,In_474);
nor U963 (N_963,In_788,In_108);
or U964 (N_964,In_915,In_344);
and U965 (N_965,In_27,In_362);
or U966 (N_966,In_391,In_787);
or U967 (N_967,In_128,In_125);
nor U968 (N_968,In_941,In_2);
and U969 (N_969,In_57,In_444);
and U970 (N_970,In_442,In_180);
nor U971 (N_971,In_209,In_621);
or U972 (N_972,In_703,In_618);
and U973 (N_973,In_373,In_219);
xnor U974 (N_974,In_102,In_917);
and U975 (N_975,In_766,In_160);
and U976 (N_976,In_512,In_907);
nand U977 (N_977,In_806,In_373);
nand U978 (N_978,In_384,In_612);
nand U979 (N_979,In_57,In_914);
nand U980 (N_980,In_565,In_480);
nand U981 (N_981,In_440,In_408);
nor U982 (N_982,In_251,In_473);
nor U983 (N_983,In_29,In_233);
or U984 (N_984,In_110,In_475);
nor U985 (N_985,In_438,In_632);
xor U986 (N_986,In_877,In_946);
nor U987 (N_987,In_819,In_105);
nand U988 (N_988,In_953,In_227);
nand U989 (N_989,In_867,In_148);
or U990 (N_990,In_14,In_476);
xor U991 (N_991,In_224,In_126);
nor U992 (N_992,In_132,In_782);
nand U993 (N_993,In_972,In_65);
or U994 (N_994,In_833,In_692);
nor U995 (N_995,In_727,In_298);
nor U996 (N_996,In_484,In_344);
or U997 (N_997,In_538,In_855);
and U998 (N_998,In_486,In_470);
nand U999 (N_999,In_583,In_103);
nand U1000 (N_1000,In_174,In_237);
or U1001 (N_1001,In_675,In_727);
nand U1002 (N_1002,In_699,In_20);
or U1003 (N_1003,In_46,In_980);
xnor U1004 (N_1004,In_859,In_791);
nor U1005 (N_1005,In_57,In_88);
nand U1006 (N_1006,In_967,In_503);
nor U1007 (N_1007,In_473,In_758);
xor U1008 (N_1008,In_439,In_600);
and U1009 (N_1009,In_220,In_294);
or U1010 (N_1010,In_938,In_939);
nand U1011 (N_1011,In_498,In_289);
nor U1012 (N_1012,In_123,In_249);
nor U1013 (N_1013,In_651,In_808);
or U1014 (N_1014,In_805,In_920);
nor U1015 (N_1015,In_437,In_181);
and U1016 (N_1016,In_292,In_299);
and U1017 (N_1017,In_365,In_340);
or U1018 (N_1018,In_9,In_584);
xnor U1019 (N_1019,In_9,In_353);
nor U1020 (N_1020,In_682,In_214);
nor U1021 (N_1021,In_809,In_7);
nand U1022 (N_1022,In_637,In_989);
nor U1023 (N_1023,In_646,In_761);
nand U1024 (N_1024,In_131,In_685);
nand U1025 (N_1025,In_127,In_790);
and U1026 (N_1026,In_270,In_703);
or U1027 (N_1027,In_911,In_499);
nor U1028 (N_1028,In_708,In_894);
and U1029 (N_1029,In_458,In_188);
and U1030 (N_1030,In_308,In_120);
xor U1031 (N_1031,In_776,In_291);
nor U1032 (N_1032,In_2,In_83);
and U1033 (N_1033,In_142,In_570);
and U1034 (N_1034,In_18,In_988);
or U1035 (N_1035,In_331,In_828);
nand U1036 (N_1036,In_348,In_245);
nor U1037 (N_1037,In_803,In_127);
nand U1038 (N_1038,In_569,In_578);
nor U1039 (N_1039,In_997,In_989);
or U1040 (N_1040,In_196,In_334);
or U1041 (N_1041,In_692,In_445);
or U1042 (N_1042,In_327,In_475);
or U1043 (N_1043,In_563,In_692);
nor U1044 (N_1044,In_176,In_286);
nor U1045 (N_1045,In_5,In_211);
and U1046 (N_1046,In_823,In_423);
or U1047 (N_1047,In_463,In_225);
nand U1048 (N_1048,In_143,In_90);
and U1049 (N_1049,In_196,In_292);
nand U1050 (N_1050,In_151,In_493);
or U1051 (N_1051,In_217,In_480);
nand U1052 (N_1052,In_461,In_454);
or U1053 (N_1053,In_938,In_160);
and U1054 (N_1054,In_785,In_72);
or U1055 (N_1055,In_123,In_214);
and U1056 (N_1056,In_771,In_67);
nand U1057 (N_1057,In_418,In_947);
nand U1058 (N_1058,In_203,In_196);
xnor U1059 (N_1059,In_440,In_173);
or U1060 (N_1060,In_711,In_343);
nor U1061 (N_1061,In_532,In_7);
and U1062 (N_1062,In_709,In_614);
nor U1063 (N_1063,In_657,In_621);
or U1064 (N_1064,In_550,In_551);
nand U1065 (N_1065,In_286,In_338);
nand U1066 (N_1066,In_611,In_623);
nand U1067 (N_1067,In_685,In_671);
nand U1068 (N_1068,In_835,In_395);
and U1069 (N_1069,In_252,In_798);
and U1070 (N_1070,In_675,In_853);
or U1071 (N_1071,In_939,In_720);
or U1072 (N_1072,In_723,In_466);
and U1073 (N_1073,In_251,In_286);
nor U1074 (N_1074,In_252,In_744);
or U1075 (N_1075,In_865,In_228);
and U1076 (N_1076,In_31,In_573);
nand U1077 (N_1077,In_290,In_734);
and U1078 (N_1078,In_400,In_958);
nor U1079 (N_1079,In_37,In_29);
nor U1080 (N_1080,In_793,In_409);
nor U1081 (N_1081,In_558,In_183);
nand U1082 (N_1082,In_829,In_518);
nand U1083 (N_1083,In_408,In_612);
or U1084 (N_1084,In_783,In_45);
nand U1085 (N_1085,In_893,In_154);
nor U1086 (N_1086,In_116,In_492);
and U1087 (N_1087,In_845,In_210);
or U1088 (N_1088,In_684,In_774);
nor U1089 (N_1089,In_609,In_389);
and U1090 (N_1090,In_957,In_750);
or U1091 (N_1091,In_314,In_5);
xnor U1092 (N_1092,In_122,In_728);
nor U1093 (N_1093,In_454,In_495);
or U1094 (N_1094,In_862,In_379);
nand U1095 (N_1095,In_972,In_768);
or U1096 (N_1096,In_114,In_901);
and U1097 (N_1097,In_428,In_749);
or U1098 (N_1098,In_260,In_764);
nand U1099 (N_1099,In_862,In_78);
nor U1100 (N_1100,In_687,In_200);
or U1101 (N_1101,In_838,In_646);
nor U1102 (N_1102,In_260,In_191);
and U1103 (N_1103,In_647,In_513);
nand U1104 (N_1104,In_667,In_363);
nand U1105 (N_1105,In_504,In_403);
or U1106 (N_1106,In_495,In_862);
or U1107 (N_1107,In_395,In_791);
nand U1108 (N_1108,In_768,In_608);
or U1109 (N_1109,In_532,In_837);
and U1110 (N_1110,In_374,In_698);
nor U1111 (N_1111,In_394,In_816);
or U1112 (N_1112,In_455,In_101);
or U1113 (N_1113,In_948,In_406);
and U1114 (N_1114,In_351,In_462);
nor U1115 (N_1115,In_408,In_496);
nand U1116 (N_1116,In_99,In_436);
and U1117 (N_1117,In_42,In_68);
or U1118 (N_1118,In_347,In_47);
xnor U1119 (N_1119,In_891,In_251);
and U1120 (N_1120,In_38,In_144);
or U1121 (N_1121,In_794,In_460);
or U1122 (N_1122,In_101,In_156);
nand U1123 (N_1123,In_314,In_142);
or U1124 (N_1124,In_725,In_304);
nand U1125 (N_1125,In_407,In_199);
nor U1126 (N_1126,In_351,In_72);
or U1127 (N_1127,In_843,In_599);
nand U1128 (N_1128,In_841,In_244);
nand U1129 (N_1129,In_795,In_834);
nand U1130 (N_1130,In_213,In_198);
and U1131 (N_1131,In_62,In_604);
and U1132 (N_1132,In_325,In_781);
nand U1133 (N_1133,In_868,In_156);
and U1134 (N_1134,In_475,In_795);
or U1135 (N_1135,In_733,In_449);
nand U1136 (N_1136,In_690,In_509);
nand U1137 (N_1137,In_21,In_629);
nand U1138 (N_1138,In_18,In_421);
nor U1139 (N_1139,In_635,In_91);
and U1140 (N_1140,In_456,In_720);
xnor U1141 (N_1141,In_132,In_216);
or U1142 (N_1142,In_432,In_266);
nand U1143 (N_1143,In_734,In_8);
and U1144 (N_1144,In_140,In_476);
nand U1145 (N_1145,In_676,In_342);
nor U1146 (N_1146,In_864,In_800);
or U1147 (N_1147,In_465,In_992);
nor U1148 (N_1148,In_676,In_240);
or U1149 (N_1149,In_926,In_378);
or U1150 (N_1150,In_835,In_211);
nor U1151 (N_1151,In_488,In_462);
and U1152 (N_1152,In_206,In_889);
or U1153 (N_1153,In_159,In_945);
and U1154 (N_1154,In_828,In_656);
nor U1155 (N_1155,In_458,In_996);
nand U1156 (N_1156,In_197,In_683);
or U1157 (N_1157,In_632,In_992);
xor U1158 (N_1158,In_787,In_418);
and U1159 (N_1159,In_921,In_599);
nand U1160 (N_1160,In_315,In_86);
nand U1161 (N_1161,In_972,In_292);
nand U1162 (N_1162,In_745,In_736);
nand U1163 (N_1163,In_889,In_524);
xor U1164 (N_1164,In_630,In_120);
nand U1165 (N_1165,In_865,In_332);
xor U1166 (N_1166,In_310,In_532);
or U1167 (N_1167,In_124,In_82);
or U1168 (N_1168,In_66,In_495);
nand U1169 (N_1169,In_42,In_557);
or U1170 (N_1170,In_991,In_344);
and U1171 (N_1171,In_399,In_230);
nand U1172 (N_1172,In_988,In_119);
or U1173 (N_1173,In_436,In_386);
nor U1174 (N_1174,In_1,In_902);
and U1175 (N_1175,In_434,In_570);
nand U1176 (N_1176,In_840,In_632);
nor U1177 (N_1177,In_121,In_313);
and U1178 (N_1178,In_994,In_284);
nor U1179 (N_1179,In_586,In_977);
nor U1180 (N_1180,In_65,In_320);
xnor U1181 (N_1181,In_707,In_29);
xor U1182 (N_1182,In_106,In_915);
or U1183 (N_1183,In_830,In_553);
nand U1184 (N_1184,In_499,In_869);
nand U1185 (N_1185,In_122,In_444);
and U1186 (N_1186,In_31,In_527);
nor U1187 (N_1187,In_746,In_81);
nor U1188 (N_1188,In_691,In_545);
xnor U1189 (N_1189,In_955,In_81);
or U1190 (N_1190,In_270,In_460);
nor U1191 (N_1191,In_222,In_293);
xnor U1192 (N_1192,In_696,In_938);
and U1193 (N_1193,In_155,In_596);
and U1194 (N_1194,In_820,In_755);
nor U1195 (N_1195,In_909,In_996);
nand U1196 (N_1196,In_409,In_363);
xor U1197 (N_1197,In_20,In_364);
and U1198 (N_1198,In_245,In_94);
nand U1199 (N_1199,In_277,In_904);
nor U1200 (N_1200,In_101,In_957);
nor U1201 (N_1201,In_570,In_267);
or U1202 (N_1202,In_345,In_330);
and U1203 (N_1203,In_779,In_799);
xor U1204 (N_1204,In_507,In_951);
and U1205 (N_1205,In_495,In_698);
xnor U1206 (N_1206,In_823,In_953);
nand U1207 (N_1207,In_588,In_13);
xor U1208 (N_1208,In_703,In_310);
xnor U1209 (N_1209,In_549,In_511);
nor U1210 (N_1210,In_362,In_618);
nand U1211 (N_1211,In_348,In_878);
nor U1212 (N_1212,In_648,In_524);
or U1213 (N_1213,In_593,In_845);
or U1214 (N_1214,In_453,In_194);
xor U1215 (N_1215,In_129,In_303);
nor U1216 (N_1216,In_650,In_192);
or U1217 (N_1217,In_208,In_309);
xor U1218 (N_1218,In_105,In_767);
and U1219 (N_1219,In_179,In_631);
nand U1220 (N_1220,In_853,In_489);
and U1221 (N_1221,In_369,In_284);
nand U1222 (N_1222,In_406,In_692);
nor U1223 (N_1223,In_602,In_347);
or U1224 (N_1224,In_389,In_446);
nand U1225 (N_1225,In_290,In_440);
nor U1226 (N_1226,In_89,In_565);
nor U1227 (N_1227,In_456,In_230);
or U1228 (N_1228,In_574,In_142);
nand U1229 (N_1229,In_77,In_249);
and U1230 (N_1230,In_243,In_300);
or U1231 (N_1231,In_346,In_285);
nor U1232 (N_1232,In_199,In_593);
and U1233 (N_1233,In_950,In_228);
and U1234 (N_1234,In_520,In_13);
and U1235 (N_1235,In_598,In_67);
and U1236 (N_1236,In_256,In_699);
xor U1237 (N_1237,In_596,In_919);
nand U1238 (N_1238,In_206,In_26);
nand U1239 (N_1239,In_523,In_140);
nor U1240 (N_1240,In_850,In_861);
or U1241 (N_1241,In_328,In_176);
and U1242 (N_1242,In_367,In_548);
xnor U1243 (N_1243,In_558,In_957);
and U1244 (N_1244,In_61,In_14);
or U1245 (N_1245,In_778,In_308);
and U1246 (N_1246,In_123,In_791);
nand U1247 (N_1247,In_525,In_446);
and U1248 (N_1248,In_763,In_696);
and U1249 (N_1249,In_6,In_530);
and U1250 (N_1250,In_709,In_582);
and U1251 (N_1251,In_974,In_139);
or U1252 (N_1252,In_473,In_390);
nor U1253 (N_1253,In_655,In_59);
nor U1254 (N_1254,In_861,In_84);
nor U1255 (N_1255,In_548,In_973);
or U1256 (N_1256,In_246,In_543);
xnor U1257 (N_1257,In_994,In_177);
and U1258 (N_1258,In_844,In_160);
xnor U1259 (N_1259,In_934,In_461);
nor U1260 (N_1260,In_604,In_321);
and U1261 (N_1261,In_223,In_27);
nand U1262 (N_1262,In_269,In_760);
nand U1263 (N_1263,In_400,In_414);
or U1264 (N_1264,In_321,In_629);
nor U1265 (N_1265,In_124,In_671);
and U1266 (N_1266,In_292,In_861);
or U1267 (N_1267,In_586,In_773);
nand U1268 (N_1268,In_749,In_937);
and U1269 (N_1269,In_509,In_151);
and U1270 (N_1270,In_168,In_624);
nor U1271 (N_1271,In_973,In_845);
or U1272 (N_1272,In_953,In_773);
nor U1273 (N_1273,In_550,In_970);
nand U1274 (N_1274,In_685,In_234);
or U1275 (N_1275,In_66,In_287);
nand U1276 (N_1276,In_40,In_907);
nand U1277 (N_1277,In_730,In_934);
and U1278 (N_1278,In_189,In_853);
nor U1279 (N_1279,In_60,In_397);
nor U1280 (N_1280,In_550,In_355);
nor U1281 (N_1281,In_200,In_910);
or U1282 (N_1282,In_551,In_267);
or U1283 (N_1283,In_336,In_406);
or U1284 (N_1284,In_85,In_572);
nand U1285 (N_1285,In_690,In_541);
or U1286 (N_1286,In_503,In_411);
nand U1287 (N_1287,In_232,In_482);
or U1288 (N_1288,In_687,In_901);
and U1289 (N_1289,In_136,In_608);
and U1290 (N_1290,In_661,In_282);
nor U1291 (N_1291,In_541,In_561);
and U1292 (N_1292,In_944,In_100);
nor U1293 (N_1293,In_165,In_371);
or U1294 (N_1294,In_731,In_88);
and U1295 (N_1295,In_681,In_11);
or U1296 (N_1296,In_949,In_256);
and U1297 (N_1297,In_965,In_161);
xnor U1298 (N_1298,In_907,In_792);
nand U1299 (N_1299,In_799,In_53);
xor U1300 (N_1300,In_893,In_106);
or U1301 (N_1301,In_809,In_774);
and U1302 (N_1302,In_239,In_535);
and U1303 (N_1303,In_704,In_368);
or U1304 (N_1304,In_64,In_289);
and U1305 (N_1305,In_113,In_419);
and U1306 (N_1306,In_893,In_620);
nor U1307 (N_1307,In_901,In_427);
nand U1308 (N_1308,In_915,In_96);
and U1309 (N_1309,In_3,In_761);
and U1310 (N_1310,In_315,In_371);
and U1311 (N_1311,In_661,In_421);
or U1312 (N_1312,In_8,In_422);
nand U1313 (N_1313,In_2,In_119);
nand U1314 (N_1314,In_382,In_67);
nor U1315 (N_1315,In_815,In_731);
or U1316 (N_1316,In_796,In_677);
nand U1317 (N_1317,In_674,In_721);
nor U1318 (N_1318,In_310,In_368);
nor U1319 (N_1319,In_479,In_628);
nand U1320 (N_1320,In_170,In_319);
nand U1321 (N_1321,In_702,In_578);
nand U1322 (N_1322,In_235,In_145);
nand U1323 (N_1323,In_329,In_834);
or U1324 (N_1324,In_964,In_147);
or U1325 (N_1325,In_477,In_951);
xor U1326 (N_1326,In_994,In_64);
nand U1327 (N_1327,In_935,In_360);
nor U1328 (N_1328,In_485,In_16);
or U1329 (N_1329,In_945,In_740);
nor U1330 (N_1330,In_971,In_707);
nor U1331 (N_1331,In_536,In_875);
or U1332 (N_1332,In_396,In_168);
or U1333 (N_1333,In_84,In_663);
nor U1334 (N_1334,In_172,In_919);
nand U1335 (N_1335,In_724,In_873);
or U1336 (N_1336,In_868,In_365);
xnor U1337 (N_1337,In_817,In_335);
nor U1338 (N_1338,In_382,In_909);
or U1339 (N_1339,In_647,In_231);
and U1340 (N_1340,In_703,In_837);
nor U1341 (N_1341,In_828,In_483);
and U1342 (N_1342,In_607,In_428);
nor U1343 (N_1343,In_313,In_983);
nand U1344 (N_1344,In_575,In_566);
xnor U1345 (N_1345,In_787,In_387);
xnor U1346 (N_1346,In_972,In_656);
and U1347 (N_1347,In_650,In_707);
nor U1348 (N_1348,In_313,In_600);
and U1349 (N_1349,In_272,In_919);
and U1350 (N_1350,In_603,In_121);
or U1351 (N_1351,In_177,In_984);
and U1352 (N_1352,In_897,In_670);
nand U1353 (N_1353,In_282,In_524);
nor U1354 (N_1354,In_834,In_439);
and U1355 (N_1355,In_207,In_745);
nand U1356 (N_1356,In_543,In_3);
nor U1357 (N_1357,In_321,In_377);
nor U1358 (N_1358,In_429,In_459);
or U1359 (N_1359,In_684,In_188);
nand U1360 (N_1360,In_995,In_535);
and U1361 (N_1361,In_935,In_576);
and U1362 (N_1362,In_985,In_302);
nor U1363 (N_1363,In_163,In_421);
xnor U1364 (N_1364,In_689,In_382);
nand U1365 (N_1365,In_677,In_1);
nor U1366 (N_1366,In_147,In_478);
or U1367 (N_1367,In_386,In_927);
nor U1368 (N_1368,In_331,In_547);
and U1369 (N_1369,In_783,In_638);
and U1370 (N_1370,In_392,In_282);
and U1371 (N_1371,In_502,In_723);
or U1372 (N_1372,In_713,In_938);
xor U1373 (N_1373,In_426,In_477);
and U1374 (N_1374,In_362,In_868);
or U1375 (N_1375,In_819,In_634);
and U1376 (N_1376,In_61,In_647);
and U1377 (N_1377,In_441,In_702);
nor U1378 (N_1378,In_700,In_951);
and U1379 (N_1379,In_127,In_118);
or U1380 (N_1380,In_335,In_918);
nor U1381 (N_1381,In_254,In_239);
nand U1382 (N_1382,In_155,In_276);
nor U1383 (N_1383,In_386,In_268);
nor U1384 (N_1384,In_445,In_890);
or U1385 (N_1385,In_68,In_629);
and U1386 (N_1386,In_595,In_597);
or U1387 (N_1387,In_46,In_789);
nor U1388 (N_1388,In_851,In_707);
xor U1389 (N_1389,In_980,In_951);
or U1390 (N_1390,In_92,In_581);
xor U1391 (N_1391,In_242,In_496);
and U1392 (N_1392,In_342,In_10);
xnor U1393 (N_1393,In_299,In_93);
xnor U1394 (N_1394,In_707,In_214);
nor U1395 (N_1395,In_741,In_136);
or U1396 (N_1396,In_326,In_144);
nor U1397 (N_1397,In_528,In_892);
nand U1398 (N_1398,In_989,In_157);
nand U1399 (N_1399,In_172,In_710);
or U1400 (N_1400,In_181,In_8);
and U1401 (N_1401,In_853,In_880);
and U1402 (N_1402,In_170,In_946);
nand U1403 (N_1403,In_272,In_690);
or U1404 (N_1404,In_848,In_692);
nand U1405 (N_1405,In_555,In_541);
or U1406 (N_1406,In_638,In_775);
and U1407 (N_1407,In_300,In_556);
nor U1408 (N_1408,In_387,In_447);
nor U1409 (N_1409,In_946,In_542);
or U1410 (N_1410,In_462,In_702);
and U1411 (N_1411,In_280,In_711);
or U1412 (N_1412,In_405,In_157);
or U1413 (N_1413,In_846,In_509);
nor U1414 (N_1414,In_921,In_867);
xor U1415 (N_1415,In_863,In_261);
and U1416 (N_1416,In_967,In_552);
nor U1417 (N_1417,In_923,In_879);
nor U1418 (N_1418,In_375,In_272);
or U1419 (N_1419,In_785,In_824);
nand U1420 (N_1420,In_226,In_700);
and U1421 (N_1421,In_408,In_517);
or U1422 (N_1422,In_710,In_238);
or U1423 (N_1423,In_576,In_760);
nand U1424 (N_1424,In_881,In_546);
nand U1425 (N_1425,In_533,In_911);
and U1426 (N_1426,In_468,In_742);
or U1427 (N_1427,In_877,In_881);
nand U1428 (N_1428,In_971,In_96);
and U1429 (N_1429,In_643,In_622);
nor U1430 (N_1430,In_474,In_670);
and U1431 (N_1431,In_667,In_6);
nor U1432 (N_1432,In_90,In_659);
nor U1433 (N_1433,In_395,In_696);
and U1434 (N_1434,In_187,In_390);
or U1435 (N_1435,In_260,In_511);
xor U1436 (N_1436,In_153,In_228);
or U1437 (N_1437,In_783,In_262);
xor U1438 (N_1438,In_593,In_839);
and U1439 (N_1439,In_328,In_272);
nor U1440 (N_1440,In_66,In_490);
and U1441 (N_1441,In_242,In_494);
nor U1442 (N_1442,In_854,In_462);
nor U1443 (N_1443,In_405,In_309);
or U1444 (N_1444,In_739,In_250);
or U1445 (N_1445,In_46,In_503);
nand U1446 (N_1446,In_877,In_613);
or U1447 (N_1447,In_767,In_57);
and U1448 (N_1448,In_700,In_754);
nand U1449 (N_1449,In_569,In_555);
nand U1450 (N_1450,In_743,In_436);
and U1451 (N_1451,In_143,In_464);
nor U1452 (N_1452,In_823,In_938);
and U1453 (N_1453,In_963,In_231);
nor U1454 (N_1454,In_403,In_264);
nor U1455 (N_1455,In_789,In_849);
and U1456 (N_1456,In_248,In_591);
or U1457 (N_1457,In_27,In_35);
and U1458 (N_1458,In_313,In_738);
xor U1459 (N_1459,In_242,In_360);
or U1460 (N_1460,In_501,In_810);
or U1461 (N_1461,In_912,In_8);
and U1462 (N_1462,In_915,In_990);
nand U1463 (N_1463,In_653,In_717);
nand U1464 (N_1464,In_351,In_15);
nor U1465 (N_1465,In_746,In_929);
or U1466 (N_1466,In_839,In_936);
and U1467 (N_1467,In_259,In_667);
nand U1468 (N_1468,In_223,In_996);
and U1469 (N_1469,In_822,In_332);
nand U1470 (N_1470,In_725,In_59);
xnor U1471 (N_1471,In_343,In_544);
nor U1472 (N_1472,In_345,In_979);
nand U1473 (N_1473,In_615,In_856);
nand U1474 (N_1474,In_864,In_115);
nor U1475 (N_1475,In_381,In_586);
nor U1476 (N_1476,In_968,In_702);
xor U1477 (N_1477,In_523,In_251);
xor U1478 (N_1478,In_94,In_596);
nor U1479 (N_1479,In_957,In_722);
xor U1480 (N_1480,In_742,In_799);
nand U1481 (N_1481,In_775,In_404);
nor U1482 (N_1482,In_350,In_518);
nand U1483 (N_1483,In_128,In_808);
nor U1484 (N_1484,In_50,In_394);
and U1485 (N_1485,In_670,In_399);
and U1486 (N_1486,In_839,In_560);
and U1487 (N_1487,In_493,In_811);
and U1488 (N_1488,In_905,In_899);
nand U1489 (N_1489,In_857,In_545);
xnor U1490 (N_1490,In_926,In_729);
or U1491 (N_1491,In_637,In_995);
nand U1492 (N_1492,In_836,In_704);
and U1493 (N_1493,In_610,In_869);
nand U1494 (N_1494,In_586,In_203);
or U1495 (N_1495,In_988,In_117);
or U1496 (N_1496,In_763,In_690);
and U1497 (N_1497,In_341,In_282);
nor U1498 (N_1498,In_324,In_734);
nand U1499 (N_1499,In_151,In_932);
or U1500 (N_1500,In_662,In_902);
or U1501 (N_1501,In_782,In_816);
xor U1502 (N_1502,In_194,In_585);
or U1503 (N_1503,In_205,In_262);
or U1504 (N_1504,In_299,In_674);
xnor U1505 (N_1505,In_524,In_814);
and U1506 (N_1506,In_522,In_297);
and U1507 (N_1507,In_635,In_689);
nor U1508 (N_1508,In_557,In_578);
and U1509 (N_1509,In_400,In_249);
xor U1510 (N_1510,In_631,In_394);
xor U1511 (N_1511,In_757,In_318);
nor U1512 (N_1512,In_221,In_941);
and U1513 (N_1513,In_519,In_771);
nand U1514 (N_1514,In_399,In_643);
nor U1515 (N_1515,In_320,In_101);
and U1516 (N_1516,In_952,In_131);
or U1517 (N_1517,In_948,In_232);
xor U1518 (N_1518,In_168,In_806);
nand U1519 (N_1519,In_620,In_751);
or U1520 (N_1520,In_517,In_294);
or U1521 (N_1521,In_919,In_263);
nand U1522 (N_1522,In_469,In_20);
or U1523 (N_1523,In_73,In_766);
or U1524 (N_1524,In_727,In_45);
and U1525 (N_1525,In_659,In_546);
and U1526 (N_1526,In_404,In_316);
or U1527 (N_1527,In_551,In_156);
or U1528 (N_1528,In_885,In_490);
nand U1529 (N_1529,In_989,In_323);
nand U1530 (N_1530,In_725,In_869);
nor U1531 (N_1531,In_450,In_195);
and U1532 (N_1532,In_943,In_98);
nor U1533 (N_1533,In_572,In_769);
or U1534 (N_1534,In_71,In_762);
and U1535 (N_1535,In_965,In_474);
xnor U1536 (N_1536,In_568,In_899);
nand U1537 (N_1537,In_958,In_891);
nand U1538 (N_1538,In_85,In_196);
nor U1539 (N_1539,In_46,In_534);
nor U1540 (N_1540,In_508,In_555);
or U1541 (N_1541,In_836,In_867);
nand U1542 (N_1542,In_486,In_513);
or U1543 (N_1543,In_205,In_756);
xor U1544 (N_1544,In_855,In_220);
and U1545 (N_1545,In_448,In_269);
nand U1546 (N_1546,In_813,In_752);
nor U1547 (N_1547,In_848,In_858);
nand U1548 (N_1548,In_344,In_418);
nor U1549 (N_1549,In_755,In_251);
or U1550 (N_1550,In_149,In_839);
xnor U1551 (N_1551,In_768,In_774);
and U1552 (N_1552,In_220,In_346);
nand U1553 (N_1553,In_181,In_557);
nor U1554 (N_1554,In_864,In_412);
and U1555 (N_1555,In_432,In_979);
and U1556 (N_1556,In_308,In_980);
and U1557 (N_1557,In_165,In_173);
and U1558 (N_1558,In_891,In_475);
nor U1559 (N_1559,In_914,In_316);
or U1560 (N_1560,In_93,In_591);
and U1561 (N_1561,In_544,In_340);
or U1562 (N_1562,In_800,In_393);
and U1563 (N_1563,In_256,In_754);
nand U1564 (N_1564,In_93,In_903);
and U1565 (N_1565,In_814,In_42);
and U1566 (N_1566,In_450,In_952);
xnor U1567 (N_1567,In_491,In_921);
or U1568 (N_1568,In_772,In_885);
and U1569 (N_1569,In_988,In_753);
nand U1570 (N_1570,In_277,In_352);
and U1571 (N_1571,In_339,In_951);
or U1572 (N_1572,In_913,In_841);
nand U1573 (N_1573,In_386,In_888);
and U1574 (N_1574,In_642,In_31);
nor U1575 (N_1575,In_130,In_783);
nor U1576 (N_1576,In_803,In_358);
or U1577 (N_1577,In_248,In_216);
nor U1578 (N_1578,In_202,In_278);
nor U1579 (N_1579,In_794,In_642);
nand U1580 (N_1580,In_577,In_476);
or U1581 (N_1581,In_811,In_793);
xor U1582 (N_1582,In_659,In_605);
nor U1583 (N_1583,In_725,In_847);
nor U1584 (N_1584,In_529,In_457);
nor U1585 (N_1585,In_632,In_761);
nand U1586 (N_1586,In_135,In_426);
nand U1587 (N_1587,In_487,In_437);
nand U1588 (N_1588,In_333,In_497);
or U1589 (N_1589,In_585,In_25);
nor U1590 (N_1590,In_362,In_7);
nor U1591 (N_1591,In_293,In_481);
nor U1592 (N_1592,In_335,In_841);
nor U1593 (N_1593,In_670,In_892);
xor U1594 (N_1594,In_855,In_982);
or U1595 (N_1595,In_180,In_301);
nor U1596 (N_1596,In_773,In_965);
nand U1597 (N_1597,In_483,In_201);
or U1598 (N_1598,In_359,In_99);
and U1599 (N_1599,In_41,In_481);
and U1600 (N_1600,In_401,In_668);
or U1601 (N_1601,In_325,In_809);
nor U1602 (N_1602,In_754,In_172);
nand U1603 (N_1603,In_689,In_926);
and U1604 (N_1604,In_319,In_580);
or U1605 (N_1605,In_983,In_456);
nor U1606 (N_1606,In_925,In_820);
and U1607 (N_1607,In_41,In_621);
and U1608 (N_1608,In_214,In_754);
and U1609 (N_1609,In_814,In_721);
and U1610 (N_1610,In_320,In_311);
or U1611 (N_1611,In_116,In_426);
and U1612 (N_1612,In_431,In_413);
and U1613 (N_1613,In_716,In_917);
nand U1614 (N_1614,In_577,In_582);
and U1615 (N_1615,In_372,In_114);
nand U1616 (N_1616,In_927,In_52);
or U1617 (N_1617,In_628,In_707);
or U1618 (N_1618,In_274,In_51);
and U1619 (N_1619,In_285,In_303);
xor U1620 (N_1620,In_976,In_137);
and U1621 (N_1621,In_221,In_118);
nand U1622 (N_1622,In_268,In_699);
and U1623 (N_1623,In_467,In_681);
nand U1624 (N_1624,In_201,In_81);
nand U1625 (N_1625,In_48,In_657);
and U1626 (N_1626,In_360,In_91);
nand U1627 (N_1627,In_171,In_41);
nand U1628 (N_1628,In_59,In_123);
nand U1629 (N_1629,In_64,In_25);
nor U1630 (N_1630,In_966,In_197);
nor U1631 (N_1631,In_827,In_517);
or U1632 (N_1632,In_819,In_986);
nor U1633 (N_1633,In_837,In_664);
nor U1634 (N_1634,In_790,In_336);
xor U1635 (N_1635,In_155,In_368);
or U1636 (N_1636,In_538,In_857);
nor U1637 (N_1637,In_45,In_436);
nand U1638 (N_1638,In_545,In_605);
nand U1639 (N_1639,In_228,In_603);
or U1640 (N_1640,In_20,In_772);
and U1641 (N_1641,In_306,In_584);
and U1642 (N_1642,In_72,In_939);
and U1643 (N_1643,In_195,In_994);
and U1644 (N_1644,In_586,In_117);
xnor U1645 (N_1645,In_40,In_592);
and U1646 (N_1646,In_253,In_573);
nor U1647 (N_1647,In_209,In_904);
and U1648 (N_1648,In_549,In_939);
nand U1649 (N_1649,In_691,In_276);
nor U1650 (N_1650,In_660,In_72);
xor U1651 (N_1651,In_228,In_316);
and U1652 (N_1652,In_711,In_767);
nor U1653 (N_1653,In_851,In_538);
nor U1654 (N_1654,In_106,In_845);
or U1655 (N_1655,In_900,In_553);
or U1656 (N_1656,In_427,In_953);
nand U1657 (N_1657,In_311,In_953);
nand U1658 (N_1658,In_135,In_938);
nor U1659 (N_1659,In_798,In_620);
nand U1660 (N_1660,In_240,In_325);
and U1661 (N_1661,In_597,In_755);
nand U1662 (N_1662,In_751,In_76);
xnor U1663 (N_1663,In_238,In_598);
nor U1664 (N_1664,In_88,In_381);
nor U1665 (N_1665,In_527,In_127);
or U1666 (N_1666,In_901,In_843);
nand U1667 (N_1667,In_779,In_44);
and U1668 (N_1668,In_99,In_269);
nand U1669 (N_1669,In_49,In_111);
or U1670 (N_1670,In_83,In_15);
or U1671 (N_1671,In_870,In_318);
nand U1672 (N_1672,In_696,In_97);
nor U1673 (N_1673,In_250,In_410);
and U1674 (N_1674,In_218,In_905);
and U1675 (N_1675,In_919,In_245);
nand U1676 (N_1676,In_846,In_31);
nor U1677 (N_1677,In_553,In_249);
nor U1678 (N_1678,In_170,In_59);
or U1679 (N_1679,In_892,In_368);
or U1680 (N_1680,In_252,In_512);
or U1681 (N_1681,In_52,In_832);
or U1682 (N_1682,In_94,In_114);
or U1683 (N_1683,In_351,In_313);
and U1684 (N_1684,In_0,In_48);
or U1685 (N_1685,In_748,In_620);
nor U1686 (N_1686,In_440,In_668);
nor U1687 (N_1687,In_272,In_701);
xor U1688 (N_1688,In_780,In_356);
nand U1689 (N_1689,In_441,In_39);
or U1690 (N_1690,In_253,In_943);
xor U1691 (N_1691,In_570,In_482);
nor U1692 (N_1692,In_764,In_790);
xor U1693 (N_1693,In_370,In_903);
or U1694 (N_1694,In_280,In_686);
or U1695 (N_1695,In_894,In_611);
or U1696 (N_1696,In_234,In_425);
or U1697 (N_1697,In_544,In_9);
or U1698 (N_1698,In_13,In_540);
and U1699 (N_1699,In_237,In_883);
or U1700 (N_1700,In_894,In_423);
xor U1701 (N_1701,In_325,In_625);
or U1702 (N_1702,In_728,In_885);
and U1703 (N_1703,In_678,In_250);
nand U1704 (N_1704,In_588,In_900);
nand U1705 (N_1705,In_210,In_899);
nor U1706 (N_1706,In_306,In_630);
xnor U1707 (N_1707,In_269,In_148);
or U1708 (N_1708,In_536,In_226);
or U1709 (N_1709,In_875,In_484);
nand U1710 (N_1710,In_280,In_15);
or U1711 (N_1711,In_497,In_866);
xor U1712 (N_1712,In_408,In_680);
or U1713 (N_1713,In_123,In_390);
nand U1714 (N_1714,In_807,In_118);
nand U1715 (N_1715,In_956,In_519);
and U1716 (N_1716,In_42,In_884);
nor U1717 (N_1717,In_37,In_189);
and U1718 (N_1718,In_581,In_921);
xnor U1719 (N_1719,In_530,In_509);
or U1720 (N_1720,In_188,In_64);
nor U1721 (N_1721,In_447,In_285);
nor U1722 (N_1722,In_248,In_29);
nand U1723 (N_1723,In_733,In_645);
nor U1724 (N_1724,In_12,In_699);
nor U1725 (N_1725,In_756,In_355);
nand U1726 (N_1726,In_463,In_584);
nand U1727 (N_1727,In_662,In_533);
nand U1728 (N_1728,In_242,In_726);
nand U1729 (N_1729,In_363,In_174);
nand U1730 (N_1730,In_185,In_944);
or U1731 (N_1731,In_559,In_635);
xnor U1732 (N_1732,In_700,In_225);
and U1733 (N_1733,In_77,In_825);
or U1734 (N_1734,In_603,In_543);
nand U1735 (N_1735,In_589,In_515);
nor U1736 (N_1736,In_122,In_681);
and U1737 (N_1737,In_482,In_889);
nor U1738 (N_1738,In_460,In_117);
nor U1739 (N_1739,In_433,In_798);
or U1740 (N_1740,In_635,In_302);
xnor U1741 (N_1741,In_619,In_291);
or U1742 (N_1742,In_112,In_497);
and U1743 (N_1743,In_775,In_99);
xor U1744 (N_1744,In_89,In_432);
nand U1745 (N_1745,In_443,In_777);
or U1746 (N_1746,In_353,In_255);
or U1747 (N_1747,In_560,In_450);
nor U1748 (N_1748,In_25,In_896);
or U1749 (N_1749,In_504,In_813);
or U1750 (N_1750,In_862,In_195);
or U1751 (N_1751,In_237,In_943);
and U1752 (N_1752,In_559,In_857);
or U1753 (N_1753,In_747,In_684);
nand U1754 (N_1754,In_689,In_289);
or U1755 (N_1755,In_692,In_344);
or U1756 (N_1756,In_555,In_829);
and U1757 (N_1757,In_969,In_360);
or U1758 (N_1758,In_200,In_470);
or U1759 (N_1759,In_367,In_772);
nor U1760 (N_1760,In_507,In_879);
xnor U1761 (N_1761,In_653,In_228);
and U1762 (N_1762,In_809,In_740);
nor U1763 (N_1763,In_697,In_843);
or U1764 (N_1764,In_3,In_751);
nand U1765 (N_1765,In_553,In_952);
nand U1766 (N_1766,In_962,In_542);
or U1767 (N_1767,In_175,In_538);
nand U1768 (N_1768,In_639,In_591);
nand U1769 (N_1769,In_625,In_571);
xor U1770 (N_1770,In_935,In_219);
nand U1771 (N_1771,In_777,In_537);
nand U1772 (N_1772,In_551,In_236);
nor U1773 (N_1773,In_978,In_824);
nand U1774 (N_1774,In_947,In_477);
xor U1775 (N_1775,In_645,In_801);
nor U1776 (N_1776,In_337,In_247);
nand U1777 (N_1777,In_995,In_463);
or U1778 (N_1778,In_883,In_307);
and U1779 (N_1779,In_492,In_656);
or U1780 (N_1780,In_37,In_58);
xor U1781 (N_1781,In_761,In_848);
or U1782 (N_1782,In_883,In_391);
nand U1783 (N_1783,In_474,In_944);
and U1784 (N_1784,In_323,In_379);
or U1785 (N_1785,In_642,In_851);
nand U1786 (N_1786,In_46,In_164);
nand U1787 (N_1787,In_239,In_417);
and U1788 (N_1788,In_811,In_526);
nand U1789 (N_1789,In_762,In_995);
nor U1790 (N_1790,In_182,In_215);
or U1791 (N_1791,In_636,In_429);
or U1792 (N_1792,In_992,In_554);
nand U1793 (N_1793,In_127,In_212);
or U1794 (N_1794,In_934,In_165);
nor U1795 (N_1795,In_559,In_883);
xor U1796 (N_1796,In_187,In_694);
nand U1797 (N_1797,In_524,In_842);
and U1798 (N_1798,In_414,In_779);
nor U1799 (N_1799,In_629,In_486);
xor U1800 (N_1800,In_182,In_801);
and U1801 (N_1801,In_119,In_610);
and U1802 (N_1802,In_561,In_471);
or U1803 (N_1803,In_836,In_686);
nand U1804 (N_1804,In_866,In_311);
nor U1805 (N_1805,In_835,In_465);
and U1806 (N_1806,In_534,In_965);
nor U1807 (N_1807,In_861,In_129);
nor U1808 (N_1808,In_689,In_895);
nand U1809 (N_1809,In_930,In_638);
or U1810 (N_1810,In_702,In_399);
nand U1811 (N_1811,In_757,In_879);
nand U1812 (N_1812,In_316,In_78);
or U1813 (N_1813,In_560,In_847);
or U1814 (N_1814,In_270,In_992);
nor U1815 (N_1815,In_499,In_444);
nor U1816 (N_1816,In_88,In_658);
or U1817 (N_1817,In_57,In_290);
and U1818 (N_1818,In_248,In_399);
nand U1819 (N_1819,In_73,In_426);
or U1820 (N_1820,In_963,In_375);
nor U1821 (N_1821,In_709,In_171);
nor U1822 (N_1822,In_250,In_144);
nand U1823 (N_1823,In_663,In_894);
nor U1824 (N_1824,In_747,In_404);
nand U1825 (N_1825,In_160,In_495);
or U1826 (N_1826,In_78,In_660);
nor U1827 (N_1827,In_370,In_457);
and U1828 (N_1828,In_134,In_511);
or U1829 (N_1829,In_734,In_352);
nor U1830 (N_1830,In_155,In_988);
nor U1831 (N_1831,In_537,In_621);
nor U1832 (N_1832,In_876,In_897);
nor U1833 (N_1833,In_879,In_849);
xnor U1834 (N_1834,In_494,In_673);
or U1835 (N_1835,In_969,In_25);
nor U1836 (N_1836,In_676,In_595);
and U1837 (N_1837,In_194,In_716);
nand U1838 (N_1838,In_977,In_474);
or U1839 (N_1839,In_791,In_971);
or U1840 (N_1840,In_81,In_807);
nor U1841 (N_1841,In_601,In_215);
nand U1842 (N_1842,In_130,In_451);
and U1843 (N_1843,In_235,In_779);
or U1844 (N_1844,In_968,In_59);
and U1845 (N_1845,In_805,In_171);
nor U1846 (N_1846,In_110,In_894);
xnor U1847 (N_1847,In_456,In_761);
nand U1848 (N_1848,In_606,In_707);
nor U1849 (N_1849,In_857,In_904);
xnor U1850 (N_1850,In_267,In_894);
or U1851 (N_1851,In_727,In_218);
xnor U1852 (N_1852,In_329,In_847);
or U1853 (N_1853,In_674,In_325);
nand U1854 (N_1854,In_78,In_590);
and U1855 (N_1855,In_102,In_760);
and U1856 (N_1856,In_745,In_493);
nand U1857 (N_1857,In_718,In_76);
or U1858 (N_1858,In_214,In_285);
and U1859 (N_1859,In_666,In_899);
nand U1860 (N_1860,In_107,In_606);
nand U1861 (N_1861,In_893,In_522);
nand U1862 (N_1862,In_957,In_633);
nand U1863 (N_1863,In_586,In_735);
nor U1864 (N_1864,In_9,In_934);
nor U1865 (N_1865,In_768,In_703);
or U1866 (N_1866,In_557,In_243);
nor U1867 (N_1867,In_529,In_452);
or U1868 (N_1868,In_771,In_563);
and U1869 (N_1869,In_440,In_768);
nor U1870 (N_1870,In_119,In_769);
and U1871 (N_1871,In_566,In_71);
and U1872 (N_1872,In_560,In_671);
and U1873 (N_1873,In_498,In_823);
xnor U1874 (N_1874,In_754,In_451);
nand U1875 (N_1875,In_526,In_592);
nor U1876 (N_1876,In_178,In_467);
and U1877 (N_1877,In_964,In_288);
nor U1878 (N_1878,In_600,In_261);
and U1879 (N_1879,In_499,In_637);
nand U1880 (N_1880,In_663,In_991);
nor U1881 (N_1881,In_98,In_731);
or U1882 (N_1882,In_833,In_473);
nand U1883 (N_1883,In_156,In_365);
nand U1884 (N_1884,In_99,In_942);
nor U1885 (N_1885,In_275,In_641);
and U1886 (N_1886,In_914,In_793);
xnor U1887 (N_1887,In_543,In_354);
nor U1888 (N_1888,In_183,In_940);
xnor U1889 (N_1889,In_793,In_252);
and U1890 (N_1890,In_435,In_406);
and U1891 (N_1891,In_84,In_236);
or U1892 (N_1892,In_128,In_447);
nand U1893 (N_1893,In_456,In_496);
nand U1894 (N_1894,In_660,In_848);
or U1895 (N_1895,In_714,In_951);
nand U1896 (N_1896,In_748,In_553);
and U1897 (N_1897,In_524,In_789);
xor U1898 (N_1898,In_572,In_652);
nor U1899 (N_1899,In_913,In_305);
nand U1900 (N_1900,In_416,In_314);
and U1901 (N_1901,In_632,In_630);
or U1902 (N_1902,In_516,In_512);
nand U1903 (N_1903,In_786,In_43);
and U1904 (N_1904,In_753,In_740);
nor U1905 (N_1905,In_395,In_765);
and U1906 (N_1906,In_511,In_850);
nand U1907 (N_1907,In_526,In_103);
or U1908 (N_1908,In_670,In_946);
nand U1909 (N_1909,In_769,In_805);
xor U1910 (N_1910,In_527,In_874);
xor U1911 (N_1911,In_667,In_705);
and U1912 (N_1912,In_438,In_128);
or U1913 (N_1913,In_369,In_182);
nand U1914 (N_1914,In_770,In_297);
and U1915 (N_1915,In_777,In_361);
nand U1916 (N_1916,In_414,In_389);
and U1917 (N_1917,In_885,In_268);
and U1918 (N_1918,In_88,In_106);
or U1919 (N_1919,In_573,In_586);
or U1920 (N_1920,In_322,In_835);
nand U1921 (N_1921,In_416,In_262);
nand U1922 (N_1922,In_551,In_813);
nand U1923 (N_1923,In_668,In_847);
nand U1924 (N_1924,In_92,In_938);
and U1925 (N_1925,In_117,In_174);
nor U1926 (N_1926,In_878,In_141);
and U1927 (N_1927,In_682,In_314);
nor U1928 (N_1928,In_467,In_943);
or U1929 (N_1929,In_814,In_843);
or U1930 (N_1930,In_234,In_8);
nor U1931 (N_1931,In_318,In_195);
or U1932 (N_1932,In_823,In_845);
nand U1933 (N_1933,In_69,In_316);
or U1934 (N_1934,In_984,In_297);
nor U1935 (N_1935,In_638,In_175);
or U1936 (N_1936,In_291,In_233);
nand U1937 (N_1937,In_142,In_601);
or U1938 (N_1938,In_259,In_270);
and U1939 (N_1939,In_18,In_711);
and U1940 (N_1940,In_874,In_159);
nor U1941 (N_1941,In_860,In_0);
nand U1942 (N_1942,In_361,In_267);
nor U1943 (N_1943,In_274,In_806);
or U1944 (N_1944,In_845,In_467);
and U1945 (N_1945,In_186,In_832);
or U1946 (N_1946,In_21,In_966);
and U1947 (N_1947,In_922,In_791);
nor U1948 (N_1948,In_805,In_7);
and U1949 (N_1949,In_534,In_285);
nand U1950 (N_1950,In_554,In_659);
nor U1951 (N_1951,In_728,In_288);
and U1952 (N_1952,In_993,In_366);
or U1953 (N_1953,In_781,In_910);
nor U1954 (N_1954,In_593,In_753);
or U1955 (N_1955,In_322,In_924);
and U1956 (N_1956,In_270,In_699);
xor U1957 (N_1957,In_646,In_841);
or U1958 (N_1958,In_562,In_193);
or U1959 (N_1959,In_860,In_409);
and U1960 (N_1960,In_388,In_238);
nor U1961 (N_1961,In_570,In_392);
nor U1962 (N_1962,In_348,In_113);
nor U1963 (N_1963,In_844,In_718);
and U1964 (N_1964,In_704,In_738);
and U1965 (N_1965,In_307,In_305);
or U1966 (N_1966,In_685,In_991);
nor U1967 (N_1967,In_335,In_346);
nand U1968 (N_1968,In_730,In_408);
nand U1969 (N_1969,In_275,In_473);
or U1970 (N_1970,In_991,In_453);
xor U1971 (N_1971,In_399,In_874);
nor U1972 (N_1972,In_279,In_126);
xor U1973 (N_1973,In_702,In_811);
or U1974 (N_1974,In_708,In_403);
nor U1975 (N_1975,In_208,In_968);
nand U1976 (N_1976,In_113,In_353);
nor U1977 (N_1977,In_303,In_344);
or U1978 (N_1978,In_320,In_102);
or U1979 (N_1979,In_236,In_933);
nand U1980 (N_1980,In_986,In_310);
xor U1981 (N_1981,In_237,In_698);
xor U1982 (N_1982,In_968,In_5);
nand U1983 (N_1983,In_968,In_482);
or U1984 (N_1984,In_283,In_612);
nor U1985 (N_1985,In_133,In_449);
and U1986 (N_1986,In_418,In_600);
nor U1987 (N_1987,In_696,In_776);
nor U1988 (N_1988,In_667,In_8);
and U1989 (N_1989,In_210,In_129);
or U1990 (N_1990,In_922,In_599);
nor U1991 (N_1991,In_404,In_39);
nor U1992 (N_1992,In_700,In_141);
and U1993 (N_1993,In_327,In_383);
and U1994 (N_1994,In_859,In_107);
or U1995 (N_1995,In_820,In_838);
and U1996 (N_1996,In_449,In_696);
or U1997 (N_1997,In_153,In_869);
or U1998 (N_1998,In_386,In_443);
xor U1999 (N_1999,In_818,In_32);
or U2000 (N_2000,In_93,In_70);
nor U2001 (N_2001,In_426,In_126);
and U2002 (N_2002,In_640,In_562);
nor U2003 (N_2003,In_589,In_697);
nor U2004 (N_2004,In_914,In_391);
and U2005 (N_2005,In_237,In_406);
xnor U2006 (N_2006,In_194,In_226);
nor U2007 (N_2007,In_656,In_765);
nand U2008 (N_2008,In_846,In_49);
or U2009 (N_2009,In_229,In_929);
nor U2010 (N_2010,In_171,In_184);
and U2011 (N_2011,In_393,In_392);
or U2012 (N_2012,In_125,In_451);
nor U2013 (N_2013,In_753,In_838);
nor U2014 (N_2014,In_503,In_612);
nor U2015 (N_2015,In_671,In_167);
nor U2016 (N_2016,In_415,In_111);
and U2017 (N_2017,In_373,In_31);
and U2018 (N_2018,In_154,In_132);
and U2019 (N_2019,In_334,In_742);
and U2020 (N_2020,In_377,In_935);
nor U2021 (N_2021,In_873,In_156);
nor U2022 (N_2022,In_191,In_315);
nand U2023 (N_2023,In_629,In_981);
nor U2024 (N_2024,In_762,In_972);
or U2025 (N_2025,In_770,In_314);
or U2026 (N_2026,In_810,In_354);
nor U2027 (N_2027,In_155,In_666);
nand U2028 (N_2028,In_852,In_421);
and U2029 (N_2029,In_569,In_988);
and U2030 (N_2030,In_804,In_112);
nand U2031 (N_2031,In_224,In_791);
nand U2032 (N_2032,In_693,In_163);
and U2033 (N_2033,In_28,In_413);
or U2034 (N_2034,In_421,In_822);
nor U2035 (N_2035,In_869,In_853);
and U2036 (N_2036,In_615,In_393);
xor U2037 (N_2037,In_553,In_270);
or U2038 (N_2038,In_684,In_612);
or U2039 (N_2039,In_348,In_600);
nand U2040 (N_2040,In_734,In_881);
xor U2041 (N_2041,In_213,In_400);
nand U2042 (N_2042,In_78,In_103);
or U2043 (N_2043,In_886,In_777);
and U2044 (N_2044,In_660,In_755);
and U2045 (N_2045,In_465,In_468);
or U2046 (N_2046,In_112,In_947);
or U2047 (N_2047,In_567,In_254);
nand U2048 (N_2048,In_783,In_582);
nor U2049 (N_2049,In_647,In_744);
and U2050 (N_2050,In_948,In_641);
nand U2051 (N_2051,In_333,In_139);
nor U2052 (N_2052,In_549,In_221);
and U2053 (N_2053,In_986,In_218);
nor U2054 (N_2054,In_858,In_49);
nand U2055 (N_2055,In_31,In_687);
nand U2056 (N_2056,In_448,In_586);
nor U2057 (N_2057,In_15,In_174);
and U2058 (N_2058,In_284,In_130);
xor U2059 (N_2059,In_243,In_633);
xor U2060 (N_2060,In_46,In_457);
nand U2061 (N_2061,In_987,In_477);
and U2062 (N_2062,In_857,In_890);
nand U2063 (N_2063,In_772,In_459);
and U2064 (N_2064,In_66,In_126);
nand U2065 (N_2065,In_960,In_367);
and U2066 (N_2066,In_477,In_112);
or U2067 (N_2067,In_661,In_575);
or U2068 (N_2068,In_904,In_37);
and U2069 (N_2069,In_563,In_940);
and U2070 (N_2070,In_105,In_573);
or U2071 (N_2071,In_478,In_807);
or U2072 (N_2072,In_16,In_328);
and U2073 (N_2073,In_512,In_860);
xor U2074 (N_2074,In_649,In_61);
or U2075 (N_2075,In_146,In_892);
and U2076 (N_2076,In_981,In_261);
nand U2077 (N_2077,In_491,In_163);
or U2078 (N_2078,In_974,In_308);
nor U2079 (N_2079,In_703,In_890);
nand U2080 (N_2080,In_957,In_617);
nand U2081 (N_2081,In_265,In_277);
nand U2082 (N_2082,In_619,In_463);
and U2083 (N_2083,In_259,In_353);
or U2084 (N_2084,In_486,In_49);
nand U2085 (N_2085,In_749,In_4);
nor U2086 (N_2086,In_580,In_61);
and U2087 (N_2087,In_227,In_556);
or U2088 (N_2088,In_546,In_696);
nor U2089 (N_2089,In_38,In_566);
nor U2090 (N_2090,In_419,In_125);
nor U2091 (N_2091,In_813,In_978);
and U2092 (N_2092,In_677,In_764);
nand U2093 (N_2093,In_847,In_667);
xor U2094 (N_2094,In_235,In_928);
and U2095 (N_2095,In_460,In_91);
or U2096 (N_2096,In_251,In_917);
nor U2097 (N_2097,In_116,In_840);
nand U2098 (N_2098,In_783,In_515);
and U2099 (N_2099,In_466,In_331);
and U2100 (N_2100,In_561,In_726);
xor U2101 (N_2101,In_505,In_790);
nor U2102 (N_2102,In_236,In_894);
or U2103 (N_2103,In_558,In_125);
nor U2104 (N_2104,In_848,In_662);
nand U2105 (N_2105,In_101,In_17);
nor U2106 (N_2106,In_761,In_810);
or U2107 (N_2107,In_901,In_367);
nor U2108 (N_2108,In_516,In_900);
or U2109 (N_2109,In_9,In_260);
nand U2110 (N_2110,In_669,In_790);
nand U2111 (N_2111,In_729,In_676);
xnor U2112 (N_2112,In_28,In_838);
or U2113 (N_2113,In_25,In_96);
or U2114 (N_2114,In_33,In_353);
and U2115 (N_2115,In_550,In_639);
or U2116 (N_2116,In_906,In_194);
nand U2117 (N_2117,In_110,In_828);
xor U2118 (N_2118,In_125,In_792);
nand U2119 (N_2119,In_525,In_684);
nor U2120 (N_2120,In_854,In_724);
and U2121 (N_2121,In_598,In_828);
nand U2122 (N_2122,In_153,In_509);
and U2123 (N_2123,In_401,In_844);
nor U2124 (N_2124,In_509,In_692);
and U2125 (N_2125,In_666,In_281);
nor U2126 (N_2126,In_331,In_964);
or U2127 (N_2127,In_86,In_222);
nor U2128 (N_2128,In_4,In_508);
nor U2129 (N_2129,In_534,In_274);
and U2130 (N_2130,In_65,In_989);
nor U2131 (N_2131,In_85,In_283);
nand U2132 (N_2132,In_759,In_955);
and U2133 (N_2133,In_654,In_754);
or U2134 (N_2134,In_296,In_208);
xor U2135 (N_2135,In_158,In_834);
nand U2136 (N_2136,In_11,In_577);
and U2137 (N_2137,In_716,In_94);
and U2138 (N_2138,In_948,In_268);
nand U2139 (N_2139,In_771,In_997);
xnor U2140 (N_2140,In_302,In_149);
or U2141 (N_2141,In_721,In_316);
nor U2142 (N_2142,In_850,In_170);
nor U2143 (N_2143,In_519,In_105);
nand U2144 (N_2144,In_941,In_329);
nand U2145 (N_2145,In_646,In_842);
nor U2146 (N_2146,In_439,In_3);
and U2147 (N_2147,In_501,In_226);
or U2148 (N_2148,In_901,In_929);
xnor U2149 (N_2149,In_882,In_713);
or U2150 (N_2150,In_272,In_470);
or U2151 (N_2151,In_428,In_55);
nand U2152 (N_2152,In_762,In_933);
and U2153 (N_2153,In_122,In_317);
nor U2154 (N_2154,In_100,In_318);
nand U2155 (N_2155,In_692,In_685);
and U2156 (N_2156,In_563,In_846);
nand U2157 (N_2157,In_20,In_244);
xnor U2158 (N_2158,In_600,In_793);
nor U2159 (N_2159,In_258,In_453);
xnor U2160 (N_2160,In_922,In_873);
and U2161 (N_2161,In_52,In_326);
nor U2162 (N_2162,In_533,In_119);
nor U2163 (N_2163,In_542,In_537);
or U2164 (N_2164,In_392,In_286);
and U2165 (N_2165,In_686,In_644);
or U2166 (N_2166,In_182,In_797);
nor U2167 (N_2167,In_811,In_373);
or U2168 (N_2168,In_562,In_639);
nor U2169 (N_2169,In_571,In_462);
nand U2170 (N_2170,In_73,In_489);
nor U2171 (N_2171,In_644,In_723);
nor U2172 (N_2172,In_130,In_291);
xnor U2173 (N_2173,In_515,In_765);
or U2174 (N_2174,In_250,In_829);
nand U2175 (N_2175,In_592,In_323);
xnor U2176 (N_2176,In_411,In_278);
and U2177 (N_2177,In_768,In_971);
or U2178 (N_2178,In_125,In_462);
or U2179 (N_2179,In_688,In_22);
or U2180 (N_2180,In_322,In_229);
and U2181 (N_2181,In_348,In_236);
or U2182 (N_2182,In_367,In_521);
or U2183 (N_2183,In_689,In_88);
or U2184 (N_2184,In_499,In_672);
nand U2185 (N_2185,In_801,In_598);
and U2186 (N_2186,In_399,In_733);
xor U2187 (N_2187,In_53,In_643);
nand U2188 (N_2188,In_399,In_906);
nand U2189 (N_2189,In_334,In_493);
or U2190 (N_2190,In_520,In_167);
nand U2191 (N_2191,In_66,In_99);
or U2192 (N_2192,In_837,In_431);
nand U2193 (N_2193,In_175,In_967);
and U2194 (N_2194,In_851,In_163);
nor U2195 (N_2195,In_560,In_914);
nor U2196 (N_2196,In_745,In_136);
nand U2197 (N_2197,In_203,In_646);
nor U2198 (N_2198,In_473,In_24);
or U2199 (N_2199,In_585,In_968);
or U2200 (N_2200,In_357,In_935);
nand U2201 (N_2201,In_256,In_478);
nor U2202 (N_2202,In_831,In_464);
nand U2203 (N_2203,In_118,In_510);
and U2204 (N_2204,In_115,In_754);
nor U2205 (N_2205,In_68,In_348);
and U2206 (N_2206,In_813,In_403);
and U2207 (N_2207,In_792,In_160);
or U2208 (N_2208,In_703,In_581);
nor U2209 (N_2209,In_329,In_153);
or U2210 (N_2210,In_304,In_610);
and U2211 (N_2211,In_134,In_311);
and U2212 (N_2212,In_984,In_422);
nor U2213 (N_2213,In_68,In_249);
or U2214 (N_2214,In_657,In_292);
or U2215 (N_2215,In_696,In_484);
nand U2216 (N_2216,In_983,In_878);
and U2217 (N_2217,In_315,In_104);
and U2218 (N_2218,In_627,In_246);
or U2219 (N_2219,In_787,In_338);
nor U2220 (N_2220,In_262,In_932);
and U2221 (N_2221,In_849,In_793);
or U2222 (N_2222,In_630,In_784);
or U2223 (N_2223,In_708,In_604);
xnor U2224 (N_2224,In_919,In_231);
nand U2225 (N_2225,In_212,In_3);
nor U2226 (N_2226,In_608,In_215);
or U2227 (N_2227,In_735,In_289);
nand U2228 (N_2228,In_80,In_481);
or U2229 (N_2229,In_753,In_237);
nor U2230 (N_2230,In_770,In_990);
nand U2231 (N_2231,In_543,In_727);
and U2232 (N_2232,In_806,In_971);
or U2233 (N_2233,In_638,In_497);
and U2234 (N_2234,In_530,In_460);
and U2235 (N_2235,In_712,In_170);
nand U2236 (N_2236,In_179,In_928);
and U2237 (N_2237,In_23,In_313);
and U2238 (N_2238,In_89,In_183);
nor U2239 (N_2239,In_318,In_780);
and U2240 (N_2240,In_790,In_927);
nand U2241 (N_2241,In_563,In_671);
xor U2242 (N_2242,In_886,In_888);
nor U2243 (N_2243,In_469,In_145);
xnor U2244 (N_2244,In_93,In_57);
and U2245 (N_2245,In_862,In_754);
nor U2246 (N_2246,In_428,In_278);
and U2247 (N_2247,In_281,In_276);
nor U2248 (N_2248,In_724,In_398);
and U2249 (N_2249,In_770,In_878);
xor U2250 (N_2250,In_84,In_196);
and U2251 (N_2251,In_872,In_846);
and U2252 (N_2252,In_706,In_871);
xnor U2253 (N_2253,In_254,In_325);
nor U2254 (N_2254,In_291,In_659);
nand U2255 (N_2255,In_631,In_169);
nand U2256 (N_2256,In_895,In_837);
nand U2257 (N_2257,In_141,In_839);
and U2258 (N_2258,In_600,In_361);
and U2259 (N_2259,In_891,In_391);
nand U2260 (N_2260,In_323,In_731);
and U2261 (N_2261,In_604,In_56);
and U2262 (N_2262,In_925,In_19);
or U2263 (N_2263,In_423,In_294);
and U2264 (N_2264,In_45,In_614);
and U2265 (N_2265,In_251,In_11);
nor U2266 (N_2266,In_6,In_291);
nand U2267 (N_2267,In_493,In_760);
or U2268 (N_2268,In_29,In_471);
nand U2269 (N_2269,In_687,In_810);
or U2270 (N_2270,In_977,In_994);
and U2271 (N_2271,In_621,In_278);
or U2272 (N_2272,In_935,In_25);
and U2273 (N_2273,In_214,In_950);
and U2274 (N_2274,In_143,In_438);
nand U2275 (N_2275,In_580,In_71);
or U2276 (N_2276,In_66,In_959);
and U2277 (N_2277,In_921,In_238);
nor U2278 (N_2278,In_603,In_308);
nor U2279 (N_2279,In_670,In_63);
or U2280 (N_2280,In_60,In_52);
nor U2281 (N_2281,In_370,In_73);
nand U2282 (N_2282,In_969,In_643);
nor U2283 (N_2283,In_475,In_227);
and U2284 (N_2284,In_29,In_903);
and U2285 (N_2285,In_913,In_283);
or U2286 (N_2286,In_764,In_975);
or U2287 (N_2287,In_207,In_204);
or U2288 (N_2288,In_797,In_889);
and U2289 (N_2289,In_966,In_620);
nand U2290 (N_2290,In_643,In_391);
nor U2291 (N_2291,In_552,In_867);
nand U2292 (N_2292,In_352,In_758);
xor U2293 (N_2293,In_507,In_597);
nand U2294 (N_2294,In_630,In_569);
and U2295 (N_2295,In_603,In_745);
or U2296 (N_2296,In_670,In_770);
and U2297 (N_2297,In_222,In_633);
nor U2298 (N_2298,In_875,In_348);
xor U2299 (N_2299,In_623,In_64);
xnor U2300 (N_2300,In_880,In_845);
nand U2301 (N_2301,In_775,In_791);
xnor U2302 (N_2302,In_721,In_799);
nor U2303 (N_2303,In_460,In_883);
nor U2304 (N_2304,In_128,In_673);
nand U2305 (N_2305,In_858,In_806);
or U2306 (N_2306,In_859,In_932);
or U2307 (N_2307,In_58,In_539);
nand U2308 (N_2308,In_133,In_91);
nor U2309 (N_2309,In_666,In_847);
or U2310 (N_2310,In_587,In_552);
nand U2311 (N_2311,In_775,In_601);
nor U2312 (N_2312,In_171,In_455);
nor U2313 (N_2313,In_68,In_684);
nor U2314 (N_2314,In_516,In_146);
and U2315 (N_2315,In_127,In_15);
or U2316 (N_2316,In_990,In_178);
or U2317 (N_2317,In_248,In_260);
nand U2318 (N_2318,In_336,In_187);
nor U2319 (N_2319,In_30,In_7);
xnor U2320 (N_2320,In_80,In_784);
and U2321 (N_2321,In_812,In_884);
or U2322 (N_2322,In_132,In_353);
nor U2323 (N_2323,In_199,In_137);
xnor U2324 (N_2324,In_939,In_875);
nand U2325 (N_2325,In_200,In_619);
and U2326 (N_2326,In_43,In_591);
and U2327 (N_2327,In_840,In_873);
and U2328 (N_2328,In_417,In_912);
and U2329 (N_2329,In_338,In_902);
or U2330 (N_2330,In_750,In_747);
or U2331 (N_2331,In_112,In_114);
nor U2332 (N_2332,In_629,In_714);
nand U2333 (N_2333,In_471,In_969);
nand U2334 (N_2334,In_185,In_793);
nor U2335 (N_2335,In_60,In_823);
and U2336 (N_2336,In_884,In_247);
xnor U2337 (N_2337,In_895,In_22);
and U2338 (N_2338,In_124,In_547);
nand U2339 (N_2339,In_433,In_390);
or U2340 (N_2340,In_197,In_390);
or U2341 (N_2341,In_359,In_612);
and U2342 (N_2342,In_680,In_211);
nor U2343 (N_2343,In_515,In_340);
nand U2344 (N_2344,In_915,In_151);
or U2345 (N_2345,In_49,In_205);
nor U2346 (N_2346,In_646,In_132);
or U2347 (N_2347,In_550,In_581);
nor U2348 (N_2348,In_877,In_375);
xnor U2349 (N_2349,In_999,In_942);
or U2350 (N_2350,In_387,In_889);
or U2351 (N_2351,In_893,In_313);
and U2352 (N_2352,In_797,In_774);
and U2353 (N_2353,In_478,In_513);
or U2354 (N_2354,In_778,In_312);
and U2355 (N_2355,In_492,In_434);
or U2356 (N_2356,In_489,In_115);
and U2357 (N_2357,In_63,In_967);
nor U2358 (N_2358,In_119,In_954);
nor U2359 (N_2359,In_411,In_583);
nand U2360 (N_2360,In_309,In_252);
or U2361 (N_2361,In_889,In_711);
nor U2362 (N_2362,In_796,In_390);
or U2363 (N_2363,In_390,In_198);
nor U2364 (N_2364,In_539,In_475);
or U2365 (N_2365,In_609,In_770);
and U2366 (N_2366,In_773,In_750);
nor U2367 (N_2367,In_634,In_999);
xor U2368 (N_2368,In_724,In_532);
and U2369 (N_2369,In_468,In_143);
or U2370 (N_2370,In_708,In_419);
nor U2371 (N_2371,In_914,In_305);
and U2372 (N_2372,In_968,In_366);
or U2373 (N_2373,In_469,In_987);
nand U2374 (N_2374,In_756,In_485);
nor U2375 (N_2375,In_965,In_199);
and U2376 (N_2376,In_462,In_160);
nand U2377 (N_2377,In_23,In_467);
or U2378 (N_2378,In_689,In_201);
nor U2379 (N_2379,In_358,In_80);
nand U2380 (N_2380,In_426,In_892);
and U2381 (N_2381,In_494,In_374);
and U2382 (N_2382,In_976,In_241);
and U2383 (N_2383,In_127,In_816);
nand U2384 (N_2384,In_92,In_463);
and U2385 (N_2385,In_165,In_168);
nand U2386 (N_2386,In_149,In_169);
xnor U2387 (N_2387,In_639,In_754);
or U2388 (N_2388,In_138,In_354);
and U2389 (N_2389,In_330,In_567);
xnor U2390 (N_2390,In_540,In_201);
xor U2391 (N_2391,In_251,In_125);
nand U2392 (N_2392,In_822,In_747);
nand U2393 (N_2393,In_617,In_536);
xor U2394 (N_2394,In_508,In_205);
and U2395 (N_2395,In_863,In_621);
nor U2396 (N_2396,In_869,In_860);
nand U2397 (N_2397,In_546,In_284);
nand U2398 (N_2398,In_595,In_231);
and U2399 (N_2399,In_498,In_413);
nor U2400 (N_2400,In_414,In_142);
or U2401 (N_2401,In_916,In_658);
and U2402 (N_2402,In_459,In_553);
and U2403 (N_2403,In_454,In_557);
nor U2404 (N_2404,In_441,In_673);
or U2405 (N_2405,In_696,In_56);
or U2406 (N_2406,In_67,In_492);
nand U2407 (N_2407,In_683,In_458);
nand U2408 (N_2408,In_677,In_549);
or U2409 (N_2409,In_945,In_529);
xnor U2410 (N_2410,In_835,In_826);
nor U2411 (N_2411,In_117,In_672);
and U2412 (N_2412,In_514,In_37);
and U2413 (N_2413,In_739,In_294);
or U2414 (N_2414,In_907,In_160);
nor U2415 (N_2415,In_596,In_291);
xnor U2416 (N_2416,In_137,In_862);
and U2417 (N_2417,In_541,In_537);
nand U2418 (N_2418,In_100,In_745);
nand U2419 (N_2419,In_45,In_878);
nand U2420 (N_2420,In_133,In_658);
xor U2421 (N_2421,In_664,In_261);
nor U2422 (N_2422,In_264,In_809);
or U2423 (N_2423,In_429,In_871);
or U2424 (N_2424,In_386,In_152);
nor U2425 (N_2425,In_628,In_646);
nor U2426 (N_2426,In_418,In_867);
nand U2427 (N_2427,In_348,In_823);
or U2428 (N_2428,In_835,In_444);
nand U2429 (N_2429,In_695,In_476);
and U2430 (N_2430,In_378,In_445);
or U2431 (N_2431,In_204,In_314);
and U2432 (N_2432,In_13,In_181);
nand U2433 (N_2433,In_660,In_179);
nand U2434 (N_2434,In_709,In_309);
nand U2435 (N_2435,In_127,In_680);
xor U2436 (N_2436,In_910,In_637);
nor U2437 (N_2437,In_933,In_646);
xnor U2438 (N_2438,In_364,In_455);
nor U2439 (N_2439,In_647,In_760);
or U2440 (N_2440,In_676,In_925);
nand U2441 (N_2441,In_417,In_426);
nor U2442 (N_2442,In_804,In_59);
nand U2443 (N_2443,In_92,In_641);
or U2444 (N_2444,In_188,In_397);
and U2445 (N_2445,In_508,In_261);
nand U2446 (N_2446,In_898,In_706);
or U2447 (N_2447,In_274,In_129);
and U2448 (N_2448,In_456,In_154);
nand U2449 (N_2449,In_829,In_926);
or U2450 (N_2450,In_163,In_240);
xor U2451 (N_2451,In_506,In_818);
nor U2452 (N_2452,In_337,In_285);
xor U2453 (N_2453,In_329,In_266);
and U2454 (N_2454,In_326,In_44);
and U2455 (N_2455,In_158,In_115);
nor U2456 (N_2456,In_613,In_507);
and U2457 (N_2457,In_407,In_967);
nor U2458 (N_2458,In_91,In_586);
or U2459 (N_2459,In_559,In_744);
nor U2460 (N_2460,In_600,In_415);
and U2461 (N_2461,In_337,In_826);
and U2462 (N_2462,In_265,In_219);
and U2463 (N_2463,In_819,In_590);
and U2464 (N_2464,In_983,In_555);
and U2465 (N_2465,In_59,In_502);
and U2466 (N_2466,In_760,In_691);
or U2467 (N_2467,In_5,In_457);
xor U2468 (N_2468,In_985,In_663);
nor U2469 (N_2469,In_479,In_796);
nor U2470 (N_2470,In_709,In_970);
nor U2471 (N_2471,In_333,In_513);
or U2472 (N_2472,In_935,In_230);
nor U2473 (N_2473,In_673,In_375);
nor U2474 (N_2474,In_439,In_832);
xor U2475 (N_2475,In_16,In_667);
nand U2476 (N_2476,In_288,In_225);
nor U2477 (N_2477,In_63,In_442);
nand U2478 (N_2478,In_43,In_485);
or U2479 (N_2479,In_833,In_153);
nor U2480 (N_2480,In_197,In_29);
or U2481 (N_2481,In_978,In_419);
nand U2482 (N_2482,In_251,In_327);
nand U2483 (N_2483,In_893,In_882);
nor U2484 (N_2484,In_326,In_324);
and U2485 (N_2485,In_76,In_899);
nand U2486 (N_2486,In_577,In_721);
nand U2487 (N_2487,In_960,In_117);
or U2488 (N_2488,In_931,In_659);
xnor U2489 (N_2489,In_364,In_148);
nand U2490 (N_2490,In_914,In_748);
or U2491 (N_2491,In_992,In_0);
or U2492 (N_2492,In_458,In_598);
or U2493 (N_2493,In_604,In_386);
and U2494 (N_2494,In_990,In_978);
nand U2495 (N_2495,In_157,In_789);
nor U2496 (N_2496,In_613,In_931);
nor U2497 (N_2497,In_960,In_991);
and U2498 (N_2498,In_494,In_679);
or U2499 (N_2499,In_217,In_772);
xor U2500 (N_2500,N_2442,N_1404);
and U2501 (N_2501,N_1625,N_2193);
xnor U2502 (N_2502,N_370,N_544);
nand U2503 (N_2503,N_1275,N_2123);
nand U2504 (N_2504,N_1400,N_1862);
or U2505 (N_2505,N_1469,N_1656);
nor U2506 (N_2506,N_2225,N_386);
nand U2507 (N_2507,N_712,N_581);
nor U2508 (N_2508,N_1326,N_1977);
xnor U2509 (N_2509,N_625,N_1238);
and U2510 (N_2510,N_909,N_1287);
or U2511 (N_2511,N_1421,N_1127);
or U2512 (N_2512,N_2400,N_1848);
nand U2513 (N_2513,N_1813,N_528);
or U2514 (N_2514,N_1909,N_2095);
and U2515 (N_2515,N_2086,N_311);
or U2516 (N_2516,N_2151,N_526);
or U2517 (N_2517,N_1787,N_1117);
nand U2518 (N_2518,N_1626,N_315);
or U2519 (N_2519,N_2424,N_1752);
xor U2520 (N_2520,N_1145,N_680);
or U2521 (N_2521,N_1286,N_551);
and U2522 (N_2522,N_2322,N_1415);
or U2523 (N_2523,N_966,N_2468);
nand U2524 (N_2524,N_1964,N_202);
nand U2525 (N_2525,N_749,N_1191);
or U2526 (N_2526,N_233,N_1076);
xor U2527 (N_2527,N_732,N_572);
or U2528 (N_2528,N_613,N_1083);
nand U2529 (N_2529,N_1256,N_49);
or U2530 (N_2530,N_1785,N_21);
and U2531 (N_2531,N_1241,N_1913);
nor U2532 (N_2532,N_574,N_1587);
nor U2533 (N_2533,N_675,N_1673);
nor U2534 (N_2534,N_2447,N_1726);
or U2535 (N_2535,N_1381,N_1608);
nand U2536 (N_2536,N_449,N_1430);
nand U2537 (N_2537,N_2002,N_1288);
nor U2538 (N_2538,N_2155,N_2279);
nor U2539 (N_2539,N_1747,N_1619);
or U2540 (N_2540,N_100,N_542);
nor U2541 (N_2541,N_145,N_1249);
nor U2542 (N_2542,N_2104,N_501);
nor U2543 (N_2543,N_2334,N_1121);
or U2544 (N_2544,N_1259,N_1035);
nor U2545 (N_2545,N_231,N_986);
nand U2546 (N_2546,N_2194,N_18);
nand U2547 (N_2547,N_1302,N_2197);
or U2548 (N_2548,N_663,N_1480);
nand U2549 (N_2549,N_1571,N_2412);
xnor U2550 (N_2550,N_1953,N_1552);
or U2551 (N_2551,N_1272,N_1965);
or U2552 (N_2552,N_1152,N_652);
nand U2553 (N_2553,N_1359,N_2467);
or U2554 (N_2554,N_2379,N_2129);
nand U2555 (N_2555,N_2287,N_1081);
nand U2556 (N_2556,N_277,N_2061);
and U2557 (N_2557,N_2032,N_1473);
xnor U2558 (N_2558,N_890,N_1157);
xnor U2559 (N_2559,N_1589,N_1845);
nand U2560 (N_2560,N_842,N_320);
nand U2561 (N_2561,N_855,N_2212);
or U2562 (N_2562,N_1350,N_1684);
and U2563 (N_2563,N_1703,N_460);
nand U2564 (N_2564,N_352,N_1522);
nand U2565 (N_2565,N_785,N_1910);
nand U2566 (N_2566,N_1919,N_2219);
xnor U2567 (N_2567,N_2049,N_838);
or U2568 (N_2568,N_2033,N_885);
and U2569 (N_2569,N_760,N_371);
or U2570 (N_2570,N_863,N_1495);
nor U2571 (N_2571,N_390,N_467);
and U2572 (N_2572,N_281,N_183);
nor U2573 (N_2573,N_2016,N_951);
and U2574 (N_2574,N_1979,N_1820);
nor U2575 (N_2575,N_2476,N_942);
or U2576 (N_2576,N_223,N_331);
nand U2577 (N_2577,N_1050,N_201);
xnor U2578 (N_2578,N_235,N_1038);
nor U2579 (N_2579,N_2118,N_1100);
or U2580 (N_2580,N_2485,N_631);
and U2581 (N_2581,N_1023,N_37);
or U2582 (N_2582,N_679,N_2135);
nand U2583 (N_2583,N_1044,N_102);
nor U2584 (N_2584,N_2042,N_2472);
and U2585 (N_2585,N_1190,N_1055);
and U2586 (N_2586,N_546,N_784);
and U2587 (N_2587,N_23,N_2186);
nand U2588 (N_2588,N_534,N_744);
or U2589 (N_2589,N_2143,N_128);
and U2590 (N_2590,N_975,N_729);
nor U2591 (N_2591,N_1576,N_1304);
nand U2592 (N_2592,N_1340,N_2388);
and U2593 (N_2593,N_820,N_1941);
xor U2594 (N_2594,N_766,N_1823);
and U2595 (N_2595,N_2237,N_1322);
nand U2596 (N_2596,N_1908,N_595);
nand U2597 (N_2597,N_2222,N_219);
nand U2598 (N_2598,N_2463,N_126);
and U2599 (N_2599,N_374,N_1419);
or U2600 (N_2600,N_1770,N_105);
or U2601 (N_2601,N_358,N_213);
nand U2602 (N_2602,N_2304,N_398);
nand U2603 (N_2603,N_670,N_1349);
and U2604 (N_2604,N_834,N_2266);
xor U2605 (N_2605,N_167,N_565);
nor U2606 (N_2606,N_1889,N_997);
nand U2607 (N_2607,N_1895,N_416);
or U2608 (N_2608,N_43,N_1344);
or U2609 (N_2609,N_336,N_661);
xnor U2610 (N_2610,N_718,N_653);
and U2611 (N_2611,N_2403,N_1174);
xnor U2612 (N_2612,N_249,N_893);
or U2613 (N_2613,N_697,N_2183);
or U2614 (N_2614,N_1244,N_739);
xnor U2615 (N_2615,N_271,N_1519);
or U2616 (N_2616,N_1338,N_1637);
xnor U2617 (N_2617,N_1588,N_2167);
nor U2618 (N_2618,N_2305,N_2079);
or U2619 (N_2619,N_1666,N_112);
nand U2620 (N_2620,N_325,N_1330);
or U2621 (N_2621,N_2383,N_1741);
or U2622 (N_2622,N_1939,N_89);
or U2623 (N_2623,N_547,N_907);
nand U2624 (N_2624,N_500,N_1136);
nor U2625 (N_2625,N_304,N_1636);
nand U2626 (N_2626,N_672,N_269);
and U2627 (N_2627,N_1798,N_1396);
and U2628 (N_2628,N_1137,N_506);
nand U2629 (N_2629,N_1971,N_1857);
and U2630 (N_2630,N_961,N_2202);
nor U2631 (N_2631,N_68,N_455);
nand U2632 (N_2632,N_2105,N_751);
nor U2633 (N_2633,N_1943,N_1745);
and U2634 (N_2634,N_1166,N_867);
nor U2635 (N_2635,N_545,N_2432);
xor U2636 (N_2636,N_916,N_1450);
xor U2637 (N_2637,N_1026,N_1643);
or U2638 (N_2638,N_1371,N_2441);
or U2639 (N_2639,N_1692,N_1661);
and U2640 (N_2640,N_97,N_2445);
xnor U2641 (N_2641,N_794,N_1245);
nand U2642 (N_2642,N_273,N_1449);
or U2643 (N_2643,N_848,N_619);
nor U2644 (N_2644,N_2234,N_793);
and U2645 (N_2645,N_1200,N_441);
nand U2646 (N_2646,N_1825,N_1700);
or U2647 (N_2647,N_195,N_1078);
xnor U2648 (N_2648,N_287,N_1432);
nand U2649 (N_2649,N_155,N_2122);
or U2650 (N_2650,N_705,N_1868);
or U2651 (N_2651,N_1187,N_2091);
xnor U2652 (N_2652,N_2165,N_2177);
or U2653 (N_2653,N_1921,N_146);
nor U2654 (N_2654,N_15,N_138);
nand U2655 (N_2655,N_1053,N_873);
xnor U2656 (N_2656,N_1882,N_969);
and U2657 (N_2657,N_400,N_504);
nand U2658 (N_2658,N_2270,N_99);
nor U2659 (N_2659,N_1309,N_2075);
nand U2660 (N_2660,N_1107,N_394);
nand U2661 (N_2661,N_952,N_556);
or U2662 (N_2662,N_1377,N_2131);
nand U2663 (N_2663,N_836,N_1967);
and U2664 (N_2664,N_839,N_1151);
or U2665 (N_2665,N_1268,N_477);
nor U2666 (N_2666,N_5,N_920);
nand U2667 (N_2667,N_1520,N_849);
nor U2668 (N_2668,N_1585,N_754);
and U2669 (N_2669,N_148,N_1277);
nand U2670 (N_2670,N_2337,N_2093);
nand U2671 (N_2671,N_1952,N_1655);
xnor U2672 (N_2672,N_987,N_2340);
and U2673 (N_2673,N_1793,N_1602);
or U2674 (N_2674,N_442,N_2101);
or U2675 (N_2675,N_2036,N_1954);
and U2676 (N_2676,N_826,N_1790);
nand U2677 (N_2677,N_965,N_1887);
nor U2678 (N_2678,N_87,N_1129);
and U2679 (N_2679,N_1273,N_2206);
nand U2680 (N_2680,N_1586,N_354);
nor U2681 (N_2681,N_59,N_512);
nand U2682 (N_2682,N_771,N_177);
nand U2683 (N_2683,N_45,N_1912);
and U2684 (N_2684,N_445,N_1120);
nand U2685 (N_2685,N_140,N_1958);
or U2686 (N_2686,N_1826,N_2452);
and U2687 (N_2687,N_1392,N_310);
nor U2688 (N_2688,N_2319,N_1080);
nor U2689 (N_2689,N_2189,N_1250);
nor U2690 (N_2690,N_1156,N_1111);
and U2691 (N_2691,N_1267,N_383);
xor U2692 (N_2692,N_735,N_1240);
and U2693 (N_2693,N_648,N_1527);
nand U2694 (N_2694,N_696,N_1056);
or U2695 (N_2695,N_1850,N_1412);
nor U2696 (N_2696,N_483,N_2241);
xnor U2697 (N_2697,N_1968,N_1598);
nand U2698 (N_2698,N_1861,N_421);
and U2699 (N_2699,N_438,N_1257);
and U2700 (N_2700,N_1583,N_2116);
nand U2701 (N_2701,N_2423,N_2088);
nand U2702 (N_2702,N_65,N_2242);
or U2703 (N_2703,N_1175,N_40);
or U2704 (N_2704,N_1718,N_31);
xnor U2705 (N_2705,N_292,N_1017);
and U2706 (N_2706,N_994,N_2026);
or U2707 (N_2707,N_154,N_1994);
and U2708 (N_2708,N_1754,N_568);
and U2709 (N_2709,N_1006,N_2339);
nand U2710 (N_2710,N_900,N_1369);
nor U2711 (N_2711,N_2057,N_1009);
xor U2712 (N_2712,N_1126,N_1292);
and U2713 (N_2713,N_1409,N_2208);
nand U2714 (N_2714,N_2048,N_1761);
nand U2715 (N_2715,N_426,N_403);
and U2716 (N_2716,N_1573,N_1030);
or U2717 (N_2717,N_185,N_2050);
nor U2718 (N_2718,N_588,N_577);
xnor U2719 (N_2719,N_1561,N_270);
nand U2720 (N_2720,N_1883,N_659);
or U2721 (N_2721,N_104,N_762);
and U2722 (N_2722,N_698,N_655);
nor U2723 (N_2723,N_466,N_962);
nor U2724 (N_2724,N_2195,N_758);
and U2725 (N_2725,N_2273,N_2271);
nand U2726 (N_2726,N_1990,N_73);
and U2727 (N_2727,N_1033,N_2469);
or U2728 (N_2728,N_2176,N_2331);
nand U2729 (N_2729,N_1372,N_1512);
and U2730 (N_2730,N_768,N_1041);
nor U2731 (N_2731,N_567,N_404);
or U2732 (N_2732,N_626,N_1526);
nor U2733 (N_2733,N_1569,N_1539);
or U2734 (N_2734,N_2115,N_1496);
and U2735 (N_2735,N_1847,N_1840);
or U2736 (N_2736,N_2170,N_1416);
nand U2737 (N_2737,N_1841,N_1983);
nor U2738 (N_2738,N_630,N_1976);
nand U2739 (N_2739,N_1015,N_800);
nor U2740 (N_2740,N_607,N_1310);
or U2741 (N_2741,N_543,N_131);
nand U2742 (N_2742,N_921,N_1417);
or U2743 (N_2743,N_1834,N_2295);
or U2744 (N_2744,N_737,N_2418);
xnor U2745 (N_2745,N_1091,N_1905);
or U2746 (N_2746,N_472,N_1969);
and U2747 (N_2747,N_2417,N_452);
and U2748 (N_2748,N_1631,N_2025);
or U2749 (N_2749,N_2492,N_2133);
or U2750 (N_2750,N_985,N_2462);
and U2751 (N_2751,N_850,N_726);
and U2752 (N_2752,N_1867,N_368);
or U2753 (N_2753,N_1686,N_1186);
nor U2754 (N_2754,N_107,N_1319);
and U2755 (N_2755,N_1125,N_1960);
nor U2756 (N_2756,N_2196,N_2020);
xor U2757 (N_2757,N_1486,N_773);
nand U2758 (N_2758,N_899,N_1494);
nand U2759 (N_2759,N_2327,N_2415);
nand U2760 (N_2760,N_989,N_578);
and U2761 (N_2761,N_2309,N_509);
and U2762 (N_2762,N_1707,N_1558);
or U2763 (N_2763,N_2479,N_2045);
or U2764 (N_2764,N_1165,N_1390);
xor U2765 (N_2765,N_1182,N_275);
nand U2766 (N_2766,N_2354,N_1690);
nor U2767 (N_2767,N_817,N_2422);
nor U2768 (N_2768,N_523,N_622);
and U2769 (N_2769,N_1713,N_159);
nand U2770 (N_2770,N_349,N_996);
and U2771 (N_2771,N_313,N_1163);
or U2772 (N_2772,N_462,N_1947);
nand U2773 (N_2773,N_247,N_1815);
and U2774 (N_2774,N_2307,N_1032);
nand U2775 (N_2775,N_289,N_2343);
and U2776 (N_2776,N_1581,N_1940);
and U2777 (N_2777,N_2360,N_602);
and U2778 (N_2778,N_927,N_33);
nand U2779 (N_2779,N_98,N_1298);
or U2780 (N_2780,N_1510,N_576);
nand U2781 (N_2781,N_1755,N_1075);
nand U2782 (N_2782,N_878,N_1515);
nor U2783 (N_2783,N_41,N_1158);
nand U2784 (N_2784,N_2265,N_232);
or U2785 (N_2785,N_0,N_2041);
nor U2786 (N_2786,N_67,N_2076);
nand U2787 (N_2787,N_1594,N_127);
nor U2788 (N_2788,N_1742,N_456);
or U2789 (N_2789,N_1639,N_2142);
nand U2790 (N_2790,N_589,N_1169);
or U2791 (N_2791,N_1523,N_1410);
or U2792 (N_2792,N_1963,N_1209);
nand U2793 (N_2793,N_2067,N_1460);
nand U2794 (N_2794,N_662,N_250);
or U2795 (N_2795,N_660,N_2277);
nand U2796 (N_2796,N_2014,N_10);
xnor U2797 (N_2797,N_295,N_606);
and U2798 (N_2798,N_1048,N_1838);
xor U2799 (N_2799,N_937,N_2128);
nand U2800 (N_2800,N_2372,N_1462);
nand U2801 (N_2801,N_1061,N_1386);
nand U2802 (N_2802,N_2156,N_2288);
and U2803 (N_2803,N_284,N_1103);
nand U2804 (N_2804,N_1630,N_388);
xor U2805 (N_2805,N_66,N_1442);
nand U2806 (N_2806,N_2480,N_2436);
and U2807 (N_2807,N_1955,N_1870);
and U2808 (N_2808,N_396,N_1856);
nor U2809 (N_2809,N_2437,N_2444);
nor U2810 (N_2810,N_555,N_51);
or U2811 (N_2811,N_1489,N_479);
nor U2812 (N_2812,N_731,N_1433);
or U2813 (N_2813,N_586,N_1067);
and U2814 (N_2814,N_1414,N_1064);
and U2815 (N_2815,N_134,N_593);
xnor U2816 (N_2816,N_833,N_406);
and U2817 (N_2817,N_53,N_12);
nor U2818 (N_2818,N_1384,N_1685);
or U2819 (N_2819,N_1063,N_429);
nand U2820 (N_2820,N_1247,N_1524);
nor U2821 (N_2821,N_716,N_1938);
nor U2822 (N_2822,N_1234,N_956);
xnor U2823 (N_2823,N_355,N_1226);
and U2824 (N_2824,N_2096,N_877);
xnor U2825 (N_2825,N_803,N_915);
or U2826 (N_2826,N_901,N_1819);
xor U2827 (N_2827,N_2280,N_95);
nand U2828 (N_2828,N_2450,N_1229);
and U2829 (N_2829,N_1730,N_1457);
or U2830 (N_2830,N_366,N_1642);
nor U2831 (N_2831,N_537,N_1459);
nor U2832 (N_2832,N_1476,N_64);
and U2833 (N_2833,N_16,N_1760);
and U2834 (N_2834,N_640,N_2268);
and U2835 (N_2835,N_1317,N_204);
and U2836 (N_2836,N_470,N_481);
nand U2837 (N_2837,N_529,N_1766);
nor U2838 (N_2838,N_1154,N_1572);
nor U2839 (N_2839,N_843,N_1222);
or U2840 (N_2840,N_1231,N_255);
and U2841 (N_2841,N_2090,N_1663);
nor U2842 (N_2842,N_1500,N_1935);
nor U2843 (N_2843,N_2037,N_1816);
and U2844 (N_2844,N_1957,N_891);
nand U2845 (N_2845,N_1366,N_853);
nand U2846 (N_2846,N_2120,N_22);
nand U2847 (N_2847,N_1949,N_1809);
and U2848 (N_2848,N_747,N_88);
nor U2849 (N_2849,N_787,N_83);
nand U2850 (N_2850,N_1346,N_2464);
nand U2851 (N_2851,N_1328,N_2204);
xor U2852 (N_2852,N_367,N_1058);
xnor U2853 (N_2853,N_720,N_714);
or U2854 (N_2854,N_1759,N_1708);
or U2855 (N_2855,N_2429,N_1985);
nand U2856 (N_2856,N_1618,N_1808);
nor U2857 (N_2857,N_276,N_559);
nor U2858 (N_2858,N_260,N_972);
or U2859 (N_2859,N_2017,N_1688);
or U2860 (N_2860,N_945,N_261);
nor U2861 (N_2861,N_2394,N_611);
or U2862 (N_2862,N_173,N_2164);
or U2863 (N_2863,N_1150,N_933);
nor U2864 (N_2864,N_955,N_2362);
nand U2865 (N_2865,N_1052,N_874);
or U2866 (N_2866,N_225,N_733);
and U2867 (N_2867,N_1914,N_1559);
or U2868 (N_2868,N_496,N_2098);
nand U2869 (N_2869,N_2365,N_116);
nand U2870 (N_2870,N_582,N_919);
and U2871 (N_2871,N_1271,N_750);
and U2872 (N_2872,N_391,N_2117);
nand U2873 (N_2873,N_62,N_1299);
nand U2874 (N_2874,N_924,N_333);
nand U2875 (N_2875,N_1477,N_647);
or U2876 (N_2876,N_2493,N_2300);
nor U2877 (N_2877,N_1096,N_81);
and U2878 (N_2878,N_2284,N_1915);
nand U2879 (N_2879,N_34,N_1474);
nor U2880 (N_2880,N_1482,N_1852);
nor U2881 (N_2881,N_738,N_1835);
xor U2882 (N_2882,N_1365,N_1719);
and U2883 (N_2883,N_38,N_175);
or U2884 (N_2884,N_609,N_2405);
and U2885 (N_2885,N_1903,N_2063);
and U2886 (N_2886,N_2312,N_1109);
nand U2887 (N_2887,N_306,N_591);
nand U2888 (N_2888,N_2232,N_1475);
and U2889 (N_2889,N_695,N_82);
and U2890 (N_2890,N_813,N_889);
or U2891 (N_2891,N_601,N_1363);
xnor U2892 (N_2892,N_816,N_1998);
nor U2893 (N_2893,N_2495,N_291);
nand U2894 (N_2894,N_558,N_1361);
nor U2895 (N_2895,N_753,N_928);
nor U2896 (N_2896,N_290,N_1612);
nand U2897 (N_2897,N_769,N_286);
and U2898 (N_2898,N_415,N_658);
nand U2899 (N_2899,N_904,N_1590);
nor U2900 (N_2900,N_1525,N_1781);
and U2901 (N_2901,N_564,N_1394);
nand U2902 (N_2902,N_1606,N_1528);
or U2903 (N_2903,N_1398,N_2457);
xor U2904 (N_2904,N_827,N_1827);
and U2905 (N_2905,N_1004,N_36);
nor U2906 (N_2906,N_991,N_360);
and U2907 (N_2907,N_74,N_594);
nor U2908 (N_2908,N_1786,N_2488);
and U2909 (N_2909,N_599,N_1227);
or U2910 (N_2910,N_1314,N_1018);
nor U2911 (N_2911,N_2243,N_690);
and U2912 (N_2912,N_327,N_515);
nor U2913 (N_2913,N_180,N_2293);
and U2914 (N_2914,N_603,N_1731);
or U2915 (N_2915,N_2127,N_2201);
or U2916 (N_2916,N_220,N_1633);
or U2917 (N_2917,N_2171,N_585);
nand U2918 (N_2918,N_495,N_1451);
nor U2919 (N_2919,N_1828,N_114);
nand U2920 (N_2920,N_1095,N_2150);
nor U2921 (N_2921,N_1746,N_147);
and U2922 (N_2922,N_142,N_1213);
and U2923 (N_2923,N_1201,N_1944);
nand U2924 (N_2924,N_2065,N_777);
nor U2925 (N_2925,N_801,N_2274);
and U2926 (N_2926,N_728,N_1418);
and U2927 (N_2927,N_1436,N_665);
nand U2928 (N_2928,N_1720,N_1927);
and U2929 (N_2929,N_1024,N_2477);
or U2930 (N_2930,N_2182,N_2078);
xor U2931 (N_2931,N_982,N_2113);
xor U2932 (N_2932,N_121,N_1353);
nor U2933 (N_2933,N_1920,N_2438);
and U2934 (N_2934,N_992,N_520);
nor U2935 (N_2935,N_797,N_1456);
and U2936 (N_2936,N_256,N_447);
nor U2937 (N_2937,N_1822,N_1047);
nand U2938 (N_2938,N_984,N_228);
nand U2939 (N_2939,N_791,N_120);
nor U2940 (N_2940,N_399,N_1888);
xor U2941 (N_2941,N_1677,N_1934);
nand U2942 (N_2942,N_436,N_1463);
xor U2943 (N_2943,N_633,N_1836);
or U2944 (N_2944,N_932,N_494);
nand U2945 (N_2945,N_666,N_866);
or U2946 (N_2946,N_770,N_979);
and U2947 (N_2947,N_1144,N_1767);
and U2948 (N_2948,N_882,N_1783);
xor U2949 (N_2949,N_1665,N_1206);
or U2950 (N_2950,N_1104,N_1093);
nor U2951 (N_2951,N_1925,N_2148);
nor U2952 (N_2952,N_2338,N_2499);
nor U2953 (N_2953,N_1195,N_2426);
or U2954 (N_2954,N_2,N_2221);
nand U2955 (N_2955,N_338,N_119);
nand U2956 (N_2956,N_2303,N_1570);
nand U2957 (N_2957,N_819,N_1776);
nor U2958 (N_2958,N_2427,N_2217);
nor U2959 (N_2959,N_2374,N_689);
nand U2960 (N_2960,N_1866,N_1795);
nor U2961 (N_2961,N_2391,N_499);
and U2962 (N_2962,N_1027,N_1470);
xor U2963 (N_2963,N_70,N_242);
and U2964 (N_2964,N_959,N_1370);
and U2965 (N_2965,N_230,N_628);
and U2966 (N_2966,N_490,N_63);
or U2967 (N_2967,N_123,N_150);
xnor U2968 (N_2968,N_1248,N_2200);
xor U2969 (N_2969,N_1147,N_1728);
nand U2970 (N_2970,N_493,N_654);
nand U2971 (N_2971,N_886,N_1135);
and U2972 (N_2972,N_1694,N_1336);
nor U2973 (N_2973,N_303,N_929);
and U2974 (N_2974,N_1305,N_1654);
xnor U2975 (N_2975,N_322,N_1045);
nand U2976 (N_2976,N_239,N_2344);
nor U2977 (N_2977,N_617,N_691);
nand U2978 (N_2978,N_1695,N_1995);
nand U2979 (N_2979,N_392,N_1114);
xor U2980 (N_2980,N_6,N_2137);
and U2981 (N_2981,N_2132,N_1548);
nand U2982 (N_2982,N_1034,N_1620);
or U2983 (N_2983,N_590,N_527);
xnor U2984 (N_2984,N_1540,N_47);
nand U2985 (N_2985,N_2019,N_1853);
and U2986 (N_2986,N_1161,N_1005);
or U2987 (N_2987,N_297,N_2056);
or U2988 (N_2988,N_1333,N_27);
and U2989 (N_2989,N_1562,N_1875);
and U2990 (N_2990,N_432,N_381);
and U2991 (N_2991,N_153,N_1832);
xnor U2992 (N_2992,N_993,N_106);
or U2993 (N_2993,N_1205,N_293);
xnor U2994 (N_2994,N_2461,N_1007);
nand U2995 (N_2995,N_1427,N_688);
nand U2996 (N_2996,N_823,N_274);
nand U2997 (N_2997,N_1514,N_300);
or U2998 (N_2998,N_2489,N_1975);
nor U2999 (N_2999,N_2373,N_1087);
or U3000 (N_3000,N_1233,N_1542);
nor U3001 (N_3001,N_1863,N_85);
or U3002 (N_3002,N_1948,N_702);
or U3003 (N_3003,N_1901,N_1556);
and U3004 (N_3004,N_736,N_434);
nor U3005 (N_3005,N_393,N_944);
nor U3006 (N_3006,N_1517,N_330);
nor U3007 (N_3007,N_324,N_1072);
nand U3008 (N_3008,N_2336,N_1907);
xor U3009 (N_3009,N_1898,N_1904);
or U3010 (N_3010,N_1070,N_2404);
nand U3011 (N_3011,N_1753,N_1662);
or U3012 (N_3012,N_1097,N_1490);
and U3013 (N_3013,N_1734,N_463);
or U3014 (N_3014,N_1321,N_2203);
and U3015 (N_3015,N_1253,N_491);
nand U3016 (N_3016,N_2267,N_1203);
nor U3017 (N_3017,N_717,N_857);
or U3018 (N_3018,N_669,N_1276);
nor U3019 (N_3019,N_748,N_1036);
and U3020 (N_3020,N_2326,N_2341);
nand U3021 (N_3021,N_2420,N_387);
and U3022 (N_3022,N_1282,N_1183);
nand U3023 (N_3023,N_664,N_583);
nor U3024 (N_3024,N_2281,N_922);
nand U3025 (N_3025,N_1942,N_1604);
nor U3026 (N_3026,N_1683,N_1580);
nand U3027 (N_3027,N_1262,N_1008);
xnor U3028 (N_3028,N_369,N_755);
nand U3029 (N_3029,N_2074,N_1444);
nor U3030 (N_3030,N_2024,N_1928);
nor U3031 (N_3031,N_1999,N_1763);
nand U3032 (N_3032,N_1323,N_90);
or U3033 (N_3033,N_869,N_531);
xor U3034 (N_3034,N_1143,N_492);
nor U3035 (N_3035,N_2181,N_55);
nand U3036 (N_3036,N_1593,N_1173);
or U3037 (N_3037,N_1518,N_1303);
nand U3038 (N_3038,N_251,N_1748);
nor U3039 (N_3039,N_1375,N_782);
nor U3040 (N_3040,N_629,N_641);
xnor U3041 (N_3041,N_2385,N_1906);
and U3042 (N_3042,N_686,N_1221);
nor U3043 (N_3043,N_517,N_1071);
nor U3044 (N_3044,N_1917,N_157);
and U3045 (N_3045,N_2000,N_1218);
nor U3046 (N_3046,N_846,N_1031);
nor U3047 (N_3047,N_1911,N_548);
and U3048 (N_3048,N_1382,N_348);
xor U3049 (N_3049,N_2077,N_1830);
or U3050 (N_3050,N_1886,N_1613);
xnor U3051 (N_3051,N_1021,N_1884);
or U3052 (N_3052,N_1634,N_1356);
and U3053 (N_3053,N_895,N_1453);
nand U3054 (N_3054,N_143,N_1797);
and U3055 (N_3055,N_612,N_347);
xor U3056 (N_3056,N_521,N_1973);
or U3057 (N_3057,N_2357,N_179);
or U3058 (N_3058,N_192,N_911);
and U3059 (N_3059,N_1341,N_1782);
or U3060 (N_3060,N_344,N_375);
nand U3061 (N_3061,N_1491,N_516);
xor U3062 (N_3062,N_1123,N_1387);
and U3063 (N_3063,N_203,N_1119);
xor U3064 (N_3064,N_2275,N_743);
nor U3065 (N_3065,N_914,N_598);
or U3066 (N_3066,N_1258,N_831);
and U3067 (N_3067,N_1022,N_566);
or U3068 (N_3068,N_1575,N_2276);
nor U3069 (N_3069,N_1729,N_910);
nor U3070 (N_3070,N_2446,N_2190);
nand U3071 (N_3071,N_335,N_1821);
and U3072 (N_3072,N_2184,N_1931);
or U3073 (N_3073,N_419,N_637);
nand U3074 (N_3074,N_860,N_262);
and U3075 (N_3075,N_502,N_418);
nor U3076 (N_3076,N_1374,N_1278);
nor U3077 (N_3077,N_2395,N_1263);
and U3078 (N_3078,N_2358,N_1181);
or U3079 (N_3079,N_2085,N_267);
nand U3080 (N_3080,N_2387,N_199);
nand U3081 (N_3081,N_1498,N_2218);
or U3082 (N_3082,N_1956,N_883);
nor U3083 (N_3083,N_1531,N_1002);
nor U3084 (N_3084,N_756,N_2286);
and U3085 (N_3085,N_1640,N_2229);
nand U3086 (N_3086,N_1290,N_592);
xnor U3087 (N_3087,N_1749,N_923);
and U3088 (N_3088,N_2013,N_86);
nor U3089 (N_3089,N_710,N_524);
or U3090 (N_3090,N_1084,N_1621);
nand U3091 (N_3091,N_765,N_380);
nand U3092 (N_3092,N_1784,N_1246);
and U3093 (N_3093,N_1878,N_187);
or U3094 (N_3094,N_1771,N_194);
xnor U3095 (N_3095,N_562,N_1142);
nor U3096 (N_3096,N_906,N_94);
nand U3097 (N_3097,N_1810,N_1077);
xor U3098 (N_3098,N_118,N_217);
nor U3099 (N_3099,N_1582,N_1364);
and U3100 (N_3100,N_378,N_957);
nor U3101 (N_3101,N_2145,N_1959);
and U3102 (N_3102,N_570,N_1725);
nor U3103 (N_3103,N_2130,N_540);
and U3104 (N_3104,N_1829,N_954);
or U3105 (N_3105,N_1487,N_1347);
and U3106 (N_3106,N_1854,N_1428);
or U3107 (N_3107,N_1550,N_2435);
or U3108 (N_3108,N_96,N_2253);
and U3109 (N_3109,N_1220,N_656);
or U3110 (N_3110,N_1115,N_1224);
or U3111 (N_3111,N_1407,N_1059);
and U3112 (N_3112,N_2185,N_1717);
and U3113 (N_3113,N_25,N_1946);
or U3114 (N_3114,N_999,N_1122);
and U3115 (N_3115,N_1446,N_197);
or U3116 (N_3116,N_1578,N_448);
xor U3117 (N_3117,N_2240,N_2214);
nor U3118 (N_3118,N_182,N_474);
or U3119 (N_3119,N_2470,N_623);
or U3120 (N_3120,N_1441,N_774);
or U3121 (N_3121,N_783,N_2313);
or U3122 (N_3122,N_1902,N_636);
nand U3123 (N_3123,N_779,N_2060);
or U3124 (N_3124,N_1073,N_608);
and U3125 (N_3125,N_807,N_2416);
and U3126 (N_3126,N_580,N_363);
nand U3127 (N_3127,N_1989,N_1153);
and U3128 (N_3128,N_2003,N_998);
nor U3129 (N_3129,N_35,N_2306);
nor U3130 (N_3130,N_265,N_761);
nor U3131 (N_3131,N_571,N_1176);
xnor U3132 (N_3132,N_2138,N_2175);
nand U3133 (N_3133,N_328,N_822);
or U3134 (N_3134,N_2325,N_1802);
or U3135 (N_3135,N_1926,N_587);
nor U3136 (N_3136,N_1454,N_2272);
nand U3137 (N_3137,N_1029,N_317);
nand U3138 (N_3138,N_2099,N_1697);
or U3139 (N_3139,N_2398,N_2459);
nand U3140 (N_3140,N_353,N_1443);
nor U3141 (N_3141,N_405,N_1085);
or U3142 (N_3142,N_539,N_2486);
or U3143 (N_3143,N_1843,N_20);
nand U3144 (N_3144,N_1132,N_1984);
nor U3145 (N_3145,N_409,N_2369);
or U3146 (N_3146,N_1001,N_1987);
and U3147 (N_3147,N_2301,N_1974);
nand U3148 (N_3148,N_1596,N_263);
and U3149 (N_3149,N_1060,N_2001);
xnor U3150 (N_3150,N_2371,N_763);
xnor U3151 (N_3151,N_511,N_1614);
and U3152 (N_3152,N_2066,N_2051);
and U3153 (N_3153,N_1650,N_2294);
and U3154 (N_3154,N_775,N_1877);
and U3155 (N_3155,N_1422,N_258);
nor U3156 (N_3156,N_2456,N_2278);
and U3157 (N_3157,N_795,N_428);
xnor U3158 (N_3158,N_1189,N_2147);
xnor U3159 (N_3159,N_2261,N_1624);
and U3160 (N_3160,N_1508,N_788);
nand U3161 (N_3161,N_1533,N_643);
nand U3162 (N_3162,N_1230,N_78);
nor U3163 (N_3163,N_2152,N_14);
and U3164 (N_3164,N_156,N_1339);
or U3165 (N_3165,N_2269,N_1773);
nand U3166 (N_3166,N_135,N_2252);
nand U3167 (N_3167,N_1799,N_1664);
nor U3168 (N_3168,N_1335,N_569);
nor U3169 (N_3169,N_1709,N_172);
nor U3170 (N_3170,N_584,N_646);
or U3171 (N_3171,N_809,N_1627);
xnor U3172 (N_3172,N_382,N_615);
and U3173 (N_3173,N_888,N_497);
nand U3174 (N_3174,N_475,N_2377);
nor U3175 (N_3175,N_1171,N_305);
or U3176 (N_3176,N_1358,N_1289);
nand U3177 (N_3177,N_1758,N_917);
nor U3178 (N_3178,N_2149,N_288);
or U3179 (N_3179,N_1814,N_964);
nor U3180 (N_3180,N_2481,N_958);
nor U3181 (N_3181,N_638,N_1452);
xor U3182 (N_3182,N_149,N_1197);
nand U3183 (N_3183,N_1332,N_776);
nor U3184 (N_3184,N_2482,N_1354);
nand U3185 (N_3185,N_222,N_2005);
nand U3186 (N_3186,N_1879,N_1733);
or U3187 (N_3187,N_184,N_1140);
nand U3188 (N_3188,N_395,N_2297);
nor U3189 (N_3189,N_1178,N_1090);
and U3190 (N_3190,N_26,N_898);
or U3191 (N_3191,N_2038,N_767);
and U3192 (N_3192,N_1865,N_926);
or U3193 (N_3193,N_254,N_402);
nor U3194 (N_3194,N_2140,N_2397);
nor U3195 (N_3195,N_2125,N_1116);
nor U3196 (N_3196,N_790,N_1529);
nor U3197 (N_3197,N_974,N_510);
or U3198 (N_3198,N_1676,N_1807);
or U3199 (N_3199,N_2257,N_514);
xnor U3200 (N_3200,N_210,N_1768);
xnor U3201 (N_3201,N_746,N_1551);
xor U3202 (N_3202,N_812,N_77);
xnor U3203 (N_3203,N_1484,N_2384);
xnor U3204 (N_3204,N_1266,N_1281);
nor U3205 (N_3205,N_1180,N_968);
nand U3206 (N_3206,N_294,N_1704);
nand U3207 (N_3207,N_2043,N_1448);
and U3208 (N_3208,N_1874,N_2169);
and U3209 (N_3209,N_236,N_108);
nand U3210 (N_3210,N_1069,N_2069);
nor U3211 (N_3211,N_2350,N_2291);
and U3212 (N_3212,N_1859,N_465);
and U3213 (N_3213,N_431,N_458);
nand U3214 (N_3214,N_682,N_1871);
nand U3215 (N_3215,N_136,N_2064);
or U3216 (N_3216,N_1264,N_875);
or U3217 (N_3217,N_1893,N_2453);
xor U3218 (N_3218,N_1671,N_700);
or U3219 (N_3219,N_1803,N_541);
and U3220 (N_3220,N_1680,N_329);
and U3221 (N_3221,N_913,N_439);
nand U3222 (N_3222,N_1629,N_1343);
or U3223 (N_3223,N_1014,N_2433);
nor U3224 (N_3224,N_1337,N_894);
nand U3225 (N_3225,N_2141,N_1675);
and U3226 (N_3226,N_1003,N_2323);
or U3227 (N_3227,N_2381,N_1812);
nand U3228 (N_3228,N_711,N_2407);
xnor U3229 (N_3229,N_1435,N_575);
and U3230 (N_3230,N_1579,N_605);
nand U3231 (N_3231,N_508,N_811);
nor U3232 (N_3232,N_2044,N_946);
or U3233 (N_3233,N_518,N_433);
or U3234 (N_3234,N_1483,N_1373);
or U3235 (N_3235,N_2409,N_1839);
or U3236 (N_3236,N_2249,N_1738);
or U3237 (N_3237,N_2239,N_1735);
nand U3238 (N_3238,N_2213,N_624);
or U3239 (N_3239,N_218,N_1873);
and U3240 (N_3240,N_1046,N_139);
and U3241 (N_3241,N_868,N_1236);
and U3242 (N_3242,N_2178,N_80);
nand U3243 (N_3243,N_1817,N_1113);
nand U3244 (N_3244,N_1139,N_489);
or U3245 (N_3245,N_708,N_2159);
or U3246 (N_3246,N_1280,N_1916);
nand U3247 (N_3247,N_478,N_2483);
xor U3248 (N_3248,N_2364,N_1623);
nand U3249 (N_3249,N_1455,N_1855);
or U3250 (N_3250,N_2315,N_3);
xnor U3251 (N_3251,N_2352,N_2192);
or U3252 (N_3252,N_1837,N_1493);
nand U3253 (N_3253,N_1403,N_2144);
xor U3254 (N_3254,N_519,N_379);
nand U3255 (N_3255,N_1601,N_257);
nor U3256 (N_3256,N_1294,N_1043);
or U3257 (N_3257,N_334,N_1744);
and U3258 (N_3258,N_2114,N_2109);
and U3259 (N_3259,N_2389,N_634);
nand U3260 (N_3260,N_1479,N_58);
nor U3261 (N_3261,N_326,N_2233);
xnor U3262 (N_3262,N_610,N_532);
and U3263 (N_3263,N_208,N_1405);
nor U3264 (N_3264,N_13,N_2430);
nand U3265 (N_3265,N_1239,N_684);
nor U3266 (N_3266,N_1563,N_1544);
nand U3267 (N_3267,N_1481,N_407);
and U3268 (N_3268,N_2496,N_1638);
nand U3269 (N_3269,N_814,N_1367);
xor U3270 (N_3270,N_1788,N_1811);
or U3271 (N_3271,N_2345,N_1922);
nor U3272 (N_3272,N_1284,N_1401);
nor U3273 (N_3273,N_420,N_1232);
or U3274 (N_3274,N_2174,N_804);
and U3275 (N_3275,N_498,N_1897);
xor U3276 (N_3276,N_1124,N_2283);
nand U3277 (N_3277,N_2168,N_224);
or U3278 (N_3278,N_870,N_1880);
nand U3279 (N_3279,N_487,N_2107);
and U3280 (N_3280,N_1660,N_2317);
xnor U3281 (N_3281,N_981,N_1890);
and U3282 (N_3282,N_600,N_216);
xor U3283 (N_3283,N_1645,N_1413);
nand U3284 (N_3284,N_1794,N_938);
nand U3285 (N_3285,N_1019,N_2363);
and U3286 (N_3286,N_1846,N_28);
nand U3287 (N_3287,N_1610,N_238);
nand U3288 (N_3288,N_596,N_1488);
nor U3289 (N_3289,N_1389,N_2314);
nand U3290 (N_3290,N_1425,N_1212);
xnor U3291 (N_3291,N_1860,N_1108);
nor U3292 (N_3292,N_164,N_2134);
nor U3293 (N_3293,N_786,N_854);
or U3294 (N_3294,N_1751,N_1521);
xnor U3295 (N_3295,N_266,N_2220);
or U3296 (N_3296,N_1391,N_1997);
nor U3297 (N_3297,N_978,N_141);
nor U3298 (N_3298,N_667,N_1308);
or U3299 (N_3299,N_1217,N_1194);
and U3300 (N_3300,N_1252,N_1198);
and U3301 (N_3301,N_2399,N_2191);
nor U3302 (N_3302,N_427,N_1141);
or U3303 (N_3303,N_1465,N_152);
nand U3304 (N_3304,N_451,N_2355);
nand U3305 (N_3305,N_372,N_1789);
xor U3306 (N_3306,N_158,N_2348);
nand U3307 (N_3307,N_1426,N_1283);
nand U3308 (N_3308,N_1682,N_469);
or U3309 (N_3309,N_2126,N_1062);
xnor U3310 (N_3310,N_2298,N_2259);
and U3311 (N_3311,N_2100,N_1167);
nor U3312 (N_3312,N_1805,N_2121);
or U3313 (N_3313,N_865,N_444);
nor U3314 (N_3314,N_2081,N_1670);
or U3315 (N_3315,N_196,N_1932);
nor U3316 (N_3316,N_1307,N_1251);
or U3317 (N_3317,N_30,N_1532);
and U3318 (N_3318,N_46,N_453);
xnor U3319 (N_3319,N_2161,N_845);
nor U3320 (N_3320,N_285,N_2473);
or U3321 (N_3321,N_1237,N_2072);
xnor U3322 (N_3322,N_2092,N_1159);
nor U3323 (N_3323,N_1177,N_2497);
nor U3324 (N_3324,N_824,N_2040);
or U3325 (N_3325,N_1993,N_1568);
nor U3326 (N_3326,N_1536,N_2258);
nor U3327 (N_3327,N_757,N_725);
nand U3328 (N_3328,N_1057,N_2419);
or U3329 (N_3329,N_2228,N_2368);
and U3330 (N_3330,N_2474,N_742);
or U3331 (N_3331,N_1219,N_1223);
nor U3332 (N_3332,N_2421,N_2347);
xnor U3333 (N_3333,N_841,N_471);
nor U3334 (N_3334,N_1698,N_563);
nand U3335 (N_3335,N_29,N_282);
xor U3336 (N_3336,N_54,N_1513);
nor U3337 (N_3337,N_934,N_1778);
or U3338 (N_3338,N_1105,N_253);
or U3339 (N_3339,N_91,N_424);
or U3340 (N_3340,N_745,N_947);
and U3341 (N_3341,N_1691,N_2089);
nor U3342 (N_3342,N_2211,N_2443);
or U3343 (N_3343,N_1193,N_963);
and U3344 (N_3344,N_111,N_1806);
nor U3345 (N_3345,N_1600,N_1208);
xor U3346 (N_3346,N_312,N_109);
nand U3347 (N_3347,N_113,N_741);
nor U3348 (N_3348,N_2223,N_2180);
and U3349 (N_3349,N_2335,N_162);
or U3350 (N_3350,N_1507,N_1693);
or U3351 (N_3351,N_1543,N_1849);
and U3352 (N_3352,N_828,N_341);
nor U3353 (N_3353,N_1546,N_1617);
and U3354 (N_3354,N_245,N_789);
nand U3355 (N_3355,N_2484,N_103);
xnor U3356 (N_3356,N_181,N_677);
or U3357 (N_3357,N_694,N_2227);
nor U3358 (N_3358,N_549,N_1869);
and U3359 (N_3359,N_1199,N_1936);
nand U3360 (N_3360,N_92,N_376);
or U3361 (N_3361,N_198,N_1501);
nand U3362 (N_3362,N_189,N_649);
or U3363 (N_3363,N_2353,N_2454);
and U3364 (N_3364,N_2428,N_1687);
nand U3365 (N_3365,N_1696,N_1986);
and U3366 (N_3366,N_2256,N_967);
nor U3367 (N_3367,N_1678,N_936);
or U3368 (N_3368,N_160,N_268);
nand U3369 (N_3369,N_1352,N_226);
or U3370 (N_3370,N_1553,N_1133);
nor U3371 (N_3371,N_1864,N_1736);
nand U3372 (N_3372,N_1214,N_1651);
nor U3373 (N_3373,N_1591,N_1134);
xnor U3374 (N_3374,N_1715,N_129);
xnor U3375 (N_3375,N_799,N_522);
and U3376 (N_3376,N_1196,N_1599);
or U3377 (N_3377,N_651,N_1972);
xnor U3378 (N_3378,N_1439,N_2022);
nor U3379 (N_3379,N_1440,N_316);
xor U3380 (N_3380,N_446,N_19);
and U3381 (N_3381,N_635,N_681);
or U3382 (N_3382,N_815,N_2402);
and U3383 (N_3383,N_903,N_1592);
or U3384 (N_3384,N_2351,N_1721);
nor U3385 (N_3385,N_976,N_345);
nand U3386 (N_3386,N_2458,N_48);
and U3387 (N_3387,N_1025,N_1584);
nand U3388 (N_3388,N_166,N_780);
nor U3389 (N_3389,N_1011,N_186);
nor U3390 (N_3390,N_2006,N_2254);
and U3391 (N_3391,N_674,N_42);
nor U3392 (N_3392,N_227,N_1635);
nor U3393 (N_3393,N_1669,N_2390);
nand U3394 (N_3394,N_925,N_552);
or U3395 (N_3395,N_1780,N_1285);
nand U3396 (N_3396,N_1054,N_1255);
xnor U3397 (N_3397,N_1541,N_1503);
or U3398 (N_3398,N_2491,N_597);
xor U3399 (N_3399,N_844,N_168);
or U3400 (N_3400,N_259,N_2226);
or U3401 (N_3401,N_234,N_1485);
nor U3402 (N_3402,N_1723,N_983);
and U3403 (N_3403,N_618,N_2111);
nor U3404 (N_3404,N_340,N_1458);
or U3405 (N_3405,N_2009,N_193);
and U3406 (N_3406,N_879,N_2205);
or U3407 (N_3407,N_11,N_1743);
or U3408 (N_3408,N_205,N_1210);
nor U3409 (N_3409,N_450,N_2320);
nor U3410 (N_3410,N_2332,N_1710);
nand U3411 (N_3411,N_2008,N_1311);
nand U3412 (N_3412,N_408,N_117);
and U3413 (N_3413,N_2021,N_1988);
and U3414 (N_3414,N_513,N_1896);
nand U3415 (N_3415,N_2172,N_1378);
xnor U3416 (N_3416,N_410,N_1327);
and U3417 (N_3417,N_2264,N_1885);
xnor U3418 (N_3418,N_60,N_960);
nor U3419 (N_3419,N_2244,N_2311);
and U3420 (N_3420,N_1574,N_79);
nor U3421 (N_3421,N_693,N_1492);
and U3422 (N_3422,N_1334,N_296);
and U3423 (N_3423,N_1402,N_137);
xor U3424 (N_3424,N_673,N_1437);
nor U3425 (N_3425,N_1506,N_1554);
xor U3426 (N_3426,N_1088,N_171);
and U3427 (N_3427,N_52,N_2367);
and U3428 (N_3428,N_115,N_949);
nand U3429 (N_3429,N_1652,N_482);
nand U3430 (N_3430,N_301,N_307);
nand U3431 (N_3431,N_1567,N_2166);
xor U3432 (N_3432,N_1099,N_56);
nand U3433 (N_3433,N_1261,N_727);
and U3434 (N_3434,N_1380,N_351);
xnor U3435 (N_3435,N_1040,N_1118);
xnor U3436 (N_3436,N_1155,N_2034);
nor U3437 (N_3437,N_2027,N_2012);
nor U3438 (N_3438,N_1478,N_1978);
or U3439 (N_3439,N_1970,N_39);
or U3440 (N_3440,N_715,N_1146);
and U3441 (N_3441,N_939,N_830);
or U3442 (N_3442,N_1622,N_1607);
nor U3443 (N_3443,N_342,N_2080);
or U3444 (N_3444,N_2393,N_414);
nand U3445 (N_3445,N_530,N_248);
nor U3446 (N_3446,N_361,N_1010);
or U3447 (N_3447,N_1411,N_1318);
or U3448 (N_3448,N_778,N_93);
nand U3449 (N_3449,N_2052,N_1894);
nand U3450 (N_3450,N_1566,N_2046);
or U3451 (N_3451,N_1800,N_2349);
nor U3452 (N_3452,N_2316,N_1647);
nor U3453 (N_3453,N_525,N_2285);
and U3454 (N_3454,N_443,N_144);
nand U3455 (N_3455,N_1648,N_1424);
and U3456 (N_3456,N_2328,N_832);
and U3457 (N_3457,N_1597,N_1899);
nor U3458 (N_3458,N_2460,N_1385);
xor U3459 (N_3459,N_488,N_2282);
nand U3460 (N_3460,N_650,N_214);
and U3461 (N_3461,N_2255,N_1945);
or U3462 (N_3462,N_2110,N_178);
nand U3463 (N_3463,N_1397,N_1992);
nand U3464 (N_3464,N_425,N_1564);
nand U3465 (N_3465,N_2356,N_174);
nor U3466 (N_3466,N_461,N_1966);
nor U3467 (N_3467,N_389,N_151);
xor U3468 (N_3468,N_1534,N_722);
and U3469 (N_3469,N_1732,N_798);
or U3470 (N_3470,N_215,N_2028);
xnor U3471 (N_3471,N_1722,N_2408);
xor U3472 (N_3472,N_1471,N_2246);
nand U3473 (N_3473,N_1705,N_169);
xor U3474 (N_3474,N_422,N_2366);
nor U3475 (N_3475,N_69,N_279);
nor U3476 (N_3476,N_2414,N_699);
or U3477 (N_3477,N_852,N_616);
or U3478 (N_3478,N_299,N_892);
xor U3479 (N_3479,N_2448,N_321);
and U3480 (N_3480,N_1668,N_808);
and U3481 (N_3481,N_2290,N_2187);
and U3482 (N_3482,N_124,N_1331);
xor U3483 (N_3483,N_1549,N_1254);
nand U3484 (N_3484,N_1641,N_897);
nor U3485 (N_3485,N_759,N_2260);
and U3486 (N_3486,N_1138,N_2154);
nand U3487 (N_3487,N_1933,N_1172);
or U3488 (N_3488,N_2173,N_413);
and U3489 (N_3489,N_851,N_2030);
nor U3490 (N_3490,N_435,N_1737);
nor U3491 (N_3491,N_357,N_332);
nand U3492 (N_3492,N_1689,N_1089);
nor U3493 (N_3493,N_1094,N_377);
xnor U3494 (N_3494,N_2245,N_76);
and U3495 (N_3495,N_1270,N_1068);
and U3496 (N_3496,N_359,N_884);
or U3497 (N_3497,N_1716,N_988);
xor U3498 (N_3498,N_188,N_246);
nor U3499 (N_3499,N_1605,N_1362);
and U3500 (N_3500,N_1900,N_829);
or U3501 (N_3501,N_1012,N_430);
xor U3502 (N_3502,N_876,N_309);
or U3503 (N_3503,N_1243,N_1842);
nand U3504 (N_3504,N_692,N_1079);
nor U3505 (N_3505,N_1779,N_2119);
nand U3506 (N_3506,N_802,N_440);
and U3507 (N_3507,N_620,N_1306);
or U3508 (N_3508,N_503,N_2318);
or U3509 (N_3509,N_1962,N_1164);
nor U3510 (N_3510,N_1545,N_930);
nor U3511 (N_3511,N_533,N_2380);
or U3512 (N_3512,N_190,N_1724);
nor U3513 (N_3513,N_1312,N_1184);
and U3514 (N_3514,N_1297,N_713);
and U3515 (N_3515,N_2330,N_2210);
or U3516 (N_3516,N_840,N_2475);
and U3517 (N_3517,N_454,N_1609);
nor U3518 (N_3518,N_2010,N_2073);
or U3519 (N_3519,N_2023,N_1982);
nand U3520 (N_3520,N_2455,N_1611);
nor U3521 (N_3521,N_2035,N_1274);
and U3522 (N_3522,N_1324,N_1438);
and U3523 (N_3523,N_734,N_1739);
and U3524 (N_3524,N_990,N_264);
nand U3525 (N_3525,N_1702,N_560);
nand U3526 (N_3526,N_730,N_1149);
nand U3527 (N_3527,N_1065,N_283);
nor U3528 (N_3528,N_1892,N_1557);
nor U3529 (N_3529,N_2094,N_318);
nand U3530 (N_3530,N_1086,N_1923);
nor U3531 (N_3531,N_1066,N_464);
and U3532 (N_3532,N_1774,N_1659);
or U3533 (N_3533,N_298,N_1646);
and U3534 (N_3534,N_1565,N_1188);
nor U3535 (N_3535,N_1148,N_1818);
nand U3536 (N_3536,N_1616,N_858);
nand U3537 (N_3537,N_1351,N_2434);
or U3538 (N_3538,N_339,N_8);
nand U3539 (N_3539,N_350,N_314);
or U3540 (N_3540,N_1537,N_1406);
nor U3541 (N_3541,N_1357,N_821);
nor U3542 (N_3542,N_2059,N_1013);
and U3543 (N_3543,N_772,N_2160);
nor U3544 (N_3544,N_2163,N_970);
and U3545 (N_3545,N_561,N_621);
nor U3546 (N_3546,N_241,N_2198);
nand U3547 (N_3547,N_2296,N_1360);
or U3548 (N_3548,N_980,N_1316);
xnor U3549 (N_3549,N_2299,N_2083);
nand U3550 (N_3550,N_1329,N_2216);
or U3551 (N_3551,N_280,N_457);
nor U3552 (N_3552,N_337,N_995);
xor U3553 (N_3553,N_110,N_1296);
and U3554 (N_3554,N_810,N_1764);
nor U3555 (N_3555,N_1632,N_362);
xnor U3556 (N_3556,N_2292,N_1260);
nor U3557 (N_3557,N_423,N_2238);
nand U3558 (N_3558,N_887,N_75);
and U3559 (N_3559,N_2487,N_2490);
xor U3560 (N_3560,N_2102,N_2359);
and U3561 (N_3561,N_1102,N_701);
nor U3562 (N_3562,N_905,N_2396);
nor U3563 (N_3563,N_2250,N_724);
nand U3564 (N_3564,N_2209,N_44);
or U3565 (N_3565,N_1844,N_1468);
nand U3566 (N_3566,N_931,N_1981);
xor U3567 (N_3567,N_1497,N_2413);
nor U3568 (N_3568,N_1657,N_212);
or U3569 (N_3569,N_2015,N_706);
nor U3570 (N_3570,N_1530,N_1714);
xor U3571 (N_3571,N_2449,N_4);
nor U3572 (N_3572,N_2153,N_943);
nand U3573 (N_3573,N_1301,N_1215);
nand U3574 (N_3574,N_825,N_240);
and U3575 (N_3575,N_536,N_1851);
nand U3576 (N_3576,N_1429,N_1037);
and U3577 (N_3577,N_2386,N_2054);
and U3578 (N_3578,N_861,N_1395);
nand U3579 (N_3579,N_781,N_871);
nor U3580 (N_3580,N_2136,N_229);
nor U3581 (N_3581,N_2310,N_2425);
and U3582 (N_3582,N_476,N_2047);
or U3583 (N_3583,N_209,N_1765);
nor U3584 (N_3584,N_1876,N_1207);
and U3585 (N_3585,N_1615,N_1769);
or U3586 (N_3586,N_1315,N_397);
and U3587 (N_3587,N_1295,N_505);
and U3588 (N_3588,N_918,N_796);
and U3589 (N_3589,N_237,N_2302);
xor U3590 (N_3590,N_7,N_343);
xor U3591 (N_3591,N_864,N_2370);
or U3592 (N_3592,N_165,N_1872);
and U3593 (N_3593,N_1881,N_1918);
or U3594 (N_3594,N_221,N_356);
nand U3595 (N_3595,N_1279,N_1701);
and U3596 (N_3596,N_480,N_657);
nor U3597 (N_3597,N_642,N_953);
nor U3598 (N_3598,N_1937,N_2440);
and U3599 (N_3599,N_1991,N_72);
nand U3600 (N_3600,N_1472,N_557);
and U3601 (N_3601,N_719,N_614);
nor U3602 (N_3602,N_507,N_1291);
nand U3603 (N_3603,N_1547,N_2011);
xnor U3604 (N_3604,N_632,N_2466);
nand U3605 (N_3605,N_1577,N_2465);
nor U3606 (N_3606,N_740,N_535);
nand U3607 (N_3607,N_704,N_908);
nand U3608 (N_3608,N_411,N_2158);
and U3609 (N_3609,N_1225,N_1667);
and U3610 (N_3610,N_473,N_2162);
nand U3611 (N_3611,N_1112,N_1269);
or U3612 (N_3612,N_2308,N_1170);
or U3613 (N_3613,N_707,N_1431);
and U3614 (N_3614,N_2146,N_50);
and U3615 (N_3615,N_2097,N_856);
and U3616 (N_3616,N_2431,N_365);
xnor U3617 (N_3617,N_538,N_550);
and U3618 (N_3618,N_880,N_244);
and U3619 (N_3619,N_2375,N_2157);
or U3620 (N_3620,N_792,N_2333);
xor U3621 (N_3621,N_2324,N_1216);
and U3622 (N_3622,N_1681,N_553);
nand U3623 (N_3623,N_644,N_2058);
nand U3624 (N_3624,N_1750,N_2478);
nor U3625 (N_3625,N_1595,N_2071);
or U3626 (N_3626,N_1712,N_1467);
xnor U3627 (N_3627,N_1016,N_2498);
nand U3628 (N_3628,N_1464,N_2103);
nand U3629 (N_3629,N_1192,N_2018);
or U3630 (N_3630,N_1051,N_207);
and U3631 (N_3631,N_1511,N_806);
xnor U3632 (N_3632,N_1342,N_835);
and U3633 (N_3633,N_2004,N_721);
or U3634 (N_3634,N_1772,N_24);
nor U3635 (N_3635,N_2231,N_2262);
nand U3636 (N_3636,N_1777,N_1538);
and U3637 (N_3637,N_862,N_1740);
nor U3638 (N_3638,N_1466,N_1762);
or U3639 (N_3639,N_1202,N_912);
nand U3640 (N_3640,N_1603,N_573);
xnor U3641 (N_3641,N_1320,N_2411);
nand U3642 (N_3642,N_2139,N_554);
nor U3643 (N_3643,N_2230,N_437);
nand U3644 (N_3644,N_752,N_941);
and U3645 (N_3645,N_671,N_1833);
and U3646 (N_3646,N_2070,N_2263);
nor U3647 (N_3647,N_1801,N_1628);
nand U3648 (N_3648,N_1831,N_1423);
nor U3649 (N_3649,N_1235,N_1447);
and U3650 (N_3650,N_384,N_2406);
nor U3651 (N_3651,N_176,N_125);
nand U3652 (N_3652,N_71,N_805);
nor U3653 (N_3653,N_1388,N_1325);
xor U3654 (N_3654,N_1535,N_319);
and U3655 (N_3655,N_1293,N_948);
and U3656 (N_3656,N_243,N_1110);
nand U3657 (N_3657,N_1757,N_1649);
or U3658 (N_3658,N_1434,N_1504);
nor U3659 (N_3659,N_364,N_1658);
and U3660 (N_3660,N_1160,N_2361);
xnor U3661 (N_3661,N_1502,N_2235);
and U3662 (N_3662,N_1049,N_1092);
xor U3663 (N_3663,N_1000,N_1891);
or U3664 (N_3664,N_1699,N_1355);
or U3665 (N_3665,N_639,N_1348);
and U3666 (N_3666,N_1300,N_133);
or U3667 (N_3667,N_459,N_2112);
or U3668 (N_3668,N_1345,N_2439);
nor U3669 (N_3669,N_1509,N_678);
or U3670 (N_3670,N_191,N_84);
nand U3671 (N_3671,N_2329,N_130);
nand U3672 (N_3672,N_2471,N_940);
nor U3673 (N_3673,N_1929,N_1775);
nor U3674 (N_3674,N_896,N_1858);
nor U3675 (N_3675,N_2376,N_1098);
and U3676 (N_3676,N_2062,N_1131);
or U3677 (N_3677,N_1499,N_1930);
nand U3678 (N_3678,N_2382,N_645);
nor U3679 (N_3679,N_872,N_412);
nor U3680 (N_3680,N_61,N_2055);
or U3681 (N_3681,N_2179,N_485);
nor U3682 (N_3682,N_2494,N_935);
and U3683 (N_3683,N_1980,N_1644);
xor U3684 (N_3684,N_1951,N_1824);
or U3685 (N_3685,N_1368,N_2124);
and U3686 (N_3686,N_484,N_1804);
nor U3687 (N_3687,N_683,N_1399);
or U3688 (N_3688,N_837,N_1461);
nor U3689 (N_3689,N_1242,N_2207);
and U3690 (N_3690,N_977,N_1074);
nor U3691 (N_3691,N_1039,N_859);
nand U3692 (N_3692,N_847,N_1792);
xnor U3693 (N_3693,N_1924,N_2236);
nand U3694 (N_3694,N_1711,N_1393);
nor U3695 (N_3695,N_1706,N_687);
xor U3696 (N_3696,N_2248,N_1672);
nand U3697 (N_3697,N_211,N_1756);
xor U3698 (N_3698,N_1679,N_272);
nor U3699 (N_3699,N_1185,N_579);
nor U3700 (N_3700,N_17,N_1020);
nor U3701 (N_3701,N_2087,N_1445);
and U3702 (N_3702,N_1,N_2084);
nand U3703 (N_3703,N_1211,N_1950);
and U3704 (N_3704,N_973,N_2108);
nand U3705 (N_3705,N_1383,N_417);
and U3706 (N_3706,N_385,N_132);
nor U3707 (N_3707,N_685,N_206);
and U3708 (N_3708,N_308,N_1555);
or U3709 (N_3709,N_1560,N_2401);
nor U3710 (N_3710,N_2029,N_1516);
nand U3711 (N_3711,N_1408,N_1674);
or U3712 (N_3712,N_668,N_486);
nand U3713 (N_3713,N_468,N_278);
nor U3714 (N_3714,N_1376,N_373);
nor U3715 (N_3715,N_1106,N_200);
nor U3716 (N_3716,N_2247,N_2031);
or U3717 (N_3717,N_9,N_1653);
and U3718 (N_3718,N_1101,N_1228);
or U3719 (N_3719,N_2346,N_902);
or U3720 (N_3720,N_1082,N_2068);
and U3721 (N_3721,N_2410,N_32);
and U3722 (N_3722,N_1042,N_818);
and U3723 (N_3723,N_2199,N_703);
and U3724 (N_3724,N_2251,N_2342);
nor U3725 (N_3725,N_57,N_2451);
nand U3726 (N_3726,N_1168,N_604);
xor U3727 (N_3727,N_1996,N_163);
nand U3728 (N_3728,N_1961,N_2082);
and U3729 (N_3729,N_1265,N_2321);
nor U3730 (N_3730,N_302,N_346);
xnor U3731 (N_3731,N_881,N_101);
nand U3732 (N_3732,N_2188,N_2378);
and U3733 (N_3733,N_723,N_2224);
nor U3734 (N_3734,N_2039,N_950);
or U3735 (N_3735,N_676,N_1204);
xor U3736 (N_3736,N_1128,N_122);
xnor U3737 (N_3737,N_252,N_709);
and U3738 (N_3738,N_627,N_2007);
and U3739 (N_3739,N_764,N_1791);
nor U3740 (N_3740,N_2053,N_1379);
nor U3741 (N_3741,N_1727,N_1028);
xor U3742 (N_3742,N_971,N_1313);
xor U3743 (N_3743,N_1130,N_2106);
xnor U3744 (N_3744,N_2289,N_401);
nand U3745 (N_3745,N_1420,N_1505);
nor U3746 (N_3746,N_161,N_2215);
or U3747 (N_3747,N_2392,N_323);
and U3748 (N_3748,N_1179,N_170);
nand U3749 (N_3749,N_1162,N_1796);
nand U3750 (N_3750,N_935,N_2223);
nand U3751 (N_3751,N_1796,N_1100);
nor U3752 (N_3752,N_1360,N_1517);
nand U3753 (N_3753,N_469,N_1381);
nand U3754 (N_3754,N_245,N_2150);
or U3755 (N_3755,N_677,N_1825);
nand U3756 (N_3756,N_1567,N_1990);
nand U3757 (N_3757,N_1015,N_2378);
or U3758 (N_3758,N_757,N_142);
or U3759 (N_3759,N_918,N_2435);
or U3760 (N_3760,N_1109,N_2302);
and U3761 (N_3761,N_332,N_880);
or U3762 (N_3762,N_2432,N_2056);
xnor U3763 (N_3763,N_475,N_263);
nor U3764 (N_3764,N_229,N_790);
xnor U3765 (N_3765,N_1867,N_228);
xnor U3766 (N_3766,N_2,N_1089);
nand U3767 (N_3767,N_335,N_2011);
and U3768 (N_3768,N_1028,N_2441);
nor U3769 (N_3769,N_1914,N_1680);
and U3770 (N_3770,N_1686,N_657);
nor U3771 (N_3771,N_1171,N_1593);
nor U3772 (N_3772,N_1218,N_1221);
nor U3773 (N_3773,N_475,N_99);
and U3774 (N_3774,N_162,N_1497);
nand U3775 (N_3775,N_1676,N_796);
and U3776 (N_3776,N_1422,N_286);
or U3777 (N_3777,N_1824,N_255);
nand U3778 (N_3778,N_1896,N_1328);
nand U3779 (N_3779,N_2278,N_1141);
and U3780 (N_3780,N_427,N_627);
nor U3781 (N_3781,N_492,N_643);
and U3782 (N_3782,N_456,N_678);
or U3783 (N_3783,N_537,N_1491);
nor U3784 (N_3784,N_752,N_1169);
or U3785 (N_3785,N_1574,N_1727);
and U3786 (N_3786,N_1507,N_444);
or U3787 (N_3787,N_1936,N_1406);
nor U3788 (N_3788,N_834,N_1115);
nand U3789 (N_3789,N_2276,N_1747);
nand U3790 (N_3790,N_650,N_1102);
and U3791 (N_3791,N_198,N_493);
nand U3792 (N_3792,N_350,N_728);
nand U3793 (N_3793,N_134,N_189);
or U3794 (N_3794,N_762,N_1539);
and U3795 (N_3795,N_1147,N_1193);
or U3796 (N_3796,N_1709,N_92);
nand U3797 (N_3797,N_1269,N_1267);
and U3798 (N_3798,N_236,N_981);
nand U3799 (N_3799,N_2437,N_1190);
nand U3800 (N_3800,N_718,N_1415);
or U3801 (N_3801,N_372,N_1693);
or U3802 (N_3802,N_189,N_2379);
nand U3803 (N_3803,N_2409,N_1519);
xor U3804 (N_3804,N_1540,N_175);
nor U3805 (N_3805,N_1160,N_1436);
nor U3806 (N_3806,N_299,N_2439);
or U3807 (N_3807,N_1265,N_530);
xnor U3808 (N_3808,N_2332,N_2158);
or U3809 (N_3809,N_349,N_21);
xor U3810 (N_3810,N_1896,N_644);
nand U3811 (N_3811,N_2118,N_1781);
nor U3812 (N_3812,N_2405,N_1103);
nor U3813 (N_3813,N_2473,N_2349);
or U3814 (N_3814,N_867,N_1593);
nand U3815 (N_3815,N_1341,N_2187);
and U3816 (N_3816,N_2042,N_1226);
or U3817 (N_3817,N_1912,N_963);
nand U3818 (N_3818,N_410,N_1366);
and U3819 (N_3819,N_15,N_1190);
and U3820 (N_3820,N_1543,N_1547);
or U3821 (N_3821,N_1000,N_1982);
nand U3822 (N_3822,N_2242,N_2244);
nand U3823 (N_3823,N_856,N_1361);
and U3824 (N_3824,N_2149,N_1236);
nand U3825 (N_3825,N_463,N_2406);
or U3826 (N_3826,N_2003,N_58);
nor U3827 (N_3827,N_1463,N_2443);
and U3828 (N_3828,N_2081,N_128);
nor U3829 (N_3829,N_1204,N_2410);
and U3830 (N_3830,N_2370,N_2420);
and U3831 (N_3831,N_1756,N_2042);
xnor U3832 (N_3832,N_1590,N_2209);
and U3833 (N_3833,N_1613,N_1778);
or U3834 (N_3834,N_500,N_1392);
or U3835 (N_3835,N_1098,N_2231);
nand U3836 (N_3836,N_583,N_1447);
nor U3837 (N_3837,N_1485,N_222);
or U3838 (N_3838,N_1508,N_221);
nor U3839 (N_3839,N_1391,N_1808);
and U3840 (N_3840,N_1286,N_2414);
xor U3841 (N_3841,N_776,N_2221);
nor U3842 (N_3842,N_2409,N_1645);
and U3843 (N_3843,N_2467,N_924);
nor U3844 (N_3844,N_2320,N_2354);
or U3845 (N_3845,N_2452,N_923);
or U3846 (N_3846,N_232,N_595);
nand U3847 (N_3847,N_1452,N_417);
and U3848 (N_3848,N_1289,N_512);
or U3849 (N_3849,N_73,N_1454);
nand U3850 (N_3850,N_212,N_1835);
nand U3851 (N_3851,N_2293,N_1573);
nand U3852 (N_3852,N_1361,N_2358);
nor U3853 (N_3853,N_1825,N_712);
or U3854 (N_3854,N_819,N_1012);
and U3855 (N_3855,N_420,N_2064);
nor U3856 (N_3856,N_267,N_1377);
xnor U3857 (N_3857,N_235,N_315);
and U3858 (N_3858,N_1170,N_1300);
nor U3859 (N_3859,N_407,N_1990);
nand U3860 (N_3860,N_2013,N_2440);
or U3861 (N_3861,N_2155,N_1808);
xor U3862 (N_3862,N_923,N_1833);
nand U3863 (N_3863,N_2074,N_1661);
nor U3864 (N_3864,N_249,N_2313);
nor U3865 (N_3865,N_1005,N_1692);
and U3866 (N_3866,N_2147,N_1387);
or U3867 (N_3867,N_133,N_572);
and U3868 (N_3868,N_903,N_1220);
and U3869 (N_3869,N_844,N_1330);
nand U3870 (N_3870,N_960,N_1397);
and U3871 (N_3871,N_1266,N_1820);
xor U3872 (N_3872,N_189,N_2484);
and U3873 (N_3873,N_1333,N_1717);
nand U3874 (N_3874,N_1215,N_534);
or U3875 (N_3875,N_941,N_614);
nor U3876 (N_3876,N_1231,N_1316);
nand U3877 (N_3877,N_1122,N_719);
nor U3878 (N_3878,N_2153,N_511);
or U3879 (N_3879,N_182,N_159);
nand U3880 (N_3880,N_1515,N_1666);
and U3881 (N_3881,N_2341,N_775);
or U3882 (N_3882,N_1617,N_834);
xnor U3883 (N_3883,N_2331,N_823);
nor U3884 (N_3884,N_564,N_146);
nor U3885 (N_3885,N_2356,N_1282);
xor U3886 (N_3886,N_337,N_12);
and U3887 (N_3887,N_1703,N_621);
and U3888 (N_3888,N_1329,N_1381);
nand U3889 (N_3889,N_917,N_1381);
xor U3890 (N_3890,N_787,N_1103);
nor U3891 (N_3891,N_469,N_305);
or U3892 (N_3892,N_1051,N_247);
or U3893 (N_3893,N_2298,N_1023);
xor U3894 (N_3894,N_2483,N_1268);
nor U3895 (N_3895,N_1466,N_745);
nand U3896 (N_3896,N_646,N_472);
xnor U3897 (N_3897,N_1697,N_228);
xnor U3898 (N_3898,N_2467,N_28);
or U3899 (N_3899,N_1270,N_1266);
or U3900 (N_3900,N_1848,N_1587);
or U3901 (N_3901,N_1231,N_724);
xor U3902 (N_3902,N_689,N_813);
or U3903 (N_3903,N_1223,N_1809);
and U3904 (N_3904,N_1028,N_2110);
nor U3905 (N_3905,N_2390,N_1162);
and U3906 (N_3906,N_2346,N_1881);
nand U3907 (N_3907,N_1504,N_1457);
and U3908 (N_3908,N_2128,N_372);
or U3909 (N_3909,N_466,N_708);
xnor U3910 (N_3910,N_1905,N_951);
nand U3911 (N_3911,N_744,N_1930);
nor U3912 (N_3912,N_317,N_178);
nor U3913 (N_3913,N_2040,N_46);
xnor U3914 (N_3914,N_935,N_1974);
or U3915 (N_3915,N_1419,N_2398);
or U3916 (N_3916,N_1425,N_325);
and U3917 (N_3917,N_2222,N_2051);
or U3918 (N_3918,N_1301,N_1012);
and U3919 (N_3919,N_127,N_1377);
nor U3920 (N_3920,N_1352,N_2442);
or U3921 (N_3921,N_1814,N_34);
and U3922 (N_3922,N_408,N_1315);
and U3923 (N_3923,N_986,N_2025);
nand U3924 (N_3924,N_1359,N_794);
and U3925 (N_3925,N_767,N_2267);
and U3926 (N_3926,N_1211,N_807);
nor U3927 (N_3927,N_1365,N_715);
nor U3928 (N_3928,N_1979,N_1855);
xnor U3929 (N_3929,N_2450,N_814);
nand U3930 (N_3930,N_2227,N_1290);
or U3931 (N_3931,N_407,N_2212);
xnor U3932 (N_3932,N_814,N_2254);
nand U3933 (N_3933,N_1566,N_1949);
and U3934 (N_3934,N_1931,N_203);
and U3935 (N_3935,N_1976,N_1561);
and U3936 (N_3936,N_1250,N_1471);
and U3937 (N_3937,N_1000,N_703);
and U3938 (N_3938,N_1604,N_251);
or U3939 (N_3939,N_2244,N_2297);
and U3940 (N_3940,N_1663,N_1175);
and U3941 (N_3941,N_2495,N_1217);
or U3942 (N_3942,N_2187,N_741);
nand U3943 (N_3943,N_647,N_917);
nand U3944 (N_3944,N_1938,N_1039);
nor U3945 (N_3945,N_1193,N_2486);
nor U3946 (N_3946,N_2461,N_427);
nand U3947 (N_3947,N_798,N_1935);
and U3948 (N_3948,N_2288,N_282);
and U3949 (N_3949,N_1093,N_29);
nor U3950 (N_3950,N_963,N_1384);
nand U3951 (N_3951,N_1039,N_2322);
nand U3952 (N_3952,N_1810,N_2005);
nor U3953 (N_3953,N_2195,N_29);
and U3954 (N_3954,N_2470,N_853);
nor U3955 (N_3955,N_391,N_392);
nor U3956 (N_3956,N_563,N_23);
xnor U3957 (N_3957,N_1731,N_2112);
or U3958 (N_3958,N_354,N_1398);
or U3959 (N_3959,N_1436,N_1523);
xnor U3960 (N_3960,N_1603,N_2014);
or U3961 (N_3961,N_2468,N_1587);
and U3962 (N_3962,N_2323,N_2136);
nand U3963 (N_3963,N_368,N_833);
nor U3964 (N_3964,N_571,N_316);
or U3965 (N_3965,N_1091,N_1128);
nor U3966 (N_3966,N_805,N_1876);
nand U3967 (N_3967,N_504,N_2293);
or U3968 (N_3968,N_1251,N_2351);
and U3969 (N_3969,N_1128,N_2002);
nand U3970 (N_3970,N_2197,N_1963);
and U3971 (N_3971,N_578,N_1621);
nand U3972 (N_3972,N_1831,N_1535);
or U3973 (N_3973,N_1568,N_1976);
xor U3974 (N_3974,N_938,N_647);
and U3975 (N_3975,N_498,N_2318);
and U3976 (N_3976,N_1446,N_1625);
nor U3977 (N_3977,N_364,N_1255);
xor U3978 (N_3978,N_822,N_577);
and U3979 (N_3979,N_2242,N_1876);
nor U3980 (N_3980,N_1601,N_467);
or U3981 (N_3981,N_1943,N_450);
nand U3982 (N_3982,N_1254,N_858);
and U3983 (N_3983,N_532,N_1164);
nor U3984 (N_3984,N_621,N_600);
and U3985 (N_3985,N_2305,N_102);
or U3986 (N_3986,N_1418,N_683);
nor U3987 (N_3987,N_846,N_590);
nor U3988 (N_3988,N_1189,N_2347);
and U3989 (N_3989,N_1468,N_2305);
or U3990 (N_3990,N_1173,N_704);
nor U3991 (N_3991,N_254,N_2495);
or U3992 (N_3992,N_850,N_1883);
nand U3993 (N_3993,N_1445,N_468);
or U3994 (N_3994,N_245,N_2454);
and U3995 (N_3995,N_2032,N_7);
and U3996 (N_3996,N_2182,N_1761);
and U3997 (N_3997,N_690,N_1423);
and U3998 (N_3998,N_1468,N_1370);
and U3999 (N_3999,N_976,N_215);
nand U4000 (N_4000,N_543,N_1963);
or U4001 (N_4001,N_387,N_2265);
nor U4002 (N_4002,N_732,N_709);
xnor U4003 (N_4003,N_1741,N_1737);
nor U4004 (N_4004,N_598,N_317);
or U4005 (N_4005,N_1369,N_1951);
and U4006 (N_4006,N_2070,N_2484);
nor U4007 (N_4007,N_1076,N_1465);
nor U4008 (N_4008,N_671,N_939);
or U4009 (N_4009,N_429,N_1626);
and U4010 (N_4010,N_2424,N_885);
nor U4011 (N_4011,N_1551,N_695);
nand U4012 (N_4012,N_1667,N_213);
nor U4013 (N_4013,N_100,N_2033);
nor U4014 (N_4014,N_2446,N_1633);
nand U4015 (N_4015,N_2330,N_1576);
or U4016 (N_4016,N_373,N_732);
or U4017 (N_4017,N_674,N_1202);
or U4018 (N_4018,N_1345,N_1020);
nand U4019 (N_4019,N_1211,N_36);
nor U4020 (N_4020,N_36,N_1176);
or U4021 (N_4021,N_27,N_1811);
nand U4022 (N_4022,N_897,N_2436);
and U4023 (N_4023,N_1180,N_1957);
and U4024 (N_4024,N_13,N_2047);
or U4025 (N_4025,N_273,N_1160);
or U4026 (N_4026,N_2380,N_1298);
or U4027 (N_4027,N_691,N_1107);
xnor U4028 (N_4028,N_607,N_2066);
xnor U4029 (N_4029,N_42,N_704);
and U4030 (N_4030,N_1442,N_2278);
nand U4031 (N_4031,N_869,N_1463);
and U4032 (N_4032,N_1606,N_804);
and U4033 (N_4033,N_1779,N_166);
xor U4034 (N_4034,N_659,N_1251);
nor U4035 (N_4035,N_336,N_2117);
nor U4036 (N_4036,N_1131,N_679);
nor U4037 (N_4037,N_2470,N_1161);
nand U4038 (N_4038,N_113,N_525);
nand U4039 (N_4039,N_282,N_357);
and U4040 (N_4040,N_2012,N_793);
nand U4041 (N_4041,N_754,N_931);
nor U4042 (N_4042,N_1472,N_419);
nor U4043 (N_4043,N_1322,N_2124);
and U4044 (N_4044,N_462,N_395);
nand U4045 (N_4045,N_414,N_418);
or U4046 (N_4046,N_1222,N_1769);
xnor U4047 (N_4047,N_582,N_329);
xnor U4048 (N_4048,N_666,N_2150);
nand U4049 (N_4049,N_1863,N_1486);
xnor U4050 (N_4050,N_1038,N_1717);
or U4051 (N_4051,N_294,N_1899);
nand U4052 (N_4052,N_282,N_1210);
or U4053 (N_4053,N_2481,N_2295);
xor U4054 (N_4054,N_256,N_1365);
or U4055 (N_4055,N_2458,N_2383);
and U4056 (N_4056,N_2383,N_2266);
xnor U4057 (N_4057,N_1120,N_1306);
and U4058 (N_4058,N_233,N_905);
nand U4059 (N_4059,N_235,N_1849);
and U4060 (N_4060,N_902,N_79);
nand U4061 (N_4061,N_983,N_2245);
xnor U4062 (N_4062,N_2077,N_207);
xor U4063 (N_4063,N_1402,N_1714);
nand U4064 (N_4064,N_1283,N_1243);
nand U4065 (N_4065,N_1894,N_1413);
or U4066 (N_4066,N_724,N_255);
nand U4067 (N_4067,N_2333,N_1681);
or U4068 (N_4068,N_631,N_1264);
and U4069 (N_4069,N_2269,N_1545);
nor U4070 (N_4070,N_821,N_1192);
and U4071 (N_4071,N_362,N_1442);
nand U4072 (N_4072,N_1641,N_1959);
nor U4073 (N_4073,N_2294,N_344);
nor U4074 (N_4074,N_197,N_1882);
and U4075 (N_4075,N_1398,N_2433);
nor U4076 (N_4076,N_1844,N_146);
nand U4077 (N_4077,N_661,N_682);
nor U4078 (N_4078,N_149,N_1416);
nor U4079 (N_4079,N_789,N_1401);
and U4080 (N_4080,N_785,N_1344);
and U4081 (N_4081,N_2371,N_2318);
nand U4082 (N_4082,N_195,N_426);
and U4083 (N_4083,N_1578,N_640);
nor U4084 (N_4084,N_2454,N_292);
and U4085 (N_4085,N_1513,N_313);
or U4086 (N_4086,N_758,N_623);
nand U4087 (N_4087,N_1271,N_824);
xor U4088 (N_4088,N_1920,N_1686);
nor U4089 (N_4089,N_572,N_1284);
nand U4090 (N_4090,N_102,N_201);
nand U4091 (N_4091,N_789,N_1134);
nand U4092 (N_4092,N_1074,N_1958);
or U4093 (N_4093,N_408,N_865);
and U4094 (N_4094,N_1371,N_608);
nand U4095 (N_4095,N_1383,N_2178);
and U4096 (N_4096,N_1787,N_501);
and U4097 (N_4097,N_520,N_1188);
and U4098 (N_4098,N_2350,N_749);
or U4099 (N_4099,N_2196,N_1705);
nand U4100 (N_4100,N_1566,N_353);
or U4101 (N_4101,N_404,N_1947);
nand U4102 (N_4102,N_2329,N_2083);
or U4103 (N_4103,N_647,N_2132);
nand U4104 (N_4104,N_1787,N_228);
or U4105 (N_4105,N_1872,N_173);
xor U4106 (N_4106,N_108,N_909);
xnor U4107 (N_4107,N_279,N_2078);
nor U4108 (N_4108,N_1110,N_2130);
xnor U4109 (N_4109,N_602,N_1275);
and U4110 (N_4110,N_2283,N_227);
nor U4111 (N_4111,N_5,N_2408);
and U4112 (N_4112,N_1418,N_2464);
nand U4113 (N_4113,N_1215,N_1783);
or U4114 (N_4114,N_1230,N_1486);
and U4115 (N_4115,N_1465,N_1647);
and U4116 (N_4116,N_1911,N_192);
and U4117 (N_4117,N_1236,N_416);
xnor U4118 (N_4118,N_956,N_1444);
nand U4119 (N_4119,N_94,N_2317);
or U4120 (N_4120,N_2381,N_616);
and U4121 (N_4121,N_1354,N_1349);
nand U4122 (N_4122,N_389,N_1082);
nand U4123 (N_4123,N_1987,N_2408);
and U4124 (N_4124,N_1847,N_688);
nand U4125 (N_4125,N_340,N_602);
or U4126 (N_4126,N_1261,N_458);
or U4127 (N_4127,N_1532,N_346);
nor U4128 (N_4128,N_434,N_41);
nor U4129 (N_4129,N_1101,N_572);
and U4130 (N_4130,N_1903,N_2260);
nand U4131 (N_4131,N_1727,N_2474);
and U4132 (N_4132,N_2072,N_223);
nor U4133 (N_4133,N_2371,N_2233);
nand U4134 (N_4134,N_564,N_388);
xnor U4135 (N_4135,N_544,N_2175);
nand U4136 (N_4136,N_485,N_954);
nor U4137 (N_4137,N_968,N_1824);
and U4138 (N_4138,N_1239,N_2454);
and U4139 (N_4139,N_110,N_1204);
and U4140 (N_4140,N_28,N_2247);
nand U4141 (N_4141,N_1990,N_2198);
and U4142 (N_4142,N_2393,N_843);
and U4143 (N_4143,N_1512,N_1039);
and U4144 (N_4144,N_1092,N_1125);
and U4145 (N_4145,N_274,N_1528);
or U4146 (N_4146,N_854,N_1585);
or U4147 (N_4147,N_1392,N_1499);
and U4148 (N_4148,N_2319,N_2432);
or U4149 (N_4149,N_1998,N_1463);
nor U4150 (N_4150,N_466,N_175);
or U4151 (N_4151,N_1980,N_5);
nor U4152 (N_4152,N_2421,N_2108);
or U4153 (N_4153,N_1682,N_1434);
and U4154 (N_4154,N_230,N_343);
nand U4155 (N_4155,N_2309,N_278);
and U4156 (N_4156,N_1847,N_1391);
nand U4157 (N_4157,N_226,N_948);
nor U4158 (N_4158,N_1176,N_1728);
nor U4159 (N_4159,N_981,N_2224);
or U4160 (N_4160,N_520,N_1593);
nor U4161 (N_4161,N_2226,N_1645);
nand U4162 (N_4162,N_918,N_1089);
or U4163 (N_4163,N_220,N_1512);
and U4164 (N_4164,N_643,N_2485);
nand U4165 (N_4165,N_442,N_526);
and U4166 (N_4166,N_968,N_847);
nor U4167 (N_4167,N_2297,N_2299);
and U4168 (N_4168,N_2144,N_1684);
or U4169 (N_4169,N_1762,N_1239);
and U4170 (N_4170,N_1055,N_1704);
and U4171 (N_4171,N_2127,N_43);
and U4172 (N_4172,N_559,N_685);
nor U4173 (N_4173,N_817,N_1108);
nor U4174 (N_4174,N_1305,N_735);
or U4175 (N_4175,N_242,N_2237);
or U4176 (N_4176,N_1347,N_2077);
or U4177 (N_4177,N_1337,N_1602);
nor U4178 (N_4178,N_2142,N_9);
or U4179 (N_4179,N_275,N_1387);
or U4180 (N_4180,N_1741,N_2088);
nor U4181 (N_4181,N_1051,N_1020);
and U4182 (N_4182,N_2014,N_999);
nor U4183 (N_4183,N_265,N_1502);
nor U4184 (N_4184,N_2404,N_1687);
or U4185 (N_4185,N_128,N_337);
or U4186 (N_4186,N_2201,N_369);
xnor U4187 (N_4187,N_311,N_1034);
and U4188 (N_4188,N_1412,N_1993);
nand U4189 (N_4189,N_2142,N_1974);
and U4190 (N_4190,N_1180,N_1806);
or U4191 (N_4191,N_1816,N_1444);
and U4192 (N_4192,N_1955,N_1023);
xor U4193 (N_4193,N_742,N_1545);
and U4194 (N_4194,N_1833,N_1476);
and U4195 (N_4195,N_1466,N_208);
or U4196 (N_4196,N_553,N_1902);
or U4197 (N_4197,N_870,N_2229);
nor U4198 (N_4198,N_2475,N_280);
and U4199 (N_4199,N_2093,N_497);
nand U4200 (N_4200,N_240,N_2195);
and U4201 (N_4201,N_998,N_1452);
and U4202 (N_4202,N_462,N_1487);
and U4203 (N_4203,N_2201,N_1635);
and U4204 (N_4204,N_1735,N_1838);
nor U4205 (N_4205,N_1523,N_1273);
nand U4206 (N_4206,N_1772,N_430);
or U4207 (N_4207,N_2331,N_1738);
xor U4208 (N_4208,N_2374,N_1451);
nand U4209 (N_4209,N_2046,N_1455);
xor U4210 (N_4210,N_191,N_2049);
nand U4211 (N_4211,N_2386,N_8);
nor U4212 (N_4212,N_1009,N_1329);
or U4213 (N_4213,N_2334,N_2047);
nand U4214 (N_4214,N_1813,N_141);
nor U4215 (N_4215,N_2355,N_2193);
nor U4216 (N_4216,N_1518,N_1225);
nor U4217 (N_4217,N_168,N_2198);
or U4218 (N_4218,N_1313,N_2222);
or U4219 (N_4219,N_271,N_2042);
nor U4220 (N_4220,N_1186,N_850);
nand U4221 (N_4221,N_724,N_1100);
nand U4222 (N_4222,N_772,N_661);
and U4223 (N_4223,N_2307,N_1013);
nand U4224 (N_4224,N_843,N_1984);
nand U4225 (N_4225,N_2058,N_2282);
or U4226 (N_4226,N_2338,N_2072);
or U4227 (N_4227,N_84,N_247);
nand U4228 (N_4228,N_1736,N_1375);
or U4229 (N_4229,N_1284,N_245);
or U4230 (N_4230,N_1249,N_342);
and U4231 (N_4231,N_422,N_134);
and U4232 (N_4232,N_1551,N_423);
and U4233 (N_4233,N_436,N_1739);
and U4234 (N_4234,N_91,N_67);
or U4235 (N_4235,N_157,N_1933);
xor U4236 (N_4236,N_2263,N_1428);
or U4237 (N_4237,N_1562,N_1352);
xor U4238 (N_4238,N_1489,N_1203);
xor U4239 (N_4239,N_1199,N_1168);
xnor U4240 (N_4240,N_1982,N_228);
nand U4241 (N_4241,N_1726,N_1077);
nand U4242 (N_4242,N_483,N_1088);
xnor U4243 (N_4243,N_1812,N_1108);
and U4244 (N_4244,N_691,N_1224);
or U4245 (N_4245,N_822,N_1393);
or U4246 (N_4246,N_1479,N_2198);
xnor U4247 (N_4247,N_617,N_777);
nor U4248 (N_4248,N_28,N_2187);
or U4249 (N_4249,N_443,N_2094);
nor U4250 (N_4250,N_1842,N_1228);
nor U4251 (N_4251,N_905,N_2326);
nand U4252 (N_4252,N_1464,N_1831);
and U4253 (N_4253,N_664,N_1548);
xnor U4254 (N_4254,N_2206,N_1501);
or U4255 (N_4255,N_1018,N_1183);
nand U4256 (N_4256,N_1934,N_386);
or U4257 (N_4257,N_269,N_2421);
nand U4258 (N_4258,N_643,N_1469);
xor U4259 (N_4259,N_2109,N_1990);
nand U4260 (N_4260,N_2323,N_342);
nand U4261 (N_4261,N_2280,N_1153);
nand U4262 (N_4262,N_1049,N_2388);
nand U4263 (N_4263,N_1922,N_2154);
nor U4264 (N_4264,N_1871,N_1357);
and U4265 (N_4265,N_423,N_309);
and U4266 (N_4266,N_905,N_225);
nand U4267 (N_4267,N_1837,N_1503);
or U4268 (N_4268,N_713,N_301);
nand U4269 (N_4269,N_440,N_1549);
nand U4270 (N_4270,N_132,N_2237);
nor U4271 (N_4271,N_1855,N_2414);
or U4272 (N_4272,N_1757,N_1988);
and U4273 (N_4273,N_1138,N_1851);
nor U4274 (N_4274,N_194,N_1542);
nand U4275 (N_4275,N_2374,N_1502);
nor U4276 (N_4276,N_1913,N_1785);
nor U4277 (N_4277,N_1983,N_1576);
or U4278 (N_4278,N_1417,N_219);
or U4279 (N_4279,N_1943,N_2287);
nor U4280 (N_4280,N_1022,N_715);
or U4281 (N_4281,N_1210,N_2419);
nand U4282 (N_4282,N_384,N_1051);
or U4283 (N_4283,N_1475,N_2413);
nor U4284 (N_4284,N_2412,N_1364);
or U4285 (N_4285,N_1028,N_692);
nor U4286 (N_4286,N_647,N_832);
and U4287 (N_4287,N_1315,N_1327);
and U4288 (N_4288,N_1544,N_2369);
nand U4289 (N_4289,N_136,N_1034);
or U4290 (N_4290,N_994,N_508);
xnor U4291 (N_4291,N_2084,N_1436);
and U4292 (N_4292,N_805,N_1646);
and U4293 (N_4293,N_1137,N_252);
and U4294 (N_4294,N_2447,N_900);
or U4295 (N_4295,N_2399,N_924);
nand U4296 (N_4296,N_2139,N_61);
and U4297 (N_4297,N_2135,N_1069);
or U4298 (N_4298,N_1541,N_743);
nor U4299 (N_4299,N_410,N_1399);
or U4300 (N_4300,N_1661,N_238);
nand U4301 (N_4301,N_1499,N_1319);
and U4302 (N_4302,N_856,N_309);
nor U4303 (N_4303,N_1080,N_1539);
nor U4304 (N_4304,N_1101,N_1549);
or U4305 (N_4305,N_2147,N_1222);
and U4306 (N_4306,N_165,N_1223);
and U4307 (N_4307,N_1352,N_2063);
and U4308 (N_4308,N_656,N_1916);
nor U4309 (N_4309,N_2436,N_131);
nor U4310 (N_4310,N_1622,N_2481);
and U4311 (N_4311,N_2388,N_469);
nor U4312 (N_4312,N_1417,N_1495);
nor U4313 (N_4313,N_593,N_797);
nor U4314 (N_4314,N_989,N_1016);
nor U4315 (N_4315,N_1013,N_1466);
and U4316 (N_4316,N_2098,N_2142);
or U4317 (N_4317,N_1681,N_290);
and U4318 (N_4318,N_1036,N_364);
and U4319 (N_4319,N_1297,N_1661);
nand U4320 (N_4320,N_107,N_911);
and U4321 (N_4321,N_493,N_865);
and U4322 (N_4322,N_511,N_1961);
xor U4323 (N_4323,N_1932,N_1266);
and U4324 (N_4324,N_1991,N_1771);
nor U4325 (N_4325,N_1649,N_1441);
nor U4326 (N_4326,N_2458,N_957);
nand U4327 (N_4327,N_47,N_576);
nand U4328 (N_4328,N_1584,N_2274);
nor U4329 (N_4329,N_1899,N_830);
nor U4330 (N_4330,N_616,N_2016);
nand U4331 (N_4331,N_2305,N_2347);
or U4332 (N_4332,N_957,N_1531);
nor U4333 (N_4333,N_950,N_1098);
nand U4334 (N_4334,N_2352,N_2136);
xor U4335 (N_4335,N_842,N_858);
nor U4336 (N_4336,N_2492,N_903);
xnor U4337 (N_4337,N_1724,N_107);
or U4338 (N_4338,N_2302,N_1446);
or U4339 (N_4339,N_2033,N_2208);
and U4340 (N_4340,N_1026,N_349);
nand U4341 (N_4341,N_587,N_2303);
and U4342 (N_4342,N_1217,N_916);
nor U4343 (N_4343,N_712,N_2325);
or U4344 (N_4344,N_645,N_368);
and U4345 (N_4345,N_1980,N_2038);
nor U4346 (N_4346,N_848,N_371);
and U4347 (N_4347,N_1452,N_822);
or U4348 (N_4348,N_676,N_1355);
nor U4349 (N_4349,N_615,N_2136);
or U4350 (N_4350,N_2010,N_996);
and U4351 (N_4351,N_1123,N_385);
and U4352 (N_4352,N_347,N_2078);
nand U4353 (N_4353,N_939,N_224);
and U4354 (N_4354,N_1558,N_874);
nor U4355 (N_4355,N_1091,N_2243);
or U4356 (N_4356,N_921,N_1757);
or U4357 (N_4357,N_723,N_2140);
xor U4358 (N_4358,N_1169,N_2263);
nand U4359 (N_4359,N_800,N_974);
or U4360 (N_4360,N_2372,N_1009);
and U4361 (N_4361,N_2195,N_2411);
nand U4362 (N_4362,N_318,N_1664);
and U4363 (N_4363,N_1720,N_2415);
nand U4364 (N_4364,N_2002,N_1044);
nor U4365 (N_4365,N_1761,N_1178);
xor U4366 (N_4366,N_1364,N_1547);
nor U4367 (N_4367,N_1166,N_1233);
and U4368 (N_4368,N_815,N_1693);
nor U4369 (N_4369,N_1364,N_1421);
nand U4370 (N_4370,N_1095,N_1711);
xor U4371 (N_4371,N_403,N_1903);
nand U4372 (N_4372,N_715,N_1955);
and U4373 (N_4373,N_1779,N_2080);
nor U4374 (N_4374,N_994,N_954);
nand U4375 (N_4375,N_2126,N_311);
or U4376 (N_4376,N_291,N_1358);
nor U4377 (N_4377,N_392,N_754);
or U4378 (N_4378,N_1671,N_1968);
and U4379 (N_4379,N_508,N_2182);
nor U4380 (N_4380,N_1839,N_868);
or U4381 (N_4381,N_1183,N_1779);
or U4382 (N_4382,N_344,N_10);
or U4383 (N_4383,N_2390,N_622);
or U4384 (N_4384,N_2020,N_132);
and U4385 (N_4385,N_1873,N_2084);
nand U4386 (N_4386,N_1387,N_740);
nor U4387 (N_4387,N_523,N_2305);
or U4388 (N_4388,N_1460,N_1763);
and U4389 (N_4389,N_2011,N_1122);
and U4390 (N_4390,N_1380,N_1568);
or U4391 (N_4391,N_1158,N_516);
and U4392 (N_4392,N_1303,N_1845);
nor U4393 (N_4393,N_1038,N_1294);
and U4394 (N_4394,N_2317,N_1836);
nand U4395 (N_4395,N_58,N_1122);
nand U4396 (N_4396,N_1433,N_1059);
or U4397 (N_4397,N_59,N_1464);
nor U4398 (N_4398,N_2178,N_120);
nor U4399 (N_4399,N_1563,N_219);
nor U4400 (N_4400,N_2288,N_549);
xor U4401 (N_4401,N_1826,N_1278);
nor U4402 (N_4402,N_1859,N_1719);
or U4403 (N_4403,N_1981,N_2271);
nor U4404 (N_4404,N_1540,N_744);
nor U4405 (N_4405,N_1176,N_1015);
or U4406 (N_4406,N_756,N_1281);
and U4407 (N_4407,N_797,N_1608);
nand U4408 (N_4408,N_1650,N_37);
and U4409 (N_4409,N_1345,N_747);
xor U4410 (N_4410,N_1930,N_2351);
nand U4411 (N_4411,N_659,N_1428);
or U4412 (N_4412,N_396,N_415);
or U4413 (N_4413,N_669,N_0);
nand U4414 (N_4414,N_498,N_1346);
and U4415 (N_4415,N_216,N_532);
and U4416 (N_4416,N_2016,N_995);
or U4417 (N_4417,N_2477,N_1825);
and U4418 (N_4418,N_724,N_2381);
nor U4419 (N_4419,N_2080,N_550);
and U4420 (N_4420,N_1964,N_2232);
nand U4421 (N_4421,N_1770,N_538);
nor U4422 (N_4422,N_1310,N_1890);
and U4423 (N_4423,N_1902,N_1033);
and U4424 (N_4424,N_2412,N_466);
and U4425 (N_4425,N_1619,N_920);
or U4426 (N_4426,N_2240,N_1406);
nor U4427 (N_4427,N_710,N_797);
xnor U4428 (N_4428,N_43,N_1368);
nor U4429 (N_4429,N_841,N_2071);
nand U4430 (N_4430,N_1196,N_402);
nand U4431 (N_4431,N_2056,N_477);
or U4432 (N_4432,N_2041,N_1877);
and U4433 (N_4433,N_921,N_531);
and U4434 (N_4434,N_195,N_889);
and U4435 (N_4435,N_787,N_28);
xor U4436 (N_4436,N_1934,N_2074);
nor U4437 (N_4437,N_2418,N_403);
nor U4438 (N_4438,N_292,N_1571);
nand U4439 (N_4439,N_1691,N_1906);
or U4440 (N_4440,N_1844,N_1529);
and U4441 (N_4441,N_308,N_567);
and U4442 (N_4442,N_499,N_1571);
nor U4443 (N_4443,N_1090,N_29);
or U4444 (N_4444,N_1425,N_2271);
nand U4445 (N_4445,N_8,N_675);
nand U4446 (N_4446,N_2485,N_644);
or U4447 (N_4447,N_454,N_955);
or U4448 (N_4448,N_877,N_962);
nor U4449 (N_4449,N_1724,N_2212);
and U4450 (N_4450,N_668,N_1631);
xor U4451 (N_4451,N_377,N_1290);
nand U4452 (N_4452,N_499,N_1951);
xnor U4453 (N_4453,N_2180,N_2165);
and U4454 (N_4454,N_2405,N_1938);
nor U4455 (N_4455,N_882,N_2147);
and U4456 (N_4456,N_1576,N_530);
nand U4457 (N_4457,N_1271,N_1981);
nand U4458 (N_4458,N_448,N_1150);
xnor U4459 (N_4459,N_1719,N_1792);
or U4460 (N_4460,N_1588,N_851);
nand U4461 (N_4461,N_83,N_81);
nor U4462 (N_4462,N_382,N_441);
nand U4463 (N_4463,N_1257,N_891);
nor U4464 (N_4464,N_160,N_2142);
nand U4465 (N_4465,N_1020,N_1891);
nand U4466 (N_4466,N_1262,N_511);
or U4467 (N_4467,N_933,N_1691);
nor U4468 (N_4468,N_1113,N_958);
nand U4469 (N_4469,N_1318,N_119);
nand U4470 (N_4470,N_1307,N_191);
or U4471 (N_4471,N_942,N_1349);
and U4472 (N_4472,N_50,N_2025);
nand U4473 (N_4473,N_30,N_451);
nor U4474 (N_4474,N_1840,N_1019);
or U4475 (N_4475,N_33,N_1837);
and U4476 (N_4476,N_1156,N_1976);
nand U4477 (N_4477,N_1820,N_313);
nand U4478 (N_4478,N_1825,N_364);
nand U4479 (N_4479,N_2407,N_2424);
xnor U4480 (N_4480,N_137,N_1219);
nor U4481 (N_4481,N_1627,N_377);
nor U4482 (N_4482,N_2435,N_2171);
nor U4483 (N_4483,N_512,N_350);
xnor U4484 (N_4484,N_839,N_1152);
and U4485 (N_4485,N_1750,N_1524);
nor U4486 (N_4486,N_2147,N_2112);
or U4487 (N_4487,N_1231,N_1037);
or U4488 (N_4488,N_1501,N_1996);
or U4489 (N_4489,N_1414,N_425);
or U4490 (N_4490,N_626,N_769);
or U4491 (N_4491,N_403,N_813);
or U4492 (N_4492,N_1489,N_16);
or U4493 (N_4493,N_1451,N_2213);
and U4494 (N_4494,N_1887,N_706);
xnor U4495 (N_4495,N_2042,N_1125);
nor U4496 (N_4496,N_508,N_2068);
nor U4497 (N_4497,N_1822,N_360);
nand U4498 (N_4498,N_2323,N_432);
and U4499 (N_4499,N_443,N_2120);
nand U4500 (N_4500,N_638,N_1606);
and U4501 (N_4501,N_2453,N_1451);
nand U4502 (N_4502,N_2459,N_1933);
or U4503 (N_4503,N_2459,N_1625);
nor U4504 (N_4504,N_1321,N_1040);
nand U4505 (N_4505,N_1898,N_29);
nand U4506 (N_4506,N_900,N_1175);
nand U4507 (N_4507,N_1926,N_1809);
or U4508 (N_4508,N_1366,N_129);
nor U4509 (N_4509,N_1882,N_21);
and U4510 (N_4510,N_1761,N_1471);
or U4511 (N_4511,N_2275,N_957);
or U4512 (N_4512,N_1363,N_556);
nand U4513 (N_4513,N_2389,N_948);
or U4514 (N_4514,N_2382,N_2034);
nor U4515 (N_4515,N_346,N_1304);
nor U4516 (N_4516,N_311,N_2142);
nand U4517 (N_4517,N_1228,N_749);
and U4518 (N_4518,N_1901,N_2250);
and U4519 (N_4519,N_1903,N_2267);
nor U4520 (N_4520,N_1116,N_1230);
nand U4521 (N_4521,N_2344,N_2278);
or U4522 (N_4522,N_1246,N_355);
nand U4523 (N_4523,N_740,N_914);
and U4524 (N_4524,N_776,N_2469);
nand U4525 (N_4525,N_1924,N_1938);
and U4526 (N_4526,N_1047,N_1399);
nor U4527 (N_4527,N_2096,N_222);
or U4528 (N_4528,N_236,N_282);
xnor U4529 (N_4529,N_651,N_231);
nand U4530 (N_4530,N_2486,N_877);
or U4531 (N_4531,N_2168,N_952);
xor U4532 (N_4532,N_276,N_932);
nor U4533 (N_4533,N_1560,N_1887);
xnor U4534 (N_4534,N_2448,N_86);
and U4535 (N_4535,N_1128,N_846);
nand U4536 (N_4536,N_819,N_1533);
or U4537 (N_4537,N_1801,N_2459);
nor U4538 (N_4538,N_1875,N_87);
nor U4539 (N_4539,N_2187,N_2101);
nor U4540 (N_4540,N_83,N_663);
nand U4541 (N_4541,N_1865,N_1638);
and U4542 (N_4542,N_271,N_315);
and U4543 (N_4543,N_1587,N_2405);
nand U4544 (N_4544,N_2437,N_1912);
or U4545 (N_4545,N_2492,N_640);
nand U4546 (N_4546,N_2022,N_422);
nor U4547 (N_4547,N_375,N_1969);
or U4548 (N_4548,N_252,N_1183);
xnor U4549 (N_4549,N_1712,N_2345);
or U4550 (N_4550,N_1612,N_1708);
or U4551 (N_4551,N_885,N_2281);
and U4552 (N_4552,N_2447,N_883);
xor U4553 (N_4553,N_1899,N_262);
xnor U4554 (N_4554,N_1015,N_477);
or U4555 (N_4555,N_836,N_2144);
nor U4556 (N_4556,N_1669,N_2289);
nor U4557 (N_4557,N_1977,N_2321);
nor U4558 (N_4558,N_2243,N_662);
nor U4559 (N_4559,N_2448,N_1041);
and U4560 (N_4560,N_1914,N_704);
nor U4561 (N_4561,N_2029,N_1854);
nand U4562 (N_4562,N_380,N_1451);
nand U4563 (N_4563,N_2225,N_1026);
xnor U4564 (N_4564,N_1231,N_1310);
nor U4565 (N_4565,N_1713,N_1018);
nor U4566 (N_4566,N_1122,N_885);
nor U4567 (N_4567,N_2164,N_1245);
and U4568 (N_4568,N_83,N_1043);
and U4569 (N_4569,N_713,N_2169);
or U4570 (N_4570,N_353,N_1906);
nor U4571 (N_4571,N_1557,N_996);
nand U4572 (N_4572,N_1815,N_2269);
and U4573 (N_4573,N_2458,N_89);
or U4574 (N_4574,N_1859,N_318);
and U4575 (N_4575,N_806,N_386);
xnor U4576 (N_4576,N_1743,N_2364);
xnor U4577 (N_4577,N_1336,N_1179);
or U4578 (N_4578,N_1462,N_1727);
nor U4579 (N_4579,N_971,N_553);
or U4580 (N_4580,N_1825,N_889);
xor U4581 (N_4581,N_2438,N_943);
nor U4582 (N_4582,N_114,N_85);
and U4583 (N_4583,N_2071,N_2079);
nor U4584 (N_4584,N_619,N_1473);
xor U4585 (N_4585,N_2163,N_1977);
xor U4586 (N_4586,N_129,N_802);
xnor U4587 (N_4587,N_715,N_2035);
and U4588 (N_4588,N_86,N_1261);
and U4589 (N_4589,N_1503,N_2304);
nand U4590 (N_4590,N_47,N_1085);
or U4591 (N_4591,N_484,N_2070);
nor U4592 (N_4592,N_2191,N_937);
xnor U4593 (N_4593,N_1963,N_1593);
and U4594 (N_4594,N_1832,N_2267);
nand U4595 (N_4595,N_2279,N_878);
or U4596 (N_4596,N_2411,N_815);
nand U4597 (N_4597,N_1008,N_141);
and U4598 (N_4598,N_852,N_1555);
and U4599 (N_4599,N_507,N_2466);
or U4600 (N_4600,N_1920,N_2376);
nand U4601 (N_4601,N_1966,N_1434);
nand U4602 (N_4602,N_1045,N_1104);
xor U4603 (N_4603,N_464,N_1234);
xor U4604 (N_4604,N_1141,N_779);
nor U4605 (N_4605,N_927,N_2170);
xnor U4606 (N_4606,N_2404,N_1005);
nand U4607 (N_4607,N_1084,N_2102);
and U4608 (N_4608,N_1577,N_1197);
nand U4609 (N_4609,N_804,N_1026);
nand U4610 (N_4610,N_1527,N_1524);
nor U4611 (N_4611,N_1064,N_1441);
and U4612 (N_4612,N_1716,N_597);
or U4613 (N_4613,N_975,N_701);
nor U4614 (N_4614,N_1735,N_1835);
or U4615 (N_4615,N_1552,N_17);
nand U4616 (N_4616,N_2134,N_196);
or U4617 (N_4617,N_1048,N_1063);
or U4618 (N_4618,N_2273,N_1622);
or U4619 (N_4619,N_1280,N_1882);
and U4620 (N_4620,N_666,N_367);
nor U4621 (N_4621,N_1186,N_807);
nor U4622 (N_4622,N_2217,N_448);
xnor U4623 (N_4623,N_476,N_862);
or U4624 (N_4624,N_1181,N_932);
nand U4625 (N_4625,N_2354,N_2181);
and U4626 (N_4626,N_2160,N_111);
xnor U4627 (N_4627,N_232,N_2078);
nor U4628 (N_4628,N_211,N_1427);
nor U4629 (N_4629,N_2301,N_317);
or U4630 (N_4630,N_1576,N_816);
nand U4631 (N_4631,N_655,N_619);
nand U4632 (N_4632,N_1370,N_285);
or U4633 (N_4633,N_1618,N_2352);
nand U4634 (N_4634,N_1058,N_26);
nor U4635 (N_4635,N_1678,N_541);
nand U4636 (N_4636,N_1612,N_2002);
nand U4637 (N_4637,N_719,N_2363);
or U4638 (N_4638,N_640,N_635);
and U4639 (N_4639,N_2301,N_2363);
nor U4640 (N_4640,N_1515,N_1421);
nand U4641 (N_4641,N_1323,N_2166);
or U4642 (N_4642,N_488,N_96);
and U4643 (N_4643,N_854,N_2205);
and U4644 (N_4644,N_1649,N_2037);
nand U4645 (N_4645,N_220,N_2004);
or U4646 (N_4646,N_493,N_2211);
and U4647 (N_4647,N_728,N_2090);
or U4648 (N_4648,N_910,N_200);
xor U4649 (N_4649,N_1790,N_715);
and U4650 (N_4650,N_1146,N_2010);
and U4651 (N_4651,N_900,N_1213);
and U4652 (N_4652,N_2488,N_1727);
and U4653 (N_4653,N_2321,N_357);
nand U4654 (N_4654,N_1428,N_2237);
or U4655 (N_4655,N_345,N_431);
nor U4656 (N_4656,N_215,N_1280);
or U4657 (N_4657,N_1130,N_689);
or U4658 (N_4658,N_1118,N_3);
and U4659 (N_4659,N_1140,N_565);
nor U4660 (N_4660,N_1909,N_11);
or U4661 (N_4661,N_2425,N_1339);
nand U4662 (N_4662,N_1380,N_2254);
or U4663 (N_4663,N_2463,N_1838);
nand U4664 (N_4664,N_2276,N_313);
and U4665 (N_4665,N_1649,N_1512);
and U4666 (N_4666,N_1640,N_2193);
and U4667 (N_4667,N_1864,N_163);
or U4668 (N_4668,N_100,N_2240);
xnor U4669 (N_4669,N_1297,N_1354);
nand U4670 (N_4670,N_606,N_2181);
nor U4671 (N_4671,N_769,N_2282);
or U4672 (N_4672,N_1623,N_1347);
nand U4673 (N_4673,N_2254,N_399);
and U4674 (N_4674,N_1171,N_943);
and U4675 (N_4675,N_1375,N_2209);
nand U4676 (N_4676,N_136,N_2327);
nand U4677 (N_4677,N_686,N_101);
nor U4678 (N_4678,N_2034,N_1365);
and U4679 (N_4679,N_1167,N_659);
nand U4680 (N_4680,N_1567,N_731);
nor U4681 (N_4681,N_589,N_1221);
and U4682 (N_4682,N_2485,N_345);
nor U4683 (N_4683,N_176,N_632);
and U4684 (N_4684,N_1164,N_542);
nand U4685 (N_4685,N_1785,N_1170);
xnor U4686 (N_4686,N_1924,N_100);
or U4687 (N_4687,N_900,N_2121);
nor U4688 (N_4688,N_1304,N_1661);
nor U4689 (N_4689,N_1351,N_2059);
and U4690 (N_4690,N_1923,N_1597);
or U4691 (N_4691,N_2260,N_1050);
or U4692 (N_4692,N_1180,N_1046);
or U4693 (N_4693,N_165,N_2157);
nor U4694 (N_4694,N_358,N_1345);
nor U4695 (N_4695,N_476,N_390);
or U4696 (N_4696,N_1073,N_1267);
nand U4697 (N_4697,N_22,N_1731);
and U4698 (N_4698,N_2425,N_341);
nor U4699 (N_4699,N_1610,N_1386);
and U4700 (N_4700,N_2309,N_1511);
or U4701 (N_4701,N_251,N_1960);
and U4702 (N_4702,N_1178,N_284);
or U4703 (N_4703,N_492,N_1281);
nand U4704 (N_4704,N_2444,N_22);
or U4705 (N_4705,N_1838,N_472);
and U4706 (N_4706,N_1649,N_349);
and U4707 (N_4707,N_1961,N_1333);
and U4708 (N_4708,N_1617,N_1267);
nand U4709 (N_4709,N_1241,N_2460);
xor U4710 (N_4710,N_2304,N_2021);
nor U4711 (N_4711,N_828,N_1946);
or U4712 (N_4712,N_285,N_330);
or U4713 (N_4713,N_2073,N_2465);
nor U4714 (N_4714,N_2222,N_250);
nand U4715 (N_4715,N_1112,N_326);
nand U4716 (N_4716,N_2355,N_502);
and U4717 (N_4717,N_1344,N_2465);
and U4718 (N_4718,N_2219,N_441);
nor U4719 (N_4719,N_332,N_1519);
nor U4720 (N_4720,N_359,N_543);
and U4721 (N_4721,N_1842,N_1293);
xor U4722 (N_4722,N_1579,N_1253);
nor U4723 (N_4723,N_1343,N_912);
nand U4724 (N_4724,N_2162,N_1927);
xor U4725 (N_4725,N_2083,N_1490);
nand U4726 (N_4726,N_1218,N_553);
nor U4727 (N_4727,N_603,N_733);
and U4728 (N_4728,N_1825,N_1536);
and U4729 (N_4729,N_1070,N_40);
and U4730 (N_4730,N_79,N_625);
nand U4731 (N_4731,N_852,N_450);
nand U4732 (N_4732,N_67,N_2342);
nor U4733 (N_4733,N_1717,N_1054);
nor U4734 (N_4734,N_2354,N_490);
or U4735 (N_4735,N_2007,N_500);
and U4736 (N_4736,N_424,N_482);
and U4737 (N_4737,N_1050,N_2438);
and U4738 (N_4738,N_2404,N_727);
and U4739 (N_4739,N_845,N_965);
nand U4740 (N_4740,N_791,N_984);
xnor U4741 (N_4741,N_714,N_2035);
and U4742 (N_4742,N_2232,N_4);
nor U4743 (N_4743,N_2444,N_254);
nand U4744 (N_4744,N_895,N_55);
or U4745 (N_4745,N_1220,N_1397);
nor U4746 (N_4746,N_926,N_5);
nand U4747 (N_4747,N_1780,N_2430);
xnor U4748 (N_4748,N_2478,N_279);
and U4749 (N_4749,N_2096,N_759);
and U4750 (N_4750,N_1999,N_438);
nand U4751 (N_4751,N_833,N_1443);
or U4752 (N_4752,N_1427,N_1635);
nor U4753 (N_4753,N_1129,N_2245);
nor U4754 (N_4754,N_1587,N_2209);
nand U4755 (N_4755,N_821,N_1102);
or U4756 (N_4756,N_574,N_216);
and U4757 (N_4757,N_2462,N_1483);
nand U4758 (N_4758,N_46,N_2375);
and U4759 (N_4759,N_2011,N_827);
nor U4760 (N_4760,N_17,N_1333);
or U4761 (N_4761,N_468,N_1552);
nor U4762 (N_4762,N_2018,N_1888);
nand U4763 (N_4763,N_1769,N_944);
xor U4764 (N_4764,N_2268,N_2399);
or U4765 (N_4765,N_2209,N_24);
or U4766 (N_4766,N_2424,N_2382);
and U4767 (N_4767,N_1415,N_1030);
or U4768 (N_4768,N_1339,N_1426);
nand U4769 (N_4769,N_1650,N_133);
nand U4770 (N_4770,N_561,N_895);
and U4771 (N_4771,N_728,N_1205);
and U4772 (N_4772,N_120,N_2388);
or U4773 (N_4773,N_845,N_613);
and U4774 (N_4774,N_2242,N_1759);
and U4775 (N_4775,N_2005,N_2009);
xnor U4776 (N_4776,N_1385,N_708);
nand U4777 (N_4777,N_954,N_781);
xor U4778 (N_4778,N_2131,N_1867);
and U4779 (N_4779,N_344,N_1637);
or U4780 (N_4780,N_1998,N_1881);
or U4781 (N_4781,N_978,N_1855);
and U4782 (N_4782,N_2099,N_276);
or U4783 (N_4783,N_636,N_2424);
nand U4784 (N_4784,N_1071,N_1327);
or U4785 (N_4785,N_2450,N_202);
xnor U4786 (N_4786,N_511,N_2089);
nand U4787 (N_4787,N_1645,N_1478);
or U4788 (N_4788,N_254,N_1577);
or U4789 (N_4789,N_2201,N_2392);
nand U4790 (N_4790,N_2042,N_141);
nand U4791 (N_4791,N_15,N_2360);
xnor U4792 (N_4792,N_1051,N_1453);
nand U4793 (N_4793,N_1191,N_46);
nand U4794 (N_4794,N_115,N_172);
or U4795 (N_4795,N_667,N_1550);
and U4796 (N_4796,N_928,N_942);
nor U4797 (N_4797,N_634,N_70);
or U4798 (N_4798,N_1226,N_2136);
nand U4799 (N_4799,N_113,N_428);
xor U4800 (N_4800,N_2479,N_1945);
or U4801 (N_4801,N_1544,N_1873);
nand U4802 (N_4802,N_950,N_1814);
and U4803 (N_4803,N_1237,N_742);
or U4804 (N_4804,N_2178,N_820);
and U4805 (N_4805,N_1160,N_1006);
nor U4806 (N_4806,N_1110,N_1045);
nand U4807 (N_4807,N_85,N_1741);
nor U4808 (N_4808,N_26,N_251);
nor U4809 (N_4809,N_1986,N_1321);
and U4810 (N_4810,N_1819,N_672);
nor U4811 (N_4811,N_2402,N_916);
or U4812 (N_4812,N_436,N_2490);
and U4813 (N_4813,N_2148,N_1296);
nand U4814 (N_4814,N_1289,N_1677);
nor U4815 (N_4815,N_1434,N_2474);
nor U4816 (N_4816,N_1799,N_910);
and U4817 (N_4817,N_262,N_1169);
and U4818 (N_4818,N_423,N_660);
nor U4819 (N_4819,N_1138,N_1550);
nor U4820 (N_4820,N_299,N_936);
nand U4821 (N_4821,N_1478,N_786);
nand U4822 (N_4822,N_2284,N_977);
or U4823 (N_4823,N_1844,N_2466);
nand U4824 (N_4824,N_2153,N_173);
or U4825 (N_4825,N_475,N_1248);
nor U4826 (N_4826,N_1733,N_2420);
or U4827 (N_4827,N_620,N_460);
or U4828 (N_4828,N_1336,N_765);
or U4829 (N_4829,N_1428,N_594);
nor U4830 (N_4830,N_1049,N_593);
nor U4831 (N_4831,N_422,N_301);
nor U4832 (N_4832,N_1837,N_2228);
and U4833 (N_4833,N_192,N_2368);
and U4834 (N_4834,N_1829,N_228);
nand U4835 (N_4835,N_1953,N_68);
and U4836 (N_4836,N_1311,N_1127);
nor U4837 (N_4837,N_1962,N_1353);
nor U4838 (N_4838,N_2448,N_686);
nand U4839 (N_4839,N_1263,N_694);
and U4840 (N_4840,N_1768,N_889);
nand U4841 (N_4841,N_2104,N_2397);
and U4842 (N_4842,N_2408,N_209);
xor U4843 (N_4843,N_1584,N_2392);
or U4844 (N_4844,N_886,N_1032);
xor U4845 (N_4845,N_536,N_1022);
xnor U4846 (N_4846,N_2040,N_31);
xnor U4847 (N_4847,N_193,N_413);
and U4848 (N_4848,N_1428,N_1930);
xor U4849 (N_4849,N_101,N_926);
or U4850 (N_4850,N_1606,N_534);
or U4851 (N_4851,N_2276,N_2428);
nor U4852 (N_4852,N_989,N_1739);
xnor U4853 (N_4853,N_721,N_1817);
nor U4854 (N_4854,N_651,N_1461);
nand U4855 (N_4855,N_2048,N_279);
and U4856 (N_4856,N_2215,N_2149);
and U4857 (N_4857,N_1600,N_962);
nand U4858 (N_4858,N_2405,N_2025);
nand U4859 (N_4859,N_2126,N_2187);
xnor U4860 (N_4860,N_788,N_375);
and U4861 (N_4861,N_2426,N_1470);
or U4862 (N_4862,N_1698,N_2413);
and U4863 (N_4863,N_1089,N_1515);
nor U4864 (N_4864,N_1775,N_1026);
or U4865 (N_4865,N_1846,N_2163);
or U4866 (N_4866,N_281,N_1335);
or U4867 (N_4867,N_2097,N_286);
nand U4868 (N_4868,N_1704,N_183);
or U4869 (N_4869,N_44,N_291);
nor U4870 (N_4870,N_1328,N_651);
nor U4871 (N_4871,N_451,N_2022);
or U4872 (N_4872,N_1455,N_1348);
and U4873 (N_4873,N_815,N_62);
nor U4874 (N_4874,N_1269,N_737);
or U4875 (N_4875,N_721,N_716);
nand U4876 (N_4876,N_1833,N_1057);
or U4877 (N_4877,N_509,N_1261);
or U4878 (N_4878,N_2016,N_718);
nor U4879 (N_4879,N_60,N_956);
nand U4880 (N_4880,N_1644,N_909);
xnor U4881 (N_4881,N_1039,N_176);
nand U4882 (N_4882,N_279,N_232);
xnor U4883 (N_4883,N_62,N_618);
and U4884 (N_4884,N_303,N_359);
and U4885 (N_4885,N_2307,N_2249);
nor U4886 (N_4886,N_2271,N_1471);
or U4887 (N_4887,N_2463,N_802);
or U4888 (N_4888,N_339,N_947);
and U4889 (N_4889,N_381,N_869);
nand U4890 (N_4890,N_2056,N_1037);
and U4891 (N_4891,N_1514,N_2094);
or U4892 (N_4892,N_1555,N_1858);
nor U4893 (N_4893,N_97,N_634);
and U4894 (N_4894,N_508,N_2062);
and U4895 (N_4895,N_1596,N_915);
or U4896 (N_4896,N_1250,N_971);
or U4897 (N_4897,N_2249,N_1042);
and U4898 (N_4898,N_150,N_2436);
or U4899 (N_4899,N_0,N_1425);
nand U4900 (N_4900,N_644,N_605);
or U4901 (N_4901,N_1871,N_2200);
nor U4902 (N_4902,N_2059,N_1741);
and U4903 (N_4903,N_1395,N_2342);
xor U4904 (N_4904,N_898,N_636);
and U4905 (N_4905,N_1466,N_2342);
or U4906 (N_4906,N_2218,N_147);
nor U4907 (N_4907,N_2321,N_2014);
and U4908 (N_4908,N_146,N_2235);
and U4909 (N_4909,N_27,N_1420);
nor U4910 (N_4910,N_2297,N_1018);
nor U4911 (N_4911,N_1936,N_1449);
nor U4912 (N_4912,N_1350,N_1145);
nor U4913 (N_4913,N_2085,N_532);
and U4914 (N_4914,N_45,N_1140);
or U4915 (N_4915,N_891,N_1728);
nand U4916 (N_4916,N_895,N_200);
or U4917 (N_4917,N_535,N_734);
nor U4918 (N_4918,N_709,N_1197);
nor U4919 (N_4919,N_681,N_1230);
and U4920 (N_4920,N_1449,N_1300);
and U4921 (N_4921,N_1137,N_2269);
xnor U4922 (N_4922,N_1472,N_1237);
nor U4923 (N_4923,N_1486,N_285);
and U4924 (N_4924,N_1797,N_1750);
xor U4925 (N_4925,N_152,N_2036);
or U4926 (N_4926,N_242,N_1722);
nand U4927 (N_4927,N_1262,N_1151);
xor U4928 (N_4928,N_1941,N_1263);
or U4929 (N_4929,N_2187,N_1587);
or U4930 (N_4930,N_489,N_2217);
nand U4931 (N_4931,N_1558,N_2303);
nor U4932 (N_4932,N_153,N_1681);
or U4933 (N_4933,N_1496,N_2484);
nor U4934 (N_4934,N_41,N_1824);
and U4935 (N_4935,N_2356,N_1586);
and U4936 (N_4936,N_1078,N_1569);
nor U4937 (N_4937,N_1688,N_2119);
or U4938 (N_4938,N_2226,N_1677);
nor U4939 (N_4939,N_2153,N_982);
and U4940 (N_4940,N_1115,N_349);
or U4941 (N_4941,N_1033,N_1449);
nand U4942 (N_4942,N_623,N_1091);
and U4943 (N_4943,N_1325,N_592);
and U4944 (N_4944,N_549,N_1279);
or U4945 (N_4945,N_2016,N_1779);
xnor U4946 (N_4946,N_2262,N_1458);
xnor U4947 (N_4947,N_2014,N_210);
nor U4948 (N_4948,N_2052,N_2411);
xor U4949 (N_4949,N_737,N_354);
nand U4950 (N_4950,N_1725,N_619);
nor U4951 (N_4951,N_777,N_49);
nand U4952 (N_4952,N_1684,N_1133);
nand U4953 (N_4953,N_374,N_1763);
nor U4954 (N_4954,N_2434,N_2492);
nor U4955 (N_4955,N_1763,N_1279);
nand U4956 (N_4956,N_2151,N_1080);
nor U4957 (N_4957,N_406,N_2130);
nand U4958 (N_4958,N_889,N_561);
nor U4959 (N_4959,N_1061,N_1406);
nand U4960 (N_4960,N_2139,N_1383);
or U4961 (N_4961,N_1269,N_2488);
nor U4962 (N_4962,N_1438,N_543);
nand U4963 (N_4963,N_67,N_1102);
xnor U4964 (N_4964,N_2474,N_834);
nor U4965 (N_4965,N_599,N_2172);
xor U4966 (N_4966,N_756,N_1290);
xnor U4967 (N_4967,N_931,N_1266);
nand U4968 (N_4968,N_2116,N_2063);
nand U4969 (N_4969,N_2263,N_218);
xor U4970 (N_4970,N_952,N_1787);
xor U4971 (N_4971,N_2030,N_519);
nor U4972 (N_4972,N_1966,N_1927);
xnor U4973 (N_4973,N_357,N_2312);
or U4974 (N_4974,N_1570,N_1763);
nand U4975 (N_4975,N_542,N_2216);
and U4976 (N_4976,N_703,N_1384);
nor U4977 (N_4977,N_1145,N_299);
and U4978 (N_4978,N_2137,N_2378);
or U4979 (N_4979,N_2263,N_2340);
or U4980 (N_4980,N_2212,N_1856);
nand U4981 (N_4981,N_898,N_286);
or U4982 (N_4982,N_706,N_316);
nor U4983 (N_4983,N_1279,N_1949);
or U4984 (N_4984,N_2462,N_651);
nor U4985 (N_4985,N_665,N_1955);
nand U4986 (N_4986,N_356,N_461);
nor U4987 (N_4987,N_1688,N_1226);
and U4988 (N_4988,N_2119,N_1624);
or U4989 (N_4989,N_675,N_306);
nor U4990 (N_4990,N_2259,N_2205);
nor U4991 (N_4991,N_130,N_2266);
nor U4992 (N_4992,N_680,N_311);
nor U4993 (N_4993,N_1703,N_2287);
or U4994 (N_4994,N_1819,N_2256);
xor U4995 (N_4995,N_1453,N_431);
nand U4996 (N_4996,N_1977,N_1405);
nor U4997 (N_4997,N_1098,N_1878);
or U4998 (N_4998,N_29,N_1465);
nand U4999 (N_4999,N_1859,N_1961);
nand U5000 (N_5000,N_4299,N_2825);
nand U5001 (N_5001,N_4908,N_2605);
xnor U5002 (N_5002,N_2717,N_3555);
or U5003 (N_5003,N_3463,N_2658);
or U5004 (N_5004,N_2673,N_3224);
nand U5005 (N_5005,N_3832,N_4181);
nand U5006 (N_5006,N_4965,N_4117);
nor U5007 (N_5007,N_3856,N_3389);
nor U5008 (N_5008,N_4550,N_3802);
xor U5009 (N_5009,N_2538,N_3203);
and U5010 (N_5010,N_3040,N_3951);
and U5011 (N_5011,N_2970,N_3714);
xnor U5012 (N_5012,N_3523,N_4253);
nand U5013 (N_5013,N_3573,N_2517);
and U5014 (N_5014,N_4764,N_4477);
or U5015 (N_5015,N_2807,N_3993);
or U5016 (N_5016,N_2952,N_3088);
nor U5017 (N_5017,N_4622,N_3287);
or U5018 (N_5018,N_4015,N_3265);
nand U5019 (N_5019,N_4857,N_3569);
or U5020 (N_5020,N_2915,N_2880);
nor U5021 (N_5021,N_4686,N_4656);
and U5022 (N_5022,N_4192,N_3734);
nor U5023 (N_5023,N_4544,N_3613);
or U5024 (N_5024,N_4966,N_4238);
xnor U5025 (N_5025,N_4692,N_2627);
and U5026 (N_5026,N_3860,N_4823);
and U5027 (N_5027,N_3139,N_4964);
nor U5028 (N_5028,N_4900,N_3415);
nor U5029 (N_5029,N_4601,N_4996);
or U5030 (N_5030,N_3290,N_3214);
and U5031 (N_5031,N_3600,N_3949);
and U5032 (N_5032,N_2743,N_3687);
xor U5033 (N_5033,N_3520,N_2847);
nand U5034 (N_5034,N_4731,N_4715);
or U5035 (N_5035,N_3901,N_2913);
or U5036 (N_5036,N_3409,N_4531);
nand U5037 (N_5037,N_3202,N_4241);
nor U5038 (N_5038,N_2729,N_4394);
nand U5039 (N_5039,N_4811,N_3410);
xor U5040 (N_5040,N_4927,N_4779);
and U5041 (N_5041,N_3103,N_3177);
nand U5042 (N_5042,N_4157,N_3731);
nand U5043 (N_5043,N_3748,N_3775);
and U5044 (N_5044,N_3508,N_2587);
nor U5045 (N_5045,N_3417,N_2916);
xnor U5046 (N_5046,N_3208,N_4329);
nor U5047 (N_5047,N_3743,N_2945);
nor U5048 (N_5048,N_3007,N_2867);
nand U5049 (N_5049,N_4075,N_4197);
nand U5050 (N_5050,N_4953,N_3027);
nand U5051 (N_5051,N_3215,N_4828);
and U5052 (N_5052,N_3848,N_2999);
xnor U5053 (N_5053,N_4429,N_2996);
nand U5054 (N_5054,N_2507,N_4146);
or U5055 (N_5055,N_4184,N_4650);
xnor U5056 (N_5056,N_4579,N_2565);
nor U5057 (N_5057,N_4213,N_3703);
and U5058 (N_5058,N_4442,N_2555);
nor U5059 (N_5059,N_3403,N_3124);
and U5060 (N_5060,N_4577,N_3161);
nand U5061 (N_5061,N_4695,N_3312);
or U5062 (N_5062,N_3201,N_4462);
nand U5063 (N_5063,N_4841,N_4364);
xnor U5064 (N_5064,N_2794,N_3930);
and U5065 (N_5065,N_2643,N_2875);
nor U5066 (N_5066,N_3019,N_4406);
or U5067 (N_5067,N_3533,N_3054);
or U5068 (N_5068,N_3707,N_4112);
nand U5069 (N_5069,N_2621,N_3671);
or U5070 (N_5070,N_4278,N_3099);
and U5071 (N_5071,N_3699,N_3246);
nand U5072 (N_5072,N_4138,N_3242);
nor U5073 (N_5073,N_3275,N_4991);
and U5074 (N_5074,N_4711,N_3333);
xnor U5075 (N_5075,N_2854,N_3359);
and U5076 (N_5076,N_3401,N_3777);
nor U5077 (N_5077,N_3763,N_3022);
or U5078 (N_5078,N_4786,N_2509);
and U5079 (N_5079,N_2602,N_4418);
nor U5080 (N_5080,N_4600,N_4613);
and U5081 (N_5081,N_3596,N_2693);
nor U5082 (N_5082,N_4982,N_3116);
or U5083 (N_5083,N_3504,N_3990);
xor U5084 (N_5084,N_3962,N_3293);
nand U5085 (N_5085,N_4549,N_2628);
nand U5086 (N_5086,N_4688,N_3388);
and U5087 (N_5087,N_4268,N_2540);
xor U5088 (N_5088,N_2888,N_3123);
or U5089 (N_5089,N_2561,N_3324);
nor U5090 (N_5090,N_3711,N_3952);
or U5091 (N_5091,N_3840,N_3647);
nor U5092 (N_5092,N_4759,N_3467);
and U5093 (N_5093,N_4926,N_3446);
nor U5094 (N_5094,N_2823,N_3051);
or U5095 (N_5095,N_4814,N_4645);
nor U5096 (N_5096,N_3392,N_3753);
or U5097 (N_5097,N_4553,N_3279);
nor U5098 (N_5098,N_4099,N_3634);
or U5099 (N_5099,N_2819,N_2719);
or U5100 (N_5100,N_2747,N_4317);
or U5101 (N_5101,N_4773,N_3209);
or U5102 (N_5102,N_4451,N_4551);
nor U5103 (N_5103,N_4165,N_3579);
and U5104 (N_5104,N_4744,N_4678);
xor U5105 (N_5105,N_3999,N_2938);
nand U5106 (N_5106,N_4776,N_3673);
nor U5107 (N_5107,N_4237,N_3805);
or U5108 (N_5108,N_4658,N_2813);
nand U5109 (N_5109,N_4279,N_3193);
or U5110 (N_5110,N_2615,N_4320);
or U5111 (N_5111,N_4855,N_2535);
xor U5112 (N_5112,N_4296,N_3919);
nand U5113 (N_5113,N_2626,N_3241);
or U5114 (N_5114,N_3571,N_3631);
and U5115 (N_5115,N_3567,N_4851);
nor U5116 (N_5116,N_3618,N_3000);
nand U5117 (N_5117,N_3319,N_3747);
and U5118 (N_5118,N_4662,N_4272);
and U5119 (N_5119,N_3517,N_4460);
nand U5120 (N_5120,N_3853,N_4143);
nand U5121 (N_5121,N_4830,N_3922);
or U5122 (N_5122,N_4298,N_3510);
nand U5123 (N_5123,N_4382,N_3666);
nand U5124 (N_5124,N_3781,N_4103);
or U5125 (N_5125,N_4751,N_4447);
and U5126 (N_5126,N_4998,N_3348);
nand U5127 (N_5127,N_3304,N_4159);
and U5128 (N_5128,N_4772,N_3439);
xor U5129 (N_5129,N_4990,N_3150);
or U5130 (N_5130,N_4264,N_2769);
nand U5131 (N_5131,N_2527,N_2775);
nor U5132 (N_5132,N_4957,N_4979);
nor U5133 (N_5133,N_2560,N_4370);
nand U5134 (N_5134,N_4952,N_3329);
and U5135 (N_5135,N_2849,N_3334);
nand U5136 (N_5136,N_3238,N_4540);
xnor U5137 (N_5137,N_3768,N_4217);
or U5138 (N_5138,N_4829,N_3250);
nor U5139 (N_5139,N_4351,N_4417);
nor U5140 (N_5140,N_3710,N_3119);
or U5141 (N_5141,N_4604,N_3609);
or U5142 (N_5142,N_4737,N_4621);
and U5143 (N_5143,N_2618,N_4722);
and U5144 (N_5144,N_4959,N_3969);
or U5145 (N_5145,N_3746,N_4535);
and U5146 (N_5146,N_3806,N_4361);
nor U5147 (N_5147,N_4465,N_4562);
nor U5148 (N_5148,N_2539,N_3098);
nand U5149 (N_5149,N_4457,N_3542);
and U5150 (N_5150,N_3918,N_3872);
and U5151 (N_5151,N_2569,N_3190);
nand U5152 (N_5152,N_3667,N_3495);
nor U5153 (N_5153,N_3380,N_2537);
nand U5154 (N_5154,N_4865,N_4387);
nor U5155 (N_5155,N_2832,N_4897);
nand U5156 (N_5156,N_2589,N_3948);
and U5157 (N_5157,N_4022,N_3128);
nand U5158 (N_5158,N_3036,N_3063);
xor U5159 (N_5159,N_3016,N_3411);
nand U5160 (N_5160,N_3166,N_4592);
nor U5161 (N_5161,N_3791,N_4742);
nor U5162 (N_5162,N_3692,N_4520);
nor U5163 (N_5163,N_3301,N_2787);
nand U5164 (N_5164,N_3732,N_3065);
nand U5165 (N_5165,N_3736,N_3628);
nor U5166 (N_5166,N_3331,N_4790);
or U5167 (N_5167,N_2919,N_3669);
and U5168 (N_5168,N_4794,N_3965);
and U5169 (N_5169,N_4256,N_3986);
or U5170 (N_5170,N_2637,N_3082);
xnor U5171 (N_5171,N_4974,N_4791);
nand U5172 (N_5172,N_3725,N_4120);
nand U5173 (N_5173,N_4205,N_2646);
or U5174 (N_5174,N_3658,N_4866);
and U5175 (N_5175,N_4559,N_4992);
nand U5176 (N_5176,N_4190,N_3869);
nand U5177 (N_5177,N_3830,N_4511);
and U5178 (N_5178,N_4523,N_4726);
nand U5179 (N_5179,N_4856,N_3838);
or U5180 (N_5180,N_3767,N_4142);
nand U5181 (N_5181,N_3844,N_4978);
xnor U5182 (N_5182,N_3055,N_3408);
nand U5183 (N_5183,N_3820,N_4440);
and U5184 (N_5184,N_3044,N_2607);
nor U5185 (N_5185,N_2511,N_3390);
xnor U5186 (N_5186,N_3010,N_2796);
nand U5187 (N_5187,N_3985,N_2765);
or U5188 (N_5188,N_3247,N_4066);
or U5189 (N_5189,N_2632,N_4479);
nand U5190 (N_5190,N_3213,N_3366);
and U5191 (N_5191,N_3911,N_3770);
or U5192 (N_5192,N_4193,N_3852);
and U5193 (N_5193,N_3896,N_4188);
or U5194 (N_5194,N_4698,N_2963);
nand U5195 (N_5195,N_4603,N_3189);
nor U5196 (N_5196,N_3198,N_3701);
nor U5197 (N_5197,N_4221,N_3910);
or U5198 (N_5198,N_3636,N_2922);
nor U5199 (N_5199,N_4547,N_4774);
nor U5200 (N_5200,N_3737,N_3079);
xor U5201 (N_5201,N_4100,N_4259);
xor U5202 (N_5202,N_4132,N_3525);
and U5203 (N_5203,N_2649,N_2793);
nor U5204 (N_5204,N_3998,N_3894);
xnor U5205 (N_5205,N_3369,N_3210);
nand U5206 (N_5206,N_4290,N_4407);
or U5207 (N_5207,N_3811,N_4231);
nand U5208 (N_5208,N_3109,N_2550);
and U5209 (N_5209,N_2519,N_3788);
nor U5210 (N_5210,N_2672,N_2834);
xor U5211 (N_5211,N_2756,N_3130);
or U5212 (N_5212,N_3289,N_3527);
and U5213 (N_5213,N_3738,N_2824);
or U5214 (N_5214,N_3170,N_2840);
nor U5215 (N_5215,N_4064,N_2577);
and U5216 (N_5216,N_2795,N_4166);
and U5217 (N_5217,N_4212,N_4567);
nand U5218 (N_5218,N_3438,N_3477);
xor U5219 (N_5219,N_4044,N_4373);
xor U5220 (N_5220,N_4614,N_2506);
and U5221 (N_5221,N_3457,N_3778);
nand U5222 (N_5222,N_3378,N_4476);
or U5223 (N_5223,N_3705,N_2651);
and U5224 (N_5224,N_2966,N_3807);
and U5225 (N_5225,N_3167,N_2781);
nor U5226 (N_5226,N_2644,N_4246);
nand U5227 (N_5227,N_4162,N_2500);
xor U5228 (N_5228,N_3184,N_4057);
or U5229 (N_5229,N_3306,N_4254);
and U5230 (N_5230,N_3696,N_4867);
nor U5231 (N_5231,N_4420,N_3970);
nand U5232 (N_5232,N_3263,N_3858);
and U5233 (N_5233,N_3940,N_3288);
and U5234 (N_5234,N_3133,N_4527);
xnor U5235 (N_5235,N_4145,N_3352);
nand U5236 (N_5236,N_2901,N_2726);
nand U5237 (N_5237,N_3792,N_4310);
xnor U5238 (N_5238,N_3994,N_3062);
or U5239 (N_5239,N_4948,N_4795);
xor U5240 (N_5240,N_3988,N_3323);
or U5241 (N_5241,N_4110,N_3262);
and U5242 (N_5242,N_4950,N_3783);
nor U5243 (N_5243,N_4338,N_3914);
nor U5244 (N_5244,N_4029,N_4854);
or U5245 (N_5245,N_4243,N_2751);
nor U5246 (N_5246,N_3982,N_4788);
nor U5247 (N_5247,N_3078,N_3363);
and U5248 (N_5248,N_2689,N_2883);
nor U5249 (N_5249,N_2778,N_2549);
xnor U5250 (N_5250,N_3780,N_2653);
or U5251 (N_5251,N_4904,N_2805);
nor U5252 (N_5252,N_2905,N_3344);
xor U5253 (N_5253,N_4881,N_2714);
nand U5254 (N_5254,N_3897,N_4833);
xnor U5255 (N_5255,N_3440,N_3039);
or U5256 (N_5256,N_3585,N_4609);
nand U5257 (N_5257,N_2852,N_4532);
or U5258 (N_5258,N_4853,N_4326);
and U5259 (N_5259,N_3235,N_2924);
and U5260 (N_5260,N_3456,N_4089);
and U5261 (N_5261,N_3603,N_3419);
nor U5262 (N_5262,N_2856,N_4670);
xor U5263 (N_5263,N_3772,N_3393);
nor U5264 (N_5264,N_4422,N_3566);
or U5265 (N_5265,N_4409,N_3338);
or U5266 (N_5266,N_4739,N_2655);
nor U5267 (N_5267,N_4333,N_3434);
and U5268 (N_5268,N_3169,N_3505);
xor U5269 (N_5269,N_3524,N_3248);
nand U5270 (N_5270,N_4566,N_3207);
nand U5271 (N_5271,N_3679,N_3612);
nand U5272 (N_5272,N_3361,N_3833);
nand U5273 (N_5273,N_4706,N_4104);
or U5274 (N_5274,N_3360,N_4675);
and U5275 (N_5275,N_3158,N_3286);
and U5276 (N_5276,N_3642,N_4195);
xor U5277 (N_5277,N_4458,N_4247);
or U5278 (N_5278,N_4931,N_3905);
nand U5279 (N_5279,N_2700,N_3164);
and U5280 (N_5280,N_3113,N_2923);
xnor U5281 (N_5281,N_4514,N_4710);
nand U5282 (N_5282,N_4702,N_3989);
and U5283 (N_5283,N_3580,N_2745);
nand U5284 (N_5284,N_4886,N_3817);
nor U5285 (N_5285,N_3118,N_4993);
and U5286 (N_5286,N_2884,N_4892);
xnor U5287 (N_5287,N_4199,N_4727);
nand U5288 (N_5288,N_2701,N_3066);
and U5289 (N_5289,N_2675,N_3627);
nand U5290 (N_5290,N_3583,N_3387);
or U5291 (N_5291,N_3377,N_4176);
and U5292 (N_5292,N_4825,N_3857);
and U5293 (N_5293,N_4115,N_3451);
nor U5294 (N_5294,N_4280,N_2936);
nor U5295 (N_5295,N_4501,N_4983);
and U5296 (N_5296,N_3195,N_4515);
xor U5297 (N_5297,N_4081,N_3625);
xnor U5298 (N_5298,N_3244,N_3528);
nand U5299 (N_5299,N_4034,N_3966);
nand U5300 (N_5300,N_2810,N_4425);
and U5301 (N_5301,N_2677,N_2528);
or U5302 (N_5302,N_3511,N_3796);
nor U5303 (N_5303,N_3432,N_4718);
and U5304 (N_5304,N_4464,N_4906);
nor U5305 (N_5305,N_2845,N_3095);
xnor U5306 (N_5306,N_3336,N_3887);
nand U5307 (N_5307,N_4557,N_3519);
xor U5308 (N_5308,N_2815,N_3509);
or U5309 (N_5309,N_4879,N_3633);
and U5310 (N_5310,N_3353,N_3216);
or U5311 (N_5311,N_3947,N_3006);
nand U5312 (N_5312,N_2948,N_4250);
xor U5313 (N_5313,N_3229,N_4976);
or U5314 (N_5314,N_3154,N_4385);
nand U5315 (N_5315,N_4219,N_3159);
nor U5316 (N_5316,N_3452,N_4587);
nor U5317 (N_5317,N_3882,N_4914);
and U5318 (N_5318,N_4466,N_2788);
nand U5319 (N_5319,N_4118,N_3649);
or U5320 (N_5320,N_3971,N_3426);
or U5321 (N_5321,N_4070,N_4661);
nor U5322 (N_5322,N_4173,N_3089);
or U5323 (N_5323,N_3147,N_4270);
or U5324 (N_5324,N_3535,N_4378);
and U5325 (N_5325,N_4597,N_3662);
nor U5326 (N_5326,N_2648,N_2954);
and U5327 (N_5327,N_3429,N_4659);
or U5328 (N_5328,N_4139,N_3141);
or U5329 (N_5329,N_3597,N_3757);
or U5330 (N_5330,N_3871,N_2908);
and U5331 (N_5331,N_4301,N_3266);
or U5332 (N_5332,N_4043,N_4304);
xnor U5333 (N_5333,N_2839,N_4655);
and U5334 (N_5334,N_3604,N_4505);
and U5335 (N_5335,N_4619,N_4668);
nor U5336 (N_5336,N_4168,N_3582);
and U5337 (N_5337,N_3398,N_3367);
and U5338 (N_5338,N_3956,N_3764);
or U5339 (N_5339,N_3050,N_3494);
or U5340 (N_5340,N_3812,N_3889);
nand U5341 (N_5341,N_4454,N_4723);
nand U5342 (N_5342,N_4391,N_2721);
nand U5343 (N_5343,N_4743,N_4623);
nor U5344 (N_5344,N_3346,N_4463);
nor U5345 (N_5345,N_2898,N_3760);
or U5346 (N_5346,N_3385,N_4348);
nor U5347 (N_5347,N_4988,N_3131);
and U5348 (N_5348,N_3491,N_4970);
or U5349 (N_5349,N_4494,N_3482);
nor U5350 (N_5350,N_3974,N_2592);
and U5351 (N_5351,N_3249,N_3194);
xor U5352 (N_5352,N_3181,N_4491);
nand U5353 (N_5353,N_2711,N_4151);
and U5354 (N_5354,N_2516,N_4318);
nor U5355 (N_5355,N_4666,N_4654);
or U5356 (N_5356,N_4339,N_3162);
nand U5357 (N_5357,N_3120,N_3867);
and U5358 (N_5358,N_3005,N_2917);
nor U5359 (N_5359,N_3358,N_4092);
nor U5360 (N_5360,N_3521,N_4350);
nor U5361 (N_5361,N_4905,N_4560);
or U5362 (N_5362,N_4677,N_3942);
nor U5363 (N_5363,N_3761,N_4288);
nand U5364 (N_5364,N_2568,N_4080);
nand U5365 (N_5365,N_4049,N_3593);
or U5366 (N_5366,N_2989,N_4431);
nor U5367 (N_5367,N_4397,N_2513);
and U5368 (N_5368,N_4332,N_3294);
nor U5369 (N_5369,N_3012,N_3908);
or U5370 (N_5370,N_3218,N_3906);
nand U5371 (N_5371,N_4760,N_3675);
or U5372 (N_5372,N_4660,N_3719);
or U5373 (N_5373,N_3332,N_4369);
nand U5374 (N_5374,N_4203,N_2613);
or U5375 (N_5375,N_2777,N_3471);
and U5376 (N_5376,N_2541,N_3616);
xnor U5377 (N_5377,N_4876,N_3973);
nand U5378 (N_5378,N_2720,N_3048);
xnor U5379 (N_5379,N_4487,N_4191);
and U5380 (N_5380,N_3093,N_2877);
nor U5381 (N_5381,N_3588,N_2739);
nor U5382 (N_5382,N_4512,N_2891);
or U5383 (N_5383,N_3728,N_3898);
nand U5384 (N_5384,N_4712,N_2993);
and U5385 (N_5385,N_2635,N_3236);
nor U5386 (N_5386,N_4210,N_4933);
and U5387 (N_5387,N_2508,N_4360);
and U5388 (N_5388,N_4135,N_2725);
nand U5389 (N_5389,N_3926,N_3543);
nand U5390 (N_5390,N_3683,N_3056);
nor U5391 (N_5391,N_3067,N_4522);
and U5392 (N_5392,N_4632,N_2681);
xnor U5393 (N_5393,N_4482,N_4311);
nand U5394 (N_5394,N_2960,N_3694);
and U5395 (N_5395,N_3977,N_4229);
xor U5396 (N_5396,N_3232,N_3292);
and U5397 (N_5397,N_4664,N_4025);
xnor U5398 (N_5398,N_3061,N_3976);
nand U5399 (N_5399,N_3371,N_4365);
and U5400 (N_5400,N_3615,N_2683);
and U5401 (N_5401,N_4041,N_3379);
or U5402 (N_5402,N_2780,N_3859);
nand U5403 (N_5403,N_3485,N_3670);
nand U5404 (N_5404,N_3002,N_4438);
nor U5405 (N_5405,N_3723,N_4835);
nor U5406 (N_5406,N_3476,N_4273);
nand U5407 (N_5407,N_2616,N_4810);
and U5408 (N_5408,N_4345,N_2552);
or U5409 (N_5409,N_4721,N_4123);
and U5410 (N_5410,N_4050,N_4060);
nand U5411 (N_5411,N_3572,N_4058);
nand U5412 (N_5412,N_4745,N_3621);
nand U5413 (N_5413,N_2978,N_3865);
nand U5414 (N_5414,N_2744,N_2737);
or U5415 (N_5415,N_2962,N_4691);
nand U5416 (N_5416,N_3021,N_3255);
and U5417 (N_5417,N_4344,N_2665);
nor U5418 (N_5418,N_4647,N_4975);
and U5419 (N_5419,N_3839,N_3529);
xor U5420 (N_5420,N_3690,N_3008);
nor U5421 (N_5421,N_3325,N_2790);
xnor U5422 (N_5422,N_2678,N_3726);
and U5423 (N_5423,N_4673,N_2973);
or U5424 (N_5424,N_2782,N_3256);
nor U5425 (N_5425,N_3739,N_3205);
or U5426 (N_5426,N_4574,N_3818);
and U5427 (N_5427,N_3316,N_3716);
and U5428 (N_5428,N_4873,N_2706);
and U5429 (N_5429,N_4985,N_3490);
xor U5430 (N_5430,N_4230,N_3094);
nand U5431 (N_5431,N_3327,N_3253);
and U5432 (N_5432,N_4021,N_4657);
nor U5433 (N_5433,N_4082,N_3225);
nand U5434 (N_5434,N_4469,N_4672);
or U5435 (N_5435,N_4258,N_2520);
xor U5436 (N_5436,N_2708,N_4428);
and U5437 (N_5437,N_3272,N_3240);
nand U5438 (N_5438,N_3427,N_4942);
nor U5439 (N_5439,N_4196,N_4434);
nor U5440 (N_5440,N_4837,N_3594);
nand U5441 (N_5441,N_3500,N_4340);
nand U5442 (N_5442,N_4822,N_4618);
nand U5443 (N_5443,N_3657,N_4068);
or U5444 (N_5444,N_4643,N_4831);
or U5445 (N_5445,N_4214,N_3721);
and U5446 (N_5446,N_3171,N_4433);
xor U5447 (N_5447,N_4870,N_3557);
nor U5448 (N_5448,N_3766,N_3168);
nor U5449 (N_5449,N_3932,N_4697);
nor U5450 (N_5450,N_2902,N_4306);
nand U5451 (N_5451,N_4252,N_3605);
xor U5452 (N_5452,N_3972,N_4898);
or U5453 (N_5453,N_3587,N_4154);
xnor U5454 (N_5454,N_4938,N_3834);
nor U5455 (N_5455,N_4977,N_2588);
or U5456 (N_5456,N_3486,N_3963);
and U5457 (N_5457,N_3186,N_4999);
nand U5458 (N_5458,N_3749,N_3590);
and U5459 (N_5459,N_4808,N_3058);
and U5460 (N_5460,N_2910,N_4228);
or U5461 (N_5461,N_4152,N_3619);
or U5462 (N_5462,N_4371,N_2980);
xnor U5463 (N_5463,N_3730,N_4910);
xor U5464 (N_5464,N_4248,N_3042);
and U5465 (N_5465,N_4750,N_3473);
nand U5466 (N_5466,N_3904,N_2596);
nor U5467 (N_5467,N_3416,N_4002);
or U5468 (N_5468,N_2601,N_2502);
or U5469 (N_5469,N_4995,N_3400);
nor U5470 (N_5470,N_4072,N_4561);
or U5471 (N_5471,N_4114,N_3462);
or U5472 (N_5472,N_4923,N_3268);
xnor U5473 (N_5473,N_4335,N_2702);
and U5474 (N_5474,N_2571,N_3717);
nor U5475 (N_5475,N_2685,N_2764);
xor U5476 (N_5476,N_3992,N_4011);
nor U5477 (N_5477,N_4669,N_4374);
nor U5478 (N_5478,N_2863,N_4861);
nand U5479 (N_5479,N_3498,N_3843);
or U5480 (N_5480,N_4590,N_2946);
nand U5481 (N_5481,N_4202,N_4717);
or U5482 (N_5482,N_3004,N_4519);
nor U5483 (N_5483,N_2551,N_2894);
nor U5484 (N_5484,N_2779,N_3009);
and U5485 (N_5485,N_2734,N_4917);
or U5486 (N_5486,N_3688,N_3142);
nand U5487 (N_5487,N_2570,N_3444);
and U5488 (N_5488,N_3046,N_3630);
xor U5489 (N_5489,N_2887,N_4134);
xnor U5490 (N_5490,N_4947,N_4144);
or U5491 (N_5491,N_2827,N_3362);
or U5492 (N_5492,N_4426,N_4951);
nor U5493 (N_5493,N_4179,N_4073);
and U5494 (N_5494,N_3484,N_4328);
and U5495 (N_5495,N_4775,N_4033);
nand U5496 (N_5496,N_4172,N_3793);
nand U5497 (N_5497,N_4652,N_4239);
or U5498 (N_5498,N_4972,N_3623);
and U5499 (N_5499,N_3041,N_4513);
or U5500 (N_5500,N_3862,N_2799);
xor U5501 (N_5501,N_2650,N_4724);
and U5502 (N_5502,N_4899,N_3650);
nor U5503 (N_5503,N_4275,N_3559);
and U5504 (N_5504,N_3043,N_4872);
nor U5505 (N_5505,N_3396,N_4492);
nand U5506 (N_5506,N_4017,N_3134);
xor U5507 (N_5507,N_3206,N_2770);
xnor U5508 (N_5508,N_4411,N_3191);
and U5509 (N_5509,N_4800,N_2523);
nand U5510 (N_5510,N_3877,N_2546);
nor U5511 (N_5511,N_3789,N_2738);
nand U5512 (N_5512,N_3307,N_4709);
nand U5513 (N_5513,N_4481,N_3556);
xnor U5514 (N_5514,N_4485,N_3996);
nor U5515 (N_5515,N_4665,N_3176);
nand U5516 (N_5516,N_3469,N_2688);
and U5517 (N_5517,N_3735,N_3132);
nand U5518 (N_5518,N_4637,N_2639);
nand U5519 (N_5519,N_4486,N_2971);
nand U5520 (N_5520,N_3611,N_3337);
nand U5521 (N_5521,N_3536,N_4761);
nand U5522 (N_5522,N_4839,N_2526);
nand U5523 (N_5523,N_3665,N_3277);
or U5524 (N_5524,N_2543,N_4671);
or U5525 (N_5525,N_2547,N_2821);
nor U5526 (N_5526,N_2789,N_3945);
and U5527 (N_5527,N_2704,N_2668);
nand U5528 (N_5528,N_4546,N_4013);
xor U5529 (N_5529,N_3180,N_3878);
nor U5530 (N_5530,N_2728,N_4708);
and U5531 (N_5531,N_4321,N_4424);
xor U5532 (N_5532,N_4612,N_4455);
nand U5533 (N_5533,N_2878,N_3893);
and U5534 (N_5534,N_4018,N_3921);
nand U5535 (N_5535,N_4215,N_4322);
nand U5536 (N_5536,N_3020,N_4000);
and U5537 (N_5537,N_4740,N_4934);
nor U5538 (N_5538,N_2732,N_4539);
nor U5539 (N_5539,N_3544,N_4785);
and U5540 (N_5540,N_4380,N_3243);
and U5541 (N_5541,N_3470,N_4504);
nor U5542 (N_5542,N_3819,N_3870);
nand U5543 (N_5543,N_2975,N_3801);
or U5544 (N_5544,N_4255,N_3879);
or U5545 (N_5545,N_4768,N_2865);
nand U5546 (N_5546,N_3129,N_4834);
nor U5547 (N_5547,N_4012,N_3825);
or U5548 (N_5548,N_2949,N_3632);
or U5549 (N_5549,N_4140,N_2670);
nand U5550 (N_5550,N_4038,N_2760);
and U5551 (N_5551,N_3863,N_4909);
nor U5552 (N_5552,N_3326,N_4626);
xnor U5553 (N_5553,N_4470,N_3617);
nand U5554 (N_5554,N_3718,N_4850);
nor U5555 (N_5555,N_4780,N_4888);
and U5556 (N_5556,N_4267,N_2992);
and U5557 (N_5557,N_4689,N_4292);
nor U5558 (N_5558,N_4687,N_3328);
nand U5559 (N_5559,N_4251,N_4679);
or U5560 (N_5560,N_4836,N_4606);
nand U5561 (N_5561,N_2935,N_2792);
and U5562 (N_5562,N_2850,N_2881);
and U5563 (N_5563,N_4128,N_3924);
or U5564 (N_5564,N_3798,N_4085);
nand U5565 (N_5565,N_4071,N_3121);
xor U5566 (N_5566,N_2741,N_3927);
nor U5567 (N_5567,N_3888,N_4402);
xor U5568 (N_5568,N_3883,N_4575);
xnor U5569 (N_5569,N_3584,N_2713);
nand U5570 (N_5570,N_4962,N_3311);
nor U5571 (N_5571,N_4967,N_4094);
nand U5572 (N_5572,N_4323,N_3755);
and U5573 (N_5573,N_3297,N_3693);
xnor U5574 (N_5574,N_4175,N_3784);
nand U5575 (N_5575,N_3727,N_4838);
or U5576 (N_5576,N_4555,N_2624);
xor U5577 (N_5577,N_3345,N_4445);
xor U5578 (N_5578,N_3873,N_4300);
or U5579 (N_5579,N_3744,N_2956);
nand U5580 (N_5580,N_2666,N_4432);
or U5581 (N_5581,N_3321,N_3855);
nor U5582 (N_5582,N_2955,N_3514);
xnor U5583 (N_5583,N_4189,N_3917);
or U5584 (N_5584,N_4436,N_4459);
nand U5585 (N_5585,N_3943,N_2876);
nor U5586 (N_5586,N_4233,N_4583);
nor U5587 (N_5587,N_3779,N_3383);
or U5588 (N_5588,N_3916,N_4046);
or U5589 (N_5589,N_4807,N_4206);
nand U5590 (N_5590,N_4696,N_2967);
nand U5591 (N_5591,N_4912,N_4194);
and U5592 (N_5592,N_3902,N_3516);
or U5593 (N_5593,N_4083,N_2691);
or U5594 (N_5594,N_3866,N_4334);
and U5595 (N_5595,N_4884,N_3281);
or U5596 (N_5596,N_3231,N_2994);
or U5597 (N_5597,N_3091,N_3836);
nand U5598 (N_5598,N_4793,N_3537);
or U5599 (N_5599,N_2724,N_4804);
and U5600 (N_5600,N_4449,N_2858);
or U5601 (N_5601,N_2581,N_4153);
or U5602 (N_5602,N_4285,N_3081);
nand U5603 (N_5603,N_3175,N_3173);
nor U5604 (N_5604,N_3995,N_4414);
xnor U5605 (N_5605,N_2654,N_3964);
nor U5606 (N_5606,N_4101,N_4542);
nor U5607 (N_5607,N_4316,N_3546);
xor U5608 (N_5608,N_4367,N_4591);
xor U5609 (N_5609,N_3715,N_4016);
nor U5610 (N_5610,N_4342,N_4676);
xnor U5611 (N_5611,N_4565,N_3720);
nor U5612 (N_5612,N_2947,N_3259);
or U5613 (N_5613,N_2939,N_3083);
nor U5614 (N_5614,N_2761,N_4939);
or U5615 (N_5615,N_3394,N_4960);
nor U5616 (N_5616,N_2951,N_2515);
xor U5617 (N_5617,N_2522,N_4131);
xnor U5618 (N_5618,N_3936,N_4007);
and U5619 (N_5619,N_3531,N_3001);
nor U5620 (N_5620,N_2835,N_3540);
xor U5621 (N_5621,N_3765,N_2647);
nand U5622 (N_5622,N_4693,N_3641);
nor U5623 (N_5623,N_3450,N_4032);
or U5624 (N_5624,N_3502,N_3220);
nand U5625 (N_5625,N_3137,N_4398);
and U5626 (N_5626,N_3421,N_4536);
nor U5627 (N_5627,N_4630,N_4052);
or U5628 (N_5628,N_4663,N_4218);
or U5629 (N_5629,N_2715,N_3179);
or U5630 (N_5630,N_4062,N_2680);
nor U5631 (N_5631,N_4891,N_2785);
or U5632 (N_5632,N_3100,N_4852);
nor U5633 (N_5633,N_3032,N_3308);
and U5634 (N_5634,N_3145,N_3550);
nand U5635 (N_5635,N_4849,N_2591);
or U5636 (N_5636,N_4694,N_3909);
or U5637 (N_5637,N_3541,N_2553);
or U5638 (N_5638,N_4922,N_4347);
and U5639 (N_5639,N_4984,N_4356);
nand U5640 (N_5640,N_2829,N_3481);
xor U5641 (N_5641,N_3709,N_2853);
nor U5642 (N_5642,N_4918,N_3441);
xor U5643 (N_5643,N_4524,N_4869);
nor U5644 (N_5644,N_2752,N_3375);
or U5645 (N_5645,N_4916,N_3414);
nand U5646 (N_5646,N_4421,N_3322);
or U5647 (N_5647,N_2742,N_3545);
and U5648 (N_5648,N_2758,N_3017);
nor U5649 (N_5649,N_4077,N_3903);
xnor U5650 (N_5650,N_4207,N_3899);
nand U5651 (N_5651,N_2842,N_3851);
or U5652 (N_5652,N_3102,N_3700);
nand U5653 (N_5653,N_3565,N_4392);
nand U5654 (N_5654,N_4517,N_4249);
xor U5655 (N_5655,N_2548,N_4895);
and U5656 (N_5656,N_4483,N_3733);
nor U5657 (N_5657,N_4667,N_2892);
nor U5658 (N_5658,N_2903,N_4681);
nand U5659 (N_5659,N_4593,N_2929);
nand U5660 (N_5660,N_4354,N_4832);
and U5661 (N_5661,N_3923,N_2659);
and U5662 (N_5662,N_4404,N_3111);
nor U5663 (N_5663,N_4815,N_4295);
xor U5664 (N_5664,N_2617,N_4343);
nand U5665 (N_5665,N_4167,N_3875);
and U5666 (N_5666,N_4889,N_4627);
xnor U5667 (N_5667,N_4170,N_4161);
nor U5668 (N_5668,N_4375,N_3660);
xor U5669 (N_5669,N_2524,N_4732);
or U5670 (N_5670,N_4042,N_3372);
nand U5671 (N_5671,N_2988,N_4498);
xor U5672 (N_5672,N_4610,N_4704);
and U5673 (N_5673,N_2501,N_4578);
nor U5674 (N_5674,N_3607,N_4816);
nor U5675 (N_5675,N_3313,N_3424);
nor U5676 (N_5676,N_2690,N_3752);
nand U5677 (N_5677,N_4784,N_3568);
xor U5678 (N_5678,N_3357,N_3648);
or U5679 (N_5679,N_4163,N_2566);
or U5680 (N_5680,N_2636,N_2671);
nand U5681 (N_5681,N_3601,N_4054);
nand U5682 (N_5682,N_4389,N_3939);
nand U5683 (N_5683,N_2995,N_3075);
nand U5684 (N_5684,N_3629,N_3644);
and U5685 (N_5685,N_3551,N_3589);
xor U5686 (N_5686,N_2921,N_4448);
nand U5687 (N_5687,N_2563,N_3487);
and U5688 (N_5688,N_3447,N_3257);
nor U5689 (N_5689,N_3234,N_4882);
or U5690 (N_5690,N_4968,N_4518);
nand U5691 (N_5691,N_4955,N_3185);
or U5692 (N_5692,N_2564,N_4758);
and U5693 (N_5693,N_3845,N_3474);
nor U5694 (N_5694,N_3199,N_4051);
and U5695 (N_5695,N_3958,N_2518);
nand U5696 (N_5696,N_3049,N_3143);
nand U5697 (N_5697,N_3599,N_3900);
or U5698 (N_5698,N_3413,N_3740);
nand U5699 (N_5699,N_3298,N_3156);
and U5700 (N_5700,N_4569,N_3810);
or U5701 (N_5701,N_2869,N_4031);
nor U5702 (N_5702,N_3771,N_4509);
nor U5703 (N_5703,N_2959,N_2558);
or U5704 (N_5704,N_2979,N_3428);
nand U5705 (N_5705,N_3983,N_3854);
nand U5706 (N_5706,N_4439,N_3881);
nand U5707 (N_5707,N_4746,N_3373);
nand U5708 (N_5708,N_4495,N_4585);
or U5709 (N_5709,N_2556,N_2941);
or U5710 (N_5710,N_2983,N_2608);
nor U5711 (N_5711,N_4631,N_3892);
nor U5712 (N_5712,N_3957,N_3769);
nor U5713 (N_5713,N_4286,N_3880);
nor U5714 (N_5714,N_4187,N_4771);
or U5715 (N_5715,N_4003,N_3654);
nor U5716 (N_5716,N_2576,N_4636);
nor U5717 (N_5717,N_4047,N_4480);
nor U5718 (N_5718,N_4005,N_2981);
nand U5719 (N_5719,N_4896,N_2864);
nor U5720 (N_5720,N_3697,N_2662);
and U5721 (N_5721,N_3975,N_2731);
or U5722 (N_5722,N_2933,N_3211);
nor U5723 (N_5723,N_3674,N_3808);
or U5724 (N_5724,N_4136,N_3053);
nor U5725 (N_5725,N_4690,N_3790);
xor U5726 (N_5726,N_4707,N_2749);
nand U5727 (N_5727,N_3391,N_4753);
and U5728 (N_5728,N_3126,N_3595);
nand U5729 (N_5729,N_3638,N_2806);
nand U5730 (N_5730,N_4372,N_3980);
or U5731 (N_5731,N_3754,N_2870);
and U5732 (N_5732,N_3799,N_4358);
or U5733 (N_5733,N_2606,N_4859);
and U5734 (N_5734,N_2841,N_3152);
and U5735 (N_5735,N_4902,N_2986);
or U5736 (N_5736,N_4182,N_4271);
and U5737 (N_5737,N_3530,N_2940);
or U5738 (N_5738,N_3653,N_4324);
and U5739 (N_5739,N_2542,N_3506);
or U5740 (N_5740,N_3684,N_4584);
or U5741 (N_5741,N_2545,N_3196);
nand U5742 (N_5742,N_4736,N_3465);
or U5743 (N_5743,N_2746,N_3085);
nand U5744 (N_5744,N_3645,N_3342);
or U5745 (N_5745,N_4216,N_3096);
or U5746 (N_5746,N_4232,N_3230);
xor U5747 (N_5747,N_2836,N_2656);
nand U5748 (N_5748,N_4642,N_4616);
or U5749 (N_5749,N_4388,N_3299);
or U5750 (N_5750,N_3997,N_2657);
nand U5751 (N_5751,N_2603,N_4864);
nor U5752 (N_5752,N_4611,N_4741);
and U5753 (N_5753,N_4471,N_4452);
xor U5754 (N_5754,N_2976,N_3023);
xnor U5755 (N_5755,N_2529,N_3047);
and U5756 (N_5756,N_4700,N_3374);
xnor U5757 (N_5757,N_3460,N_2937);
and U5758 (N_5758,N_2679,N_4297);
nor U5759 (N_5759,N_4911,N_4648);
nand U5760 (N_5760,N_2802,N_4615);
or U5761 (N_5761,N_4503,N_3317);
nor U5762 (N_5762,N_3157,N_3614);
nand U5763 (N_5763,N_4019,N_3837);
nand U5764 (N_5764,N_4796,N_4149);
or U5765 (N_5765,N_3280,N_3204);
and U5766 (N_5766,N_3219,N_3822);
nand U5767 (N_5767,N_4858,N_3245);
and U5768 (N_5768,N_3135,N_3934);
or U5769 (N_5769,N_4336,N_4036);
and U5770 (N_5770,N_4521,N_3850);
nor U5771 (N_5771,N_4684,N_3912);
nand U5772 (N_5772,N_3478,N_2735);
and U5773 (N_5773,N_3826,N_3706);
or U5774 (N_5774,N_3273,N_4180);
nand U5775 (N_5775,N_4235,N_3028);
nor U5776 (N_5776,N_4699,N_4223);
and U5777 (N_5777,N_4053,N_3499);
nor U5778 (N_5778,N_3397,N_2991);
xnor U5779 (N_5779,N_3370,N_2562);
nand U5780 (N_5780,N_4801,N_4106);
or U5781 (N_5781,N_4443,N_4812);
nand U5782 (N_5782,N_2612,N_3222);
nand U5783 (N_5783,N_2818,N_3402);
or U5784 (N_5784,N_3829,N_4624);
and U5785 (N_5785,N_4113,N_3876);
or U5786 (N_5786,N_3310,N_3639);
or U5787 (N_5787,N_3678,N_4987);
nor U5788 (N_5788,N_3672,N_3305);
nor U5789 (N_5789,N_2907,N_4415);
or U5790 (N_5790,N_3045,N_3928);
and U5791 (N_5791,N_2750,N_3445);
nand U5792 (N_5792,N_3320,N_4646);
or U5793 (N_5793,N_2594,N_4291);
or U5794 (N_5794,N_4588,N_2868);
xnor U5795 (N_5795,N_3561,N_3314);
xnor U5796 (N_5796,N_3492,N_3183);
nor U5797 (N_5797,N_3064,N_3689);
or U5798 (N_5798,N_2625,N_2661);
and U5799 (N_5799,N_3895,N_3014);
nor U5800 (N_5800,N_4798,N_3269);
and U5801 (N_5801,N_4930,N_3722);
nand U5802 (N_5802,N_4961,N_3349);
nor U5803 (N_5803,N_3418,N_4625);
nor U5804 (N_5804,N_4846,N_3885);
nor U5805 (N_5805,N_2797,N_3454);
or U5806 (N_5806,N_2896,N_3512);
or U5807 (N_5807,N_4074,N_4639);
nand U5808 (N_5808,N_4594,N_4130);
nand U5809 (N_5809,N_3548,N_2866);
xnor U5810 (N_5810,N_4543,N_4940);
nand U5811 (N_5811,N_2754,N_4981);
xor U5812 (N_5812,N_4529,N_3925);
xnor U5813 (N_5813,N_3933,N_2575);
xnor U5814 (N_5814,N_3217,N_2873);
and U5815 (N_5815,N_4086,N_3685);
nand U5816 (N_5816,N_4129,N_2674);
or U5817 (N_5817,N_4122,N_4824);
or U5818 (N_5818,N_4155,N_3018);
nor U5819 (N_5819,N_2698,N_2619);
nor U5820 (N_5820,N_4674,N_4412);
or U5821 (N_5821,N_2861,N_4341);
or U5822 (N_5822,N_3578,N_4638);
or U5823 (N_5823,N_4403,N_4943);
xnor U5824 (N_5824,N_3515,N_4393);
or U5825 (N_5825,N_4729,N_4580);
nand U5826 (N_5826,N_2521,N_4789);
or U5827 (N_5827,N_3803,N_2830);
and U5828 (N_5828,N_3795,N_3562);
or U5829 (N_5829,N_4395,N_3117);
nor U5830 (N_5830,N_4986,N_4035);
xor U5831 (N_5831,N_4441,N_3635);
nand U5832 (N_5832,N_4843,N_4792);
and U5833 (N_5833,N_2953,N_3300);
nand U5834 (N_5834,N_3384,N_3591);
or U5835 (N_5835,N_4713,N_4453);
xor U5836 (N_5836,N_4929,N_3112);
and U5837 (N_5837,N_2817,N_4928);
xnor U5838 (N_5838,N_3165,N_3938);
nand U5839 (N_5839,N_3991,N_2667);
nand U5840 (N_5840,N_3526,N_2567);
and U5841 (N_5841,N_4877,N_3412);
or U5842 (N_5842,N_3024,N_3624);
nand U5843 (N_5843,N_3239,N_3350);
or U5844 (N_5844,N_3404,N_4484);
and U5845 (N_5845,N_3172,N_3513);
nand U5846 (N_5846,N_4359,N_4444);
nor U5847 (N_5847,N_2590,N_4945);
or U5848 (N_5848,N_3479,N_4763);
and U5849 (N_5849,N_4084,N_4413);
nand U5850 (N_5850,N_2800,N_3282);
nor U5851 (N_5851,N_4177,N_4878);
nand U5852 (N_5852,N_4027,N_2889);
nor U5853 (N_5853,N_4346,N_4119);
or U5854 (N_5854,N_4913,N_2893);
and U5855 (N_5855,N_3437,N_4065);
or U5856 (N_5856,N_4994,N_4738);
or U5857 (N_5857,N_3946,N_3340);
or U5858 (N_5858,N_4091,N_2530);
or U5859 (N_5859,N_4461,N_4770);
nand U5860 (N_5860,N_3258,N_3060);
nor U5861 (N_5861,N_3708,N_4269);
nand U5862 (N_5862,N_4893,N_3343);
nand U5863 (N_5863,N_3261,N_3425);
and U5864 (N_5864,N_4396,N_2914);
and U5865 (N_5865,N_4649,N_4641);
and U5866 (N_5866,N_4980,N_2772);
nor U5867 (N_5867,N_4728,N_4226);
and U5868 (N_5868,N_3035,N_3935);
and U5869 (N_5869,N_2812,N_3449);
nand U5870 (N_5870,N_2753,N_4353);
or U5871 (N_5871,N_4969,N_2890);
nand U5872 (N_5872,N_4949,N_4399);
or U5873 (N_5873,N_2645,N_3144);
or U5874 (N_5874,N_3330,N_3276);
nand U5875 (N_5875,N_2798,N_4937);
or U5876 (N_5876,N_2557,N_2642);
nand U5877 (N_5877,N_2803,N_2882);
and U5878 (N_5878,N_4303,N_3069);
nor U5879 (N_5879,N_3254,N_4234);
or U5880 (N_5880,N_4366,N_4312);
and U5881 (N_5881,N_3691,N_2997);
or U5882 (N_5882,N_2712,N_4701);
or U5883 (N_5883,N_3800,N_3759);
or U5884 (N_5884,N_4734,N_3522);
and U5885 (N_5885,N_2904,N_3037);
nand U5886 (N_5886,N_2716,N_3443);
nand U5887 (N_5887,N_4282,N_2820);
nor U5888 (N_5888,N_4944,N_3052);
and U5889 (N_5889,N_4958,N_2623);
nand U5890 (N_5890,N_3472,N_2897);
nor U5891 (N_5891,N_4919,N_4563);
or U5892 (N_5892,N_4222,N_3534);
nand U5893 (N_5893,N_3459,N_4797);
and U5894 (N_5894,N_2611,N_2580);
nand U5895 (N_5895,N_4040,N_4390);
and U5896 (N_5896,N_3376,N_2597);
or U5897 (N_5897,N_4556,N_4628);
and U5898 (N_5898,N_2748,N_3407);
or U5899 (N_5899,N_4502,N_4400);
or U5900 (N_5900,N_3115,N_3296);
nor U5901 (N_5901,N_4473,N_3646);
nor U5902 (N_5902,N_4474,N_3809);
nand U5903 (N_5903,N_2505,N_2682);
nand U5904 (N_5904,N_4024,N_2862);
xnor U5905 (N_5905,N_3355,N_4607);
and U5906 (N_5906,N_4644,N_4735);
nand U5907 (N_5907,N_3742,N_3110);
and U5908 (N_5908,N_2926,N_3077);
nand U5909 (N_5909,N_4757,N_4488);
and U5910 (N_5910,N_3381,N_2985);
or U5911 (N_5911,N_4467,N_3080);
and U5912 (N_5912,N_3953,N_4862);
and U5913 (N_5913,N_2822,N_2838);
nor U5914 (N_5914,N_3794,N_3354);
xor U5915 (N_5915,N_4330,N_2503);
xor U5916 (N_5916,N_3125,N_3797);
nor U5917 (N_5917,N_4954,N_3686);
nand U5918 (N_5918,N_3260,N_4063);
or U5919 (N_5919,N_2855,N_3013);
nor U5920 (N_5920,N_4006,N_3090);
xor U5921 (N_5921,N_4508,N_4901);
xor U5922 (N_5922,N_3070,N_4787);
nand U5923 (N_5923,N_3188,N_2920);
and U5924 (N_5924,N_3861,N_3148);
nand U5925 (N_5925,N_3138,N_3285);
or U5926 (N_5926,N_4209,N_2957);
or U5927 (N_5927,N_3197,N_2833);
or U5928 (N_5928,N_2695,N_3776);
xnor U5929 (N_5929,N_3564,N_3026);
xor U5930 (N_5930,N_3824,N_3386);
and U5931 (N_5931,N_3745,N_4548);
or U5932 (N_5932,N_4164,N_4111);
nand U5933 (N_5933,N_4534,N_4126);
and U5934 (N_5934,N_4586,N_4059);
nand U5935 (N_5935,N_4782,N_2634);
nand U5936 (N_5936,N_4493,N_4874);
or U5937 (N_5937,N_3967,N_4598);
or U5938 (N_5938,N_4570,N_4533);
or U5939 (N_5939,N_2909,N_4010);
and U5940 (N_5940,N_3864,N_3944);
nor U5941 (N_5941,N_4349,N_3318);
nor U5942 (N_5942,N_2762,N_4204);
nand U5943 (N_5943,N_4450,N_4102);
or U5944 (N_5944,N_2694,N_4069);
nand U5945 (N_5945,N_4777,N_2774);
and U5946 (N_5946,N_2525,N_2609);
nand U5947 (N_5947,N_2857,N_2660);
or U5948 (N_5948,N_3406,N_2912);
xnor U5949 (N_5949,N_3815,N_3602);
and U5950 (N_5950,N_3643,N_3104);
nand U5951 (N_5951,N_4806,N_3461);
nand U5952 (N_5952,N_4276,N_3842);
or U5953 (N_5953,N_2831,N_4564);
nor U5954 (N_5954,N_3560,N_3868);
and U5955 (N_5955,N_2598,N_4401);
or U5956 (N_5956,N_4516,N_3598);
or U5957 (N_5957,N_4496,N_3663);
or U5958 (N_5958,N_3455,N_3122);
nand U5959 (N_5959,N_3489,N_4680);
nand U5960 (N_5960,N_4963,N_3890);
nand U5961 (N_5961,N_3554,N_4174);
xnor U5962 (N_5962,N_4257,N_4186);
nor U5963 (N_5963,N_3187,N_4150);
nand U5964 (N_5964,N_4294,N_3931);
nor U5965 (N_5965,N_4629,N_3278);
nand U5966 (N_5966,N_2641,N_4121);
and U5967 (N_5967,N_3695,N_4014);
and U5968 (N_5968,N_4095,N_3774);
nor U5969 (N_5969,N_4802,N_3915);
and U5970 (N_5970,N_3072,N_4305);
and U5971 (N_5971,N_3339,N_3399);
and U5972 (N_5972,N_3011,N_3303);
and U5973 (N_5973,N_2759,N_2610);
or U5974 (N_5974,N_3029,N_3821);
or U5975 (N_5975,N_4506,N_4124);
xor U5976 (N_5976,N_4651,N_2652);
or U5977 (N_5977,N_2584,N_4827);
nand U5978 (N_5978,N_4325,N_3979);
and U5979 (N_5979,N_4236,N_4277);
nor U5980 (N_5980,N_2554,N_2755);
xor U5981 (N_5981,N_2504,N_4490);
and U5982 (N_5982,N_3816,N_3038);
or U5983 (N_5983,N_3712,N_4090);
nor U5984 (N_5984,N_4973,N_2536);
nand U5985 (N_5985,N_4098,N_4076);
nand U5986 (N_5986,N_4525,N_4093);
and U5987 (N_5987,N_3575,N_3626);
xor U5988 (N_5988,N_2586,N_2718);
or U5989 (N_5989,N_4507,N_4805);
nor U5990 (N_5990,N_4244,N_3480);
nand U5991 (N_5991,N_3950,N_4137);
nand U5992 (N_5992,N_4875,N_3108);
and U5993 (N_5993,N_4262,N_3034);
nor U5994 (N_5994,N_4274,N_4352);
nand U5995 (N_5995,N_4158,N_4840);
nand U5996 (N_5996,N_4809,N_3782);
nor U5997 (N_5997,N_4045,N_4799);
nor U5998 (N_5998,N_4860,N_4989);
or U5999 (N_5999,N_3227,N_4932);
and U6000 (N_6000,N_4437,N_3074);
and U6001 (N_6001,N_3488,N_3153);
nand U6002 (N_6002,N_4337,N_4208);
nand U6003 (N_6003,N_4653,N_3151);
xor U6004 (N_6004,N_2579,N_3563);
nand U6005 (N_6005,N_2709,N_3929);
or U6006 (N_6006,N_2773,N_4225);
nand U6007 (N_6007,N_4781,N_4705);
and U6008 (N_6008,N_2885,N_4541);
or U6009 (N_6009,N_4510,N_4227);
nor U6010 (N_6010,N_4819,N_3651);
and U6011 (N_6011,N_2931,N_4733);
nand U6012 (N_6012,N_2844,N_4456);
nand U6013 (N_6013,N_3223,N_3252);
nand U6014 (N_6014,N_2730,N_4640);
nand U6015 (N_6015,N_3827,N_4921);
xnor U6016 (N_6016,N_4078,N_4720);
nand U6017 (N_6017,N_3475,N_4571);
and U6018 (N_6018,N_4416,N_2964);
xor U6019 (N_6019,N_3228,N_4783);
or U6020 (N_6020,N_2722,N_4971);
xor U6021 (N_6021,N_4376,N_4056);
or U6022 (N_6022,N_2684,N_2533);
nand U6023 (N_6023,N_2828,N_4803);
nor U6024 (N_6024,N_2620,N_2982);
nor U6025 (N_6025,N_4133,N_2631);
nor U6026 (N_6026,N_4307,N_2801);
nand U6027 (N_6027,N_4719,N_3750);
nand U6028 (N_6028,N_3356,N_4383);
nand U6029 (N_6029,N_4281,N_4384);
nor U6030 (N_6030,N_2944,N_4526);
xor U6031 (N_6031,N_3501,N_4605);
nand U6032 (N_6032,N_2984,N_4368);
and U6033 (N_6033,N_3756,N_3814);
nand U6034 (N_6034,N_3668,N_3466);
nand U6035 (N_6035,N_2582,N_2676);
nor U6036 (N_6036,N_2578,N_2990);
and U6037 (N_6037,N_3981,N_4147);
and U6038 (N_6038,N_3785,N_4755);
or U6039 (N_6039,N_4109,N_3192);
nand U6040 (N_6040,N_3891,N_2843);
or U6041 (N_6041,N_4883,N_2510);
and U6042 (N_6042,N_2574,N_4500);
nor U6043 (N_6043,N_2692,N_4302);
nand U6044 (N_6044,N_4430,N_3106);
xor U6045 (N_6045,N_3174,N_3140);
or U6046 (N_6046,N_4820,N_2727);
nor U6047 (N_6047,N_4105,N_3608);
nand U6048 (N_6048,N_2928,N_3676);
nor U6049 (N_6049,N_3284,N_2723);
or U6050 (N_6050,N_4844,N_3913);
nand U6051 (N_6051,N_4055,N_2686);
nand U6052 (N_6052,N_3200,N_4468);
or U6053 (N_6053,N_4108,N_4756);
nor U6054 (N_6054,N_4489,N_3961);
and U6055 (N_6055,N_3640,N_4817);
xor U6056 (N_6056,N_2705,N_3652);
or U6057 (N_6057,N_2733,N_4848);
nor U6058 (N_6058,N_3105,N_2638);
and U6059 (N_6059,N_4749,N_4863);
nor U6060 (N_6060,N_3341,N_3226);
or U6061 (N_6061,N_4156,N_4997);
nor U6062 (N_6062,N_2786,N_4224);
or U6063 (N_6063,N_4682,N_3786);
nand U6064 (N_6064,N_3659,N_3233);
xor U6065 (N_6065,N_3448,N_3283);
nand U6066 (N_6066,N_3622,N_4754);
xnor U6067 (N_6067,N_3610,N_4497);
and U6068 (N_6068,N_3178,N_4183);
and U6069 (N_6069,N_3365,N_4020);
nor U6070 (N_6070,N_4331,N_3267);
xor U6071 (N_6071,N_3068,N_4200);
and U6072 (N_6072,N_3549,N_2826);
nand U6073 (N_6073,N_3420,N_3849);
or U6074 (N_6074,N_3101,N_2950);
or U6075 (N_6075,N_3212,N_2784);
nor U6076 (N_6076,N_3270,N_4552);
or U6077 (N_6077,N_3955,N_4313);
or U6078 (N_6078,N_4608,N_3264);
and U6079 (N_6079,N_3086,N_4423);
nor U6080 (N_6080,N_3987,N_2987);
xnor U6081 (N_6081,N_4410,N_3507);
nand U6082 (N_6082,N_4198,N_4030);
xnor U6083 (N_6083,N_4582,N_2811);
or U6084 (N_6084,N_2664,N_2848);
nand U6085 (N_6085,N_3960,N_4821);
and U6086 (N_6086,N_2859,N_4087);
and U6087 (N_6087,N_3309,N_3886);
or U6088 (N_6088,N_3570,N_4357);
and U6089 (N_6089,N_3874,N_4568);
nor U6090 (N_6090,N_4845,N_2977);
nand U6091 (N_6091,N_2532,N_4903);
and U6092 (N_6092,N_2629,N_4620);
or U6093 (N_6093,N_4920,N_3907);
nor U6094 (N_6094,N_3092,N_3586);
nand U6095 (N_6095,N_4703,N_4178);
nand U6096 (N_6096,N_3677,N_3497);
nand U6097 (N_6097,N_4148,N_3076);
or U6098 (N_6098,N_4240,N_2633);
and U6099 (N_6099,N_4386,N_3136);
nor U6100 (N_6100,N_3155,N_3954);
or U6101 (N_6101,N_4079,N_4185);
nand U6102 (N_6102,N_2687,N_4946);
or U6103 (N_6103,N_2969,N_2783);
nor U6104 (N_6104,N_3574,N_4956);
or U6105 (N_6105,N_4004,N_2710);
or U6106 (N_6106,N_2932,N_4026);
nor U6107 (N_6107,N_3015,N_3114);
and U6108 (N_6108,N_4160,N_4813);
nand U6109 (N_6109,N_3059,N_2906);
and U6110 (N_6110,N_2837,N_3435);
xor U6111 (N_6111,N_4602,N_3661);
nor U6112 (N_6112,N_3368,N_3831);
nand U6113 (N_6113,N_2604,N_4769);
nand U6114 (N_6114,N_3347,N_2768);
and U6115 (N_6115,N_4596,N_4868);
or U6116 (N_6116,N_3182,N_2512);
nand U6117 (N_6117,N_2640,N_2927);
nor U6118 (N_6118,N_2531,N_4907);
or U6119 (N_6119,N_2874,N_4915);
and U6120 (N_6120,N_3442,N_4308);
nor U6121 (N_6121,N_4558,N_4842);
and U6122 (N_6122,N_2514,N_3713);
and U6123 (N_6123,N_2600,N_3071);
nand U6124 (N_6124,N_4554,N_3704);
nand U6125 (N_6125,N_3030,N_2943);
or U6126 (N_6126,N_3576,N_2622);
nand U6127 (N_6127,N_3423,N_3364);
nor U6128 (N_6128,N_4125,N_2703);
nand U6129 (N_6129,N_4266,N_2740);
nand U6130 (N_6130,N_4581,N_4314);
or U6131 (N_6131,N_2583,N_4847);
and U6132 (N_6132,N_2998,N_4472);
nor U6133 (N_6133,N_2961,N_3315);
or U6134 (N_6134,N_2791,N_3978);
nand U6135 (N_6135,N_3107,N_4683);
or U6136 (N_6136,N_2595,N_2699);
and U6137 (N_6137,N_4446,N_4714);
nor U6138 (N_6138,N_4293,N_3539);
xor U6139 (N_6139,N_2808,N_3773);
nor U6140 (N_6140,N_3656,N_4362);
xnor U6141 (N_6141,N_2872,N_2707);
xor U6142 (N_6142,N_4716,N_2972);
xnor U6143 (N_6143,N_3655,N_3968);
xor U6144 (N_6144,N_4096,N_4765);
or U6145 (N_6145,N_3496,N_4530);
or U6146 (N_6146,N_3057,N_2871);
nand U6147 (N_6147,N_2776,N_2918);
nor U6148 (N_6148,N_3835,N_4752);
nor U6149 (N_6149,N_2593,N_4363);
or U6150 (N_6150,N_3751,N_3941);
nor U6151 (N_6151,N_4315,N_3828);
or U6152 (N_6152,N_3483,N_2573);
nor U6153 (N_6153,N_3804,N_4039);
and U6154 (N_6154,N_4747,N_4730);
nand U6155 (N_6155,N_3493,N_3302);
nand U6156 (N_6156,N_2809,N_4319);
or U6157 (N_6157,N_4778,N_3577);
xor U6158 (N_6158,N_4408,N_3271);
and U6159 (N_6159,N_4925,N_3430);
nand U6160 (N_6160,N_3031,N_3847);
nand U6161 (N_6161,N_3237,N_4871);
nand U6162 (N_6162,N_3422,N_3405);
nor U6163 (N_6163,N_3762,N_3884);
xnor U6164 (N_6164,N_4545,N_2736);
nor U6165 (N_6165,N_3433,N_2534);
and U6166 (N_6166,N_4008,N_4589);
or U6167 (N_6167,N_4595,N_3532);
and U6168 (N_6168,N_3698,N_4327);
or U6169 (N_6169,N_3097,N_4067);
and U6170 (N_6170,N_2767,N_2886);
nor U6171 (N_6171,N_4381,N_2942);
and U6172 (N_6172,N_3464,N_3553);
and U6173 (N_6173,N_2958,N_3395);
and U6174 (N_6174,N_2559,N_3087);
xor U6175 (N_6175,N_4419,N_3274);
nor U6176 (N_6176,N_4537,N_2860);
xnor U6177 (N_6177,N_4599,N_4725);
nand U6178 (N_6178,N_4048,N_2846);
nand U6179 (N_6179,N_4576,N_4935);
nand U6180 (N_6180,N_3518,N_3295);
nand U6181 (N_6181,N_4088,N_3084);
nor U6182 (N_6182,N_2816,N_2899);
nand U6183 (N_6183,N_4220,N_4936);
and U6184 (N_6184,N_2697,N_2599);
nand U6185 (N_6185,N_3984,N_2900);
xor U6186 (N_6186,N_3073,N_4287);
nand U6187 (N_6187,N_3841,N_4171);
xnor U6188 (N_6188,N_4633,N_3149);
and U6189 (N_6189,N_3729,N_2968);
and U6190 (N_6190,N_4617,N_4001);
or U6191 (N_6191,N_2763,N_3291);
nor U6192 (N_6192,N_2771,N_2585);
nand U6193 (N_6193,N_4427,N_4885);
or U6194 (N_6194,N_4355,N_2766);
or U6195 (N_6195,N_4762,N_4890);
nor U6196 (N_6196,N_4201,N_3453);
or U6197 (N_6197,N_4377,N_4475);
or U6198 (N_6198,N_3033,N_4061);
nand U6199 (N_6199,N_4435,N_3592);
and U6200 (N_6200,N_2614,N_3538);
nor U6201 (N_6201,N_4635,N_3146);
or U6202 (N_6202,N_4141,N_2814);
xnor U6203 (N_6203,N_4037,N_2879);
nand U6204 (N_6204,N_3741,N_4242);
or U6205 (N_6205,N_4263,N_3664);
nand U6206 (N_6206,N_3959,N_4284);
nor U6207 (N_6207,N_4009,N_4379);
nor U6208 (N_6208,N_2669,N_3351);
xnor U6209 (N_6209,N_2757,N_3547);
nand U6210 (N_6210,N_2630,N_4127);
or U6211 (N_6211,N_3758,N_4941);
and U6212 (N_6212,N_3025,N_4748);
or U6213 (N_6213,N_3813,N_4766);
xor U6214 (N_6214,N_3458,N_4023);
or U6215 (N_6215,N_3702,N_4478);
nand U6216 (N_6216,N_4289,N_4573);
or U6217 (N_6217,N_3637,N_2851);
nor U6218 (N_6218,N_4245,N_3937);
nand U6219 (N_6219,N_4116,N_3846);
or U6220 (N_6220,N_4283,N_4265);
nand U6221 (N_6221,N_4528,N_4169);
nor U6222 (N_6222,N_3436,N_4261);
and U6223 (N_6223,N_3558,N_4887);
or U6224 (N_6224,N_3581,N_3606);
nand U6225 (N_6225,N_3552,N_3003);
and U6226 (N_6226,N_2925,N_3335);
and U6227 (N_6227,N_3787,N_4107);
or U6228 (N_6228,N_4826,N_3468);
nand U6229 (N_6229,N_3127,N_3503);
nand U6230 (N_6230,N_4260,N_4097);
xnor U6231 (N_6231,N_4685,N_4572);
nor U6232 (N_6232,N_4818,N_2911);
or U6233 (N_6233,N_2572,N_4880);
nor U6234 (N_6234,N_2804,N_2544);
nand U6235 (N_6235,N_3221,N_4924);
nor U6236 (N_6236,N_3823,N_4309);
nand U6237 (N_6237,N_3680,N_3681);
nand U6238 (N_6238,N_4767,N_3620);
nor U6239 (N_6239,N_4634,N_4499);
or U6240 (N_6240,N_4211,N_2663);
xnor U6241 (N_6241,N_3251,N_2965);
nand U6242 (N_6242,N_3431,N_2696);
nand U6243 (N_6243,N_2895,N_3160);
and U6244 (N_6244,N_2974,N_2930);
and U6245 (N_6245,N_3163,N_4894);
nand U6246 (N_6246,N_3382,N_4405);
nand U6247 (N_6247,N_3920,N_2934);
or U6248 (N_6248,N_4028,N_4538);
nor U6249 (N_6249,N_3682,N_3724);
nor U6250 (N_6250,N_4156,N_4339);
or U6251 (N_6251,N_3984,N_4431);
nor U6252 (N_6252,N_2582,N_2855);
and U6253 (N_6253,N_3566,N_2526);
or U6254 (N_6254,N_4988,N_2753);
nand U6255 (N_6255,N_4850,N_3636);
nor U6256 (N_6256,N_4804,N_3249);
nor U6257 (N_6257,N_4959,N_2585);
and U6258 (N_6258,N_3266,N_3339);
nor U6259 (N_6259,N_2598,N_3017);
or U6260 (N_6260,N_3454,N_4926);
nor U6261 (N_6261,N_4409,N_3121);
nand U6262 (N_6262,N_4064,N_3764);
nor U6263 (N_6263,N_4538,N_3047);
and U6264 (N_6264,N_3076,N_4218);
nand U6265 (N_6265,N_3676,N_2545);
nor U6266 (N_6266,N_3116,N_4355);
or U6267 (N_6267,N_4902,N_4885);
nor U6268 (N_6268,N_3510,N_4070);
or U6269 (N_6269,N_3305,N_2759);
and U6270 (N_6270,N_3403,N_4169);
or U6271 (N_6271,N_2696,N_3270);
nor U6272 (N_6272,N_3764,N_3887);
and U6273 (N_6273,N_3426,N_3833);
or U6274 (N_6274,N_4072,N_3310);
or U6275 (N_6275,N_3907,N_4256);
and U6276 (N_6276,N_4971,N_3886);
and U6277 (N_6277,N_4095,N_2951);
or U6278 (N_6278,N_4055,N_2830);
nor U6279 (N_6279,N_4450,N_3536);
nor U6280 (N_6280,N_2893,N_3781);
or U6281 (N_6281,N_2675,N_3397);
xor U6282 (N_6282,N_4982,N_3620);
or U6283 (N_6283,N_4318,N_3890);
and U6284 (N_6284,N_2625,N_3130);
and U6285 (N_6285,N_2695,N_4325);
nand U6286 (N_6286,N_4590,N_3689);
nand U6287 (N_6287,N_2700,N_3556);
nor U6288 (N_6288,N_4794,N_4999);
xor U6289 (N_6289,N_3898,N_4587);
nor U6290 (N_6290,N_4971,N_4989);
nand U6291 (N_6291,N_3850,N_3035);
and U6292 (N_6292,N_4960,N_4521);
xnor U6293 (N_6293,N_4176,N_4914);
nand U6294 (N_6294,N_4465,N_2894);
and U6295 (N_6295,N_4486,N_4329);
or U6296 (N_6296,N_4653,N_3673);
nor U6297 (N_6297,N_4406,N_3735);
or U6298 (N_6298,N_2581,N_4953);
nor U6299 (N_6299,N_3562,N_3313);
xnor U6300 (N_6300,N_3036,N_4916);
or U6301 (N_6301,N_4631,N_4698);
nor U6302 (N_6302,N_3089,N_3808);
nand U6303 (N_6303,N_4447,N_3901);
xor U6304 (N_6304,N_3853,N_3258);
and U6305 (N_6305,N_3132,N_3423);
xnor U6306 (N_6306,N_2599,N_2746);
or U6307 (N_6307,N_3355,N_4709);
nand U6308 (N_6308,N_4852,N_4749);
nor U6309 (N_6309,N_2713,N_4701);
nor U6310 (N_6310,N_3784,N_3911);
nand U6311 (N_6311,N_3132,N_4626);
or U6312 (N_6312,N_3567,N_4750);
nand U6313 (N_6313,N_4163,N_4457);
nand U6314 (N_6314,N_3845,N_4482);
or U6315 (N_6315,N_4458,N_4202);
xor U6316 (N_6316,N_3712,N_2529);
and U6317 (N_6317,N_2595,N_3045);
nor U6318 (N_6318,N_2594,N_3289);
or U6319 (N_6319,N_4458,N_4100);
and U6320 (N_6320,N_3132,N_4784);
nor U6321 (N_6321,N_4272,N_3607);
and U6322 (N_6322,N_4020,N_4524);
nor U6323 (N_6323,N_2599,N_2649);
or U6324 (N_6324,N_4223,N_3612);
nor U6325 (N_6325,N_4060,N_4630);
nor U6326 (N_6326,N_4914,N_2607);
or U6327 (N_6327,N_3120,N_2648);
and U6328 (N_6328,N_2986,N_3778);
or U6329 (N_6329,N_3765,N_4791);
and U6330 (N_6330,N_4152,N_3334);
nor U6331 (N_6331,N_2772,N_4740);
xnor U6332 (N_6332,N_3573,N_2979);
nor U6333 (N_6333,N_4896,N_2779);
and U6334 (N_6334,N_2940,N_4187);
nor U6335 (N_6335,N_4127,N_4374);
nor U6336 (N_6336,N_3346,N_3844);
and U6337 (N_6337,N_4742,N_2599);
and U6338 (N_6338,N_4112,N_3627);
nor U6339 (N_6339,N_2902,N_3516);
or U6340 (N_6340,N_2959,N_3633);
xor U6341 (N_6341,N_3874,N_2880);
and U6342 (N_6342,N_3904,N_4916);
and U6343 (N_6343,N_4105,N_3681);
nand U6344 (N_6344,N_2989,N_4170);
or U6345 (N_6345,N_3182,N_3613);
nand U6346 (N_6346,N_3980,N_3918);
or U6347 (N_6347,N_4479,N_3202);
nor U6348 (N_6348,N_3740,N_3784);
nand U6349 (N_6349,N_2782,N_2879);
nor U6350 (N_6350,N_4144,N_4078);
nor U6351 (N_6351,N_3477,N_4295);
nor U6352 (N_6352,N_3597,N_4022);
nor U6353 (N_6353,N_4130,N_3734);
nor U6354 (N_6354,N_3983,N_4020);
nor U6355 (N_6355,N_4592,N_3220);
nor U6356 (N_6356,N_3459,N_4580);
or U6357 (N_6357,N_4252,N_4836);
nor U6358 (N_6358,N_2832,N_3098);
or U6359 (N_6359,N_3976,N_2831);
and U6360 (N_6360,N_3590,N_3326);
and U6361 (N_6361,N_2869,N_3469);
nand U6362 (N_6362,N_3461,N_3556);
or U6363 (N_6363,N_3925,N_4644);
or U6364 (N_6364,N_3226,N_2948);
or U6365 (N_6365,N_4486,N_4303);
or U6366 (N_6366,N_4996,N_3808);
nor U6367 (N_6367,N_2932,N_3460);
xnor U6368 (N_6368,N_3255,N_2893);
or U6369 (N_6369,N_2971,N_2981);
and U6370 (N_6370,N_3382,N_3171);
nand U6371 (N_6371,N_4972,N_2658);
nand U6372 (N_6372,N_3908,N_3082);
xnor U6373 (N_6373,N_3210,N_3502);
nor U6374 (N_6374,N_2792,N_4302);
and U6375 (N_6375,N_4724,N_3145);
or U6376 (N_6376,N_4019,N_3594);
nor U6377 (N_6377,N_4408,N_3646);
nand U6378 (N_6378,N_3029,N_4557);
nor U6379 (N_6379,N_4694,N_4957);
nand U6380 (N_6380,N_4226,N_2740);
or U6381 (N_6381,N_4809,N_3409);
nor U6382 (N_6382,N_4719,N_4562);
or U6383 (N_6383,N_4362,N_3744);
and U6384 (N_6384,N_2535,N_4924);
nor U6385 (N_6385,N_3508,N_2572);
nand U6386 (N_6386,N_3259,N_4241);
or U6387 (N_6387,N_2679,N_2658);
nor U6388 (N_6388,N_4473,N_3172);
nand U6389 (N_6389,N_3222,N_4216);
nand U6390 (N_6390,N_3936,N_4985);
nand U6391 (N_6391,N_4126,N_3279);
nand U6392 (N_6392,N_2655,N_3699);
nor U6393 (N_6393,N_3409,N_3179);
xnor U6394 (N_6394,N_4624,N_2712);
and U6395 (N_6395,N_2680,N_4861);
nand U6396 (N_6396,N_2922,N_3259);
nand U6397 (N_6397,N_2685,N_3773);
xnor U6398 (N_6398,N_3400,N_3224);
nor U6399 (N_6399,N_3970,N_3361);
and U6400 (N_6400,N_4831,N_2953);
xnor U6401 (N_6401,N_4315,N_4252);
and U6402 (N_6402,N_4514,N_3482);
or U6403 (N_6403,N_4478,N_2978);
nor U6404 (N_6404,N_2567,N_4150);
nand U6405 (N_6405,N_2682,N_4890);
nand U6406 (N_6406,N_4253,N_4197);
and U6407 (N_6407,N_4109,N_4070);
nor U6408 (N_6408,N_4957,N_3040);
and U6409 (N_6409,N_4809,N_4328);
nand U6410 (N_6410,N_2527,N_2945);
or U6411 (N_6411,N_4692,N_4728);
nand U6412 (N_6412,N_2715,N_4182);
xor U6413 (N_6413,N_2543,N_4632);
or U6414 (N_6414,N_4327,N_3741);
or U6415 (N_6415,N_2775,N_3927);
nor U6416 (N_6416,N_3487,N_4184);
and U6417 (N_6417,N_4281,N_4310);
or U6418 (N_6418,N_3567,N_3116);
xor U6419 (N_6419,N_2556,N_3267);
nand U6420 (N_6420,N_4205,N_3540);
nor U6421 (N_6421,N_2773,N_3429);
and U6422 (N_6422,N_4802,N_3970);
and U6423 (N_6423,N_4456,N_3735);
nor U6424 (N_6424,N_2551,N_2865);
or U6425 (N_6425,N_4744,N_4279);
or U6426 (N_6426,N_2634,N_3451);
or U6427 (N_6427,N_4055,N_3805);
or U6428 (N_6428,N_3678,N_4036);
and U6429 (N_6429,N_3886,N_2532);
nand U6430 (N_6430,N_3026,N_4093);
nand U6431 (N_6431,N_4580,N_3457);
or U6432 (N_6432,N_3011,N_3429);
or U6433 (N_6433,N_3577,N_4898);
or U6434 (N_6434,N_4964,N_4818);
nor U6435 (N_6435,N_2531,N_4345);
nor U6436 (N_6436,N_2941,N_4852);
nand U6437 (N_6437,N_4467,N_2889);
or U6438 (N_6438,N_2953,N_2688);
nor U6439 (N_6439,N_4108,N_2905);
or U6440 (N_6440,N_3107,N_4121);
and U6441 (N_6441,N_3016,N_4468);
nor U6442 (N_6442,N_3685,N_3737);
and U6443 (N_6443,N_2969,N_3918);
nor U6444 (N_6444,N_3785,N_3152);
nand U6445 (N_6445,N_3034,N_2776);
or U6446 (N_6446,N_3172,N_4739);
xnor U6447 (N_6447,N_4137,N_3065);
or U6448 (N_6448,N_4468,N_4015);
or U6449 (N_6449,N_3293,N_4391);
or U6450 (N_6450,N_4334,N_4206);
or U6451 (N_6451,N_3855,N_4708);
xnor U6452 (N_6452,N_3308,N_3779);
or U6453 (N_6453,N_2699,N_3104);
nand U6454 (N_6454,N_4774,N_4798);
nor U6455 (N_6455,N_4810,N_2862);
xnor U6456 (N_6456,N_4172,N_4557);
and U6457 (N_6457,N_4547,N_4379);
nand U6458 (N_6458,N_2712,N_2663);
nor U6459 (N_6459,N_3069,N_2621);
nand U6460 (N_6460,N_3416,N_3500);
nand U6461 (N_6461,N_3924,N_4192);
or U6462 (N_6462,N_3179,N_3933);
and U6463 (N_6463,N_4551,N_2737);
and U6464 (N_6464,N_3536,N_3723);
or U6465 (N_6465,N_4757,N_2508);
nor U6466 (N_6466,N_4726,N_3956);
xor U6467 (N_6467,N_2677,N_3382);
nor U6468 (N_6468,N_4654,N_4710);
and U6469 (N_6469,N_4354,N_4994);
xor U6470 (N_6470,N_3559,N_3701);
xnor U6471 (N_6471,N_4437,N_4939);
and U6472 (N_6472,N_4656,N_3915);
nand U6473 (N_6473,N_4361,N_4037);
and U6474 (N_6474,N_2858,N_3747);
nor U6475 (N_6475,N_4999,N_4963);
nor U6476 (N_6476,N_4271,N_3081);
or U6477 (N_6477,N_3076,N_3836);
nand U6478 (N_6478,N_3841,N_2524);
nor U6479 (N_6479,N_2507,N_3563);
nand U6480 (N_6480,N_3365,N_3381);
and U6481 (N_6481,N_2609,N_4640);
and U6482 (N_6482,N_3762,N_4496);
or U6483 (N_6483,N_2850,N_3762);
and U6484 (N_6484,N_3783,N_3480);
nand U6485 (N_6485,N_2862,N_3776);
or U6486 (N_6486,N_4332,N_3110);
and U6487 (N_6487,N_4723,N_4461);
or U6488 (N_6488,N_2706,N_3734);
nand U6489 (N_6489,N_3880,N_4897);
and U6490 (N_6490,N_3004,N_4189);
nand U6491 (N_6491,N_4904,N_4915);
and U6492 (N_6492,N_4209,N_4506);
nor U6493 (N_6493,N_4558,N_3727);
nor U6494 (N_6494,N_3631,N_4941);
and U6495 (N_6495,N_4082,N_4615);
nor U6496 (N_6496,N_4443,N_2707);
nor U6497 (N_6497,N_3360,N_3062);
nand U6498 (N_6498,N_4223,N_3897);
and U6499 (N_6499,N_3328,N_3640);
and U6500 (N_6500,N_3704,N_4544);
or U6501 (N_6501,N_4033,N_2817);
nand U6502 (N_6502,N_4497,N_3619);
nand U6503 (N_6503,N_4705,N_4482);
xnor U6504 (N_6504,N_4990,N_4654);
or U6505 (N_6505,N_3778,N_4558);
nand U6506 (N_6506,N_2864,N_3644);
xnor U6507 (N_6507,N_3508,N_2644);
nor U6508 (N_6508,N_4119,N_3280);
nand U6509 (N_6509,N_3785,N_2936);
nor U6510 (N_6510,N_4946,N_3316);
and U6511 (N_6511,N_4831,N_2629);
or U6512 (N_6512,N_3319,N_3554);
nor U6513 (N_6513,N_3183,N_2705);
nor U6514 (N_6514,N_4228,N_2563);
nand U6515 (N_6515,N_3776,N_4948);
and U6516 (N_6516,N_4396,N_4332);
nor U6517 (N_6517,N_4472,N_3240);
nand U6518 (N_6518,N_3029,N_4561);
and U6519 (N_6519,N_3997,N_2747);
or U6520 (N_6520,N_3407,N_4629);
nand U6521 (N_6521,N_2778,N_3199);
and U6522 (N_6522,N_3904,N_2764);
or U6523 (N_6523,N_4365,N_4399);
nand U6524 (N_6524,N_3336,N_3355);
nor U6525 (N_6525,N_2735,N_2946);
and U6526 (N_6526,N_3177,N_4299);
or U6527 (N_6527,N_4668,N_2622);
nor U6528 (N_6528,N_3047,N_3331);
and U6529 (N_6529,N_3952,N_4958);
nor U6530 (N_6530,N_3712,N_3071);
nor U6531 (N_6531,N_3341,N_4978);
or U6532 (N_6532,N_4245,N_4563);
nand U6533 (N_6533,N_4033,N_4564);
nand U6534 (N_6534,N_4118,N_4396);
and U6535 (N_6535,N_3774,N_3777);
nor U6536 (N_6536,N_3919,N_2813);
nor U6537 (N_6537,N_3391,N_4805);
or U6538 (N_6538,N_3137,N_2578);
and U6539 (N_6539,N_2511,N_4197);
and U6540 (N_6540,N_3908,N_2912);
xnor U6541 (N_6541,N_4117,N_2917);
nor U6542 (N_6542,N_4722,N_4694);
nand U6543 (N_6543,N_3025,N_4594);
xnor U6544 (N_6544,N_3447,N_3415);
or U6545 (N_6545,N_3902,N_2857);
or U6546 (N_6546,N_4380,N_3923);
xor U6547 (N_6547,N_4944,N_3455);
or U6548 (N_6548,N_4771,N_2926);
nand U6549 (N_6549,N_2633,N_4429);
and U6550 (N_6550,N_3216,N_3166);
nand U6551 (N_6551,N_4961,N_3815);
nor U6552 (N_6552,N_2654,N_2593);
nand U6553 (N_6553,N_4880,N_2598);
nor U6554 (N_6554,N_3262,N_4582);
nand U6555 (N_6555,N_3932,N_2641);
and U6556 (N_6556,N_3062,N_2634);
nand U6557 (N_6557,N_4173,N_3076);
nor U6558 (N_6558,N_3051,N_4375);
and U6559 (N_6559,N_3900,N_3541);
nor U6560 (N_6560,N_4889,N_3118);
and U6561 (N_6561,N_2798,N_4822);
nand U6562 (N_6562,N_3583,N_3853);
nand U6563 (N_6563,N_3074,N_4352);
nand U6564 (N_6564,N_2508,N_3763);
nor U6565 (N_6565,N_3656,N_4311);
nor U6566 (N_6566,N_4281,N_3818);
or U6567 (N_6567,N_2628,N_3531);
and U6568 (N_6568,N_4574,N_4596);
and U6569 (N_6569,N_3553,N_3065);
nand U6570 (N_6570,N_3289,N_4548);
and U6571 (N_6571,N_3448,N_3183);
nor U6572 (N_6572,N_2926,N_3321);
or U6573 (N_6573,N_3929,N_4042);
nor U6574 (N_6574,N_3236,N_2550);
or U6575 (N_6575,N_2706,N_2769);
and U6576 (N_6576,N_2692,N_3235);
nor U6577 (N_6577,N_4897,N_3352);
nand U6578 (N_6578,N_4188,N_4564);
or U6579 (N_6579,N_3686,N_3284);
nand U6580 (N_6580,N_2876,N_3523);
and U6581 (N_6581,N_4276,N_4477);
or U6582 (N_6582,N_4152,N_3102);
nor U6583 (N_6583,N_4416,N_2653);
nand U6584 (N_6584,N_4934,N_4140);
and U6585 (N_6585,N_2906,N_3924);
and U6586 (N_6586,N_4972,N_4349);
and U6587 (N_6587,N_2721,N_4519);
or U6588 (N_6588,N_4262,N_3229);
and U6589 (N_6589,N_3262,N_4365);
and U6590 (N_6590,N_2716,N_3295);
nor U6591 (N_6591,N_2949,N_4116);
or U6592 (N_6592,N_2975,N_4797);
xor U6593 (N_6593,N_4989,N_2684);
nor U6594 (N_6594,N_4388,N_2757);
and U6595 (N_6595,N_3616,N_3130);
nor U6596 (N_6596,N_3385,N_4872);
nor U6597 (N_6597,N_3828,N_3974);
nand U6598 (N_6598,N_2681,N_3078);
nor U6599 (N_6599,N_3415,N_2525);
and U6600 (N_6600,N_4835,N_4939);
or U6601 (N_6601,N_3186,N_3056);
and U6602 (N_6602,N_4536,N_2668);
xor U6603 (N_6603,N_4637,N_4194);
nand U6604 (N_6604,N_3363,N_3127);
nand U6605 (N_6605,N_2585,N_4775);
nand U6606 (N_6606,N_4351,N_3742);
xnor U6607 (N_6607,N_4769,N_2842);
nand U6608 (N_6608,N_3806,N_4021);
and U6609 (N_6609,N_3657,N_4010);
nand U6610 (N_6610,N_2559,N_2675);
nand U6611 (N_6611,N_3319,N_4952);
or U6612 (N_6612,N_3047,N_4117);
nand U6613 (N_6613,N_3617,N_3963);
nand U6614 (N_6614,N_3633,N_3092);
xor U6615 (N_6615,N_3949,N_2508);
and U6616 (N_6616,N_4179,N_2992);
nor U6617 (N_6617,N_3502,N_4403);
xor U6618 (N_6618,N_4411,N_4583);
xnor U6619 (N_6619,N_4673,N_3379);
xnor U6620 (N_6620,N_2555,N_2713);
and U6621 (N_6621,N_4118,N_3684);
nand U6622 (N_6622,N_3679,N_3673);
xnor U6623 (N_6623,N_4326,N_3303);
xnor U6624 (N_6624,N_2917,N_4627);
xnor U6625 (N_6625,N_2880,N_3987);
nor U6626 (N_6626,N_3353,N_4687);
or U6627 (N_6627,N_4254,N_3921);
nand U6628 (N_6628,N_4926,N_4567);
nand U6629 (N_6629,N_4981,N_2638);
nand U6630 (N_6630,N_3442,N_3941);
xor U6631 (N_6631,N_3521,N_2607);
nor U6632 (N_6632,N_4103,N_4364);
nor U6633 (N_6633,N_3963,N_3228);
nor U6634 (N_6634,N_3918,N_4226);
or U6635 (N_6635,N_3434,N_4434);
xor U6636 (N_6636,N_2990,N_4005);
or U6637 (N_6637,N_4932,N_4642);
nand U6638 (N_6638,N_3788,N_4086);
nor U6639 (N_6639,N_2768,N_4650);
nor U6640 (N_6640,N_2878,N_2779);
nor U6641 (N_6641,N_3816,N_3209);
or U6642 (N_6642,N_3732,N_3071);
nand U6643 (N_6643,N_4305,N_2552);
nor U6644 (N_6644,N_3833,N_2733);
and U6645 (N_6645,N_4943,N_3337);
and U6646 (N_6646,N_2911,N_4015);
nand U6647 (N_6647,N_4231,N_4781);
nor U6648 (N_6648,N_4104,N_3228);
or U6649 (N_6649,N_4425,N_4193);
and U6650 (N_6650,N_3828,N_4367);
xor U6651 (N_6651,N_3680,N_2693);
nor U6652 (N_6652,N_2923,N_3047);
and U6653 (N_6653,N_3285,N_2795);
nor U6654 (N_6654,N_3390,N_4880);
and U6655 (N_6655,N_4393,N_4573);
or U6656 (N_6656,N_4800,N_3231);
xnor U6657 (N_6657,N_4945,N_3877);
nor U6658 (N_6658,N_4342,N_2926);
and U6659 (N_6659,N_4446,N_3411);
and U6660 (N_6660,N_3267,N_4557);
or U6661 (N_6661,N_4643,N_4586);
nor U6662 (N_6662,N_4442,N_3809);
xor U6663 (N_6663,N_4782,N_4417);
nor U6664 (N_6664,N_4973,N_4777);
xor U6665 (N_6665,N_2652,N_4657);
nor U6666 (N_6666,N_3816,N_4565);
nor U6667 (N_6667,N_3803,N_3920);
or U6668 (N_6668,N_4048,N_3259);
nor U6669 (N_6669,N_3459,N_3694);
nor U6670 (N_6670,N_2552,N_4137);
or U6671 (N_6671,N_3409,N_2575);
nor U6672 (N_6672,N_2968,N_4376);
and U6673 (N_6673,N_3701,N_2531);
and U6674 (N_6674,N_2883,N_3730);
nor U6675 (N_6675,N_3748,N_2929);
nor U6676 (N_6676,N_3439,N_4078);
nor U6677 (N_6677,N_4666,N_4296);
xor U6678 (N_6678,N_4163,N_3616);
xor U6679 (N_6679,N_3377,N_2585);
and U6680 (N_6680,N_2905,N_3057);
or U6681 (N_6681,N_4975,N_4976);
or U6682 (N_6682,N_3136,N_3642);
or U6683 (N_6683,N_2864,N_3940);
or U6684 (N_6684,N_3787,N_3633);
and U6685 (N_6685,N_2572,N_4479);
and U6686 (N_6686,N_4362,N_3399);
nand U6687 (N_6687,N_2899,N_3415);
nor U6688 (N_6688,N_4581,N_3760);
or U6689 (N_6689,N_3625,N_3485);
nor U6690 (N_6690,N_2614,N_3269);
and U6691 (N_6691,N_4512,N_2604);
nand U6692 (N_6692,N_3217,N_3151);
nand U6693 (N_6693,N_4184,N_4104);
nor U6694 (N_6694,N_4463,N_3796);
or U6695 (N_6695,N_3028,N_3876);
or U6696 (N_6696,N_3554,N_3218);
xnor U6697 (N_6697,N_2630,N_3191);
nor U6698 (N_6698,N_3369,N_3955);
or U6699 (N_6699,N_2712,N_4390);
nand U6700 (N_6700,N_4586,N_3314);
or U6701 (N_6701,N_4311,N_3384);
nor U6702 (N_6702,N_3202,N_2631);
and U6703 (N_6703,N_3850,N_3433);
nor U6704 (N_6704,N_2633,N_2679);
and U6705 (N_6705,N_3838,N_3280);
nand U6706 (N_6706,N_2543,N_3818);
or U6707 (N_6707,N_3565,N_3787);
and U6708 (N_6708,N_4936,N_2869);
and U6709 (N_6709,N_4443,N_4690);
nor U6710 (N_6710,N_4315,N_2625);
and U6711 (N_6711,N_2552,N_2959);
and U6712 (N_6712,N_2987,N_3751);
nand U6713 (N_6713,N_4567,N_4873);
xor U6714 (N_6714,N_2745,N_3597);
nor U6715 (N_6715,N_4182,N_2770);
nor U6716 (N_6716,N_3170,N_4426);
and U6717 (N_6717,N_2672,N_4933);
and U6718 (N_6718,N_2942,N_3626);
or U6719 (N_6719,N_2670,N_4831);
nand U6720 (N_6720,N_3951,N_4426);
or U6721 (N_6721,N_3689,N_2846);
xnor U6722 (N_6722,N_4572,N_4153);
nand U6723 (N_6723,N_3444,N_4955);
or U6724 (N_6724,N_4050,N_3133);
and U6725 (N_6725,N_4753,N_4346);
nor U6726 (N_6726,N_3000,N_4388);
or U6727 (N_6727,N_4442,N_3693);
nor U6728 (N_6728,N_4276,N_4720);
or U6729 (N_6729,N_4376,N_3432);
and U6730 (N_6730,N_3540,N_2609);
and U6731 (N_6731,N_2972,N_4451);
nand U6732 (N_6732,N_4871,N_3341);
or U6733 (N_6733,N_4131,N_4667);
nand U6734 (N_6734,N_4683,N_4989);
nor U6735 (N_6735,N_3020,N_3706);
nor U6736 (N_6736,N_2616,N_4478);
xnor U6737 (N_6737,N_4806,N_3498);
nor U6738 (N_6738,N_2892,N_4575);
and U6739 (N_6739,N_4189,N_2971);
or U6740 (N_6740,N_4561,N_4704);
and U6741 (N_6741,N_2981,N_4166);
nand U6742 (N_6742,N_4074,N_4175);
nor U6743 (N_6743,N_4663,N_4569);
xor U6744 (N_6744,N_4278,N_4263);
nor U6745 (N_6745,N_2553,N_3021);
or U6746 (N_6746,N_4313,N_3835);
xnor U6747 (N_6747,N_4148,N_3330);
and U6748 (N_6748,N_2598,N_3624);
or U6749 (N_6749,N_4657,N_4744);
nand U6750 (N_6750,N_3218,N_3456);
and U6751 (N_6751,N_3113,N_3818);
or U6752 (N_6752,N_3498,N_4388);
nor U6753 (N_6753,N_4550,N_3496);
nand U6754 (N_6754,N_2510,N_2623);
nor U6755 (N_6755,N_4097,N_2708);
nor U6756 (N_6756,N_3095,N_2607);
xor U6757 (N_6757,N_4245,N_4101);
or U6758 (N_6758,N_2970,N_3295);
or U6759 (N_6759,N_4955,N_3303);
nand U6760 (N_6760,N_4472,N_4135);
or U6761 (N_6761,N_4004,N_3073);
and U6762 (N_6762,N_4296,N_3686);
and U6763 (N_6763,N_3951,N_3261);
and U6764 (N_6764,N_3169,N_3588);
nor U6765 (N_6765,N_2654,N_3937);
nor U6766 (N_6766,N_4044,N_4376);
or U6767 (N_6767,N_2784,N_2585);
nor U6768 (N_6768,N_3511,N_3850);
nand U6769 (N_6769,N_4193,N_2590);
xor U6770 (N_6770,N_2756,N_2637);
and U6771 (N_6771,N_3990,N_3878);
xor U6772 (N_6772,N_3875,N_3299);
nor U6773 (N_6773,N_2606,N_4604);
and U6774 (N_6774,N_3351,N_2681);
or U6775 (N_6775,N_3865,N_2852);
nor U6776 (N_6776,N_2985,N_4603);
xor U6777 (N_6777,N_3435,N_2538);
nor U6778 (N_6778,N_4597,N_3384);
and U6779 (N_6779,N_2539,N_3216);
and U6780 (N_6780,N_3209,N_3469);
nand U6781 (N_6781,N_2763,N_3038);
xnor U6782 (N_6782,N_4563,N_2589);
nand U6783 (N_6783,N_4301,N_3452);
or U6784 (N_6784,N_4547,N_4216);
and U6785 (N_6785,N_3474,N_4871);
and U6786 (N_6786,N_4549,N_3561);
or U6787 (N_6787,N_2581,N_3614);
nor U6788 (N_6788,N_4095,N_2969);
and U6789 (N_6789,N_3540,N_2866);
or U6790 (N_6790,N_4031,N_3583);
or U6791 (N_6791,N_4017,N_4597);
and U6792 (N_6792,N_2629,N_4614);
xor U6793 (N_6793,N_3966,N_4496);
and U6794 (N_6794,N_3528,N_4290);
nor U6795 (N_6795,N_2676,N_3164);
nand U6796 (N_6796,N_4207,N_4031);
or U6797 (N_6797,N_2632,N_4722);
or U6798 (N_6798,N_4402,N_3944);
or U6799 (N_6799,N_2591,N_3512);
nand U6800 (N_6800,N_3472,N_3745);
nand U6801 (N_6801,N_3182,N_2720);
or U6802 (N_6802,N_2638,N_3326);
xor U6803 (N_6803,N_3113,N_4994);
and U6804 (N_6804,N_3755,N_4462);
nor U6805 (N_6805,N_4888,N_2710);
nor U6806 (N_6806,N_4214,N_2727);
nand U6807 (N_6807,N_3747,N_4844);
xnor U6808 (N_6808,N_4564,N_2713);
nor U6809 (N_6809,N_4469,N_3968);
nor U6810 (N_6810,N_2638,N_2794);
or U6811 (N_6811,N_4896,N_3601);
and U6812 (N_6812,N_3052,N_3312);
xnor U6813 (N_6813,N_3908,N_4217);
or U6814 (N_6814,N_3955,N_3450);
nand U6815 (N_6815,N_2576,N_4022);
nand U6816 (N_6816,N_4421,N_3156);
or U6817 (N_6817,N_3590,N_3188);
nand U6818 (N_6818,N_4200,N_4840);
or U6819 (N_6819,N_2580,N_4527);
xor U6820 (N_6820,N_3977,N_4949);
nand U6821 (N_6821,N_2897,N_4269);
or U6822 (N_6822,N_2648,N_3861);
xnor U6823 (N_6823,N_4928,N_3210);
or U6824 (N_6824,N_4575,N_4563);
nor U6825 (N_6825,N_3190,N_3719);
or U6826 (N_6826,N_3502,N_4692);
nor U6827 (N_6827,N_2960,N_2772);
or U6828 (N_6828,N_3263,N_2522);
or U6829 (N_6829,N_3573,N_3367);
nor U6830 (N_6830,N_4742,N_3100);
and U6831 (N_6831,N_3728,N_4769);
and U6832 (N_6832,N_2608,N_4002);
or U6833 (N_6833,N_4388,N_3987);
and U6834 (N_6834,N_4675,N_2508);
or U6835 (N_6835,N_2686,N_3054);
and U6836 (N_6836,N_4709,N_4071);
and U6837 (N_6837,N_2747,N_2690);
nor U6838 (N_6838,N_4143,N_4246);
nand U6839 (N_6839,N_4377,N_3571);
xnor U6840 (N_6840,N_3392,N_4993);
xnor U6841 (N_6841,N_3311,N_3102);
or U6842 (N_6842,N_3004,N_4592);
and U6843 (N_6843,N_3305,N_3760);
nor U6844 (N_6844,N_4948,N_2695);
and U6845 (N_6845,N_2745,N_4189);
nand U6846 (N_6846,N_3597,N_2916);
and U6847 (N_6847,N_2529,N_3152);
and U6848 (N_6848,N_4428,N_2983);
and U6849 (N_6849,N_4574,N_2557);
nor U6850 (N_6850,N_3281,N_4757);
nor U6851 (N_6851,N_4718,N_4434);
nor U6852 (N_6852,N_4913,N_3203);
and U6853 (N_6853,N_3395,N_2811);
nand U6854 (N_6854,N_4234,N_4673);
and U6855 (N_6855,N_2591,N_3309);
nor U6856 (N_6856,N_3836,N_2757);
nand U6857 (N_6857,N_2896,N_4657);
nand U6858 (N_6858,N_3442,N_3431);
xnor U6859 (N_6859,N_4681,N_4492);
nand U6860 (N_6860,N_3082,N_2570);
nor U6861 (N_6861,N_2660,N_4715);
and U6862 (N_6862,N_2925,N_4246);
nand U6863 (N_6863,N_3925,N_3930);
or U6864 (N_6864,N_3901,N_4107);
xnor U6865 (N_6865,N_4739,N_2509);
and U6866 (N_6866,N_2999,N_2570);
nor U6867 (N_6867,N_4826,N_3282);
or U6868 (N_6868,N_3505,N_2909);
nor U6869 (N_6869,N_2535,N_4275);
or U6870 (N_6870,N_4285,N_3282);
xnor U6871 (N_6871,N_4323,N_2548);
xnor U6872 (N_6872,N_3250,N_3706);
xnor U6873 (N_6873,N_3554,N_4637);
nor U6874 (N_6874,N_2856,N_3525);
nor U6875 (N_6875,N_4144,N_2628);
nor U6876 (N_6876,N_4250,N_3784);
xnor U6877 (N_6877,N_4388,N_3285);
nor U6878 (N_6878,N_4330,N_4556);
nor U6879 (N_6879,N_3069,N_3461);
or U6880 (N_6880,N_3015,N_2646);
xor U6881 (N_6881,N_3946,N_2940);
nor U6882 (N_6882,N_2923,N_3517);
and U6883 (N_6883,N_4530,N_3585);
and U6884 (N_6884,N_4969,N_3742);
xnor U6885 (N_6885,N_3478,N_3508);
xor U6886 (N_6886,N_4498,N_3433);
or U6887 (N_6887,N_3787,N_4272);
nand U6888 (N_6888,N_4345,N_3722);
or U6889 (N_6889,N_4517,N_2751);
and U6890 (N_6890,N_3253,N_2511);
nand U6891 (N_6891,N_3165,N_4483);
and U6892 (N_6892,N_3807,N_4355);
and U6893 (N_6893,N_4470,N_2717);
or U6894 (N_6894,N_2504,N_3171);
or U6895 (N_6895,N_4058,N_4363);
nor U6896 (N_6896,N_2510,N_3110);
nand U6897 (N_6897,N_3213,N_4375);
and U6898 (N_6898,N_2896,N_3343);
nor U6899 (N_6899,N_3959,N_3633);
nor U6900 (N_6900,N_4134,N_4824);
nand U6901 (N_6901,N_4491,N_4390);
nor U6902 (N_6902,N_4572,N_4778);
nor U6903 (N_6903,N_2983,N_4725);
nor U6904 (N_6904,N_4000,N_4537);
nor U6905 (N_6905,N_4477,N_3303);
and U6906 (N_6906,N_3168,N_3575);
nor U6907 (N_6907,N_4867,N_2523);
xor U6908 (N_6908,N_2646,N_3613);
or U6909 (N_6909,N_3887,N_4715);
and U6910 (N_6910,N_3590,N_4256);
or U6911 (N_6911,N_3040,N_4727);
or U6912 (N_6912,N_4791,N_4483);
nor U6913 (N_6913,N_3389,N_4204);
or U6914 (N_6914,N_4616,N_3797);
nor U6915 (N_6915,N_3051,N_2737);
or U6916 (N_6916,N_3012,N_3540);
nor U6917 (N_6917,N_4010,N_4502);
xnor U6918 (N_6918,N_4590,N_3841);
or U6919 (N_6919,N_4405,N_2891);
xnor U6920 (N_6920,N_3066,N_3018);
and U6921 (N_6921,N_4656,N_3223);
or U6922 (N_6922,N_3639,N_3825);
nand U6923 (N_6923,N_3527,N_2914);
nand U6924 (N_6924,N_3810,N_4030);
and U6925 (N_6925,N_4844,N_3007);
xnor U6926 (N_6926,N_2678,N_4330);
nand U6927 (N_6927,N_2850,N_2529);
xnor U6928 (N_6928,N_3799,N_3359);
and U6929 (N_6929,N_3410,N_3089);
or U6930 (N_6930,N_3760,N_3109);
and U6931 (N_6931,N_3985,N_3737);
xor U6932 (N_6932,N_4892,N_3450);
nor U6933 (N_6933,N_4145,N_4900);
or U6934 (N_6934,N_3886,N_3894);
nor U6935 (N_6935,N_2506,N_3921);
nand U6936 (N_6936,N_4147,N_2756);
xor U6937 (N_6937,N_3296,N_4424);
nor U6938 (N_6938,N_3435,N_3805);
or U6939 (N_6939,N_3477,N_3857);
nor U6940 (N_6940,N_4565,N_3087);
xor U6941 (N_6941,N_4928,N_4977);
and U6942 (N_6942,N_3927,N_4782);
nor U6943 (N_6943,N_3581,N_2916);
or U6944 (N_6944,N_3626,N_4921);
nor U6945 (N_6945,N_2766,N_3800);
nand U6946 (N_6946,N_4994,N_3609);
and U6947 (N_6947,N_2522,N_3700);
nor U6948 (N_6948,N_2597,N_3721);
or U6949 (N_6949,N_3299,N_2778);
or U6950 (N_6950,N_3490,N_3441);
nand U6951 (N_6951,N_4376,N_2849);
nor U6952 (N_6952,N_2943,N_4814);
or U6953 (N_6953,N_3961,N_4421);
xnor U6954 (N_6954,N_3949,N_3028);
and U6955 (N_6955,N_3597,N_3824);
or U6956 (N_6956,N_4910,N_4109);
nand U6957 (N_6957,N_3919,N_3445);
nand U6958 (N_6958,N_2957,N_4447);
and U6959 (N_6959,N_3414,N_4982);
and U6960 (N_6960,N_4787,N_4805);
nor U6961 (N_6961,N_3352,N_3320);
nor U6962 (N_6962,N_3415,N_4563);
nor U6963 (N_6963,N_4688,N_4575);
nor U6964 (N_6964,N_4107,N_3744);
nor U6965 (N_6965,N_3257,N_2966);
nor U6966 (N_6966,N_4641,N_3475);
xnor U6967 (N_6967,N_4930,N_3400);
nor U6968 (N_6968,N_4231,N_3472);
and U6969 (N_6969,N_4946,N_2926);
xor U6970 (N_6970,N_4993,N_4443);
xnor U6971 (N_6971,N_3460,N_4374);
xnor U6972 (N_6972,N_3436,N_3297);
nand U6973 (N_6973,N_4000,N_2889);
and U6974 (N_6974,N_4625,N_4587);
nand U6975 (N_6975,N_4696,N_4820);
and U6976 (N_6976,N_3361,N_3388);
nor U6977 (N_6977,N_4031,N_3068);
and U6978 (N_6978,N_3034,N_4577);
nor U6979 (N_6979,N_2671,N_2807);
or U6980 (N_6980,N_4979,N_4670);
and U6981 (N_6981,N_4267,N_3459);
nand U6982 (N_6982,N_3318,N_3339);
and U6983 (N_6983,N_2909,N_3627);
nand U6984 (N_6984,N_3621,N_4368);
nand U6985 (N_6985,N_2954,N_3638);
or U6986 (N_6986,N_2660,N_2841);
and U6987 (N_6987,N_2686,N_3017);
and U6988 (N_6988,N_4459,N_2548);
nand U6989 (N_6989,N_4286,N_3627);
nand U6990 (N_6990,N_4264,N_4708);
or U6991 (N_6991,N_3578,N_2815);
and U6992 (N_6992,N_2895,N_4059);
nor U6993 (N_6993,N_4610,N_3985);
nand U6994 (N_6994,N_4656,N_4633);
nand U6995 (N_6995,N_3353,N_2802);
nor U6996 (N_6996,N_4412,N_4764);
nor U6997 (N_6997,N_3671,N_2556);
xor U6998 (N_6998,N_4284,N_4684);
or U6999 (N_6999,N_2781,N_2824);
nor U7000 (N_7000,N_4955,N_4655);
and U7001 (N_7001,N_3858,N_2856);
nand U7002 (N_7002,N_4850,N_4693);
or U7003 (N_7003,N_2965,N_3617);
and U7004 (N_7004,N_4362,N_4664);
xnor U7005 (N_7005,N_3090,N_4447);
or U7006 (N_7006,N_4928,N_3907);
nor U7007 (N_7007,N_3507,N_4297);
or U7008 (N_7008,N_3345,N_3220);
or U7009 (N_7009,N_4371,N_3241);
and U7010 (N_7010,N_4748,N_3324);
or U7011 (N_7011,N_3919,N_3107);
nor U7012 (N_7012,N_4071,N_3924);
nor U7013 (N_7013,N_2878,N_3464);
nand U7014 (N_7014,N_3434,N_2553);
xnor U7015 (N_7015,N_3145,N_3749);
xnor U7016 (N_7016,N_3580,N_3378);
nand U7017 (N_7017,N_2852,N_2574);
nand U7018 (N_7018,N_2559,N_4041);
xor U7019 (N_7019,N_4190,N_3309);
and U7020 (N_7020,N_2940,N_4594);
or U7021 (N_7021,N_2744,N_4824);
nand U7022 (N_7022,N_4143,N_4719);
nor U7023 (N_7023,N_4502,N_3526);
nor U7024 (N_7024,N_4061,N_4376);
and U7025 (N_7025,N_3902,N_3637);
nor U7026 (N_7026,N_4311,N_3973);
nor U7027 (N_7027,N_3155,N_3463);
nor U7028 (N_7028,N_4540,N_3491);
and U7029 (N_7029,N_3558,N_3431);
and U7030 (N_7030,N_3584,N_3819);
and U7031 (N_7031,N_2869,N_3520);
nor U7032 (N_7032,N_3533,N_4239);
or U7033 (N_7033,N_4116,N_4785);
or U7034 (N_7034,N_3279,N_3845);
nand U7035 (N_7035,N_3713,N_4504);
or U7036 (N_7036,N_4515,N_3047);
nand U7037 (N_7037,N_4907,N_2732);
or U7038 (N_7038,N_2751,N_4178);
nand U7039 (N_7039,N_3591,N_4474);
or U7040 (N_7040,N_3056,N_3904);
nor U7041 (N_7041,N_4348,N_3605);
nand U7042 (N_7042,N_3163,N_4352);
and U7043 (N_7043,N_4894,N_3453);
nor U7044 (N_7044,N_2658,N_3144);
and U7045 (N_7045,N_2604,N_4681);
nor U7046 (N_7046,N_4271,N_3890);
nor U7047 (N_7047,N_3686,N_3175);
and U7048 (N_7048,N_3681,N_2964);
or U7049 (N_7049,N_3554,N_3974);
nand U7050 (N_7050,N_3086,N_3286);
and U7051 (N_7051,N_3034,N_4756);
nand U7052 (N_7052,N_4649,N_4774);
and U7053 (N_7053,N_4034,N_4937);
nand U7054 (N_7054,N_2773,N_2842);
or U7055 (N_7055,N_3676,N_4097);
and U7056 (N_7056,N_2881,N_4372);
nand U7057 (N_7057,N_3882,N_3550);
and U7058 (N_7058,N_4323,N_2717);
nand U7059 (N_7059,N_4325,N_4666);
xnor U7060 (N_7060,N_3921,N_4934);
or U7061 (N_7061,N_2797,N_4056);
nand U7062 (N_7062,N_2880,N_3357);
nor U7063 (N_7063,N_2934,N_2958);
and U7064 (N_7064,N_3406,N_2923);
xor U7065 (N_7065,N_3359,N_3333);
nand U7066 (N_7066,N_3317,N_3633);
nor U7067 (N_7067,N_2866,N_4163);
and U7068 (N_7068,N_3258,N_2635);
nor U7069 (N_7069,N_2607,N_2824);
or U7070 (N_7070,N_4840,N_4804);
nor U7071 (N_7071,N_3210,N_3969);
nor U7072 (N_7072,N_2874,N_4538);
and U7073 (N_7073,N_3778,N_3384);
or U7074 (N_7074,N_4710,N_2854);
nand U7075 (N_7075,N_2818,N_3231);
or U7076 (N_7076,N_4544,N_4599);
xor U7077 (N_7077,N_3396,N_2628);
nand U7078 (N_7078,N_4755,N_4287);
nand U7079 (N_7079,N_2807,N_3029);
or U7080 (N_7080,N_3694,N_4265);
nor U7081 (N_7081,N_2637,N_3833);
or U7082 (N_7082,N_4920,N_3577);
nor U7083 (N_7083,N_3385,N_3292);
nand U7084 (N_7084,N_3724,N_2832);
nand U7085 (N_7085,N_3965,N_4935);
and U7086 (N_7086,N_3168,N_4858);
nand U7087 (N_7087,N_2506,N_3109);
or U7088 (N_7088,N_3689,N_2503);
and U7089 (N_7089,N_4350,N_3610);
and U7090 (N_7090,N_4208,N_3575);
or U7091 (N_7091,N_4200,N_3003);
nand U7092 (N_7092,N_3431,N_2649);
nand U7093 (N_7093,N_2645,N_4182);
nand U7094 (N_7094,N_2815,N_4018);
nor U7095 (N_7095,N_4687,N_4437);
nor U7096 (N_7096,N_3009,N_3194);
xnor U7097 (N_7097,N_4314,N_4044);
nor U7098 (N_7098,N_3111,N_4854);
nand U7099 (N_7099,N_3989,N_2821);
nand U7100 (N_7100,N_4254,N_3645);
xor U7101 (N_7101,N_2901,N_3672);
nor U7102 (N_7102,N_4620,N_2568);
xor U7103 (N_7103,N_2777,N_4521);
and U7104 (N_7104,N_2929,N_3637);
or U7105 (N_7105,N_2858,N_2800);
nand U7106 (N_7106,N_4188,N_3568);
nor U7107 (N_7107,N_4031,N_4380);
or U7108 (N_7108,N_2550,N_4531);
or U7109 (N_7109,N_3300,N_4424);
and U7110 (N_7110,N_4954,N_4881);
nand U7111 (N_7111,N_3204,N_4309);
or U7112 (N_7112,N_3855,N_3581);
or U7113 (N_7113,N_4673,N_4895);
xor U7114 (N_7114,N_4770,N_4157);
and U7115 (N_7115,N_2792,N_3321);
or U7116 (N_7116,N_3282,N_4315);
nor U7117 (N_7117,N_4166,N_4806);
nand U7118 (N_7118,N_2862,N_3934);
nand U7119 (N_7119,N_3655,N_4223);
or U7120 (N_7120,N_3607,N_4008);
and U7121 (N_7121,N_2635,N_4484);
nand U7122 (N_7122,N_4235,N_4613);
and U7123 (N_7123,N_2537,N_3359);
nor U7124 (N_7124,N_3142,N_3423);
and U7125 (N_7125,N_3729,N_2846);
xnor U7126 (N_7126,N_4164,N_4930);
nor U7127 (N_7127,N_3164,N_2565);
or U7128 (N_7128,N_4501,N_4865);
nand U7129 (N_7129,N_3382,N_4147);
or U7130 (N_7130,N_2826,N_4316);
or U7131 (N_7131,N_3385,N_3667);
nand U7132 (N_7132,N_2743,N_2599);
and U7133 (N_7133,N_2645,N_4031);
xor U7134 (N_7134,N_4187,N_2966);
nor U7135 (N_7135,N_3797,N_2826);
or U7136 (N_7136,N_3908,N_2830);
or U7137 (N_7137,N_4208,N_4377);
nor U7138 (N_7138,N_4347,N_4512);
nand U7139 (N_7139,N_2638,N_4441);
nand U7140 (N_7140,N_3420,N_4323);
nor U7141 (N_7141,N_3930,N_3629);
xor U7142 (N_7142,N_3369,N_4730);
and U7143 (N_7143,N_2953,N_3293);
nor U7144 (N_7144,N_3417,N_2542);
and U7145 (N_7145,N_3903,N_3324);
or U7146 (N_7146,N_4277,N_3744);
xor U7147 (N_7147,N_2678,N_3540);
nand U7148 (N_7148,N_3642,N_4873);
nand U7149 (N_7149,N_4066,N_3824);
and U7150 (N_7150,N_3074,N_4131);
or U7151 (N_7151,N_3451,N_4585);
nand U7152 (N_7152,N_3675,N_4912);
and U7153 (N_7153,N_3361,N_4586);
or U7154 (N_7154,N_4040,N_4107);
or U7155 (N_7155,N_3034,N_3768);
and U7156 (N_7156,N_3480,N_4878);
and U7157 (N_7157,N_4524,N_4111);
nor U7158 (N_7158,N_4579,N_2904);
or U7159 (N_7159,N_3672,N_3220);
or U7160 (N_7160,N_3237,N_2981);
nor U7161 (N_7161,N_4237,N_4344);
or U7162 (N_7162,N_4536,N_3991);
nand U7163 (N_7163,N_4863,N_2997);
and U7164 (N_7164,N_4971,N_3924);
nor U7165 (N_7165,N_4046,N_3093);
nand U7166 (N_7166,N_3445,N_4349);
and U7167 (N_7167,N_4828,N_3012);
nor U7168 (N_7168,N_3478,N_2514);
or U7169 (N_7169,N_4117,N_3661);
nand U7170 (N_7170,N_3311,N_3391);
nor U7171 (N_7171,N_4203,N_4178);
nor U7172 (N_7172,N_3080,N_4481);
xor U7173 (N_7173,N_3530,N_2956);
or U7174 (N_7174,N_4392,N_3684);
or U7175 (N_7175,N_2724,N_4947);
nand U7176 (N_7176,N_3859,N_3536);
nand U7177 (N_7177,N_4137,N_3338);
nor U7178 (N_7178,N_3040,N_2839);
nand U7179 (N_7179,N_4309,N_4189);
and U7180 (N_7180,N_4038,N_3430);
and U7181 (N_7181,N_2593,N_3107);
xnor U7182 (N_7182,N_4949,N_2638);
xnor U7183 (N_7183,N_3595,N_3378);
nand U7184 (N_7184,N_4734,N_4360);
and U7185 (N_7185,N_4363,N_2511);
nor U7186 (N_7186,N_3263,N_2978);
nand U7187 (N_7187,N_4423,N_3726);
nor U7188 (N_7188,N_3180,N_3347);
or U7189 (N_7189,N_4238,N_3882);
and U7190 (N_7190,N_2943,N_2510);
and U7191 (N_7191,N_4377,N_3831);
and U7192 (N_7192,N_3282,N_3336);
and U7193 (N_7193,N_2906,N_4391);
nand U7194 (N_7194,N_3451,N_4643);
or U7195 (N_7195,N_4462,N_3617);
nand U7196 (N_7196,N_2548,N_2726);
nor U7197 (N_7197,N_2966,N_2845);
or U7198 (N_7198,N_3624,N_3478);
nor U7199 (N_7199,N_4600,N_4526);
nor U7200 (N_7200,N_2939,N_4294);
nor U7201 (N_7201,N_3928,N_3974);
nor U7202 (N_7202,N_2951,N_3379);
xor U7203 (N_7203,N_2836,N_3244);
or U7204 (N_7204,N_3341,N_4150);
and U7205 (N_7205,N_2993,N_4454);
and U7206 (N_7206,N_2578,N_2593);
or U7207 (N_7207,N_4770,N_3869);
nor U7208 (N_7208,N_4438,N_4127);
and U7209 (N_7209,N_4945,N_3731);
and U7210 (N_7210,N_3205,N_4696);
or U7211 (N_7211,N_2551,N_3339);
nor U7212 (N_7212,N_4801,N_3750);
nor U7213 (N_7213,N_4754,N_2666);
or U7214 (N_7214,N_2526,N_3452);
nand U7215 (N_7215,N_4792,N_4523);
and U7216 (N_7216,N_4000,N_3443);
nand U7217 (N_7217,N_3785,N_3665);
nand U7218 (N_7218,N_4178,N_3998);
or U7219 (N_7219,N_3444,N_3129);
or U7220 (N_7220,N_3119,N_4305);
nand U7221 (N_7221,N_2771,N_4034);
nor U7222 (N_7222,N_4747,N_4621);
nand U7223 (N_7223,N_2542,N_2979);
or U7224 (N_7224,N_2920,N_3259);
nor U7225 (N_7225,N_4720,N_3778);
nor U7226 (N_7226,N_3845,N_4642);
nor U7227 (N_7227,N_3076,N_2862);
nor U7228 (N_7228,N_2726,N_3475);
and U7229 (N_7229,N_3456,N_4063);
nor U7230 (N_7230,N_3281,N_3872);
or U7231 (N_7231,N_3509,N_3875);
xor U7232 (N_7232,N_3908,N_2600);
nand U7233 (N_7233,N_2500,N_3452);
and U7234 (N_7234,N_4552,N_3380);
or U7235 (N_7235,N_4479,N_3700);
nand U7236 (N_7236,N_4554,N_3223);
and U7237 (N_7237,N_4738,N_4223);
xor U7238 (N_7238,N_3084,N_3403);
or U7239 (N_7239,N_3588,N_2860);
or U7240 (N_7240,N_4367,N_4459);
nand U7241 (N_7241,N_3930,N_3996);
xor U7242 (N_7242,N_2527,N_4147);
nor U7243 (N_7243,N_2960,N_3152);
and U7244 (N_7244,N_3936,N_3918);
nor U7245 (N_7245,N_4349,N_4470);
nand U7246 (N_7246,N_4992,N_4689);
or U7247 (N_7247,N_2675,N_4258);
nor U7248 (N_7248,N_2559,N_3779);
or U7249 (N_7249,N_4432,N_4870);
or U7250 (N_7250,N_2500,N_2806);
nand U7251 (N_7251,N_4501,N_4697);
nor U7252 (N_7252,N_2563,N_4053);
nor U7253 (N_7253,N_3853,N_4840);
nand U7254 (N_7254,N_3460,N_3379);
or U7255 (N_7255,N_4877,N_4793);
nor U7256 (N_7256,N_2849,N_3815);
and U7257 (N_7257,N_3681,N_2620);
nor U7258 (N_7258,N_4433,N_3619);
nor U7259 (N_7259,N_4469,N_3853);
nand U7260 (N_7260,N_3334,N_4195);
nor U7261 (N_7261,N_4698,N_3646);
and U7262 (N_7262,N_2917,N_4995);
nor U7263 (N_7263,N_2513,N_3232);
and U7264 (N_7264,N_3095,N_4881);
xnor U7265 (N_7265,N_3540,N_4527);
nor U7266 (N_7266,N_4215,N_3408);
or U7267 (N_7267,N_2826,N_2847);
nor U7268 (N_7268,N_2899,N_4147);
nand U7269 (N_7269,N_3377,N_2578);
and U7270 (N_7270,N_4542,N_3487);
nand U7271 (N_7271,N_4866,N_4416);
or U7272 (N_7272,N_3219,N_2865);
and U7273 (N_7273,N_3002,N_2577);
nand U7274 (N_7274,N_2896,N_4759);
nand U7275 (N_7275,N_4103,N_4406);
nor U7276 (N_7276,N_3743,N_4090);
nor U7277 (N_7277,N_4420,N_4317);
nor U7278 (N_7278,N_3620,N_4628);
nand U7279 (N_7279,N_3112,N_4275);
nand U7280 (N_7280,N_4775,N_3172);
nor U7281 (N_7281,N_3637,N_2790);
and U7282 (N_7282,N_2761,N_3016);
nand U7283 (N_7283,N_4712,N_3548);
nor U7284 (N_7284,N_3486,N_3793);
or U7285 (N_7285,N_2731,N_4300);
or U7286 (N_7286,N_4103,N_2736);
nor U7287 (N_7287,N_4566,N_4227);
or U7288 (N_7288,N_4542,N_3312);
nand U7289 (N_7289,N_4493,N_4219);
nor U7290 (N_7290,N_2819,N_3418);
xor U7291 (N_7291,N_4698,N_2582);
and U7292 (N_7292,N_3117,N_3637);
and U7293 (N_7293,N_2536,N_3025);
xor U7294 (N_7294,N_4967,N_3746);
nor U7295 (N_7295,N_3890,N_3424);
nand U7296 (N_7296,N_2942,N_3216);
and U7297 (N_7297,N_3796,N_3770);
nand U7298 (N_7298,N_2565,N_4695);
and U7299 (N_7299,N_4588,N_2541);
nand U7300 (N_7300,N_4713,N_2910);
xor U7301 (N_7301,N_4939,N_3905);
nand U7302 (N_7302,N_4812,N_4506);
or U7303 (N_7303,N_4146,N_4450);
xor U7304 (N_7304,N_4289,N_3549);
xor U7305 (N_7305,N_3166,N_2817);
or U7306 (N_7306,N_2892,N_4296);
or U7307 (N_7307,N_4026,N_3701);
and U7308 (N_7308,N_3939,N_3646);
nor U7309 (N_7309,N_4019,N_4158);
nor U7310 (N_7310,N_4991,N_2939);
or U7311 (N_7311,N_2713,N_3560);
nand U7312 (N_7312,N_3268,N_4483);
and U7313 (N_7313,N_3367,N_4894);
or U7314 (N_7314,N_3096,N_3016);
and U7315 (N_7315,N_4048,N_3188);
nand U7316 (N_7316,N_4142,N_4285);
nor U7317 (N_7317,N_2824,N_2940);
xnor U7318 (N_7318,N_4468,N_3435);
and U7319 (N_7319,N_3564,N_2931);
and U7320 (N_7320,N_4409,N_3343);
nand U7321 (N_7321,N_4539,N_3382);
nand U7322 (N_7322,N_4281,N_4048);
nand U7323 (N_7323,N_3655,N_3389);
and U7324 (N_7324,N_3075,N_3921);
and U7325 (N_7325,N_2684,N_3299);
nor U7326 (N_7326,N_2863,N_3033);
or U7327 (N_7327,N_4178,N_2669);
and U7328 (N_7328,N_3709,N_4314);
nand U7329 (N_7329,N_4962,N_3648);
or U7330 (N_7330,N_4426,N_3072);
xnor U7331 (N_7331,N_3063,N_2778);
nand U7332 (N_7332,N_2583,N_4940);
and U7333 (N_7333,N_4898,N_4163);
nand U7334 (N_7334,N_4393,N_3251);
or U7335 (N_7335,N_3581,N_4496);
xnor U7336 (N_7336,N_4585,N_3923);
and U7337 (N_7337,N_4875,N_4762);
xor U7338 (N_7338,N_2584,N_2924);
nor U7339 (N_7339,N_4032,N_2715);
xnor U7340 (N_7340,N_2807,N_3689);
nor U7341 (N_7341,N_3110,N_3615);
nand U7342 (N_7342,N_4573,N_3582);
nand U7343 (N_7343,N_3659,N_2721);
and U7344 (N_7344,N_3771,N_2657);
nand U7345 (N_7345,N_3521,N_3835);
and U7346 (N_7346,N_4767,N_2578);
nor U7347 (N_7347,N_4336,N_3254);
or U7348 (N_7348,N_4243,N_3896);
and U7349 (N_7349,N_4930,N_3955);
nand U7350 (N_7350,N_2880,N_2760);
nand U7351 (N_7351,N_4861,N_4936);
nor U7352 (N_7352,N_3090,N_4879);
or U7353 (N_7353,N_4930,N_4457);
or U7354 (N_7354,N_3366,N_3428);
or U7355 (N_7355,N_4958,N_4481);
xor U7356 (N_7356,N_2730,N_4307);
and U7357 (N_7357,N_3606,N_2959);
nand U7358 (N_7358,N_4965,N_4884);
or U7359 (N_7359,N_3809,N_2801);
and U7360 (N_7360,N_3544,N_4239);
nor U7361 (N_7361,N_2559,N_2638);
xnor U7362 (N_7362,N_2776,N_3653);
or U7363 (N_7363,N_4651,N_3305);
nand U7364 (N_7364,N_2571,N_3177);
nor U7365 (N_7365,N_3521,N_2858);
nand U7366 (N_7366,N_4962,N_3773);
or U7367 (N_7367,N_3133,N_4695);
or U7368 (N_7368,N_2596,N_3675);
and U7369 (N_7369,N_2672,N_3159);
xor U7370 (N_7370,N_3623,N_4982);
nor U7371 (N_7371,N_3123,N_3709);
or U7372 (N_7372,N_3617,N_4708);
and U7373 (N_7373,N_3668,N_3779);
or U7374 (N_7374,N_2505,N_3029);
or U7375 (N_7375,N_4162,N_3872);
nand U7376 (N_7376,N_3122,N_2887);
nor U7377 (N_7377,N_4055,N_4731);
and U7378 (N_7378,N_4563,N_3527);
and U7379 (N_7379,N_3573,N_4833);
or U7380 (N_7380,N_4321,N_2659);
nand U7381 (N_7381,N_4495,N_2662);
and U7382 (N_7382,N_2867,N_3172);
or U7383 (N_7383,N_4780,N_3401);
nor U7384 (N_7384,N_3248,N_3209);
nor U7385 (N_7385,N_4170,N_2988);
xor U7386 (N_7386,N_3968,N_4754);
or U7387 (N_7387,N_3226,N_4070);
and U7388 (N_7388,N_3084,N_4742);
or U7389 (N_7389,N_3659,N_4913);
nor U7390 (N_7390,N_3538,N_4313);
nor U7391 (N_7391,N_3634,N_3915);
and U7392 (N_7392,N_2541,N_4804);
nor U7393 (N_7393,N_3686,N_4702);
and U7394 (N_7394,N_4003,N_2708);
nor U7395 (N_7395,N_3945,N_2566);
nand U7396 (N_7396,N_2864,N_2657);
xnor U7397 (N_7397,N_3461,N_2638);
nand U7398 (N_7398,N_4427,N_2687);
nand U7399 (N_7399,N_4701,N_4352);
nor U7400 (N_7400,N_3309,N_2632);
nand U7401 (N_7401,N_4139,N_3924);
xor U7402 (N_7402,N_3039,N_2973);
nor U7403 (N_7403,N_3190,N_3134);
and U7404 (N_7404,N_4622,N_4814);
xor U7405 (N_7405,N_4547,N_4108);
and U7406 (N_7406,N_3096,N_4019);
and U7407 (N_7407,N_4173,N_3253);
nand U7408 (N_7408,N_4622,N_2914);
nor U7409 (N_7409,N_3790,N_3402);
nor U7410 (N_7410,N_4574,N_2857);
or U7411 (N_7411,N_4078,N_4218);
nor U7412 (N_7412,N_4480,N_2763);
and U7413 (N_7413,N_4269,N_4385);
nor U7414 (N_7414,N_4944,N_4494);
and U7415 (N_7415,N_4862,N_4311);
or U7416 (N_7416,N_3781,N_4974);
nor U7417 (N_7417,N_4993,N_4272);
xor U7418 (N_7418,N_3561,N_4688);
nand U7419 (N_7419,N_3362,N_4264);
and U7420 (N_7420,N_4330,N_4728);
nor U7421 (N_7421,N_4489,N_4899);
and U7422 (N_7422,N_4696,N_4536);
or U7423 (N_7423,N_2530,N_3323);
nand U7424 (N_7424,N_4429,N_4771);
or U7425 (N_7425,N_3271,N_2726);
or U7426 (N_7426,N_3973,N_3158);
nor U7427 (N_7427,N_3527,N_2580);
or U7428 (N_7428,N_4817,N_3739);
and U7429 (N_7429,N_4757,N_4122);
or U7430 (N_7430,N_3824,N_4569);
or U7431 (N_7431,N_4006,N_2561);
or U7432 (N_7432,N_4189,N_3711);
or U7433 (N_7433,N_4375,N_4121);
nand U7434 (N_7434,N_3147,N_2674);
and U7435 (N_7435,N_3603,N_4326);
or U7436 (N_7436,N_3994,N_3925);
or U7437 (N_7437,N_2929,N_3516);
nor U7438 (N_7438,N_3092,N_3342);
and U7439 (N_7439,N_2929,N_2735);
xnor U7440 (N_7440,N_4080,N_3089);
or U7441 (N_7441,N_3574,N_4938);
nor U7442 (N_7442,N_4192,N_4317);
nor U7443 (N_7443,N_4823,N_4632);
xnor U7444 (N_7444,N_4423,N_3836);
and U7445 (N_7445,N_3326,N_3365);
or U7446 (N_7446,N_3321,N_4501);
or U7447 (N_7447,N_2885,N_2639);
nor U7448 (N_7448,N_2532,N_2646);
xor U7449 (N_7449,N_3737,N_4988);
and U7450 (N_7450,N_4253,N_2550);
nor U7451 (N_7451,N_2685,N_4181);
nand U7452 (N_7452,N_3045,N_2983);
and U7453 (N_7453,N_4915,N_4896);
nand U7454 (N_7454,N_3896,N_3631);
nor U7455 (N_7455,N_3106,N_4831);
and U7456 (N_7456,N_3853,N_3848);
nand U7457 (N_7457,N_3566,N_3236);
or U7458 (N_7458,N_3937,N_2757);
or U7459 (N_7459,N_3995,N_4459);
and U7460 (N_7460,N_2636,N_3640);
nor U7461 (N_7461,N_4061,N_4729);
or U7462 (N_7462,N_3846,N_4263);
nand U7463 (N_7463,N_2863,N_3684);
and U7464 (N_7464,N_3388,N_4959);
nor U7465 (N_7465,N_4119,N_2647);
xnor U7466 (N_7466,N_4357,N_4536);
nand U7467 (N_7467,N_2683,N_2506);
nand U7468 (N_7468,N_3052,N_4177);
and U7469 (N_7469,N_2669,N_4867);
nor U7470 (N_7470,N_3377,N_2936);
nor U7471 (N_7471,N_4139,N_3099);
nand U7472 (N_7472,N_3182,N_3597);
nand U7473 (N_7473,N_2588,N_3295);
nand U7474 (N_7474,N_2824,N_3799);
xnor U7475 (N_7475,N_3145,N_4360);
nand U7476 (N_7476,N_4725,N_4167);
xor U7477 (N_7477,N_2924,N_3517);
nand U7478 (N_7478,N_3305,N_4256);
nand U7479 (N_7479,N_3763,N_2872);
xnor U7480 (N_7480,N_2974,N_2625);
or U7481 (N_7481,N_3999,N_3899);
and U7482 (N_7482,N_3722,N_3544);
nor U7483 (N_7483,N_4433,N_4139);
nand U7484 (N_7484,N_4678,N_2963);
or U7485 (N_7485,N_2527,N_4385);
and U7486 (N_7486,N_3134,N_4504);
nor U7487 (N_7487,N_4422,N_3801);
nand U7488 (N_7488,N_3338,N_2608);
nor U7489 (N_7489,N_3635,N_3583);
xor U7490 (N_7490,N_4073,N_3550);
and U7491 (N_7491,N_4159,N_4216);
or U7492 (N_7492,N_3205,N_4294);
and U7493 (N_7493,N_3626,N_3201);
or U7494 (N_7494,N_4083,N_2929);
or U7495 (N_7495,N_4282,N_2855);
or U7496 (N_7496,N_4112,N_3574);
nand U7497 (N_7497,N_2996,N_4506);
xnor U7498 (N_7498,N_3447,N_3928);
or U7499 (N_7499,N_4723,N_3477);
or U7500 (N_7500,N_5449,N_5303);
xor U7501 (N_7501,N_6998,N_6586);
and U7502 (N_7502,N_6888,N_5220);
and U7503 (N_7503,N_5556,N_5201);
and U7504 (N_7504,N_5121,N_6419);
and U7505 (N_7505,N_5743,N_5551);
or U7506 (N_7506,N_5787,N_6119);
nand U7507 (N_7507,N_5395,N_5529);
and U7508 (N_7508,N_6829,N_6861);
nand U7509 (N_7509,N_6818,N_6365);
nand U7510 (N_7510,N_7389,N_5465);
nor U7511 (N_7511,N_6088,N_7386);
nor U7512 (N_7512,N_7041,N_5888);
or U7513 (N_7513,N_7433,N_5625);
nand U7514 (N_7514,N_7240,N_6248);
and U7515 (N_7515,N_6504,N_6674);
and U7516 (N_7516,N_6233,N_6309);
nor U7517 (N_7517,N_5892,N_5213);
nor U7518 (N_7518,N_5536,N_6115);
nand U7519 (N_7519,N_6966,N_6354);
nor U7520 (N_7520,N_5764,N_5109);
or U7521 (N_7521,N_6681,N_7482);
nor U7522 (N_7522,N_5940,N_5247);
or U7523 (N_7523,N_7344,N_5950);
nand U7524 (N_7524,N_5023,N_6841);
nor U7525 (N_7525,N_6703,N_6587);
xnor U7526 (N_7526,N_5555,N_5917);
and U7527 (N_7527,N_5637,N_6224);
nand U7528 (N_7528,N_5511,N_5317);
nor U7529 (N_7529,N_6239,N_6024);
xor U7530 (N_7530,N_6219,N_5514);
or U7531 (N_7531,N_6759,N_7477);
nand U7532 (N_7532,N_5512,N_7276);
nor U7533 (N_7533,N_6750,N_7335);
and U7534 (N_7534,N_6550,N_7244);
xor U7535 (N_7535,N_7159,N_7225);
nor U7536 (N_7536,N_5645,N_7138);
or U7537 (N_7537,N_5991,N_6195);
and U7538 (N_7538,N_7031,N_5324);
xnor U7539 (N_7539,N_5834,N_5478);
nor U7540 (N_7540,N_7167,N_5338);
nand U7541 (N_7541,N_5945,N_7014);
nor U7542 (N_7542,N_6001,N_7391);
and U7543 (N_7543,N_6270,N_6461);
and U7544 (N_7544,N_6277,N_6178);
or U7545 (N_7545,N_5617,N_7088);
xor U7546 (N_7546,N_5158,N_6491);
nand U7547 (N_7547,N_5133,N_7498);
and U7548 (N_7548,N_6454,N_5733);
xor U7549 (N_7549,N_6907,N_5159);
and U7550 (N_7550,N_5634,N_5288);
or U7551 (N_7551,N_7122,N_6951);
or U7552 (N_7552,N_6968,N_6186);
nor U7553 (N_7553,N_6852,N_7441);
or U7554 (N_7554,N_5913,N_6325);
xor U7555 (N_7555,N_7497,N_6428);
xnor U7556 (N_7556,N_5624,N_5061);
nor U7557 (N_7557,N_5557,N_6409);
nor U7558 (N_7558,N_5243,N_6468);
and U7559 (N_7559,N_5662,N_5257);
or U7560 (N_7560,N_6211,N_6124);
nor U7561 (N_7561,N_5123,N_7094);
nor U7562 (N_7562,N_5573,N_5701);
nand U7563 (N_7563,N_6367,N_5825);
nor U7564 (N_7564,N_6009,N_5138);
and U7565 (N_7565,N_6886,N_5812);
and U7566 (N_7566,N_5521,N_5632);
nor U7567 (N_7567,N_5612,N_7395);
xor U7568 (N_7568,N_6305,N_5581);
nor U7569 (N_7569,N_5909,N_7376);
nand U7570 (N_7570,N_5673,N_5187);
nor U7571 (N_7571,N_6390,N_5763);
nor U7572 (N_7572,N_6081,N_5585);
or U7573 (N_7573,N_6474,N_7157);
and U7574 (N_7574,N_5746,N_7220);
nor U7575 (N_7575,N_5592,N_6969);
nand U7576 (N_7576,N_7355,N_5753);
nor U7577 (N_7577,N_5507,N_6819);
nor U7578 (N_7578,N_6971,N_5602);
and U7579 (N_7579,N_7221,N_6201);
and U7580 (N_7580,N_6440,N_7388);
nand U7581 (N_7581,N_6838,N_6007);
nor U7582 (N_7582,N_6286,N_5406);
nand U7583 (N_7583,N_6901,N_5480);
nand U7584 (N_7584,N_6814,N_6220);
or U7585 (N_7585,N_5530,N_6031);
or U7586 (N_7586,N_6486,N_6027);
nor U7587 (N_7587,N_5212,N_5941);
and U7588 (N_7588,N_6093,N_7362);
nor U7589 (N_7589,N_5967,N_7179);
and U7590 (N_7590,N_5304,N_5473);
nand U7591 (N_7591,N_6707,N_5327);
nand U7592 (N_7592,N_5183,N_7084);
or U7593 (N_7593,N_5630,N_6113);
nand U7594 (N_7594,N_6648,N_5112);
nor U7595 (N_7595,N_6417,N_5619);
nor U7596 (N_7596,N_6871,N_6231);
or U7597 (N_7597,N_7044,N_6931);
and U7598 (N_7598,N_5287,N_7439);
nand U7599 (N_7599,N_6036,N_6831);
nand U7600 (N_7600,N_6643,N_5914);
and U7601 (N_7601,N_5434,N_6222);
nor U7602 (N_7602,N_6216,N_5817);
nand U7603 (N_7603,N_6746,N_5208);
or U7604 (N_7604,N_5678,N_6920);
nand U7605 (N_7605,N_7004,N_6843);
and U7606 (N_7606,N_6565,N_5546);
nand U7607 (N_7607,N_6741,N_6539);
and U7608 (N_7608,N_6551,N_5777);
nand U7609 (N_7609,N_6116,N_5136);
nor U7610 (N_7610,N_5877,N_5562);
nor U7611 (N_7611,N_5587,N_5809);
nor U7612 (N_7612,N_6174,N_6257);
nor U7613 (N_7613,N_5631,N_6778);
and U7614 (N_7614,N_5452,N_5999);
and U7615 (N_7615,N_5383,N_5603);
nand U7616 (N_7616,N_5916,N_6061);
xnor U7617 (N_7617,N_5259,N_5608);
nand U7618 (N_7618,N_5609,N_5722);
nand U7619 (N_7619,N_6527,N_5902);
and U7620 (N_7620,N_6370,N_6312);
nor U7621 (N_7621,N_5938,N_5066);
nand U7622 (N_7622,N_6663,N_6092);
nand U7623 (N_7623,N_6884,N_5936);
and U7624 (N_7624,N_6709,N_6275);
or U7625 (N_7625,N_6290,N_5488);
xnor U7626 (N_7626,N_7414,N_6645);
nor U7627 (N_7627,N_7006,N_6531);
xor U7628 (N_7628,N_5225,N_6068);
and U7629 (N_7629,N_7491,N_6820);
and U7630 (N_7630,N_6157,N_5453);
xnor U7631 (N_7631,N_5593,N_6259);
and U7632 (N_7632,N_5696,N_5079);
nand U7633 (N_7633,N_6189,N_7351);
and U7634 (N_7634,N_5033,N_7374);
nand U7635 (N_7635,N_5508,N_5072);
and U7636 (N_7636,N_5717,N_7160);
or U7637 (N_7637,N_5790,N_7471);
or U7638 (N_7638,N_5709,N_7205);
xnor U7639 (N_7639,N_7375,N_5698);
and U7640 (N_7640,N_6604,N_6608);
or U7641 (N_7641,N_7163,N_6546);
or U7642 (N_7642,N_5328,N_5871);
nor U7643 (N_7643,N_5387,N_5782);
and U7644 (N_7644,N_7005,N_6481);
or U7645 (N_7645,N_5041,N_7145);
nand U7646 (N_7646,N_7449,N_7315);
or U7647 (N_7647,N_6251,N_7165);
or U7648 (N_7648,N_7270,N_6111);
and U7649 (N_7649,N_5081,N_5515);
and U7650 (N_7650,N_6324,N_6722);
nand U7651 (N_7651,N_7399,N_5052);
or U7652 (N_7652,N_5852,N_5160);
or U7653 (N_7653,N_6200,N_5348);
or U7654 (N_7654,N_5549,N_6571);
xor U7655 (N_7655,N_5318,N_6458);
xnor U7656 (N_7656,N_5830,N_7401);
nor U7657 (N_7657,N_5277,N_7464);
xnor U7658 (N_7658,N_5826,N_6077);
nor U7659 (N_7659,N_6577,N_5055);
and U7660 (N_7660,N_6994,N_5713);
nor U7661 (N_7661,N_5369,N_6471);
or U7662 (N_7662,N_5088,N_5657);
nand U7663 (N_7663,N_7275,N_6452);
nor U7664 (N_7664,N_7030,N_5627);
and U7665 (N_7665,N_6786,N_6755);
and U7666 (N_7666,N_7361,N_5036);
nand U7667 (N_7667,N_7092,N_5922);
or U7668 (N_7668,N_5102,N_7460);
or U7669 (N_7669,N_7372,N_6492);
nand U7670 (N_7670,N_6781,N_5094);
and U7671 (N_7671,N_5124,N_7332);
nand U7672 (N_7672,N_6505,N_5629);
or U7673 (N_7673,N_6134,N_6644);
nor U7674 (N_7674,N_5775,N_7484);
nor U7675 (N_7675,N_6448,N_5861);
and U7676 (N_7676,N_6387,N_6212);
nand U7677 (N_7677,N_7176,N_5498);
nand U7678 (N_7678,N_5975,N_5107);
nand U7679 (N_7679,N_6876,N_6521);
nor U7680 (N_7680,N_6840,N_5884);
and U7681 (N_7681,N_7095,N_7046);
nor U7682 (N_7682,N_5192,N_7191);
nor U7683 (N_7683,N_6084,N_6598);
and U7684 (N_7684,N_7305,N_5168);
nand U7685 (N_7685,N_6979,N_6334);
or U7686 (N_7686,N_6533,N_7429);
and U7687 (N_7687,N_5727,N_6333);
nand U7688 (N_7688,N_6184,N_6285);
nand U7689 (N_7689,N_7237,N_5312);
and U7690 (N_7690,N_7051,N_6183);
and U7691 (N_7691,N_6692,N_7082);
xnor U7692 (N_7692,N_6694,N_5525);
or U7693 (N_7693,N_6997,N_5228);
nor U7694 (N_7694,N_5814,N_5003);
xnor U7695 (N_7695,N_7173,N_6611);
or U7696 (N_7696,N_7017,N_7431);
nor U7697 (N_7697,N_6363,N_6427);
and U7698 (N_7698,N_6826,N_6617);
and U7699 (N_7699,N_6340,N_7156);
or U7700 (N_7700,N_5359,N_7271);
and U7701 (N_7701,N_5485,N_6097);
nor U7702 (N_7702,N_5650,N_7129);
nand U7703 (N_7703,N_6261,N_6637);
nor U7704 (N_7704,N_5930,N_6625);
nand U7705 (N_7705,N_5923,N_6105);
or U7706 (N_7706,N_6622,N_6804);
and U7707 (N_7707,N_5263,N_6591);
and U7708 (N_7708,N_7197,N_7164);
and U7709 (N_7709,N_5334,N_5151);
and U7710 (N_7710,N_7303,N_6272);
and U7711 (N_7711,N_6989,N_5035);
xnor U7712 (N_7712,N_6980,N_7474);
and U7713 (N_7713,N_5600,N_5886);
nand U7714 (N_7714,N_7309,N_6028);
nor U7715 (N_7715,N_5392,N_6131);
nor U7716 (N_7716,N_7069,N_6052);
xor U7717 (N_7717,N_6965,N_6837);
nor U7718 (N_7718,N_6519,N_5718);
nand U7719 (N_7719,N_5952,N_6535);
or U7720 (N_7720,N_5245,N_6815);
or U7721 (N_7721,N_6086,N_6547);
or U7722 (N_7722,N_6145,N_7187);
or U7723 (N_7723,N_6667,N_6213);
or U7724 (N_7724,N_7243,N_7152);
nor U7725 (N_7725,N_5011,N_5311);
xor U7726 (N_7726,N_5222,N_6520);
nor U7727 (N_7727,N_6055,N_5251);
or U7728 (N_7728,N_5497,N_6613);
and U7729 (N_7729,N_7003,N_7450);
nand U7730 (N_7730,N_5179,N_6624);
and U7731 (N_7731,N_6990,N_6580);
and U7732 (N_7732,N_6004,N_5043);
nor U7733 (N_7733,N_6863,N_5655);
or U7734 (N_7734,N_5726,N_7116);
nor U7735 (N_7735,N_5569,N_6266);
xnor U7736 (N_7736,N_7140,N_5391);
or U7737 (N_7737,N_5533,N_5248);
nand U7738 (N_7738,N_6881,N_5463);
and U7739 (N_7739,N_7043,N_6500);
nor U7740 (N_7740,N_7162,N_5792);
nand U7741 (N_7741,N_5297,N_5535);
nor U7742 (N_7742,N_6832,N_5065);
and U7743 (N_7743,N_5495,N_6414);
and U7744 (N_7744,N_5788,N_6972);
and U7745 (N_7745,N_6364,N_5882);
nand U7746 (N_7746,N_6894,N_5682);
or U7747 (N_7747,N_7045,N_5844);
nor U7748 (N_7748,N_7473,N_6745);
and U7749 (N_7749,N_7048,N_5227);
xor U7750 (N_7750,N_6293,N_5474);
nor U7751 (N_7751,N_7128,N_6225);
nand U7752 (N_7752,N_6721,N_5797);
xor U7753 (N_7753,N_5751,N_6583);
nand U7754 (N_7754,N_7462,N_5887);
nor U7755 (N_7755,N_5358,N_6715);
nand U7756 (N_7756,N_5542,N_5928);
nor U7757 (N_7757,N_7396,N_5146);
or U7758 (N_7758,N_5695,N_7324);
or U7759 (N_7759,N_7207,N_5221);
nand U7760 (N_7760,N_6317,N_5719);
or U7761 (N_7761,N_5699,N_6646);
nand U7762 (N_7762,N_5931,N_6949);
or U7763 (N_7763,N_6592,N_6253);
and U7764 (N_7764,N_5260,N_5493);
or U7765 (N_7765,N_6264,N_7360);
nand U7766 (N_7766,N_6540,N_6789);
xnor U7767 (N_7767,N_6469,N_5336);
and U7768 (N_7768,N_5639,N_6988);
or U7769 (N_7769,N_6371,N_6695);
xor U7770 (N_7770,N_7104,N_5070);
nor U7771 (N_7771,N_5285,N_6017);
nor U7772 (N_7772,N_5450,N_7049);
nand U7773 (N_7773,N_5870,N_6857);
xor U7774 (N_7774,N_7480,N_6782);
or U7775 (N_7775,N_6545,N_6210);
nor U7776 (N_7776,N_6612,N_6763);
nor U7777 (N_7777,N_6512,N_5660);
and U7778 (N_7778,N_7468,N_6634);
xnor U7779 (N_7779,N_6537,N_6578);
and U7780 (N_7780,N_5837,N_7255);
nand U7781 (N_7781,N_5890,N_7019);
nor U7782 (N_7782,N_6449,N_5527);
or U7783 (N_7783,N_5807,N_7228);
and U7784 (N_7784,N_7298,N_7203);
or U7785 (N_7785,N_6342,N_5537);
and U7786 (N_7786,N_5607,N_6557);
nand U7787 (N_7787,N_6574,N_6214);
or U7788 (N_7788,N_6725,N_6146);
and U7789 (N_7789,N_6380,N_5795);
and U7790 (N_7790,N_6553,N_5781);
xor U7791 (N_7791,N_6572,N_6422);
nor U7792 (N_7792,N_5357,N_5086);
xnor U7793 (N_7793,N_6102,N_6660);
nor U7794 (N_7794,N_5953,N_5396);
nor U7795 (N_7795,N_7039,N_6176);
nand U7796 (N_7796,N_7108,N_6675);
and U7797 (N_7797,N_5910,N_5961);
nor U7798 (N_7798,N_6022,N_5134);
or U7799 (N_7799,N_6062,N_5700);
and U7800 (N_7800,N_6398,N_7445);
or U7801 (N_7801,N_6615,N_6006);
or U7802 (N_7802,N_6875,N_5606);
or U7803 (N_7803,N_6172,N_7231);
nand U7804 (N_7804,N_5860,N_7264);
or U7805 (N_7805,N_6824,N_6727);
and U7806 (N_7806,N_7209,N_6747);
and U7807 (N_7807,N_5436,N_6262);
xnor U7808 (N_7808,N_7064,N_6784);
nor U7809 (N_7809,N_6602,N_7423);
and U7810 (N_7810,N_6835,N_5659);
xnor U7811 (N_7811,N_6700,N_6138);
and U7812 (N_7812,N_5768,N_7210);
or U7813 (N_7813,N_6827,N_5433);
nand U7814 (N_7814,N_5957,N_6299);
or U7815 (N_7815,N_5640,N_6327);
or U7816 (N_7816,N_5972,N_6282);
nand U7817 (N_7817,N_6166,N_7115);
nand U7818 (N_7818,N_6069,N_7133);
and U7819 (N_7819,N_5808,N_7118);
xor U7820 (N_7820,N_5059,N_6160);
and U7821 (N_7821,N_6271,N_6588);
or U7822 (N_7822,N_6447,N_7025);
and U7823 (N_7823,N_7038,N_6839);
nor U7824 (N_7824,N_5728,N_7499);
or U7825 (N_7825,N_6227,N_5597);
xnor U7826 (N_7826,N_6352,N_5572);
nand U7827 (N_7827,N_6767,N_7214);
or U7828 (N_7828,N_6283,N_7348);
and U7829 (N_7829,N_6413,N_5095);
and U7830 (N_7830,N_5210,N_6985);
or U7831 (N_7831,N_6952,N_5832);
nand U7832 (N_7832,N_6064,N_5841);
nor U7833 (N_7833,N_5946,N_5779);
xnor U7834 (N_7834,N_6435,N_6025);
or U7835 (N_7835,N_5384,N_5987);
xor U7836 (N_7836,N_5758,N_6517);
xor U7837 (N_7837,N_5415,N_7254);
and U7838 (N_7838,N_6381,N_5738);
nand U7839 (N_7839,N_5705,N_5047);
and U7840 (N_7840,N_5419,N_5564);
and U7841 (N_7841,N_5496,N_7454);
and U7842 (N_7842,N_5979,N_6281);
and U7843 (N_7843,N_6744,N_6676);
nand U7844 (N_7844,N_7341,N_7387);
and U7845 (N_7845,N_5799,N_5320);
and U7846 (N_7846,N_6476,N_5918);
or U7847 (N_7847,N_6473,N_6331);
and U7848 (N_7848,N_5191,N_6029);
and U7849 (N_7849,N_6045,N_5866);
and U7850 (N_7850,N_6743,N_5706);
and U7851 (N_7851,N_5424,N_5897);
or U7852 (N_7852,N_6267,N_5708);
or U7853 (N_7853,N_6601,N_6459);
or U7854 (N_7854,N_5520,N_5855);
or U7855 (N_7855,N_7493,N_6834);
xnor U7856 (N_7856,N_6563,N_5256);
nor U7857 (N_7857,N_7483,N_6377);
and U7858 (N_7858,N_5538,N_5739);
or U7859 (N_7859,N_6800,N_7380);
and U7860 (N_7860,N_5420,N_5017);
xor U7861 (N_7861,N_5876,N_5981);
nor U7862 (N_7862,N_7068,N_7343);
nor U7863 (N_7863,N_6658,N_5091);
and U7864 (N_7864,N_6696,N_7416);
and U7865 (N_7865,N_5435,N_7060);
nor U7866 (N_7866,N_6947,N_5195);
xnor U7867 (N_7867,N_5407,N_6654);
xor U7868 (N_7868,N_5301,N_5883);
nor U7869 (N_7869,N_5128,N_7170);
nor U7870 (N_7870,N_5621,N_6833);
or U7871 (N_7871,N_5197,N_5813);
or U7872 (N_7872,N_6892,N_5547);
and U7873 (N_7873,N_7093,N_5749);
and U7874 (N_7874,N_6221,N_7475);
nand U7875 (N_7875,N_6430,N_7071);
and U7876 (N_7876,N_5667,N_5594);
nand U7877 (N_7877,N_7251,N_5176);
and U7878 (N_7878,N_5315,N_6698);
and U7879 (N_7879,N_6925,N_6629);
nand U7880 (N_7880,N_7397,N_7438);
nand U7881 (N_7881,N_7467,N_5087);
nor U7882 (N_7882,N_5644,N_7404);
or U7883 (N_7883,N_5702,N_5429);
xor U7884 (N_7884,N_5058,N_5704);
xnor U7885 (N_7885,N_6974,N_6005);
nand U7886 (N_7886,N_6651,N_5255);
xnor U7887 (N_7887,N_5494,N_6347);
nand U7888 (N_7888,N_6339,N_5867);
nor U7889 (N_7889,N_5170,N_5375);
nand U7890 (N_7890,N_7317,N_6810);
and U7891 (N_7891,N_6918,N_5769);
or U7892 (N_7892,N_5097,N_6549);
and U7893 (N_7893,N_7457,N_7065);
or U7894 (N_7894,N_5729,N_6493);
or U7895 (N_7895,N_5589,N_6133);
or U7896 (N_7896,N_7072,N_6590);
nand U7897 (N_7897,N_5413,N_6243);
or U7898 (N_7898,N_5292,N_5691);
and U7899 (N_7899,N_5074,N_6060);
nor U7900 (N_7900,N_7201,N_7268);
and U7901 (N_7901,N_5965,N_6489);
xor U7902 (N_7902,N_6234,N_5130);
nor U7903 (N_7903,N_6074,N_7059);
nor U7904 (N_7904,N_5380,N_6295);
or U7905 (N_7905,N_5155,N_7009);
or U7906 (N_7906,N_7453,N_5692);
nand U7907 (N_7907,N_6779,N_6171);
nor U7908 (N_7908,N_5754,N_5284);
and U7909 (N_7909,N_6292,N_6796);
or U7910 (N_7910,N_5075,N_7121);
or U7911 (N_7911,N_5671,N_6962);
and U7912 (N_7912,N_5161,N_7110);
nand U7913 (N_7913,N_6899,N_7472);
nand U7914 (N_7914,N_7393,N_7008);
nand U7915 (N_7915,N_6506,N_6666);
nor U7916 (N_7916,N_6359,N_5446);
xor U7917 (N_7917,N_7223,N_6065);
xor U7918 (N_7918,N_5985,N_6867);
nor U7919 (N_7919,N_5492,N_7266);
and U7920 (N_7920,N_5641,N_6067);
or U7921 (N_7921,N_7026,N_5177);
and U7922 (N_7922,N_5188,N_6177);
nor U7923 (N_7923,N_5934,N_6467);
nor U7924 (N_7924,N_6303,N_7451);
and U7925 (N_7925,N_5522,N_5426);
or U7926 (N_7926,N_6627,N_7249);
nand U7927 (N_7927,N_7291,N_5793);
xor U7928 (N_7928,N_7142,N_6360);
nor U7929 (N_7929,N_5165,N_5686);
and U7930 (N_7930,N_7289,N_7461);
nand U7931 (N_7931,N_6460,N_6085);
nor U7932 (N_7932,N_5580,N_6850);
and U7933 (N_7933,N_5716,N_5531);
nor U7934 (N_7934,N_6923,N_7137);
nand U7935 (N_7935,N_6165,N_7378);
and U7936 (N_7936,N_7333,N_5150);
nor U7937 (N_7937,N_6559,N_6155);
nand U7938 (N_7938,N_7089,N_6101);
nand U7939 (N_7939,N_6144,N_5185);
and U7940 (N_7940,N_5044,N_6768);
or U7941 (N_7941,N_7306,N_7269);
or U7942 (N_7942,N_6669,N_6358);
or U7943 (N_7943,N_5172,N_5281);
and U7944 (N_7944,N_7224,N_5805);
and U7945 (N_7945,N_5076,N_6967);
or U7946 (N_7946,N_5561,N_5783);
nand U7947 (N_7947,N_5982,N_6689);
and U7948 (N_7948,N_7417,N_7486);
nand U7949 (N_7949,N_6016,N_6465);
xor U7950 (N_7950,N_6532,N_6683);
or U7951 (N_7951,N_6154,N_6349);
nor U7952 (N_7952,N_7234,N_7434);
xnor U7953 (N_7953,N_5878,N_6185);
nor U7954 (N_7954,N_5926,N_7111);
and U7955 (N_7955,N_6245,N_5924);
nand U7956 (N_7956,N_5835,N_6066);
and U7957 (N_7957,N_7284,N_6730);
nor U7958 (N_7958,N_6401,N_6437);
or U7959 (N_7959,N_6418,N_7313);
and U7960 (N_7960,N_5008,N_7412);
and U7961 (N_7961,N_7148,N_6987);
or U7962 (N_7962,N_6156,N_5163);
and U7963 (N_7963,N_5374,N_7123);
or U7964 (N_7964,N_5481,N_5850);
xor U7965 (N_7965,N_5741,N_5652);
or U7966 (N_7966,N_5845,N_5675);
or U7967 (N_7967,N_7382,N_6063);
or U7968 (N_7968,N_5037,N_6652);
xnor U7969 (N_7969,N_6020,N_5857);
xor U7970 (N_7970,N_6127,N_6953);
and U7971 (N_7971,N_6374,N_6330);
xor U7972 (N_7972,N_7358,N_5326);
nand U7973 (N_7973,N_7370,N_7010);
xor U7974 (N_7974,N_5623,N_6208);
and U7975 (N_7975,N_5500,N_6255);
and U7976 (N_7976,N_5563,N_5270);
and U7977 (N_7977,N_5765,N_6773);
nor U7978 (N_7978,N_5186,N_6217);
nor U7979 (N_7979,N_5995,N_6050);
nand U7980 (N_7980,N_5162,N_6671);
nand U7981 (N_7981,N_5411,N_5274);
nand U7982 (N_7982,N_7310,N_7099);
and U7983 (N_7983,N_6599,N_6526);
and U7984 (N_7984,N_5214,N_6351);
and U7985 (N_7985,N_6596,N_5794);
nand U7986 (N_7986,N_5278,N_7297);
nor U7987 (N_7987,N_5252,N_6302);
xnor U7988 (N_7988,N_7184,N_6335);
nand U7989 (N_7989,N_5929,N_6441);
nor U7990 (N_7990,N_7192,N_6868);
and U7991 (N_7991,N_5977,N_6757);
and U7992 (N_7992,N_6003,N_5353);
and U7993 (N_7993,N_5875,N_5108);
nor U7994 (N_7994,N_6935,N_6830);
nor U7995 (N_7995,N_5989,N_6203);
nor U7996 (N_7996,N_5745,N_6793);
or U7997 (N_7997,N_5448,N_6860);
and U7998 (N_7998,N_6278,N_5120);
nand U7999 (N_7999,N_6566,N_6497);
xnor U8000 (N_8000,N_5622,N_7288);
xnor U8001 (N_8001,N_7394,N_5819);
nor U8002 (N_8002,N_5966,N_6909);
nand U8003 (N_8003,N_6691,N_5014);
nor U8004 (N_8004,N_5171,N_7427);
nand U8005 (N_8005,N_6724,N_5628);
nand U8006 (N_8006,N_6083,N_6938);
xor U8007 (N_8007,N_6107,N_5073);
nor U8008 (N_8008,N_6382,N_7021);
or U8009 (N_8009,N_5275,N_6737);
or U8010 (N_8010,N_5042,N_5444);
nand U8011 (N_8011,N_7435,N_7035);
nor U8012 (N_8012,N_6753,N_7458);
xor U8013 (N_8013,N_7345,N_5129);
and U8014 (N_8014,N_6341,N_6880);
or U8015 (N_8015,N_5239,N_6276);
and U8016 (N_8016,N_7469,N_5648);
and U8017 (N_8017,N_5296,N_5862);
or U8018 (N_8018,N_5670,N_5026);
or U8019 (N_8019,N_5544,N_6879);
or U8020 (N_8020,N_6790,N_6343);
nor U8021 (N_8021,N_6589,N_5601);
nor U8022 (N_8022,N_7114,N_6114);
and U8023 (N_8023,N_6670,N_5021);
nor U8024 (N_8024,N_6776,N_6291);
or U8025 (N_8025,N_5636,N_5665);
and U8026 (N_8026,N_7286,N_7217);
nor U8027 (N_8027,N_7101,N_5703);
nand U8028 (N_8028,N_6405,N_6424);
or U8029 (N_8029,N_5235,N_6568);
xor U8030 (N_8030,N_5955,N_7081);
or U8031 (N_8031,N_6668,N_7202);
or U8032 (N_8032,N_5962,N_5445);
and U8033 (N_8033,N_5683,N_7096);
or U8034 (N_8034,N_6581,N_6916);
xnor U8035 (N_8035,N_5103,N_5092);
nand U8036 (N_8036,N_6560,N_5299);
nor U8037 (N_8037,N_7367,N_7278);
nand U8038 (N_8038,N_7196,N_6564);
xnor U8039 (N_8039,N_6164,N_5119);
and U8040 (N_8040,N_6326,N_6915);
nand U8041 (N_8041,N_5410,N_5828);
and U8042 (N_8042,N_5291,N_7215);
and U8043 (N_8043,N_7230,N_5182);
and U8044 (N_8044,N_6487,N_5237);
and U8045 (N_8045,N_5140,N_7347);
xnor U8046 (N_8046,N_6848,N_5829);
nand U8047 (N_8047,N_6813,N_6693);
or U8048 (N_8048,N_6429,N_6758);
or U8049 (N_8049,N_6582,N_7027);
nor U8050 (N_8050,N_6684,N_5626);
nand U8051 (N_8051,N_5258,N_5401);
or U8052 (N_8052,N_5352,N_6508);
nor U8053 (N_8053,N_7144,N_7149);
nor U8054 (N_8054,N_6269,N_7037);
nand U8055 (N_8055,N_5230,N_5441);
nand U8056 (N_8056,N_7040,N_5541);
or U8057 (N_8057,N_5344,N_6181);
nand U8058 (N_8058,N_6190,N_5135);
or U8059 (N_8059,N_5174,N_6525);
nand U8060 (N_8060,N_6209,N_6472);
and U8061 (N_8061,N_6656,N_5490);
and U8062 (N_8062,N_5646,N_6263);
or U8063 (N_8063,N_5534,N_6393);
or U8064 (N_8064,N_6984,N_5774);
xnor U8065 (N_8065,N_5851,N_5893);
nand U8066 (N_8066,N_6021,N_7316);
nand U8067 (N_8067,N_7222,N_6548);
or U8068 (N_8068,N_5018,N_5202);
or U8069 (N_8069,N_6182,N_6797);
nand U8070 (N_8070,N_6389,N_6463);
and U8071 (N_8071,N_7001,N_6847);
or U8072 (N_8072,N_6456,N_6284);
nor U8073 (N_8073,N_6619,N_6950);
nand U8074 (N_8074,N_5935,N_7011);
nor U8075 (N_8075,N_7036,N_6618);
or U8076 (N_8076,N_5757,N_6958);
nor U8077 (N_8077,N_6237,N_6502);
nor U8078 (N_8078,N_7075,N_6760);
nand U8079 (N_8079,N_6432,N_6388);
nor U8080 (N_8080,N_7314,N_5313);
or U8081 (N_8081,N_5154,N_5838);
or U8082 (N_8082,N_6594,N_7055);
xor U8083 (N_8083,N_7319,N_5149);
or U8084 (N_8084,N_5685,N_6117);
or U8085 (N_8085,N_5020,N_5001);
nand U8086 (N_8086,N_6908,N_5152);
and U8087 (N_8087,N_5679,N_6704);
and U8088 (N_8088,N_7161,N_6169);
nand U8089 (N_8089,N_6911,N_6956);
nand U8090 (N_8090,N_5464,N_5462);
nand U8091 (N_8091,N_5164,N_6632);
nand U8092 (N_8092,N_5175,N_7371);
and U8093 (N_8093,N_5471,N_5385);
and U8094 (N_8094,N_5894,N_7481);
xor U8095 (N_8095,N_5681,N_6844);
xor U8096 (N_8096,N_5853,N_5049);
nor U8097 (N_8097,N_6412,N_5314);
nor U8098 (N_8098,N_5933,N_7253);
and U8099 (N_8099,N_5246,N_5205);
and U8100 (N_8100,N_6408,N_5901);
nor U8101 (N_8101,N_6774,N_5101);
nor U8102 (N_8102,N_6123,N_5360);
nand U8103 (N_8103,N_5048,N_5340);
nor U8104 (N_8104,N_6082,N_5064);
or U8105 (N_8105,N_5083,N_7226);
and U8106 (N_8106,N_6955,N_5577);
or U8107 (N_8107,N_5242,N_5596);
and U8108 (N_8108,N_6788,N_5578);
nand U8109 (N_8109,N_5856,N_5265);
nor U8110 (N_8110,N_6173,N_5004);
nand U8111 (N_8111,N_5944,N_5132);
xnor U8112 (N_8112,N_6569,N_6954);
nand U8113 (N_8113,N_7273,N_6957);
or U8114 (N_8114,N_6103,N_5651);
nor U8115 (N_8115,N_5976,N_6900);
or U8116 (N_8116,N_5071,N_6887);
or U8117 (N_8117,N_6087,N_6982);
nand U8118 (N_8118,N_6136,N_5649);
and U8119 (N_8119,N_6049,N_5863);
or U8120 (N_8120,N_6620,N_6976);
or U8121 (N_8121,N_6012,N_5068);
and U8122 (N_8122,N_6230,N_7090);
or U8123 (N_8123,N_6945,N_6436);
and U8124 (N_8124,N_6803,N_5145);
xnor U8125 (N_8125,N_6775,N_5077);
nand U8126 (N_8126,N_6687,N_7301);
nor U8127 (N_8127,N_6672,N_6623);
nor U8128 (N_8128,N_6148,N_7024);
nor U8129 (N_8129,N_6902,N_7331);
or U8130 (N_8130,N_5664,N_5379);
nor U8131 (N_8131,N_7079,N_5219);
xor U8132 (N_8132,N_7377,N_7419);
and U8133 (N_8133,N_7368,N_7147);
nor U8134 (N_8134,N_7153,N_6927);
nand U8135 (N_8135,N_7247,N_5971);
xor U8136 (N_8136,N_7119,N_7091);
and U8137 (N_8137,N_6159,N_6242);
nand U8138 (N_8138,N_7195,N_6917);
xnor U8139 (N_8139,N_6708,N_5847);
or U8140 (N_8140,N_5811,N_6391);
xnor U8141 (N_8141,N_5421,N_7076);
or U8142 (N_8142,N_6610,N_6070);
nand U8143 (N_8143,N_7403,N_6034);
nor U8144 (N_8144,N_5349,N_5199);
nand U8145 (N_8145,N_5427,N_7489);
nand U8146 (N_8146,N_5181,N_6498);
nor U8147 (N_8147,N_5082,N_6090);
and U8148 (N_8148,N_5365,N_5414);
nand U8149 (N_8149,N_5206,N_5229);
or U8150 (N_8150,N_6718,N_6094);
or U8151 (N_8151,N_7238,N_6978);
nor U8152 (N_8152,N_5404,N_6313);
nand U8153 (N_8153,N_7109,N_7352);
xnor U8154 (N_8154,N_5968,N_6320);
nor U8155 (N_8155,N_6193,N_5381);
nor U8156 (N_8156,N_5920,N_5139);
nor U8157 (N_8157,N_7052,N_6073);
nor U8158 (N_8158,N_6575,N_7029);
and U8159 (N_8159,N_5791,N_5467);
nor U8160 (N_8160,N_7175,N_7302);
or U8161 (N_8161,N_6051,N_5428);
or U8162 (N_8162,N_6605,N_6207);
nor U8163 (N_8163,N_7402,N_6192);
and U8164 (N_8164,N_6319,N_5309);
or U8165 (N_8165,N_5361,N_6685);
nand U8166 (N_8166,N_6510,N_6383);
nand U8167 (N_8167,N_6891,N_5725);
nor U8168 (N_8168,N_7151,N_6883);
nand U8169 (N_8169,N_7290,N_5342);
and U8170 (N_8170,N_5865,N_5653);
or U8171 (N_8171,N_6350,N_5316);
or U8172 (N_8172,N_5399,N_6163);
nand U8173 (N_8173,N_6806,N_6930);
and U8174 (N_8174,N_5822,N_7105);
or U8175 (N_8175,N_5282,N_6453);
nor U8176 (N_8176,N_5254,N_5499);
nor U8177 (N_8177,N_5919,N_5057);
or U8178 (N_8178,N_5815,N_6897);
and U8179 (N_8179,N_7256,N_6158);
xnor U8180 (N_8180,N_6959,N_5800);
and U8181 (N_8181,N_7330,N_5050);
nor U8182 (N_8182,N_6141,N_7337);
nand U8183 (N_8183,N_5438,N_5661);
or U8184 (N_8184,N_6348,N_7182);
or U8185 (N_8185,N_6742,N_6026);
or U8186 (N_8186,N_6849,N_7086);
nor U8187 (N_8187,N_5302,N_5579);
or U8188 (N_8188,N_6121,N_5233);
nor U8189 (N_8189,N_7356,N_5022);
nand U8190 (N_8190,N_7185,N_6431);
and U8191 (N_8191,N_6726,N_5509);
and U8192 (N_8192,N_7465,N_6442);
and U8193 (N_8193,N_6287,N_7425);
nor U8194 (N_8194,N_6948,N_6033);
nand U8195 (N_8195,N_6764,N_7373);
and U8196 (N_8196,N_6011,N_6934);
nand U8197 (N_8197,N_5545,N_6010);
nand U8198 (N_8198,N_5350,N_7312);
and U8199 (N_8199,N_6096,N_6922);
xor U8200 (N_8200,N_6756,N_5234);
nand U8201 (N_8201,N_6944,N_7443);
nand U8202 (N_8202,N_5761,N_6630);
and U8203 (N_8203,N_7420,N_5802);
nand U8204 (N_8204,N_5460,N_7390);
and U8205 (N_8205,N_5289,N_7180);
or U8206 (N_8206,N_7177,N_6332);
nand U8207 (N_8207,N_7357,N_6478);
nor U8208 (N_8208,N_5211,N_6480);
or U8209 (N_8209,N_5431,N_6426);
xnor U8210 (N_8210,N_5322,N_5105);
and U8211 (N_8211,N_6379,N_5039);
or U8212 (N_8212,N_5540,N_6080);
xor U8213 (N_8213,N_6058,N_5409);
nor U8214 (N_8214,N_7318,N_5780);
nor U8215 (N_8215,N_5598,N_5457);
or U8216 (N_8216,N_6866,N_7078);
and U8217 (N_8217,N_5240,N_6023);
and U8218 (N_8218,N_6904,N_5784);
xnor U8219 (N_8219,N_6072,N_6162);
or U8220 (N_8220,N_5742,N_6318);
nor U8221 (N_8221,N_5030,N_6226);
or U8222 (N_8222,N_5006,N_5543);
and U8223 (N_8223,N_5824,N_6609);
and U8224 (N_8224,N_7311,N_5859);
nor U8225 (N_8225,N_5568,N_5595);
or U8226 (N_8226,N_5759,N_6541);
or U8227 (N_8227,N_5153,N_5298);
or U8228 (N_8228,N_5687,N_5519);
nand U8229 (N_8229,N_6002,N_5785);
and U8230 (N_8230,N_6496,N_6232);
or U8231 (N_8231,N_5843,N_7229);
nand U8232 (N_8232,N_5748,N_7248);
nand U8233 (N_8233,N_6483,N_5200);
or U8234 (N_8234,N_6640,N_6384);
or U8235 (N_8235,N_5267,N_6273);
or U8236 (N_8236,N_5455,N_5466);
and U8237 (N_8237,N_6905,N_5013);
nor U8238 (N_8238,N_6842,N_7350);
or U8239 (N_8239,N_6723,N_5680);
and U8240 (N_8240,N_7213,N_6252);
nand U8241 (N_8241,N_5998,N_6822);
nand U8242 (N_8242,N_6933,N_6823);
or U8243 (N_8243,N_6731,N_6941);
nand U8244 (N_8244,N_5874,N_6853);
nor U8245 (N_8245,N_6122,N_5367);
nor U8246 (N_8246,N_5707,N_6522);
nor U8247 (N_8247,N_5333,N_5548);
nand U8248 (N_8248,N_6872,N_7325);
and U8249 (N_8249,N_6037,N_6665);
nand U8250 (N_8250,N_5080,N_5276);
nand U8251 (N_8251,N_5960,N_5858);
or U8252 (N_8252,N_6929,N_6752);
nor U8253 (N_8253,N_6846,N_5907);
nor U8254 (N_8254,N_6368,N_5915);
xor U8255 (N_8255,N_6518,N_7136);
or U8256 (N_8256,N_6135,N_5654);
nor U8257 (N_8257,N_6129,N_6639);
nand U8258 (N_8258,N_5550,N_5416);
nor U8259 (N_8259,N_7428,N_6614);
and U8260 (N_8260,N_6128,N_5148);
nand U8261 (N_8261,N_6878,N_6109);
and U8262 (N_8262,N_6153,N_5341);
and U8263 (N_8263,N_6893,N_6095);
and U8264 (N_8264,N_6812,N_7418);
or U8265 (N_8265,N_6205,N_5911);
or U8266 (N_8266,N_6986,N_7424);
xnor U8267 (N_8267,N_6336,N_6711);
and U8268 (N_8268,N_6805,N_5294);
nand U8269 (N_8269,N_6919,N_6828);
nor U8270 (N_8270,N_6659,N_7018);
or U8271 (N_8271,N_5300,N_5377);
nor U8272 (N_8272,N_7100,N_5106);
nor U8273 (N_8273,N_5347,N_5881);
nor U8274 (N_8274,N_6898,N_6018);
or U8275 (N_8275,N_7134,N_7020);
nand U8276 (N_8276,N_6714,N_6678);
nor U8277 (N_8277,N_6633,N_5710);
nand U8278 (N_8278,N_6112,N_7208);
or U8279 (N_8279,N_6981,N_5051);
or U8280 (N_8280,N_6964,N_6528);
or U8281 (N_8281,N_6104,N_5586);
nor U8282 (N_8282,N_6536,N_5231);
xor U8283 (N_8283,N_5190,N_5329);
xor U8284 (N_8284,N_7295,N_5351);
and U8285 (N_8285,N_6762,N_5283);
xor U8286 (N_8286,N_5677,N_5127);
or U8287 (N_8287,N_5224,N_5560);
or U8288 (N_8288,N_5458,N_5854);
and U8289 (N_8289,N_5459,N_6250);
nor U8290 (N_8290,N_6120,N_5203);
nand U8291 (N_8291,N_6098,N_5356);
xnor U8292 (N_8292,N_5178,N_6626);
xor U8293 (N_8293,N_6228,N_7383);
or U8294 (N_8294,N_5386,N_5635);
or U8295 (N_8295,N_6555,N_5332);
xnor U8296 (N_8296,N_6375,N_7479);
or U8297 (N_8297,N_5002,N_5207);
and U8298 (N_8298,N_7308,N_5423);
or U8299 (N_8299,N_5354,N_5261);
or U8300 (N_8300,N_5939,N_6597);
nand U8301 (N_8301,N_6877,N_6513);
nand U8302 (N_8302,N_6035,N_5672);
nand U8303 (N_8303,N_6301,N_5417);
nor U8304 (N_8304,N_6785,N_5479);
and U8305 (N_8305,N_6362,N_6256);
or U8306 (N_8306,N_5089,N_5475);
or U8307 (N_8307,N_7171,N_5032);
and U8308 (N_8308,N_5715,N_7321);
and U8309 (N_8309,N_5062,N_5262);
xor U8310 (N_8310,N_5778,N_6777);
nor U8311 (N_8311,N_6046,N_6748);
and U8312 (N_8312,N_5712,N_6438);
or U8313 (N_8313,N_5552,N_5618);
and U8314 (N_8314,N_5988,N_6507);
or U8315 (N_8315,N_6197,N_5959);
nor U8316 (N_8316,N_5721,N_6139);
or U8317 (N_8317,N_6279,N_6740);
and U8318 (N_8318,N_6932,N_6446);
nand U8319 (N_8319,N_6701,N_7279);
or U8320 (N_8320,N_7061,N_6043);
nor U8321 (N_8321,N_6825,N_5997);
nor U8322 (N_8322,N_7283,N_5576);
or U8323 (N_8323,N_5482,N_5308);
and U8324 (N_8324,N_5046,N_5319);
xnor U8325 (N_8325,N_7392,N_5370);
nor U8326 (N_8326,N_6690,N_5566);
nor U8327 (N_8327,N_6013,N_5189);
or U8328 (N_8328,N_6514,N_7463);
nand U8329 (N_8329,N_6770,N_6196);
nor U8330 (N_8330,N_7227,N_5908);
or U8331 (N_8331,N_7053,N_7466);
nor U8332 (N_8332,N_6561,N_6353);
or U8333 (N_8333,N_6247,N_5925);
nand U8334 (N_8334,N_6859,N_6729);
nand U8335 (N_8335,N_7456,N_5840);
nor U8336 (N_8336,N_7280,N_6421);
or U8337 (N_8337,N_5842,N_5400);
nand U8338 (N_8338,N_7204,N_5253);
nor U8339 (N_8339,N_6712,N_6053);
nand U8340 (N_8340,N_6631,N_7354);
or U8341 (N_8341,N_5921,N_6874);
or U8342 (N_8342,N_6399,N_5388);
nor U8343 (N_8343,N_5504,N_7262);
or U8344 (N_8344,N_6673,N_5293);
nor U8345 (N_8345,N_6167,N_5964);
nand U8346 (N_8346,N_7206,N_6821);
nor U8347 (N_8347,N_7112,N_6600);
and U8348 (N_8348,N_6444,N_5232);
nor U8349 (N_8349,N_6089,N_6130);
nor U8350 (N_8350,N_5517,N_7232);
or U8351 (N_8351,N_7246,N_5196);
nand U8352 (N_8352,N_5000,N_7168);
and U8353 (N_8353,N_5582,N_6056);
and U8354 (N_8354,N_6355,N_6862);
or U8355 (N_8355,N_5054,N_6960);
and U8356 (N_8356,N_6771,N_6791);
nor U8357 (N_8357,N_5583,N_6057);
or U8358 (N_8358,N_5099,N_5373);
nor U8359 (N_8359,N_7346,N_7385);
nor U8360 (N_8360,N_6406,N_6484);
or U8361 (N_8361,N_7143,N_5331);
and U8362 (N_8362,N_5216,N_5970);
and U8363 (N_8363,N_5118,N_7032);
nor U8364 (N_8364,N_6143,N_6856);
nor U8365 (N_8365,N_7113,N_5905);
xnor U8366 (N_8366,N_5034,N_6315);
or U8367 (N_8367,N_7085,N_5025);
or U8368 (N_8368,N_6059,N_6751);
and U8369 (N_8369,N_7353,N_5472);
xnor U8370 (N_8370,N_7259,N_5831);
xnor U8371 (N_8371,N_7250,N_6511);
or U8372 (N_8372,N_5836,N_5873);
or U8373 (N_8373,N_5484,N_5752);
or U8374 (N_8374,N_5364,N_5193);
or U8375 (N_8375,N_6882,N_6524);
and U8376 (N_8376,N_5900,N_6316);
or U8377 (N_8377,N_6635,N_6584);
xor U8378 (N_8378,N_6161,N_7292);
or U8379 (N_8379,N_5590,N_5010);
or U8380 (N_8380,N_5376,N_7496);
xor U8381 (N_8381,N_6543,N_6366);
or U8382 (N_8382,N_5827,N_5408);
nor U8383 (N_8383,N_7260,N_7257);
nand U8384 (N_8384,N_5223,N_7432);
nand U8385 (N_8385,N_5218,N_6792);
nor U8386 (N_8386,N_6765,N_6662);
or U8387 (N_8387,N_7074,N_5085);
nand U8388 (N_8388,N_7296,N_6042);
and U8389 (N_8389,N_7107,N_7359);
xnor U8390 (N_8390,N_5669,N_6699);
nor U8391 (N_8391,N_5969,N_6455);
or U8392 (N_8392,N_5943,N_7409);
xnor U8393 (N_8393,N_6928,N_5801);
xor U8394 (N_8394,N_7124,N_6030);
and U8395 (N_8395,N_6556,N_5040);
xor U8396 (N_8396,N_7323,N_7186);
and U8397 (N_8397,N_5539,N_5771);
nand U8398 (N_8398,N_6274,N_7028);
nor U8399 (N_8399,N_6585,N_6246);
and U8400 (N_8400,N_6495,N_7141);
nor U8401 (N_8401,N_7442,N_6501);
or U8402 (N_8402,N_7062,N_5833);
nor U8403 (N_8403,N_7400,N_6118);
or U8404 (N_8404,N_6705,N_6268);
or U8405 (N_8405,N_6038,N_5806);
nand U8406 (N_8406,N_7277,N_6530);
nand U8407 (N_8407,N_7421,N_6152);
xor U8408 (N_8408,N_5390,N_5732);
and U8409 (N_8409,N_7379,N_6308);
nand U8410 (N_8410,N_7130,N_7073);
and U8411 (N_8411,N_6204,N_5038);
or U8412 (N_8412,N_5236,N_7307);
nand U8413 (N_8413,N_7169,N_7369);
nor U8414 (N_8414,N_5904,N_5849);
and U8415 (N_8415,N_5864,N_5658);
nor U8416 (N_8416,N_7405,N_5372);
nand U8417 (N_8417,N_5440,N_6783);
nand U8418 (N_8418,N_7272,N_6706);
nor U8419 (N_8419,N_5614,N_6260);
nand U8420 (N_8420,N_7042,N_6345);
or U8421 (N_8421,N_6329,N_6870);
and U8422 (N_8422,N_5770,N_6235);
xnor U8423 (N_8423,N_5528,N_5767);
nor U8424 (N_8424,N_6180,N_6720);
and U8425 (N_8425,N_5244,N_5575);
or U8426 (N_8426,N_7336,N_5570);
nor U8427 (N_8427,N_6297,N_7166);
xnor U8428 (N_8428,N_5776,N_5616);
or U8429 (N_8429,N_5378,N_7188);
xnor U8430 (N_8430,N_5456,N_5558);
nor U8431 (N_8431,N_7022,N_5786);
nor U8432 (N_8432,N_5060,N_6795);
and U8433 (N_8433,N_7282,N_6215);
and U8434 (N_8434,N_7194,N_5734);
or U8435 (N_8435,N_6562,N_5804);
nand U8436 (N_8436,N_5306,N_6423);
nand U8437 (N_8437,N_5009,N_5005);
nand U8438 (N_8438,N_5345,N_7245);
xor U8439 (N_8439,N_5821,N_6811);
nand U8440 (N_8440,N_5280,N_7448);
xor U8441 (N_8441,N_5869,N_6855);
nand U8442 (N_8442,N_5523,N_6710);
nor U8443 (N_8443,N_6236,N_7364);
nand U8444 (N_8444,N_7365,N_5116);
nor U8445 (N_8445,N_6150,N_6677);
and U8446 (N_8446,N_6403,N_7447);
nor U8447 (N_8447,N_5157,N_6937);
nor U8448 (N_8448,N_6048,N_5947);
xor U8449 (N_8449,N_7063,N_5167);
nor U8450 (N_8450,N_5412,N_6479);
nor U8451 (N_8451,N_7219,N_5454);
nor U8452 (N_8452,N_6126,N_5402);
nor U8453 (N_8453,N_6337,N_6780);
xnor U8454 (N_8454,N_5553,N_5565);
nand U8455 (N_8455,N_5215,N_6628);
or U8456 (N_8456,N_5588,N_6249);
nor U8457 (N_8457,N_7077,N_5425);
xnor U8458 (N_8458,N_6047,N_6218);
nand U8459 (N_8459,N_5393,N_5984);
nand U8460 (N_8460,N_7410,N_6697);
or U8461 (N_8461,N_5891,N_7328);
nor U8462 (N_8462,N_6996,N_5643);
nand U8463 (N_8463,N_5468,N_6924);
and U8464 (N_8464,N_6132,N_7407);
or U8465 (N_8465,N_5397,N_5194);
nand U8466 (N_8466,N_5803,N_5605);
nor U8467 (N_8467,N_5430,N_6682);
and U8468 (N_8468,N_5295,N_7102);
nand U8469 (N_8469,N_5974,N_5736);
and U8470 (N_8470,N_6702,N_5740);
and U8471 (N_8471,N_5007,N_5980);
nor U8472 (N_8472,N_5756,N_5335);
nor U8473 (N_8473,N_7150,N_5773);
or U8474 (N_8474,N_6992,N_6451);
xor U8475 (N_8475,N_5279,N_6344);
and U8476 (N_8476,N_5028,N_7106);
nor U8477 (N_8477,N_5737,N_6534);
nor U8478 (N_8478,N_6558,N_6869);
nand U8479 (N_8479,N_7047,N_6910);
or U8480 (N_8480,N_5518,N_6995);
nor U8481 (N_8481,N_5620,N_7125);
xor U8482 (N_8482,N_6392,N_6433);
xnor U8483 (N_8483,N_6450,N_7320);
xor U8484 (N_8484,N_6386,N_5184);
and U8485 (N_8485,N_6416,N_5217);
xor U8486 (N_8486,N_6607,N_5398);
or U8487 (N_8487,N_7193,N_6970);
nor U8488 (N_8488,N_6000,N_5986);
or U8489 (N_8489,N_6137,N_7437);
nand U8490 (N_8490,N_6199,N_7242);
nor U8491 (N_8491,N_6108,N_5330);
and U8492 (N_8492,N_5173,N_5355);
xnor U8493 (N_8493,N_6999,N_7155);
nand U8494 (N_8494,N_6490,N_6322);
and U8495 (N_8495,N_5491,N_5273);
xor U8496 (N_8496,N_6503,N_6889);
xnor U8497 (N_8497,N_6140,N_6688);
nor U8498 (N_8498,N_6921,N_6716);
and U8499 (N_8499,N_7015,N_5898);
or U8500 (N_8500,N_5647,N_7485);
or U8501 (N_8501,N_6961,N_5486);
nor U8502 (N_8502,N_6254,N_5983);
xor U8503 (N_8503,N_5615,N_6194);
nor U8504 (N_8504,N_5093,N_5432);
nand U8505 (N_8505,N_7070,N_5798);
nand U8506 (N_8506,N_6801,N_6686);
or U8507 (N_8507,N_6595,N_7183);
or U8508 (N_8508,N_6198,N_5470);
nand U8509 (N_8509,N_5405,N_5090);
and U8510 (N_8510,N_7300,N_6653);
or U8511 (N_8511,N_6523,N_5638);
nor U8512 (N_8512,N_7146,N_6914);
and U8513 (N_8513,N_6304,N_6238);
nand U8514 (N_8514,N_5027,N_5990);
or U8515 (N_8515,N_5656,N_5868);
nand U8516 (N_8516,N_6404,N_7239);
nand U8517 (N_8517,N_5180,N_5744);
or U8518 (N_8518,N_5599,N_6306);
xor U8519 (N_8519,N_6415,N_5418);
nand U8520 (N_8520,N_5321,N_7057);
and U8521 (N_8521,N_7436,N_6864);
or U8522 (N_8522,N_7198,N_5209);
nand U8523 (N_8523,N_7287,N_6397);
or U8524 (N_8524,N_6361,N_7000);
nand U8525 (N_8525,N_6499,N_6240);
and U8526 (N_8526,N_7252,N_7087);
nand U8527 (N_8527,N_7487,N_5249);
nor U8528 (N_8528,N_7050,N_7440);
nor U8529 (N_8529,N_5117,N_6661);
xnor U8530 (N_8530,N_5963,N_7274);
nand U8531 (N_8531,N_6044,N_5723);
nor U8532 (N_8532,N_5611,N_7381);
xor U8533 (N_8533,N_5343,N_7135);
and U8534 (N_8534,N_7398,N_6713);
nand U8535 (N_8535,N_7455,N_6079);
or U8536 (N_8536,N_7406,N_6940);
nand U8537 (N_8537,N_7430,N_5069);
and U8538 (N_8538,N_5731,N_5443);
or U8539 (N_8539,N_6187,N_7233);
nor U8540 (N_8540,N_7492,N_5506);
nor U8541 (N_8541,N_6395,N_7334);
nand U8542 (N_8542,N_5422,N_6509);
nand U8543 (N_8543,N_6188,N_7422);
nor U8544 (N_8544,N_6650,N_6032);
xor U8545 (N_8545,N_6772,N_6445);
and U8546 (N_8546,N_6369,N_5816);
or U8547 (N_8547,N_7098,N_5290);
nor U8548 (N_8548,N_6936,N_5442);
or U8549 (N_8549,N_5238,N_5056);
nand U8550 (N_8550,N_7103,N_5250);
nor U8551 (N_8551,N_7236,N_6054);
and U8552 (N_8552,N_5818,N_7363);
nand U8553 (N_8553,N_5142,N_5346);
xor U8554 (N_8554,N_6728,N_5571);
nand U8555 (N_8555,N_5879,N_5156);
nand U8556 (N_8556,N_6649,N_7329);
or U8557 (N_8557,N_5126,N_5899);
or U8558 (N_8558,N_6845,N_5147);
or U8559 (N_8559,N_6443,N_5169);
nor U8560 (N_8560,N_5226,N_7066);
or U8561 (N_8561,N_5954,N_6816);
and U8562 (N_8562,N_6977,N_5848);
and U8563 (N_8563,N_6655,N_7218);
or U8564 (N_8564,N_5690,N_5789);
or U8565 (N_8565,N_5016,N_5031);
nand U8566 (N_8566,N_6071,N_5362);
or U8567 (N_8567,N_6885,N_6621);
nor U8568 (N_8568,N_5389,N_5098);
nand U8569 (N_8569,N_6147,N_6394);
and U8570 (N_8570,N_7265,N_5689);
or U8571 (N_8571,N_6170,N_6019);
nor U8572 (N_8572,N_6396,N_5310);
nor U8573 (N_8573,N_5019,N_5325);
nand U8574 (N_8574,N_6638,N_5131);
or U8575 (N_8575,N_5469,N_6749);
or U8576 (N_8576,N_6078,N_5949);
and U8577 (N_8577,N_5015,N_7067);
xor U8578 (N_8578,N_7285,N_5810);
and U8579 (N_8579,N_5337,N_5477);
nor U8580 (N_8580,N_5730,N_6346);
or U8581 (N_8581,N_7490,N_7261);
nor U8582 (N_8582,N_7158,N_6457);
nand U8583 (N_8583,N_5144,N_6294);
and U8584 (N_8584,N_6142,N_6420);
and U8585 (N_8585,N_7258,N_6963);
and U8586 (N_8586,N_7459,N_5559);
xor U8587 (N_8587,N_6657,N_6616);
and U8588 (N_8588,N_5198,N_5889);
and U8589 (N_8589,N_6926,N_6943);
nor U8590 (N_8590,N_6373,N_6464);
xnor U8591 (N_8591,N_6485,N_6865);
and U8592 (N_8592,N_7200,N_6040);
nor U8593 (N_8593,N_5305,N_7154);
or U8594 (N_8594,N_5604,N_7494);
nand U8595 (N_8595,N_6206,N_5382);
nand U8596 (N_8596,N_5978,N_6895);
nor U8597 (N_8597,N_6179,N_7495);
and U8598 (N_8598,N_5711,N_5503);
and U8599 (N_8599,N_7181,N_6836);
nor U8600 (N_8600,N_6202,N_6946);
or U8601 (N_8601,N_6265,N_7216);
nor U8602 (N_8602,N_6149,N_5067);
nor U8603 (N_8603,N_5286,N_6151);
and U8604 (N_8604,N_6754,N_7294);
or U8605 (N_8605,N_6515,N_5554);
nand U8606 (N_8606,N_5932,N_6356);
nand U8607 (N_8607,N_5024,N_5676);
and U8608 (N_8608,N_6280,N_7408);
xnor U8609 (N_8609,N_7190,N_6975);
and U8610 (N_8610,N_6993,N_5724);
or U8611 (N_8611,N_7172,N_6175);
nor U8612 (N_8612,N_6738,N_5574);
xor U8613 (N_8613,N_5674,N_6376);
and U8614 (N_8614,N_5323,N_6794);
and U8615 (N_8615,N_5104,N_5668);
nor U8616 (N_8616,N_6494,N_6296);
nand U8617 (N_8617,N_7139,N_5958);
nor U8618 (N_8618,N_5307,N_7444);
xnor U8619 (N_8619,N_7327,N_7263);
or U8620 (N_8620,N_7488,N_5143);
or U8621 (N_8621,N_5750,N_5951);
or U8622 (N_8622,N_7120,N_7127);
or U8623 (N_8623,N_7476,N_5906);
and U8624 (N_8624,N_5204,N_6014);
or U8625 (N_8625,N_6890,N_5762);
xnor U8626 (N_8626,N_6357,N_5642);
or U8627 (N_8627,N_7007,N_5111);
and U8628 (N_8628,N_5264,N_5895);
nor U8629 (N_8629,N_6099,N_6439);
nor U8630 (N_8630,N_6873,N_5820);
or U8631 (N_8631,N_5693,N_7056);
nor U8632 (N_8632,N_7339,N_6809);
nand U8633 (N_8633,N_6407,N_6244);
or U8634 (N_8634,N_5012,N_6191);
nor U8635 (N_8635,N_6769,N_7054);
nor U8636 (N_8636,N_5633,N_5591);
nor U8637 (N_8637,N_5684,N_6462);
nor U8638 (N_8638,N_5368,N_6733);
and U8639 (N_8639,N_6466,N_6258);
and U8640 (N_8640,N_5122,N_5993);
nor U8641 (N_8641,N_6378,N_6679);
and U8642 (N_8642,N_5567,N_5487);
nor U8643 (N_8643,N_7002,N_7349);
xnor U8644 (N_8644,N_5613,N_5483);
nand U8645 (N_8645,N_6229,N_6576);
and U8646 (N_8646,N_5823,N_6554);
or U8647 (N_8647,N_7384,N_5942);
and U8648 (N_8648,N_6300,N_5927);
or U8649 (N_8649,N_6858,N_6732);
and U8650 (N_8650,N_7080,N_7131);
or U8651 (N_8651,N_6787,N_6425);
and U8652 (N_8652,N_5269,N_5973);
and U8653 (N_8653,N_5110,N_5839);
and U8654 (N_8654,N_6311,N_6125);
nor U8655 (N_8655,N_6896,N_6008);
nor U8656 (N_8656,N_6808,N_5271);
nand U8657 (N_8657,N_5084,N_7058);
nor U8658 (N_8658,N_6488,N_6321);
nand U8659 (N_8659,N_5437,N_6538);
and U8660 (N_8660,N_7034,N_6091);
nor U8661 (N_8661,N_5872,N_5760);
or U8662 (N_8662,N_5403,N_6647);
nor U8663 (N_8663,N_7013,N_6075);
nor U8664 (N_8664,N_7016,N_5524);
and U8665 (N_8665,N_6717,N_7023);
nand U8666 (N_8666,N_5755,N_6903);
and U8667 (N_8667,N_6851,N_6906);
nor U8668 (N_8668,N_6106,N_7097);
xor U8669 (N_8669,N_5476,N_6567);
nand U8670 (N_8670,N_6314,N_7338);
nand U8671 (N_8671,N_7470,N_6544);
xor U8672 (N_8672,N_6991,N_5584);
and U8673 (N_8673,N_6807,N_5266);
nor U8674 (N_8674,N_6168,N_7126);
or U8675 (N_8675,N_6798,N_6579);
xor U8676 (N_8676,N_5394,N_5697);
nand U8677 (N_8677,N_5688,N_6606);
and U8678 (N_8678,N_6912,N_7212);
and U8679 (N_8679,N_6939,N_7083);
xor U8680 (N_8680,N_6913,N_6734);
or U8681 (N_8681,N_5896,N_7178);
nand U8682 (N_8682,N_5846,N_5956);
and U8683 (N_8683,N_6470,N_5735);
nor U8684 (N_8684,N_5502,N_6642);
or U8685 (N_8685,N_6223,N_7322);
nor U8686 (N_8686,N_5610,N_7174);
nor U8687 (N_8687,N_7446,N_5510);
and U8688 (N_8688,N_5996,N_6983);
xnor U8689 (N_8689,N_6385,N_6400);
nor U8690 (N_8690,N_7299,N_6542);
and U8691 (N_8691,N_5505,N_6802);
nor U8692 (N_8692,N_7452,N_5666);
xor U8693 (N_8693,N_6041,N_5125);
nor U8694 (N_8694,N_5029,N_5937);
and U8695 (N_8695,N_7426,N_7293);
xnor U8696 (N_8696,N_5053,N_7342);
nand U8697 (N_8697,N_5526,N_6110);
nand U8698 (N_8698,N_6593,N_5912);
or U8699 (N_8699,N_5114,N_6310);
nor U8700 (N_8700,N_5439,N_6241);
and U8701 (N_8701,N_6328,N_5100);
and U8702 (N_8702,N_7235,N_5694);
or U8703 (N_8703,N_7132,N_5994);
and U8704 (N_8704,N_6817,N_5447);
nor U8705 (N_8705,N_5663,N_5115);
and U8706 (N_8706,N_5992,N_6410);
nor U8707 (N_8707,N_6039,N_5516);
nand U8708 (N_8708,N_7267,N_5078);
nor U8709 (N_8709,N_5339,N_6307);
and U8710 (N_8710,N_6799,N_6076);
and U8711 (N_8711,N_7415,N_5880);
and U8712 (N_8712,N_5948,N_5272);
nor U8713 (N_8713,N_6516,N_5371);
nor U8714 (N_8714,N_5489,N_6735);
or U8715 (N_8715,N_7304,N_6664);
xor U8716 (N_8716,N_5747,N_6636);
xnor U8717 (N_8717,N_6854,N_6100);
and U8718 (N_8718,N_7411,N_5096);
and U8719 (N_8719,N_6603,N_6288);
or U8720 (N_8720,N_6680,N_5513);
nor U8721 (N_8721,N_5363,N_7211);
and U8722 (N_8722,N_6015,N_5045);
nor U8723 (N_8723,N_5166,N_6411);
xnor U8724 (N_8724,N_7117,N_7281);
or U8725 (N_8725,N_5714,N_5141);
nor U8726 (N_8726,N_5113,N_5796);
nand U8727 (N_8727,N_6942,N_5241);
xor U8728 (N_8728,N_5532,N_6552);
or U8729 (N_8729,N_7413,N_6736);
or U8730 (N_8730,N_6298,N_6973);
or U8731 (N_8731,N_6482,N_7033);
nor U8732 (N_8732,N_5366,N_5885);
and U8733 (N_8733,N_5501,N_6402);
nand U8734 (N_8734,N_5772,N_6573);
or U8735 (N_8735,N_6570,N_7189);
and U8736 (N_8736,N_6719,N_6739);
nand U8737 (N_8737,N_7241,N_5137);
nand U8738 (N_8738,N_6434,N_7340);
nor U8739 (N_8739,N_5451,N_7012);
nand U8740 (N_8740,N_7199,N_6475);
and U8741 (N_8741,N_6323,N_6761);
and U8742 (N_8742,N_7366,N_5766);
and U8743 (N_8743,N_6766,N_6372);
nor U8744 (N_8744,N_6477,N_5268);
and U8745 (N_8745,N_7478,N_5461);
xor U8746 (N_8746,N_7326,N_5720);
nor U8747 (N_8747,N_5063,N_6289);
or U8748 (N_8748,N_6338,N_6641);
or U8749 (N_8749,N_5903,N_6529);
nor U8750 (N_8750,N_5556,N_5764);
and U8751 (N_8751,N_7321,N_5660);
and U8752 (N_8752,N_6209,N_6997);
or U8753 (N_8753,N_5123,N_5756);
nand U8754 (N_8754,N_5860,N_6372);
nor U8755 (N_8755,N_5646,N_5402);
nor U8756 (N_8756,N_6597,N_5204);
and U8757 (N_8757,N_5812,N_7467);
nor U8758 (N_8758,N_5960,N_6340);
and U8759 (N_8759,N_5693,N_5868);
nand U8760 (N_8760,N_7384,N_5152);
or U8761 (N_8761,N_5272,N_6376);
and U8762 (N_8762,N_5782,N_5403);
nor U8763 (N_8763,N_5683,N_6749);
or U8764 (N_8764,N_6075,N_6671);
or U8765 (N_8765,N_5528,N_5035);
nor U8766 (N_8766,N_7098,N_6025);
nor U8767 (N_8767,N_5598,N_7193);
nor U8768 (N_8768,N_7101,N_6086);
xnor U8769 (N_8769,N_5136,N_5239);
nand U8770 (N_8770,N_6598,N_5655);
and U8771 (N_8771,N_6740,N_5880);
xor U8772 (N_8772,N_5756,N_6596);
nor U8773 (N_8773,N_5940,N_5772);
nand U8774 (N_8774,N_7154,N_5092);
and U8775 (N_8775,N_5609,N_6614);
and U8776 (N_8776,N_6209,N_6021);
nor U8777 (N_8777,N_6881,N_6945);
or U8778 (N_8778,N_6461,N_6944);
and U8779 (N_8779,N_5670,N_6681);
nand U8780 (N_8780,N_5347,N_7433);
and U8781 (N_8781,N_7334,N_5964);
and U8782 (N_8782,N_6205,N_6966);
xor U8783 (N_8783,N_6233,N_6192);
nor U8784 (N_8784,N_7296,N_6326);
or U8785 (N_8785,N_5751,N_7421);
xor U8786 (N_8786,N_6553,N_5480);
and U8787 (N_8787,N_6553,N_6626);
xor U8788 (N_8788,N_7206,N_6011);
nand U8789 (N_8789,N_5217,N_5643);
and U8790 (N_8790,N_5573,N_7373);
and U8791 (N_8791,N_5670,N_5850);
nand U8792 (N_8792,N_6174,N_6629);
nor U8793 (N_8793,N_7368,N_5028);
or U8794 (N_8794,N_5321,N_7411);
nor U8795 (N_8795,N_5605,N_6938);
xnor U8796 (N_8796,N_5846,N_5157);
nand U8797 (N_8797,N_7203,N_5055);
nand U8798 (N_8798,N_7161,N_6565);
or U8799 (N_8799,N_6798,N_7238);
nand U8800 (N_8800,N_6343,N_5746);
and U8801 (N_8801,N_5256,N_5600);
or U8802 (N_8802,N_6449,N_7072);
or U8803 (N_8803,N_6719,N_6938);
nor U8804 (N_8804,N_6250,N_5709);
and U8805 (N_8805,N_5015,N_5478);
nand U8806 (N_8806,N_6658,N_7198);
xnor U8807 (N_8807,N_7312,N_5839);
nor U8808 (N_8808,N_7065,N_6233);
or U8809 (N_8809,N_6058,N_5698);
nand U8810 (N_8810,N_6318,N_5277);
nand U8811 (N_8811,N_5270,N_5037);
nor U8812 (N_8812,N_6084,N_6516);
nor U8813 (N_8813,N_6155,N_5591);
and U8814 (N_8814,N_6963,N_5803);
or U8815 (N_8815,N_6668,N_5433);
xor U8816 (N_8816,N_5336,N_5767);
or U8817 (N_8817,N_6715,N_5770);
nor U8818 (N_8818,N_6472,N_5588);
or U8819 (N_8819,N_5958,N_7020);
or U8820 (N_8820,N_7425,N_5015);
nand U8821 (N_8821,N_5837,N_6610);
nand U8822 (N_8822,N_6643,N_7172);
xnor U8823 (N_8823,N_6853,N_7372);
or U8824 (N_8824,N_7250,N_6181);
xnor U8825 (N_8825,N_5960,N_6179);
nand U8826 (N_8826,N_6469,N_7411);
xnor U8827 (N_8827,N_5364,N_6598);
and U8828 (N_8828,N_5295,N_5046);
nor U8829 (N_8829,N_5392,N_6799);
xor U8830 (N_8830,N_5392,N_6467);
and U8831 (N_8831,N_6293,N_6677);
nand U8832 (N_8832,N_6264,N_6379);
nor U8833 (N_8833,N_5103,N_6431);
nor U8834 (N_8834,N_7084,N_6035);
or U8835 (N_8835,N_6460,N_6049);
nor U8836 (N_8836,N_5452,N_6984);
nor U8837 (N_8837,N_5243,N_5893);
nand U8838 (N_8838,N_6598,N_5970);
or U8839 (N_8839,N_7076,N_5539);
and U8840 (N_8840,N_5383,N_7392);
or U8841 (N_8841,N_6297,N_5513);
and U8842 (N_8842,N_5835,N_5609);
nor U8843 (N_8843,N_5046,N_6997);
nor U8844 (N_8844,N_5844,N_5210);
and U8845 (N_8845,N_7421,N_6289);
nand U8846 (N_8846,N_6828,N_5236);
xor U8847 (N_8847,N_5135,N_5566);
and U8848 (N_8848,N_6554,N_6320);
nand U8849 (N_8849,N_6983,N_7136);
and U8850 (N_8850,N_6531,N_6458);
nor U8851 (N_8851,N_5084,N_5548);
nand U8852 (N_8852,N_7344,N_6497);
xnor U8853 (N_8853,N_5956,N_7327);
nor U8854 (N_8854,N_5401,N_5743);
and U8855 (N_8855,N_5748,N_7298);
nor U8856 (N_8856,N_7481,N_5582);
nand U8857 (N_8857,N_6036,N_6314);
nand U8858 (N_8858,N_6965,N_6072);
nor U8859 (N_8859,N_6287,N_7184);
nand U8860 (N_8860,N_6142,N_5959);
nor U8861 (N_8861,N_7216,N_6472);
nand U8862 (N_8862,N_5066,N_7012);
nand U8863 (N_8863,N_6904,N_6088);
and U8864 (N_8864,N_5377,N_5578);
and U8865 (N_8865,N_5140,N_5624);
nor U8866 (N_8866,N_7046,N_6531);
nand U8867 (N_8867,N_5555,N_6305);
and U8868 (N_8868,N_7114,N_6031);
nand U8869 (N_8869,N_5929,N_7040);
and U8870 (N_8870,N_5233,N_7229);
nor U8871 (N_8871,N_7267,N_6828);
nand U8872 (N_8872,N_7191,N_7322);
nand U8873 (N_8873,N_6305,N_5358);
xor U8874 (N_8874,N_6789,N_5427);
nor U8875 (N_8875,N_5768,N_6360);
nor U8876 (N_8876,N_6878,N_5067);
nor U8877 (N_8877,N_6683,N_5079);
nor U8878 (N_8878,N_7257,N_5910);
nor U8879 (N_8879,N_5423,N_7071);
or U8880 (N_8880,N_6468,N_5957);
or U8881 (N_8881,N_6261,N_6549);
nand U8882 (N_8882,N_7274,N_6929);
and U8883 (N_8883,N_6550,N_7272);
xnor U8884 (N_8884,N_6630,N_6513);
and U8885 (N_8885,N_5356,N_5220);
nand U8886 (N_8886,N_6365,N_5845);
or U8887 (N_8887,N_5308,N_6666);
xnor U8888 (N_8888,N_5393,N_5906);
and U8889 (N_8889,N_5053,N_6900);
and U8890 (N_8890,N_7467,N_6436);
or U8891 (N_8891,N_6172,N_5064);
nand U8892 (N_8892,N_5650,N_5889);
xor U8893 (N_8893,N_6425,N_7126);
nand U8894 (N_8894,N_6733,N_5225);
and U8895 (N_8895,N_5975,N_6537);
nand U8896 (N_8896,N_6974,N_5199);
and U8897 (N_8897,N_5534,N_5980);
nand U8898 (N_8898,N_5611,N_7323);
nand U8899 (N_8899,N_6396,N_5210);
and U8900 (N_8900,N_6417,N_5630);
nor U8901 (N_8901,N_5208,N_6836);
xor U8902 (N_8902,N_6647,N_6453);
nor U8903 (N_8903,N_5994,N_7350);
nand U8904 (N_8904,N_6903,N_5329);
or U8905 (N_8905,N_6561,N_6887);
nand U8906 (N_8906,N_5184,N_5768);
nand U8907 (N_8907,N_7399,N_5533);
xor U8908 (N_8908,N_6307,N_6224);
nand U8909 (N_8909,N_6887,N_6234);
nor U8910 (N_8910,N_7447,N_5115);
nor U8911 (N_8911,N_6576,N_6750);
nand U8912 (N_8912,N_6350,N_6890);
or U8913 (N_8913,N_7184,N_5486);
or U8914 (N_8914,N_5434,N_5194);
or U8915 (N_8915,N_7487,N_5221);
or U8916 (N_8916,N_6695,N_5301);
or U8917 (N_8917,N_5762,N_7155);
nand U8918 (N_8918,N_6619,N_7392);
nand U8919 (N_8919,N_6717,N_6165);
nor U8920 (N_8920,N_5828,N_6483);
nand U8921 (N_8921,N_6213,N_5031);
and U8922 (N_8922,N_7395,N_7237);
or U8923 (N_8923,N_6618,N_5127);
or U8924 (N_8924,N_5936,N_5565);
nand U8925 (N_8925,N_6035,N_5419);
nor U8926 (N_8926,N_6078,N_6979);
nand U8927 (N_8927,N_5100,N_6155);
nor U8928 (N_8928,N_7260,N_6888);
nand U8929 (N_8929,N_7046,N_6572);
and U8930 (N_8930,N_5089,N_7106);
nand U8931 (N_8931,N_5128,N_6251);
or U8932 (N_8932,N_6795,N_6946);
or U8933 (N_8933,N_7081,N_5585);
nor U8934 (N_8934,N_6870,N_5439);
xnor U8935 (N_8935,N_5207,N_5961);
or U8936 (N_8936,N_7256,N_6284);
nor U8937 (N_8937,N_6996,N_6918);
or U8938 (N_8938,N_6738,N_5754);
nor U8939 (N_8939,N_6435,N_6574);
nor U8940 (N_8940,N_7256,N_6665);
xor U8941 (N_8941,N_7444,N_6790);
nand U8942 (N_8942,N_6245,N_6889);
nand U8943 (N_8943,N_6701,N_7100);
nand U8944 (N_8944,N_6113,N_6048);
or U8945 (N_8945,N_5289,N_6187);
or U8946 (N_8946,N_7236,N_6430);
nand U8947 (N_8947,N_5294,N_5378);
nor U8948 (N_8948,N_7033,N_5879);
nor U8949 (N_8949,N_5347,N_6096);
nand U8950 (N_8950,N_5349,N_5764);
nand U8951 (N_8951,N_6272,N_7008);
or U8952 (N_8952,N_5058,N_6576);
nor U8953 (N_8953,N_6888,N_6192);
nand U8954 (N_8954,N_6291,N_5614);
and U8955 (N_8955,N_7366,N_6433);
or U8956 (N_8956,N_7164,N_5194);
xnor U8957 (N_8957,N_7459,N_7405);
or U8958 (N_8958,N_7324,N_6239);
and U8959 (N_8959,N_7072,N_6682);
and U8960 (N_8960,N_7279,N_7125);
or U8961 (N_8961,N_6985,N_6842);
and U8962 (N_8962,N_5481,N_6096);
nor U8963 (N_8963,N_5210,N_6603);
or U8964 (N_8964,N_5110,N_5307);
or U8965 (N_8965,N_6687,N_5855);
nand U8966 (N_8966,N_5549,N_7419);
nor U8967 (N_8967,N_5393,N_6779);
nor U8968 (N_8968,N_6708,N_6755);
or U8969 (N_8969,N_6803,N_6110);
nand U8970 (N_8970,N_5705,N_7151);
xor U8971 (N_8971,N_7456,N_5584);
nor U8972 (N_8972,N_6352,N_5170);
nand U8973 (N_8973,N_5103,N_5248);
or U8974 (N_8974,N_7187,N_6214);
and U8975 (N_8975,N_6664,N_7186);
nand U8976 (N_8976,N_7283,N_5567);
and U8977 (N_8977,N_6425,N_6264);
xnor U8978 (N_8978,N_6785,N_6494);
or U8979 (N_8979,N_5312,N_5535);
nand U8980 (N_8980,N_6642,N_7146);
nand U8981 (N_8981,N_6619,N_6154);
nand U8982 (N_8982,N_7198,N_6716);
nor U8983 (N_8983,N_6320,N_6747);
and U8984 (N_8984,N_6779,N_6619);
nor U8985 (N_8985,N_6600,N_6570);
nor U8986 (N_8986,N_6201,N_6583);
nand U8987 (N_8987,N_6201,N_5719);
and U8988 (N_8988,N_6165,N_5479);
or U8989 (N_8989,N_5541,N_5015);
and U8990 (N_8990,N_6778,N_5858);
xnor U8991 (N_8991,N_5791,N_5441);
and U8992 (N_8992,N_7496,N_5791);
nor U8993 (N_8993,N_5731,N_5696);
or U8994 (N_8994,N_5720,N_6871);
or U8995 (N_8995,N_6441,N_6899);
or U8996 (N_8996,N_5183,N_5316);
xor U8997 (N_8997,N_5458,N_7365);
and U8998 (N_8998,N_5248,N_6302);
and U8999 (N_8999,N_5815,N_5491);
nand U9000 (N_9000,N_5839,N_6472);
nor U9001 (N_9001,N_5440,N_7097);
and U9002 (N_9002,N_7410,N_5886);
or U9003 (N_9003,N_5776,N_5005);
xnor U9004 (N_9004,N_5696,N_5610);
and U9005 (N_9005,N_6907,N_7062);
xnor U9006 (N_9006,N_5601,N_5413);
and U9007 (N_9007,N_6260,N_7424);
or U9008 (N_9008,N_5307,N_7345);
nor U9009 (N_9009,N_7300,N_6121);
nand U9010 (N_9010,N_6957,N_5642);
nor U9011 (N_9011,N_5245,N_5128);
and U9012 (N_9012,N_5668,N_6948);
or U9013 (N_9013,N_6345,N_5392);
and U9014 (N_9014,N_7030,N_6966);
nor U9015 (N_9015,N_5581,N_6018);
or U9016 (N_9016,N_6450,N_6735);
xor U9017 (N_9017,N_5725,N_5791);
or U9018 (N_9018,N_5245,N_5804);
xnor U9019 (N_9019,N_5273,N_6779);
and U9020 (N_9020,N_7175,N_5059);
and U9021 (N_9021,N_6608,N_5087);
nor U9022 (N_9022,N_5030,N_6129);
or U9023 (N_9023,N_7018,N_6228);
nand U9024 (N_9024,N_5557,N_5355);
and U9025 (N_9025,N_6567,N_5576);
nor U9026 (N_9026,N_7339,N_6635);
and U9027 (N_9027,N_6750,N_7445);
or U9028 (N_9028,N_7362,N_6090);
nand U9029 (N_9029,N_6856,N_5165);
or U9030 (N_9030,N_5962,N_5456);
and U9031 (N_9031,N_7197,N_7272);
xnor U9032 (N_9032,N_5115,N_6301);
nor U9033 (N_9033,N_6606,N_6320);
or U9034 (N_9034,N_6843,N_5839);
and U9035 (N_9035,N_5712,N_7073);
nor U9036 (N_9036,N_6659,N_5796);
and U9037 (N_9037,N_6191,N_5620);
xor U9038 (N_9038,N_5988,N_6901);
nor U9039 (N_9039,N_6742,N_7477);
nand U9040 (N_9040,N_6354,N_7381);
nand U9041 (N_9041,N_5711,N_6517);
and U9042 (N_9042,N_6438,N_6394);
nand U9043 (N_9043,N_5907,N_7454);
nor U9044 (N_9044,N_6576,N_5778);
nor U9045 (N_9045,N_6984,N_7363);
nand U9046 (N_9046,N_6226,N_7411);
or U9047 (N_9047,N_5482,N_7116);
nand U9048 (N_9048,N_5340,N_5343);
and U9049 (N_9049,N_6109,N_6339);
nand U9050 (N_9050,N_6957,N_7035);
or U9051 (N_9051,N_6380,N_6912);
and U9052 (N_9052,N_6465,N_6346);
xor U9053 (N_9053,N_5875,N_7294);
nand U9054 (N_9054,N_7145,N_5432);
and U9055 (N_9055,N_6232,N_5761);
nor U9056 (N_9056,N_6648,N_5529);
or U9057 (N_9057,N_6960,N_7484);
or U9058 (N_9058,N_7303,N_7237);
nand U9059 (N_9059,N_6577,N_5167);
or U9060 (N_9060,N_6813,N_7190);
nand U9061 (N_9061,N_5722,N_5865);
or U9062 (N_9062,N_6689,N_6621);
and U9063 (N_9063,N_6860,N_5153);
nand U9064 (N_9064,N_6047,N_6845);
and U9065 (N_9065,N_7116,N_6156);
nor U9066 (N_9066,N_7037,N_6172);
and U9067 (N_9067,N_6978,N_6548);
nand U9068 (N_9068,N_7297,N_5865);
xor U9069 (N_9069,N_6019,N_6541);
and U9070 (N_9070,N_6542,N_6970);
nor U9071 (N_9071,N_6900,N_5343);
nor U9072 (N_9072,N_5292,N_6363);
nor U9073 (N_9073,N_5488,N_6305);
nor U9074 (N_9074,N_6569,N_7390);
or U9075 (N_9075,N_7037,N_5639);
or U9076 (N_9076,N_6861,N_5286);
or U9077 (N_9077,N_6308,N_7114);
nor U9078 (N_9078,N_7247,N_6336);
nor U9079 (N_9079,N_5332,N_6448);
nand U9080 (N_9080,N_6296,N_6288);
or U9081 (N_9081,N_6855,N_6621);
nor U9082 (N_9082,N_5062,N_5866);
nand U9083 (N_9083,N_5931,N_6163);
nor U9084 (N_9084,N_6984,N_6954);
nand U9085 (N_9085,N_5796,N_5976);
and U9086 (N_9086,N_6882,N_6679);
and U9087 (N_9087,N_6674,N_5000);
nand U9088 (N_9088,N_6376,N_5956);
nand U9089 (N_9089,N_5238,N_5407);
and U9090 (N_9090,N_7070,N_7269);
or U9091 (N_9091,N_6457,N_5572);
nand U9092 (N_9092,N_6747,N_7344);
xor U9093 (N_9093,N_6775,N_6601);
nor U9094 (N_9094,N_6562,N_6186);
nand U9095 (N_9095,N_5101,N_6523);
and U9096 (N_9096,N_5219,N_5036);
and U9097 (N_9097,N_6271,N_6436);
nor U9098 (N_9098,N_5586,N_5668);
nand U9099 (N_9099,N_6200,N_5676);
nor U9100 (N_9100,N_5210,N_6983);
or U9101 (N_9101,N_7375,N_6912);
and U9102 (N_9102,N_6029,N_5460);
and U9103 (N_9103,N_5609,N_7182);
nand U9104 (N_9104,N_5461,N_5469);
nor U9105 (N_9105,N_6285,N_5569);
nor U9106 (N_9106,N_6358,N_6993);
or U9107 (N_9107,N_6132,N_5913);
and U9108 (N_9108,N_5020,N_5866);
nor U9109 (N_9109,N_6676,N_7198);
nand U9110 (N_9110,N_5448,N_5977);
nor U9111 (N_9111,N_5941,N_7015);
nand U9112 (N_9112,N_6049,N_6884);
xnor U9113 (N_9113,N_7447,N_6351);
and U9114 (N_9114,N_6496,N_5826);
nand U9115 (N_9115,N_6210,N_5470);
or U9116 (N_9116,N_5611,N_6853);
nor U9117 (N_9117,N_6602,N_6807);
nand U9118 (N_9118,N_6716,N_5143);
or U9119 (N_9119,N_6997,N_6842);
and U9120 (N_9120,N_7147,N_5709);
or U9121 (N_9121,N_5650,N_6986);
nor U9122 (N_9122,N_5391,N_7239);
and U9123 (N_9123,N_5882,N_5351);
nand U9124 (N_9124,N_5571,N_7323);
nand U9125 (N_9125,N_5200,N_7130);
nor U9126 (N_9126,N_6652,N_6815);
nand U9127 (N_9127,N_5550,N_6110);
xor U9128 (N_9128,N_5843,N_7348);
nor U9129 (N_9129,N_6653,N_6881);
nand U9130 (N_9130,N_6850,N_5458);
and U9131 (N_9131,N_7367,N_6464);
nand U9132 (N_9132,N_7109,N_5080);
and U9133 (N_9133,N_6908,N_5867);
nand U9134 (N_9134,N_6693,N_5129);
or U9135 (N_9135,N_5694,N_6260);
nand U9136 (N_9136,N_6322,N_6161);
nor U9137 (N_9137,N_5054,N_6559);
xnor U9138 (N_9138,N_7001,N_7350);
nand U9139 (N_9139,N_6249,N_5132);
nand U9140 (N_9140,N_6931,N_7251);
or U9141 (N_9141,N_7111,N_5596);
or U9142 (N_9142,N_5976,N_7284);
nor U9143 (N_9143,N_6805,N_6658);
nand U9144 (N_9144,N_6403,N_6105);
xor U9145 (N_9145,N_6275,N_6167);
nand U9146 (N_9146,N_7130,N_6727);
nor U9147 (N_9147,N_7091,N_7156);
nor U9148 (N_9148,N_6703,N_5965);
xnor U9149 (N_9149,N_5671,N_7081);
xor U9150 (N_9150,N_5302,N_5645);
or U9151 (N_9151,N_5415,N_5078);
and U9152 (N_9152,N_7384,N_5107);
xor U9153 (N_9153,N_7036,N_6436);
nor U9154 (N_9154,N_6531,N_5701);
or U9155 (N_9155,N_5141,N_7416);
and U9156 (N_9156,N_5710,N_6056);
and U9157 (N_9157,N_5687,N_7277);
nand U9158 (N_9158,N_6668,N_6331);
and U9159 (N_9159,N_5628,N_7109);
or U9160 (N_9160,N_5021,N_5412);
nor U9161 (N_9161,N_7000,N_5182);
or U9162 (N_9162,N_7324,N_7458);
nor U9163 (N_9163,N_7051,N_5276);
nand U9164 (N_9164,N_5361,N_5441);
or U9165 (N_9165,N_5066,N_6560);
nor U9166 (N_9166,N_5378,N_5695);
or U9167 (N_9167,N_5679,N_6670);
nor U9168 (N_9168,N_7207,N_7428);
nor U9169 (N_9169,N_7023,N_7089);
nand U9170 (N_9170,N_7459,N_5266);
nor U9171 (N_9171,N_5276,N_5535);
nor U9172 (N_9172,N_6468,N_6512);
or U9173 (N_9173,N_6281,N_7132);
nor U9174 (N_9174,N_6911,N_5495);
nor U9175 (N_9175,N_7249,N_5095);
or U9176 (N_9176,N_5009,N_6471);
nand U9177 (N_9177,N_5131,N_6796);
xnor U9178 (N_9178,N_6686,N_5267);
and U9179 (N_9179,N_7418,N_6197);
xnor U9180 (N_9180,N_5079,N_7027);
nor U9181 (N_9181,N_6303,N_6685);
nor U9182 (N_9182,N_5192,N_6891);
nor U9183 (N_9183,N_6790,N_5506);
and U9184 (N_9184,N_5429,N_5682);
xor U9185 (N_9185,N_5171,N_6033);
nor U9186 (N_9186,N_7383,N_6928);
nand U9187 (N_9187,N_5047,N_5912);
nor U9188 (N_9188,N_6968,N_7393);
nor U9189 (N_9189,N_6481,N_6748);
nor U9190 (N_9190,N_6248,N_7350);
nor U9191 (N_9191,N_6089,N_5412);
xor U9192 (N_9192,N_6521,N_5090);
and U9193 (N_9193,N_5871,N_7373);
or U9194 (N_9194,N_7087,N_5455);
and U9195 (N_9195,N_6382,N_6211);
and U9196 (N_9196,N_7436,N_5001);
or U9197 (N_9197,N_6428,N_5419);
nand U9198 (N_9198,N_5699,N_6098);
nand U9199 (N_9199,N_5060,N_5374);
nor U9200 (N_9200,N_6051,N_7344);
and U9201 (N_9201,N_5065,N_6274);
xnor U9202 (N_9202,N_5679,N_5732);
or U9203 (N_9203,N_5085,N_6714);
nand U9204 (N_9204,N_7255,N_6354);
nor U9205 (N_9205,N_5492,N_5317);
nand U9206 (N_9206,N_6655,N_5646);
or U9207 (N_9207,N_7215,N_6983);
nand U9208 (N_9208,N_6112,N_6263);
nor U9209 (N_9209,N_6338,N_5515);
xor U9210 (N_9210,N_6230,N_5987);
nor U9211 (N_9211,N_6412,N_5315);
and U9212 (N_9212,N_5623,N_7492);
nand U9213 (N_9213,N_6852,N_6925);
nand U9214 (N_9214,N_6844,N_7178);
and U9215 (N_9215,N_5367,N_5671);
nand U9216 (N_9216,N_5075,N_5707);
or U9217 (N_9217,N_5221,N_6549);
nor U9218 (N_9218,N_5280,N_6564);
xnor U9219 (N_9219,N_5144,N_6061);
and U9220 (N_9220,N_6702,N_6733);
nand U9221 (N_9221,N_7193,N_7167);
nand U9222 (N_9222,N_6577,N_7097);
and U9223 (N_9223,N_5866,N_7446);
or U9224 (N_9224,N_7094,N_6000);
or U9225 (N_9225,N_6573,N_6761);
and U9226 (N_9226,N_5618,N_7394);
nor U9227 (N_9227,N_6348,N_6076);
nor U9228 (N_9228,N_5076,N_7436);
and U9229 (N_9229,N_7158,N_6504);
and U9230 (N_9230,N_7170,N_6576);
and U9231 (N_9231,N_5743,N_5762);
or U9232 (N_9232,N_5634,N_5575);
or U9233 (N_9233,N_5482,N_5456);
or U9234 (N_9234,N_6338,N_6874);
or U9235 (N_9235,N_7142,N_5332);
nor U9236 (N_9236,N_5653,N_7254);
nand U9237 (N_9237,N_5007,N_5269);
and U9238 (N_9238,N_7096,N_7331);
nand U9239 (N_9239,N_7302,N_6836);
nor U9240 (N_9240,N_5111,N_6417);
nand U9241 (N_9241,N_6722,N_6871);
or U9242 (N_9242,N_5302,N_5900);
and U9243 (N_9243,N_5404,N_6980);
and U9244 (N_9244,N_5084,N_5997);
or U9245 (N_9245,N_7449,N_6274);
xor U9246 (N_9246,N_7430,N_6382);
nor U9247 (N_9247,N_5773,N_5224);
xor U9248 (N_9248,N_6349,N_6737);
xor U9249 (N_9249,N_5893,N_6183);
and U9250 (N_9250,N_5535,N_6137);
nor U9251 (N_9251,N_5011,N_6598);
xor U9252 (N_9252,N_6498,N_5571);
nand U9253 (N_9253,N_7057,N_5684);
nand U9254 (N_9254,N_7467,N_6931);
nor U9255 (N_9255,N_6291,N_5393);
and U9256 (N_9256,N_6703,N_5481);
nor U9257 (N_9257,N_6120,N_5580);
or U9258 (N_9258,N_5434,N_6045);
nand U9259 (N_9259,N_5911,N_6396);
or U9260 (N_9260,N_5218,N_5711);
nand U9261 (N_9261,N_7291,N_7114);
or U9262 (N_9262,N_5534,N_5873);
nand U9263 (N_9263,N_5697,N_6936);
nor U9264 (N_9264,N_5211,N_6007);
or U9265 (N_9265,N_5154,N_5871);
and U9266 (N_9266,N_6879,N_6017);
and U9267 (N_9267,N_5540,N_7347);
xnor U9268 (N_9268,N_6896,N_6659);
xor U9269 (N_9269,N_5012,N_5946);
xor U9270 (N_9270,N_7162,N_5721);
or U9271 (N_9271,N_5554,N_5802);
nor U9272 (N_9272,N_7389,N_7151);
xor U9273 (N_9273,N_5620,N_7077);
nor U9274 (N_9274,N_6566,N_6535);
or U9275 (N_9275,N_6996,N_5583);
xnor U9276 (N_9276,N_7235,N_7150);
or U9277 (N_9277,N_5042,N_5263);
and U9278 (N_9278,N_6475,N_5015);
nor U9279 (N_9279,N_6349,N_5433);
nor U9280 (N_9280,N_6285,N_6033);
nor U9281 (N_9281,N_6848,N_5141);
nand U9282 (N_9282,N_5082,N_5695);
xor U9283 (N_9283,N_6554,N_6809);
nor U9284 (N_9284,N_5812,N_5792);
and U9285 (N_9285,N_5639,N_6853);
nor U9286 (N_9286,N_7144,N_7178);
nand U9287 (N_9287,N_6961,N_5148);
nand U9288 (N_9288,N_7112,N_6117);
or U9289 (N_9289,N_6020,N_6342);
xnor U9290 (N_9290,N_6340,N_6622);
xor U9291 (N_9291,N_6584,N_5627);
or U9292 (N_9292,N_5616,N_6707);
nor U9293 (N_9293,N_6328,N_6052);
nor U9294 (N_9294,N_6104,N_6052);
nand U9295 (N_9295,N_7438,N_6997);
nor U9296 (N_9296,N_6147,N_5695);
and U9297 (N_9297,N_7171,N_6529);
nor U9298 (N_9298,N_6769,N_6562);
nand U9299 (N_9299,N_7263,N_6449);
nor U9300 (N_9300,N_6046,N_6207);
and U9301 (N_9301,N_7033,N_5478);
nand U9302 (N_9302,N_6707,N_6705);
nand U9303 (N_9303,N_6525,N_7375);
nand U9304 (N_9304,N_5889,N_5259);
or U9305 (N_9305,N_5979,N_7044);
or U9306 (N_9306,N_6079,N_5315);
or U9307 (N_9307,N_7011,N_5174);
nor U9308 (N_9308,N_6170,N_5221);
and U9309 (N_9309,N_6577,N_5821);
nor U9310 (N_9310,N_5028,N_5372);
nand U9311 (N_9311,N_7134,N_6506);
nor U9312 (N_9312,N_6636,N_5119);
nor U9313 (N_9313,N_6535,N_5650);
or U9314 (N_9314,N_7496,N_6852);
or U9315 (N_9315,N_5144,N_5206);
or U9316 (N_9316,N_5792,N_6739);
nor U9317 (N_9317,N_5595,N_6749);
and U9318 (N_9318,N_5966,N_6864);
nor U9319 (N_9319,N_5735,N_6747);
nand U9320 (N_9320,N_5084,N_6110);
nand U9321 (N_9321,N_6246,N_7331);
nand U9322 (N_9322,N_5715,N_5717);
nand U9323 (N_9323,N_5766,N_6660);
nor U9324 (N_9324,N_6474,N_5994);
nand U9325 (N_9325,N_6098,N_5417);
and U9326 (N_9326,N_6458,N_7050);
nand U9327 (N_9327,N_6194,N_6794);
or U9328 (N_9328,N_5955,N_6492);
and U9329 (N_9329,N_6992,N_7084);
and U9330 (N_9330,N_5162,N_6574);
or U9331 (N_9331,N_5133,N_6346);
and U9332 (N_9332,N_7190,N_7182);
or U9333 (N_9333,N_6613,N_6963);
nor U9334 (N_9334,N_5091,N_5385);
nand U9335 (N_9335,N_6252,N_5904);
and U9336 (N_9336,N_5552,N_6979);
nor U9337 (N_9337,N_5568,N_6711);
and U9338 (N_9338,N_6123,N_7098);
nor U9339 (N_9339,N_5795,N_5937);
xor U9340 (N_9340,N_6417,N_6689);
or U9341 (N_9341,N_5738,N_6617);
nand U9342 (N_9342,N_5132,N_7061);
and U9343 (N_9343,N_5259,N_5536);
nor U9344 (N_9344,N_5240,N_5092);
nor U9345 (N_9345,N_6424,N_6017);
xnor U9346 (N_9346,N_7414,N_6529);
nor U9347 (N_9347,N_5789,N_6592);
nand U9348 (N_9348,N_5820,N_6273);
nor U9349 (N_9349,N_5706,N_7076);
nor U9350 (N_9350,N_7211,N_6836);
nand U9351 (N_9351,N_5030,N_6825);
nor U9352 (N_9352,N_5624,N_7496);
and U9353 (N_9353,N_5646,N_5260);
nor U9354 (N_9354,N_6836,N_7070);
xor U9355 (N_9355,N_6808,N_7427);
nand U9356 (N_9356,N_6032,N_5290);
xnor U9357 (N_9357,N_7491,N_6924);
nand U9358 (N_9358,N_5572,N_7051);
and U9359 (N_9359,N_5577,N_7213);
nand U9360 (N_9360,N_7260,N_6543);
or U9361 (N_9361,N_6007,N_6051);
nor U9362 (N_9362,N_5524,N_6806);
nor U9363 (N_9363,N_7137,N_7030);
nand U9364 (N_9364,N_5060,N_6335);
and U9365 (N_9365,N_5957,N_6466);
nand U9366 (N_9366,N_6414,N_5275);
nand U9367 (N_9367,N_7319,N_6016);
or U9368 (N_9368,N_5059,N_6486);
and U9369 (N_9369,N_6456,N_6271);
nor U9370 (N_9370,N_6284,N_6718);
and U9371 (N_9371,N_7276,N_6687);
nand U9372 (N_9372,N_6474,N_6937);
nor U9373 (N_9373,N_7009,N_6931);
nand U9374 (N_9374,N_7064,N_6805);
nor U9375 (N_9375,N_5856,N_6626);
or U9376 (N_9376,N_7339,N_5379);
nor U9377 (N_9377,N_7185,N_7352);
nor U9378 (N_9378,N_5753,N_7040);
nand U9379 (N_9379,N_6794,N_5729);
nor U9380 (N_9380,N_7221,N_5731);
nor U9381 (N_9381,N_5683,N_7451);
nand U9382 (N_9382,N_5633,N_5551);
and U9383 (N_9383,N_7234,N_7148);
or U9384 (N_9384,N_6767,N_6781);
nand U9385 (N_9385,N_6007,N_6510);
or U9386 (N_9386,N_5461,N_5259);
and U9387 (N_9387,N_5363,N_5566);
and U9388 (N_9388,N_5985,N_5153);
and U9389 (N_9389,N_6817,N_5230);
nand U9390 (N_9390,N_5100,N_5336);
and U9391 (N_9391,N_5259,N_5768);
xor U9392 (N_9392,N_6872,N_5504);
xnor U9393 (N_9393,N_6962,N_6394);
nor U9394 (N_9394,N_5132,N_5198);
nor U9395 (N_9395,N_5686,N_6312);
and U9396 (N_9396,N_7264,N_7373);
nand U9397 (N_9397,N_6304,N_5757);
and U9398 (N_9398,N_6089,N_6446);
xor U9399 (N_9399,N_6973,N_7272);
nand U9400 (N_9400,N_6058,N_5367);
nand U9401 (N_9401,N_6854,N_6253);
nor U9402 (N_9402,N_6691,N_7128);
nand U9403 (N_9403,N_7444,N_7180);
nand U9404 (N_9404,N_7346,N_5660);
nand U9405 (N_9405,N_5053,N_5775);
and U9406 (N_9406,N_6953,N_5464);
or U9407 (N_9407,N_5406,N_6659);
and U9408 (N_9408,N_6576,N_5826);
nand U9409 (N_9409,N_6940,N_5904);
and U9410 (N_9410,N_5345,N_6196);
and U9411 (N_9411,N_6974,N_5445);
nor U9412 (N_9412,N_6817,N_6560);
nand U9413 (N_9413,N_7117,N_7040);
nor U9414 (N_9414,N_5568,N_6010);
or U9415 (N_9415,N_6218,N_7378);
nor U9416 (N_9416,N_6305,N_5353);
and U9417 (N_9417,N_5642,N_5609);
and U9418 (N_9418,N_5489,N_7148);
nor U9419 (N_9419,N_5512,N_5120);
and U9420 (N_9420,N_5789,N_5955);
nor U9421 (N_9421,N_5429,N_7381);
nor U9422 (N_9422,N_5797,N_7435);
nor U9423 (N_9423,N_6040,N_7442);
and U9424 (N_9424,N_6140,N_5283);
nor U9425 (N_9425,N_6667,N_6945);
or U9426 (N_9426,N_5654,N_6247);
nand U9427 (N_9427,N_6171,N_6398);
xnor U9428 (N_9428,N_6917,N_5954);
and U9429 (N_9429,N_6866,N_5862);
or U9430 (N_9430,N_5837,N_7323);
nor U9431 (N_9431,N_7026,N_6501);
nand U9432 (N_9432,N_6985,N_5274);
or U9433 (N_9433,N_6851,N_6112);
nand U9434 (N_9434,N_5038,N_7331);
or U9435 (N_9435,N_7229,N_6586);
and U9436 (N_9436,N_6868,N_5534);
nand U9437 (N_9437,N_7465,N_7362);
nand U9438 (N_9438,N_5894,N_5273);
and U9439 (N_9439,N_6278,N_5142);
nand U9440 (N_9440,N_6436,N_6903);
and U9441 (N_9441,N_5272,N_6358);
xnor U9442 (N_9442,N_5132,N_5071);
or U9443 (N_9443,N_6168,N_7016);
and U9444 (N_9444,N_5712,N_6212);
xor U9445 (N_9445,N_5433,N_5156);
and U9446 (N_9446,N_5666,N_5325);
nand U9447 (N_9447,N_7414,N_7194);
nor U9448 (N_9448,N_6048,N_7118);
nand U9449 (N_9449,N_5580,N_5729);
nor U9450 (N_9450,N_7103,N_6368);
nand U9451 (N_9451,N_5728,N_6340);
nand U9452 (N_9452,N_5339,N_7264);
or U9453 (N_9453,N_5653,N_5242);
or U9454 (N_9454,N_5046,N_6089);
nand U9455 (N_9455,N_6227,N_6146);
nor U9456 (N_9456,N_6702,N_5349);
nor U9457 (N_9457,N_6643,N_5032);
and U9458 (N_9458,N_5235,N_5257);
nand U9459 (N_9459,N_7255,N_6007);
nor U9460 (N_9460,N_7400,N_6873);
nor U9461 (N_9461,N_5460,N_5014);
nand U9462 (N_9462,N_6352,N_5531);
nor U9463 (N_9463,N_6404,N_6473);
or U9464 (N_9464,N_7427,N_7388);
and U9465 (N_9465,N_5887,N_7270);
nor U9466 (N_9466,N_5481,N_7493);
or U9467 (N_9467,N_5874,N_6095);
or U9468 (N_9468,N_5612,N_5346);
nand U9469 (N_9469,N_6671,N_6517);
or U9470 (N_9470,N_7316,N_5947);
or U9471 (N_9471,N_6748,N_5610);
or U9472 (N_9472,N_7214,N_5716);
nor U9473 (N_9473,N_7025,N_6038);
or U9474 (N_9474,N_6326,N_5440);
nor U9475 (N_9475,N_7327,N_5542);
nor U9476 (N_9476,N_5363,N_6538);
nand U9477 (N_9477,N_6163,N_5035);
nor U9478 (N_9478,N_5760,N_5124);
nand U9479 (N_9479,N_6641,N_6465);
nor U9480 (N_9480,N_6532,N_6369);
and U9481 (N_9481,N_6175,N_5573);
nor U9482 (N_9482,N_6068,N_7394);
or U9483 (N_9483,N_6632,N_7434);
xnor U9484 (N_9484,N_5347,N_6660);
nand U9485 (N_9485,N_5625,N_6504);
nand U9486 (N_9486,N_6889,N_7222);
or U9487 (N_9487,N_7042,N_7228);
or U9488 (N_9488,N_5132,N_5619);
nor U9489 (N_9489,N_7350,N_5519);
or U9490 (N_9490,N_6686,N_6072);
nand U9491 (N_9491,N_5325,N_5059);
nand U9492 (N_9492,N_5260,N_6539);
nand U9493 (N_9493,N_5930,N_6431);
or U9494 (N_9494,N_5850,N_7250);
and U9495 (N_9495,N_6059,N_6559);
nand U9496 (N_9496,N_6953,N_5038);
nor U9497 (N_9497,N_7474,N_7266);
nor U9498 (N_9498,N_5667,N_6519);
nand U9499 (N_9499,N_5149,N_7005);
and U9500 (N_9500,N_7135,N_5781);
nor U9501 (N_9501,N_6386,N_7483);
nand U9502 (N_9502,N_5711,N_5231);
nor U9503 (N_9503,N_6169,N_6394);
or U9504 (N_9504,N_5646,N_5827);
xor U9505 (N_9505,N_5917,N_6011);
or U9506 (N_9506,N_5871,N_5336);
or U9507 (N_9507,N_6415,N_6962);
nor U9508 (N_9508,N_6949,N_5179);
nand U9509 (N_9509,N_5908,N_5772);
nor U9510 (N_9510,N_5823,N_6492);
or U9511 (N_9511,N_5494,N_7261);
and U9512 (N_9512,N_5936,N_6090);
or U9513 (N_9513,N_6163,N_7275);
and U9514 (N_9514,N_6965,N_6526);
and U9515 (N_9515,N_6933,N_5448);
and U9516 (N_9516,N_6526,N_7468);
nor U9517 (N_9517,N_5817,N_5464);
nor U9518 (N_9518,N_6062,N_5975);
nand U9519 (N_9519,N_5286,N_5143);
or U9520 (N_9520,N_7083,N_6058);
nor U9521 (N_9521,N_5636,N_7051);
or U9522 (N_9522,N_7417,N_6694);
nor U9523 (N_9523,N_7450,N_5537);
nand U9524 (N_9524,N_5239,N_5683);
and U9525 (N_9525,N_5975,N_7385);
or U9526 (N_9526,N_7318,N_6766);
nand U9527 (N_9527,N_6954,N_6561);
nand U9528 (N_9528,N_5671,N_5831);
nor U9529 (N_9529,N_5617,N_5928);
xnor U9530 (N_9530,N_7374,N_6414);
or U9531 (N_9531,N_5386,N_7091);
and U9532 (N_9532,N_6647,N_6494);
nand U9533 (N_9533,N_5396,N_5101);
nand U9534 (N_9534,N_6260,N_5959);
xor U9535 (N_9535,N_5825,N_7084);
or U9536 (N_9536,N_5794,N_5329);
or U9537 (N_9537,N_6600,N_5539);
or U9538 (N_9538,N_6949,N_6486);
or U9539 (N_9539,N_7436,N_7074);
nor U9540 (N_9540,N_6990,N_6255);
nand U9541 (N_9541,N_7214,N_5814);
or U9542 (N_9542,N_6206,N_5879);
and U9543 (N_9543,N_6583,N_5819);
nor U9544 (N_9544,N_5463,N_6169);
and U9545 (N_9545,N_7049,N_5645);
nand U9546 (N_9546,N_6000,N_5438);
nand U9547 (N_9547,N_5634,N_6658);
nor U9548 (N_9548,N_5886,N_7385);
or U9549 (N_9549,N_5817,N_5401);
and U9550 (N_9550,N_5599,N_6529);
or U9551 (N_9551,N_6801,N_7271);
and U9552 (N_9552,N_7051,N_6854);
nor U9553 (N_9553,N_6618,N_5231);
nor U9554 (N_9554,N_5106,N_5696);
nor U9555 (N_9555,N_7458,N_7344);
and U9556 (N_9556,N_5953,N_5142);
and U9557 (N_9557,N_5457,N_6503);
nor U9558 (N_9558,N_5522,N_7389);
and U9559 (N_9559,N_5864,N_6816);
and U9560 (N_9560,N_6912,N_6228);
or U9561 (N_9561,N_5013,N_5442);
nand U9562 (N_9562,N_6418,N_6648);
nor U9563 (N_9563,N_5466,N_5419);
and U9564 (N_9564,N_5542,N_7028);
or U9565 (N_9565,N_5938,N_7139);
nand U9566 (N_9566,N_5953,N_5848);
nor U9567 (N_9567,N_6615,N_5201);
and U9568 (N_9568,N_5269,N_5939);
nor U9569 (N_9569,N_7371,N_6986);
nor U9570 (N_9570,N_6426,N_7007);
xnor U9571 (N_9571,N_7436,N_7265);
or U9572 (N_9572,N_6239,N_5639);
nand U9573 (N_9573,N_5219,N_6111);
nand U9574 (N_9574,N_6307,N_5741);
nand U9575 (N_9575,N_5019,N_6929);
nor U9576 (N_9576,N_6851,N_5426);
or U9577 (N_9577,N_7312,N_6343);
nor U9578 (N_9578,N_5295,N_5311);
and U9579 (N_9579,N_5280,N_6631);
xnor U9580 (N_9580,N_5599,N_6157);
nor U9581 (N_9581,N_5116,N_5969);
nor U9582 (N_9582,N_7030,N_7378);
and U9583 (N_9583,N_5473,N_5433);
nand U9584 (N_9584,N_5810,N_6393);
nand U9585 (N_9585,N_7365,N_5115);
nand U9586 (N_9586,N_5402,N_5782);
or U9587 (N_9587,N_6271,N_5971);
nor U9588 (N_9588,N_7148,N_6255);
nor U9589 (N_9589,N_5346,N_6762);
or U9590 (N_9590,N_5543,N_5392);
nand U9591 (N_9591,N_5770,N_6006);
nand U9592 (N_9592,N_7204,N_6325);
or U9593 (N_9593,N_6604,N_5570);
nand U9594 (N_9594,N_6673,N_5485);
xnor U9595 (N_9595,N_5021,N_5531);
nand U9596 (N_9596,N_5171,N_5941);
and U9597 (N_9597,N_5151,N_5557);
nand U9598 (N_9598,N_5487,N_6359);
or U9599 (N_9599,N_5942,N_7439);
and U9600 (N_9600,N_6281,N_5741);
and U9601 (N_9601,N_5437,N_6665);
nor U9602 (N_9602,N_5488,N_6996);
and U9603 (N_9603,N_5462,N_7003);
and U9604 (N_9604,N_5441,N_6164);
and U9605 (N_9605,N_5870,N_6010);
nor U9606 (N_9606,N_5371,N_6099);
or U9607 (N_9607,N_6932,N_6535);
or U9608 (N_9608,N_6204,N_5175);
nor U9609 (N_9609,N_6611,N_5047);
or U9610 (N_9610,N_7170,N_6961);
nand U9611 (N_9611,N_6023,N_6314);
and U9612 (N_9612,N_5886,N_6886);
or U9613 (N_9613,N_7489,N_7139);
nor U9614 (N_9614,N_6889,N_7002);
nand U9615 (N_9615,N_5288,N_6452);
xor U9616 (N_9616,N_5446,N_6123);
nor U9617 (N_9617,N_5631,N_6158);
xnor U9618 (N_9618,N_6149,N_6749);
and U9619 (N_9619,N_6242,N_7185);
and U9620 (N_9620,N_5294,N_7069);
and U9621 (N_9621,N_5303,N_5287);
and U9622 (N_9622,N_5515,N_6129);
and U9623 (N_9623,N_5905,N_6886);
nand U9624 (N_9624,N_6509,N_7407);
nor U9625 (N_9625,N_7187,N_6090);
or U9626 (N_9626,N_5977,N_5778);
xor U9627 (N_9627,N_7443,N_7075);
and U9628 (N_9628,N_5152,N_7249);
or U9629 (N_9629,N_5176,N_6258);
nand U9630 (N_9630,N_6542,N_7362);
and U9631 (N_9631,N_6256,N_5222);
nor U9632 (N_9632,N_6891,N_5416);
nand U9633 (N_9633,N_5786,N_7208);
and U9634 (N_9634,N_6556,N_5476);
nand U9635 (N_9635,N_5434,N_5627);
and U9636 (N_9636,N_5699,N_5363);
or U9637 (N_9637,N_6013,N_5090);
and U9638 (N_9638,N_7051,N_6476);
and U9639 (N_9639,N_7333,N_6341);
nor U9640 (N_9640,N_5465,N_6975);
nand U9641 (N_9641,N_6318,N_6721);
nor U9642 (N_9642,N_6105,N_6193);
nor U9643 (N_9643,N_6045,N_5437);
and U9644 (N_9644,N_7372,N_7340);
and U9645 (N_9645,N_6559,N_6177);
and U9646 (N_9646,N_6128,N_6200);
and U9647 (N_9647,N_5961,N_5447);
nor U9648 (N_9648,N_6654,N_6439);
nand U9649 (N_9649,N_5322,N_6423);
xnor U9650 (N_9650,N_5117,N_5948);
or U9651 (N_9651,N_5242,N_5226);
and U9652 (N_9652,N_6473,N_6031);
nor U9653 (N_9653,N_6578,N_5479);
nand U9654 (N_9654,N_6697,N_7303);
or U9655 (N_9655,N_7000,N_6332);
xor U9656 (N_9656,N_5067,N_5564);
xnor U9657 (N_9657,N_5166,N_6476);
nor U9658 (N_9658,N_5619,N_6787);
and U9659 (N_9659,N_7084,N_6960);
nor U9660 (N_9660,N_7163,N_6967);
nor U9661 (N_9661,N_5173,N_6083);
and U9662 (N_9662,N_6743,N_5666);
nand U9663 (N_9663,N_7416,N_7069);
xnor U9664 (N_9664,N_6762,N_6360);
and U9665 (N_9665,N_6972,N_5907);
and U9666 (N_9666,N_5339,N_7098);
xor U9667 (N_9667,N_6994,N_6658);
nor U9668 (N_9668,N_5549,N_5233);
nor U9669 (N_9669,N_6841,N_6500);
and U9670 (N_9670,N_5012,N_6617);
or U9671 (N_9671,N_7460,N_6850);
nor U9672 (N_9672,N_7099,N_5780);
nand U9673 (N_9673,N_6890,N_6989);
nor U9674 (N_9674,N_6716,N_7057);
nand U9675 (N_9675,N_5873,N_7057);
nand U9676 (N_9676,N_7414,N_5277);
or U9677 (N_9677,N_5336,N_7251);
or U9678 (N_9678,N_6114,N_6302);
xor U9679 (N_9679,N_5949,N_5944);
and U9680 (N_9680,N_5633,N_7290);
or U9681 (N_9681,N_6692,N_7268);
and U9682 (N_9682,N_5502,N_6936);
nand U9683 (N_9683,N_6548,N_5310);
and U9684 (N_9684,N_7222,N_7442);
or U9685 (N_9685,N_5746,N_5677);
nand U9686 (N_9686,N_5578,N_6807);
or U9687 (N_9687,N_6384,N_6000);
xnor U9688 (N_9688,N_7445,N_6721);
and U9689 (N_9689,N_6653,N_5035);
or U9690 (N_9690,N_5280,N_5085);
nor U9691 (N_9691,N_6857,N_6389);
nand U9692 (N_9692,N_5744,N_6743);
and U9693 (N_9693,N_6095,N_6397);
nand U9694 (N_9694,N_6445,N_7107);
xnor U9695 (N_9695,N_7454,N_6410);
or U9696 (N_9696,N_5388,N_6477);
and U9697 (N_9697,N_5735,N_5985);
xnor U9698 (N_9698,N_7420,N_7355);
or U9699 (N_9699,N_5861,N_6120);
and U9700 (N_9700,N_6126,N_5484);
nand U9701 (N_9701,N_5962,N_5591);
and U9702 (N_9702,N_5562,N_5423);
or U9703 (N_9703,N_6078,N_6176);
nand U9704 (N_9704,N_6107,N_5753);
and U9705 (N_9705,N_6705,N_6983);
or U9706 (N_9706,N_6201,N_6702);
nor U9707 (N_9707,N_6216,N_7277);
nor U9708 (N_9708,N_6618,N_7030);
nand U9709 (N_9709,N_5703,N_5600);
nor U9710 (N_9710,N_5922,N_6679);
and U9711 (N_9711,N_5670,N_6157);
nor U9712 (N_9712,N_5668,N_6282);
and U9713 (N_9713,N_5558,N_6969);
xor U9714 (N_9714,N_6201,N_5647);
or U9715 (N_9715,N_7422,N_7216);
and U9716 (N_9716,N_5070,N_6825);
nand U9717 (N_9717,N_6206,N_6317);
nand U9718 (N_9718,N_6548,N_6707);
or U9719 (N_9719,N_5778,N_6176);
nor U9720 (N_9720,N_5111,N_6887);
and U9721 (N_9721,N_5259,N_6187);
or U9722 (N_9722,N_7296,N_5552);
and U9723 (N_9723,N_6343,N_7148);
or U9724 (N_9724,N_5009,N_7082);
and U9725 (N_9725,N_5292,N_6438);
nor U9726 (N_9726,N_5226,N_5357);
or U9727 (N_9727,N_5656,N_6636);
or U9728 (N_9728,N_7059,N_5264);
or U9729 (N_9729,N_5904,N_6905);
and U9730 (N_9730,N_7284,N_5995);
or U9731 (N_9731,N_5320,N_5976);
or U9732 (N_9732,N_6274,N_5300);
nand U9733 (N_9733,N_6445,N_6636);
nor U9734 (N_9734,N_7117,N_7015);
xnor U9735 (N_9735,N_6859,N_6025);
nand U9736 (N_9736,N_7235,N_6678);
and U9737 (N_9737,N_5783,N_5780);
and U9738 (N_9738,N_6704,N_7035);
nor U9739 (N_9739,N_6824,N_5742);
nor U9740 (N_9740,N_6641,N_5139);
or U9741 (N_9741,N_5612,N_7485);
or U9742 (N_9742,N_7082,N_6153);
and U9743 (N_9743,N_7298,N_7268);
xor U9744 (N_9744,N_6270,N_5106);
nand U9745 (N_9745,N_6081,N_5495);
xor U9746 (N_9746,N_5446,N_5957);
or U9747 (N_9747,N_6667,N_6044);
or U9748 (N_9748,N_7279,N_6515);
nand U9749 (N_9749,N_5250,N_5185);
xor U9750 (N_9750,N_6213,N_6521);
nor U9751 (N_9751,N_5048,N_7197);
or U9752 (N_9752,N_6534,N_5149);
nand U9753 (N_9753,N_7233,N_7335);
nand U9754 (N_9754,N_6189,N_7385);
or U9755 (N_9755,N_7433,N_7497);
and U9756 (N_9756,N_6489,N_6736);
xnor U9757 (N_9757,N_5148,N_7323);
nor U9758 (N_9758,N_6848,N_7046);
or U9759 (N_9759,N_7370,N_5008);
and U9760 (N_9760,N_6066,N_6617);
and U9761 (N_9761,N_7377,N_6092);
or U9762 (N_9762,N_7004,N_6967);
nand U9763 (N_9763,N_6595,N_7310);
nor U9764 (N_9764,N_5496,N_5063);
xor U9765 (N_9765,N_6690,N_5818);
and U9766 (N_9766,N_6178,N_6761);
nand U9767 (N_9767,N_5194,N_5994);
xor U9768 (N_9768,N_5809,N_5860);
or U9769 (N_9769,N_5414,N_7249);
nor U9770 (N_9770,N_5164,N_5552);
nand U9771 (N_9771,N_5043,N_5436);
and U9772 (N_9772,N_5535,N_6639);
xor U9773 (N_9773,N_7159,N_7453);
nor U9774 (N_9774,N_5800,N_7412);
nor U9775 (N_9775,N_6522,N_6345);
and U9776 (N_9776,N_7030,N_6146);
nand U9777 (N_9777,N_7120,N_5518);
or U9778 (N_9778,N_5958,N_5718);
xor U9779 (N_9779,N_7408,N_7019);
or U9780 (N_9780,N_7295,N_5484);
or U9781 (N_9781,N_5753,N_6437);
or U9782 (N_9782,N_6325,N_6107);
nand U9783 (N_9783,N_6130,N_7124);
or U9784 (N_9784,N_7394,N_5742);
and U9785 (N_9785,N_5124,N_6237);
and U9786 (N_9786,N_6484,N_7464);
nand U9787 (N_9787,N_6161,N_5350);
and U9788 (N_9788,N_5605,N_5329);
nor U9789 (N_9789,N_6125,N_6424);
nor U9790 (N_9790,N_7114,N_6709);
nand U9791 (N_9791,N_5315,N_7136);
nor U9792 (N_9792,N_6106,N_7266);
nor U9793 (N_9793,N_6851,N_5308);
and U9794 (N_9794,N_7188,N_7184);
nand U9795 (N_9795,N_6976,N_6519);
nor U9796 (N_9796,N_5073,N_5038);
and U9797 (N_9797,N_7277,N_7189);
or U9798 (N_9798,N_7052,N_6824);
xor U9799 (N_9799,N_7167,N_7451);
nor U9800 (N_9800,N_7107,N_5199);
or U9801 (N_9801,N_6556,N_5216);
and U9802 (N_9802,N_5074,N_6619);
and U9803 (N_9803,N_5352,N_5546);
nor U9804 (N_9804,N_5411,N_5749);
nand U9805 (N_9805,N_5958,N_6692);
nand U9806 (N_9806,N_6732,N_7441);
and U9807 (N_9807,N_6647,N_5512);
and U9808 (N_9808,N_5783,N_5074);
nand U9809 (N_9809,N_5145,N_6415);
nand U9810 (N_9810,N_6461,N_6102);
and U9811 (N_9811,N_5163,N_5251);
nor U9812 (N_9812,N_6085,N_5931);
and U9813 (N_9813,N_7209,N_5888);
nand U9814 (N_9814,N_6140,N_6954);
nor U9815 (N_9815,N_5772,N_7043);
xor U9816 (N_9816,N_5874,N_7099);
or U9817 (N_9817,N_5941,N_5743);
xnor U9818 (N_9818,N_5275,N_6690);
nand U9819 (N_9819,N_7159,N_6809);
nor U9820 (N_9820,N_7407,N_7419);
or U9821 (N_9821,N_5189,N_5666);
nand U9822 (N_9822,N_7357,N_6762);
and U9823 (N_9823,N_5035,N_7415);
xor U9824 (N_9824,N_6264,N_5163);
nor U9825 (N_9825,N_7498,N_5257);
and U9826 (N_9826,N_5287,N_5333);
nand U9827 (N_9827,N_5333,N_6976);
nand U9828 (N_9828,N_5915,N_7075);
nand U9829 (N_9829,N_6856,N_5254);
nor U9830 (N_9830,N_6168,N_5829);
xnor U9831 (N_9831,N_5116,N_7195);
or U9832 (N_9832,N_5800,N_7118);
and U9833 (N_9833,N_6957,N_6403);
and U9834 (N_9834,N_6029,N_7085);
nor U9835 (N_9835,N_6736,N_7085);
xnor U9836 (N_9836,N_6099,N_5681);
or U9837 (N_9837,N_6984,N_6804);
or U9838 (N_9838,N_6486,N_6900);
or U9839 (N_9839,N_5166,N_6103);
nand U9840 (N_9840,N_7152,N_7464);
or U9841 (N_9841,N_5416,N_6680);
or U9842 (N_9842,N_6784,N_5172);
and U9843 (N_9843,N_6207,N_6379);
or U9844 (N_9844,N_5465,N_6337);
xnor U9845 (N_9845,N_6590,N_5782);
nor U9846 (N_9846,N_5963,N_6512);
or U9847 (N_9847,N_5015,N_7097);
nand U9848 (N_9848,N_6709,N_5708);
nand U9849 (N_9849,N_7373,N_5602);
xnor U9850 (N_9850,N_5102,N_6300);
nand U9851 (N_9851,N_6536,N_5094);
or U9852 (N_9852,N_7174,N_7463);
or U9853 (N_9853,N_7220,N_6494);
nor U9854 (N_9854,N_5818,N_5179);
nand U9855 (N_9855,N_5909,N_5675);
nor U9856 (N_9856,N_5772,N_5419);
nor U9857 (N_9857,N_6761,N_5857);
and U9858 (N_9858,N_6835,N_7310);
or U9859 (N_9859,N_6563,N_5759);
nand U9860 (N_9860,N_5674,N_7295);
or U9861 (N_9861,N_5533,N_7077);
or U9862 (N_9862,N_5788,N_5287);
nor U9863 (N_9863,N_5770,N_5913);
nand U9864 (N_9864,N_5687,N_5129);
nand U9865 (N_9865,N_6784,N_6310);
nand U9866 (N_9866,N_5144,N_6105);
or U9867 (N_9867,N_7048,N_6269);
nor U9868 (N_9868,N_5091,N_5458);
nor U9869 (N_9869,N_5380,N_6321);
nand U9870 (N_9870,N_7208,N_5818);
nand U9871 (N_9871,N_6888,N_5147);
or U9872 (N_9872,N_5873,N_7237);
and U9873 (N_9873,N_7294,N_6607);
and U9874 (N_9874,N_5888,N_6779);
nor U9875 (N_9875,N_5335,N_5485);
and U9876 (N_9876,N_5577,N_6398);
nand U9877 (N_9877,N_5509,N_5152);
or U9878 (N_9878,N_6191,N_6427);
or U9879 (N_9879,N_7384,N_6269);
nor U9880 (N_9880,N_7259,N_6545);
or U9881 (N_9881,N_6850,N_6695);
xnor U9882 (N_9882,N_6687,N_6032);
nor U9883 (N_9883,N_6151,N_5354);
nand U9884 (N_9884,N_5641,N_5237);
nand U9885 (N_9885,N_5141,N_6709);
or U9886 (N_9886,N_6790,N_5758);
and U9887 (N_9887,N_5511,N_7346);
nor U9888 (N_9888,N_7438,N_5990);
and U9889 (N_9889,N_5459,N_6777);
nor U9890 (N_9890,N_7472,N_7042);
xor U9891 (N_9891,N_6541,N_5506);
and U9892 (N_9892,N_6053,N_6643);
xnor U9893 (N_9893,N_6181,N_7288);
nand U9894 (N_9894,N_7356,N_5401);
nand U9895 (N_9895,N_6892,N_7289);
nand U9896 (N_9896,N_6807,N_7349);
nand U9897 (N_9897,N_6428,N_7277);
nor U9898 (N_9898,N_7246,N_6237);
or U9899 (N_9899,N_5582,N_6664);
nand U9900 (N_9900,N_7255,N_6437);
or U9901 (N_9901,N_7090,N_5642);
nor U9902 (N_9902,N_6864,N_6709);
nor U9903 (N_9903,N_6828,N_5411);
and U9904 (N_9904,N_6292,N_6623);
nand U9905 (N_9905,N_5692,N_6566);
nor U9906 (N_9906,N_6907,N_6801);
nand U9907 (N_9907,N_7229,N_7456);
nor U9908 (N_9908,N_5481,N_6838);
nor U9909 (N_9909,N_6963,N_5275);
nand U9910 (N_9910,N_6757,N_6925);
nor U9911 (N_9911,N_6710,N_5069);
or U9912 (N_9912,N_5359,N_5416);
xnor U9913 (N_9913,N_6659,N_6377);
and U9914 (N_9914,N_6519,N_6765);
nand U9915 (N_9915,N_7400,N_6025);
nand U9916 (N_9916,N_5715,N_5955);
nand U9917 (N_9917,N_6492,N_5198);
and U9918 (N_9918,N_6282,N_5261);
nor U9919 (N_9919,N_5873,N_5680);
nand U9920 (N_9920,N_6601,N_7341);
nand U9921 (N_9921,N_5607,N_6377);
and U9922 (N_9922,N_6746,N_5389);
or U9923 (N_9923,N_6880,N_6646);
and U9924 (N_9924,N_7060,N_5441);
or U9925 (N_9925,N_6286,N_5211);
nor U9926 (N_9926,N_6476,N_6624);
xnor U9927 (N_9927,N_6286,N_6205);
and U9928 (N_9928,N_5745,N_6737);
nor U9929 (N_9929,N_5256,N_6055);
xor U9930 (N_9930,N_6276,N_6895);
nand U9931 (N_9931,N_5751,N_6418);
nand U9932 (N_9932,N_6205,N_5084);
nand U9933 (N_9933,N_5397,N_6035);
and U9934 (N_9934,N_7384,N_6204);
xnor U9935 (N_9935,N_6312,N_5312);
nand U9936 (N_9936,N_6556,N_5809);
xor U9937 (N_9937,N_6756,N_5122);
or U9938 (N_9938,N_6001,N_5697);
nor U9939 (N_9939,N_6371,N_5248);
nand U9940 (N_9940,N_7156,N_6699);
xor U9941 (N_9941,N_6764,N_6901);
nor U9942 (N_9942,N_6308,N_6141);
or U9943 (N_9943,N_6047,N_5194);
nor U9944 (N_9944,N_5142,N_6558);
nand U9945 (N_9945,N_6800,N_5341);
or U9946 (N_9946,N_6128,N_5632);
and U9947 (N_9947,N_6199,N_5832);
and U9948 (N_9948,N_6955,N_6724);
nand U9949 (N_9949,N_5644,N_7290);
xor U9950 (N_9950,N_6333,N_6605);
or U9951 (N_9951,N_6999,N_6101);
nand U9952 (N_9952,N_5311,N_6970);
xnor U9953 (N_9953,N_6647,N_5666);
xor U9954 (N_9954,N_5483,N_6233);
nor U9955 (N_9955,N_6719,N_6530);
xor U9956 (N_9956,N_5223,N_5638);
nand U9957 (N_9957,N_6029,N_6563);
nor U9958 (N_9958,N_6438,N_7167);
or U9959 (N_9959,N_5949,N_5063);
nor U9960 (N_9960,N_7372,N_5715);
nand U9961 (N_9961,N_5804,N_7473);
nand U9962 (N_9962,N_6198,N_5488);
nand U9963 (N_9963,N_6497,N_7247);
nand U9964 (N_9964,N_6484,N_5859);
or U9965 (N_9965,N_7499,N_6588);
or U9966 (N_9966,N_6801,N_6628);
nand U9967 (N_9967,N_6082,N_5370);
xnor U9968 (N_9968,N_6757,N_5551);
nor U9969 (N_9969,N_7072,N_7461);
nand U9970 (N_9970,N_5785,N_5819);
and U9971 (N_9971,N_6025,N_6478);
and U9972 (N_9972,N_5283,N_5645);
or U9973 (N_9973,N_7481,N_5308);
and U9974 (N_9974,N_5014,N_5911);
nand U9975 (N_9975,N_5852,N_7203);
nor U9976 (N_9976,N_5157,N_5345);
nand U9977 (N_9977,N_5875,N_5865);
nor U9978 (N_9978,N_5357,N_5598);
and U9979 (N_9979,N_5008,N_6061);
nor U9980 (N_9980,N_7081,N_5741);
xnor U9981 (N_9981,N_6724,N_6515);
nor U9982 (N_9982,N_6593,N_6676);
or U9983 (N_9983,N_5277,N_6837);
and U9984 (N_9984,N_6716,N_6394);
nand U9985 (N_9985,N_5900,N_7412);
and U9986 (N_9986,N_5983,N_5837);
or U9987 (N_9987,N_6940,N_5785);
nor U9988 (N_9988,N_5754,N_6358);
or U9989 (N_9989,N_5462,N_6696);
or U9990 (N_9990,N_5814,N_5178);
nand U9991 (N_9991,N_5925,N_5415);
xor U9992 (N_9992,N_5415,N_6558);
and U9993 (N_9993,N_6290,N_6499);
nor U9994 (N_9994,N_6804,N_5610);
xor U9995 (N_9995,N_5588,N_5011);
or U9996 (N_9996,N_5124,N_5352);
and U9997 (N_9997,N_5818,N_5840);
nand U9998 (N_9998,N_6905,N_5031);
nand U9999 (N_9999,N_5427,N_5634);
or UO_0 (O_0,N_9200,N_8601);
or UO_1 (O_1,N_9551,N_9541);
nor UO_2 (O_2,N_9353,N_9907);
nor UO_3 (O_3,N_8094,N_8118);
xor UO_4 (O_4,N_8827,N_9799);
xnor UO_5 (O_5,N_9729,N_7612);
or UO_6 (O_6,N_7999,N_9593);
nor UO_7 (O_7,N_7972,N_8719);
and UO_8 (O_8,N_9757,N_8133);
or UO_9 (O_9,N_7556,N_8990);
or UO_10 (O_10,N_9616,N_9554);
xor UO_11 (O_11,N_8607,N_7554);
and UO_12 (O_12,N_8101,N_9693);
and UO_13 (O_13,N_7930,N_8218);
nand UO_14 (O_14,N_9039,N_8735);
nor UO_15 (O_15,N_8233,N_9118);
nor UO_16 (O_16,N_8934,N_7818);
nand UO_17 (O_17,N_8740,N_9932);
or UO_18 (O_18,N_8380,N_9972);
nand UO_19 (O_19,N_7873,N_8314);
or UO_20 (O_20,N_9034,N_7949);
and UO_21 (O_21,N_9140,N_9001);
and UO_22 (O_22,N_9243,N_8170);
nor UO_23 (O_23,N_7919,N_8142);
nand UO_24 (O_24,N_9030,N_8761);
or UO_25 (O_25,N_7503,N_9369);
and UO_26 (O_26,N_8364,N_8005);
nor UO_27 (O_27,N_7705,N_9281);
or UO_28 (O_28,N_9786,N_9559);
or UO_29 (O_29,N_9056,N_8489);
xor UO_30 (O_30,N_8894,N_8409);
or UO_31 (O_31,N_8302,N_9457);
and UO_32 (O_32,N_9330,N_7931);
xor UO_33 (O_33,N_9208,N_7951);
and UO_34 (O_34,N_7526,N_9100);
xnor UO_35 (O_35,N_9071,N_9536);
or UO_36 (O_36,N_9015,N_8394);
and UO_37 (O_37,N_8125,N_7610);
nand UO_38 (O_38,N_9641,N_9189);
xnor UO_39 (O_39,N_9721,N_7959);
xnor UO_40 (O_40,N_7865,N_8940);
and UO_41 (O_41,N_7740,N_8199);
and UO_42 (O_42,N_9918,N_9890);
and UO_43 (O_43,N_8318,N_7805);
xor UO_44 (O_44,N_9855,N_8109);
nor UO_45 (O_45,N_7633,N_9660);
xor UO_46 (O_46,N_8344,N_9453);
nand UO_47 (O_47,N_8405,N_8611);
and UO_48 (O_48,N_8411,N_8555);
and UO_49 (O_49,N_9094,N_8419);
or UO_50 (O_50,N_7917,N_9321);
or UO_51 (O_51,N_8643,N_8596);
or UO_52 (O_52,N_7994,N_7542);
nor UO_53 (O_53,N_8283,N_8279);
and UO_54 (O_54,N_9807,N_7684);
xor UO_55 (O_55,N_7769,N_9405);
and UO_56 (O_56,N_9632,N_9078);
or UO_57 (O_57,N_8184,N_7574);
nor UO_58 (O_58,N_7774,N_9867);
or UO_59 (O_59,N_8134,N_7978);
nand UO_60 (O_60,N_8182,N_7726);
or UO_61 (O_61,N_8424,N_7946);
and UO_62 (O_62,N_9154,N_7651);
and UO_63 (O_63,N_7541,N_9639);
and UO_64 (O_64,N_8996,N_9575);
nand UO_65 (O_65,N_9132,N_7645);
nand UO_66 (O_66,N_9813,N_9626);
nor UO_67 (O_67,N_8030,N_7883);
or UO_68 (O_68,N_8738,N_8725);
and UO_69 (O_69,N_9089,N_8703);
or UO_70 (O_70,N_9621,N_7591);
nand UO_71 (O_71,N_8259,N_9199);
xnor UO_72 (O_72,N_8965,N_9506);
nand UO_73 (O_73,N_8228,N_9422);
nand UO_74 (O_74,N_7785,N_8463);
or UO_75 (O_75,N_7636,N_9215);
or UO_76 (O_76,N_8169,N_8888);
and UO_77 (O_77,N_9230,N_9274);
nand UO_78 (O_78,N_7665,N_8048);
nor UO_79 (O_79,N_9882,N_7844);
or UO_80 (O_80,N_9066,N_8285);
nand UO_81 (O_81,N_9017,N_9194);
xor UO_82 (O_82,N_7950,N_9112);
or UO_83 (O_83,N_7565,N_9964);
nor UO_84 (O_84,N_9360,N_9863);
or UO_85 (O_85,N_7581,N_9682);
and UO_86 (O_86,N_8253,N_8350);
and UO_87 (O_87,N_7657,N_9550);
nor UO_88 (O_88,N_9052,N_9270);
nor UO_89 (O_89,N_9432,N_9679);
nor UO_90 (O_90,N_9856,N_8274);
nand UO_91 (O_91,N_7830,N_7587);
and UO_92 (O_92,N_9691,N_8771);
nand UO_93 (O_93,N_8426,N_8494);
nand UO_94 (O_94,N_9012,N_8904);
nand UO_95 (O_95,N_9183,N_9257);
and UO_96 (O_96,N_8537,N_9700);
or UO_97 (O_97,N_9305,N_8053);
or UO_98 (O_98,N_7788,N_7906);
and UO_99 (O_99,N_8924,N_8869);
and UO_100 (O_100,N_9595,N_7647);
or UO_101 (O_101,N_7653,N_8078);
nor UO_102 (O_102,N_9351,N_9553);
nand UO_103 (O_103,N_9149,N_9563);
nor UO_104 (O_104,N_9711,N_9607);
xor UO_105 (O_105,N_8251,N_9436);
nor UO_106 (O_106,N_9180,N_8821);
or UO_107 (O_107,N_8986,N_8379);
nor UO_108 (O_108,N_7870,N_9776);
nor UO_109 (O_109,N_7695,N_9887);
nor UO_110 (O_110,N_9759,N_8785);
nor UO_111 (O_111,N_9386,N_8363);
nor UO_112 (O_112,N_8261,N_9143);
nor UO_113 (O_113,N_9620,N_9343);
and UO_114 (O_114,N_8993,N_8896);
and UO_115 (O_115,N_8187,N_8640);
and UO_116 (O_116,N_8820,N_8324);
xnor UO_117 (O_117,N_9892,N_8520);
nand UO_118 (O_118,N_9467,N_9894);
and UO_119 (O_119,N_8626,N_7558);
xnor UO_120 (O_120,N_9710,N_9774);
nand UO_121 (O_121,N_8576,N_7583);
nand UO_122 (O_122,N_7842,N_8737);
nor UO_123 (O_123,N_8296,N_8544);
xor UO_124 (O_124,N_9528,N_9852);
and UO_125 (O_125,N_9433,N_8646);
nor UO_126 (O_126,N_9440,N_8083);
nor UO_127 (O_127,N_7517,N_8110);
and UO_128 (O_128,N_9081,N_9673);
xor UO_129 (O_129,N_9513,N_8830);
xor UO_130 (O_130,N_7791,N_9771);
or UO_131 (O_131,N_9119,N_7613);
nand UO_132 (O_132,N_9950,N_8009);
and UO_133 (O_133,N_9372,N_8875);
nand UO_134 (O_134,N_8399,N_8977);
nor UO_135 (O_135,N_9597,N_8967);
or UO_136 (O_136,N_8167,N_9323);
nor UO_137 (O_137,N_7758,N_8683);
and UO_138 (O_138,N_7981,N_8829);
nor UO_139 (O_139,N_7660,N_8352);
nor UO_140 (O_140,N_7577,N_7955);
nor UO_141 (O_141,N_8981,N_8443);
or UO_142 (O_142,N_9058,N_9242);
or UO_143 (O_143,N_7886,N_7545);
nor UO_144 (O_144,N_7929,N_9451);
xor UO_145 (O_145,N_7736,N_7845);
and UO_146 (O_146,N_7685,N_9581);
or UO_147 (O_147,N_9051,N_7979);
or UO_148 (O_148,N_9619,N_9886);
and UO_149 (O_149,N_8839,N_7520);
nand UO_150 (O_150,N_7834,N_8526);
or UO_151 (O_151,N_9308,N_9885);
nand UO_152 (O_152,N_8024,N_7802);
or UO_153 (O_153,N_7722,N_9955);
and UO_154 (O_154,N_9625,N_8874);
and UO_155 (O_155,N_9198,N_9136);
nor UO_156 (O_156,N_7836,N_8288);
nor UO_157 (O_157,N_7773,N_9831);
nand UO_158 (O_158,N_9511,N_7719);
or UO_159 (O_159,N_9879,N_8408);
nand UO_160 (O_160,N_8516,N_8256);
nand UO_161 (O_161,N_8201,N_8868);
nor UO_162 (O_162,N_9333,N_9121);
nor UO_163 (O_163,N_9181,N_8211);
or UO_164 (O_164,N_8151,N_9135);
or UO_165 (O_165,N_8594,N_7553);
or UO_166 (O_166,N_9795,N_8480);
xor UO_167 (O_167,N_9901,N_9168);
nor UO_168 (O_168,N_9779,N_9310);
or UO_169 (O_169,N_8268,N_8698);
and UO_170 (O_170,N_8770,N_7627);
nand UO_171 (O_171,N_8671,N_8615);
nand UO_172 (O_172,N_9289,N_8673);
and UO_173 (O_173,N_8695,N_9127);
nand UO_174 (O_174,N_8776,N_9778);
nor UO_175 (O_175,N_9772,N_9096);
nand UO_176 (O_176,N_9296,N_8124);
nor UO_177 (O_177,N_9787,N_8402);
and UO_178 (O_178,N_8921,N_8326);
nor UO_179 (O_179,N_9282,N_8734);
nand UO_180 (O_180,N_9941,N_7888);
and UO_181 (O_181,N_8747,N_8759);
and UO_182 (O_182,N_9789,N_8714);
nor UO_183 (O_183,N_9961,N_7837);
or UO_184 (O_184,N_8027,N_8751);
nand UO_185 (O_185,N_9104,N_9000);
or UO_186 (O_186,N_8926,N_8997);
or UO_187 (O_187,N_9207,N_8858);
and UO_188 (O_188,N_8081,N_8205);
nor UO_189 (O_189,N_7913,N_7884);
nand UO_190 (O_190,N_8757,N_7743);
and UO_191 (O_191,N_8389,N_9830);
nand UO_192 (O_192,N_9288,N_9611);
or UO_193 (O_193,N_9615,N_9072);
nor UO_194 (O_194,N_7829,N_8107);
or UO_195 (O_195,N_8456,N_9917);
nand UO_196 (O_196,N_8286,N_7516);
nor UO_197 (O_197,N_9490,N_8885);
nand UO_198 (O_198,N_8597,N_8100);
or UO_199 (O_199,N_8795,N_9283);
and UO_200 (O_200,N_9010,N_7815);
nor UO_201 (O_201,N_7759,N_9820);
xnor UO_202 (O_202,N_8964,N_7625);
or UO_203 (O_203,N_9500,N_9426);
or UO_204 (O_204,N_9661,N_8119);
nand UO_205 (O_205,N_9290,N_8447);
nor UO_206 (O_206,N_8844,N_8095);
nor UO_207 (O_207,N_8928,N_9322);
nand UO_208 (O_208,N_8741,N_9853);
xnor UO_209 (O_209,N_8733,N_8828);
and UO_210 (O_210,N_9562,N_9249);
nor UO_211 (O_211,N_7847,N_9319);
nand UO_212 (O_212,N_8299,N_7854);
nor UO_213 (O_213,N_7808,N_9683);
nand UO_214 (O_214,N_8250,N_9442);
or UO_215 (O_215,N_7980,N_8451);
xor UO_216 (O_216,N_8814,N_8290);
nand UO_217 (O_217,N_9148,N_8718);
and UO_218 (O_218,N_9746,N_7650);
and UO_219 (O_219,N_9702,N_7717);
nor UO_220 (O_220,N_8649,N_7857);
or UO_221 (O_221,N_7954,N_8912);
and UO_222 (O_222,N_8680,N_9416);
nor UO_223 (O_223,N_9601,N_8598);
and UO_224 (O_224,N_7973,N_9443);
and UO_225 (O_225,N_9745,N_9508);
and UO_226 (O_226,N_9291,N_7760);
or UO_227 (O_227,N_7535,N_8554);
and UO_228 (O_228,N_7851,N_9124);
nor UO_229 (O_229,N_8907,N_9596);
and UO_230 (O_230,N_7524,N_8152);
and UO_231 (O_231,N_7895,N_8386);
or UO_232 (O_232,N_7598,N_9927);
nand UO_233 (O_233,N_8758,N_9473);
and UO_234 (O_234,N_9864,N_7504);
nor UO_235 (O_235,N_7661,N_9031);
nand UO_236 (O_236,N_9828,N_9099);
or UO_237 (O_237,N_8841,N_7920);
or UO_238 (O_238,N_8323,N_7584);
xnor UO_239 (O_239,N_8700,N_9184);
or UO_240 (O_240,N_7536,N_8273);
and UO_241 (O_241,N_8730,N_9752);
and UO_242 (O_242,N_8238,N_8836);
nand UO_243 (O_243,N_9086,N_9401);
or UO_244 (O_244,N_9061,N_9365);
or UO_245 (O_245,N_9966,N_8879);
or UO_246 (O_246,N_9874,N_8944);
or UO_247 (O_247,N_9331,N_9994);
nand UO_248 (O_248,N_7778,N_9675);
nand UO_249 (O_249,N_8085,N_8023);
nand UO_250 (O_250,N_7751,N_8739);
and UO_251 (O_251,N_9672,N_8724);
or UO_252 (O_252,N_8527,N_9743);
nor UO_253 (O_253,N_9507,N_9431);
or UO_254 (O_254,N_9793,N_9413);
or UO_255 (O_255,N_9999,N_9712);
nor UO_256 (O_256,N_8754,N_8383);
and UO_257 (O_257,N_9844,N_9638);
nor UO_258 (O_258,N_8635,N_7640);
nor UO_259 (O_259,N_7654,N_9279);
and UO_260 (O_260,N_8662,N_8374);
and UO_261 (O_261,N_8307,N_8400);
nor UO_262 (O_262,N_8512,N_9465);
or UO_263 (O_263,N_9047,N_9788);
nand UO_264 (O_264,N_9872,N_7995);
nand UO_265 (O_265,N_7694,N_7668);
or UO_266 (O_266,N_8128,N_9007);
and UO_267 (O_267,N_9841,N_8452);
or UO_268 (O_268,N_9309,N_9042);
and UO_269 (O_269,N_9583,N_8701);
or UO_270 (O_270,N_9839,N_8353);
nand UO_271 (O_271,N_8528,N_9750);
nand UO_272 (O_272,N_8331,N_9645);
or UO_273 (O_273,N_9258,N_9904);
nand UO_274 (O_274,N_7772,N_9880);
nand UO_275 (O_275,N_7875,N_7820);
and UO_276 (O_276,N_8854,N_9307);
xnor UO_277 (O_277,N_9128,N_7700);
or UO_278 (O_278,N_8506,N_9354);
nor UO_279 (O_279,N_9598,N_8316);
nor UO_280 (O_280,N_9824,N_8864);
or UO_281 (O_281,N_8059,N_7643);
or UO_282 (O_282,N_8974,N_9400);
nor UO_283 (O_283,N_7666,N_9898);
or UO_284 (O_284,N_7530,N_7787);
or UO_285 (O_285,N_7605,N_9387);
nor UO_286 (O_286,N_9869,N_9582);
or UO_287 (O_287,N_8918,N_7702);
and UO_288 (O_288,N_8441,N_8049);
or UO_289 (O_289,N_8459,N_8599);
or UO_290 (O_290,N_8750,N_8391);
nor UO_291 (O_291,N_9870,N_9805);
nand UO_292 (O_292,N_8393,N_8946);
or UO_293 (O_293,N_8280,N_9566);
and UO_294 (O_294,N_8521,N_9133);
nand UO_295 (O_295,N_9934,N_8219);
or UO_296 (O_296,N_8255,N_9816);
nand UO_297 (O_297,N_7992,N_8927);
or UO_298 (O_298,N_7540,N_7988);
or UO_299 (O_299,N_8191,N_8123);
nor UO_300 (O_300,N_8689,N_8901);
or UO_301 (O_301,N_9647,N_7589);
nor UO_302 (O_302,N_8158,N_8265);
or UO_303 (O_303,N_7925,N_7531);
nand UO_304 (O_304,N_8478,N_8705);
nor UO_305 (O_305,N_8475,N_9464);
nor UO_306 (O_306,N_9669,N_7922);
nor UO_307 (O_307,N_9804,N_8312);
nor UO_308 (O_308,N_7623,N_8486);
and UO_309 (O_309,N_8192,N_9263);
and UO_310 (O_310,N_9703,N_8315);
or UO_311 (O_311,N_7877,N_9951);
xnor UO_312 (O_312,N_7916,N_7548);
nand UO_313 (O_313,N_9106,N_8444);
nand UO_314 (O_314,N_9605,N_8498);
nand UO_315 (O_315,N_9614,N_7576);
nor UO_316 (O_316,N_9476,N_9460);
or UO_317 (O_317,N_7986,N_9916);
nor UO_318 (O_318,N_8212,N_9299);
xnor UO_319 (O_319,N_9969,N_9547);
nor UO_320 (O_320,N_7699,N_9130);
nor UO_321 (O_321,N_8668,N_9809);
nand UO_322 (O_322,N_7510,N_9923);
nor UO_323 (O_323,N_8726,N_9285);
nand UO_324 (O_324,N_9744,N_8214);
nand UO_325 (O_325,N_8018,N_8873);
nand UO_326 (O_326,N_8077,N_9742);
xor UO_327 (O_327,N_9835,N_8347);
nor UO_328 (O_328,N_9618,N_8306);
and UO_329 (O_329,N_9803,N_9722);
xor UO_330 (O_330,N_8710,N_9740);
nand UO_331 (O_331,N_8473,N_8271);
and UO_332 (O_332,N_9568,N_9931);
nor UO_333 (O_333,N_9524,N_9990);
or UO_334 (O_334,N_9849,N_7745);
nand UO_335 (O_335,N_8849,N_9069);
nand UO_336 (O_336,N_9084,N_7567);
or UO_337 (O_337,N_9585,N_7855);
or UO_338 (O_338,N_7741,N_7659);
and UO_339 (O_339,N_8210,N_8566);
or UO_340 (O_340,N_8417,N_7638);
nor UO_341 (O_341,N_8308,N_8482);
and UO_342 (O_342,N_9261,N_8064);
nand UO_343 (O_343,N_9439,N_8908);
nand UO_344 (O_344,N_8106,N_9512);
nor UO_345 (O_345,N_7796,N_8816);
or UO_346 (O_346,N_9032,N_9093);
and UO_347 (O_347,N_9138,N_9810);
and UO_348 (O_348,N_8588,N_8242);
nand UO_349 (O_349,N_9687,N_9197);
or UO_350 (O_350,N_9662,N_7572);
nor UO_351 (O_351,N_9948,N_7580);
nand UO_352 (O_352,N_9062,N_8509);
nand UO_353 (O_353,N_9264,N_9794);
nand UO_354 (O_354,N_7593,N_8621);
and UO_355 (O_355,N_9876,N_7761);
and UO_356 (O_356,N_9303,N_9812);
and UO_357 (O_357,N_8434,N_7770);
nor UO_358 (O_358,N_8892,N_8044);
nand UO_359 (O_359,N_8975,N_8295);
xnor UO_360 (O_360,N_9371,N_7826);
nor UO_361 (O_361,N_8817,N_8179);
xor UO_362 (O_362,N_9368,N_8942);
or UO_363 (O_363,N_9156,N_7846);
nand UO_364 (O_364,N_8507,N_8088);
nor UO_365 (O_365,N_8970,N_7506);
or UO_366 (O_366,N_9067,N_7940);
nor UO_367 (O_367,N_9602,N_8999);
nand UO_368 (O_368,N_8254,N_8641);
nand UO_369 (O_369,N_8846,N_8438);
nor UO_370 (O_370,N_7944,N_7961);
or UO_371 (O_371,N_8608,N_9250);
nor UO_372 (O_372,N_9385,N_9642);
or UO_373 (O_373,N_9760,N_9908);
nand UO_374 (O_374,N_9983,N_9748);
or UO_375 (O_375,N_9680,N_8861);
and UO_376 (O_376,N_9022,N_7968);
and UO_377 (O_377,N_7667,N_7914);
and UO_378 (O_378,N_8373,N_8867);
or UO_379 (O_379,N_9195,N_8960);
nand UO_380 (O_380,N_9185,N_8232);
nand UO_381 (O_381,N_9196,N_7566);
or UO_382 (O_382,N_9228,N_8462);
and UO_383 (O_383,N_9122,N_9463);
xor UO_384 (O_384,N_9609,N_8209);
and UO_385 (O_385,N_9686,N_8230);
nor UO_386 (O_386,N_8222,N_8881);
and UO_387 (O_387,N_8172,N_7910);
or UO_388 (O_388,N_8782,N_9026);
nor UO_389 (O_389,N_7941,N_9373);
and UO_390 (O_390,N_8863,N_8831);
nor UO_391 (O_391,N_8072,N_8160);
and UO_392 (O_392,N_9651,N_8269);
or UO_393 (O_393,N_9718,N_7676);
and UO_394 (O_394,N_9589,N_9671);
and UO_395 (O_395,N_9260,N_9091);
and UO_396 (O_396,N_9569,N_8382);
and UO_397 (O_397,N_9986,N_8040);
xnor UO_398 (O_398,N_9978,N_9311);
xor UO_399 (O_399,N_8173,N_9244);
or UO_400 (O_400,N_7849,N_7915);
nor UO_401 (O_401,N_8272,N_9800);
nand UO_402 (O_402,N_8561,N_9201);
and UO_403 (O_403,N_9688,N_8045);
nor UO_404 (O_404,N_9977,N_8529);
or UO_405 (O_405,N_8213,N_8291);
nor UO_406 (O_406,N_8181,N_9781);
and UO_407 (O_407,N_8345,N_9095);
nand UO_408 (O_408,N_8141,N_8017);
nor UO_409 (O_409,N_8633,N_7544);
or UO_410 (O_410,N_7555,N_9998);
or UO_411 (O_411,N_9957,N_8859);
or UO_412 (O_412,N_8050,N_9161);
nor UO_413 (O_413,N_9306,N_8574);
and UO_414 (O_414,N_9499,N_7756);
xnor UO_415 (O_415,N_9477,N_7711);
nand UO_416 (O_416,N_8356,N_9796);
nand UO_417 (O_417,N_8978,N_7797);
and UO_418 (O_418,N_9170,N_8126);
or UO_419 (O_419,N_7786,N_8398);
or UO_420 (O_420,N_9806,N_8385);
nor UO_421 (O_421,N_9576,N_9048);
or UO_422 (O_422,N_7840,N_9055);
nor UO_423 (O_423,N_9173,N_8440);
or UO_424 (O_424,N_8342,N_7742);
or UO_425 (O_425,N_9151,N_7579);
or UO_426 (O_426,N_8371,N_9006);
xor UO_427 (O_427,N_7943,N_9734);
nand UO_428 (O_428,N_8401,N_9738);
or UO_429 (O_429,N_8721,N_8029);
nor UO_430 (O_430,N_8736,N_7532);
nand UO_431 (O_431,N_9783,N_9259);
nand UO_432 (O_432,N_8013,N_7853);
or UO_433 (O_433,N_8973,N_9802);
and UO_434 (O_434,N_8466,N_7880);
nand UO_435 (O_435,N_8235,N_9418);
or UO_436 (O_436,N_8267,N_7582);
nand UO_437 (O_437,N_8961,N_7921);
nor UO_438 (O_438,N_9267,N_9567);
and UO_439 (O_439,N_8546,N_9224);
or UO_440 (O_440,N_8176,N_9177);
nand UO_441 (O_441,N_9580,N_9574);
nand UO_442 (O_442,N_8129,N_8573);
nor UO_443 (O_443,N_9921,N_8991);
or UO_444 (O_444,N_9954,N_8247);
nor UO_445 (O_445,N_7814,N_8805);
nand UO_446 (O_446,N_7551,N_8925);
or UO_447 (O_447,N_8629,N_9819);
and UO_448 (O_448,N_8772,N_7680);
and UO_449 (O_449,N_8847,N_9176);
and UO_450 (O_450,N_9340,N_8972);
nand UO_451 (O_451,N_7908,N_9233);
and UO_452 (O_452,N_7681,N_7896);
nand UO_453 (O_453,N_8749,N_9367);
or UO_454 (O_454,N_7527,N_8204);
nand UO_455 (O_455,N_7618,N_7990);
and UO_456 (O_456,N_9236,N_7969);
and UO_457 (O_457,N_8038,N_9226);
or UO_458 (O_458,N_9996,N_8582);
nor UO_459 (O_459,N_7858,N_9797);
or UO_460 (O_460,N_9544,N_8073);
nor UO_461 (O_461,N_8403,N_9204);
xor UO_462 (O_462,N_8800,N_7804);
nand UO_463 (O_463,N_9667,N_9469);
nand UO_464 (O_464,N_8609,N_9868);
and UO_465 (O_465,N_9036,N_9696);
and UO_466 (O_466,N_8369,N_9773);
xor UO_467 (O_467,N_8556,N_9492);
nand UO_468 (O_468,N_8062,N_9107);
xnor UO_469 (O_469,N_9801,N_9137);
or UO_470 (O_470,N_8500,N_9145);
and UO_471 (O_471,N_8012,N_7869);
nand UO_472 (O_472,N_8667,N_9389);
nor UO_473 (O_473,N_8939,N_8819);
nand UO_474 (O_474,N_8935,N_9613);
and UO_475 (O_475,N_7856,N_9504);
xor UO_476 (O_476,N_9527,N_8390);
and UO_477 (O_477,N_7885,N_8055);
nand UO_478 (O_478,N_7771,N_7909);
xnor UO_479 (O_479,N_9262,N_9848);
and UO_480 (O_480,N_9780,N_7614);
or UO_481 (O_481,N_9540,N_8810);
and UO_482 (O_482,N_7515,N_9555);
or UO_483 (O_483,N_7603,N_8445);
nand UO_484 (O_484,N_8697,N_8485);
nor UO_485 (O_485,N_9903,N_7803);
or UO_486 (O_486,N_7655,N_8327);
xor UO_487 (O_487,N_8508,N_7575);
and UO_488 (O_488,N_9014,N_8684);
and UO_489 (O_489,N_8548,N_8190);
or UO_490 (O_490,N_9029,N_9650);
and UO_491 (O_491,N_9142,N_7521);
nor UO_492 (O_492,N_9753,N_9754);
or UO_493 (O_493,N_8889,N_8499);
nand UO_494 (O_494,N_8876,N_8784);
xnor UO_495 (O_495,N_9286,N_7891);
and UO_496 (O_496,N_9287,N_9798);
and UO_497 (O_497,N_9939,N_9370);
xnor UO_498 (O_498,N_9792,N_8430);
and UO_499 (O_499,N_8992,N_9505);
nor UO_500 (O_500,N_9097,N_8769);
and UO_501 (O_501,N_9345,N_8033);
and UO_502 (O_502,N_8026,N_9973);
nor UO_503 (O_503,N_9116,N_8808);
nand UO_504 (O_504,N_9294,N_7731);
nand UO_505 (O_505,N_8429,N_9775);
and UO_506 (O_506,N_7790,N_7958);
and UO_507 (O_507,N_9732,N_9277);
nor UO_508 (O_508,N_8098,N_8571);
nand UO_509 (O_509,N_8605,N_8835);
nand UO_510 (O_510,N_9946,N_9967);
nor UO_511 (O_511,N_8407,N_9493);
nand UO_512 (O_512,N_9486,N_9355);
or UO_513 (O_513,N_9325,N_8037);
nand UO_514 (O_514,N_7898,N_9338);
and UO_515 (O_515,N_8843,N_9393);
nand UO_516 (O_516,N_9412,N_8897);
nand UO_517 (O_517,N_9944,N_9989);
xnor UO_518 (O_518,N_9980,N_9942);
nand UO_519 (O_519,N_7674,N_7887);
or UO_520 (O_520,N_8616,N_9375);
nor UO_521 (O_521,N_8263,N_8144);
nand UO_522 (O_522,N_8905,N_8663);
or UO_523 (O_523,N_9063,N_8577);
xnor UO_524 (O_524,N_7528,N_8236);
or UO_525 (O_525,N_7635,N_8852);
xor UO_526 (O_526,N_8166,N_7936);
or UO_527 (O_527,N_9475,N_8822);
and UO_528 (O_528,N_9975,N_9157);
nand UO_529 (O_529,N_8781,N_9077);
xnor UO_530 (O_530,N_9214,N_9455);
nor UO_531 (O_531,N_8948,N_9211);
and UO_532 (O_532,N_7683,N_9068);
nor UO_533 (O_533,N_8976,N_9182);
nor UO_534 (O_534,N_9139,N_8448);
nor UO_535 (O_535,N_9163,N_8837);
nand UO_536 (O_536,N_9737,N_7689);
nand UO_537 (O_537,N_8479,N_9899);
nor UO_538 (O_538,N_8681,N_8322);
nor UO_539 (O_539,N_9704,N_9314);
nor UO_540 (O_540,N_8748,N_9021);
nand UO_541 (O_541,N_9708,N_9720);
or UO_542 (O_542,N_8047,N_8336);
and UO_543 (O_543,N_7718,N_8234);
nand UO_544 (O_544,N_7724,N_9845);
nor UO_545 (O_545,N_7996,N_8541);
nand UO_546 (O_546,N_8774,N_9008);
nor UO_547 (O_547,N_9390,N_9922);
nor UO_548 (O_548,N_9266,N_9115);
or UO_549 (O_549,N_8636,N_8370);
nand UO_550 (O_550,N_8161,N_7586);
nor UO_551 (O_551,N_8777,N_9024);
or UO_552 (O_552,N_8330,N_8941);
nor UO_553 (O_553,N_9350,N_9947);
or UO_554 (O_554,N_9357,N_8414);
and UO_555 (O_555,N_9044,N_8922);
nand UO_556 (O_556,N_9377,N_7983);
and UO_557 (O_557,N_9222,N_9730);
or UO_558 (O_558,N_8538,N_9076);
and UO_559 (O_559,N_7902,N_7602);
and UO_560 (O_560,N_8533,N_8021);
and UO_561 (O_561,N_9040,N_7500);
or UO_562 (O_562,N_9352,N_8226);
and UO_563 (O_563,N_7867,N_8131);
nand UO_564 (O_564,N_9991,N_9216);
or UO_565 (O_565,N_7890,N_8560);
nor UO_566 (O_566,N_8593,N_7632);
nor UO_567 (O_567,N_9186,N_9103);
nor UO_568 (O_568,N_8804,N_9035);
or UO_569 (O_569,N_9082,N_9612);
or UO_570 (O_570,N_8058,N_9764);
nand UO_571 (O_571,N_9060,N_7809);
nand UO_572 (O_572,N_8900,N_8642);
xor UO_573 (O_573,N_8792,N_8620);
and UO_574 (O_574,N_9080,N_9846);
nor UO_575 (O_575,N_9817,N_8378);
or UO_576 (O_576,N_9891,N_8084);
or UO_577 (O_577,N_8959,N_8206);
nor UO_578 (O_578,N_8449,N_8054);
nand UO_579 (O_579,N_8360,N_8634);
nand UO_580 (O_580,N_9971,N_9328);
and UO_581 (O_581,N_9420,N_9984);
and UO_582 (O_582,N_9379,N_8632);
or UO_583 (O_583,N_8693,N_8335);
or UO_584 (O_584,N_8262,N_8034);
nor UO_585 (O_585,N_9041,N_7713);
and UO_586 (O_586,N_9153,N_9573);
and UO_587 (O_587,N_9532,N_8534);
and UO_588 (O_588,N_9239,N_9016);
and UO_589 (O_589,N_8971,N_7518);
nand UO_590 (O_590,N_9397,N_9374);
nand UO_591 (O_591,N_7701,N_8000);
nand UO_592 (O_592,N_8916,N_9529);
nor UO_593 (O_593,N_8917,N_8032);
and UO_594 (O_594,N_8148,N_9920);
nor UO_595 (O_595,N_9491,N_7606);
nand UO_596 (O_596,N_9866,N_8862);
xor UO_597 (O_597,N_8060,N_8592);
nor UO_598 (O_598,N_9326,N_7889);
and UO_599 (O_599,N_8174,N_7952);
and UO_600 (O_600,N_7573,N_8604);
and UO_601 (O_601,N_8035,N_7905);
nor UO_602 (O_602,N_8276,N_8791);
or UO_603 (O_603,N_9538,N_7646);
nor UO_604 (O_604,N_8461,N_7799);
xnor UO_605 (O_605,N_8984,N_9447);
and UO_606 (O_606,N_8687,N_8711);
or UO_607 (O_607,N_8303,N_8264);
and UO_608 (O_608,N_7843,N_9509);
or UO_609 (O_609,N_7671,N_8224);
nand UO_610 (O_610,N_8305,N_9533);
and UO_611 (O_611,N_9535,N_9495);
and UO_612 (O_612,N_8328,N_8146);
nor UO_613 (O_613,N_9109,N_9050);
nor UO_614 (O_614,N_9915,N_8248);
and UO_615 (O_615,N_8982,N_7947);
nor UO_616 (O_616,N_8911,N_9152);
and UO_617 (O_617,N_8071,N_9826);
nor UO_618 (O_618,N_8937,N_8183);
or UO_619 (O_619,N_7562,N_9640);
xor UO_620 (O_620,N_7817,N_8783);
or UO_621 (O_621,N_9456,N_8956);
nand UO_622 (O_622,N_8707,N_9965);
nand UO_623 (O_623,N_7609,N_9292);
nor UO_624 (O_624,N_7993,N_9560);
and UO_625 (O_625,N_7833,N_9502);
or UO_626 (O_626,N_7879,N_9902);
and UO_627 (O_627,N_8117,N_8292);
nor UO_628 (O_628,N_9111,N_9543);
and UO_629 (O_629,N_8065,N_7714);
nor UO_630 (O_630,N_7729,N_7823);
nor UO_631 (O_631,N_8731,N_8833);
nor UO_632 (O_632,N_9425,N_7734);
and UO_633 (O_633,N_8773,N_9192);
nor UO_634 (O_634,N_8838,N_8715);
nor UO_635 (O_635,N_8717,N_8557);
or UO_636 (O_636,N_7764,N_9539);
nor UO_637 (O_637,N_9485,N_9537);
xnor UO_638 (O_638,N_8428,N_7942);
nor UO_639 (O_639,N_8502,N_7537);
nand UO_640 (O_640,N_9938,N_8493);
nand UO_641 (O_641,N_7578,N_9087);
nor UO_642 (O_642,N_8293,N_8834);
xnor UO_643 (O_643,N_8627,N_8171);
nand UO_644 (O_644,N_8229,N_9976);
nand UO_645 (O_645,N_9677,N_9606);
xor UO_646 (O_646,N_8872,N_7876);
nor UO_647 (O_647,N_7564,N_8439);
xor UO_648 (O_648,N_9516,N_8648);
or UO_649 (O_649,N_7766,N_8614);
and UO_650 (O_650,N_8909,N_9234);
nand UO_651 (O_651,N_9689,N_9335);
or UO_652 (O_652,N_9430,N_8969);
and UO_653 (O_653,N_9468,N_9332);
nor UO_654 (O_654,N_9295,N_9818);
nand UO_655 (O_655,N_8052,N_8732);
xnor UO_656 (O_656,N_8366,N_7864);
nor UO_657 (O_657,N_9404,N_9329);
or UO_658 (O_658,N_7596,N_8531);
and UO_659 (O_659,N_8240,N_7715);
or UO_660 (O_660,N_9896,N_7810);
nand UO_661 (O_661,N_8468,N_8583);
nor UO_662 (O_662,N_9437,N_9346);
nor UO_663 (O_663,N_9318,N_9755);
nor UO_664 (O_664,N_8082,N_9462);
nor UO_665 (O_665,N_8079,N_8309);
nor UO_666 (O_666,N_7686,N_8138);
or UO_667 (O_667,N_9349,N_8780);
nor UO_668 (O_668,N_7508,N_9565);
or UO_669 (O_669,N_8674,N_9479);
and UO_670 (O_670,N_8664,N_9248);
or UO_671 (O_671,N_7934,N_8850);
and UO_672 (O_672,N_9150,N_8551);
nand UO_673 (O_673,N_8678,N_8388);
and UO_674 (O_674,N_9587,N_9815);
and UO_675 (O_675,N_8676,N_7639);
nand UO_676 (O_676,N_8728,N_8216);
and UO_677 (O_677,N_8985,N_8137);
and UO_678 (O_678,N_9503,N_8584);
nand UO_679 (O_679,N_9247,N_8763);
and UO_680 (O_680,N_8069,N_8579);
or UO_681 (O_681,N_8086,N_8767);
nor UO_682 (O_682,N_8865,N_9488);
and UO_683 (O_683,N_7502,N_8099);
or UO_684 (O_684,N_8797,N_9603);
nand UO_685 (O_685,N_8421,N_9843);
or UO_686 (O_686,N_7819,N_9217);
nand UO_687 (O_687,N_9952,N_9736);
and UO_688 (O_688,N_7670,N_8105);
nand UO_689 (O_689,N_8910,N_8530);
or UO_690 (O_690,N_8252,N_7893);
nor UO_691 (O_691,N_9785,N_8660);
and UO_692 (O_692,N_8963,N_9827);
nor UO_693 (O_693,N_7511,N_9459);
nor UO_694 (O_694,N_8121,N_7512);
or UO_695 (O_695,N_9220,N_9699);
or UO_696 (O_696,N_8022,N_7776);
and UO_697 (O_697,N_7704,N_8351);
and UO_698 (O_698,N_9716,N_8497);
or UO_699 (O_699,N_8031,N_9070);
nand UO_700 (O_700,N_8578,N_9079);
and UO_701 (O_701,N_8416,N_9435);
and UO_702 (O_702,N_8727,N_8061);
nor UO_703 (O_703,N_8706,N_8188);
nand UO_704 (O_704,N_9438,N_8692);
or UO_705 (O_705,N_8657,N_9428);
nor UO_706 (O_706,N_9735,N_9271);
nand UO_707 (O_707,N_7514,N_7737);
nor UO_708 (O_708,N_7534,N_8540);
and UO_709 (O_709,N_8798,N_8275);
and UO_710 (O_710,N_9454,N_9458);
and UO_711 (O_711,N_8310,N_9594);
and UO_712 (O_712,N_9893,N_8647);
or UO_713 (O_713,N_8041,N_9557);
xnor UO_714 (O_714,N_9275,N_7757);
and UO_715 (O_715,N_9963,N_9359);
or UO_716 (O_716,N_8329,N_7801);
nand UO_717 (O_717,N_7827,N_8207);
nand UO_718 (O_718,N_8930,N_9019);
nor UO_719 (O_719,N_8289,N_9945);
and UO_720 (O_720,N_9770,N_9391);
nor UO_721 (O_721,N_8756,N_8655);
nand UO_722 (O_722,N_7522,N_8460);
nor UO_723 (O_723,N_8477,N_9510);
or UO_724 (O_724,N_8260,N_9085);
nand UO_725 (O_725,N_9162,N_8622);
xor UO_726 (O_726,N_7881,N_8492);
or UO_727 (O_727,N_9668,N_7529);
nand UO_728 (O_728,N_9579,N_9147);
and UO_729 (O_729,N_9501,N_8650);
nand UO_730 (O_730,N_9429,N_9530);
and UO_731 (O_731,N_8565,N_7648);
or UO_732 (O_732,N_7782,N_9655);
nand UO_733 (O_733,N_8523,N_9125);
or UO_734 (O_734,N_9376,N_9304);
and UO_735 (O_735,N_8337,N_7546);
nand UO_736 (O_736,N_7703,N_9825);
or UO_737 (O_737,N_8418,N_7821);
nor UO_738 (O_738,N_9993,N_9466);
xnor UO_739 (O_739,N_9474,N_9895);
or UO_740 (O_740,N_8185,N_7991);
and UO_741 (O_741,N_9909,N_8752);
or UO_742 (O_742,N_9424,N_9223);
nand UO_743 (O_743,N_8368,N_8422);
or UO_744 (O_744,N_9949,N_8003);
xnor UO_745 (O_745,N_7693,N_9758);
and UO_746 (O_746,N_8704,N_8656);
and UO_747 (O_747,N_9378,N_7629);
and UO_748 (O_748,N_7569,N_9556);
nor UO_749 (O_749,N_8481,N_8610);
xor UO_750 (O_750,N_8890,N_7677);
nand UO_751 (O_751,N_8938,N_7927);
nand UO_752 (O_752,N_8197,N_8087);
or UO_753 (O_753,N_8425,N_9448);
or UO_754 (O_754,N_7621,N_7746);
nor UO_755 (O_755,N_8458,N_9630);
xor UO_756 (O_756,N_8962,N_7707);
nor UO_757 (O_757,N_7767,N_9246);
nor UO_758 (O_758,N_9850,N_7811);
nand UO_759 (O_759,N_9525,N_7539);
nand UO_760 (O_760,N_9985,N_7594);
or UO_761 (O_761,N_8281,N_8690);
and UO_762 (O_762,N_8920,N_8221);
or UO_763 (O_763,N_7900,N_7904);
or UO_764 (O_764,N_7533,N_9713);
and UO_765 (O_765,N_8568,N_8535);
or UO_766 (O_766,N_9570,N_7557);
or UO_767 (O_767,N_7903,N_8474);
and UO_768 (O_768,N_9727,N_7617);
nand UO_769 (O_769,N_9608,N_9470);
or UO_770 (O_770,N_9883,N_7507);
nor UO_771 (O_771,N_7779,N_8539);
nand UO_772 (O_772,N_8665,N_9427);
xnor UO_773 (O_773,N_8090,N_8338);
nand UO_774 (O_774,N_8745,N_8760);
xor UO_775 (O_775,N_8321,N_9496);
or UO_776 (O_776,N_9114,N_8848);
or UO_777 (O_777,N_8536,N_9414);
nor UO_778 (O_778,N_8702,N_9232);
nand UO_779 (O_779,N_8755,N_9497);
and UO_780 (O_780,N_9756,N_9861);
xnor UO_781 (O_781,N_9862,N_8341);
xnor UO_782 (O_782,N_7798,N_9784);
nor UO_783 (O_783,N_9045,N_8433);
and UO_784 (O_784,N_8708,N_7732);
and UO_785 (O_785,N_8454,N_7607);
nor UO_786 (O_786,N_9191,N_9705);
nand UO_787 (O_787,N_9146,N_9252);
nand UO_788 (O_788,N_7987,N_9765);
and UO_789 (O_789,N_9237,N_9715);
or UO_790 (O_790,N_9255,N_9417);
nor UO_791 (O_791,N_8004,N_8672);
nor UO_792 (O_792,N_9578,N_9273);
nor UO_793 (O_793,N_8168,N_9494);
and UO_794 (O_794,N_8949,N_9698);
nor UO_795 (O_795,N_9187,N_7848);
nor UO_796 (O_796,N_9717,N_8287);
or UO_797 (O_797,N_8149,N_7622);
nor UO_798 (O_798,N_9751,N_8688);
or UO_799 (O_799,N_8779,N_9212);
nand UO_800 (O_800,N_8801,N_9654);
nor UO_801 (O_801,N_8068,N_8006);
nand UO_802 (O_802,N_7784,N_7728);
xnor UO_803 (O_803,N_8524,N_8947);
and UO_804 (O_804,N_8423,N_9483);
xor UO_805 (O_805,N_9073,N_9723);
and UO_806 (O_806,N_9623,N_9160);
or UO_807 (O_807,N_8397,N_8572);
and UO_808 (O_808,N_9004,N_9545);
or UO_809 (O_809,N_8104,N_8122);
and UO_810 (O_810,N_7730,N_9900);
and UO_811 (O_811,N_8504,N_8547);
or UO_812 (O_812,N_9202,N_9415);
or UO_813 (O_813,N_9808,N_9617);
or UO_814 (O_814,N_9518,N_9498);
nand UO_815 (O_815,N_7692,N_9167);
nor UO_816 (O_816,N_8076,N_8880);
or UO_817 (O_817,N_8567,N_8933);
or UO_818 (O_818,N_8015,N_9117);
nand UO_819 (O_819,N_8070,N_8487);
xnor UO_820 (O_820,N_9053,N_8856);
and UO_821 (O_821,N_8612,N_9213);
nor UO_822 (O_822,N_9384,N_7965);
nor UO_823 (O_823,N_7560,N_9179);
and UO_824 (O_824,N_9919,N_9933);
and UO_825 (O_825,N_9591,N_8215);
nor UO_826 (O_826,N_9171,N_7828);
nor UO_827 (O_827,N_8446,N_8699);
nand UO_828 (O_828,N_8659,N_8130);
nor UO_829 (O_829,N_8175,N_8147);
nand UO_830 (O_830,N_9395,N_8789);
and UO_831 (O_831,N_9043,N_8359);
nand UO_832 (O_832,N_9126,N_9854);
and UO_833 (O_833,N_8115,N_9449);
or UO_834 (O_834,N_7822,N_7727);
nor UO_835 (O_835,N_8644,N_8712);
nand UO_836 (O_836,N_8613,N_8136);
or UO_837 (O_837,N_8164,N_8325);
and UO_838 (O_838,N_7971,N_8066);
and UO_839 (O_839,N_7841,N_8348);
nand UO_840 (O_840,N_8595,N_7525);
or UO_841 (O_841,N_9013,N_8899);
or UO_842 (O_842,N_7571,N_9571);
nand UO_843 (O_843,N_7813,N_9166);
or UO_844 (O_844,N_8813,N_9480);
nor UO_845 (O_845,N_9388,N_8806);
nand UO_846 (O_846,N_9684,N_9564);
xor UO_847 (O_847,N_9878,N_7832);
or UO_848 (O_848,N_8513,N_8395);
or UO_849 (O_849,N_8958,N_9144);
or UO_850 (O_850,N_9225,N_7747);
or UO_851 (O_851,N_7616,N_8645);
nand UO_852 (O_852,N_7604,N_8339);
and UO_853 (O_853,N_9158,N_9123);
nor UO_854 (O_854,N_7644,N_9175);
and UO_855 (O_855,N_8766,N_9419);
or UO_856 (O_856,N_7982,N_9877);
nor UO_857 (O_857,N_9546,N_9633);
or UO_858 (O_858,N_8367,N_8787);
nor UO_859 (O_859,N_9120,N_8679);
nor UO_860 (O_860,N_8120,N_9837);
nand UO_861 (O_861,N_8957,N_8853);
and UO_862 (O_862,N_7709,N_8915);
or UO_863 (O_863,N_8510,N_9937);
and UO_864 (O_864,N_8437,N_9622);
or UO_865 (O_865,N_7775,N_9251);
nand UO_866 (O_866,N_8812,N_8624);
or UO_867 (O_867,N_9873,N_7956);
and UO_868 (O_868,N_8096,N_8143);
nand UO_869 (O_869,N_7675,N_8108);
xnor UO_870 (O_870,N_8016,N_9659);
and UO_871 (O_871,N_9670,N_7563);
and UO_872 (O_872,N_9728,N_7871);
or UO_873 (O_873,N_9858,N_9658);
or UO_874 (O_874,N_9600,N_8796);
nor UO_875 (O_875,N_9206,N_8694);
and UO_876 (O_876,N_9134,N_9241);
nand UO_877 (O_877,N_9871,N_8723);
or UO_878 (O_878,N_8159,N_7637);
and UO_879 (O_879,N_9635,N_8011);
nor UO_880 (O_880,N_8768,N_7924);
nand UO_881 (O_881,N_9749,N_9960);
xor UO_882 (O_882,N_7783,N_9763);
xor UO_883 (O_883,N_9534,N_8282);
and UO_884 (O_884,N_8270,N_8637);
or UO_885 (O_885,N_8135,N_7907);
xnor UO_886 (O_886,N_8413,N_8488);
nor UO_887 (O_887,N_9707,N_8628);
nand UO_888 (O_888,N_8127,N_9790);
nor UO_889 (O_889,N_9714,N_8112);
and UO_890 (O_890,N_9542,N_8455);
or UO_891 (O_891,N_8617,N_9782);
or UO_892 (O_892,N_7619,N_9218);
or UO_893 (O_893,N_8802,N_8332);
xnor UO_894 (O_894,N_8471,N_8923);
nor UO_895 (O_895,N_8845,N_7825);
nor UO_896 (O_896,N_7592,N_8818);
or UO_897 (O_897,N_8762,N_7777);
nand UO_898 (O_898,N_7899,N_9090);
and UO_899 (O_899,N_9974,N_9381);
xnor UO_900 (O_900,N_9982,N_9092);
or UO_901 (O_901,N_8998,N_9690);
xnor UO_902 (O_902,N_8929,N_8132);
or UO_903 (O_903,N_9240,N_8484);
and UO_904 (O_904,N_8691,N_8193);
and UO_905 (O_905,N_9652,N_9366);
nor UO_906 (O_906,N_8075,N_7698);
and UO_907 (O_907,N_9113,N_9958);
xor UO_908 (O_908,N_9884,N_8936);
xnor UO_909 (O_909,N_8898,N_7620);
nand UO_910 (O_910,N_9777,N_8377);
nor UO_911 (O_911,N_7552,N_8177);
and UO_912 (O_912,N_9685,N_7860);
or UO_913 (O_913,N_9724,N_7662);
or UO_914 (O_914,N_9472,N_9762);
and UO_915 (O_915,N_8300,N_9694);
nor UO_916 (O_916,N_7935,N_7800);
or UO_917 (O_917,N_9471,N_7866);
nand UO_918 (O_918,N_9231,N_7624);
or UO_919 (O_919,N_9159,N_8476);
and UO_920 (O_920,N_9356,N_9209);
or UO_921 (O_921,N_8415,N_8196);
nor UO_922 (O_922,N_8882,N_8361);
or UO_923 (O_923,N_9098,N_9558);
and UO_924 (O_924,N_9320,N_7977);
nand UO_925 (O_925,N_7682,N_9190);
and UO_926 (O_926,N_8505,N_9924);
and UO_927 (O_927,N_8340,N_8580);
nand UO_928 (O_928,N_7696,N_7669);
xor UO_929 (O_929,N_7824,N_8319);
and UO_930 (O_930,N_8658,N_7652);
and UO_931 (O_931,N_9174,N_7831);
nor UO_932 (O_932,N_8317,N_9347);
nand UO_933 (O_933,N_9995,N_8840);
or UO_934 (O_934,N_8490,N_8165);
or UO_935 (O_935,N_8884,N_9300);
nand UO_936 (O_936,N_9968,N_9636);
and UO_937 (O_937,N_9656,N_7505);
nand UO_938 (O_938,N_8102,N_7549);
and UO_939 (O_939,N_8542,N_9697);
or UO_940 (O_940,N_7806,N_7945);
or UO_941 (O_941,N_9410,N_8155);
or UO_942 (O_942,N_8056,N_9588);
or UO_943 (O_943,N_8581,N_7733);
nand UO_944 (O_944,N_8951,N_9674);
nor UO_945 (O_945,N_8294,N_9889);
nor UO_946 (O_946,N_9037,N_7748);
nor UO_947 (O_947,N_8113,N_9337);
or UO_948 (O_948,N_8775,N_8720);
and UO_949 (O_949,N_7750,N_9521);
nor UO_950 (O_950,N_9522,N_8298);
nor UO_951 (O_951,N_9268,N_8435);
or UO_952 (O_952,N_9926,N_9444);
and UO_953 (O_953,N_8189,N_8020);
or UO_954 (O_954,N_9131,N_9407);
nor UO_955 (O_955,N_8284,N_9101);
and UO_956 (O_956,N_9382,N_9398);
or UO_957 (O_957,N_8010,N_7874);
xnor UO_958 (O_958,N_9577,N_9649);
nor UO_959 (O_959,N_9421,N_8931);
nor UO_960 (O_960,N_8220,N_9905);
and UO_961 (O_961,N_8051,N_8682);
nand UO_962 (O_962,N_8223,N_7708);
nor UO_963 (O_963,N_7588,N_8586);
xor UO_964 (O_964,N_7568,N_9906);
and UO_965 (O_965,N_9910,N_8729);
xnor UO_966 (O_966,N_8803,N_8569);
xor UO_967 (O_967,N_7816,N_7762);
nor UO_968 (O_968,N_9881,N_8217);
nand UO_969 (O_969,N_8543,N_7754);
and UO_970 (O_970,N_8570,N_8995);
nand UO_971 (O_971,N_8677,N_7868);
or UO_972 (O_972,N_7679,N_8713);
xnor UO_973 (O_973,N_8313,N_7673);
or UO_974 (O_974,N_8431,N_9678);
and UO_975 (O_975,N_9484,N_8346);
xor UO_976 (O_976,N_7812,N_7523);
and UO_977 (O_977,N_9461,N_9912);
nor UO_978 (O_978,N_7912,N_8522);
and UO_979 (O_979,N_9627,N_7585);
or UO_980 (O_980,N_8764,N_8587);
xnor UO_981 (O_981,N_8525,N_7656);
and UO_982 (O_982,N_9992,N_9832);
or UO_983 (O_983,N_8815,N_7725);
and UO_984 (O_984,N_9065,N_7780);
or UO_985 (O_985,N_8007,N_8811);
and UO_986 (O_986,N_9188,N_9666);
nand UO_987 (O_987,N_7501,N_7911);
nor UO_988 (O_988,N_8950,N_7957);
nand UO_989 (O_989,N_9327,N_7835);
or UO_990 (O_990,N_8799,N_8495);
nor UO_991 (O_991,N_9851,N_9833);
nor UO_992 (O_992,N_9269,N_9074);
nor UO_993 (O_993,N_7710,N_8245);
nor UO_994 (O_994,N_8793,N_9836);
nor UO_995 (O_995,N_7649,N_8427);
nand UO_996 (O_996,N_7795,N_8406);
and UO_997 (O_997,N_9033,N_9489);
or UO_998 (O_998,N_7852,N_8832);
xor UO_999 (O_999,N_9011,N_8661);
xnor UO_1000 (O_1000,N_8375,N_8150);
nand UO_1001 (O_1001,N_8778,N_9701);
nor UO_1002 (O_1002,N_9731,N_9105);
and UO_1003 (O_1003,N_9059,N_9075);
xor UO_1004 (O_1004,N_8093,N_9361);
nand UO_1005 (O_1005,N_8716,N_9434);
or UO_1006 (O_1006,N_8953,N_9997);
nor UO_1007 (O_1007,N_9324,N_9057);
or UO_1008 (O_1008,N_9811,N_9129);
nor UO_1009 (O_1009,N_9719,N_8465);
xor UO_1010 (O_1010,N_8381,N_9838);
and UO_1011 (O_1011,N_9219,N_8914);
and UO_1012 (O_1012,N_8412,N_9364);
nor UO_1013 (O_1013,N_7975,N_9411);
or UO_1014 (O_1014,N_9888,N_7976);
nor UO_1015 (O_1015,N_7600,N_8025);
nand UO_1016 (O_1016,N_9561,N_8932);
and UO_1017 (O_1017,N_8686,N_8866);
or UO_1018 (O_1018,N_9339,N_8008);
nor UO_1019 (O_1019,N_9814,N_9403);
and UO_1020 (O_1020,N_8063,N_9875);
nor UO_1021 (O_1021,N_7753,N_8036);
nor UO_1022 (O_1022,N_9312,N_8968);
nand UO_1023 (O_1023,N_9834,N_8491);
or UO_1024 (O_1024,N_8392,N_9298);
xor UO_1025 (O_1025,N_7998,N_8955);
nand UO_1026 (O_1026,N_9929,N_7739);
or UO_1027 (O_1027,N_9930,N_7690);
nand UO_1028 (O_1028,N_9979,N_9519);
xnor UO_1029 (O_1029,N_7626,N_7631);
xor UO_1030 (O_1030,N_9747,N_9383);
and UO_1031 (O_1031,N_8067,N_8154);
or UO_1032 (O_1032,N_9478,N_8619);
or UO_1033 (O_1033,N_9631,N_9766);
nand UO_1034 (O_1034,N_7839,N_8563);
or UO_1035 (O_1035,N_8517,N_8194);
nand UO_1036 (O_1036,N_8623,N_9610);
nor UO_1037 (O_1037,N_8744,N_8590);
or UO_1038 (O_1038,N_8826,N_8410);
or UO_1039 (O_1039,N_8809,N_7989);
and UO_1040 (O_1040,N_9653,N_7630);
nand UO_1041 (O_1041,N_8195,N_9165);
nand UO_1042 (O_1042,N_9238,N_9396);
or UO_1043 (O_1043,N_8532,N_9637);
nand UO_1044 (O_1044,N_8111,N_8092);
xnor UO_1045 (O_1045,N_9842,N_7597);
nand UO_1046 (O_1046,N_9695,N_7933);
and UO_1047 (O_1047,N_8870,N_7720);
or UO_1048 (O_1048,N_8603,N_9399);
or UO_1049 (O_1049,N_8943,N_9003);
nand UO_1050 (O_1050,N_9083,N_8983);
or UO_1051 (O_1051,N_9038,N_7781);
nor UO_1052 (O_1052,N_7892,N_9341);
and UO_1053 (O_1053,N_8585,N_7964);
xor UO_1054 (O_1054,N_9970,N_9987);
nand UO_1055 (O_1055,N_7561,N_8602);
or UO_1056 (O_1056,N_8722,N_9023);
and UO_1057 (O_1057,N_8652,N_9344);
and UO_1058 (O_1058,N_8631,N_8186);
nand UO_1059 (O_1059,N_8358,N_8301);
xnor UO_1060 (O_1060,N_8362,N_9394);
and UO_1061 (O_1061,N_9108,N_8200);
or UO_1062 (O_1062,N_8472,N_9221);
nand UO_1063 (O_1063,N_9302,N_9859);
or UO_1064 (O_1064,N_8297,N_9392);
and UO_1065 (O_1065,N_8266,N_8355);
and UO_1066 (O_1066,N_7878,N_8618);
xor UO_1067 (O_1067,N_9590,N_8945);
or UO_1068 (O_1068,N_7763,N_7901);
or UO_1069 (O_1069,N_7861,N_9005);
xnor UO_1070 (O_1070,N_8675,N_7664);
xnor UO_1071 (O_1071,N_7663,N_7749);
nand UO_1072 (O_1072,N_8157,N_8638);
nand UO_1073 (O_1073,N_8919,N_9002);
nor UO_1074 (O_1074,N_9336,N_9681);
nor UO_1075 (O_1075,N_7706,N_8753);
and UO_1076 (O_1076,N_8420,N_9334);
and UO_1077 (O_1077,N_9768,N_9054);
or UO_1078 (O_1078,N_8042,N_9726);
and UO_1079 (O_1079,N_8562,N_8788);
and UO_1080 (O_1080,N_7960,N_9531);
and UO_1081 (O_1081,N_9523,N_8320);
nor UO_1082 (O_1082,N_8243,N_9205);
nand UO_1083 (O_1083,N_9925,N_9769);
xnor UO_1084 (O_1084,N_8989,N_8824);
or UO_1085 (O_1085,N_9028,N_8515);
xor UO_1086 (O_1086,N_7789,N_9709);
and UO_1087 (O_1087,N_8503,N_7538);
nor UO_1088 (O_1088,N_8354,N_8074);
nand UO_1089 (O_1089,N_9599,N_9110);
or UO_1090 (O_1090,N_7974,N_8891);
nand UO_1091 (O_1091,N_8871,N_9914);
nand UO_1092 (O_1092,N_9018,N_9928);
nor UO_1093 (O_1093,N_8043,N_9940);
and UO_1094 (O_1094,N_8514,N_7697);
nand UO_1095 (O_1095,N_9821,N_9276);
nor UO_1096 (O_1096,N_8227,N_9936);
and UO_1097 (O_1097,N_8954,N_8246);
nand UO_1098 (O_1098,N_8842,N_7672);
nor UO_1099 (O_1099,N_8913,N_9648);
xnor UO_1100 (O_1100,N_7918,N_8387);
xnor UO_1101 (O_1101,N_7948,N_9317);
nand UO_1102 (O_1102,N_8002,N_8855);
and UO_1103 (O_1103,N_8442,N_9229);
and UO_1104 (O_1104,N_8333,N_8825);
and UO_1105 (O_1105,N_9064,N_9840);
nand UO_1106 (O_1106,N_8028,N_9646);
nor UO_1107 (O_1107,N_8046,N_8483);
nor UO_1108 (O_1108,N_7590,N_9254);
nor UO_1109 (O_1109,N_9245,N_9409);
nand UO_1110 (O_1110,N_8887,N_9141);
nand UO_1111 (O_1111,N_7628,N_8278);
and UO_1112 (O_1112,N_8496,N_7938);
or UO_1113 (O_1113,N_9913,N_8786);
or UO_1114 (O_1114,N_8966,N_9515);
and UO_1115 (O_1115,N_9102,N_7966);
or UO_1116 (O_1116,N_8553,N_8591);
and UO_1117 (O_1117,N_9009,N_8878);
or UO_1118 (O_1118,N_7970,N_9278);
nand UO_1119 (O_1119,N_9342,N_8153);
and UO_1120 (O_1120,N_9860,N_8343);
and UO_1121 (O_1121,N_7985,N_8670);
nor UO_1122 (O_1122,N_8666,N_7519);
nor UO_1123 (O_1123,N_8349,N_8039);
xor UO_1124 (O_1124,N_8860,N_7687);
nor UO_1125 (O_1125,N_9358,N_9592);
and UO_1126 (O_1126,N_7608,N_9548);
and UO_1127 (O_1127,N_8396,N_8019);
or UO_1128 (O_1128,N_7926,N_8198);
or UO_1129 (O_1129,N_8180,N_8883);
or UO_1130 (O_1130,N_9301,N_8501);
nand UO_1131 (O_1131,N_7615,N_9959);
nor UO_1132 (O_1132,N_8208,N_8987);
nor UO_1133 (O_1133,N_8511,N_8549);
nor UO_1134 (O_1134,N_9911,N_7550);
and UO_1135 (O_1135,N_8902,N_8080);
or UO_1136 (O_1136,N_8372,N_7738);
nor UO_1137 (O_1137,N_9897,N_9604);
and UO_1138 (O_1138,N_8857,N_7658);
and UO_1139 (O_1139,N_9741,N_8980);
or UO_1140 (O_1140,N_9088,N_7939);
or UO_1141 (O_1141,N_9445,N_8014);
or UO_1142 (O_1142,N_9935,N_9441);
xnor UO_1143 (O_1143,N_9549,N_8794);
nand UO_1144 (O_1144,N_9450,N_8225);
and UO_1145 (O_1145,N_8384,N_7543);
nor UO_1146 (O_1146,N_8651,N_7547);
nor UO_1147 (O_1147,N_7642,N_8453);
nor UO_1148 (O_1148,N_9847,N_8630);
and UO_1149 (O_1149,N_7932,N_8163);
nor UO_1150 (O_1150,N_8162,N_8625);
and UO_1151 (O_1151,N_8746,N_8575);
and UO_1152 (O_1152,N_9761,N_8519);
and UO_1153 (O_1153,N_9172,N_9981);
xnor UO_1154 (O_1154,N_9293,N_9227);
nor UO_1155 (O_1155,N_7928,N_9315);
nand UO_1156 (O_1156,N_9235,N_9584);
and UO_1157 (O_1157,N_8807,N_8241);
and UO_1158 (O_1158,N_9164,N_7723);
nand UO_1159 (O_1159,N_7634,N_7678);
nor UO_1160 (O_1160,N_9253,N_9169);
nor UO_1161 (O_1161,N_7793,N_9178);
or UO_1162 (O_1162,N_7599,N_9956);
and UO_1163 (O_1163,N_9663,N_9676);
or UO_1164 (O_1164,N_8545,N_9193);
nor UO_1165 (O_1165,N_8237,N_8450);
or UO_1166 (O_1166,N_9210,N_8231);
nand UO_1167 (O_1167,N_9514,N_8559);
or UO_1168 (O_1168,N_8765,N_9348);
or UO_1169 (O_1169,N_8558,N_9572);
nand UO_1170 (O_1170,N_8139,N_9423);
nand UO_1171 (O_1171,N_8464,N_9552);
nand UO_1172 (O_1172,N_8304,N_9865);
nor UO_1173 (O_1173,N_8089,N_8685);
xor UO_1174 (O_1174,N_9526,N_9025);
and UO_1175 (O_1175,N_8518,N_9706);
nor UO_1176 (O_1176,N_8114,N_7601);
nand UO_1177 (O_1177,N_8001,N_9586);
xnor UO_1178 (O_1178,N_9297,N_7744);
and UO_1179 (O_1179,N_8893,N_8669);
nor UO_1180 (O_1180,N_9272,N_9643);
or UO_1181 (O_1181,N_9049,N_8906);
nor UO_1182 (O_1182,N_8357,N_9446);
nand UO_1183 (O_1183,N_7712,N_9953);
nand UO_1184 (O_1184,N_8654,N_8696);
nand UO_1185 (O_1185,N_8257,N_8552);
nand UO_1186 (O_1186,N_8249,N_9155);
nor UO_1187 (O_1187,N_7963,N_8116);
nand UO_1188 (O_1188,N_8877,N_9020);
xnor UO_1189 (O_1189,N_7859,N_8952);
xor UO_1190 (O_1190,N_7559,N_8145);
nor UO_1191 (O_1191,N_8404,N_8258);
nand UO_1192 (O_1192,N_7838,N_8277);
xnor UO_1193 (O_1193,N_9256,N_8823);
nor UO_1194 (O_1194,N_8091,N_7882);
and UO_1195 (O_1195,N_7691,N_8886);
xnor UO_1196 (O_1196,N_7721,N_9988);
nor UO_1197 (O_1197,N_8790,N_8470);
nand UO_1198 (O_1198,N_9634,N_8436);
nand UO_1199 (O_1199,N_7997,N_7688);
xnor UO_1200 (O_1200,N_8550,N_8589);
and UO_1201 (O_1201,N_8639,N_9767);
and UO_1202 (O_1202,N_8097,N_9380);
or UO_1203 (O_1203,N_7735,N_7872);
and UO_1204 (O_1204,N_9402,N_7984);
nor UO_1205 (O_1205,N_9027,N_8653);
and UO_1206 (O_1206,N_9284,N_9517);
nor UO_1207 (O_1207,N_9406,N_7937);
nor UO_1208 (O_1208,N_9316,N_8709);
and UO_1209 (O_1209,N_8178,N_8103);
nor UO_1210 (O_1210,N_8467,N_8742);
nand UO_1211 (O_1211,N_9943,N_8334);
nand UO_1212 (O_1212,N_7894,N_8851);
and UO_1213 (O_1213,N_9823,N_8564);
and UO_1214 (O_1214,N_8988,N_7765);
xnor UO_1215 (O_1215,N_9481,N_8743);
or UO_1216 (O_1216,N_9313,N_7513);
and UO_1217 (O_1217,N_7863,N_7641);
or UO_1218 (O_1218,N_7768,N_7953);
and UO_1219 (O_1219,N_8365,N_9046);
and UO_1220 (O_1220,N_8311,N_8432);
nand UO_1221 (O_1221,N_8376,N_8239);
and UO_1222 (O_1222,N_7752,N_8203);
nor UO_1223 (O_1223,N_7897,N_8469);
xnor UO_1224 (O_1224,N_9203,N_9725);
or UO_1225 (O_1225,N_9362,N_9822);
or UO_1226 (O_1226,N_7923,N_7807);
nand UO_1227 (O_1227,N_7716,N_8994);
and UO_1228 (O_1228,N_9733,N_8606);
xnor UO_1229 (O_1229,N_8979,N_9482);
or UO_1230 (O_1230,N_9265,N_7792);
nand UO_1231 (O_1231,N_8057,N_9739);
nand UO_1232 (O_1232,N_8202,N_9692);
nor UO_1233 (O_1233,N_7509,N_9624);
nand UO_1234 (O_1234,N_9520,N_9857);
and UO_1235 (O_1235,N_8156,N_9664);
and UO_1236 (O_1236,N_7755,N_8903);
nor UO_1237 (O_1237,N_9962,N_9280);
and UO_1238 (O_1238,N_7570,N_8457);
and UO_1239 (O_1239,N_7611,N_8244);
nor UO_1240 (O_1240,N_7794,N_9363);
or UO_1241 (O_1241,N_7967,N_8140);
or UO_1242 (O_1242,N_9829,N_9628);
xnor UO_1243 (O_1243,N_8600,N_7862);
xnor UO_1244 (O_1244,N_9644,N_9791);
nand UO_1245 (O_1245,N_8895,N_9629);
nor UO_1246 (O_1246,N_9408,N_9487);
or UO_1247 (O_1247,N_9657,N_7962);
xnor UO_1248 (O_1248,N_9665,N_9452);
or UO_1249 (O_1249,N_7595,N_7850);
or UO_1250 (O_1250,N_7893,N_9083);
and UO_1251 (O_1251,N_9287,N_8187);
or UO_1252 (O_1252,N_9101,N_8676);
nor UO_1253 (O_1253,N_9082,N_9007);
nand UO_1254 (O_1254,N_9600,N_9559);
nand UO_1255 (O_1255,N_9466,N_9183);
nor UO_1256 (O_1256,N_8036,N_9622);
or UO_1257 (O_1257,N_7917,N_7674);
nand UO_1258 (O_1258,N_9067,N_8428);
xnor UO_1259 (O_1259,N_8172,N_9536);
or UO_1260 (O_1260,N_9854,N_7917);
nor UO_1261 (O_1261,N_9788,N_8946);
nand UO_1262 (O_1262,N_8092,N_7728);
nand UO_1263 (O_1263,N_9668,N_9170);
nor UO_1264 (O_1264,N_9838,N_9708);
xnor UO_1265 (O_1265,N_9107,N_9188);
or UO_1266 (O_1266,N_8825,N_8507);
or UO_1267 (O_1267,N_8718,N_8240);
or UO_1268 (O_1268,N_9119,N_9412);
nor UO_1269 (O_1269,N_8712,N_9866);
nor UO_1270 (O_1270,N_8883,N_7900);
and UO_1271 (O_1271,N_8978,N_8547);
and UO_1272 (O_1272,N_8275,N_7976);
nand UO_1273 (O_1273,N_9840,N_8975);
nor UO_1274 (O_1274,N_8002,N_7860);
and UO_1275 (O_1275,N_8212,N_9903);
and UO_1276 (O_1276,N_8243,N_9057);
nand UO_1277 (O_1277,N_8165,N_8039);
or UO_1278 (O_1278,N_8288,N_9191);
nor UO_1279 (O_1279,N_8446,N_7737);
nor UO_1280 (O_1280,N_8690,N_8841);
or UO_1281 (O_1281,N_8934,N_9637);
xor UO_1282 (O_1282,N_7858,N_8791);
and UO_1283 (O_1283,N_8515,N_8969);
xnor UO_1284 (O_1284,N_9603,N_9590);
nor UO_1285 (O_1285,N_7603,N_9540);
nand UO_1286 (O_1286,N_9349,N_8241);
and UO_1287 (O_1287,N_8771,N_8170);
and UO_1288 (O_1288,N_9505,N_9707);
nor UO_1289 (O_1289,N_8349,N_7844);
and UO_1290 (O_1290,N_8346,N_7778);
and UO_1291 (O_1291,N_8851,N_7914);
nand UO_1292 (O_1292,N_7519,N_9166);
and UO_1293 (O_1293,N_9435,N_9584);
nand UO_1294 (O_1294,N_7788,N_7831);
or UO_1295 (O_1295,N_9366,N_9103);
nor UO_1296 (O_1296,N_9715,N_8297);
nor UO_1297 (O_1297,N_8834,N_8623);
nor UO_1298 (O_1298,N_9639,N_7924);
xnor UO_1299 (O_1299,N_9939,N_9145);
nor UO_1300 (O_1300,N_9265,N_7648);
nand UO_1301 (O_1301,N_9381,N_7533);
nand UO_1302 (O_1302,N_7704,N_9950);
nor UO_1303 (O_1303,N_8499,N_8274);
nor UO_1304 (O_1304,N_9355,N_7898);
nor UO_1305 (O_1305,N_9968,N_8174);
xnor UO_1306 (O_1306,N_9631,N_8599);
or UO_1307 (O_1307,N_9728,N_8875);
nor UO_1308 (O_1308,N_9332,N_7607);
nor UO_1309 (O_1309,N_8092,N_8826);
nor UO_1310 (O_1310,N_7645,N_7696);
nand UO_1311 (O_1311,N_8931,N_9514);
or UO_1312 (O_1312,N_7928,N_9746);
xnor UO_1313 (O_1313,N_9757,N_8658);
nor UO_1314 (O_1314,N_9854,N_9846);
xor UO_1315 (O_1315,N_9367,N_9926);
nor UO_1316 (O_1316,N_8812,N_8515);
nand UO_1317 (O_1317,N_7964,N_8140);
and UO_1318 (O_1318,N_9420,N_9418);
or UO_1319 (O_1319,N_8251,N_9677);
or UO_1320 (O_1320,N_8788,N_9494);
nand UO_1321 (O_1321,N_9720,N_9239);
or UO_1322 (O_1322,N_9759,N_7942);
nor UO_1323 (O_1323,N_8643,N_8020);
nand UO_1324 (O_1324,N_7872,N_7574);
nor UO_1325 (O_1325,N_8790,N_9158);
or UO_1326 (O_1326,N_8000,N_9789);
nor UO_1327 (O_1327,N_8118,N_9098);
and UO_1328 (O_1328,N_8610,N_8516);
nand UO_1329 (O_1329,N_8635,N_8518);
and UO_1330 (O_1330,N_8655,N_9675);
and UO_1331 (O_1331,N_7665,N_9106);
nor UO_1332 (O_1332,N_9235,N_8373);
xnor UO_1333 (O_1333,N_8351,N_7975);
nand UO_1334 (O_1334,N_9756,N_9516);
or UO_1335 (O_1335,N_8507,N_8888);
and UO_1336 (O_1336,N_8137,N_7910);
xor UO_1337 (O_1337,N_9801,N_8971);
or UO_1338 (O_1338,N_8492,N_7721);
nor UO_1339 (O_1339,N_8359,N_8228);
or UO_1340 (O_1340,N_9598,N_7888);
xnor UO_1341 (O_1341,N_8728,N_8734);
and UO_1342 (O_1342,N_8648,N_7529);
nand UO_1343 (O_1343,N_7989,N_9825);
and UO_1344 (O_1344,N_9135,N_7872);
xnor UO_1345 (O_1345,N_8691,N_8570);
nor UO_1346 (O_1346,N_9644,N_7902);
or UO_1347 (O_1347,N_8942,N_8047);
nor UO_1348 (O_1348,N_9174,N_9346);
or UO_1349 (O_1349,N_9024,N_9664);
and UO_1350 (O_1350,N_8593,N_8151);
xnor UO_1351 (O_1351,N_8451,N_8873);
or UO_1352 (O_1352,N_7743,N_8105);
and UO_1353 (O_1353,N_9696,N_7652);
or UO_1354 (O_1354,N_9162,N_8880);
or UO_1355 (O_1355,N_7613,N_8586);
nand UO_1356 (O_1356,N_8723,N_7615);
nor UO_1357 (O_1357,N_7776,N_9428);
and UO_1358 (O_1358,N_9615,N_9959);
or UO_1359 (O_1359,N_7872,N_9771);
and UO_1360 (O_1360,N_7997,N_7866);
and UO_1361 (O_1361,N_8177,N_8576);
xor UO_1362 (O_1362,N_8668,N_7791);
and UO_1363 (O_1363,N_8821,N_8376);
and UO_1364 (O_1364,N_7583,N_8922);
and UO_1365 (O_1365,N_8796,N_9731);
and UO_1366 (O_1366,N_9126,N_7990);
nor UO_1367 (O_1367,N_8699,N_7607);
or UO_1368 (O_1368,N_9378,N_8008);
nand UO_1369 (O_1369,N_9054,N_7780);
nand UO_1370 (O_1370,N_7942,N_9656);
xor UO_1371 (O_1371,N_8926,N_8741);
nor UO_1372 (O_1372,N_8759,N_8729);
and UO_1373 (O_1373,N_8295,N_8729);
and UO_1374 (O_1374,N_9654,N_8496);
xnor UO_1375 (O_1375,N_9315,N_8255);
or UO_1376 (O_1376,N_9339,N_8948);
nor UO_1377 (O_1377,N_7984,N_8771);
nand UO_1378 (O_1378,N_9681,N_8003);
or UO_1379 (O_1379,N_7638,N_8467);
nand UO_1380 (O_1380,N_9426,N_8523);
and UO_1381 (O_1381,N_8558,N_8081);
and UO_1382 (O_1382,N_7938,N_8406);
nand UO_1383 (O_1383,N_9250,N_9102);
nand UO_1384 (O_1384,N_7567,N_8662);
and UO_1385 (O_1385,N_8866,N_9126);
nand UO_1386 (O_1386,N_8537,N_8516);
and UO_1387 (O_1387,N_9981,N_8393);
or UO_1388 (O_1388,N_9044,N_9015);
or UO_1389 (O_1389,N_9478,N_9538);
nand UO_1390 (O_1390,N_9151,N_7812);
or UO_1391 (O_1391,N_9700,N_9437);
nor UO_1392 (O_1392,N_7762,N_8034);
xor UO_1393 (O_1393,N_7687,N_8112);
xor UO_1394 (O_1394,N_9378,N_9087);
nand UO_1395 (O_1395,N_9972,N_7978);
xor UO_1396 (O_1396,N_8024,N_9606);
nand UO_1397 (O_1397,N_9829,N_8328);
nor UO_1398 (O_1398,N_8381,N_9528);
nand UO_1399 (O_1399,N_9148,N_8447);
and UO_1400 (O_1400,N_8359,N_9659);
xnor UO_1401 (O_1401,N_8013,N_7818);
or UO_1402 (O_1402,N_7684,N_7891);
or UO_1403 (O_1403,N_8034,N_9225);
and UO_1404 (O_1404,N_8375,N_8085);
nand UO_1405 (O_1405,N_9993,N_9551);
nor UO_1406 (O_1406,N_9342,N_8146);
and UO_1407 (O_1407,N_7615,N_8591);
nor UO_1408 (O_1408,N_9300,N_9629);
xnor UO_1409 (O_1409,N_8187,N_8160);
or UO_1410 (O_1410,N_7755,N_9415);
and UO_1411 (O_1411,N_8105,N_9267);
and UO_1412 (O_1412,N_7850,N_7692);
nand UO_1413 (O_1413,N_9893,N_8590);
or UO_1414 (O_1414,N_7939,N_9901);
and UO_1415 (O_1415,N_9838,N_9642);
nor UO_1416 (O_1416,N_9552,N_9380);
xnor UO_1417 (O_1417,N_7522,N_7635);
and UO_1418 (O_1418,N_9140,N_9542);
and UO_1419 (O_1419,N_9307,N_9735);
xnor UO_1420 (O_1420,N_9077,N_8121);
and UO_1421 (O_1421,N_9688,N_7826);
and UO_1422 (O_1422,N_8373,N_9320);
or UO_1423 (O_1423,N_8393,N_9086);
or UO_1424 (O_1424,N_9011,N_9594);
or UO_1425 (O_1425,N_9466,N_8041);
nor UO_1426 (O_1426,N_8813,N_9543);
and UO_1427 (O_1427,N_9043,N_9444);
and UO_1428 (O_1428,N_8761,N_8194);
and UO_1429 (O_1429,N_9818,N_7898);
nor UO_1430 (O_1430,N_9386,N_8968);
and UO_1431 (O_1431,N_9630,N_8247);
and UO_1432 (O_1432,N_7527,N_7580);
nor UO_1433 (O_1433,N_9641,N_8879);
nand UO_1434 (O_1434,N_8639,N_7635);
nand UO_1435 (O_1435,N_9464,N_9227);
nor UO_1436 (O_1436,N_9050,N_9048);
and UO_1437 (O_1437,N_8380,N_9470);
xor UO_1438 (O_1438,N_9555,N_8699);
and UO_1439 (O_1439,N_7595,N_8221);
or UO_1440 (O_1440,N_9461,N_9649);
or UO_1441 (O_1441,N_7918,N_8774);
or UO_1442 (O_1442,N_9727,N_7777);
nor UO_1443 (O_1443,N_9402,N_9946);
nand UO_1444 (O_1444,N_9864,N_9103);
xnor UO_1445 (O_1445,N_8345,N_7621);
and UO_1446 (O_1446,N_9621,N_7574);
or UO_1447 (O_1447,N_9152,N_9832);
and UO_1448 (O_1448,N_9700,N_7622);
or UO_1449 (O_1449,N_8102,N_8091);
nor UO_1450 (O_1450,N_9363,N_9250);
nor UO_1451 (O_1451,N_8631,N_8964);
nor UO_1452 (O_1452,N_7609,N_8853);
nand UO_1453 (O_1453,N_8227,N_9967);
or UO_1454 (O_1454,N_8774,N_7509);
or UO_1455 (O_1455,N_9585,N_7792);
xor UO_1456 (O_1456,N_7562,N_8972);
xnor UO_1457 (O_1457,N_7590,N_8766);
nor UO_1458 (O_1458,N_9503,N_8272);
xor UO_1459 (O_1459,N_8994,N_7631);
xor UO_1460 (O_1460,N_7509,N_9237);
or UO_1461 (O_1461,N_9602,N_8411);
nand UO_1462 (O_1462,N_9434,N_8715);
nor UO_1463 (O_1463,N_7505,N_8641);
or UO_1464 (O_1464,N_7792,N_9939);
nand UO_1465 (O_1465,N_7743,N_8078);
xor UO_1466 (O_1466,N_7641,N_7557);
nand UO_1467 (O_1467,N_8953,N_9733);
or UO_1468 (O_1468,N_8874,N_7893);
and UO_1469 (O_1469,N_8181,N_8685);
or UO_1470 (O_1470,N_9462,N_7841);
nor UO_1471 (O_1471,N_7875,N_9821);
or UO_1472 (O_1472,N_7569,N_7583);
nand UO_1473 (O_1473,N_8127,N_8970);
nor UO_1474 (O_1474,N_8864,N_9117);
or UO_1475 (O_1475,N_9881,N_9535);
and UO_1476 (O_1476,N_9165,N_8384);
and UO_1477 (O_1477,N_9021,N_9922);
nand UO_1478 (O_1478,N_9467,N_9826);
and UO_1479 (O_1479,N_9990,N_9828);
or UO_1480 (O_1480,N_8556,N_9881);
or UO_1481 (O_1481,N_9353,N_8265);
xnor UO_1482 (O_1482,N_9885,N_8761);
nand UO_1483 (O_1483,N_9995,N_8954);
nand UO_1484 (O_1484,N_8075,N_7710);
or UO_1485 (O_1485,N_8576,N_9846);
nor UO_1486 (O_1486,N_9603,N_7797);
xnor UO_1487 (O_1487,N_8769,N_8298);
nand UO_1488 (O_1488,N_7862,N_8353);
and UO_1489 (O_1489,N_9889,N_9119);
or UO_1490 (O_1490,N_8766,N_8871);
and UO_1491 (O_1491,N_8454,N_8722);
or UO_1492 (O_1492,N_9283,N_8887);
and UO_1493 (O_1493,N_8864,N_9852);
xnor UO_1494 (O_1494,N_7667,N_8340);
nor UO_1495 (O_1495,N_9920,N_9869);
or UO_1496 (O_1496,N_8398,N_8880);
nand UO_1497 (O_1497,N_9421,N_8762);
or UO_1498 (O_1498,N_7649,N_7637);
nand UO_1499 (O_1499,N_8839,N_9344);
endmodule