module basic_2000_20000_2500_80_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1997,In_1570);
nand U1 (N_1,In_1067,In_867);
or U2 (N_2,In_880,In_797);
or U3 (N_3,In_1486,In_67);
or U4 (N_4,In_1422,In_191);
and U5 (N_5,In_466,In_61);
and U6 (N_6,In_1169,In_429);
and U7 (N_7,In_111,In_1758);
and U8 (N_8,In_733,In_1701);
and U9 (N_9,In_1365,In_1960);
nor U10 (N_10,In_113,In_1256);
or U11 (N_11,In_236,In_1465);
nor U12 (N_12,In_1407,In_1456);
or U13 (N_13,In_905,In_785);
nor U14 (N_14,In_1111,In_95);
nor U15 (N_15,In_625,In_655);
nand U16 (N_16,In_1041,In_748);
or U17 (N_17,In_281,In_1385);
nor U18 (N_18,In_1438,In_1770);
nor U19 (N_19,In_842,In_904);
or U20 (N_20,In_1370,In_304);
and U21 (N_21,In_603,In_528);
and U22 (N_22,In_1588,In_1112);
and U23 (N_23,In_1810,In_977);
or U24 (N_24,In_1278,In_1102);
nor U25 (N_25,In_205,In_1554);
nor U26 (N_26,In_18,In_1396);
or U27 (N_27,In_1194,In_162);
or U28 (N_28,In_1190,In_902);
nor U29 (N_29,In_1583,In_317);
nand U30 (N_30,In_632,In_815);
or U31 (N_31,In_1730,In_935);
xnor U32 (N_32,In_1377,In_138);
nor U33 (N_33,In_915,In_1917);
and U34 (N_34,In_13,In_1604);
xnor U35 (N_35,In_523,In_402);
and U36 (N_36,In_1900,In_1071);
or U37 (N_37,In_37,In_1320);
and U38 (N_38,In_1606,In_270);
nand U39 (N_39,In_389,In_1276);
nand U40 (N_40,In_371,In_1781);
or U41 (N_41,In_1192,In_1752);
and U42 (N_42,In_1417,In_1675);
or U43 (N_43,In_810,In_1507);
or U44 (N_44,In_1506,In_386);
and U45 (N_45,In_586,In_519);
nor U46 (N_46,In_1318,In_744);
and U47 (N_47,In_708,In_376);
nand U48 (N_48,In_1187,In_1130);
nand U49 (N_49,In_1826,In_1533);
or U50 (N_50,In_10,In_1799);
nor U51 (N_51,In_1193,In_1938);
nor U52 (N_52,In_241,In_1467);
xnor U53 (N_53,In_1116,In_17);
and U54 (N_54,In_1766,In_231);
nand U55 (N_55,In_722,In_1366);
nor U56 (N_56,In_1692,In_457);
nand U57 (N_57,In_1515,In_1052);
nand U58 (N_58,In_524,In_578);
nand U59 (N_59,In_1633,In_858);
nor U60 (N_60,In_1670,In_1346);
nand U61 (N_61,In_463,In_1062);
or U62 (N_62,In_1085,In_1735);
or U63 (N_63,In_1906,In_151);
nand U64 (N_64,In_1270,In_1844);
xnor U65 (N_65,In_1895,In_1402);
or U66 (N_66,In_57,In_734);
nor U67 (N_67,In_1827,In_984);
nand U68 (N_68,In_1977,In_154);
nand U69 (N_69,In_606,In_213);
xnor U70 (N_70,In_1206,In_1860);
nand U71 (N_71,In_1672,In_1108);
or U72 (N_72,In_1277,In_1582);
or U73 (N_73,In_732,In_366);
and U74 (N_74,In_729,In_1995);
and U75 (N_75,In_547,In_1143);
or U76 (N_76,In_1249,In_653);
and U77 (N_77,In_527,In_594);
or U78 (N_78,In_1879,In_152);
and U79 (N_79,In_752,In_561);
xor U80 (N_80,In_1654,In_484);
nor U81 (N_81,In_778,In_131);
or U82 (N_82,In_1122,In_1261);
nor U83 (N_83,In_1316,In_1949);
nand U84 (N_84,In_677,In_1914);
and U85 (N_85,In_787,In_1403);
and U86 (N_86,In_1980,In_1065);
xnor U87 (N_87,In_1331,In_1353);
nand U88 (N_88,In_1232,In_828);
nand U89 (N_89,In_1129,In_799);
and U90 (N_90,In_983,In_197);
nand U91 (N_91,In_793,In_1535);
or U92 (N_92,In_830,In_1901);
nand U93 (N_93,In_1907,In_1598);
nor U94 (N_94,In_1473,In_1708);
and U95 (N_95,In_1703,In_1098);
or U96 (N_96,In_177,In_262);
nor U97 (N_97,In_1158,In_588);
or U98 (N_98,In_1452,In_1630);
and U99 (N_99,In_1559,In_1220);
or U100 (N_100,In_1020,In_1514);
or U101 (N_101,In_1090,In_607);
nand U102 (N_102,In_692,In_275);
or U103 (N_103,In_314,In_1354);
nand U104 (N_104,In_1406,In_1739);
and U105 (N_105,In_694,In_1121);
nand U106 (N_106,In_1723,In_1266);
and U107 (N_107,In_1873,In_605);
and U108 (N_108,In_772,In_1940);
nor U109 (N_109,In_1573,In_1419);
or U110 (N_110,In_637,In_1092);
and U111 (N_111,In_763,In_237);
nor U112 (N_112,In_1610,In_1449);
nor U113 (N_113,In_1607,In_203);
and U114 (N_114,In_1254,In_453);
xnor U115 (N_115,In_1771,In_760);
and U116 (N_116,In_602,In_1077);
or U117 (N_117,In_1455,In_1795);
and U118 (N_118,In_503,In_207);
or U119 (N_119,In_1728,In_308);
nor U120 (N_120,In_333,In_367);
xnor U121 (N_121,In_1373,In_1155);
or U122 (N_122,In_1942,In_1344);
and U123 (N_123,In_1055,In_1843);
nand U124 (N_124,In_368,In_1897);
nand U125 (N_125,In_1482,In_1841);
and U126 (N_126,In_1097,In_933);
nand U127 (N_127,In_1680,In_344);
or U128 (N_128,In_397,In_633);
nand U129 (N_129,In_516,In_1293);
nand U130 (N_130,In_352,In_1699);
and U131 (N_131,In_265,In_1778);
nor U132 (N_132,In_496,In_592);
and U133 (N_133,In_351,In_583);
and U134 (N_134,In_730,In_318);
and U135 (N_135,In_220,In_669);
nor U136 (N_136,In_914,In_652);
and U137 (N_137,In_341,In_1659);
nor U138 (N_138,In_826,In_409);
nor U139 (N_139,In_443,In_69);
nor U140 (N_140,In_631,In_522);
or U141 (N_141,In_865,In_1773);
nor U142 (N_142,In_1282,In_1528);
and U143 (N_143,In_1635,In_1484);
nand U144 (N_144,In_932,In_992);
nand U145 (N_145,In_1836,In_1095);
and U146 (N_146,In_343,In_767);
nor U147 (N_147,In_814,In_357);
xor U148 (N_148,In_1070,In_739);
nand U149 (N_149,In_1846,In_273);
and U150 (N_150,In_401,In_590);
nand U151 (N_151,In_951,In_1073);
nand U152 (N_152,In_1264,In_1027);
nand U153 (N_153,In_1991,In_1557);
nor U154 (N_154,In_460,In_601);
nand U155 (N_155,In_1265,In_41);
nor U156 (N_156,In_1530,In_1740);
and U157 (N_157,In_1848,In_129);
or U158 (N_158,In_2,In_1527);
or U159 (N_159,In_636,In_1596);
and U160 (N_160,In_664,In_1267);
nor U161 (N_161,In_1896,In_469);
nand U162 (N_162,In_845,In_1600);
xnor U163 (N_163,In_83,In_981);
nand U164 (N_164,In_358,In_1859);
nor U165 (N_165,In_1998,In_1875);
nor U166 (N_166,In_206,In_937);
or U167 (N_167,In_1364,In_759);
or U168 (N_168,In_1281,In_1247);
or U169 (N_169,In_1114,In_1817);
or U170 (N_170,In_1829,In_841);
and U171 (N_171,In_1823,In_1732);
or U172 (N_172,In_78,In_1593);
nand U173 (N_173,In_1315,In_1156);
or U174 (N_174,In_1488,In_682);
nor U175 (N_175,In_155,In_1880);
nor U176 (N_176,In_1602,In_209);
nor U177 (N_177,In_1031,In_577);
nand U178 (N_178,In_1555,In_1919);
or U179 (N_179,In_135,In_657);
xor U180 (N_180,In_1953,In_1131);
nor U181 (N_181,In_986,In_1168);
nor U182 (N_182,In_1054,In_892);
and U183 (N_183,In_1626,In_967);
nor U184 (N_184,In_1132,In_1671);
nor U185 (N_185,In_1648,In_699);
and U186 (N_186,In_611,In_1170);
nand U187 (N_187,In_32,In_824);
and U188 (N_188,In_1549,In_189);
nor U189 (N_189,In_736,In_1024);
xor U190 (N_190,In_1093,In_1500);
nand U191 (N_191,In_753,In_264);
or U192 (N_192,In_1814,In_1704);
nor U193 (N_193,In_1234,In_383);
or U194 (N_194,In_19,In_1013);
nor U195 (N_195,In_473,In_369);
nor U196 (N_196,In_179,In_678);
nor U197 (N_197,In_340,In_1337);
and U198 (N_198,In_1718,In_1138);
and U199 (N_199,In_321,In_1012);
and U200 (N_200,In_1433,In_640);
or U201 (N_201,In_579,In_142);
and U202 (N_202,In_1483,In_1695);
or U203 (N_203,In_1432,In_1601);
nor U204 (N_204,In_966,In_998);
nor U205 (N_205,In_1975,In_844);
and U206 (N_206,In_1643,In_1151);
nand U207 (N_207,In_261,In_315);
nor U208 (N_208,In_1462,In_582);
nor U209 (N_209,In_1308,In_1595);
nor U210 (N_210,In_1043,In_29);
or U211 (N_211,In_1404,In_1461);
nor U212 (N_212,In_489,In_741);
or U213 (N_213,In_1618,In_1932);
xnor U214 (N_214,In_1279,In_1477);
nor U215 (N_215,In_809,In_596);
and U216 (N_216,In_1401,In_1259);
nor U217 (N_217,In_755,In_1238);
or U218 (N_218,In_724,In_433);
or U219 (N_219,In_1059,In_122);
nand U220 (N_220,In_481,In_1979);
nor U221 (N_221,In_866,In_1136);
or U222 (N_222,In_1755,In_773);
nor U223 (N_223,In_686,In_299);
and U224 (N_224,In_477,In_656);
nand U225 (N_225,In_1390,In_768);
or U226 (N_226,In_379,In_249);
and U227 (N_227,In_1541,In_1683);
and U228 (N_228,In_170,In_1805);
or U229 (N_229,In_544,In_1513);
xnor U230 (N_230,In_1963,In_1457);
nand U231 (N_231,In_1288,In_423);
nor U232 (N_232,In_584,In_1894);
xnor U233 (N_233,In_1305,In_491);
nor U234 (N_234,In_1923,In_1347);
nor U235 (N_235,In_923,In_1439);
nor U236 (N_236,In_838,In_794);
nand U237 (N_237,In_176,In_1831);
nor U238 (N_238,In_520,In_1566);
or U239 (N_239,In_1840,In_1682);
xor U240 (N_240,In_202,In_894);
and U241 (N_241,In_381,In_1273);
nor U242 (N_242,In_1389,In_660);
or U243 (N_243,In_46,In_16);
nor U244 (N_244,In_1522,In_1818);
or U245 (N_245,In_167,In_1258);
and U246 (N_246,In_257,In_1984);
and U247 (N_247,In_118,In_1524);
nand U248 (N_248,In_1792,In_1580);
or U249 (N_249,In_913,In_372);
and U250 (N_250,In_1434,In_926);
or U251 (N_251,In_1948,In_836);
or U252 (N_252,In_1519,In_1430);
nand U253 (N_253,N_117,In_28);
or U254 (N_254,In_1287,In_898);
nor U255 (N_255,In_1191,N_96);
nor U256 (N_256,In_438,In_34);
nand U257 (N_257,N_140,In_1222);
and U258 (N_258,In_1145,In_1415);
nand U259 (N_259,In_1357,In_662);
nand U260 (N_260,In_1036,In_919);
nor U261 (N_261,N_190,In_159);
or U262 (N_262,In_1471,In_311);
or U263 (N_263,In_499,In_1691);
or U264 (N_264,In_1291,In_1444);
xor U265 (N_265,In_1117,N_63);
or U266 (N_266,In_948,N_149);
nand U267 (N_267,In_1800,In_307);
or U268 (N_268,In_1028,In_1378);
or U269 (N_269,In_1684,In_1006);
or U270 (N_270,In_303,In_1994);
and U271 (N_271,In_1319,In_1207);
and U272 (N_272,In_235,In_971);
nor U273 (N_273,N_118,N_45);
nor U274 (N_274,In_1050,N_243);
nand U275 (N_275,In_1309,In_965);
or U276 (N_276,In_994,In_1849);
nor U277 (N_277,In_467,In_705);
nand U278 (N_278,N_206,In_1391);
and U279 (N_279,In_1871,In_1971);
nor U280 (N_280,In_1985,In_1216);
and U281 (N_281,In_1908,In_886);
nand U282 (N_282,In_1982,In_1416);
nand U283 (N_283,In_1173,In_556);
xor U284 (N_284,N_27,In_1436);
nand U285 (N_285,In_80,In_1460);
nand U286 (N_286,In_860,In_1321);
nor U287 (N_287,In_475,In_1887);
nand U288 (N_288,N_39,In_1748);
nand U289 (N_289,In_1180,N_110);
nand U290 (N_290,In_156,In_493);
or U291 (N_291,In_294,In_743);
nand U292 (N_292,N_183,In_1233);
or U293 (N_293,In_570,In_181);
and U294 (N_294,N_26,In_1147);
or U295 (N_295,In_1497,In_1516);
and U296 (N_296,In_1140,In_406);
xnor U297 (N_297,In_1904,In_818);
xnor U298 (N_298,N_207,In_765);
or U299 (N_299,In_1165,N_56);
nor U300 (N_300,In_1546,In_171);
or U301 (N_301,In_254,In_897);
and U302 (N_302,In_576,In_574);
or U303 (N_303,In_1218,In_1328);
or U304 (N_304,In_431,In_1197);
and U305 (N_305,In_1023,In_1693);
and U306 (N_306,In_1387,N_22);
nor U307 (N_307,In_1727,In_1240);
or U308 (N_308,In_136,In_250);
or U309 (N_309,In_859,In_1733);
and U310 (N_310,In_1118,In_1186);
or U311 (N_311,In_1983,In_1010);
nand U312 (N_312,In_100,In_1105);
nor U313 (N_313,In_1313,In_1548);
and U314 (N_314,In_791,In_1368);
and U315 (N_315,In_148,In_245);
or U316 (N_316,In_827,In_326);
or U317 (N_317,In_1198,N_228);
or U318 (N_318,In_153,In_959);
nand U319 (N_319,In_690,In_23);
and U320 (N_320,In_20,In_626);
nor U321 (N_321,In_1981,In_702);
nand U322 (N_322,In_840,In_110);
nor U323 (N_323,N_3,In_328);
and U324 (N_324,In_747,In_160);
nand U325 (N_325,In_1664,In_1395);
xnor U326 (N_326,In_1577,In_1639);
or U327 (N_327,In_1411,In_1784);
nand U328 (N_328,In_1824,N_11);
nor U329 (N_329,In_901,In_829);
nor U330 (N_330,In_1174,In_1251);
and U331 (N_331,In_1476,In_881);
or U332 (N_332,In_12,In_931);
or U333 (N_333,In_1736,In_1531);
nor U334 (N_334,In_1958,In_1526);
nor U335 (N_335,In_1177,In_486);
nor U336 (N_336,In_1567,In_373);
nor U337 (N_337,In_239,In_116);
or U338 (N_338,In_1161,N_173);
xnor U339 (N_339,In_1351,N_220);
and U340 (N_340,In_1756,In_1341);
or U341 (N_341,In_444,N_236);
or U342 (N_342,In_24,In_1665);
or U343 (N_343,In_1474,In_1058);
nand U344 (N_344,In_1620,N_144);
and U345 (N_345,In_542,In_1295);
nor U346 (N_346,In_1362,N_104);
and U347 (N_347,In_1493,In_1628);
and U348 (N_348,N_88,N_92);
or U349 (N_349,In_408,In_1806);
xnor U350 (N_350,In_1517,In_1081);
nand U351 (N_351,N_204,In_876);
nand U352 (N_352,In_1941,In_801);
nor U353 (N_353,In_1296,In_929);
and U354 (N_354,In_1892,In_1412);
or U355 (N_355,In_1657,In_1463);
nor U356 (N_356,In_1154,N_152);
nand U357 (N_357,In_1615,N_178);
or U358 (N_358,In_4,In_508);
nor U359 (N_359,In_953,In_449);
xnor U360 (N_360,In_310,In_244);
and U361 (N_361,In_1821,In_109);
or U362 (N_362,N_121,In_297);
nor U363 (N_363,N_8,In_364);
and U364 (N_364,N_54,In_30);
nand U365 (N_365,In_64,In_1509);
and U366 (N_366,In_506,In_703);
and U367 (N_367,In_121,In_541);
nor U368 (N_368,In_356,In_941);
nor U369 (N_369,In_993,In_713);
nor U370 (N_370,In_618,In_1889);
or U371 (N_371,In_1934,In_192);
and U372 (N_372,N_66,In_661);
xor U373 (N_373,In_305,In_1001);
nor U374 (N_374,In_81,N_94);
and U375 (N_375,In_127,N_115);
or U376 (N_376,N_62,In_790);
or U377 (N_377,N_79,In_232);
nor U378 (N_378,In_101,N_87);
nor U379 (N_379,In_1414,N_86);
nand U380 (N_380,N_160,In_1518);
nand U381 (N_381,N_10,In_320);
or U382 (N_382,In_471,N_161);
or U383 (N_383,In_1888,In_1134);
xor U384 (N_384,N_0,In_396);
and U385 (N_385,In_667,N_237);
and U386 (N_386,N_131,In_1274);
or U387 (N_387,In_1584,In_1275);
nor U388 (N_388,In_857,In_1033);
and U389 (N_389,In_925,In_862);
and U390 (N_390,In_454,In_1864);
nor U391 (N_391,In_1687,In_884);
or U392 (N_392,N_145,In_419);
nand U393 (N_393,In_1891,In_715);
and U394 (N_394,In_956,In_1585);
nand U395 (N_395,In_365,In_1564);
and U396 (N_396,In_658,In_852);
or U397 (N_397,In_1804,In_595);
nand U398 (N_398,In_1830,In_621);
xor U399 (N_399,In_1525,In_1427);
nor U400 (N_400,In_1791,In_1819);
nor U401 (N_401,In_1290,In_492);
or U402 (N_402,In_494,In_1646);
nand U403 (N_403,In_821,In_1492);
nand U404 (N_404,N_102,In_665);
nor U405 (N_405,In_742,In_1969);
or U406 (N_406,In_711,In_1150);
xnor U407 (N_407,In_1721,In_1747);
nand U408 (N_408,In_1236,In_1409);
xnor U409 (N_409,In_624,In_437);
or U410 (N_410,In_726,In_385);
nand U411 (N_411,In_1100,In_921);
and U412 (N_412,In_1424,In_1230);
and U413 (N_413,In_1512,In_482);
and U414 (N_414,N_143,In_1650);
or U415 (N_415,In_1119,In_422);
or U416 (N_416,N_136,In_816);
or U417 (N_417,N_176,In_639);
or U418 (N_418,In_456,In_887);
or U419 (N_419,In_780,In_1712);
or U420 (N_420,In_73,In_1420);
nor U421 (N_421,In_461,In_1552);
or U422 (N_422,In_485,N_23);
nor U423 (N_423,In_1835,In_1044);
nand U424 (N_424,In_1418,In_1213);
nor U425 (N_425,In_1196,In_1679);
or U426 (N_426,In_1631,In_330);
nor U427 (N_427,N_189,N_21);
nand U428 (N_428,In_674,In_681);
nand U429 (N_429,In_1060,In_1634);
or U430 (N_430,In_1008,In_483);
nor U431 (N_431,In_784,In_1211);
xor U432 (N_432,In_1710,In_987);
nand U433 (N_433,In_1208,In_1480);
and U434 (N_434,In_608,In_1042);
nand U435 (N_435,N_109,In_1468);
nor U436 (N_436,In_764,In_944);
and U437 (N_437,N_212,In_1749);
nand U438 (N_438,In_1022,In_1903);
and U439 (N_439,In_172,In_1974);
or U440 (N_440,In_1886,In_1597);
nand U441 (N_441,In_1454,In_1939);
nand U442 (N_442,N_98,In_1361);
or U443 (N_443,In_638,N_97);
xor U444 (N_444,In_659,In_282);
nand U445 (N_445,In_1045,In_1965);
nand U446 (N_446,In_92,In_548);
nor U447 (N_447,In_947,In_1992);
nor U448 (N_448,In_55,In_1113);
nand U449 (N_449,In_480,In_1340);
and U450 (N_450,N_116,N_55);
nor U451 (N_451,In_1883,N_49);
nor U452 (N_452,In_1976,In_871);
and U453 (N_453,In_969,In_1440);
xor U454 (N_454,In_1744,In_267);
or U455 (N_455,In_150,In_1080);
nand U456 (N_456,In_1523,In_98);
or U457 (N_457,In_403,In_511);
nand U458 (N_458,In_585,In_188);
nor U459 (N_459,In_1016,In_1591);
and U460 (N_460,N_67,In_1009);
and U461 (N_461,In_1303,In_1774);
and U462 (N_462,N_181,In_644);
and U463 (N_463,In_393,N_169);
or U464 (N_464,In_1820,In_786);
nand U465 (N_465,In_916,In_960);
or U466 (N_466,In_1408,In_455);
nand U467 (N_467,In_173,N_226);
and U468 (N_468,N_241,In_600);
nand U469 (N_469,N_155,In_962);
and U470 (N_470,In_1088,In_688);
xor U471 (N_471,In_1561,In_900);
nor U472 (N_472,In_1990,In_1061);
nand U473 (N_473,In_709,In_1645);
xnor U474 (N_474,In_1210,In_120);
and U475 (N_475,In_717,In_293);
nand U476 (N_476,In_1759,In_349);
nand U477 (N_477,In_276,In_1837);
xor U478 (N_478,In_0,In_1632);
xor U479 (N_479,In_1812,In_1709);
xor U480 (N_480,In_700,In_1702);
xor U481 (N_481,In_347,In_1334);
and U482 (N_482,In_566,N_245);
and U483 (N_483,In_1429,In_1694);
or U484 (N_484,In_139,In_327);
or U485 (N_485,In_1280,In_1263);
and U486 (N_486,In_1698,N_168);
xor U487 (N_487,In_1576,In_1825);
xor U488 (N_488,N_47,N_157);
nor U489 (N_489,In_1076,In_545);
or U490 (N_490,In_228,In_1957);
or U491 (N_491,In_805,In_360);
xnor U492 (N_492,In_622,N_127);
xnor U493 (N_493,N_230,N_34);
and U494 (N_494,In_266,In_974);
nand U495 (N_495,In_970,In_218);
and U496 (N_496,In_134,In_9);
nand U497 (N_497,In_609,N_195);
nor U498 (N_498,In_704,In_1120);
nand U499 (N_499,In_927,In_387);
or U500 (N_500,In_201,In_104);
or U501 (N_501,In_641,In_1039);
or U502 (N_502,In_1532,In_1026);
nor U503 (N_503,In_11,In_1929);
or U504 (N_504,In_1157,In_240);
nand U505 (N_505,In_613,N_358);
and U506 (N_506,In_554,In_750);
and U507 (N_507,N_467,N_38);
and U508 (N_508,In_855,N_210);
nand U509 (N_509,In_1543,In_1126);
nand U510 (N_510,N_421,In_184);
or U511 (N_511,N_232,In_446);
or U512 (N_512,In_1360,N_71);
and U513 (N_513,In_689,In_629);
and U514 (N_514,In_164,N_163);
xor U515 (N_515,N_400,N_423);
or U516 (N_516,In_391,In_1272);
nand U517 (N_517,In_147,N_36);
or U518 (N_518,In_1536,In_1030);
or U519 (N_519,N_307,N_130);
and U520 (N_520,In_946,N_167);
or U521 (N_521,In_335,In_1014);
nor U522 (N_522,In_348,In_350);
nor U523 (N_523,In_1753,N_355);
or U524 (N_524,In_1437,In_1171);
and U525 (N_525,In_1123,In_1973);
nand U526 (N_526,N_6,In_117);
xnor U527 (N_527,N_246,N_303);
or U528 (N_528,N_327,In_889);
or U529 (N_529,N_271,In_93);
nand U530 (N_530,In_1246,N_128);
nand U531 (N_531,In_3,In_1032);
nand U532 (N_532,N_330,In_1002);
and U533 (N_533,In_1181,In_543);
nand U534 (N_534,In_573,In_1343);
and U535 (N_535,In_1470,In_501);
and U536 (N_536,In_1967,In_90);
nor U537 (N_537,In_292,In_1955);
nand U538 (N_538,In_82,In_627);
and U539 (N_539,In_883,In_1394);
nor U540 (N_540,N_337,In_291);
nand U541 (N_541,In_377,In_647);
nor U542 (N_542,N_171,N_219);
nand U543 (N_543,In_199,In_1215);
nor U544 (N_544,In_512,In_399);
or U545 (N_545,N_377,In_1807);
xnor U546 (N_546,In_918,In_1481);
and U547 (N_547,In_518,In_33);
nand U548 (N_548,In_1299,In_137);
nor U549 (N_549,N_250,N_446);
and U550 (N_550,In_263,In_31);
nand U551 (N_551,In_899,In_1371);
nand U552 (N_552,In_450,In_572);
or U553 (N_553,N_286,In_663);
and U554 (N_554,N_216,In_1229);
and U555 (N_555,In_873,In_108);
xnor U556 (N_556,In_329,In_260);
xnor U557 (N_557,In_1164,In_1666);
and U558 (N_558,In_510,In_1782);
nand U559 (N_559,In_551,N_33);
or U560 (N_560,N_148,N_396);
nor U561 (N_561,In_243,In_757);
or U562 (N_562,In_1428,In_1271);
nor U563 (N_563,In_1760,N_442);
nand U564 (N_564,In_27,N_135);
or U565 (N_565,In_1928,In_1605);
nor U566 (N_566,N_52,N_69);
or U567 (N_567,In_771,N_479);
xnor U568 (N_568,In_1874,N_319);
or U569 (N_569,N_420,N_499);
or U570 (N_570,N_388,In_975);
and U571 (N_571,N_64,In_1838);
nand U572 (N_572,In_1135,In_22);
and U573 (N_573,In_1950,In_1269);
and U574 (N_574,In_124,In_737);
or U575 (N_575,In_1858,In_107);
nand U576 (N_576,In_1877,In_1363);
or U577 (N_577,In_58,In_672);
nor U578 (N_578,In_1376,N_434);
or U579 (N_579,In_1005,In_680);
and U580 (N_580,In_313,N_222);
nand U581 (N_581,N_199,In_1681);
or U582 (N_582,In_1209,N_424);
or U583 (N_583,In_1617,In_1624);
nor U584 (N_584,In_1326,N_114);
and U585 (N_585,In_978,N_346);
or U586 (N_586,In_1336,N_187);
and U587 (N_587,In_1446,N_248);
or U588 (N_588,N_493,N_441);
nor U589 (N_589,In_339,In_1450);
nor U590 (N_590,In_1731,N_12);
nor U591 (N_591,N_277,In_353);
nor U592 (N_592,In_1185,In_1930);
or U593 (N_593,In_465,In_445);
and U594 (N_594,N_380,N_122);
or U595 (N_595,In_670,N_449);
nand U596 (N_596,N_411,In_846);
nor U597 (N_597,In_448,In_280);
nor U598 (N_598,In_1775,In_1547);
nand U599 (N_599,In_26,In_1018);
xor U600 (N_600,In_666,In_1183);
nand U601 (N_601,In_416,N_14);
and U602 (N_602,In_1927,In_1542);
and U603 (N_603,In_930,In_1999);
xor U604 (N_604,In_684,In_230);
or U605 (N_605,In_1302,In_1426);
and U606 (N_606,In_378,In_1653);
xor U607 (N_607,In_559,N_74);
nand U608 (N_608,N_105,In_806);
or U609 (N_609,In_500,In_6);
nand U610 (N_610,In_370,N_208);
nand U611 (N_611,N_414,In_319);
nor U612 (N_612,In_1647,N_344);
nand U613 (N_613,N_452,In_1865);
or U614 (N_614,In_1642,In_65);
xor U615 (N_615,In_88,In_1338);
and U616 (N_616,In_1936,In_1380);
and U617 (N_617,N_90,In_563);
nor U618 (N_618,In_1911,In_1324);
xnor U619 (N_619,N_99,In_650);
or U620 (N_620,In_1294,In_823);
nor U621 (N_621,In_1329,N_78);
or U622 (N_622,N_153,N_399);
nand U623 (N_623,In_424,In_1785);
nor U624 (N_624,N_188,In_1574);
nand U625 (N_625,In_15,In_1828);
or U626 (N_626,In_1015,In_720);
and U627 (N_627,N_261,In_1890);
nand U628 (N_628,In_256,In_1069);
and U629 (N_629,In_1084,In_850);
nor U630 (N_630,In_1099,In_1332);
nor U631 (N_631,In_1978,In_97);
and U632 (N_632,In_502,N_431);
or U633 (N_633,In_1163,N_274);
or U634 (N_634,In_298,In_1619);
nor U635 (N_635,In_803,In_1913);
xor U636 (N_636,In_1811,In_1757);
and U637 (N_637,N_427,In_922);
nand U638 (N_638,In_1764,In_407);
and U639 (N_639,N_42,In_169);
xor U640 (N_640,N_375,In_1350);
nor U641 (N_641,N_360,In_549);
xor U642 (N_642,In_76,N_459);
nor U643 (N_643,N_356,N_287);
nor U644 (N_644,In_1188,In_1690);
nand U645 (N_645,In_1487,N_306);
and U646 (N_646,N_439,In_1590);
or U647 (N_647,In_945,In_936);
nor U648 (N_648,N_300,In_1839);
and U649 (N_649,In_848,In_1832);
or U650 (N_650,N_325,N_259);
nor U651 (N_651,N_72,In_568);
and U652 (N_652,In_1918,In_1729);
and U653 (N_653,In_1356,In_792);
nand U654 (N_654,In_864,In_1856);
nor U655 (N_655,In_1179,In_1383);
nor U656 (N_656,In_552,N_132);
nor U657 (N_657,In_783,In_1529);
and U658 (N_658,In_1040,N_59);
nand U659 (N_659,In_362,In_1219);
nor U660 (N_660,In_415,In_128);
or U661 (N_661,In_1201,In_706);
or U662 (N_662,In_1707,In_322);
nand U663 (N_663,In_1104,In_1110);
and U664 (N_664,N_395,In_891);
nor U665 (N_665,N_343,In_1255);
or U666 (N_666,N_269,N_80);
xnor U667 (N_667,In_957,In_979);
nand U668 (N_668,In_1310,In_851);
nor U669 (N_669,N_235,In_1711);
and U670 (N_670,In_834,In_1551);
or U671 (N_671,In_288,In_77);
or U672 (N_672,N_276,In_1352);
nor U673 (N_673,In_1779,In_1751);
or U674 (N_674,In_598,In_1490);
nand U675 (N_675,In_1285,N_448);
xor U676 (N_676,In_1638,In_597);
nand U677 (N_677,In_50,In_825);
and U678 (N_678,In_1772,In_1115);
nand U679 (N_679,In_1786,N_315);
nand U680 (N_680,In_1951,In_1926);
and U681 (N_681,N_326,In_54);
nand U682 (N_682,In_166,In_1459);
nand U683 (N_683,In_434,In_53);
or U684 (N_684,N_314,N_106);
and U685 (N_685,In_521,In_1797);
nand U686 (N_686,In_36,In_697);
and U687 (N_687,In_487,In_165);
nand U688 (N_688,In_1393,N_416);
nor U689 (N_689,N_46,In_234);
nor U690 (N_690,In_1075,In_1469);
xnor U691 (N_691,In_211,N_378);
nand U692 (N_692,N_29,In_163);
or U693 (N_693,In_675,In_1074);
or U694 (N_694,In_1046,In_145);
nor U695 (N_695,In_515,In_1413);
nand U696 (N_696,In_890,In_721);
and U697 (N_697,In_258,N_363);
xnor U698 (N_698,In_1558,In_1861);
xnor U699 (N_699,In_404,N_367);
nor U700 (N_700,In_1538,In_560);
or U701 (N_701,N_83,In_782);
nand U702 (N_702,N_223,In_1625);
and U703 (N_703,N_304,N_408);
nand U704 (N_704,In_1677,In_1922);
nor U705 (N_705,In_1925,In_1149);
nand U706 (N_706,N_445,In_776);
nand U707 (N_707,In_1443,In_1478);
nor U708 (N_708,N_422,In_968);
or U709 (N_709,N_255,In_1783);
and U710 (N_710,N_9,In_382);
nand U711 (N_711,In_1262,N_382);
nor U712 (N_712,N_495,In_229);
and U713 (N_713,In_1268,In_835);
and U714 (N_714,In_144,In_1325);
xnor U715 (N_715,N_266,In_1038);
nor U716 (N_716,N_194,N_256);
nor U717 (N_717,In_813,In_45);
nand U718 (N_718,In_1944,In_571);
or U719 (N_719,In_72,N_438);
nand U720 (N_720,In_847,In_812);
xnor U721 (N_721,In_761,In_430);
nand U722 (N_722,In_1734,In_47);
nor U723 (N_723,In_1794,N_25);
nand U724 (N_724,N_457,N_345);
xor U725 (N_725,In_1968,In_1946);
nor U726 (N_726,In_212,In_995);
or U727 (N_727,In_1063,In_1575);
xor U728 (N_728,In_648,In_934);
and U729 (N_729,In_687,In_996);
or U730 (N_730,In_869,In_1924);
nor U731 (N_731,In_289,N_218);
or U732 (N_732,In_985,In_777);
or U733 (N_733,N_81,In_1935);
nor U734 (N_734,In_468,In_226);
nor U735 (N_735,In_991,N_231);
nand U736 (N_736,N_381,In_1884);
nand U737 (N_737,N_125,In_1204);
and U738 (N_738,In_1544,N_417);
nor U739 (N_739,N_24,In_187);
and U740 (N_740,N_316,In_1304);
or U741 (N_741,In_1599,In_811);
nand U742 (N_742,In_1521,In_290);
nor U743 (N_743,In_1715,In_283);
or U744 (N_744,N_247,In_950);
nand U745 (N_745,In_119,N_1);
xor U746 (N_746,N_175,In_1662);
nor U747 (N_747,In_1212,In_1815);
and U748 (N_748,In_1,N_494);
or U749 (N_749,In_1064,In_221);
and U750 (N_750,N_321,In_1822);
xnor U751 (N_751,In_1809,In_1550);
and U752 (N_752,N_119,In_428);
xnor U753 (N_753,N_588,N_469);
nand U754 (N_754,In_695,N_682);
or U755 (N_755,In_839,In_617);
nand U756 (N_756,N_518,In_1945);
and U757 (N_757,N_450,N_557);
and U758 (N_758,N_564,In_1056);
and U759 (N_759,In_1505,In_146);
and U760 (N_760,N_713,N_293);
and U761 (N_761,N_526,N_348);
or U762 (N_762,N_488,N_731);
nor U763 (N_763,In_964,In_43);
nor U764 (N_764,In_1148,In_1252);
nand U765 (N_765,In_478,In_854);
xnor U766 (N_766,N_500,N_260);
nand U767 (N_767,In_1244,N_569);
nor U768 (N_768,In_1195,N_656);
or U769 (N_769,In_247,N_44);
and U770 (N_770,N_224,N_107);
and U771 (N_771,In_710,N_100);
nand U772 (N_772,N_695,N_308);
and U773 (N_773,In_345,N_697);
or U774 (N_774,In_804,N_402);
and U775 (N_775,N_565,In_1475);
nand U776 (N_776,N_252,In_939);
nand U777 (N_777,In_1359,In_130);
or U778 (N_778,N_392,N_586);
and U779 (N_779,In_1902,N_470);
xnor U780 (N_780,In_1769,In_745);
nor U781 (N_781,In_271,In_476);
and U782 (N_782,N_738,N_141);
or U783 (N_783,In_1609,N_95);
nor U784 (N_784,N_607,In_8);
nor U785 (N_785,N_735,N_65);
nor U786 (N_786,In_912,N_462);
nor U787 (N_787,In_587,In_1563);
and U788 (N_788,N_700,In_749);
and U789 (N_789,N_619,In_414);
and U790 (N_790,In_1689,In_1226);
and U791 (N_791,N_587,In_1250);
and U792 (N_792,N_368,In_798);
nor U793 (N_793,In_1954,In_1349);
or U794 (N_794,N_727,In_1594);
and U795 (N_795,In_1613,N_523);
nor U796 (N_796,In_1479,In_346);
or U797 (N_797,N_322,In_1388);
nor U798 (N_798,N_318,In_398);
nor U799 (N_799,N_599,N_542);
nand U800 (N_800,N_585,In_1754);
or U801 (N_801,N_671,N_721);
nand U802 (N_802,N_298,In_849);
nor U803 (N_803,In_462,N_180);
nor U804 (N_804,In_623,N_548);
nor U805 (N_805,N_340,N_609);
nor U806 (N_806,In_517,N_649);
xnor U807 (N_807,N_133,N_387);
or U808 (N_808,In_405,N_379);
and U809 (N_809,N_112,N_606);
and U810 (N_810,N_748,N_556);
or U811 (N_811,N_366,In_1007);
or U812 (N_812,In_86,N_407);
or U813 (N_813,N_20,N_629);
nor U814 (N_814,In_1726,N_323);
nand U815 (N_815,In_440,In_1224);
nor U816 (N_816,In_1448,In_1592);
nor U817 (N_817,N_635,In_1964);
and U818 (N_818,In_1636,N_594);
or U819 (N_819,N_405,In_1472);
nand U820 (N_820,In_1725,In_1676);
or U821 (N_821,In_762,In_1700);
xnor U822 (N_822,In_550,In_1813);
and U823 (N_823,In_224,In_843);
and U824 (N_824,In_1655,In_312);
or U825 (N_825,N_507,In_800);
or U826 (N_826,In_1696,N_460);
nand U827 (N_827,In_616,In_1768);
or U828 (N_828,In_928,In_712);
or U829 (N_829,In_123,N_528);
xor U830 (N_830,In_630,In_89);
nor U831 (N_831,In_775,In_972);
nand U832 (N_832,N_61,In_673);
nand U833 (N_833,In_1510,In_1400);
nor U834 (N_834,N_156,In_222);
xnor U835 (N_835,In_68,In_279);
nand U836 (N_836,N_544,In_1669);
or U837 (N_837,In_361,N_113);
nand U838 (N_838,In_1166,In_1189);
or U839 (N_839,N_383,N_262);
nor U840 (N_840,N_618,In_1386);
and U841 (N_841,In_436,In_820);
and U842 (N_842,In_400,In_719);
or U843 (N_843,N_174,N_679);
and U844 (N_844,N_626,In_1581);
nand U845 (N_845,N_570,In_1504);
or U846 (N_846,In_819,N_15);
nand U847 (N_847,In_1139,In_1909);
nand U848 (N_848,In_1881,In_1724);
nor U849 (N_849,In_1621,In_676);
nand U850 (N_850,N_257,In_447);
nor U851 (N_851,In_1614,In_1893);
nand U852 (N_852,In_1237,N_709);
nor U853 (N_853,In_459,N_657);
nand U854 (N_854,In_817,N_623);
or U855 (N_855,In_390,N_684);
and U856 (N_856,N_693,N_253);
nor U857 (N_857,N_455,N_593);
nand U858 (N_858,In_470,In_285);
nand U859 (N_859,In_1947,In_1298);
or U860 (N_860,In_204,In_781);
nor U861 (N_861,N_279,In_770);
xor U862 (N_862,In_161,In_1242);
nor U863 (N_863,In_1553,N_481);
or U864 (N_864,N_554,N_35);
nand U865 (N_865,In_1987,In_1317);
or U866 (N_866,N_608,In_1431);
or U867 (N_867,N_221,In_1537);
or U868 (N_868,In_1952,In_1398);
nor U869 (N_869,In_300,In_718);
nand U870 (N_870,In_1916,N_370);
xnor U871 (N_871,N_409,In_175);
nor U872 (N_872,In_42,N_737);
nor U873 (N_873,N_497,In_532);
nor U874 (N_874,N_553,In_1765);
xnor U875 (N_875,N_349,In_1962);
nand U876 (N_876,N_461,N_137);
xor U877 (N_877,In_907,N_389);
nor U878 (N_878,In_882,In_40);
nor U879 (N_879,In_252,N_390);
nand U880 (N_880,In_1231,In_1616);
and U881 (N_881,N_611,N_82);
or U882 (N_882,In_363,N_234);
nor U883 (N_883,N_7,N_444);
nand U884 (N_884,N_524,N_664);
nor U885 (N_885,In_1260,In_1306);
or U886 (N_886,In_472,In_1392);
nand U887 (N_887,In_140,In_1572);
nand U888 (N_888,In_1802,In_668);
or U889 (N_889,In_628,In_112);
nand U890 (N_890,In_1789,In_1961);
or U891 (N_891,N_333,In_1589);
or U892 (N_892,N_458,In_1656);
nor U893 (N_893,N_205,In_1738);
and U894 (N_894,In_911,N_749);
or U895 (N_895,In_863,N_701);
or U896 (N_896,In_1688,N_336);
and U897 (N_897,N_668,In_420);
or U898 (N_898,In_558,In_1144);
nor U899 (N_899,N_703,In_1637);
nor U900 (N_900,N_690,N_386);
xor U901 (N_901,In_1674,In_1142);
nor U902 (N_902,In_1034,In_1066);
and U903 (N_903,In_60,In_1214);
nor U904 (N_904,In_614,In_1986);
nand U905 (N_905,In_1501,N_515);
or U906 (N_906,N_294,N_48);
nand U907 (N_907,In_1627,In_1342);
nor U908 (N_908,In_537,In_620);
xor U909 (N_909,In_1200,N_331);
xnor U910 (N_910,N_284,N_320);
and U911 (N_911,N_589,In_497);
and U912 (N_912,In_1556,N_715);
nand U913 (N_913,N_443,In_973);
nor U914 (N_914,N_642,N_590);
or U915 (N_915,N_698,In_48);
and U916 (N_916,N_734,N_562);
xnor U917 (N_917,N_631,In_555);
nand U918 (N_918,In_1053,In_1899);
nand U919 (N_919,In_529,N_743);
nand U920 (N_920,N_705,In_1107);
and U921 (N_921,In_332,In_619);
xnor U922 (N_922,In_180,N_617);
or U923 (N_923,N_616,In_1203);
nand U924 (N_924,In_1746,In_1989);
and U925 (N_925,In_268,N_512);
nand U926 (N_926,N_487,N_288);
or U927 (N_927,N_475,N_673);
nor U928 (N_928,N_742,N_372);
and U929 (N_929,In_1777,N_60);
nand U930 (N_930,In_822,In_1245);
xnor U931 (N_931,In_198,N_91);
xnor U932 (N_932,N_678,In_432);
nor U933 (N_933,N_89,N_275);
nand U934 (N_934,N_254,In_1381);
nand U935 (N_935,N_660,In_1087);
nand U936 (N_936,N_520,In_1579);
or U937 (N_937,N_747,N_621);
nand U938 (N_938,In_1851,N_572);
or U939 (N_939,N_650,N_413);
xor U940 (N_940,In_1993,In_1697);
nor U941 (N_941,In_79,N_600);
and U942 (N_942,In_920,N_415);
nand U943 (N_943,In_1788,In_1397);
or U944 (N_944,In_1852,N_490);
xnor U945 (N_945,In_1399,N_70);
or U946 (N_946,In_1384,In_1146);
or U947 (N_947,In_738,N_696);
xnor U948 (N_948,N_555,In_1466);
and U949 (N_949,In_635,In_1159);
nor U950 (N_950,N_614,In_417);
nor U951 (N_951,In_539,N_484);
and U952 (N_952,N_93,N_648);
nand U953 (N_953,In_1124,N_301);
nor U954 (N_954,In_1182,In_1652);
nand U955 (N_955,In_392,N_401);
or U956 (N_956,N_634,In_1569);
or U957 (N_957,In_1868,In_1798);
and U958 (N_958,In_1495,N_683);
nor U959 (N_959,In_49,In_302);
nand U960 (N_960,N_311,In_488);
nor U961 (N_961,In_513,N_640);
or U962 (N_962,N_329,In_186);
and U963 (N_963,N_440,In_375);
or U964 (N_964,In_355,In_1741);
and U965 (N_965,In_1017,In_102);
and U966 (N_966,In_1348,N_312);
nor U967 (N_967,In_1101,N_525);
and U968 (N_968,N_313,In_498);
or U969 (N_969,In_751,In_325);
nand U970 (N_970,N_165,N_547);
nor U971 (N_971,In_1355,In_531);
nand U972 (N_972,N_559,N_632);
or U973 (N_973,In_394,N_177);
and U974 (N_974,In_569,In_44);
or U975 (N_975,In_1870,N_214);
nor U976 (N_976,In_1421,In_219);
nor U977 (N_977,In_779,In_1578);
nor U978 (N_978,In_324,In_426);
or U979 (N_979,N_101,N_108);
or U980 (N_980,In_727,N_332);
xor U981 (N_981,N_432,In_106);
nand U982 (N_982,In_540,N_192);
and U983 (N_983,In_1743,In_246);
or U984 (N_984,In_877,N_672);
nand U985 (N_985,In_1228,N_674);
nor U986 (N_986,N_483,N_17);
xnor U987 (N_987,N_258,In_553);
or U988 (N_988,In_1307,N_265);
nor U989 (N_989,N_397,In_1453);
and U990 (N_990,In_195,N_273);
and U991 (N_991,In_1441,In_833);
nand U992 (N_992,N_489,In_1503);
xnor U993 (N_993,In_610,N_209);
nand U994 (N_994,In_509,In_940);
and U995 (N_995,In_604,N_530);
nor U996 (N_996,N_32,N_706);
nor U997 (N_997,In_1491,N_40);
nand U998 (N_998,N_339,N_394);
and U999 (N_999,N_663,In_1956);
and U1000 (N_1000,In_309,N_211);
or U1001 (N_1001,In_1327,N_347);
and U1002 (N_1002,N_198,N_850);
nand U1003 (N_1003,N_999,N_964);
and U1004 (N_1004,N_848,N_579);
nor U1005 (N_1005,In_1047,N_295);
nand U1006 (N_1006,N_838,In_958);
and U1007 (N_1007,In_643,N_932);
xor U1008 (N_1008,N_763,In_193);
and U1009 (N_1009,N_688,N_376);
nor U1010 (N_1010,In_1021,N_430);
and U1011 (N_1011,In_39,In_227);
xnor U1012 (N_1012,N_73,N_426);
nor U1013 (N_1013,In_1172,N_956);
xor U1014 (N_1014,N_857,N_781);
xor U1015 (N_1015,In_114,In_1025);
or U1016 (N_1016,N_43,N_662);
nand U1017 (N_1017,N_945,N_900);
xnor U1018 (N_1018,N_861,In_190);
nand U1019 (N_1019,N_784,In_1217);
nor U1020 (N_1020,In_1623,N_710);
or U1021 (N_1021,N_844,N_724);
nor U1022 (N_1022,N_711,N_787);
or U1023 (N_1023,In_942,N_971);
xnor U1024 (N_1024,N_403,In_868);
xor U1025 (N_1025,N_474,In_1966);
nor U1026 (N_1026,N_806,N_595);
and U1027 (N_1027,N_874,N_369);
and U1028 (N_1028,N_558,N_815);
or U1029 (N_1029,N_604,N_539);
nand U1030 (N_1030,N_645,In_85);
nand U1031 (N_1031,In_1051,N_921);
and U1032 (N_1032,N_753,In_1937);
nor U1033 (N_1033,In_893,N_215);
nand U1034 (N_1034,In_651,N_227);
and U1035 (N_1035,N_371,N_305);
nor U1036 (N_1036,N_940,In_1072);
nor U1037 (N_1037,In_910,In_395);
nor U1038 (N_1038,N_571,N_504);
nor U1039 (N_1039,N_817,In_1867);
or U1040 (N_1040,N_702,N_856);
nand U1041 (N_1041,N_661,N_761);
nor U1042 (N_1042,N_916,In_1106);
or U1043 (N_1043,In_185,N_30);
nand U1044 (N_1044,N_755,In_1089);
and U1045 (N_1045,N_406,N_685);
and U1046 (N_1046,N_882,In_530);
nand U1047 (N_1047,In_1660,N_2);
nor U1048 (N_1048,In_1442,In_593);
nand U1049 (N_1049,N_597,N_637);
xnor U1050 (N_1050,In_1289,N_926);
nor U1051 (N_1051,N_53,In_1761);
and U1052 (N_1052,N_890,N_691);
or U1053 (N_1053,N_436,N_918);
xor U1054 (N_1054,N_624,In_642);
and U1055 (N_1055,N_816,N_404);
nor U1056 (N_1056,N_796,N_789);
nand U1057 (N_1057,N_847,N_859);
nor U1058 (N_1058,N_774,In_1790);
nor U1059 (N_1059,In_62,N_986);
nand U1060 (N_1060,N_839,N_982);
or U1061 (N_1061,In_990,In_1793);
or U1062 (N_1062,In_75,N_855);
nand U1063 (N_1063,N_268,In_1283);
and U1064 (N_1064,N_726,In_1855);
nand U1065 (N_1065,In_1845,N_270);
or U1066 (N_1066,N_788,N_584);
or U1067 (N_1067,In_795,In_441);
nand U1068 (N_1068,In_1375,In_70);
or U1069 (N_1069,N_798,In_1435);
nand U1070 (N_1070,In_1943,N_159);
or U1071 (N_1071,In_411,N_983);
xor U1072 (N_1072,In_1447,In_1176);
or U1073 (N_1073,In_435,N_994);
nand U1074 (N_1074,N_574,In_1000);
nand U1075 (N_1075,In_1776,N_85);
nor U1076 (N_1076,N_988,N_927);
nor U1077 (N_1077,N_84,In_284);
or U1078 (N_1078,In_413,N_767);
and U1079 (N_1079,N_545,In_1658);
or U1080 (N_1080,In_1312,In_507);
nand U1081 (N_1081,N_677,N_264);
or U1082 (N_1082,In_223,In_789);
nor U1083 (N_1083,In_1833,N_773);
nor U1084 (N_1084,N_338,N_797);
xnor U1085 (N_1085,N_953,N_533);
nand U1086 (N_1086,N_906,In_909);
xor U1087 (N_1087,In_1750,N_393);
and U1088 (N_1088,N_516,N_233);
or U1089 (N_1089,N_915,In_1808);
xnor U1090 (N_1090,N_299,In_105);
or U1091 (N_1091,N_581,In_1629);
and U1092 (N_1092,N_884,N_919);
nor U1093 (N_1093,N_760,In_1004);
xnor U1094 (N_1094,N_799,N_675);
and U1095 (N_1095,N_473,N_454);
nor U1096 (N_1096,In_754,N_733);
and U1097 (N_1097,N_123,N_653);
and U1098 (N_1098,In_1498,N_745);
nand U1099 (N_1099,N_566,In_1763);
or U1100 (N_1100,In_575,In_1178);
xor U1101 (N_1101,N_943,In_954);
or U1102 (N_1102,In_1345,N_361);
nor U1103 (N_1103,N_759,N_667);
or U1104 (N_1104,N_827,In_1857);
nand U1105 (N_1105,N_795,In_1128);
and U1106 (N_1106,In_1539,In_1912);
xnor U1107 (N_1107,In_56,In_1540);
nand U1108 (N_1108,In_1876,N_730);
or U1109 (N_1109,In_103,In_1405);
xor U1110 (N_1110,In_5,N_802);
nor U1111 (N_1111,N_151,N_942);
nor U1112 (N_1112,In_989,N_843);
or U1113 (N_1113,N_692,N_923);
nor U1114 (N_1114,N_418,N_717);
nor U1115 (N_1115,N_578,N_567);
and U1116 (N_1116,N_238,N_831);
xor U1117 (N_1117,N_292,In_1959);
and U1118 (N_1118,N_804,In_215);
or U1119 (N_1119,N_689,In_714);
and U1120 (N_1120,In_691,N_996);
and U1121 (N_1121,N_842,In_210);
nand U1122 (N_1122,N_981,N_718);
and U1123 (N_1123,N_891,N_908);
and U1124 (N_1124,N_948,N_828);
and U1125 (N_1125,In_99,N_466);
xnor U1126 (N_1126,N_998,N_636);
and U1127 (N_1127,In_384,N_782);
and U1128 (N_1128,In_1425,N_950);
or U1129 (N_1129,In_961,N_858);
or U1130 (N_1130,In_949,In_269);
nand U1131 (N_1131,N_851,In_1372);
nor U1132 (N_1132,N_465,In_1933);
and U1133 (N_1133,N_757,In_336);
or U1134 (N_1134,In_646,In_525);
or U1135 (N_1135,N_471,In_1878);
nor U1136 (N_1136,In_1037,N_193);
nand U1137 (N_1137,In_581,In_1608);
nor U1138 (N_1138,In_1464,N_139);
and U1139 (N_1139,N_750,N_510);
xnor U1140 (N_1140,N_546,In_591);
or U1141 (N_1141,In_334,N_979);
nor U1142 (N_1142,In_1603,N_583);
nor U1143 (N_1143,N_728,In_725);
nand U1144 (N_1144,In_157,In_1496);
or U1145 (N_1145,N_888,In_380);
xor U1146 (N_1146,In_91,N_324);
and U1147 (N_1147,N_203,N_941);
or U1148 (N_1148,N_962,In_1678);
or U1149 (N_1149,N_768,In_141);
and U1150 (N_1150,In_546,In_615);
and U1151 (N_1151,In_1885,In_1011);
xor U1152 (N_1152,In_1239,N_704);
or U1153 (N_1153,In_1520,In_1996);
and U1154 (N_1154,In_837,In_255);
nor U1155 (N_1155,In_1410,N_522);
and U1156 (N_1156,In_233,In_96);
and U1157 (N_1157,N_560,N_937);
or U1158 (N_1158,N_892,In_1029);
and U1159 (N_1159,In_1141,In_1673);
nand U1160 (N_1160,N_852,In_802);
nand U1161 (N_1161,N_754,N_317);
nand U1162 (N_1162,N_707,In_567);
nor U1163 (N_1163,N_786,N_876);
or U1164 (N_1164,In_888,N_561);
xor U1165 (N_1165,In_274,N_714);
nand U1166 (N_1166,N_641,In_878);
nor U1167 (N_1167,N_687,In_1742);
and U1168 (N_1168,N_741,In_1667);
nor U1169 (N_1169,In_683,In_374);
or U1170 (N_1170,N_643,In_796);
nor U1171 (N_1171,In_25,N_766);
and U1172 (N_1172,In_1292,N_756);
or U1173 (N_1173,N_746,In_1571);
or U1174 (N_1174,In_1301,N_719);
nand U1175 (N_1175,In_1205,N_901);
or U1176 (N_1176,In_562,In_976);
or U1177 (N_1177,In_526,N_76);
nand U1178 (N_1178,In_885,N_509);
or U1179 (N_1179,In_1705,In_1803);
or U1180 (N_1180,In_1847,N_162);
nand U1181 (N_1181,N_803,In_1719);
xnor U1182 (N_1182,N_535,In_645);
nand U1183 (N_1183,In_178,In_1339);
nand U1184 (N_1184,In_1716,N_818);
or U1185 (N_1185,In_514,N_592);
nor U1186 (N_1186,N_723,N_335);
and U1187 (N_1187,N_666,N_503);
or U1188 (N_1188,In_1184,N_834);
or U1189 (N_1189,N_809,N_811);
or U1190 (N_1190,N_771,N_960);
or U1191 (N_1191,N_917,In_1663);
or U1192 (N_1192,In_1787,N_867);
nor U1193 (N_1193,N_77,In_1722);
and U1194 (N_1194,In_479,N_521);
xor U1195 (N_1195,In_599,N_980);
nand U1196 (N_1196,In_1127,In_1862);
nand U1197 (N_1197,In_1586,In_774);
nor U1198 (N_1198,N_612,In_63);
nand U1199 (N_1199,In_287,In_1622);
xnor U1200 (N_1200,In_425,N_935);
and U1201 (N_1201,N_751,N_453);
nand U1202 (N_1202,N_527,In_671);
and U1203 (N_1203,In_861,In_1767);
nand U1204 (N_1204,N_37,N_716);
nand U1205 (N_1205,N_832,N_615);
or U1206 (N_1206,N_914,In_908);
or U1207 (N_1207,In_1109,N_739);
or U1208 (N_1208,In_685,N_922);
or U1209 (N_1209,N_138,N_909);
or U1210 (N_1210,N_961,N_573);
nor U1211 (N_1211,In_1612,In_1866);
nand U1212 (N_1212,In_1323,In_1094);
nand U1213 (N_1213,In_696,In_1369);
nand U1214 (N_1214,In_505,In_728);
or U1215 (N_1215,N_712,N_374);
and U1216 (N_1216,N_824,In_1227);
nand U1217 (N_1217,In_451,N_854);
nor U1218 (N_1218,N_837,N_875);
nand U1219 (N_1219,In_1685,In_1297);
nor U1220 (N_1220,N_864,N_870);
nand U1221 (N_1221,In_59,N_353);
nand U1222 (N_1222,N_352,In_533);
nor U1223 (N_1223,In_980,N_164);
and U1224 (N_1224,N_18,In_740);
nor U1225 (N_1225,N_647,In_1311);
nand U1226 (N_1226,N_866,In_769);
and U1227 (N_1227,N_708,N_536);
and U1228 (N_1228,N_877,N_873);
nand U1229 (N_1229,N_938,N_291);
nand U1230 (N_1230,N_896,N_830);
nor U1231 (N_1231,N_244,In_1920);
and U1232 (N_1232,N_758,N_947);
and U1233 (N_1233,In_1850,N_965);
xnor U1234 (N_1234,N_147,N_862);
or U1235 (N_1235,In_1499,N_776);
nor U1236 (N_1236,In_84,N_865);
and U1237 (N_1237,In_21,N_872);
and U1238 (N_1238,In_217,In_158);
nand U1239 (N_1239,In_1379,In_1445);
or U1240 (N_1240,N_531,N_184);
and U1241 (N_1241,In_649,N_897);
nor U1242 (N_1242,In_1035,N_620);
and U1243 (N_1243,N_41,N_541);
nand U1244 (N_1244,In_766,In_125);
nand U1245 (N_1245,N_974,N_580);
nor U1246 (N_1246,N_903,In_870);
and U1247 (N_1247,In_149,In_1451);
and U1248 (N_1248,N_791,In_988);
nor U1249 (N_1249,N_532,In_1068);
nor U1250 (N_1250,N_1077,N_285);
and U1251 (N_1251,N_103,N_50);
and U1252 (N_1252,N_967,N_951);
nor U1253 (N_1253,In_1649,N_166);
or U1254 (N_1254,In_1562,N_362);
and U1255 (N_1255,N_1179,In_1717);
nor U1256 (N_1256,N_482,N_959);
or U1257 (N_1257,In_1915,N_1103);
nand U1258 (N_1258,In_538,N_1215);
nor U1259 (N_1259,N_638,N_1230);
or U1260 (N_1260,N_534,N_1191);
or U1261 (N_1261,N_801,N_384);
or U1262 (N_1262,N_1117,In_807);
or U1263 (N_1263,N_491,N_835);
nor U1264 (N_1264,N_829,N_899);
nor U1265 (N_1265,N_736,N_1159);
nand U1266 (N_1266,N_1130,N_517);
and U1267 (N_1267,N_812,N_1050);
xor U1268 (N_1268,In_1202,N_1248);
and U1269 (N_1269,In_1083,N_1161);
xnor U1270 (N_1270,N_764,In_1737);
nand U1271 (N_1271,N_1137,N_1056);
nor U1272 (N_1272,N_1058,In_1745);
nand U1273 (N_1273,N_225,In_580);
and U1274 (N_1274,N_1175,N_1151);
or U1275 (N_1275,N_984,N_1220);
and U1276 (N_1276,N_1008,N_1125);
or U1277 (N_1277,N_428,N_1210);
nand U1278 (N_1278,N_577,In_331);
or U1279 (N_1279,N_1106,In_1078);
nand U1280 (N_1280,N_5,N_1089);
and U1281 (N_1281,N_1177,N_1239);
xnor U1282 (N_1282,N_502,In_208);
or U1283 (N_1283,In_1358,N_309);
nor U1284 (N_1284,N_1073,In_296);
nand U1285 (N_1285,N_239,In_1560);
xnor U1286 (N_1286,In_1863,In_536);
nand U1287 (N_1287,N_1176,N_1240);
and U1288 (N_1288,N_334,N_1232);
or U1289 (N_1289,N_1084,N_1123);
nor U1290 (N_1290,N_342,In_182);
xnor U1291 (N_1291,N_1134,N_1012);
or U1292 (N_1292,N_783,N_1133);
and U1293 (N_1293,In_295,In_756);
nand U1294 (N_1294,In_410,N_1102);
nor U1295 (N_1295,N_625,In_1153);
and U1296 (N_1296,N_1242,N_1066);
xor U1297 (N_1297,In_1079,In_903);
nor U1298 (N_1298,In_1720,In_1988);
and U1299 (N_1299,N_477,N_1227);
nand U1300 (N_1300,N_1040,N_1092);
nand U1301 (N_1301,N_1249,N_1153);
nor U1302 (N_1302,N_283,In_1314);
xnor U1303 (N_1303,N_785,In_504);
nor U1304 (N_1304,N_1088,N_598);
and U1305 (N_1305,N_1083,N_1141);
or U1306 (N_1306,N_911,N_1039);
and U1307 (N_1307,N_1054,N_1035);
or U1308 (N_1308,N_485,N_1079);
nand U1309 (N_1309,In_1248,N_977);
nor U1310 (N_1310,In_7,In_421);
or U1311 (N_1311,N_364,N_1162);
nor U1312 (N_1312,In_1367,N_551);
nor U1313 (N_1313,In_74,In_1086);
nand U1314 (N_1314,N_1051,In_66);
nor U1315 (N_1315,N_591,In_1137);
xnor U1316 (N_1316,N_1096,N_1075);
nor U1317 (N_1317,In_301,N_575);
or U1318 (N_1318,N_1140,In_242);
or U1319 (N_1319,N_437,N_1033);
and U1320 (N_1320,In_565,N_993);
and U1321 (N_1321,In_557,N_821);
xnor U1322 (N_1322,N_792,N_576);
and U1323 (N_1323,N_770,N_1048);
nand U1324 (N_1324,In_1651,N_514);
nor U1325 (N_1325,N_134,N_1150);
nand U1326 (N_1326,N_251,N_1241);
nand U1327 (N_1327,N_1104,N_354);
nand U1328 (N_1328,In_1167,N_68);
nand U1329 (N_1329,N_860,N_267);
nor U1330 (N_1330,In_253,In_707);
nand U1331 (N_1331,N_1010,In_495);
or U1332 (N_1332,N_952,N_563);
and U1333 (N_1333,N_846,In_693);
or U1334 (N_1334,N_840,In_1458);
nand U1335 (N_1335,In_875,In_35);
xor U1336 (N_1336,N_111,N_825);
nor U1337 (N_1337,In_194,N_1028);
nand U1338 (N_1338,N_549,In_306);
nand U1339 (N_1339,In_612,N_1086);
nor U1340 (N_1340,N_1041,N_823);
xor U1341 (N_1341,N_836,N_1112);
nor U1342 (N_1342,N_1098,In_1489);
nor U1343 (N_1343,N_1032,N_1234);
or U1344 (N_1344,N_1065,N_1168);
or U1345 (N_1345,In_174,N_278);
nor U1346 (N_1346,In_1162,N_492);
nor U1347 (N_1347,N_456,In_464);
nand U1348 (N_1348,N_486,N_1166);
nor U1349 (N_1349,N_425,N_1223);
nand U1350 (N_1350,N_568,N_644);
nand U1351 (N_1351,N_1085,In_1816);
nand U1352 (N_1352,N_814,N_19);
xnor U1353 (N_1353,In_354,N_191);
nand U1354 (N_1354,In_52,N_582);
or U1355 (N_1355,In_1921,N_433);
nand U1356 (N_1356,In_1641,N_1091);
or U1357 (N_1357,N_1113,N_1205);
xor U1358 (N_1358,N_725,In_87);
nor U1359 (N_1359,In_214,N_681);
nor U1360 (N_1360,In_906,N_478);
and U1361 (N_1361,N_1059,In_735);
or U1362 (N_1362,N_1093,In_1284);
nand U1363 (N_1363,N_1030,N_1131);
or U1364 (N_1364,In_534,N_893);
xnor U1365 (N_1365,In_490,N_1067);
nand U1366 (N_1366,N_780,In_1286);
xnor U1367 (N_1367,N_537,In_896);
nand U1368 (N_1368,N_1029,N_654);
nor U1369 (N_1369,In_278,N_1064);
or U1370 (N_1370,N_1170,N_1146);
and U1371 (N_1371,N_1148,N_242);
nor U1372 (N_1372,N_686,N_1026);
nand U1373 (N_1373,N_808,N_1174);
nor U1374 (N_1374,N_841,N_1023);
or U1375 (N_1375,In_1714,In_1494);
or U1376 (N_1376,N_1221,N_894);
xor U1377 (N_1377,N_1228,In_277);
nand U1378 (N_1378,In_746,N_1024);
and U1379 (N_1379,In_879,In_200);
nor U1380 (N_1380,In_589,N_120);
or U1381 (N_1381,In_701,N_596);
xor U1382 (N_1382,N_622,N_249);
nor U1383 (N_1383,N_398,N_805);
and U1384 (N_1384,In_316,In_1057);
or U1385 (N_1385,N_513,N_126);
or U1386 (N_1386,N_1018,N_1081);
or U1387 (N_1387,N_1087,N_1114);
and U1388 (N_1388,In_1931,N_357);
nor U1389 (N_1389,N_385,N_987);
nand U1390 (N_1390,In_442,N_28);
or U1391 (N_1391,In_853,N_954);
nand U1392 (N_1392,In_427,N_296);
xnor U1393 (N_1393,N_412,N_869);
and U1394 (N_1394,N_655,N_778);
and U1395 (N_1395,In_1661,N_51);
nor U1396 (N_1396,In_808,In_439);
or U1397 (N_1397,N_1057,N_341);
nor U1398 (N_1398,N_968,N_1129);
nand U1399 (N_1399,In_388,In_1225);
and U1400 (N_1400,N_1155,N_772);
and U1401 (N_1401,N_472,N_476);
or U1402 (N_1402,N_1198,N_146);
or U1403 (N_1403,N_1017,N_613);
nor U1404 (N_1404,N_793,N_1235);
or U1405 (N_1405,In_338,In_133);
nand U1406 (N_1406,N_464,In_1970);
nand U1407 (N_1407,N_1007,N_1244);
xnor U1408 (N_1408,N_1072,N_1216);
and U1409 (N_1409,N_1208,In_1644);
and U1410 (N_1410,N_651,N_958);
nor U1411 (N_1411,N_819,In_238);
xor U1412 (N_1412,N_912,N_1124);
or U1413 (N_1413,N_263,In_1221);
nor U1414 (N_1414,In_342,N_902);
nand U1415 (N_1415,N_179,In_1485);
nand U1416 (N_1416,N_1178,In_94);
and U1417 (N_1417,N_1013,N_895);
and U1418 (N_1418,N_605,N_975);
nand U1419 (N_1419,N_669,N_1052);
or U1420 (N_1420,In_1382,N_185);
nor U1421 (N_1421,In_788,N_765);
nor U1422 (N_1422,N_1211,N_543);
or U1423 (N_1423,In_679,N_944);
or U1424 (N_1424,N_410,N_1144);
nand U1425 (N_1425,N_480,N_1003);
nor U1426 (N_1426,N_1108,N_762);
or U1427 (N_1427,N_447,In_917);
or U1428 (N_1428,In_196,In_698);
and U1429 (N_1429,In_1854,N_129);
nand U1430 (N_1430,N_538,N_124);
or U1431 (N_1431,N_1009,N_1199);
or U1432 (N_1432,N_1021,N_1207);
xnor U1433 (N_1433,N_868,N_881);
or U1434 (N_1434,In_1335,N_652);
and U1435 (N_1435,N_924,N_752);
nand U1436 (N_1436,N_602,N_297);
or U1437 (N_1437,N_391,In_1322);
nand U1438 (N_1438,N_740,In_999);
nand U1439 (N_1439,N_779,N_1184);
nand U1440 (N_1440,In_564,In_1125);
nor U1441 (N_1441,N_976,N_601);
or U1442 (N_1442,N_934,N_1193);
nand U1443 (N_1443,N_1145,N_883);
or U1444 (N_1444,N_1213,N_540);
xor U1445 (N_1445,In_1640,N_905);
nor U1446 (N_1446,N_1107,N_630);
and U1447 (N_1447,N_670,N_744);
and U1448 (N_1448,N_887,N_200);
xnor U1449 (N_1449,N_904,N_1233);
or U1450 (N_1450,N_1080,In_952);
nor U1451 (N_1451,In_1103,N_929);
or U1452 (N_1452,N_603,N_1187);
nor U1453 (N_1453,In_938,N_1042);
and U1454 (N_1454,N_511,N_863);
xor U1455 (N_1455,N_1231,In_963);
or U1456 (N_1456,N_1061,N_1095);
and U1457 (N_1457,N_928,N_1180);
nand U1458 (N_1458,N_879,N_1025);
and U1459 (N_1459,N_57,N_978);
and U1460 (N_1460,N_939,N_1015);
nor U1461 (N_1461,In_183,N_1225);
or U1462 (N_1462,N_272,In_1568);
nand U1463 (N_1463,N_1120,N_197);
and U1464 (N_1464,N_550,In_1257);
and U1465 (N_1465,In_132,In_831);
and U1466 (N_1466,In_1898,N_1245);
xnor U1467 (N_1467,N_990,N_1060);
and U1468 (N_1468,In_924,In_758);
nand U1469 (N_1469,In_216,N_880);
nand U1470 (N_1470,N_289,N_946);
nor U1471 (N_1471,In_1762,In_1796);
nand U1472 (N_1472,In_943,N_1094);
nor U1473 (N_1473,N_16,In_115);
nor U1474 (N_1474,N_1063,In_1853);
or U1475 (N_1475,N_186,N_1229);
nor U1476 (N_1476,N_328,N_1062);
or U1477 (N_1477,N_1111,N_790);
nor U1478 (N_1478,In_1511,N_1069);
xor U1479 (N_1479,N_646,In_1003);
or U1480 (N_1480,N_913,N_31);
and U1481 (N_1481,In_955,N_694);
and U1482 (N_1482,N_506,N_302);
or U1483 (N_1483,N_1090,N_182);
or U1484 (N_1484,In_1152,N_290);
nand U1485 (N_1485,N_1194,In_458);
xnor U1486 (N_1486,N_676,In_1019);
nor U1487 (N_1487,N_1217,N_665);
or U1488 (N_1488,In_832,In_143);
nand U1489 (N_1489,N_1158,In_259);
or U1490 (N_1490,In_418,N_969);
and U1491 (N_1491,N_807,In_251);
nand U1492 (N_1492,N_1157,N_1004);
and U1493 (N_1493,In_1869,In_895);
nand U1494 (N_1494,N_158,In_1300);
and U1495 (N_1495,In_286,N_1099);
xnor U1496 (N_1496,N_989,In_1423);
and U1497 (N_1497,In_1091,N_1147);
nor U1498 (N_1498,N_1139,N_170);
or U1499 (N_1499,N_1183,N_1047);
nor U1500 (N_1500,N_1373,N_1493);
xnor U1501 (N_1501,N_1045,In_1545);
or U1502 (N_1502,N_1399,N_1014);
and U1503 (N_1503,N_775,N_1238);
nor U1504 (N_1504,N_1261,N_1381);
nor U1505 (N_1505,N_1423,N_196);
nand U1506 (N_1506,N_1353,N_995);
nand U1507 (N_1507,N_777,N_505);
nand U1508 (N_1508,N_1407,N_1386);
nor U1509 (N_1509,N_498,N_963);
xnor U1510 (N_1510,N_435,In_359);
and U1511 (N_1511,N_1326,In_1910);
nand U1512 (N_1512,N_1189,N_1218);
xor U1513 (N_1513,N_1222,N_1446);
or U1514 (N_1514,N_1396,N_1377);
and U1515 (N_1515,N_1343,In_1706);
nor U1516 (N_1516,N_1331,N_1404);
and U1517 (N_1517,N_1408,N_1195);
nor U1518 (N_1518,N_1055,In_1686);
and U1519 (N_1519,N_1119,In_654);
or U1520 (N_1520,N_1308,N_1302);
nand U1521 (N_1521,N_1101,N_1348);
and U1522 (N_1522,N_1031,In_1882);
nand U1523 (N_1523,N_1169,N_722);
nor U1524 (N_1524,N_973,In_1160);
nor U1525 (N_1525,In_1872,N_1280);
nand U1526 (N_1526,N_1226,N_1132);
and U1527 (N_1527,In_1082,N_1477);
or U1528 (N_1528,N_1478,N_351);
nor U1529 (N_1529,N_1305,N_1461);
nand U1530 (N_1530,N_1451,N_1224);
nor U1531 (N_1531,N_1398,N_1285);
or U1532 (N_1532,N_1277,In_997);
and U1533 (N_1533,N_878,N_1078);
nand U1534 (N_1534,In_1668,N_1206);
nand U1535 (N_1535,In_1199,In_1611);
nand U1536 (N_1536,N_1254,N_1071);
nor U1537 (N_1537,N_1273,N_373);
nand U1538 (N_1538,N_1251,N_1459);
nor U1539 (N_1539,N_1259,N_1068);
and U1540 (N_1540,N_1264,N_281);
and U1541 (N_1541,N_1363,N_1383);
and U1542 (N_1542,N_1143,N_202);
nor U1543 (N_1543,N_1197,N_633);
and U1544 (N_1544,In_1333,N_970);
nand U1545 (N_1545,N_1447,N_1289);
and U1546 (N_1546,N_1488,N_898);
nor U1547 (N_1547,N_1214,In_272);
nor U1548 (N_1548,N_1304,N_1498);
nor U1549 (N_1549,N_1299,N_508);
or U1550 (N_1550,N_1483,N_1118);
nand U1551 (N_1551,N_1499,N_1345);
or U1552 (N_1552,N_1374,N_1414);
nand U1553 (N_1553,N_1329,N_1318);
or U1554 (N_1554,N_1434,N_1371);
or U1555 (N_1555,N_1460,N_1444);
and U1556 (N_1556,In_126,N_1163);
or U1557 (N_1557,In_1330,N_1246);
nor U1558 (N_1558,N_1171,N_1422);
xnor U1559 (N_1559,N_1384,N_1327);
and U1560 (N_1560,N_1458,N_529);
nor U1561 (N_1561,N_1209,In_634);
nand U1562 (N_1562,N_1173,N_820);
and U1563 (N_1563,In_1801,N_1445);
and U1564 (N_1564,N_1385,N_1260);
nand U1565 (N_1565,N_1367,N_1462);
or U1566 (N_1566,N_1387,N_1351);
nor U1567 (N_1567,N_1270,N_1036);
and U1568 (N_1568,N_1271,N_1418);
nor U1569 (N_1569,N_949,In_1972);
nor U1570 (N_1570,N_1037,N_1294);
or U1571 (N_1571,N_229,In_1534);
and U1572 (N_1572,N_1312,N_1027);
and U1573 (N_1573,N_1400,N_732);
xor U1574 (N_1574,N_729,N_1201);
and U1575 (N_1575,N_1243,N_1473);
xnor U1576 (N_1576,N_4,N_1466);
and U1577 (N_1577,N_1164,N_1441);
nand U1578 (N_1578,N_849,N_1338);
and U1579 (N_1579,N_853,N_1339);
nand U1580 (N_1580,N_1272,N_985);
xnor U1581 (N_1581,N_1410,N_1278);
or U1582 (N_1582,In_1502,N_1265);
nand U1583 (N_1583,N_1456,N_1049);
nand U1584 (N_1584,N_658,N_1463);
nand U1585 (N_1585,N_1464,N_1297);
nand U1586 (N_1586,N_886,N_1282);
nor U1587 (N_1587,N_150,N_1350);
nand U1588 (N_1588,N_822,N_1333);
nand U1589 (N_1589,N_1300,N_463);
nand U1590 (N_1590,N_1469,N_1496);
or U1591 (N_1591,N_992,N_1330);
nor U1592 (N_1592,N_552,N_1420);
nand U1593 (N_1593,N_1472,N_826);
xnor U1594 (N_1594,N_1255,N_1307);
and U1595 (N_1595,N_813,N_1165);
nand U1596 (N_1596,N_419,N_910);
or U1597 (N_1597,N_1480,N_845);
and U1598 (N_1598,In_1133,N_1324);
and U1599 (N_1599,N_1354,N_1303);
nor U1600 (N_1600,N_1253,N_936);
nand U1601 (N_1601,N_1346,N_1403);
and U1602 (N_1602,N_1484,N_800);
or U1603 (N_1603,N_1368,N_1274);
and U1604 (N_1604,N_1154,In_1048);
or U1605 (N_1605,In_1587,N_1430);
or U1606 (N_1606,N_720,N_1428);
or U1607 (N_1607,N_1448,N_997);
xnor U1608 (N_1608,N_1136,N_1156);
or U1609 (N_1609,N_1236,N_75);
and U1610 (N_1610,N_1293,N_1311);
and U1611 (N_1611,In_1508,N_1290);
and U1612 (N_1612,N_1122,N_1135);
xnor U1613 (N_1613,N_1167,In_1842);
nor U1614 (N_1614,N_933,In_474);
nor U1615 (N_1615,N_1370,N_1449);
and U1616 (N_1616,N_1355,In_1905);
and U1617 (N_1617,N_1453,N_201);
nor U1618 (N_1618,In_1713,N_1389);
nand U1619 (N_1619,N_991,N_1126);
or U1620 (N_1620,N_1405,N_1316);
and U1621 (N_1621,N_1347,N_1203);
nand U1622 (N_1622,N_1436,N_1314);
nand U1623 (N_1623,N_1313,N_1283);
or U1624 (N_1624,N_1391,N_1497);
xor U1625 (N_1625,N_1247,N_1252);
and U1626 (N_1626,N_359,N_1421);
nand U1627 (N_1627,N_1020,N_1409);
nor U1628 (N_1628,N_1002,N_794);
nor U1629 (N_1629,N_1328,N_1425);
and U1630 (N_1630,N_1429,In_731);
nor U1631 (N_1631,N_639,N_1366);
nor U1632 (N_1632,N_1397,In_856);
nor U1633 (N_1633,N_280,N_1358);
nand U1634 (N_1634,N_1127,N_1298);
nand U1635 (N_1635,N_1301,N_310);
and U1636 (N_1636,N_1019,In_248);
nor U1637 (N_1637,N_627,N_1279);
nand U1638 (N_1638,N_1188,N_217);
or U1639 (N_1639,N_1100,N_1263);
nor U1640 (N_1640,N_1186,N_1142);
or U1641 (N_1641,N_1288,In_716);
or U1642 (N_1642,N_1250,N_1426);
or U1643 (N_1643,N_1412,N_920);
and U1644 (N_1644,N_1401,In_1241);
nand U1645 (N_1645,In_723,N_1492);
nand U1646 (N_1646,N_1292,N_1435);
nand U1647 (N_1647,N_1276,N_1364);
or U1648 (N_1648,N_1378,N_1196);
nor U1649 (N_1649,In_1565,N_1262);
and U1650 (N_1650,N_1237,N_1415);
nor U1651 (N_1651,N_1306,N_1190);
nor U1652 (N_1652,N_957,N_501);
nand U1653 (N_1653,N_1392,N_1138);
nand U1654 (N_1654,N_1485,N_1471);
nor U1655 (N_1655,N_1432,N_1390);
nor U1656 (N_1656,N_1006,N_1320);
nand U1657 (N_1657,N_1382,N_1487);
nand U1658 (N_1658,In_1223,N_1424);
nand U1659 (N_1659,N_1388,N_1417);
nand U1660 (N_1660,N_1212,N_1431);
and U1661 (N_1661,N_1110,N_1437);
or U1662 (N_1662,N_1105,N_1433);
xnor U1663 (N_1663,N_1044,N_1411);
nor U1664 (N_1664,N_1475,N_1267);
xnor U1665 (N_1665,N_931,N_1481);
nor U1666 (N_1666,In_1780,N_1393);
nand U1667 (N_1667,In_1049,N_1349);
and U1668 (N_1668,N_1467,N_1286);
or U1669 (N_1669,N_889,N_350);
or U1670 (N_1670,N_1321,N_1257);
nor U1671 (N_1671,N_172,In_1235);
nand U1672 (N_1672,N_1309,N_1319);
nand U1673 (N_1673,N_1185,N_1005);
xnor U1674 (N_1674,N_1332,N_1325);
or U1675 (N_1675,N_1340,N_1457);
or U1676 (N_1676,N_1315,N_1001);
nand U1677 (N_1677,N_1256,N_1356);
or U1678 (N_1678,In_225,N_1016);
nor U1679 (N_1679,N_1317,N_1310);
nand U1680 (N_1680,N_885,N_1360);
or U1681 (N_1681,N_1287,N_1082);
nand U1682 (N_1682,N_1336,N_972);
or U1683 (N_1683,N_142,In_1834);
nor U1684 (N_1684,N_1070,N_1439);
or U1685 (N_1685,N_1352,N_1097);
or U1686 (N_1686,N_1474,N_810);
and U1687 (N_1687,N_1258,N_519);
nor U1688 (N_1688,N_1490,N_1116);
nor U1689 (N_1689,N_955,N_1269);
or U1690 (N_1690,In_872,In_168);
xnor U1691 (N_1691,N_1375,N_1034);
xnor U1692 (N_1692,N_1275,N_1491);
nor U1693 (N_1693,N_1323,N_1043);
or U1694 (N_1694,N_907,N_1341);
nand U1695 (N_1695,In_535,N_1115);
nand U1696 (N_1696,N_1172,N_1402);
xnor U1697 (N_1697,N_930,N_1416);
nand U1698 (N_1698,N_1266,N_628);
nor U1699 (N_1699,N_1204,In_1374);
nand U1700 (N_1700,N_1342,In_337);
or U1701 (N_1701,N_154,In_71);
and U1702 (N_1702,N_680,N_1121);
nand U1703 (N_1703,N_1494,N_966);
xnor U1704 (N_1704,N_1486,In_323);
and U1705 (N_1705,In_1253,In_412);
or U1706 (N_1706,N_1470,In_982);
nand U1707 (N_1707,N_769,N_1365);
xnor U1708 (N_1708,N_1395,N_240);
nand U1709 (N_1709,N_1443,In_14);
nor U1710 (N_1710,N_1489,N_1053);
xor U1711 (N_1711,N_468,N_1046);
nand U1712 (N_1712,N_1284,N_1022);
or U1713 (N_1713,N_1011,N_610);
and U1714 (N_1714,N_451,In_452);
nor U1715 (N_1715,N_1476,N_1192);
nand U1716 (N_1716,N_1291,N_1482);
or U1717 (N_1717,N_1376,N_1357);
xnor U1718 (N_1718,N_1419,N_1362);
nand U1719 (N_1719,In_1096,N_1344);
nor U1720 (N_1720,N_1413,N_833);
and U1721 (N_1721,N_1406,N_925);
nand U1722 (N_1722,N_1465,N_1479);
nor U1723 (N_1723,N_13,N_1152);
nand U1724 (N_1724,N_659,N_1200);
nand U1725 (N_1725,N_1219,N_1268);
nor U1726 (N_1726,N_1468,N_1322);
or U1727 (N_1727,N_1394,N_1455);
nor U1728 (N_1728,In_38,N_213);
nand U1729 (N_1729,N_1128,In_874);
xor U1730 (N_1730,N_1334,N_1450);
and U1731 (N_1731,N_58,N_1372);
and U1732 (N_1732,N_1369,N_1109);
or U1733 (N_1733,N_1454,In_51);
nor U1734 (N_1734,N_1149,N_1452);
nand U1735 (N_1735,N_1160,N_282);
nand U1736 (N_1736,N_1295,N_1076);
xor U1737 (N_1737,N_871,N_1442);
and U1738 (N_1738,N_1038,N_365);
and U1739 (N_1739,N_1379,In_1243);
xnor U1740 (N_1740,N_1495,N_496);
xor U1741 (N_1741,N_1000,N_1335);
and U1742 (N_1742,N_1182,N_1440);
nor U1743 (N_1743,N_1380,N_1181);
or U1744 (N_1744,N_1361,N_1202);
nand U1745 (N_1745,N_699,N_1337);
or U1746 (N_1746,N_1427,N_1438);
and U1747 (N_1747,N_1074,N_1359);
nor U1748 (N_1748,N_1281,N_429);
and U1749 (N_1749,In_1175,N_1296);
or U1750 (N_1750,N_1651,N_1528);
or U1751 (N_1751,N_1516,N_1514);
or U1752 (N_1752,N_1653,N_1619);
nor U1753 (N_1753,N_1676,N_1584);
nand U1754 (N_1754,N_1596,N_1644);
and U1755 (N_1755,N_1592,N_1606);
and U1756 (N_1756,N_1590,N_1525);
or U1757 (N_1757,N_1522,N_1695);
and U1758 (N_1758,N_1730,N_1721);
nand U1759 (N_1759,N_1690,N_1501);
nand U1760 (N_1760,N_1569,N_1649);
and U1761 (N_1761,N_1663,N_1685);
nor U1762 (N_1762,N_1684,N_1616);
or U1763 (N_1763,N_1548,N_1586);
or U1764 (N_1764,N_1518,N_1531);
and U1765 (N_1765,N_1521,N_1669);
nor U1766 (N_1766,N_1538,N_1739);
or U1767 (N_1767,N_1723,N_1541);
or U1768 (N_1768,N_1603,N_1642);
nor U1769 (N_1769,N_1577,N_1626);
xnor U1770 (N_1770,N_1713,N_1503);
nor U1771 (N_1771,N_1561,N_1720);
nor U1772 (N_1772,N_1706,N_1562);
xor U1773 (N_1773,N_1623,N_1542);
xnor U1774 (N_1774,N_1563,N_1637);
or U1775 (N_1775,N_1575,N_1696);
nor U1776 (N_1776,N_1520,N_1735);
and U1777 (N_1777,N_1677,N_1634);
nor U1778 (N_1778,N_1682,N_1574);
and U1779 (N_1779,N_1661,N_1741);
nor U1780 (N_1780,N_1728,N_1727);
nand U1781 (N_1781,N_1511,N_1567);
xnor U1782 (N_1782,N_1745,N_1607);
and U1783 (N_1783,N_1698,N_1549);
and U1784 (N_1784,N_1578,N_1565);
and U1785 (N_1785,N_1658,N_1533);
nand U1786 (N_1786,N_1620,N_1704);
nor U1787 (N_1787,N_1570,N_1654);
and U1788 (N_1788,N_1614,N_1517);
nand U1789 (N_1789,N_1504,N_1641);
or U1790 (N_1790,N_1609,N_1679);
or U1791 (N_1791,N_1568,N_1532);
nor U1792 (N_1792,N_1710,N_1546);
and U1793 (N_1793,N_1559,N_1582);
xnor U1794 (N_1794,N_1736,N_1711);
nand U1795 (N_1795,N_1618,N_1712);
or U1796 (N_1796,N_1699,N_1656);
xnor U1797 (N_1797,N_1600,N_1645);
nand U1798 (N_1798,N_1719,N_1724);
nand U1799 (N_1799,N_1508,N_1675);
nand U1800 (N_1800,N_1547,N_1691);
or U1801 (N_1801,N_1558,N_1689);
and U1802 (N_1802,N_1500,N_1572);
nor U1803 (N_1803,N_1680,N_1709);
or U1804 (N_1804,N_1673,N_1581);
and U1805 (N_1805,N_1513,N_1705);
nand U1806 (N_1806,N_1560,N_1718);
xnor U1807 (N_1807,N_1657,N_1613);
nand U1808 (N_1808,N_1536,N_1544);
nor U1809 (N_1809,N_1640,N_1507);
xor U1810 (N_1810,N_1509,N_1707);
xnor U1811 (N_1811,N_1540,N_1693);
and U1812 (N_1812,N_1744,N_1672);
nand U1813 (N_1813,N_1612,N_1697);
or U1814 (N_1814,N_1556,N_1597);
nor U1815 (N_1815,N_1716,N_1725);
and U1816 (N_1816,N_1633,N_1650);
nand U1817 (N_1817,N_1551,N_1731);
nor U1818 (N_1818,N_1740,N_1576);
nor U1819 (N_1819,N_1608,N_1545);
nand U1820 (N_1820,N_1628,N_1598);
nand U1821 (N_1821,N_1733,N_1749);
and U1822 (N_1822,N_1692,N_1638);
nor U1823 (N_1823,N_1646,N_1652);
and U1824 (N_1824,N_1564,N_1585);
and U1825 (N_1825,N_1694,N_1587);
or U1826 (N_1826,N_1671,N_1665);
nand U1827 (N_1827,N_1535,N_1664);
and U1828 (N_1828,N_1553,N_1687);
nand U1829 (N_1829,N_1539,N_1571);
or U1830 (N_1830,N_1742,N_1523);
nor U1831 (N_1831,N_1670,N_1660);
nor U1832 (N_1832,N_1537,N_1593);
nand U1833 (N_1833,N_1737,N_1519);
or U1834 (N_1834,N_1550,N_1595);
and U1835 (N_1835,N_1583,N_1580);
and U1836 (N_1836,N_1747,N_1717);
or U1837 (N_1837,N_1636,N_1529);
or U1838 (N_1838,N_1502,N_1617);
or U1839 (N_1839,N_1611,N_1715);
nor U1840 (N_1840,N_1674,N_1630);
or U1841 (N_1841,N_1534,N_1743);
and U1842 (N_1842,N_1621,N_1594);
or U1843 (N_1843,N_1734,N_1635);
nor U1844 (N_1844,N_1667,N_1668);
or U1845 (N_1845,N_1588,N_1708);
and U1846 (N_1846,N_1659,N_1748);
nand U1847 (N_1847,N_1515,N_1624);
xnor U1848 (N_1848,N_1554,N_1732);
nor U1849 (N_1849,N_1589,N_1599);
and U1850 (N_1850,N_1530,N_1681);
nor U1851 (N_1851,N_1566,N_1622);
xor U1852 (N_1852,N_1639,N_1543);
or U1853 (N_1853,N_1746,N_1527);
or U1854 (N_1854,N_1510,N_1648);
nor U1855 (N_1855,N_1647,N_1601);
nor U1856 (N_1856,N_1625,N_1512);
and U1857 (N_1857,N_1683,N_1591);
xor U1858 (N_1858,N_1662,N_1573);
nor U1859 (N_1859,N_1738,N_1714);
nor U1860 (N_1860,N_1703,N_1700);
or U1861 (N_1861,N_1686,N_1643);
nor U1862 (N_1862,N_1655,N_1631);
or U1863 (N_1863,N_1701,N_1678);
or U1864 (N_1864,N_1506,N_1666);
or U1865 (N_1865,N_1602,N_1557);
and U1866 (N_1866,N_1605,N_1610);
xnor U1867 (N_1867,N_1552,N_1579);
or U1868 (N_1868,N_1629,N_1615);
and U1869 (N_1869,N_1604,N_1688);
nand U1870 (N_1870,N_1505,N_1632);
nor U1871 (N_1871,N_1729,N_1722);
or U1872 (N_1872,N_1555,N_1627);
nor U1873 (N_1873,N_1726,N_1702);
and U1874 (N_1874,N_1526,N_1524);
nand U1875 (N_1875,N_1642,N_1605);
nor U1876 (N_1876,N_1515,N_1726);
and U1877 (N_1877,N_1503,N_1656);
or U1878 (N_1878,N_1663,N_1658);
xor U1879 (N_1879,N_1622,N_1640);
xor U1880 (N_1880,N_1589,N_1580);
or U1881 (N_1881,N_1709,N_1556);
xor U1882 (N_1882,N_1665,N_1609);
nor U1883 (N_1883,N_1507,N_1605);
nand U1884 (N_1884,N_1621,N_1606);
xor U1885 (N_1885,N_1728,N_1627);
xor U1886 (N_1886,N_1555,N_1701);
nand U1887 (N_1887,N_1688,N_1676);
nand U1888 (N_1888,N_1738,N_1626);
nand U1889 (N_1889,N_1746,N_1647);
nor U1890 (N_1890,N_1688,N_1706);
and U1891 (N_1891,N_1674,N_1571);
or U1892 (N_1892,N_1576,N_1738);
xnor U1893 (N_1893,N_1669,N_1661);
xnor U1894 (N_1894,N_1539,N_1578);
or U1895 (N_1895,N_1644,N_1605);
nand U1896 (N_1896,N_1654,N_1583);
and U1897 (N_1897,N_1703,N_1643);
or U1898 (N_1898,N_1598,N_1561);
nand U1899 (N_1899,N_1686,N_1584);
or U1900 (N_1900,N_1570,N_1529);
nand U1901 (N_1901,N_1694,N_1545);
or U1902 (N_1902,N_1743,N_1635);
and U1903 (N_1903,N_1653,N_1610);
nand U1904 (N_1904,N_1509,N_1719);
nand U1905 (N_1905,N_1712,N_1748);
nor U1906 (N_1906,N_1729,N_1577);
and U1907 (N_1907,N_1721,N_1716);
nor U1908 (N_1908,N_1558,N_1641);
or U1909 (N_1909,N_1636,N_1732);
nand U1910 (N_1910,N_1591,N_1590);
nor U1911 (N_1911,N_1709,N_1601);
or U1912 (N_1912,N_1748,N_1574);
nand U1913 (N_1913,N_1670,N_1692);
or U1914 (N_1914,N_1642,N_1503);
and U1915 (N_1915,N_1656,N_1612);
nor U1916 (N_1916,N_1646,N_1575);
and U1917 (N_1917,N_1670,N_1656);
or U1918 (N_1918,N_1698,N_1740);
or U1919 (N_1919,N_1565,N_1746);
or U1920 (N_1920,N_1565,N_1538);
or U1921 (N_1921,N_1559,N_1602);
or U1922 (N_1922,N_1507,N_1639);
nor U1923 (N_1923,N_1504,N_1578);
nand U1924 (N_1924,N_1562,N_1651);
or U1925 (N_1925,N_1535,N_1587);
nor U1926 (N_1926,N_1700,N_1729);
or U1927 (N_1927,N_1589,N_1686);
nor U1928 (N_1928,N_1659,N_1604);
or U1929 (N_1929,N_1545,N_1638);
nand U1930 (N_1930,N_1622,N_1623);
or U1931 (N_1931,N_1743,N_1680);
nand U1932 (N_1932,N_1664,N_1643);
xnor U1933 (N_1933,N_1571,N_1701);
nor U1934 (N_1934,N_1607,N_1723);
nor U1935 (N_1935,N_1558,N_1713);
nand U1936 (N_1936,N_1603,N_1585);
nand U1937 (N_1937,N_1648,N_1600);
or U1938 (N_1938,N_1552,N_1530);
xor U1939 (N_1939,N_1729,N_1571);
or U1940 (N_1940,N_1541,N_1546);
nand U1941 (N_1941,N_1585,N_1544);
nand U1942 (N_1942,N_1662,N_1747);
nor U1943 (N_1943,N_1585,N_1723);
nor U1944 (N_1944,N_1644,N_1507);
and U1945 (N_1945,N_1658,N_1734);
and U1946 (N_1946,N_1649,N_1727);
nor U1947 (N_1947,N_1588,N_1694);
or U1948 (N_1948,N_1723,N_1603);
nand U1949 (N_1949,N_1720,N_1617);
nor U1950 (N_1950,N_1558,N_1500);
and U1951 (N_1951,N_1661,N_1675);
or U1952 (N_1952,N_1522,N_1587);
nand U1953 (N_1953,N_1741,N_1574);
nand U1954 (N_1954,N_1620,N_1594);
nor U1955 (N_1955,N_1608,N_1544);
nand U1956 (N_1956,N_1605,N_1681);
xor U1957 (N_1957,N_1581,N_1505);
nand U1958 (N_1958,N_1611,N_1574);
or U1959 (N_1959,N_1740,N_1629);
nor U1960 (N_1960,N_1694,N_1600);
or U1961 (N_1961,N_1538,N_1506);
and U1962 (N_1962,N_1541,N_1675);
nor U1963 (N_1963,N_1598,N_1583);
nor U1964 (N_1964,N_1564,N_1624);
and U1965 (N_1965,N_1515,N_1533);
or U1966 (N_1966,N_1713,N_1658);
nor U1967 (N_1967,N_1527,N_1532);
nor U1968 (N_1968,N_1594,N_1517);
or U1969 (N_1969,N_1660,N_1743);
and U1970 (N_1970,N_1714,N_1556);
nor U1971 (N_1971,N_1545,N_1616);
and U1972 (N_1972,N_1552,N_1647);
or U1973 (N_1973,N_1689,N_1667);
and U1974 (N_1974,N_1641,N_1531);
nand U1975 (N_1975,N_1632,N_1552);
or U1976 (N_1976,N_1734,N_1678);
nand U1977 (N_1977,N_1644,N_1725);
nor U1978 (N_1978,N_1633,N_1553);
nor U1979 (N_1979,N_1699,N_1587);
nor U1980 (N_1980,N_1724,N_1514);
nor U1981 (N_1981,N_1594,N_1667);
nand U1982 (N_1982,N_1525,N_1565);
nor U1983 (N_1983,N_1669,N_1743);
or U1984 (N_1984,N_1728,N_1692);
or U1985 (N_1985,N_1620,N_1541);
or U1986 (N_1986,N_1623,N_1626);
or U1987 (N_1987,N_1512,N_1724);
nand U1988 (N_1988,N_1686,N_1601);
nand U1989 (N_1989,N_1578,N_1538);
xor U1990 (N_1990,N_1639,N_1662);
or U1991 (N_1991,N_1526,N_1680);
nor U1992 (N_1992,N_1736,N_1661);
and U1993 (N_1993,N_1629,N_1580);
or U1994 (N_1994,N_1605,N_1620);
or U1995 (N_1995,N_1536,N_1699);
or U1996 (N_1996,N_1666,N_1534);
and U1997 (N_1997,N_1631,N_1643);
xor U1998 (N_1998,N_1745,N_1609);
xor U1999 (N_1999,N_1544,N_1520);
nand U2000 (N_2000,N_1842,N_1882);
or U2001 (N_2001,N_1754,N_1894);
nand U2002 (N_2002,N_1824,N_1815);
and U2003 (N_2003,N_1865,N_1752);
nand U2004 (N_2004,N_1839,N_1972);
xnor U2005 (N_2005,N_1834,N_1887);
and U2006 (N_2006,N_1927,N_1876);
or U2007 (N_2007,N_1860,N_1869);
nand U2008 (N_2008,N_1909,N_1758);
nor U2009 (N_2009,N_1976,N_1949);
nand U2010 (N_2010,N_1837,N_1898);
nand U2011 (N_2011,N_1796,N_1942);
nor U2012 (N_2012,N_1954,N_1995);
and U2013 (N_2013,N_1872,N_1757);
and U2014 (N_2014,N_1917,N_1870);
nor U2015 (N_2015,N_1924,N_1926);
nand U2016 (N_2016,N_1801,N_1921);
or U2017 (N_2017,N_1750,N_1768);
nand U2018 (N_2018,N_1775,N_1868);
nand U2019 (N_2019,N_1897,N_1987);
xnor U2020 (N_2020,N_1878,N_1845);
or U2021 (N_2021,N_1885,N_1804);
nand U2022 (N_2022,N_1879,N_1829);
nor U2023 (N_2023,N_1975,N_1831);
nor U2024 (N_2024,N_1998,N_1895);
and U2025 (N_2025,N_1828,N_1938);
or U2026 (N_2026,N_1812,N_1814);
nand U2027 (N_2027,N_1763,N_1803);
nand U2028 (N_2028,N_1772,N_1899);
and U2029 (N_2029,N_1910,N_1859);
nand U2030 (N_2030,N_1993,N_1939);
or U2031 (N_2031,N_1985,N_1811);
nor U2032 (N_2032,N_1932,N_1858);
xnor U2033 (N_2033,N_1988,N_1816);
xor U2034 (N_2034,N_1918,N_1767);
nand U2035 (N_2035,N_1861,N_1905);
nand U2036 (N_2036,N_1820,N_1959);
nor U2037 (N_2037,N_1990,N_1992);
nand U2038 (N_2038,N_1777,N_1883);
nor U2039 (N_2039,N_1760,N_1904);
and U2040 (N_2040,N_1956,N_1780);
nor U2041 (N_2041,N_1892,N_1840);
nor U2042 (N_2042,N_1886,N_1914);
nor U2043 (N_2043,N_1806,N_1844);
nand U2044 (N_2044,N_1873,N_1854);
nor U2045 (N_2045,N_1986,N_1761);
nand U2046 (N_2046,N_1929,N_1912);
and U2047 (N_2047,N_1769,N_1962);
nor U2048 (N_2048,N_1863,N_1771);
nand U2049 (N_2049,N_1825,N_1821);
nor U2050 (N_2050,N_1934,N_1981);
and U2051 (N_2051,N_1849,N_1784);
and U2052 (N_2052,N_1984,N_1953);
nor U2053 (N_2053,N_1813,N_1817);
nand U2054 (N_2054,N_1838,N_1915);
or U2055 (N_2055,N_1792,N_1952);
and U2056 (N_2056,N_1908,N_1770);
xnor U2057 (N_2057,N_1843,N_1787);
xor U2058 (N_2058,N_1928,N_1874);
or U2059 (N_2059,N_1794,N_1805);
and U2060 (N_2060,N_1946,N_1864);
or U2061 (N_2061,N_1753,N_1862);
nor U2062 (N_2062,N_1857,N_1989);
and U2063 (N_2063,N_1818,N_1835);
xor U2064 (N_2064,N_1901,N_1789);
nor U2065 (N_2065,N_1919,N_1766);
and U2066 (N_2066,N_1936,N_1931);
nand U2067 (N_2067,N_1965,N_1967);
nor U2068 (N_2068,N_1877,N_1977);
xnor U2069 (N_2069,N_1955,N_1798);
nor U2070 (N_2070,N_1832,N_1791);
or U2071 (N_2071,N_1764,N_1880);
xor U2072 (N_2072,N_1994,N_1925);
or U2073 (N_2073,N_1997,N_1996);
and U2074 (N_2074,N_1855,N_1999);
nand U2075 (N_2075,N_1937,N_1871);
nor U2076 (N_2076,N_1891,N_1762);
or U2077 (N_2077,N_1916,N_1941);
nor U2078 (N_2078,N_1948,N_1782);
or U2079 (N_2079,N_1776,N_1822);
nor U2080 (N_2080,N_1779,N_1961);
nand U2081 (N_2081,N_1795,N_1866);
xor U2082 (N_2082,N_1846,N_1841);
and U2083 (N_2083,N_1807,N_1968);
nand U2084 (N_2084,N_1833,N_1896);
and U2085 (N_2085,N_1852,N_1759);
nor U2086 (N_2086,N_1793,N_1935);
or U2087 (N_2087,N_1923,N_1930);
nor U2088 (N_2088,N_1893,N_1964);
or U2089 (N_2089,N_1907,N_1920);
nor U2090 (N_2090,N_1980,N_1966);
and U2091 (N_2091,N_1951,N_1853);
or U2092 (N_2092,N_1950,N_1808);
nand U2093 (N_2093,N_1755,N_1957);
xnor U2094 (N_2094,N_1756,N_1851);
xor U2095 (N_2095,N_1970,N_1790);
and U2096 (N_2096,N_1971,N_1765);
nand U2097 (N_2097,N_1922,N_1960);
and U2098 (N_2098,N_1800,N_1799);
xnor U2099 (N_2099,N_1963,N_1826);
or U2100 (N_2100,N_1786,N_1943);
xor U2101 (N_2101,N_1848,N_1773);
nor U2102 (N_2102,N_1850,N_1983);
and U2103 (N_2103,N_1781,N_1969);
and U2104 (N_2104,N_1774,N_1778);
xor U2105 (N_2105,N_1884,N_1900);
nand U2106 (N_2106,N_1973,N_1830);
xnor U2107 (N_2107,N_1856,N_1785);
nor U2108 (N_2108,N_1902,N_1978);
or U2109 (N_2109,N_1906,N_1889);
or U2110 (N_2110,N_1783,N_1947);
nand U2111 (N_2111,N_1958,N_1911);
or U2112 (N_2112,N_1881,N_1819);
nand U2113 (N_2113,N_1974,N_1979);
or U2114 (N_2114,N_1890,N_1944);
and U2115 (N_2115,N_1751,N_1888);
or U2116 (N_2116,N_1867,N_1788);
or U2117 (N_2117,N_1913,N_1991);
and U2118 (N_2118,N_1810,N_1802);
or U2119 (N_2119,N_1823,N_1847);
nand U2120 (N_2120,N_1940,N_1982);
or U2121 (N_2121,N_1836,N_1827);
nor U2122 (N_2122,N_1933,N_1797);
xnor U2123 (N_2123,N_1875,N_1903);
and U2124 (N_2124,N_1945,N_1809);
nor U2125 (N_2125,N_1886,N_1840);
nor U2126 (N_2126,N_1906,N_1860);
and U2127 (N_2127,N_1782,N_1997);
nor U2128 (N_2128,N_1769,N_1798);
and U2129 (N_2129,N_1849,N_1824);
nand U2130 (N_2130,N_1997,N_1761);
nand U2131 (N_2131,N_1848,N_1963);
nand U2132 (N_2132,N_1825,N_1779);
and U2133 (N_2133,N_1853,N_1868);
and U2134 (N_2134,N_1974,N_1881);
nor U2135 (N_2135,N_1810,N_1884);
nor U2136 (N_2136,N_1980,N_1989);
nor U2137 (N_2137,N_1906,N_1916);
xor U2138 (N_2138,N_1834,N_1796);
and U2139 (N_2139,N_1977,N_1994);
and U2140 (N_2140,N_1780,N_1931);
nor U2141 (N_2141,N_1912,N_1938);
nor U2142 (N_2142,N_1881,N_1846);
nor U2143 (N_2143,N_1886,N_1862);
nand U2144 (N_2144,N_1914,N_1878);
and U2145 (N_2145,N_1964,N_1925);
or U2146 (N_2146,N_1795,N_1935);
or U2147 (N_2147,N_1832,N_1888);
or U2148 (N_2148,N_1910,N_1832);
and U2149 (N_2149,N_1898,N_1856);
and U2150 (N_2150,N_1861,N_1776);
and U2151 (N_2151,N_1986,N_1768);
nor U2152 (N_2152,N_1854,N_1821);
and U2153 (N_2153,N_1809,N_1873);
nor U2154 (N_2154,N_1910,N_1775);
or U2155 (N_2155,N_1868,N_1917);
nor U2156 (N_2156,N_1802,N_1888);
nor U2157 (N_2157,N_1907,N_1992);
and U2158 (N_2158,N_1872,N_1920);
and U2159 (N_2159,N_1974,N_1799);
nand U2160 (N_2160,N_1889,N_1791);
and U2161 (N_2161,N_1955,N_1814);
and U2162 (N_2162,N_1960,N_1989);
nand U2163 (N_2163,N_1953,N_1931);
nand U2164 (N_2164,N_1980,N_1792);
or U2165 (N_2165,N_1814,N_1950);
nor U2166 (N_2166,N_1908,N_1973);
and U2167 (N_2167,N_1861,N_1834);
and U2168 (N_2168,N_1958,N_1791);
nor U2169 (N_2169,N_1845,N_1859);
nand U2170 (N_2170,N_1817,N_1836);
and U2171 (N_2171,N_1994,N_1970);
and U2172 (N_2172,N_1908,N_1889);
nor U2173 (N_2173,N_1899,N_1794);
or U2174 (N_2174,N_1804,N_1853);
or U2175 (N_2175,N_1819,N_1861);
nand U2176 (N_2176,N_1856,N_1800);
and U2177 (N_2177,N_1768,N_1887);
nor U2178 (N_2178,N_1789,N_1900);
xnor U2179 (N_2179,N_1761,N_1754);
and U2180 (N_2180,N_1768,N_1815);
nand U2181 (N_2181,N_1781,N_1821);
or U2182 (N_2182,N_1752,N_1915);
or U2183 (N_2183,N_1783,N_1821);
nor U2184 (N_2184,N_1878,N_1805);
or U2185 (N_2185,N_1931,N_1774);
nor U2186 (N_2186,N_1876,N_1806);
nand U2187 (N_2187,N_1786,N_1829);
nand U2188 (N_2188,N_1920,N_1756);
nand U2189 (N_2189,N_1754,N_1824);
nor U2190 (N_2190,N_1951,N_1989);
nor U2191 (N_2191,N_1929,N_1907);
and U2192 (N_2192,N_1955,N_1816);
nand U2193 (N_2193,N_1944,N_1838);
nand U2194 (N_2194,N_1810,N_1987);
or U2195 (N_2195,N_1974,N_1789);
or U2196 (N_2196,N_1751,N_1954);
or U2197 (N_2197,N_1923,N_1835);
or U2198 (N_2198,N_1971,N_1780);
or U2199 (N_2199,N_1874,N_1985);
and U2200 (N_2200,N_1962,N_1823);
or U2201 (N_2201,N_1948,N_1813);
or U2202 (N_2202,N_1932,N_1928);
and U2203 (N_2203,N_1853,N_1824);
and U2204 (N_2204,N_1898,N_1889);
nor U2205 (N_2205,N_1827,N_1772);
nor U2206 (N_2206,N_1847,N_1935);
and U2207 (N_2207,N_1894,N_1871);
nor U2208 (N_2208,N_1855,N_1813);
or U2209 (N_2209,N_1886,N_1851);
xor U2210 (N_2210,N_1898,N_1839);
nand U2211 (N_2211,N_1947,N_1831);
nor U2212 (N_2212,N_1911,N_1990);
or U2213 (N_2213,N_1878,N_1843);
nand U2214 (N_2214,N_1791,N_1790);
nor U2215 (N_2215,N_1853,N_1825);
or U2216 (N_2216,N_1786,N_1861);
nor U2217 (N_2217,N_1923,N_1984);
or U2218 (N_2218,N_1754,N_1774);
or U2219 (N_2219,N_1814,N_1898);
nor U2220 (N_2220,N_1985,N_1933);
or U2221 (N_2221,N_1837,N_1885);
and U2222 (N_2222,N_1899,N_1982);
xnor U2223 (N_2223,N_1990,N_1903);
xor U2224 (N_2224,N_1951,N_1995);
xor U2225 (N_2225,N_1846,N_1923);
xnor U2226 (N_2226,N_1937,N_1988);
nand U2227 (N_2227,N_1901,N_1940);
nor U2228 (N_2228,N_1854,N_1929);
and U2229 (N_2229,N_1937,N_1961);
nor U2230 (N_2230,N_1757,N_1810);
nand U2231 (N_2231,N_1800,N_1828);
xnor U2232 (N_2232,N_1760,N_1993);
or U2233 (N_2233,N_1904,N_1881);
or U2234 (N_2234,N_1781,N_1800);
nor U2235 (N_2235,N_1780,N_1995);
nand U2236 (N_2236,N_1915,N_1909);
nor U2237 (N_2237,N_1891,N_1857);
and U2238 (N_2238,N_1904,N_1809);
nand U2239 (N_2239,N_1867,N_1884);
and U2240 (N_2240,N_1957,N_1874);
and U2241 (N_2241,N_1849,N_1962);
nand U2242 (N_2242,N_1997,N_1951);
and U2243 (N_2243,N_1956,N_1810);
nand U2244 (N_2244,N_1782,N_1911);
and U2245 (N_2245,N_1799,N_1946);
or U2246 (N_2246,N_1999,N_1924);
nor U2247 (N_2247,N_1812,N_1933);
or U2248 (N_2248,N_1912,N_1765);
nand U2249 (N_2249,N_1991,N_1858);
and U2250 (N_2250,N_2066,N_2101);
or U2251 (N_2251,N_2238,N_2207);
xor U2252 (N_2252,N_2201,N_2085);
nor U2253 (N_2253,N_2186,N_2034);
or U2254 (N_2254,N_2022,N_2227);
or U2255 (N_2255,N_2188,N_2202);
or U2256 (N_2256,N_2082,N_2129);
and U2257 (N_2257,N_2136,N_2194);
and U2258 (N_2258,N_2065,N_2014);
nor U2259 (N_2259,N_2028,N_2067);
or U2260 (N_2260,N_2025,N_2209);
xnor U2261 (N_2261,N_2117,N_2193);
or U2262 (N_2262,N_2245,N_2061);
nor U2263 (N_2263,N_2051,N_2023);
nand U2264 (N_2264,N_2010,N_2153);
xnor U2265 (N_2265,N_2037,N_2174);
or U2266 (N_2266,N_2086,N_2070);
and U2267 (N_2267,N_2189,N_2103);
or U2268 (N_2268,N_2029,N_2217);
nand U2269 (N_2269,N_2011,N_2033);
and U2270 (N_2270,N_2096,N_2111);
or U2271 (N_2271,N_2246,N_2148);
and U2272 (N_2272,N_2050,N_2038);
or U2273 (N_2273,N_2046,N_2159);
or U2274 (N_2274,N_2183,N_2146);
nor U2275 (N_2275,N_2184,N_2178);
nand U2276 (N_2276,N_2237,N_2091);
and U2277 (N_2277,N_2035,N_2204);
or U2278 (N_2278,N_2080,N_2171);
nor U2279 (N_2279,N_2017,N_2230);
nor U2280 (N_2280,N_2241,N_2212);
and U2281 (N_2281,N_2208,N_2163);
nand U2282 (N_2282,N_2090,N_2100);
xor U2283 (N_2283,N_2239,N_2125);
nand U2284 (N_2284,N_2205,N_2141);
and U2285 (N_2285,N_2248,N_2223);
or U2286 (N_2286,N_2021,N_2197);
nand U2287 (N_2287,N_2057,N_2190);
or U2288 (N_2288,N_2001,N_2226);
and U2289 (N_2289,N_2095,N_2078);
or U2290 (N_2290,N_2094,N_2043);
or U2291 (N_2291,N_2048,N_2047);
nor U2292 (N_2292,N_2076,N_2236);
xnor U2293 (N_2293,N_2004,N_2191);
nand U2294 (N_2294,N_2087,N_2151);
nand U2295 (N_2295,N_2018,N_2147);
or U2296 (N_2296,N_2053,N_2064);
nor U2297 (N_2297,N_2114,N_2181);
nor U2298 (N_2298,N_2106,N_2072);
xor U2299 (N_2299,N_2030,N_2052);
nor U2300 (N_2300,N_2128,N_2122);
or U2301 (N_2301,N_2231,N_2016);
nand U2302 (N_2302,N_2112,N_2088);
nor U2303 (N_2303,N_2196,N_2131);
nand U2304 (N_2304,N_2039,N_2177);
and U2305 (N_2305,N_2124,N_2221);
nand U2306 (N_2306,N_2060,N_2150);
nor U2307 (N_2307,N_2247,N_2019);
nor U2308 (N_2308,N_2149,N_2195);
nor U2309 (N_2309,N_2092,N_2121);
nand U2310 (N_2310,N_2002,N_2249);
or U2311 (N_2311,N_2008,N_2135);
xor U2312 (N_2312,N_2185,N_2118);
nand U2313 (N_2313,N_2225,N_2099);
or U2314 (N_2314,N_2003,N_2026);
and U2315 (N_2315,N_2215,N_2134);
nor U2316 (N_2316,N_2055,N_2058);
and U2317 (N_2317,N_2044,N_2182);
nor U2318 (N_2318,N_2170,N_2127);
and U2319 (N_2319,N_2109,N_2213);
nor U2320 (N_2320,N_2219,N_2000);
or U2321 (N_2321,N_2007,N_2075);
nor U2322 (N_2322,N_2105,N_2126);
or U2323 (N_2323,N_2040,N_2045);
and U2324 (N_2324,N_2108,N_2027);
nand U2325 (N_2325,N_2123,N_2083);
nand U2326 (N_2326,N_2013,N_2012);
nor U2327 (N_2327,N_2168,N_2200);
nor U2328 (N_2328,N_2049,N_2119);
and U2329 (N_2329,N_2089,N_2240);
nand U2330 (N_2330,N_2180,N_2155);
nand U2331 (N_2331,N_2211,N_2113);
and U2332 (N_2332,N_2071,N_2132);
nand U2333 (N_2333,N_2224,N_2120);
and U2334 (N_2334,N_2152,N_2142);
or U2335 (N_2335,N_2074,N_2069);
and U2336 (N_2336,N_2220,N_2140);
nand U2337 (N_2337,N_2199,N_2005);
or U2338 (N_2338,N_2009,N_2102);
nand U2339 (N_2339,N_2166,N_2158);
nor U2340 (N_2340,N_2081,N_2218);
nor U2341 (N_2341,N_2203,N_2160);
nor U2342 (N_2342,N_2235,N_2244);
and U2343 (N_2343,N_2130,N_2156);
nand U2344 (N_2344,N_2192,N_2176);
nor U2345 (N_2345,N_2110,N_2042);
or U2346 (N_2346,N_2229,N_2165);
or U2347 (N_2347,N_2169,N_2115);
xor U2348 (N_2348,N_2198,N_2228);
or U2349 (N_2349,N_2162,N_2243);
and U2350 (N_2350,N_2161,N_2097);
nand U2351 (N_2351,N_2063,N_2098);
or U2352 (N_2352,N_2172,N_2222);
nand U2353 (N_2353,N_2242,N_2056);
nand U2354 (N_2354,N_2214,N_2167);
xor U2355 (N_2355,N_2145,N_2139);
and U2356 (N_2356,N_2006,N_2079);
and U2357 (N_2357,N_2206,N_2059);
xor U2358 (N_2358,N_2210,N_2233);
nor U2359 (N_2359,N_2187,N_2234);
and U2360 (N_2360,N_2144,N_2073);
and U2361 (N_2361,N_2133,N_2107);
nor U2362 (N_2362,N_2031,N_2032);
xnor U2363 (N_2363,N_2084,N_2093);
nand U2364 (N_2364,N_2179,N_2015);
or U2365 (N_2365,N_2054,N_2024);
and U2366 (N_2366,N_2068,N_2138);
and U2367 (N_2367,N_2216,N_2175);
or U2368 (N_2368,N_2157,N_2020);
nor U2369 (N_2369,N_2116,N_2232);
or U2370 (N_2370,N_2137,N_2173);
nor U2371 (N_2371,N_2041,N_2164);
nor U2372 (N_2372,N_2036,N_2077);
or U2373 (N_2373,N_2143,N_2154);
and U2374 (N_2374,N_2104,N_2062);
nand U2375 (N_2375,N_2030,N_2070);
or U2376 (N_2376,N_2218,N_2155);
or U2377 (N_2377,N_2118,N_2232);
nor U2378 (N_2378,N_2137,N_2193);
nand U2379 (N_2379,N_2064,N_2201);
and U2380 (N_2380,N_2101,N_2092);
nor U2381 (N_2381,N_2199,N_2081);
or U2382 (N_2382,N_2126,N_2012);
nand U2383 (N_2383,N_2198,N_2225);
or U2384 (N_2384,N_2247,N_2142);
or U2385 (N_2385,N_2175,N_2197);
nor U2386 (N_2386,N_2082,N_2069);
nor U2387 (N_2387,N_2242,N_2148);
xnor U2388 (N_2388,N_2170,N_2014);
nor U2389 (N_2389,N_2073,N_2045);
nand U2390 (N_2390,N_2214,N_2089);
nor U2391 (N_2391,N_2060,N_2110);
xnor U2392 (N_2392,N_2116,N_2061);
nand U2393 (N_2393,N_2115,N_2070);
and U2394 (N_2394,N_2023,N_2207);
nand U2395 (N_2395,N_2001,N_2125);
and U2396 (N_2396,N_2174,N_2077);
and U2397 (N_2397,N_2087,N_2023);
or U2398 (N_2398,N_2108,N_2177);
nor U2399 (N_2399,N_2033,N_2170);
xnor U2400 (N_2400,N_2230,N_2194);
nand U2401 (N_2401,N_2211,N_2168);
and U2402 (N_2402,N_2156,N_2226);
nand U2403 (N_2403,N_2171,N_2036);
nor U2404 (N_2404,N_2163,N_2070);
nand U2405 (N_2405,N_2045,N_2183);
nor U2406 (N_2406,N_2081,N_2125);
or U2407 (N_2407,N_2144,N_2142);
nor U2408 (N_2408,N_2150,N_2097);
and U2409 (N_2409,N_2164,N_2165);
and U2410 (N_2410,N_2140,N_2203);
or U2411 (N_2411,N_2077,N_2018);
nor U2412 (N_2412,N_2004,N_2100);
nand U2413 (N_2413,N_2033,N_2179);
and U2414 (N_2414,N_2184,N_2097);
nand U2415 (N_2415,N_2164,N_2169);
and U2416 (N_2416,N_2050,N_2195);
and U2417 (N_2417,N_2128,N_2115);
nor U2418 (N_2418,N_2182,N_2132);
or U2419 (N_2419,N_2103,N_2229);
or U2420 (N_2420,N_2017,N_2078);
and U2421 (N_2421,N_2053,N_2056);
and U2422 (N_2422,N_2026,N_2051);
or U2423 (N_2423,N_2187,N_2116);
nor U2424 (N_2424,N_2019,N_2162);
and U2425 (N_2425,N_2059,N_2172);
nand U2426 (N_2426,N_2162,N_2109);
and U2427 (N_2427,N_2033,N_2065);
nor U2428 (N_2428,N_2170,N_2178);
nand U2429 (N_2429,N_2158,N_2218);
nor U2430 (N_2430,N_2101,N_2000);
or U2431 (N_2431,N_2167,N_2012);
nand U2432 (N_2432,N_2185,N_2074);
and U2433 (N_2433,N_2182,N_2151);
or U2434 (N_2434,N_2172,N_2030);
nor U2435 (N_2435,N_2070,N_2020);
nand U2436 (N_2436,N_2003,N_2220);
and U2437 (N_2437,N_2013,N_2097);
or U2438 (N_2438,N_2104,N_2051);
and U2439 (N_2439,N_2118,N_2128);
nor U2440 (N_2440,N_2232,N_2007);
nor U2441 (N_2441,N_2094,N_2023);
and U2442 (N_2442,N_2248,N_2204);
xnor U2443 (N_2443,N_2056,N_2189);
or U2444 (N_2444,N_2109,N_2238);
and U2445 (N_2445,N_2056,N_2154);
or U2446 (N_2446,N_2209,N_2065);
or U2447 (N_2447,N_2126,N_2149);
nor U2448 (N_2448,N_2001,N_2168);
nand U2449 (N_2449,N_2030,N_2205);
or U2450 (N_2450,N_2238,N_2180);
nor U2451 (N_2451,N_2242,N_2243);
nand U2452 (N_2452,N_2069,N_2145);
nand U2453 (N_2453,N_2079,N_2148);
or U2454 (N_2454,N_2212,N_2033);
or U2455 (N_2455,N_2223,N_2042);
and U2456 (N_2456,N_2169,N_2042);
nor U2457 (N_2457,N_2175,N_2022);
nor U2458 (N_2458,N_2213,N_2157);
nand U2459 (N_2459,N_2177,N_2032);
xnor U2460 (N_2460,N_2102,N_2167);
nand U2461 (N_2461,N_2169,N_2215);
nor U2462 (N_2462,N_2083,N_2139);
or U2463 (N_2463,N_2034,N_2050);
and U2464 (N_2464,N_2030,N_2142);
nand U2465 (N_2465,N_2173,N_2054);
nand U2466 (N_2466,N_2014,N_2113);
nand U2467 (N_2467,N_2113,N_2009);
and U2468 (N_2468,N_2210,N_2246);
nand U2469 (N_2469,N_2082,N_2134);
nand U2470 (N_2470,N_2248,N_2171);
nand U2471 (N_2471,N_2026,N_2127);
and U2472 (N_2472,N_2094,N_2123);
or U2473 (N_2473,N_2002,N_2030);
nor U2474 (N_2474,N_2128,N_2249);
nor U2475 (N_2475,N_2074,N_2155);
and U2476 (N_2476,N_2212,N_2124);
or U2477 (N_2477,N_2154,N_2156);
or U2478 (N_2478,N_2244,N_2199);
or U2479 (N_2479,N_2108,N_2064);
nor U2480 (N_2480,N_2118,N_2062);
xor U2481 (N_2481,N_2068,N_2066);
nor U2482 (N_2482,N_2164,N_2087);
or U2483 (N_2483,N_2110,N_2231);
xnor U2484 (N_2484,N_2063,N_2121);
or U2485 (N_2485,N_2194,N_2203);
or U2486 (N_2486,N_2030,N_2019);
nand U2487 (N_2487,N_2165,N_2081);
nor U2488 (N_2488,N_2235,N_2068);
and U2489 (N_2489,N_2144,N_2015);
and U2490 (N_2490,N_2100,N_2040);
nor U2491 (N_2491,N_2067,N_2203);
or U2492 (N_2492,N_2121,N_2159);
nand U2493 (N_2493,N_2126,N_2004);
or U2494 (N_2494,N_2226,N_2040);
nor U2495 (N_2495,N_2175,N_2158);
nor U2496 (N_2496,N_2068,N_2012);
nand U2497 (N_2497,N_2173,N_2143);
xor U2498 (N_2498,N_2005,N_2196);
nor U2499 (N_2499,N_2053,N_2137);
or U2500 (N_2500,N_2321,N_2271);
and U2501 (N_2501,N_2297,N_2439);
or U2502 (N_2502,N_2442,N_2263);
or U2503 (N_2503,N_2307,N_2315);
nor U2504 (N_2504,N_2371,N_2281);
or U2505 (N_2505,N_2302,N_2454);
nor U2506 (N_2506,N_2483,N_2385);
nand U2507 (N_2507,N_2346,N_2438);
nand U2508 (N_2508,N_2251,N_2416);
or U2509 (N_2509,N_2389,N_2278);
nand U2510 (N_2510,N_2421,N_2407);
nand U2511 (N_2511,N_2490,N_2375);
and U2512 (N_2512,N_2434,N_2276);
nor U2513 (N_2513,N_2358,N_2482);
and U2514 (N_2514,N_2255,N_2456);
or U2515 (N_2515,N_2402,N_2425);
xnor U2516 (N_2516,N_2269,N_2467);
nor U2517 (N_2517,N_2461,N_2360);
xor U2518 (N_2518,N_2260,N_2447);
nor U2519 (N_2519,N_2440,N_2384);
nor U2520 (N_2520,N_2399,N_2361);
nand U2521 (N_2521,N_2418,N_2303);
and U2522 (N_2522,N_2353,N_2441);
or U2523 (N_2523,N_2462,N_2391);
nand U2524 (N_2524,N_2471,N_2277);
and U2525 (N_2525,N_2350,N_2436);
and U2526 (N_2526,N_2468,N_2465);
or U2527 (N_2527,N_2314,N_2422);
or U2528 (N_2528,N_2379,N_2400);
or U2529 (N_2529,N_2344,N_2295);
or U2530 (N_2530,N_2300,N_2347);
nor U2531 (N_2531,N_2287,N_2320);
and U2532 (N_2532,N_2362,N_2279);
nand U2533 (N_2533,N_2472,N_2444);
and U2534 (N_2534,N_2488,N_2481);
or U2535 (N_2535,N_2274,N_2426);
nand U2536 (N_2536,N_2448,N_2257);
or U2537 (N_2537,N_2337,N_2311);
and U2538 (N_2538,N_2417,N_2312);
nor U2539 (N_2539,N_2419,N_2394);
nand U2540 (N_2540,N_2405,N_2289);
nand U2541 (N_2541,N_2397,N_2477);
and U2542 (N_2542,N_2460,N_2290);
or U2543 (N_2543,N_2406,N_2395);
nor U2544 (N_2544,N_2497,N_2334);
nand U2545 (N_2545,N_2331,N_2386);
nor U2546 (N_2546,N_2363,N_2427);
nand U2547 (N_2547,N_2301,N_2259);
nand U2548 (N_2548,N_2415,N_2252);
nand U2549 (N_2549,N_2332,N_2273);
nand U2550 (N_2550,N_2306,N_2499);
and U2551 (N_2551,N_2487,N_2494);
and U2552 (N_2552,N_2285,N_2430);
or U2553 (N_2553,N_2359,N_2339);
nor U2554 (N_2554,N_2318,N_2414);
nand U2555 (N_2555,N_2390,N_2413);
xnor U2556 (N_2556,N_2366,N_2449);
nor U2557 (N_2557,N_2294,N_2403);
and U2558 (N_2558,N_2450,N_2495);
nor U2559 (N_2559,N_2378,N_2489);
and U2560 (N_2560,N_2412,N_2473);
nor U2561 (N_2561,N_2453,N_2451);
xnor U2562 (N_2562,N_2299,N_2475);
or U2563 (N_2563,N_2492,N_2280);
or U2564 (N_2564,N_2329,N_2420);
xor U2565 (N_2565,N_2404,N_2322);
and U2566 (N_2566,N_2335,N_2408);
nor U2567 (N_2567,N_2327,N_2478);
nand U2568 (N_2568,N_2387,N_2298);
nor U2569 (N_2569,N_2463,N_2310);
nand U2570 (N_2570,N_2382,N_2326);
xor U2571 (N_2571,N_2338,N_2459);
nor U2572 (N_2572,N_2372,N_2293);
and U2573 (N_2573,N_2357,N_2401);
or U2574 (N_2574,N_2484,N_2368);
xor U2575 (N_2575,N_2431,N_2396);
and U2576 (N_2576,N_2262,N_2275);
and U2577 (N_2577,N_2253,N_2340);
nor U2578 (N_2578,N_2429,N_2393);
nor U2579 (N_2579,N_2496,N_2474);
nand U2580 (N_2580,N_2345,N_2313);
or U2581 (N_2581,N_2486,N_2336);
or U2582 (N_2582,N_2261,N_2469);
nor U2583 (N_2583,N_2491,N_2466);
nor U2584 (N_2584,N_2352,N_2479);
and U2585 (N_2585,N_2342,N_2341);
nand U2586 (N_2586,N_2433,N_2268);
nand U2587 (N_2587,N_2284,N_2367);
nor U2588 (N_2588,N_2333,N_2376);
nor U2589 (N_2589,N_2258,N_2286);
and U2590 (N_2590,N_2288,N_2325);
nand U2591 (N_2591,N_2356,N_2354);
or U2592 (N_2592,N_2351,N_2270);
or U2593 (N_2593,N_2493,N_2296);
and U2594 (N_2594,N_2498,N_2381);
and U2595 (N_2595,N_2324,N_2377);
nand U2596 (N_2596,N_2316,N_2256);
nor U2597 (N_2597,N_2445,N_2343);
nand U2598 (N_2598,N_2374,N_2264);
nor U2599 (N_2599,N_2443,N_2452);
nand U2600 (N_2600,N_2317,N_2464);
nor U2601 (N_2601,N_2411,N_2364);
or U2602 (N_2602,N_2283,N_2458);
and U2603 (N_2603,N_2323,N_2485);
nand U2604 (N_2604,N_2410,N_2388);
nor U2605 (N_2605,N_2254,N_2328);
and U2606 (N_2606,N_2355,N_2250);
nand U2607 (N_2607,N_2432,N_2476);
xor U2608 (N_2608,N_2305,N_2282);
and U2609 (N_2609,N_2428,N_2424);
or U2610 (N_2610,N_2309,N_2266);
and U2611 (N_2611,N_2455,N_2267);
nand U2612 (N_2612,N_2291,N_2370);
nand U2613 (N_2613,N_2392,N_2348);
or U2614 (N_2614,N_2308,N_2437);
and U2615 (N_2615,N_2383,N_2265);
nor U2616 (N_2616,N_2480,N_2365);
nand U2617 (N_2617,N_2446,N_2435);
nor U2618 (N_2618,N_2470,N_2398);
nor U2619 (N_2619,N_2349,N_2319);
xor U2620 (N_2620,N_2292,N_2272);
nor U2621 (N_2621,N_2330,N_2304);
and U2622 (N_2622,N_2409,N_2380);
nor U2623 (N_2623,N_2369,N_2457);
and U2624 (N_2624,N_2373,N_2423);
nand U2625 (N_2625,N_2324,N_2250);
or U2626 (N_2626,N_2418,N_2470);
xor U2627 (N_2627,N_2296,N_2389);
nand U2628 (N_2628,N_2459,N_2272);
or U2629 (N_2629,N_2250,N_2409);
nand U2630 (N_2630,N_2260,N_2428);
and U2631 (N_2631,N_2260,N_2320);
and U2632 (N_2632,N_2366,N_2318);
nand U2633 (N_2633,N_2355,N_2339);
nand U2634 (N_2634,N_2400,N_2332);
or U2635 (N_2635,N_2465,N_2447);
or U2636 (N_2636,N_2473,N_2291);
nand U2637 (N_2637,N_2498,N_2447);
and U2638 (N_2638,N_2330,N_2274);
nor U2639 (N_2639,N_2268,N_2366);
xor U2640 (N_2640,N_2318,N_2341);
nand U2641 (N_2641,N_2388,N_2397);
or U2642 (N_2642,N_2464,N_2343);
xor U2643 (N_2643,N_2281,N_2295);
and U2644 (N_2644,N_2301,N_2337);
or U2645 (N_2645,N_2484,N_2489);
and U2646 (N_2646,N_2426,N_2302);
or U2647 (N_2647,N_2290,N_2394);
and U2648 (N_2648,N_2318,N_2413);
nand U2649 (N_2649,N_2481,N_2435);
or U2650 (N_2650,N_2324,N_2440);
and U2651 (N_2651,N_2322,N_2305);
nor U2652 (N_2652,N_2382,N_2279);
nor U2653 (N_2653,N_2471,N_2489);
nor U2654 (N_2654,N_2313,N_2470);
xor U2655 (N_2655,N_2471,N_2499);
and U2656 (N_2656,N_2317,N_2485);
or U2657 (N_2657,N_2284,N_2354);
nand U2658 (N_2658,N_2346,N_2293);
nor U2659 (N_2659,N_2387,N_2468);
nor U2660 (N_2660,N_2272,N_2481);
nor U2661 (N_2661,N_2355,N_2301);
xor U2662 (N_2662,N_2388,N_2295);
nor U2663 (N_2663,N_2389,N_2335);
and U2664 (N_2664,N_2279,N_2440);
nand U2665 (N_2665,N_2456,N_2400);
nand U2666 (N_2666,N_2385,N_2363);
nand U2667 (N_2667,N_2486,N_2333);
and U2668 (N_2668,N_2444,N_2284);
or U2669 (N_2669,N_2490,N_2382);
nor U2670 (N_2670,N_2369,N_2381);
and U2671 (N_2671,N_2493,N_2354);
or U2672 (N_2672,N_2365,N_2373);
nand U2673 (N_2673,N_2346,N_2491);
nor U2674 (N_2674,N_2366,N_2400);
xor U2675 (N_2675,N_2344,N_2262);
nand U2676 (N_2676,N_2295,N_2257);
or U2677 (N_2677,N_2496,N_2254);
and U2678 (N_2678,N_2310,N_2287);
and U2679 (N_2679,N_2251,N_2478);
nand U2680 (N_2680,N_2325,N_2418);
nand U2681 (N_2681,N_2319,N_2310);
and U2682 (N_2682,N_2470,N_2490);
xor U2683 (N_2683,N_2320,N_2468);
xor U2684 (N_2684,N_2285,N_2405);
xnor U2685 (N_2685,N_2488,N_2461);
or U2686 (N_2686,N_2458,N_2456);
and U2687 (N_2687,N_2391,N_2398);
nand U2688 (N_2688,N_2309,N_2469);
nand U2689 (N_2689,N_2428,N_2349);
nor U2690 (N_2690,N_2348,N_2318);
and U2691 (N_2691,N_2408,N_2478);
nand U2692 (N_2692,N_2413,N_2443);
nand U2693 (N_2693,N_2467,N_2288);
nor U2694 (N_2694,N_2313,N_2317);
and U2695 (N_2695,N_2286,N_2285);
nand U2696 (N_2696,N_2485,N_2313);
nor U2697 (N_2697,N_2276,N_2268);
and U2698 (N_2698,N_2250,N_2495);
and U2699 (N_2699,N_2340,N_2463);
nand U2700 (N_2700,N_2356,N_2308);
and U2701 (N_2701,N_2384,N_2255);
nand U2702 (N_2702,N_2337,N_2344);
nand U2703 (N_2703,N_2422,N_2441);
xor U2704 (N_2704,N_2368,N_2369);
nand U2705 (N_2705,N_2298,N_2349);
nor U2706 (N_2706,N_2321,N_2255);
and U2707 (N_2707,N_2351,N_2340);
nand U2708 (N_2708,N_2447,N_2364);
xnor U2709 (N_2709,N_2419,N_2475);
nor U2710 (N_2710,N_2496,N_2313);
nand U2711 (N_2711,N_2361,N_2352);
and U2712 (N_2712,N_2347,N_2342);
or U2713 (N_2713,N_2428,N_2419);
or U2714 (N_2714,N_2343,N_2495);
or U2715 (N_2715,N_2334,N_2338);
nand U2716 (N_2716,N_2427,N_2492);
xnor U2717 (N_2717,N_2277,N_2386);
and U2718 (N_2718,N_2282,N_2316);
or U2719 (N_2719,N_2415,N_2423);
xor U2720 (N_2720,N_2259,N_2319);
or U2721 (N_2721,N_2322,N_2340);
and U2722 (N_2722,N_2406,N_2383);
nand U2723 (N_2723,N_2310,N_2403);
nor U2724 (N_2724,N_2459,N_2495);
nor U2725 (N_2725,N_2365,N_2356);
nor U2726 (N_2726,N_2294,N_2475);
nand U2727 (N_2727,N_2338,N_2414);
nor U2728 (N_2728,N_2441,N_2321);
or U2729 (N_2729,N_2316,N_2383);
nand U2730 (N_2730,N_2346,N_2407);
nor U2731 (N_2731,N_2492,N_2394);
and U2732 (N_2732,N_2372,N_2329);
and U2733 (N_2733,N_2438,N_2444);
xnor U2734 (N_2734,N_2337,N_2378);
nor U2735 (N_2735,N_2260,N_2438);
and U2736 (N_2736,N_2260,N_2332);
nand U2737 (N_2737,N_2429,N_2484);
xor U2738 (N_2738,N_2443,N_2297);
and U2739 (N_2739,N_2408,N_2283);
and U2740 (N_2740,N_2329,N_2338);
or U2741 (N_2741,N_2394,N_2280);
nand U2742 (N_2742,N_2265,N_2481);
nand U2743 (N_2743,N_2405,N_2356);
nand U2744 (N_2744,N_2387,N_2406);
nand U2745 (N_2745,N_2493,N_2368);
nor U2746 (N_2746,N_2261,N_2316);
or U2747 (N_2747,N_2471,N_2334);
nand U2748 (N_2748,N_2359,N_2373);
nand U2749 (N_2749,N_2363,N_2412);
nor U2750 (N_2750,N_2655,N_2533);
and U2751 (N_2751,N_2541,N_2738);
and U2752 (N_2752,N_2685,N_2593);
xnor U2753 (N_2753,N_2604,N_2514);
and U2754 (N_2754,N_2729,N_2693);
and U2755 (N_2755,N_2575,N_2644);
xor U2756 (N_2756,N_2614,N_2612);
or U2757 (N_2757,N_2547,N_2714);
or U2758 (N_2758,N_2726,N_2699);
and U2759 (N_2759,N_2584,N_2734);
and U2760 (N_2760,N_2694,N_2641);
nand U2761 (N_2761,N_2717,N_2572);
or U2762 (N_2762,N_2608,N_2739);
and U2763 (N_2763,N_2585,N_2667);
xnor U2764 (N_2764,N_2646,N_2586);
xnor U2765 (N_2765,N_2559,N_2749);
nand U2766 (N_2766,N_2536,N_2510);
and U2767 (N_2767,N_2731,N_2682);
or U2768 (N_2768,N_2643,N_2532);
nand U2769 (N_2769,N_2562,N_2552);
nand U2770 (N_2770,N_2511,N_2660);
and U2771 (N_2771,N_2578,N_2635);
and U2772 (N_2772,N_2589,N_2550);
nor U2773 (N_2773,N_2709,N_2544);
nand U2774 (N_2774,N_2568,N_2623);
or U2775 (N_2775,N_2513,N_2560);
or U2776 (N_2776,N_2590,N_2565);
or U2777 (N_2777,N_2727,N_2733);
and U2778 (N_2778,N_2702,N_2705);
and U2779 (N_2779,N_2658,N_2588);
or U2780 (N_2780,N_2622,N_2645);
or U2781 (N_2781,N_2557,N_2665);
and U2782 (N_2782,N_2602,N_2615);
or U2783 (N_2783,N_2554,N_2583);
nand U2784 (N_2784,N_2521,N_2748);
or U2785 (N_2785,N_2689,N_2522);
xnor U2786 (N_2786,N_2553,N_2592);
nand U2787 (N_2787,N_2708,N_2524);
or U2788 (N_2788,N_2677,N_2692);
and U2789 (N_2789,N_2613,N_2549);
and U2790 (N_2790,N_2620,N_2636);
nand U2791 (N_2791,N_2728,N_2618);
or U2792 (N_2792,N_2698,N_2691);
and U2793 (N_2793,N_2642,N_2587);
and U2794 (N_2794,N_2629,N_2570);
or U2795 (N_2795,N_2741,N_2518);
and U2796 (N_2796,N_2519,N_2540);
xnor U2797 (N_2797,N_2504,N_2579);
nor U2798 (N_2798,N_2580,N_2680);
and U2799 (N_2799,N_2687,N_2581);
nor U2800 (N_2800,N_2515,N_2672);
nor U2801 (N_2801,N_2664,N_2747);
and U2802 (N_2802,N_2577,N_2516);
nand U2803 (N_2803,N_2526,N_2517);
or U2804 (N_2804,N_2656,N_2529);
or U2805 (N_2805,N_2610,N_2599);
and U2806 (N_2806,N_2663,N_2527);
nand U2807 (N_2807,N_2647,N_2649);
nand U2808 (N_2808,N_2505,N_2591);
xor U2809 (N_2809,N_2601,N_2670);
or U2810 (N_2810,N_2594,N_2648);
nor U2811 (N_2811,N_2697,N_2509);
and U2812 (N_2812,N_2528,N_2501);
nand U2813 (N_2813,N_2707,N_2523);
or U2814 (N_2814,N_2574,N_2722);
and U2815 (N_2815,N_2624,N_2661);
nor U2816 (N_2816,N_2743,N_2662);
and U2817 (N_2817,N_2546,N_2595);
and U2818 (N_2818,N_2531,N_2634);
nand U2819 (N_2819,N_2673,N_2558);
and U2820 (N_2820,N_2678,N_2628);
or U2821 (N_2821,N_2563,N_2617);
nor U2822 (N_2822,N_2545,N_2520);
nor U2823 (N_2823,N_2730,N_2639);
or U2824 (N_2824,N_2696,N_2569);
and U2825 (N_2825,N_2582,N_2551);
nand U2826 (N_2826,N_2571,N_2525);
xnor U2827 (N_2827,N_2711,N_2710);
xnor U2828 (N_2828,N_2605,N_2503);
nor U2829 (N_2829,N_2632,N_2745);
nor U2830 (N_2830,N_2506,N_2681);
nand U2831 (N_2831,N_2548,N_2671);
or U2832 (N_2832,N_2651,N_2742);
and U2833 (N_2833,N_2674,N_2659);
nand U2834 (N_2834,N_2626,N_2721);
and U2835 (N_2835,N_2735,N_2718);
nor U2836 (N_2836,N_2638,N_2744);
nor U2837 (N_2837,N_2537,N_2538);
or U2838 (N_2838,N_2668,N_2566);
nor U2839 (N_2839,N_2679,N_2627);
and U2840 (N_2840,N_2713,N_2561);
nor U2841 (N_2841,N_2573,N_2576);
nand U2842 (N_2842,N_2704,N_2686);
and U2843 (N_2843,N_2669,N_2640);
nor U2844 (N_2844,N_2684,N_2683);
nor U2845 (N_2845,N_2706,N_2597);
nand U2846 (N_2846,N_2596,N_2712);
nand U2847 (N_2847,N_2695,N_2690);
xnor U2848 (N_2848,N_2719,N_2736);
or U2849 (N_2849,N_2746,N_2534);
nor U2850 (N_2850,N_2621,N_2507);
nand U2851 (N_2851,N_2609,N_2542);
nand U2852 (N_2852,N_2688,N_2703);
nand U2853 (N_2853,N_2724,N_2567);
or U2854 (N_2854,N_2619,N_2723);
or U2855 (N_2855,N_2633,N_2631);
nor U2856 (N_2856,N_2676,N_2611);
xor U2857 (N_2857,N_2500,N_2539);
and U2858 (N_2858,N_2732,N_2637);
and U2859 (N_2859,N_2715,N_2543);
nand U2860 (N_2860,N_2555,N_2607);
xor U2861 (N_2861,N_2630,N_2616);
or U2862 (N_2862,N_2720,N_2508);
and U2863 (N_2863,N_2535,N_2654);
nor U2864 (N_2864,N_2603,N_2657);
nand U2865 (N_2865,N_2598,N_2512);
nand U2866 (N_2866,N_2700,N_2653);
nor U2867 (N_2867,N_2652,N_2606);
nand U2868 (N_2868,N_2737,N_2666);
and U2869 (N_2869,N_2530,N_2701);
nor U2870 (N_2870,N_2650,N_2740);
or U2871 (N_2871,N_2564,N_2625);
or U2872 (N_2872,N_2600,N_2675);
or U2873 (N_2873,N_2502,N_2716);
nand U2874 (N_2874,N_2556,N_2725);
xor U2875 (N_2875,N_2510,N_2625);
nor U2876 (N_2876,N_2542,N_2657);
or U2877 (N_2877,N_2709,N_2591);
nor U2878 (N_2878,N_2550,N_2617);
or U2879 (N_2879,N_2529,N_2672);
nand U2880 (N_2880,N_2653,N_2504);
nand U2881 (N_2881,N_2739,N_2632);
or U2882 (N_2882,N_2678,N_2573);
and U2883 (N_2883,N_2638,N_2515);
or U2884 (N_2884,N_2713,N_2719);
and U2885 (N_2885,N_2732,N_2682);
or U2886 (N_2886,N_2632,N_2543);
nor U2887 (N_2887,N_2550,N_2729);
nor U2888 (N_2888,N_2607,N_2649);
or U2889 (N_2889,N_2665,N_2700);
nor U2890 (N_2890,N_2661,N_2682);
nor U2891 (N_2891,N_2518,N_2598);
nor U2892 (N_2892,N_2700,N_2523);
nand U2893 (N_2893,N_2545,N_2701);
nor U2894 (N_2894,N_2607,N_2715);
xor U2895 (N_2895,N_2500,N_2732);
and U2896 (N_2896,N_2523,N_2618);
or U2897 (N_2897,N_2636,N_2584);
and U2898 (N_2898,N_2536,N_2526);
nor U2899 (N_2899,N_2574,N_2568);
nand U2900 (N_2900,N_2643,N_2718);
nor U2901 (N_2901,N_2642,N_2541);
nor U2902 (N_2902,N_2658,N_2702);
nand U2903 (N_2903,N_2591,N_2565);
xor U2904 (N_2904,N_2559,N_2692);
or U2905 (N_2905,N_2543,N_2608);
nand U2906 (N_2906,N_2654,N_2579);
nor U2907 (N_2907,N_2528,N_2723);
nor U2908 (N_2908,N_2684,N_2704);
nand U2909 (N_2909,N_2740,N_2512);
nor U2910 (N_2910,N_2679,N_2741);
or U2911 (N_2911,N_2706,N_2684);
and U2912 (N_2912,N_2503,N_2618);
nor U2913 (N_2913,N_2732,N_2712);
and U2914 (N_2914,N_2632,N_2533);
nand U2915 (N_2915,N_2716,N_2678);
or U2916 (N_2916,N_2658,N_2621);
nand U2917 (N_2917,N_2506,N_2605);
and U2918 (N_2918,N_2635,N_2706);
nor U2919 (N_2919,N_2523,N_2514);
and U2920 (N_2920,N_2730,N_2686);
and U2921 (N_2921,N_2547,N_2739);
nor U2922 (N_2922,N_2728,N_2704);
or U2923 (N_2923,N_2723,N_2541);
and U2924 (N_2924,N_2662,N_2514);
nand U2925 (N_2925,N_2564,N_2680);
nor U2926 (N_2926,N_2646,N_2706);
nand U2927 (N_2927,N_2532,N_2624);
or U2928 (N_2928,N_2597,N_2642);
nand U2929 (N_2929,N_2694,N_2718);
xor U2930 (N_2930,N_2670,N_2648);
nor U2931 (N_2931,N_2539,N_2672);
or U2932 (N_2932,N_2530,N_2567);
and U2933 (N_2933,N_2692,N_2574);
and U2934 (N_2934,N_2680,N_2618);
nor U2935 (N_2935,N_2576,N_2744);
nand U2936 (N_2936,N_2571,N_2711);
and U2937 (N_2937,N_2592,N_2680);
or U2938 (N_2938,N_2543,N_2549);
or U2939 (N_2939,N_2547,N_2519);
nand U2940 (N_2940,N_2537,N_2525);
and U2941 (N_2941,N_2587,N_2715);
nand U2942 (N_2942,N_2576,N_2524);
or U2943 (N_2943,N_2651,N_2559);
and U2944 (N_2944,N_2563,N_2530);
nand U2945 (N_2945,N_2624,N_2549);
and U2946 (N_2946,N_2731,N_2580);
nand U2947 (N_2947,N_2595,N_2696);
and U2948 (N_2948,N_2508,N_2569);
and U2949 (N_2949,N_2666,N_2545);
and U2950 (N_2950,N_2617,N_2663);
and U2951 (N_2951,N_2579,N_2577);
nor U2952 (N_2952,N_2649,N_2734);
and U2953 (N_2953,N_2507,N_2569);
nand U2954 (N_2954,N_2615,N_2732);
nand U2955 (N_2955,N_2507,N_2503);
and U2956 (N_2956,N_2695,N_2534);
nor U2957 (N_2957,N_2681,N_2547);
or U2958 (N_2958,N_2625,N_2574);
and U2959 (N_2959,N_2748,N_2588);
or U2960 (N_2960,N_2596,N_2622);
or U2961 (N_2961,N_2711,N_2522);
nand U2962 (N_2962,N_2539,N_2532);
nand U2963 (N_2963,N_2514,N_2728);
nand U2964 (N_2964,N_2564,N_2729);
nand U2965 (N_2965,N_2682,N_2720);
nor U2966 (N_2966,N_2694,N_2567);
or U2967 (N_2967,N_2746,N_2704);
xor U2968 (N_2968,N_2538,N_2540);
nand U2969 (N_2969,N_2615,N_2684);
xnor U2970 (N_2970,N_2749,N_2606);
nand U2971 (N_2971,N_2682,N_2536);
nand U2972 (N_2972,N_2678,N_2647);
and U2973 (N_2973,N_2606,N_2539);
or U2974 (N_2974,N_2530,N_2572);
xor U2975 (N_2975,N_2515,N_2514);
xor U2976 (N_2976,N_2651,N_2704);
or U2977 (N_2977,N_2601,N_2727);
nor U2978 (N_2978,N_2608,N_2564);
or U2979 (N_2979,N_2714,N_2502);
nand U2980 (N_2980,N_2687,N_2637);
or U2981 (N_2981,N_2587,N_2566);
and U2982 (N_2982,N_2570,N_2598);
and U2983 (N_2983,N_2611,N_2684);
nand U2984 (N_2984,N_2599,N_2511);
nor U2985 (N_2985,N_2607,N_2706);
and U2986 (N_2986,N_2710,N_2557);
or U2987 (N_2987,N_2670,N_2708);
nand U2988 (N_2988,N_2589,N_2612);
nand U2989 (N_2989,N_2545,N_2504);
nor U2990 (N_2990,N_2573,N_2721);
or U2991 (N_2991,N_2738,N_2514);
nand U2992 (N_2992,N_2730,N_2637);
or U2993 (N_2993,N_2660,N_2519);
or U2994 (N_2994,N_2694,N_2518);
nand U2995 (N_2995,N_2583,N_2630);
or U2996 (N_2996,N_2729,N_2705);
and U2997 (N_2997,N_2655,N_2652);
or U2998 (N_2998,N_2599,N_2749);
nor U2999 (N_2999,N_2630,N_2599);
or U3000 (N_3000,N_2869,N_2766);
nand U3001 (N_3001,N_2937,N_2752);
nand U3002 (N_3002,N_2870,N_2972);
and U3003 (N_3003,N_2979,N_2873);
or U3004 (N_3004,N_2864,N_2816);
and U3005 (N_3005,N_2913,N_2848);
nor U3006 (N_3006,N_2986,N_2973);
nand U3007 (N_3007,N_2838,N_2855);
and U3008 (N_3008,N_2961,N_2952);
and U3009 (N_3009,N_2755,N_2878);
or U3010 (N_3010,N_2910,N_2798);
nand U3011 (N_3011,N_2962,N_2888);
or U3012 (N_3012,N_2803,N_2750);
nand U3013 (N_3013,N_2835,N_2868);
xnor U3014 (N_3014,N_2851,N_2974);
and U3015 (N_3015,N_2906,N_2898);
nand U3016 (N_3016,N_2886,N_2753);
xnor U3017 (N_3017,N_2780,N_2783);
nor U3018 (N_3018,N_2762,N_2921);
or U3019 (N_3019,N_2936,N_2957);
nand U3020 (N_3020,N_2953,N_2925);
nand U3021 (N_3021,N_2944,N_2789);
nand U3022 (N_3022,N_2796,N_2949);
nand U3023 (N_3023,N_2996,N_2820);
nor U3024 (N_3024,N_2940,N_2993);
nor U3025 (N_3025,N_2779,N_2751);
xnor U3026 (N_3026,N_2861,N_2985);
or U3027 (N_3027,N_2824,N_2997);
nor U3028 (N_3028,N_2769,N_2988);
or U3029 (N_3029,N_2929,N_2982);
xnor U3030 (N_3030,N_2860,N_2811);
nor U3031 (N_3031,N_2915,N_2950);
and U3032 (N_3032,N_2806,N_2881);
or U3033 (N_3033,N_2884,N_2852);
or U3034 (N_3034,N_2939,N_2772);
nand U3035 (N_3035,N_2856,N_2989);
nor U3036 (N_3036,N_2760,N_2866);
or U3037 (N_3037,N_2920,N_2914);
or U3038 (N_3038,N_2872,N_2963);
nand U3039 (N_3039,N_2799,N_2976);
and U3040 (N_3040,N_2951,N_2904);
nor U3041 (N_3041,N_2823,N_2810);
or U3042 (N_3042,N_2923,N_2966);
and U3043 (N_3043,N_2825,N_2850);
nand U3044 (N_3044,N_2801,N_2858);
or U3045 (N_3045,N_2770,N_2968);
and U3046 (N_3046,N_2812,N_2773);
or U3047 (N_3047,N_2827,N_2896);
nor U3048 (N_3048,N_2882,N_2809);
and U3049 (N_3049,N_2894,N_2918);
nor U3050 (N_3050,N_2931,N_2756);
nor U3051 (N_3051,N_2943,N_2761);
nor U3052 (N_3052,N_2831,N_2849);
xnor U3053 (N_3053,N_2828,N_2900);
nor U3054 (N_3054,N_2916,N_2836);
nor U3055 (N_3055,N_2768,N_2975);
nor U3056 (N_3056,N_2792,N_2908);
nor U3057 (N_3057,N_2984,N_2797);
or U3058 (N_3058,N_2948,N_2905);
and U3059 (N_3059,N_2774,N_2790);
nor U3060 (N_3060,N_2782,N_2965);
or U3061 (N_3061,N_2771,N_2793);
nor U3062 (N_3062,N_2917,N_2967);
or U3063 (N_3063,N_2791,N_2947);
nor U3064 (N_3064,N_2969,N_2839);
or U3065 (N_3065,N_2991,N_2871);
xnor U3066 (N_3066,N_2874,N_2909);
nor U3067 (N_3067,N_2822,N_2837);
nor U3068 (N_3068,N_2971,N_2814);
and U3069 (N_3069,N_2958,N_2880);
nand U3070 (N_3070,N_2767,N_2844);
nor U3071 (N_3071,N_2758,N_2785);
and U3072 (N_3072,N_2899,N_2826);
or U3073 (N_3073,N_2890,N_2926);
nor U3074 (N_3074,N_2875,N_2912);
or U3075 (N_3075,N_2842,N_2887);
nor U3076 (N_3076,N_2841,N_2757);
xor U3077 (N_3077,N_2981,N_2955);
or U3078 (N_3078,N_2935,N_2843);
and U3079 (N_3079,N_2859,N_2922);
nand U3080 (N_3080,N_2832,N_2932);
nand U3081 (N_3081,N_2795,N_2754);
nor U3082 (N_3082,N_2863,N_2765);
nor U3083 (N_3083,N_2777,N_2802);
or U3084 (N_3084,N_2857,N_2960);
xnor U3085 (N_3085,N_2891,N_2885);
and U3086 (N_3086,N_2794,N_2964);
or U3087 (N_3087,N_2845,N_2992);
nor U3088 (N_3088,N_2883,N_2980);
nor U3089 (N_3089,N_2867,N_2786);
nand U3090 (N_3090,N_2897,N_2805);
nor U3091 (N_3091,N_2903,N_2759);
nand U3092 (N_3092,N_2817,N_2959);
nor U3093 (N_3093,N_2854,N_2876);
and U3094 (N_3094,N_2800,N_2763);
and U3095 (N_3095,N_2804,N_2933);
nand U3096 (N_3096,N_2840,N_2987);
nand U3097 (N_3097,N_2781,N_2977);
and U3098 (N_3098,N_2778,N_2990);
nand U3099 (N_3099,N_2998,N_2877);
and U3100 (N_3100,N_2927,N_2893);
or U3101 (N_3101,N_2787,N_2919);
nand U3102 (N_3102,N_2970,N_2846);
nor U3103 (N_3103,N_2930,N_2853);
and U3104 (N_3104,N_2928,N_2829);
nand U3105 (N_3105,N_2821,N_2946);
nor U3106 (N_3106,N_2924,N_2945);
xnor U3107 (N_3107,N_2954,N_2819);
or U3108 (N_3108,N_2995,N_2775);
nor U3109 (N_3109,N_2983,N_2895);
or U3110 (N_3110,N_2911,N_2808);
and U3111 (N_3111,N_2941,N_2815);
or U3112 (N_3112,N_2813,N_2834);
and U3113 (N_3113,N_2999,N_2902);
or U3114 (N_3114,N_2784,N_2788);
nor U3115 (N_3115,N_2978,N_2830);
nand U3116 (N_3116,N_2934,N_2889);
and U3117 (N_3117,N_2879,N_2956);
xnor U3118 (N_3118,N_2807,N_2892);
or U3119 (N_3119,N_2907,N_2818);
nor U3120 (N_3120,N_2862,N_2942);
nand U3121 (N_3121,N_2833,N_2764);
and U3122 (N_3122,N_2901,N_2938);
nor U3123 (N_3123,N_2865,N_2847);
and U3124 (N_3124,N_2994,N_2776);
nand U3125 (N_3125,N_2772,N_2998);
xor U3126 (N_3126,N_2907,N_2795);
and U3127 (N_3127,N_2794,N_2770);
nor U3128 (N_3128,N_2947,N_2978);
nor U3129 (N_3129,N_2897,N_2784);
nor U3130 (N_3130,N_2891,N_2864);
nand U3131 (N_3131,N_2774,N_2934);
nor U3132 (N_3132,N_2903,N_2970);
and U3133 (N_3133,N_2828,N_2764);
xnor U3134 (N_3134,N_2764,N_2768);
nand U3135 (N_3135,N_2833,N_2934);
nand U3136 (N_3136,N_2836,N_2883);
nand U3137 (N_3137,N_2967,N_2913);
or U3138 (N_3138,N_2833,N_2780);
nand U3139 (N_3139,N_2773,N_2870);
or U3140 (N_3140,N_2862,N_2829);
and U3141 (N_3141,N_2926,N_2873);
nand U3142 (N_3142,N_2917,N_2982);
and U3143 (N_3143,N_2983,N_2996);
and U3144 (N_3144,N_2770,N_2791);
nand U3145 (N_3145,N_2752,N_2873);
and U3146 (N_3146,N_2798,N_2882);
nand U3147 (N_3147,N_2957,N_2828);
nand U3148 (N_3148,N_2818,N_2910);
or U3149 (N_3149,N_2954,N_2804);
nor U3150 (N_3150,N_2797,N_2953);
nor U3151 (N_3151,N_2773,N_2892);
nand U3152 (N_3152,N_2916,N_2766);
xnor U3153 (N_3153,N_2851,N_2970);
or U3154 (N_3154,N_2925,N_2915);
or U3155 (N_3155,N_2911,N_2758);
nor U3156 (N_3156,N_2858,N_2852);
and U3157 (N_3157,N_2907,N_2886);
nand U3158 (N_3158,N_2903,N_2910);
or U3159 (N_3159,N_2963,N_2937);
xnor U3160 (N_3160,N_2952,N_2832);
or U3161 (N_3161,N_2770,N_2797);
or U3162 (N_3162,N_2964,N_2856);
nand U3163 (N_3163,N_2970,N_2777);
or U3164 (N_3164,N_2812,N_2788);
or U3165 (N_3165,N_2928,N_2813);
xor U3166 (N_3166,N_2899,N_2766);
nor U3167 (N_3167,N_2977,N_2793);
xor U3168 (N_3168,N_2828,N_2887);
and U3169 (N_3169,N_2992,N_2756);
xnor U3170 (N_3170,N_2946,N_2779);
nand U3171 (N_3171,N_2782,N_2937);
nand U3172 (N_3172,N_2960,N_2786);
or U3173 (N_3173,N_2841,N_2984);
nand U3174 (N_3174,N_2984,N_2753);
nand U3175 (N_3175,N_2766,N_2873);
nand U3176 (N_3176,N_2885,N_2844);
and U3177 (N_3177,N_2837,N_2978);
nand U3178 (N_3178,N_2876,N_2859);
nor U3179 (N_3179,N_2866,N_2995);
nand U3180 (N_3180,N_2838,N_2754);
nand U3181 (N_3181,N_2814,N_2837);
nor U3182 (N_3182,N_2851,N_2788);
nor U3183 (N_3183,N_2842,N_2964);
and U3184 (N_3184,N_2900,N_2824);
or U3185 (N_3185,N_2799,N_2977);
nor U3186 (N_3186,N_2875,N_2986);
or U3187 (N_3187,N_2958,N_2859);
and U3188 (N_3188,N_2871,N_2947);
and U3189 (N_3189,N_2773,N_2973);
nor U3190 (N_3190,N_2756,N_2927);
nor U3191 (N_3191,N_2880,N_2927);
or U3192 (N_3192,N_2799,N_2870);
and U3193 (N_3193,N_2904,N_2935);
and U3194 (N_3194,N_2860,N_2859);
or U3195 (N_3195,N_2900,N_2982);
and U3196 (N_3196,N_2839,N_2780);
nand U3197 (N_3197,N_2769,N_2851);
nand U3198 (N_3198,N_2961,N_2814);
or U3199 (N_3199,N_2988,N_2806);
and U3200 (N_3200,N_2879,N_2767);
and U3201 (N_3201,N_2903,N_2911);
or U3202 (N_3202,N_2849,N_2873);
or U3203 (N_3203,N_2989,N_2819);
or U3204 (N_3204,N_2844,N_2854);
and U3205 (N_3205,N_2997,N_2818);
nand U3206 (N_3206,N_2762,N_2972);
or U3207 (N_3207,N_2810,N_2830);
nand U3208 (N_3208,N_2929,N_2834);
nor U3209 (N_3209,N_2863,N_2819);
nand U3210 (N_3210,N_2902,N_2963);
or U3211 (N_3211,N_2808,N_2790);
nor U3212 (N_3212,N_2846,N_2792);
nand U3213 (N_3213,N_2907,N_2924);
or U3214 (N_3214,N_2993,N_2768);
nand U3215 (N_3215,N_2995,N_2985);
or U3216 (N_3216,N_2826,N_2767);
or U3217 (N_3217,N_2768,N_2931);
nand U3218 (N_3218,N_2873,N_2974);
and U3219 (N_3219,N_2770,N_2890);
nor U3220 (N_3220,N_2846,N_2853);
and U3221 (N_3221,N_2817,N_2900);
xnor U3222 (N_3222,N_2943,N_2824);
and U3223 (N_3223,N_2854,N_2953);
nor U3224 (N_3224,N_2947,N_2815);
nor U3225 (N_3225,N_2783,N_2857);
nand U3226 (N_3226,N_2951,N_2983);
xor U3227 (N_3227,N_2925,N_2870);
nand U3228 (N_3228,N_2877,N_2885);
xnor U3229 (N_3229,N_2801,N_2897);
nand U3230 (N_3230,N_2866,N_2816);
or U3231 (N_3231,N_2948,N_2886);
and U3232 (N_3232,N_2866,N_2847);
and U3233 (N_3233,N_2922,N_2998);
and U3234 (N_3234,N_2942,N_2915);
and U3235 (N_3235,N_2974,N_2794);
nor U3236 (N_3236,N_2813,N_2800);
nand U3237 (N_3237,N_2842,N_2943);
or U3238 (N_3238,N_2885,N_2775);
and U3239 (N_3239,N_2817,N_2884);
nand U3240 (N_3240,N_2974,N_2930);
xor U3241 (N_3241,N_2882,N_2933);
xnor U3242 (N_3242,N_2975,N_2859);
nand U3243 (N_3243,N_2954,N_2880);
nor U3244 (N_3244,N_2955,N_2971);
nor U3245 (N_3245,N_2785,N_2794);
nand U3246 (N_3246,N_2926,N_2921);
nor U3247 (N_3247,N_2908,N_2866);
and U3248 (N_3248,N_2797,N_2909);
or U3249 (N_3249,N_2896,N_2964);
nor U3250 (N_3250,N_3074,N_3150);
or U3251 (N_3251,N_3008,N_3036);
nor U3252 (N_3252,N_3088,N_3192);
or U3253 (N_3253,N_3232,N_3046);
nor U3254 (N_3254,N_3238,N_3098);
xnor U3255 (N_3255,N_3018,N_3083);
and U3256 (N_3256,N_3109,N_3133);
nor U3257 (N_3257,N_3168,N_3114);
or U3258 (N_3258,N_3241,N_3171);
and U3259 (N_3259,N_3089,N_3041);
nand U3260 (N_3260,N_3182,N_3155);
or U3261 (N_3261,N_3131,N_3203);
nand U3262 (N_3262,N_3196,N_3124);
and U3263 (N_3263,N_3009,N_3006);
nor U3264 (N_3264,N_3211,N_3186);
nor U3265 (N_3265,N_3123,N_3176);
and U3266 (N_3266,N_3095,N_3043);
or U3267 (N_3267,N_3126,N_3161);
and U3268 (N_3268,N_3027,N_3197);
nor U3269 (N_3269,N_3082,N_3184);
and U3270 (N_3270,N_3115,N_3188);
or U3271 (N_3271,N_3069,N_3075);
nor U3272 (N_3272,N_3227,N_3142);
nor U3273 (N_3273,N_3042,N_3034);
nand U3274 (N_3274,N_3217,N_3084);
and U3275 (N_3275,N_3249,N_3038);
xor U3276 (N_3276,N_3064,N_3050);
nor U3277 (N_3277,N_3057,N_3121);
nand U3278 (N_3278,N_3056,N_3230);
nor U3279 (N_3279,N_3097,N_3245);
xor U3280 (N_3280,N_3206,N_3180);
nand U3281 (N_3281,N_3116,N_3012);
and U3282 (N_3282,N_3086,N_3135);
nor U3283 (N_3283,N_3237,N_3139);
or U3284 (N_3284,N_3029,N_3146);
nor U3285 (N_3285,N_3159,N_3017);
and U3286 (N_3286,N_3165,N_3215);
or U3287 (N_3287,N_3066,N_3059);
or U3288 (N_3288,N_3175,N_3226);
xor U3289 (N_3289,N_3191,N_3201);
nand U3290 (N_3290,N_3242,N_3080);
nand U3291 (N_3291,N_3070,N_3032);
nand U3292 (N_3292,N_3223,N_3187);
nor U3293 (N_3293,N_3147,N_3216);
nor U3294 (N_3294,N_3235,N_3140);
nor U3295 (N_3295,N_3096,N_3243);
nand U3296 (N_3296,N_3119,N_3212);
nor U3297 (N_3297,N_3055,N_3170);
or U3298 (N_3298,N_3222,N_3156);
nor U3299 (N_3299,N_3033,N_3177);
nor U3300 (N_3300,N_3007,N_3094);
nor U3301 (N_3301,N_3127,N_3077);
nor U3302 (N_3302,N_3103,N_3058);
or U3303 (N_3303,N_3138,N_3051);
xor U3304 (N_3304,N_3221,N_3193);
nand U3305 (N_3305,N_3183,N_3048);
nand U3306 (N_3306,N_3053,N_3002);
nand U3307 (N_3307,N_3153,N_3169);
nand U3308 (N_3308,N_3072,N_3167);
or U3309 (N_3309,N_3151,N_3166);
or U3310 (N_3310,N_3076,N_3093);
or U3311 (N_3311,N_3078,N_3229);
nand U3312 (N_3312,N_3125,N_3154);
nand U3313 (N_3313,N_3035,N_3195);
nor U3314 (N_3314,N_3107,N_3039);
and U3315 (N_3315,N_3218,N_3157);
nor U3316 (N_3316,N_3152,N_3202);
nor U3317 (N_3317,N_3079,N_3248);
or U3318 (N_3318,N_3025,N_3073);
nand U3319 (N_3319,N_3105,N_3129);
or U3320 (N_3320,N_3185,N_3200);
nand U3321 (N_3321,N_3141,N_3021);
nand U3322 (N_3322,N_3011,N_3030);
or U3323 (N_3323,N_3108,N_3052);
nor U3324 (N_3324,N_3020,N_3205);
and U3325 (N_3325,N_3061,N_3204);
nor U3326 (N_3326,N_3194,N_3010);
and U3327 (N_3327,N_3054,N_3143);
nand U3328 (N_3328,N_3209,N_3110);
and U3329 (N_3329,N_3019,N_3149);
nand U3330 (N_3330,N_3130,N_3160);
nor U3331 (N_3331,N_3207,N_3090);
and U3332 (N_3332,N_3028,N_3220);
nor U3333 (N_3333,N_3111,N_3162);
or U3334 (N_3334,N_3172,N_3190);
nor U3335 (N_3335,N_3100,N_3247);
nor U3336 (N_3336,N_3225,N_3113);
or U3337 (N_3337,N_3179,N_3022);
nand U3338 (N_3338,N_3091,N_3219);
and U3339 (N_3339,N_3174,N_3210);
xor U3340 (N_3340,N_3047,N_3016);
and U3341 (N_3341,N_3137,N_3037);
nor U3342 (N_3342,N_3044,N_3236);
xor U3343 (N_3343,N_3181,N_3013);
nand U3344 (N_3344,N_3234,N_3087);
and U3345 (N_3345,N_3060,N_3213);
and U3346 (N_3346,N_3112,N_3004);
xnor U3347 (N_3347,N_3132,N_3023);
or U3348 (N_3348,N_3228,N_3118);
nand U3349 (N_3349,N_3063,N_3101);
or U3350 (N_3350,N_3214,N_3068);
or U3351 (N_3351,N_3085,N_3040);
nand U3352 (N_3352,N_3244,N_3233);
nor U3353 (N_3353,N_3099,N_3065);
or U3354 (N_3354,N_3158,N_3198);
xnor U3355 (N_3355,N_3128,N_3024);
nand U3356 (N_3356,N_3173,N_3120);
xnor U3357 (N_3357,N_3231,N_3026);
xnor U3358 (N_3358,N_3062,N_3145);
or U3359 (N_3359,N_3208,N_3163);
or U3360 (N_3360,N_3106,N_3067);
nor U3361 (N_3361,N_3000,N_3102);
or U3362 (N_3362,N_3117,N_3240);
nor U3363 (N_3363,N_3164,N_3092);
or U3364 (N_3364,N_3134,N_3014);
or U3365 (N_3365,N_3049,N_3189);
and U3366 (N_3366,N_3122,N_3144);
nand U3367 (N_3367,N_3001,N_3199);
xor U3368 (N_3368,N_3246,N_3015);
nor U3369 (N_3369,N_3071,N_3045);
and U3370 (N_3370,N_3224,N_3136);
or U3371 (N_3371,N_3239,N_3104);
and U3372 (N_3372,N_3178,N_3005);
and U3373 (N_3373,N_3003,N_3081);
nor U3374 (N_3374,N_3031,N_3148);
or U3375 (N_3375,N_3017,N_3019);
nor U3376 (N_3376,N_3191,N_3102);
xnor U3377 (N_3377,N_3145,N_3022);
xor U3378 (N_3378,N_3032,N_3054);
nor U3379 (N_3379,N_3017,N_3238);
nor U3380 (N_3380,N_3167,N_3186);
or U3381 (N_3381,N_3151,N_3056);
and U3382 (N_3382,N_3212,N_3040);
nand U3383 (N_3383,N_3071,N_3008);
and U3384 (N_3384,N_3043,N_3126);
and U3385 (N_3385,N_3038,N_3024);
nor U3386 (N_3386,N_3221,N_3235);
nand U3387 (N_3387,N_3246,N_3232);
and U3388 (N_3388,N_3216,N_3178);
nor U3389 (N_3389,N_3232,N_3132);
nand U3390 (N_3390,N_3209,N_3177);
and U3391 (N_3391,N_3204,N_3123);
and U3392 (N_3392,N_3197,N_3035);
nor U3393 (N_3393,N_3060,N_3184);
nor U3394 (N_3394,N_3052,N_3082);
and U3395 (N_3395,N_3229,N_3115);
nand U3396 (N_3396,N_3223,N_3115);
xnor U3397 (N_3397,N_3032,N_3116);
or U3398 (N_3398,N_3002,N_3174);
xnor U3399 (N_3399,N_3094,N_3058);
xnor U3400 (N_3400,N_3211,N_3024);
nor U3401 (N_3401,N_3051,N_3066);
or U3402 (N_3402,N_3119,N_3180);
nand U3403 (N_3403,N_3185,N_3032);
and U3404 (N_3404,N_3230,N_3020);
xnor U3405 (N_3405,N_3052,N_3206);
or U3406 (N_3406,N_3105,N_3094);
and U3407 (N_3407,N_3115,N_3237);
and U3408 (N_3408,N_3151,N_3101);
xnor U3409 (N_3409,N_3009,N_3016);
and U3410 (N_3410,N_3069,N_3219);
nand U3411 (N_3411,N_3120,N_3109);
xor U3412 (N_3412,N_3089,N_3108);
or U3413 (N_3413,N_3092,N_3237);
xor U3414 (N_3414,N_3111,N_3046);
and U3415 (N_3415,N_3246,N_3223);
or U3416 (N_3416,N_3184,N_3033);
nor U3417 (N_3417,N_3007,N_3194);
nand U3418 (N_3418,N_3106,N_3022);
or U3419 (N_3419,N_3067,N_3120);
xnor U3420 (N_3420,N_3043,N_3114);
nand U3421 (N_3421,N_3022,N_3092);
or U3422 (N_3422,N_3224,N_3130);
xor U3423 (N_3423,N_3133,N_3025);
nor U3424 (N_3424,N_3064,N_3128);
nand U3425 (N_3425,N_3226,N_3124);
or U3426 (N_3426,N_3037,N_3080);
and U3427 (N_3427,N_3133,N_3028);
xnor U3428 (N_3428,N_3056,N_3215);
nor U3429 (N_3429,N_3040,N_3216);
nand U3430 (N_3430,N_3223,N_3225);
nand U3431 (N_3431,N_3089,N_3198);
xnor U3432 (N_3432,N_3091,N_3181);
nand U3433 (N_3433,N_3193,N_3184);
or U3434 (N_3434,N_3056,N_3039);
nor U3435 (N_3435,N_3216,N_3017);
or U3436 (N_3436,N_3088,N_3027);
and U3437 (N_3437,N_3177,N_3039);
nor U3438 (N_3438,N_3055,N_3127);
xor U3439 (N_3439,N_3056,N_3224);
and U3440 (N_3440,N_3038,N_3070);
nand U3441 (N_3441,N_3148,N_3059);
xnor U3442 (N_3442,N_3185,N_3158);
nand U3443 (N_3443,N_3176,N_3213);
xor U3444 (N_3444,N_3226,N_3068);
nor U3445 (N_3445,N_3148,N_3245);
nand U3446 (N_3446,N_3157,N_3174);
and U3447 (N_3447,N_3098,N_3232);
or U3448 (N_3448,N_3021,N_3046);
nor U3449 (N_3449,N_3149,N_3177);
xnor U3450 (N_3450,N_3167,N_3240);
nand U3451 (N_3451,N_3232,N_3153);
and U3452 (N_3452,N_3107,N_3016);
nor U3453 (N_3453,N_3033,N_3189);
or U3454 (N_3454,N_3207,N_3123);
nor U3455 (N_3455,N_3073,N_3156);
nor U3456 (N_3456,N_3118,N_3009);
or U3457 (N_3457,N_3018,N_3084);
and U3458 (N_3458,N_3050,N_3226);
nand U3459 (N_3459,N_3106,N_3026);
or U3460 (N_3460,N_3129,N_3157);
nor U3461 (N_3461,N_3118,N_3044);
xnor U3462 (N_3462,N_3149,N_3219);
nand U3463 (N_3463,N_3150,N_3236);
or U3464 (N_3464,N_3079,N_3016);
and U3465 (N_3465,N_3151,N_3161);
and U3466 (N_3466,N_3083,N_3161);
or U3467 (N_3467,N_3129,N_3192);
or U3468 (N_3468,N_3092,N_3234);
or U3469 (N_3469,N_3107,N_3015);
or U3470 (N_3470,N_3052,N_3012);
nand U3471 (N_3471,N_3123,N_3177);
xnor U3472 (N_3472,N_3023,N_3082);
nor U3473 (N_3473,N_3139,N_3010);
or U3474 (N_3474,N_3051,N_3199);
and U3475 (N_3475,N_3229,N_3061);
or U3476 (N_3476,N_3220,N_3137);
nand U3477 (N_3477,N_3134,N_3119);
nor U3478 (N_3478,N_3055,N_3209);
nand U3479 (N_3479,N_3191,N_3235);
nor U3480 (N_3480,N_3115,N_3152);
nor U3481 (N_3481,N_3181,N_3216);
and U3482 (N_3482,N_3183,N_3152);
and U3483 (N_3483,N_3093,N_3081);
nand U3484 (N_3484,N_3026,N_3050);
nand U3485 (N_3485,N_3148,N_3208);
or U3486 (N_3486,N_3188,N_3099);
or U3487 (N_3487,N_3119,N_3012);
or U3488 (N_3488,N_3032,N_3154);
nor U3489 (N_3489,N_3214,N_3200);
nor U3490 (N_3490,N_3051,N_3149);
and U3491 (N_3491,N_3178,N_3166);
nor U3492 (N_3492,N_3158,N_3197);
nand U3493 (N_3493,N_3184,N_3079);
and U3494 (N_3494,N_3118,N_3091);
nand U3495 (N_3495,N_3131,N_3149);
nand U3496 (N_3496,N_3211,N_3041);
xnor U3497 (N_3497,N_3189,N_3239);
and U3498 (N_3498,N_3241,N_3041);
and U3499 (N_3499,N_3152,N_3194);
nand U3500 (N_3500,N_3381,N_3366);
or U3501 (N_3501,N_3490,N_3299);
and U3502 (N_3502,N_3474,N_3318);
nand U3503 (N_3503,N_3413,N_3497);
and U3504 (N_3504,N_3275,N_3287);
xor U3505 (N_3505,N_3444,N_3423);
nor U3506 (N_3506,N_3254,N_3262);
nor U3507 (N_3507,N_3293,N_3315);
and U3508 (N_3508,N_3492,N_3274);
nor U3509 (N_3509,N_3377,N_3445);
or U3510 (N_3510,N_3295,N_3402);
nand U3511 (N_3511,N_3464,N_3322);
or U3512 (N_3512,N_3371,N_3364);
nor U3513 (N_3513,N_3498,N_3272);
nor U3514 (N_3514,N_3278,N_3338);
and U3515 (N_3515,N_3294,N_3326);
nor U3516 (N_3516,N_3394,N_3325);
and U3517 (N_3517,N_3431,N_3347);
nand U3518 (N_3518,N_3283,N_3449);
or U3519 (N_3519,N_3340,N_3428);
xnor U3520 (N_3520,N_3432,N_3410);
nor U3521 (N_3521,N_3436,N_3470);
and U3522 (N_3522,N_3267,N_3403);
xor U3523 (N_3523,N_3344,N_3456);
nand U3524 (N_3524,N_3312,N_3458);
and U3525 (N_3525,N_3300,N_3285);
nor U3526 (N_3526,N_3466,N_3425);
nand U3527 (N_3527,N_3407,N_3361);
or U3528 (N_3528,N_3412,N_3332);
or U3529 (N_3529,N_3487,N_3405);
or U3530 (N_3530,N_3307,N_3457);
xnor U3531 (N_3531,N_3292,N_3453);
or U3532 (N_3532,N_3454,N_3303);
or U3533 (N_3533,N_3400,N_3393);
xor U3534 (N_3534,N_3495,N_3319);
xnor U3535 (N_3535,N_3380,N_3341);
or U3536 (N_3536,N_3335,N_3424);
nand U3537 (N_3537,N_3486,N_3485);
nand U3538 (N_3538,N_3468,N_3313);
and U3539 (N_3539,N_3404,N_3376);
and U3540 (N_3540,N_3258,N_3397);
or U3541 (N_3541,N_3308,N_3346);
and U3542 (N_3542,N_3416,N_3280);
nand U3543 (N_3543,N_3396,N_3320);
nor U3544 (N_3544,N_3460,N_3337);
nor U3545 (N_3545,N_3391,N_3336);
or U3546 (N_3546,N_3384,N_3378);
and U3547 (N_3547,N_3309,N_3443);
or U3548 (N_3548,N_3417,N_3450);
nor U3549 (N_3549,N_3289,N_3465);
nand U3550 (N_3550,N_3469,N_3399);
and U3551 (N_3551,N_3351,N_3379);
xor U3552 (N_3552,N_3284,N_3477);
and U3553 (N_3553,N_3479,N_3388);
xnor U3554 (N_3554,N_3448,N_3463);
and U3555 (N_3555,N_3296,N_3355);
nand U3556 (N_3556,N_3250,N_3348);
nand U3557 (N_3557,N_3433,N_3323);
nor U3558 (N_3558,N_3499,N_3387);
nand U3559 (N_3559,N_3421,N_3451);
nand U3560 (N_3560,N_3420,N_3252);
nand U3561 (N_3561,N_3447,N_3398);
or U3562 (N_3562,N_3392,N_3491);
nand U3563 (N_3563,N_3365,N_3430);
nor U3564 (N_3564,N_3476,N_3268);
or U3565 (N_3565,N_3418,N_3304);
nand U3566 (N_3566,N_3419,N_3415);
xnor U3567 (N_3567,N_3406,N_3298);
or U3568 (N_3568,N_3343,N_3368);
nor U3569 (N_3569,N_3459,N_3281);
nor U3570 (N_3570,N_3302,N_3446);
nor U3571 (N_3571,N_3261,N_3256);
nand U3572 (N_3572,N_3467,N_3321);
nor U3573 (N_3573,N_3494,N_3435);
nand U3574 (N_3574,N_3440,N_3310);
and U3575 (N_3575,N_3342,N_3473);
nor U3576 (N_3576,N_3266,N_3265);
or U3577 (N_3577,N_3375,N_3286);
nor U3578 (N_3578,N_3314,N_3434);
and U3579 (N_3579,N_3386,N_3408);
xor U3580 (N_3580,N_3306,N_3349);
nand U3581 (N_3581,N_3462,N_3442);
or U3582 (N_3582,N_3354,N_3409);
nand U3583 (N_3583,N_3264,N_3363);
and U3584 (N_3584,N_3471,N_3483);
and U3585 (N_3585,N_3277,N_3263);
or U3586 (N_3586,N_3350,N_3369);
nor U3587 (N_3587,N_3273,N_3270);
and U3588 (N_3588,N_3455,N_3269);
nor U3589 (N_3589,N_3484,N_3411);
nand U3590 (N_3590,N_3279,N_3426);
or U3591 (N_3591,N_3390,N_3367);
nand U3592 (N_3592,N_3330,N_3282);
xnor U3593 (N_3593,N_3288,N_3481);
nor U3594 (N_3594,N_3290,N_3356);
nor U3595 (N_3595,N_3276,N_3489);
and U3596 (N_3596,N_3480,N_3329);
and U3597 (N_3597,N_3328,N_3260);
and U3598 (N_3598,N_3383,N_3482);
nor U3599 (N_3599,N_3357,N_3331);
and U3600 (N_3600,N_3452,N_3334);
or U3601 (N_3601,N_3374,N_3401);
nor U3602 (N_3602,N_3382,N_3360);
or U3603 (N_3603,N_3301,N_3461);
nor U3604 (N_3604,N_3389,N_3427);
or U3605 (N_3605,N_3305,N_3373);
or U3606 (N_3606,N_3327,N_3439);
and U3607 (N_3607,N_3345,N_3317);
nand U3608 (N_3608,N_3475,N_3257);
or U3609 (N_3609,N_3311,N_3271);
nor U3610 (N_3610,N_3478,N_3362);
nor U3611 (N_3611,N_3259,N_3395);
nand U3612 (N_3612,N_3372,N_3437);
and U3613 (N_3613,N_3353,N_3438);
nand U3614 (N_3614,N_3370,N_3414);
or U3615 (N_3615,N_3429,N_3324);
and U3616 (N_3616,N_3352,N_3316);
nand U3617 (N_3617,N_3488,N_3441);
nor U3618 (N_3618,N_3385,N_3422);
nand U3619 (N_3619,N_3297,N_3291);
or U3620 (N_3620,N_3472,N_3358);
or U3621 (N_3621,N_3496,N_3255);
and U3622 (N_3622,N_3251,N_3359);
nand U3623 (N_3623,N_3253,N_3493);
or U3624 (N_3624,N_3333,N_3339);
or U3625 (N_3625,N_3409,N_3457);
nand U3626 (N_3626,N_3453,N_3416);
or U3627 (N_3627,N_3258,N_3289);
nand U3628 (N_3628,N_3458,N_3311);
nor U3629 (N_3629,N_3298,N_3337);
nor U3630 (N_3630,N_3485,N_3322);
or U3631 (N_3631,N_3437,N_3284);
and U3632 (N_3632,N_3285,N_3448);
or U3633 (N_3633,N_3276,N_3328);
and U3634 (N_3634,N_3310,N_3414);
nor U3635 (N_3635,N_3391,N_3329);
nand U3636 (N_3636,N_3471,N_3442);
and U3637 (N_3637,N_3318,N_3331);
or U3638 (N_3638,N_3472,N_3357);
and U3639 (N_3639,N_3312,N_3488);
nand U3640 (N_3640,N_3433,N_3350);
nor U3641 (N_3641,N_3456,N_3288);
nor U3642 (N_3642,N_3462,N_3293);
or U3643 (N_3643,N_3363,N_3300);
or U3644 (N_3644,N_3410,N_3333);
or U3645 (N_3645,N_3358,N_3465);
and U3646 (N_3646,N_3496,N_3473);
and U3647 (N_3647,N_3372,N_3289);
nand U3648 (N_3648,N_3364,N_3323);
nand U3649 (N_3649,N_3446,N_3394);
and U3650 (N_3650,N_3302,N_3450);
nor U3651 (N_3651,N_3285,N_3280);
or U3652 (N_3652,N_3314,N_3346);
nand U3653 (N_3653,N_3294,N_3446);
xnor U3654 (N_3654,N_3408,N_3478);
nand U3655 (N_3655,N_3435,N_3255);
or U3656 (N_3656,N_3320,N_3337);
and U3657 (N_3657,N_3476,N_3317);
nand U3658 (N_3658,N_3323,N_3392);
and U3659 (N_3659,N_3349,N_3400);
nor U3660 (N_3660,N_3396,N_3316);
nand U3661 (N_3661,N_3444,N_3391);
or U3662 (N_3662,N_3464,N_3308);
xnor U3663 (N_3663,N_3358,N_3442);
nand U3664 (N_3664,N_3416,N_3253);
nor U3665 (N_3665,N_3442,N_3265);
or U3666 (N_3666,N_3301,N_3463);
and U3667 (N_3667,N_3421,N_3433);
or U3668 (N_3668,N_3412,N_3292);
and U3669 (N_3669,N_3428,N_3477);
or U3670 (N_3670,N_3259,N_3314);
or U3671 (N_3671,N_3412,N_3360);
xnor U3672 (N_3672,N_3453,N_3255);
xor U3673 (N_3673,N_3428,N_3455);
nor U3674 (N_3674,N_3257,N_3439);
nor U3675 (N_3675,N_3465,N_3371);
or U3676 (N_3676,N_3385,N_3379);
nor U3677 (N_3677,N_3405,N_3400);
nor U3678 (N_3678,N_3381,N_3314);
nor U3679 (N_3679,N_3350,N_3413);
nand U3680 (N_3680,N_3358,N_3335);
xnor U3681 (N_3681,N_3361,N_3274);
and U3682 (N_3682,N_3496,N_3465);
xor U3683 (N_3683,N_3322,N_3280);
nor U3684 (N_3684,N_3340,N_3430);
and U3685 (N_3685,N_3494,N_3272);
xor U3686 (N_3686,N_3319,N_3406);
nor U3687 (N_3687,N_3259,N_3257);
nor U3688 (N_3688,N_3395,N_3412);
nand U3689 (N_3689,N_3451,N_3324);
and U3690 (N_3690,N_3259,N_3487);
xnor U3691 (N_3691,N_3484,N_3288);
xnor U3692 (N_3692,N_3422,N_3302);
or U3693 (N_3693,N_3327,N_3254);
nor U3694 (N_3694,N_3391,N_3412);
nor U3695 (N_3695,N_3498,N_3296);
nand U3696 (N_3696,N_3302,N_3389);
nor U3697 (N_3697,N_3489,N_3498);
nand U3698 (N_3698,N_3263,N_3438);
and U3699 (N_3699,N_3461,N_3358);
xnor U3700 (N_3700,N_3479,N_3447);
and U3701 (N_3701,N_3460,N_3251);
xnor U3702 (N_3702,N_3322,N_3294);
nand U3703 (N_3703,N_3344,N_3325);
nor U3704 (N_3704,N_3282,N_3484);
and U3705 (N_3705,N_3367,N_3365);
or U3706 (N_3706,N_3414,N_3426);
nor U3707 (N_3707,N_3363,N_3480);
nand U3708 (N_3708,N_3332,N_3316);
nor U3709 (N_3709,N_3422,N_3289);
xnor U3710 (N_3710,N_3456,N_3353);
or U3711 (N_3711,N_3341,N_3284);
or U3712 (N_3712,N_3367,N_3495);
nor U3713 (N_3713,N_3292,N_3470);
nor U3714 (N_3714,N_3400,N_3489);
nor U3715 (N_3715,N_3458,N_3498);
or U3716 (N_3716,N_3317,N_3372);
nand U3717 (N_3717,N_3411,N_3348);
xnor U3718 (N_3718,N_3406,N_3480);
nand U3719 (N_3719,N_3403,N_3311);
and U3720 (N_3720,N_3250,N_3291);
nand U3721 (N_3721,N_3333,N_3292);
nor U3722 (N_3722,N_3457,N_3479);
nand U3723 (N_3723,N_3280,N_3414);
xor U3724 (N_3724,N_3415,N_3432);
nor U3725 (N_3725,N_3423,N_3372);
nand U3726 (N_3726,N_3279,N_3360);
or U3727 (N_3727,N_3484,N_3439);
xnor U3728 (N_3728,N_3419,N_3401);
nor U3729 (N_3729,N_3370,N_3272);
and U3730 (N_3730,N_3340,N_3362);
or U3731 (N_3731,N_3320,N_3486);
and U3732 (N_3732,N_3481,N_3329);
xor U3733 (N_3733,N_3297,N_3457);
or U3734 (N_3734,N_3375,N_3355);
nand U3735 (N_3735,N_3373,N_3464);
nand U3736 (N_3736,N_3295,N_3304);
nor U3737 (N_3737,N_3414,N_3465);
or U3738 (N_3738,N_3490,N_3341);
nand U3739 (N_3739,N_3371,N_3399);
nor U3740 (N_3740,N_3493,N_3375);
and U3741 (N_3741,N_3318,N_3338);
or U3742 (N_3742,N_3377,N_3385);
or U3743 (N_3743,N_3402,N_3391);
or U3744 (N_3744,N_3312,N_3490);
nor U3745 (N_3745,N_3307,N_3298);
nand U3746 (N_3746,N_3499,N_3304);
nor U3747 (N_3747,N_3377,N_3414);
nor U3748 (N_3748,N_3428,N_3346);
nor U3749 (N_3749,N_3320,N_3386);
nor U3750 (N_3750,N_3559,N_3608);
nor U3751 (N_3751,N_3692,N_3554);
nand U3752 (N_3752,N_3556,N_3683);
or U3753 (N_3753,N_3714,N_3731);
nor U3754 (N_3754,N_3569,N_3504);
or U3755 (N_3755,N_3696,N_3733);
and U3756 (N_3756,N_3663,N_3667);
and U3757 (N_3757,N_3720,N_3526);
nand U3758 (N_3758,N_3558,N_3678);
and U3759 (N_3759,N_3599,N_3594);
and U3760 (N_3760,N_3681,N_3536);
nor U3761 (N_3761,N_3735,N_3549);
nor U3762 (N_3762,N_3575,N_3564);
and U3763 (N_3763,N_3617,N_3747);
or U3764 (N_3764,N_3623,N_3650);
or U3765 (N_3765,N_3621,N_3545);
nand U3766 (N_3766,N_3652,N_3719);
and U3767 (N_3767,N_3689,N_3567);
nand U3768 (N_3768,N_3505,N_3518);
nand U3769 (N_3769,N_3664,N_3609);
nand U3770 (N_3770,N_3618,N_3588);
or U3771 (N_3771,N_3710,N_3568);
or U3772 (N_3772,N_3613,N_3566);
nand U3773 (N_3773,N_3627,N_3723);
nor U3774 (N_3774,N_3637,N_3532);
xor U3775 (N_3775,N_3639,N_3745);
and U3776 (N_3776,N_3573,N_3534);
or U3777 (N_3777,N_3645,N_3516);
nor U3778 (N_3778,N_3682,N_3749);
and U3779 (N_3779,N_3711,N_3501);
nand U3780 (N_3780,N_3625,N_3700);
and U3781 (N_3781,N_3633,N_3661);
or U3782 (N_3782,N_3697,N_3699);
nand U3783 (N_3783,N_3514,N_3522);
or U3784 (N_3784,N_3541,N_3595);
nor U3785 (N_3785,N_3644,N_3548);
nor U3786 (N_3786,N_3523,N_3676);
or U3787 (N_3787,N_3726,N_3744);
or U3788 (N_3788,N_3748,N_3631);
and U3789 (N_3789,N_3651,N_3668);
and U3790 (N_3790,N_3643,N_3592);
or U3791 (N_3791,N_3602,N_3646);
or U3792 (N_3792,N_3725,N_3597);
and U3793 (N_3793,N_3641,N_3611);
nor U3794 (N_3794,N_3677,N_3574);
and U3795 (N_3795,N_3578,N_3691);
and U3796 (N_3796,N_3557,N_3553);
and U3797 (N_3797,N_3738,N_3584);
and U3798 (N_3798,N_3577,N_3622);
nand U3799 (N_3799,N_3603,N_3674);
and U3800 (N_3800,N_3743,N_3620);
nor U3801 (N_3801,N_3734,N_3636);
nor U3802 (N_3802,N_3737,N_3552);
xnor U3803 (N_3803,N_3724,N_3590);
nand U3804 (N_3804,N_3629,N_3693);
nand U3805 (N_3805,N_3585,N_3528);
nand U3806 (N_3806,N_3741,N_3601);
nor U3807 (N_3807,N_3600,N_3510);
or U3808 (N_3808,N_3686,N_3647);
nor U3809 (N_3809,N_3571,N_3730);
nor U3810 (N_3810,N_3687,N_3517);
nor U3811 (N_3811,N_3746,N_3721);
or U3812 (N_3812,N_3648,N_3582);
nand U3813 (N_3813,N_3593,N_3628);
nor U3814 (N_3814,N_3565,N_3708);
nand U3815 (N_3815,N_3580,N_3550);
nor U3816 (N_3816,N_3685,N_3511);
or U3817 (N_3817,N_3722,N_3515);
xor U3818 (N_3818,N_3519,N_3576);
nand U3819 (N_3819,N_3665,N_3598);
nor U3820 (N_3820,N_3736,N_3537);
or U3821 (N_3821,N_3655,N_3555);
nand U3822 (N_3822,N_3521,N_3702);
nand U3823 (N_3823,N_3589,N_3539);
or U3824 (N_3824,N_3562,N_3704);
and U3825 (N_3825,N_3642,N_3507);
and U3826 (N_3826,N_3503,N_3560);
or U3827 (N_3827,N_3531,N_3551);
and U3828 (N_3828,N_3508,N_3561);
nand U3829 (N_3829,N_3690,N_3701);
or U3830 (N_3830,N_3624,N_3524);
nand U3831 (N_3831,N_3614,N_3707);
nor U3832 (N_3832,N_3649,N_3538);
xor U3833 (N_3833,N_3583,N_3640);
or U3834 (N_3834,N_3657,N_3672);
nand U3835 (N_3835,N_3610,N_3671);
or U3836 (N_3836,N_3506,N_3713);
nor U3837 (N_3837,N_3616,N_3688);
and U3838 (N_3838,N_3679,N_3654);
nand U3839 (N_3839,N_3615,N_3572);
nor U3840 (N_3840,N_3675,N_3729);
nand U3841 (N_3841,N_3509,N_3604);
and U3842 (N_3842,N_3695,N_3732);
or U3843 (N_3843,N_3543,N_3706);
xnor U3844 (N_3844,N_3638,N_3634);
and U3845 (N_3845,N_3658,N_3540);
or U3846 (N_3846,N_3742,N_3513);
or U3847 (N_3847,N_3606,N_3612);
nand U3848 (N_3848,N_3662,N_3666);
xnor U3849 (N_3849,N_3669,N_3717);
nor U3850 (N_3850,N_3563,N_3533);
xnor U3851 (N_3851,N_3596,N_3512);
or U3852 (N_3852,N_3535,N_3739);
or U3853 (N_3853,N_3659,N_3709);
and U3854 (N_3854,N_3626,N_3716);
xnor U3855 (N_3855,N_3547,N_3656);
xor U3856 (N_3856,N_3712,N_3607);
nor U3857 (N_3857,N_3591,N_3698);
nand U3858 (N_3858,N_3619,N_3605);
and U3859 (N_3859,N_3630,N_3529);
and U3860 (N_3860,N_3544,N_3546);
and U3861 (N_3861,N_3740,N_3670);
or U3862 (N_3862,N_3694,N_3705);
or U3863 (N_3863,N_3570,N_3715);
and U3864 (N_3864,N_3520,N_3530);
or U3865 (N_3865,N_3718,N_3635);
or U3866 (N_3866,N_3673,N_3542);
and U3867 (N_3867,N_3632,N_3502);
and U3868 (N_3868,N_3581,N_3579);
and U3869 (N_3869,N_3527,N_3525);
or U3870 (N_3870,N_3680,N_3500);
or U3871 (N_3871,N_3703,N_3684);
and U3872 (N_3872,N_3586,N_3727);
or U3873 (N_3873,N_3653,N_3587);
nand U3874 (N_3874,N_3728,N_3660);
nor U3875 (N_3875,N_3586,N_3747);
nor U3876 (N_3876,N_3744,N_3557);
nor U3877 (N_3877,N_3585,N_3563);
and U3878 (N_3878,N_3685,N_3590);
xnor U3879 (N_3879,N_3681,N_3654);
nor U3880 (N_3880,N_3505,N_3644);
nand U3881 (N_3881,N_3605,N_3637);
nand U3882 (N_3882,N_3668,N_3720);
or U3883 (N_3883,N_3727,N_3559);
or U3884 (N_3884,N_3537,N_3684);
nand U3885 (N_3885,N_3546,N_3647);
or U3886 (N_3886,N_3742,N_3565);
nor U3887 (N_3887,N_3631,N_3599);
or U3888 (N_3888,N_3534,N_3675);
xnor U3889 (N_3889,N_3637,N_3727);
or U3890 (N_3890,N_3601,N_3553);
xnor U3891 (N_3891,N_3693,N_3612);
xor U3892 (N_3892,N_3547,N_3628);
or U3893 (N_3893,N_3688,N_3500);
nor U3894 (N_3894,N_3580,N_3651);
xnor U3895 (N_3895,N_3645,N_3699);
or U3896 (N_3896,N_3668,N_3719);
or U3897 (N_3897,N_3541,N_3669);
nand U3898 (N_3898,N_3643,N_3515);
or U3899 (N_3899,N_3703,N_3719);
and U3900 (N_3900,N_3653,N_3713);
nor U3901 (N_3901,N_3516,N_3606);
or U3902 (N_3902,N_3620,N_3740);
nand U3903 (N_3903,N_3619,N_3677);
and U3904 (N_3904,N_3553,N_3597);
nor U3905 (N_3905,N_3543,N_3533);
and U3906 (N_3906,N_3571,N_3630);
nor U3907 (N_3907,N_3746,N_3633);
nand U3908 (N_3908,N_3647,N_3629);
xor U3909 (N_3909,N_3740,N_3506);
or U3910 (N_3910,N_3629,N_3543);
or U3911 (N_3911,N_3618,N_3728);
nand U3912 (N_3912,N_3506,N_3694);
or U3913 (N_3913,N_3723,N_3567);
and U3914 (N_3914,N_3704,N_3512);
xor U3915 (N_3915,N_3573,N_3539);
nor U3916 (N_3916,N_3746,N_3523);
xor U3917 (N_3917,N_3579,N_3659);
nor U3918 (N_3918,N_3716,N_3609);
nor U3919 (N_3919,N_3557,N_3698);
nand U3920 (N_3920,N_3572,N_3521);
nor U3921 (N_3921,N_3502,N_3669);
and U3922 (N_3922,N_3653,N_3715);
or U3923 (N_3923,N_3539,N_3551);
nor U3924 (N_3924,N_3530,N_3742);
or U3925 (N_3925,N_3540,N_3523);
and U3926 (N_3926,N_3610,N_3568);
or U3927 (N_3927,N_3713,N_3740);
and U3928 (N_3928,N_3515,N_3584);
nand U3929 (N_3929,N_3537,N_3742);
and U3930 (N_3930,N_3587,N_3654);
nor U3931 (N_3931,N_3626,N_3669);
nor U3932 (N_3932,N_3563,N_3611);
nor U3933 (N_3933,N_3591,N_3616);
nor U3934 (N_3934,N_3710,N_3687);
nand U3935 (N_3935,N_3606,N_3555);
nor U3936 (N_3936,N_3589,N_3555);
nand U3937 (N_3937,N_3539,N_3683);
or U3938 (N_3938,N_3572,N_3646);
and U3939 (N_3939,N_3707,N_3535);
or U3940 (N_3940,N_3626,N_3654);
xor U3941 (N_3941,N_3647,N_3579);
or U3942 (N_3942,N_3706,N_3672);
and U3943 (N_3943,N_3626,N_3711);
and U3944 (N_3944,N_3535,N_3606);
and U3945 (N_3945,N_3653,N_3660);
or U3946 (N_3946,N_3528,N_3647);
xor U3947 (N_3947,N_3705,N_3739);
nor U3948 (N_3948,N_3725,N_3636);
nor U3949 (N_3949,N_3502,N_3723);
or U3950 (N_3950,N_3718,N_3572);
and U3951 (N_3951,N_3692,N_3721);
and U3952 (N_3952,N_3593,N_3607);
nor U3953 (N_3953,N_3646,N_3745);
nand U3954 (N_3954,N_3695,N_3650);
and U3955 (N_3955,N_3570,N_3691);
or U3956 (N_3956,N_3725,N_3557);
xnor U3957 (N_3957,N_3748,N_3663);
or U3958 (N_3958,N_3682,N_3574);
nand U3959 (N_3959,N_3546,N_3599);
nor U3960 (N_3960,N_3601,N_3663);
and U3961 (N_3961,N_3514,N_3721);
or U3962 (N_3962,N_3662,N_3676);
nand U3963 (N_3963,N_3703,N_3717);
nor U3964 (N_3964,N_3697,N_3687);
xor U3965 (N_3965,N_3565,N_3677);
nand U3966 (N_3966,N_3560,N_3739);
nand U3967 (N_3967,N_3717,N_3564);
and U3968 (N_3968,N_3506,N_3638);
nor U3969 (N_3969,N_3675,N_3688);
or U3970 (N_3970,N_3509,N_3582);
and U3971 (N_3971,N_3672,N_3678);
nor U3972 (N_3972,N_3521,N_3697);
nor U3973 (N_3973,N_3532,N_3708);
nor U3974 (N_3974,N_3611,N_3526);
nand U3975 (N_3975,N_3549,N_3626);
and U3976 (N_3976,N_3500,N_3507);
and U3977 (N_3977,N_3508,N_3618);
and U3978 (N_3978,N_3511,N_3536);
nand U3979 (N_3979,N_3574,N_3537);
nor U3980 (N_3980,N_3529,N_3589);
and U3981 (N_3981,N_3518,N_3565);
and U3982 (N_3982,N_3525,N_3540);
nand U3983 (N_3983,N_3551,N_3569);
nor U3984 (N_3984,N_3713,N_3542);
xnor U3985 (N_3985,N_3662,N_3562);
and U3986 (N_3986,N_3667,N_3634);
nor U3987 (N_3987,N_3509,N_3704);
nand U3988 (N_3988,N_3502,N_3573);
nand U3989 (N_3989,N_3517,N_3628);
and U3990 (N_3990,N_3528,N_3749);
or U3991 (N_3991,N_3653,N_3648);
and U3992 (N_3992,N_3747,N_3608);
nand U3993 (N_3993,N_3720,N_3702);
and U3994 (N_3994,N_3600,N_3743);
xor U3995 (N_3995,N_3653,N_3540);
nor U3996 (N_3996,N_3728,N_3580);
xnor U3997 (N_3997,N_3702,N_3575);
or U3998 (N_3998,N_3659,N_3695);
nor U3999 (N_3999,N_3637,N_3733);
nand U4000 (N_4000,N_3843,N_3776);
nor U4001 (N_4001,N_3811,N_3787);
nand U4002 (N_4002,N_3856,N_3880);
nand U4003 (N_4003,N_3812,N_3955);
xor U4004 (N_4004,N_3781,N_3762);
nand U4005 (N_4005,N_3930,N_3840);
and U4006 (N_4006,N_3866,N_3932);
and U4007 (N_4007,N_3879,N_3992);
nand U4008 (N_4008,N_3967,N_3792);
or U4009 (N_4009,N_3935,N_3860);
xnor U4010 (N_4010,N_3874,N_3821);
and U4011 (N_4011,N_3844,N_3814);
nor U4012 (N_4012,N_3906,N_3993);
nor U4013 (N_4013,N_3859,N_3914);
xnor U4014 (N_4014,N_3858,N_3966);
nor U4015 (N_4015,N_3928,N_3940);
nand U4016 (N_4016,N_3852,N_3757);
and U4017 (N_4017,N_3962,N_3845);
and U4018 (N_4018,N_3897,N_3803);
nand U4019 (N_4019,N_3995,N_3754);
nand U4020 (N_4020,N_3944,N_3790);
nand U4021 (N_4021,N_3875,N_3945);
nor U4022 (N_4022,N_3975,N_3828);
or U4023 (N_4023,N_3902,N_3947);
nor U4024 (N_4024,N_3881,N_3893);
nor U4025 (N_4025,N_3786,N_3989);
and U4026 (N_4026,N_3837,N_3824);
nor U4027 (N_4027,N_3861,N_3959);
nor U4028 (N_4028,N_3823,N_3931);
and U4029 (N_4029,N_3949,N_3974);
nand U4030 (N_4030,N_3951,N_3753);
nand U4031 (N_4031,N_3923,N_3789);
or U4032 (N_4032,N_3991,N_3791);
nand U4033 (N_4033,N_3808,N_3817);
nor U4034 (N_4034,N_3885,N_3954);
or U4035 (N_4035,N_3934,N_3984);
and U4036 (N_4036,N_3977,N_3976);
nor U4037 (N_4037,N_3867,N_3765);
nor U4038 (N_4038,N_3807,N_3898);
and U4039 (N_4039,N_3957,N_3756);
and U4040 (N_4040,N_3761,N_3985);
or U4041 (N_4041,N_3942,N_3848);
nor U4042 (N_4042,N_3876,N_3889);
xor U4043 (N_4043,N_3799,N_3750);
and U4044 (N_4044,N_3784,N_3963);
nand U4045 (N_4045,N_3903,N_3948);
nand U4046 (N_4046,N_3771,N_3924);
nor U4047 (N_4047,N_3982,N_3830);
nor U4048 (N_4048,N_3968,N_3895);
nor U4049 (N_4049,N_3887,N_3758);
nor U4050 (N_4050,N_3805,N_3978);
nand U4051 (N_4051,N_3904,N_3869);
nor U4052 (N_4052,N_3853,N_3990);
or U4053 (N_4053,N_3809,N_3936);
nand U4054 (N_4054,N_3846,N_3818);
xnor U4055 (N_4055,N_3788,N_3910);
or U4056 (N_4056,N_3822,N_3933);
nand U4057 (N_4057,N_3804,N_3836);
nor U4058 (N_4058,N_3892,N_3891);
and U4059 (N_4059,N_3827,N_3883);
or U4060 (N_4060,N_3922,N_3801);
nor U4061 (N_4061,N_3973,N_3868);
nand U4062 (N_4062,N_3796,N_3926);
nor U4063 (N_4063,N_3981,N_3983);
nand U4064 (N_4064,N_3829,N_3912);
and U4065 (N_4065,N_3911,N_3908);
and U4066 (N_4066,N_3873,N_3964);
and U4067 (N_4067,N_3986,N_3886);
nor U4068 (N_4068,N_3943,N_3938);
or U4069 (N_4069,N_3941,N_3939);
and U4070 (N_4070,N_3920,N_3764);
and U4071 (N_4071,N_3815,N_3970);
and U4072 (N_4072,N_3917,N_3996);
and U4073 (N_4073,N_3806,N_3839);
nor U4074 (N_4074,N_3888,N_3950);
nand U4075 (N_4075,N_3864,N_3958);
nand U4076 (N_4076,N_3820,N_3851);
or U4077 (N_4077,N_3766,N_3831);
nor U4078 (N_4078,N_3913,N_3872);
nor U4079 (N_4079,N_3863,N_3979);
and U4080 (N_4080,N_3795,N_3779);
or U4081 (N_4081,N_3797,N_3834);
xor U4082 (N_4082,N_3819,N_3921);
nor U4083 (N_4083,N_3772,N_3965);
and U4084 (N_4084,N_3751,N_3918);
or U4085 (N_4085,N_3838,N_3961);
xnor U4086 (N_4086,N_3870,N_3773);
nor U4087 (N_4087,N_3901,N_3810);
xor U4088 (N_4088,N_3915,N_3849);
nor U4089 (N_4089,N_3826,N_3907);
nand U4090 (N_4090,N_3988,N_3782);
nor U4091 (N_4091,N_3878,N_3953);
nor U4092 (N_4092,N_3850,N_3987);
and U4093 (N_4093,N_3816,N_3777);
or U4094 (N_4094,N_3835,N_3775);
or U4095 (N_4095,N_3998,N_3842);
nand U4096 (N_4096,N_3882,N_3884);
nand U4097 (N_4097,N_3800,N_3755);
nand U4098 (N_4098,N_3905,N_3952);
or U4099 (N_4099,N_3890,N_3927);
nor U4100 (N_4100,N_3929,N_3972);
and U4101 (N_4101,N_3847,N_3774);
or U4102 (N_4102,N_3862,N_3999);
and U4103 (N_4103,N_3971,N_3813);
nand U4104 (N_4104,N_3763,N_3794);
nor U4105 (N_4105,N_3937,N_3767);
and U4106 (N_4106,N_3785,N_3894);
nor U4107 (N_4107,N_3769,N_3841);
nand U4108 (N_4108,N_3798,N_3778);
xor U4109 (N_4109,N_3857,N_3997);
or U4110 (N_4110,N_3832,N_3768);
and U4111 (N_4111,N_3752,N_3871);
nor U4112 (N_4112,N_3994,N_3780);
and U4113 (N_4113,N_3802,N_3916);
nor U4114 (N_4114,N_3896,N_3899);
xnor U4115 (N_4115,N_3969,N_3759);
nor U4116 (N_4116,N_3946,N_3770);
and U4117 (N_4117,N_3855,N_3909);
nand U4118 (N_4118,N_3783,N_3925);
nand U4119 (N_4119,N_3900,N_3877);
and U4120 (N_4120,N_3980,N_3865);
or U4121 (N_4121,N_3793,N_3956);
and U4122 (N_4122,N_3825,N_3854);
nor U4123 (N_4123,N_3960,N_3919);
or U4124 (N_4124,N_3760,N_3833);
nor U4125 (N_4125,N_3890,N_3751);
or U4126 (N_4126,N_3972,N_3968);
nor U4127 (N_4127,N_3765,N_3757);
xor U4128 (N_4128,N_3754,N_3981);
nand U4129 (N_4129,N_3838,N_3975);
xnor U4130 (N_4130,N_3981,N_3915);
nand U4131 (N_4131,N_3802,N_3881);
nand U4132 (N_4132,N_3828,N_3797);
or U4133 (N_4133,N_3955,N_3866);
and U4134 (N_4134,N_3859,N_3991);
and U4135 (N_4135,N_3766,N_3849);
nand U4136 (N_4136,N_3928,N_3793);
and U4137 (N_4137,N_3752,N_3996);
or U4138 (N_4138,N_3761,N_3908);
xor U4139 (N_4139,N_3908,N_3894);
nand U4140 (N_4140,N_3847,N_3831);
nand U4141 (N_4141,N_3929,N_3962);
nor U4142 (N_4142,N_3809,N_3901);
nor U4143 (N_4143,N_3793,N_3784);
nor U4144 (N_4144,N_3891,N_3917);
xor U4145 (N_4145,N_3811,N_3842);
nand U4146 (N_4146,N_3966,N_3983);
nand U4147 (N_4147,N_3846,N_3751);
xor U4148 (N_4148,N_3819,N_3783);
nor U4149 (N_4149,N_3876,N_3917);
xor U4150 (N_4150,N_3885,N_3842);
nor U4151 (N_4151,N_3853,N_3900);
nor U4152 (N_4152,N_3833,N_3964);
or U4153 (N_4153,N_3963,N_3921);
or U4154 (N_4154,N_3806,N_3753);
and U4155 (N_4155,N_3902,N_3839);
nand U4156 (N_4156,N_3930,N_3813);
or U4157 (N_4157,N_3993,N_3945);
nor U4158 (N_4158,N_3890,N_3784);
and U4159 (N_4159,N_3992,N_3918);
nand U4160 (N_4160,N_3940,N_3936);
and U4161 (N_4161,N_3990,N_3897);
or U4162 (N_4162,N_3816,N_3849);
or U4163 (N_4163,N_3923,N_3835);
nand U4164 (N_4164,N_3821,N_3936);
nor U4165 (N_4165,N_3909,N_3946);
and U4166 (N_4166,N_3775,N_3949);
and U4167 (N_4167,N_3772,N_3951);
nor U4168 (N_4168,N_3793,N_3779);
or U4169 (N_4169,N_3934,N_3831);
or U4170 (N_4170,N_3937,N_3751);
or U4171 (N_4171,N_3850,N_3775);
nor U4172 (N_4172,N_3928,N_3809);
or U4173 (N_4173,N_3965,N_3866);
nor U4174 (N_4174,N_3980,N_3988);
and U4175 (N_4175,N_3953,N_3925);
nor U4176 (N_4176,N_3830,N_3791);
or U4177 (N_4177,N_3813,N_3866);
and U4178 (N_4178,N_3815,N_3784);
nor U4179 (N_4179,N_3856,N_3909);
or U4180 (N_4180,N_3860,N_3845);
nor U4181 (N_4181,N_3967,N_3916);
nand U4182 (N_4182,N_3854,N_3842);
nand U4183 (N_4183,N_3779,N_3756);
xor U4184 (N_4184,N_3795,N_3861);
or U4185 (N_4185,N_3936,N_3874);
nand U4186 (N_4186,N_3896,N_3973);
and U4187 (N_4187,N_3937,N_3846);
nand U4188 (N_4188,N_3930,N_3868);
or U4189 (N_4189,N_3987,N_3957);
or U4190 (N_4190,N_3820,N_3996);
nand U4191 (N_4191,N_3924,N_3995);
or U4192 (N_4192,N_3842,N_3879);
xnor U4193 (N_4193,N_3800,N_3971);
nand U4194 (N_4194,N_3927,N_3873);
nand U4195 (N_4195,N_3844,N_3811);
and U4196 (N_4196,N_3849,N_3798);
and U4197 (N_4197,N_3828,N_3830);
xor U4198 (N_4198,N_3816,N_3844);
and U4199 (N_4199,N_3857,N_3798);
or U4200 (N_4200,N_3944,N_3993);
nand U4201 (N_4201,N_3792,N_3826);
and U4202 (N_4202,N_3824,N_3895);
xnor U4203 (N_4203,N_3765,N_3773);
nor U4204 (N_4204,N_3924,N_3849);
nor U4205 (N_4205,N_3774,N_3830);
and U4206 (N_4206,N_3810,N_3758);
xor U4207 (N_4207,N_3971,N_3806);
nand U4208 (N_4208,N_3876,N_3982);
xor U4209 (N_4209,N_3859,N_3755);
or U4210 (N_4210,N_3958,N_3886);
xor U4211 (N_4211,N_3849,N_3980);
or U4212 (N_4212,N_3956,N_3891);
or U4213 (N_4213,N_3916,N_3965);
and U4214 (N_4214,N_3788,N_3829);
and U4215 (N_4215,N_3925,N_3811);
xor U4216 (N_4216,N_3862,N_3922);
or U4217 (N_4217,N_3786,N_3942);
xor U4218 (N_4218,N_3804,N_3991);
or U4219 (N_4219,N_3858,N_3962);
and U4220 (N_4220,N_3808,N_3893);
and U4221 (N_4221,N_3894,N_3838);
or U4222 (N_4222,N_3975,N_3946);
and U4223 (N_4223,N_3943,N_3793);
nand U4224 (N_4224,N_3964,N_3921);
xor U4225 (N_4225,N_3764,N_3976);
nand U4226 (N_4226,N_3793,N_3910);
nor U4227 (N_4227,N_3886,N_3940);
or U4228 (N_4228,N_3886,N_3951);
and U4229 (N_4229,N_3939,N_3909);
xnor U4230 (N_4230,N_3770,N_3907);
nand U4231 (N_4231,N_3792,N_3865);
or U4232 (N_4232,N_3892,N_3977);
or U4233 (N_4233,N_3783,N_3785);
nand U4234 (N_4234,N_3809,N_3817);
or U4235 (N_4235,N_3990,N_3936);
or U4236 (N_4236,N_3789,N_3762);
nand U4237 (N_4237,N_3929,N_3912);
or U4238 (N_4238,N_3834,N_3893);
nand U4239 (N_4239,N_3873,N_3823);
or U4240 (N_4240,N_3818,N_3990);
or U4241 (N_4241,N_3875,N_3993);
and U4242 (N_4242,N_3867,N_3988);
nor U4243 (N_4243,N_3871,N_3987);
or U4244 (N_4244,N_3957,N_3811);
nand U4245 (N_4245,N_3898,N_3966);
or U4246 (N_4246,N_3901,N_3914);
and U4247 (N_4247,N_3886,N_3907);
xor U4248 (N_4248,N_3967,N_3846);
or U4249 (N_4249,N_3810,N_3892);
nor U4250 (N_4250,N_4239,N_4090);
or U4251 (N_4251,N_4077,N_4231);
nand U4252 (N_4252,N_4111,N_4218);
nor U4253 (N_4253,N_4185,N_4027);
and U4254 (N_4254,N_4045,N_4122);
nor U4255 (N_4255,N_4242,N_4119);
and U4256 (N_4256,N_4088,N_4143);
nand U4257 (N_4257,N_4219,N_4205);
or U4258 (N_4258,N_4236,N_4189);
or U4259 (N_4259,N_4164,N_4015);
and U4260 (N_4260,N_4232,N_4136);
or U4261 (N_4261,N_4181,N_4028);
xor U4262 (N_4262,N_4041,N_4073);
nor U4263 (N_4263,N_4078,N_4179);
or U4264 (N_4264,N_4135,N_4032);
xor U4265 (N_4265,N_4156,N_4116);
nor U4266 (N_4266,N_4106,N_4142);
nor U4267 (N_4267,N_4200,N_4021);
nor U4268 (N_4268,N_4153,N_4033);
nor U4269 (N_4269,N_4139,N_4000);
nand U4270 (N_4270,N_4117,N_4210);
nor U4271 (N_4271,N_4020,N_4202);
and U4272 (N_4272,N_4040,N_4098);
or U4273 (N_4273,N_4050,N_4051);
nand U4274 (N_4274,N_4022,N_4221);
nand U4275 (N_4275,N_4230,N_4148);
or U4276 (N_4276,N_4204,N_4059);
xor U4277 (N_4277,N_4183,N_4114);
nor U4278 (N_4278,N_4245,N_4120);
and U4279 (N_4279,N_4100,N_4034);
and U4280 (N_4280,N_4154,N_4160);
xor U4281 (N_4281,N_4191,N_4223);
or U4282 (N_4282,N_4087,N_4084);
xor U4283 (N_4283,N_4099,N_4072);
xor U4284 (N_4284,N_4171,N_4151);
and U4285 (N_4285,N_4159,N_4101);
and U4286 (N_4286,N_4083,N_4125);
and U4287 (N_4287,N_4062,N_4064);
nor U4288 (N_4288,N_4080,N_4244);
and U4289 (N_4289,N_4076,N_4212);
and U4290 (N_4290,N_4203,N_4118);
and U4291 (N_4291,N_4161,N_4039);
or U4292 (N_4292,N_4158,N_4246);
nor U4293 (N_4293,N_4052,N_4126);
nand U4294 (N_4294,N_4047,N_4107);
nand U4295 (N_4295,N_4134,N_4030);
nand U4296 (N_4296,N_4197,N_4092);
or U4297 (N_4297,N_4070,N_4169);
or U4298 (N_4298,N_4056,N_4211);
and U4299 (N_4299,N_4109,N_4113);
and U4300 (N_4300,N_4140,N_4228);
or U4301 (N_4301,N_4168,N_4180);
and U4302 (N_4302,N_4121,N_4131);
and U4303 (N_4303,N_4075,N_4127);
nand U4304 (N_4304,N_4024,N_4123);
nor U4305 (N_4305,N_4137,N_4165);
nand U4306 (N_4306,N_4207,N_4178);
nand U4307 (N_4307,N_4166,N_4128);
and U4308 (N_4308,N_4152,N_4213);
or U4309 (N_4309,N_4048,N_4192);
or U4310 (N_4310,N_4019,N_4038);
nand U4311 (N_4311,N_4138,N_4014);
or U4312 (N_4312,N_4017,N_4103);
xnor U4313 (N_4313,N_4172,N_4147);
nand U4314 (N_4314,N_4155,N_4157);
or U4315 (N_4315,N_4068,N_4248);
xor U4316 (N_4316,N_4173,N_4054);
xor U4317 (N_4317,N_4074,N_4145);
or U4318 (N_4318,N_4217,N_4233);
nor U4319 (N_4319,N_4102,N_4225);
or U4320 (N_4320,N_4031,N_4081);
or U4321 (N_4321,N_4175,N_4067);
nand U4322 (N_4322,N_4141,N_4104);
nor U4323 (N_4323,N_4190,N_4243);
or U4324 (N_4324,N_4096,N_4079);
nor U4325 (N_4325,N_4177,N_4086);
nand U4326 (N_4326,N_4227,N_4133);
nand U4327 (N_4327,N_4012,N_4206);
nand U4328 (N_4328,N_4010,N_4186);
or U4329 (N_4329,N_4174,N_4201);
or U4330 (N_4330,N_4187,N_4115);
and U4331 (N_4331,N_4144,N_4044);
and U4332 (N_4332,N_4184,N_4007);
nand U4333 (N_4333,N_4235,N_4003);
xnor U4334 (N_4334,N_4105,N_4214);
or U4335 (N_4335,N_4129,N_4222);
and U4336 (N_4336,N_4193,N_4061);
nand U4337 (N_4337,N_4234,N_4237);
nor U4338 (N_4338,N_4216,N_4229);
or U4339 (N_4339,N_4240,N_4026);
xor U4340 (N_4340,N_4071,N_4198);
nor U4341 (N_4341,N_4063,N_4196);
and U4342 (N_4342,N_4001,N_4094);
nand U4343 (N_4343,N_4132,N_4009);
or U4344 (N_4344,N_4176,N_4149);
nand U4345 (N_4345,N_4209,N_4163);
nor U4346 (N_4346,N_4170,N_4167);
nand U4347 (N_4347,N_4037,N_4016);
nand U4348 (N_4348,N_4013,N_4004);
or U4349 (N_4349,N_4188,N_4005);
nor U4350 (N_4350,N_4124,N_4097);
nand U4351 (N_4351,N_4036,N_4091);
nor U4352 (N_4352,N_4042,N_4065);
xor U4353 (N_4353,N_4066,N_4162);
xnor U4354 (N_4354,N_4095,N_4008);
nand U4355 (N_4355,N_4089,N_4055);
and U4356 (N_4356,N_4215,N_4053);
and U4357 (N_4357,N_4110,N_4194);
and U4358 (N_4358,N_4057,N_4224);
nand U4359 (N_4359,N_4049,N_4035);
nor U4360 (N_4360,N_4060,N_4182);
or U4361 (N_4361,N_4043,N_4011);
and U4362 (N_4362,N_4006,N_4082);
nor U4363 (N_4363,N_4018,N_4023);
nand U4364 (N_4364,N_4069,N_4199);
or U4365 (N_4365,N_4247,N_4002);
nand U4366 (N_4366,N_4249,N_4025);
and U4367 (N_4367,N_4093,N_4058);
and U4368 (N_4368,N_4226,N_4108);
nand U4369 (N_4369,N_4241,N_4220);
and U4370 (N_4370,N_4208,N_4029);
nand U4371 (N_4371,N_4195,N_4150);
nand U4372 (N_4372,N_4238,N_4085);
nand U4373 (N_4373,N_4130,N_4046);
xor U4374 (N_4374,N_4146,N_4112);
and U4375 (N_4375,N_4018,N_4226);
and U4376 (N_4376,N_4118,N_4207);
nor U4377 (N_4377,N_4226,N_4065);
nand U4378 (N_4378,N_4170,N_4106);
nand U4379 (N_4379,N_4154,N_4074);
or U4380 (N_4380,N_4031,N_4089);
and U4381 (N_4381,N_4135,N_4003);
and U4382 (N_4382,N_4244,N_4057);
nand U4383 (N_4383,N_4020,N_4235);
nand U4384 (N_4384,N_4143,N_4065);
or U4385 (N_4385,N_4064,N_4183);
nor U4386 (N_4386,N_4063,N_4225);
xnor U4387 (N_4387,N_4076,N_4233);
and U4388 (N_4388,N_4249,N_4190);
nand U4389 (N_4389,N_4162,N_4187);
nor U4390 (N_4390,N_4149,N_4221);
nor U4391 (N_4391,N_4093,N_4050);
and U4392 (N_4392,N_4048,N_4059);
and U4393 (N_4393,N_4052,N_4212);
or U4394 (N_4394,N_4140,N_4021);
and U4395 (N_4395,N_4094,N_4220);
nor U4396 (N_4396,N_4084,N_4114);
nand U4397 (N_4397,N_4045,N_4249);
nor U4398 (N_4398,N_4197,N_4007);
nand U4399 (N_4399,N_4188,N_4126);
or U4400 (N_4400,N_4196,N_4013);
or U4401 (N_4401,N_4234,N_4058);
nand U4402 (N_4402,N_4100,N_4135);
and U4403 (N_4403,N_4217,N_4160);
or U4404 (N_4404,N_4191,N_4173);
and U4405 (N_4405,N_4162,N_4201);
nand U4406 (N_4406,N_4146,N_4217);
xor U4407 (N_4407,N_4032,N_4168);
nand U4408 (N_4408,N_4183,N_4095);
or U4409 (N_4409,N_4177,N_4145);
nand U4410 (N_4410,N_4022,N_4050);
and U4411 (N_4411,N_4092,N_4236);
and U4412 (N_4412,N_4155,N_4167);
nor U4413 (N_4413,N_4142,N_4181);
nor U4414 (N_4414,N_4008,N_4246);
nand U4415 (N_4415,N_4015,N_4084);
or U4416 (N_4416,N_4191,N_4131);
nand U4417 (N_4417,N_4110,N_4092);
nor U4418 (N_4418,N_4141,N_4066);
or U4419 (N_4419,N_4062,N_4036);
nand U4420 (N_4420,N_4160,N_4134);
and U4421 (N_4421,N_4132,N_4225);
or U4422 (N_4422,N_4227,N_4249);
nor U4423 (N_4423,N_4077,N_4138);
nand U4424 (N_4424,N_4054,N_4202);
or U4425 (N_4425,N_4065,N_4088);
nand U4426 (N_4426,N_4235,N_4148);
and U4427 (N_4427,N_4157,N_4004);
or U4428 (N_4428,N_4214,N_4240);
nor U4429 (N_4429,N_4187,N_4182);
nand U4430 (N_4430,N_4026,N_4244);
nor U4431 (N_4431,N_4193,N_4074);
nor U4432 (N_4432,N_4149,N_4227);
nor U4433 (N_4433,N_4100,N_4019);
nor U4434 (N_4434,N_4060,N_4091);
or U4435 (N_4435,N_4190,N_4231);
nor U4436 (N_4436,N_4200,N_4165);
and U4437 (N_4437,N_4213,N_4202);
nand U4438 (N_4438,N_4010,N_4062);
nand U4439 (N_4439,N_4232,N_4043);
or U4440 (N_4440,N_4062,N_4193);
nor U4441 (N_4441,N_4134,N_4149);
and U4442 (N_4442,N_4209,N_4236);
and U4443 (N_4443,N_4210,N_4172);
xnor U4444 (N_4444,N_4169,N_4073);
and U4445 (N_4445,N_4001,N_4004);
and U4446 (N_4446,N_4080,N_4167);
nor U4447 (N_4447,N_4026,N_4062);
nor U4448 (N_4448,N_4238,N_4053);
nand U4449 (N_4449,N_4153,N_4011);
nand U4450 (N_4450,N_4239,N_4005);
nand U4451 (N_4451,N_4024,N_4192);
xnor U4452 (N_4452,N_4164,N_4030);
xor U4453 (N_4453,N_4109,N_4229);
and U4454 (N_4454,N_4061,N_4223);
and U4455 (N_4455,N_4236,N_4245);
or U4456 (N_4456,N_4133,N_4244);
nor U4457 (N_4457,N_4026,N_4212);
or U4458 (N_4458,N_4089,N_4051);
or U4459 (N_4459,N_4042,N_4108);
or U4460 (N_4460,N_4076,N_4151);
or U4461 (N_4461,N_4195,N_4187);
and U4462 (N_4462,N_4059,N_4154);
and U4463 (N_4463,N_4129,N_4085);
nand U4464 (N_4464,N_4110,N_4072);
nand U4465 (N_4465,N_4038,N_4227);
nor U4466 (N_4466,N_4122,N_4152);
nor U4467 (N_4467,N_4199,N_4114);
or U4468 (N_4468,N_4047,N_4183);
nor U4469 (N_4469,N_4091,N_4198);
nor U4470 (N_4470,N_4083,N_4181);
nand U4471 (N_4471,N_4024,N_4227);
nor U4472 (N_4472,N_4011,N_4077);
or U4473 (N_4473,N_4122,N_4046);
or U4474 (N_4474,N_4075,N_4150);
and U4475 (N_4475,N_4155,N_4052);
xnor U4476 (N_4476,N_4236,N_4135);
or U4477 (N_4477,N_4147,N_4010);
nand U4478 (N_4478,N_4173,N_4194);
xor U4479 (N_4479,N_4065,N_4183);
and U4480 (N_4480,N_4091,N_4246);
nand U4481 (N_4481,N_4164,N_4132);
and U4482 (N_4482,N_4087,N_4180);
or U4483 (N_4483,N_4197,N_4223);
nor U4484 (N_4484,N_4204,N_4061);
nand U4485 (N_4485,N_4069,N_4040);
or U4486 (N_4486,N_4067,N_4144);
xnor U4487 (N_4487,N_4214,N_4122);
or U4488 (N_4488,N_4055,N_4111);
nor U4489 (N_4489,N_4120,N_4031);
or U4490 (N_4490,N_4061,N_4095);
nor U4491 (N_4491,N_4084,N_4228);
nand U4492 (N_4492,N_4116,N_4182);
nand U4493 (N_4493,N_4136,N_4048);
nand U4494 (N_4494,N_4013,N_4151);
nor U4495 (N_4495,N_4009,N_4051);
nor U4496 (N_4496,N_4091,N_4015);
nor U4497 (N_4497,N_4167,N_4025);
xnor U4498 (N_4498,N_4019,N_4142);
nand U4499 (N_4499,N_4161,N_4187);
or U4500 (N_4500,N_4485,N_4285);
and U4501 (N_4501,N_4413,N_4422);
nand U4502 (N_4502,N_4450,N_4351);
or U4503 (N_4503,N_4256,N_4324);
xnor U4504 (N_4504,N_4475,N_4266);
nand U4505 (N_4505,N_4339,N_4439);
nand U4506 (N_4506,N_4499,N_4269);
xor U4507 (N_4507,N_4265,N_4434);
nor U4508 (N_4508,N_4489,N_4441);
or U4509 (N_4509,N_4299,N_4410);
or U4510 (N_4510,N_4471,N_4494);
nand U4511 (N_4511,N_4397,N_4393);
and U4512 (N_4512,N_4480,N_4261);
xnor U4513 (N_4513,N_4257,N_4315);
nor U4514 (N_4514,N_4334,N_4448);
or U4515 (N_4515,N_4469,N_4286);
nor U4516 (N_4516,N_4320,N_4323);
or U4517 (N_4517,N_4426,N_4496);
and U4518 (N_4518,N_4411,N_4470);
xor U4519 (N_4519,N_4287,N_4417);
nand U4520 (N_4520,N_4355,N_4486);
or U4521 (N_4521,N_4383,N_4384);
and U4522 (N_4522,N_4298,N_4457);
nor U4523 (N_4523,N_4389,N_4466);
or U4524 (N_4524,N_4318,N_4380);
or U4525 (N_4525,N_4372,N_4376);
nand U4526 (N_4526,N_4278,N_4447);
and U4527 (N_4527,N_4419,N_4365);
or U4528 (N_4528,N_4373,N_4359);
nand U4529 (N_4529,N_4487,N_4335);
nor U4530 (N_4530,N_4392,N_4282);
xnor U4531 (N_4531,N_4474,N_4444);
nor U4532 (N_4532,N_4483,N_4456);
or U4533 (N_4533,N_4264,N_4352);
nand U4534 (N_4534,N_4319,N_4275);
nor U4535 (N_4535,N_4348,N_4293);
or U4536 (N_4536,N_4405,N_4387);
and U4537 (N_4537,N_4307,N_4368);
or U4538 (N_4538,N_4342,N_4358);
nand U4539 (N_4539,N_4325,N_4349);
nor U4540 (N_4540,N_4375,N_4311);
nand U4541 (N_4541,N_4366,N_4316);
nor U4542 (N_4542,N_4304,N_4404);
nor U4543 (N_4543,N_4436,N_4347);
nor U4544 (N_4544,N_4403,N_4367);
and U4545 (N_4545,N_4271,N_4267);
and U4546 (N_4546,N_4343,N_4421);
and U4547 (N_4547,N_4260,N_4498);
nand U4548 (N_4548,N_4473,N_4378);
nor U4549 (N_4549,N_4381,N_4326);
nor U4550 (N_4550,N_4251,N_4440);
and U4551 (N_4551,N_4479,N_4361);
xnor U4552 (N_4552,N_4350,N_4294);
and U4553 (N_4553,N_4445,N_4467);
nor U4554 (N_4554,N_4341,N_4482);
xnor U4555 (N_4555,N_4452,N_4281);
nor U4556 (N_4556,N_4296,N_4263);
nand U4557 (N_4557,N_4492,N_4396);
nand U4558 (N_4558,N_4306,N_4254);
or U4559 (N_4559,N_4284,N_4394);
nor U4560 (N_4560,N_4461,N_4331);
or U4561 (N_4561,N_4274,N_4344);
and U4562 (N_4562,N_4289,N_4356);
or U4563 (N_4563,N_4478,N_4268);
xnor U4564 (N_4564,N_4451,N_4462);
and U4565 (N_4565,N_4449,N_4333);
or U4566 (N_4566,N_4357,N_4338);
xor U4567 (N_4567,N_4493,N_4377);
or U4568 (N_4568,N_4312,N_4438);
and U4569 (N_4569,N_4385,N_4250);
or U4570 (N_4570,N_4458,N_4363);
nand U4571 (N_4571,N_4321,N_4277);
and U4572 (N_4572,N_4488,N_4424);
xnor U4573 (N_4573,N_4437,N_4313);
nand U4574 (N_4574,N_4330,N_4481);
or U4575 (N_4575,N_4453,N_4255);
xnor U4576 (N_4576,N_4336,N_4310);
or U4577 (N_4577,N_4252,N_4272);
and U4578 (N_4578,N_4362,N_4290);
and U4579 (N_4579,N_4346,N_4300);
nand U4580 (N_4580,N_4322,N_4433);
nand U4581 (N_4581,N_4412,N_4476);
and U4582 (N_4582,N_4429,N_4371);
nand U4583 (N_4583,N_4420,N_4345);
or U4584 (N_4584,N_4409,N_4288);
nand U4585 (N_4585,N_4314,N_4390);
nand U4586 (N_4586,N_4354,N_4491);
and U4587 (N_4587,N_4295,N_4425);
nand U4588 (N_4588,N_4364,N_4305);
xnor U4589 (N_4589,N_4262,N_4414);
or U4590 (N_4590,N_4446,N_4465);
or U4591 (N_4591,N_4353,N_4431);
or U4592 (N_4592,N_4497,N_4276);
or U4593 (N_4593,N_4279,N_4291);
nor U4594 (N_4594,N_4484,N_4297);
and U4595 (N_4595,N_4443,N_4283);
and U4596 (N_4596,N_4435,N_4407);
nand U4597 (N_4597,N_4253,N_4270);
xor U4598 (N_4598,N_4460,N_4442);
and U4599 (N_4599,N_4309,N_4428);
nand U4600 (N_4600,N_4401,N_4463);
and U4601 (N_4601,N_4454,N_4301);
or U4602 (N_4602,N_4292,N_4340);
or U4603 (N_4603,N_4402,N_4370);
nand U4604 (N_4604,N_4382,N_4406);
or U4605 (N_4605,N_4386,N_4399);
nand U4606 (N_4606,N_4369,N_4459);
and U4607 (N_4607,N_4388,N_4302);
and U4608 (N_4608,N_4415,N_4280);
xnor U4609 (N_4609,N_4379,N_4408);
nor U4610 (N_4610,N_4317,N_4398);
nand U4611 (N_4611,N_4332,N_4400);
or U4612 (N_4612,N_4430,N_4391);
and U4613 (N_4613,N_4495,N_4360);
nand U4614 (N_4614,N_4395,N_4416);
or U4615 (N_4615,N_4468,N_4464);
and U4616 (N_4616,N_4259,N_4328);
nand U4617 (N_4617,N_4472,N_4477);
and U4618 (N_4618,N_4374,N_4308);
or U4619 (N_4619,N_4337,N_4329);
or U4620 (N_4620,N_4303,N_4455);
xnor U4621 (N_4621,N_4423,N_4327);
and U4622 (N_4622,N_4427,N_4258);
and U4623 (N_4623,N_4432,N_4418);
nor U4624 (N_4624,N_4490,N_4273);
and U4625 (N_4625,N_4402,N_4489);
nand U4626 (N_4626,N_4377,N_4482);
or U4627 (N_4627,N_4470,N_4271);
xor U4628 (N_4628,N_4478,N_4307);
and U4629 (N_4629,N_4368,N_4277);
or U4630 (N_4630,N_4392,N_4483);
xnor U4631 (N_4631,N_4343,N_4266);
nand U4632 (N_4632,N_4255,N_4308);
nand U4633 (N_4633,N_4439,N_4260);
and U4634 (N_4634,N_4460,N_4373);
or U4635 (N_4635,N_4402,N_4455);
and U4636 (N_4636,N_4285,N_4288);
or U4637 (N_4637,N_4255,N_4355);
or U4638 (N_4638,N_4470,N_4444);
nand U4639 (N_4639,N_4373,N_4422);
or U4640 (N_4640,N_4449,N_4301);
nand U4641 (N_4641,N_4433,N_4289);
or U4642 (N_4642,N_4308,N_4468);
or U4643 (N_4643,N_4385,N_4369);
or U4644 (N_4644,N_4359,N_4341);
nor U4645 (N_4645,N_4482,N_4378);
nand U4646 (N_4646,N_4279,N_4365);
and U4647 (N_4647,N_4286,N_4307);
nor U4648 (N_4648,N_4301,N_4428);
nand U4649 (N_4649,N_4482,N_4328);
nand U4650 (N_4650,N_4386,N_4318);
or U4651 (N_4651,N_4460,N_4377);
nor U4652 (N_4652,N_4307,N_4425);
and U4653 (N_4653,N_4417,N_4261);
nor U4654 (N_4654,N_4285,N_4356);
nand U4655 (N_4655,N_4493,N_4369);
and U4656 (N_4656,N_4310,N_4358);
and U4657 (N_4657,N_4264,N_4251);
nand U4658 (N_4658,N_4446,N_4456);
xnor U4659 (N_4659,N_4343,N_4481);
nor U4660 (N_4660,N_4446,N_4412);
and U4661 (N_4661,N_4388,N_4297);
and U4662 (N_4662,N_4341,N_4477);
nor U4663 (N_4663,N_4331,N_4407);
nor U4664 (N_4664,N_4299,N_4387);
xnor U4665 (N_4665,N_4266,N_4362);
nor U4666 (N_4666,N_4435,N_4430);
and U4667 (N_4667,N_4384,N_4399);
nor U4668 (N_4668,N_4486,N_4452);
xor U4669 (N_4669,N_4447,N_4462);
nor U4670 (N_4670,N_4495,N_4440);
xnor U4671 (N_4671,N_4358,N_4296);
or U4672 (N_4672,N_4317,N_4484);
nor U4673 (N_4673,N_4349,N_4429);
or U4674 (N_4674,N_4486,N_4481);
nand U4675 (N_4675,N_4278,N_4448);
nand U4676 (N_4676,N_4446,N_4403);
xnor U4677 (N_4677,N_4460,N_4459);
or U4678 (N_4678,N_4429,N_4347);
or U4679 (N_4679,N_4336,N_4268);
xnor U4680 (N_4680,N_4468,N_4274);
and U4681 (N_4681,N_4250,N_4439);
xor U4682 (N_4682,N_4336,N_4382);
xnor U4683 (N_4683,N_4414,N_4259);
nor U4684 (N_4684,N_4322,N_4255);
nand U4685 (N_4685,N_4324,N_4314);
nor U4686 (N_4686,N_4291,N_4254);
nor U4687 (N_4687,N_4356,N_4310);
and U4688 (N_4688,N_4357,N_4442);
nand U4689 (N_4689,N_4393,N_4408);
or U4690 (N_4690,N_4457,N_4283);
nor U4691 (N_4691,N_4397,N_4313);
nand U4692 (N_4692,N_4290,N_4352);
nand U4693 (N_4693,N_4308,N_4254);
nor U4694 (N_4694,N_4346,N_4379);
nor U4695 (N_4695,N_4364,N_4427);
xor U4696 (N_4696,N_4286,N_4403);
and U4697 (N_4697,N_4484,N_4343);
and U4698 (N_4698,N_4369,N_4452);
xnor U4699 (N_4699,N_4391,N_4310);
nor U4700 (N_4700,N_4365,N_4328);
and U4701 (N_4701,N_4430,N_4257);
nand U4702 (N_4702,N_4330,N_4400);
nand U4703 (N_4703,N_4468,N_4461);
or U4704 (N_4704,N_4429,N_4271);
nand U4705 (N_4705,N_4365,N_4343);
and U4706 (N_4706,N_4395,N_4360);
nand U4707 (N_4707,N_4339,N_4458);
and U4708 (N_4708,N_4252,N_4359);
nor U4709 (N_4709,N_4449,N_4337);
or U4710 (N_4710,N_4325,N_4293);
and U4711 (N_4711,N_4446,N_4307);
nand U4712 (N_4712,N_4347,N_4270);
or U4713 (N_4713,N_4437,N_4322);
or U4714 (N_4714,N_4348,N_4466);
or U4715 (N_4715,N_4434,N_4360);
and U4716 (N_4716,N_4380,N_4309);
and U4717 (N_4717,N_4475,N_4430);
xnor U4718 (N_4718,N_4278,N_4445);
and U4719 (N_4719,N_4399,N_4471);
and U4720 (N_4720,N_4313,N_4270);
and U4721 (N_4721,N_4255,N_4337);
or U4722 (N_4722,N_4428,N_4305);
or U4723 (N_4723,N_4490,N_4494);
nor U4724 (N_4724,N_4472,N_4402);
xnor U4725 (N_4725,N_4325,N_4412);
or U4726 (N_4726,N_4348,N_4481);
xor U4727 (N_4727,N_4423,N_4413);
and U4728 (N_4728,N_4324,N_4461);
and U4729 (N_4729,N_4301,N_4295);
nor U4730 (N_4730,N_4280,N_4481);
xnor U4731 (N_4731,N_4370,N_4335);
nor U4732 (N_4732,N_4313,N_4382);
nor U4733 (N_4733,N_4365,N_4494);
xnor U4734 (N_4734,N_4349,N_4437);
nand U4735 (N_4735,N_4314,N_4389);
or U4736 (N_4736,N_4409,N_4492);
or U4737 (N_4737,N_4380,N_4483);
nand U4738 (N_4738,N_4254,N_4345);
and U4739 (N_4739,N_4344,N_4337);
or U4740 (N_4740,N_4339,N_4284);
and U4741 (N_4741,N_4258,N_4489);
or U4742 (N_4742,N_4352,N_4401);
or U4743 (N_4743,N_4429,N_4353);
or U4744 (N_4744,N_4419,N_4376);
and U4745 (N_4745,N_4419,N_4379);
nand U4746 (N_4746,N_4386,N_4398);
and U4747 (N_4747,N_4326,N_4469);
or U4748 (N_4748,N_4321,N_4436);
nand U4749 (N_4749,N_4376,N_4349);
or U4750 (N_4750,N_4543,N_4698);
nor U4751 (N_4751,N_4616,N_4576);
xnor U4752 (N_4752,N_4665,N_4512);
nand U4753 (N_4753,N_4714,N_4650);
or U4754 (N_4754,N_4710,N_4505);
nor U4755 (N_4755,N_4675,N_4737);
xnor U4756 (N_4756,N_4708,N_4571);
or U4757 (N_4757,N_4730,N_4717);
or U4758 (N_4758,N_4615,N_4600);
nor U4759 (N_4759,N_4736,N_4645);
and U4760 (N_4760,N_4527,N_4646);
and U4761 (N_4761,N_4703,N_4555);
nand U4762 (N_4762,N_4726,N_4599);
nor U4763 (N_4763,N_4643,N_4729);
xnor U4764 (N_4764,N_4740,N_4502);
or U4765 (N_4765,N_4504,N_4719);
and U4766 (N_4766,N_4677,N_4634);
and U4767 (N_4767,N_4689,N_4607);
nor U4768 (N_4768,N_4545,N_4541);
nor U4769 (N_4769,N_4559,N_4687);
or U4770 (N_4770,N_4733,N_4612);
nand U4771 (N_4771,N_4585,N_4518);
nand U4772 (N_4772,N_4566,N_4657);
or U4773 (N_4773,N_4648,N_4627);
or U4774 (N_4774,N_4619,N_4704);
nand U4775 (N_4775,N_4651,N_4696);
and U4776 (N_4776,N_4604,N_4538);
and U4777 (N_4777,N_4635,N_4606);
nor U4778 (N_4778,N_4629,N_4716);
and U4779 (N_4779,N_4613,N_4514);
or U4780 (N_4780,N_4544,N_4558);
and U4781 (N_4781,N_4638,N_4633);
and U4782 (N_4782,N_4739,N_4735);
nor U4783 (N_4783,N_4745,N_4670);
nor U4784 (N_4784,N_4702,N_4659);
nand U4785 (N_4785,N_4524,N_4586);
or U4786 (N_4786,N_4682,N_4501);
xnor U4787 (N_4787,N_4513,N_4692);
or U4788 (N_4788,N_4690,N_4529);
nor U4789 (N_4789,N_4738,N_4582);
or U4790 (N_4790,N_4723,N_4637);
nand U4791 (N_4791,N_4685,N_4562);
nand U4792 (N_4792,N_4668,N_4746);
and U4793 (N_4793,N_4626,N_4727);
nor U4794 (N_4794,N_4741,N_4556);
xnor U4795 (N_4795,N_4591,N_4721);
or U4796 (N_4796,N_4695,N_4597);
nand U4797 (N_4797,N_4601,N_4749);
or U4798 (N_4798,N_4530,N_4706);
nand U4799 (N_4799,N_4628,N_4532);
nor U4800 (N_4800,N_4551,N_4713);
nand U4801 (N_4801,N_4728,N_4691);
nand U4802 (N_4802,N_4693,N_4681);
or U4803 (N_4803,N_4655,N_4580);
and U4804 (N_4804,N_4653,N_4622);
xor U4805 (N_4805,N_4644,N_4718);
and U4806 (N_4806,N_4503,N_4508);
nor U4807 (N_4807,N_4656,N_4570);
and U4808 (N_4808,N_4587,N_4525);
or U4809 (N_4809,N_4747,N_4589);
nor U4810 (N_4810,N_4724,N_4748);
or U4811 (N_4811,N_4520,N_4715);
nand U4812 (N_4812,N_4534,N_4678);
nor U4813 (N_4813,N_4672,N_4709);
nand U4814 (N_4814,N_4535,N_4575);
nor U4815 (N_4815,N_4602,N_4642);
or U4816 (N_4816,N_4517,N_4515);
nand U4817 (N_4817,N_4528,N_4707);
nor U4818 (N_4818,N_4554,N_4577);
nor U4819 (N_4819,N_4509,N_4531);
nor U4820 (N_4820,N_4614,N_4547);
or U4821 (N_4821,N_4674,N_4595);
and U4822 (N_4822,N_4550,N_4663);
nand U4823 (N_4823,N_4609,N_4632);
nand U4824 (N_4824,N_4557,N_4673);
nor U4825 (N_4825,N_4583,N_4500);
nor U4826 (N_4826,N_4639,N_4573);
or U4827 (N_4827,N_4636,N_4537);
xnor U4828 (N_4828,N_4744,N_4565);
nand U4829 (N_4829,N_4567,N_4722);
and U4830 (N_4830,N_4631,N_4608);
and U4831 (N_4831,N_4590,N_4523);
nand U4832 (N_4832,N_4679,N_4579);
or U4833 (N_4833,N_4712,N_4664);
and U4834 (N_4834,N_4568,N_4688);
xor U4835 (N_4835,N_4623,N_4521);
nand U4836 (N_4836,N_4526,N_4546);
nor U4837 (N_4837,N_4540,N_4519);
or U4838 (N_4838,N_4564,N_4676);
nand U4839 (N_4839,N_4711,N_4683);
or U4840 (N_4840,N_4552,N_4617);
nor U4841 (N_4841,N_4572,N_4596);
and U4842 (N_4842,N_4720,N_4611);
nor U4843 (N_4843,N_4666,N_4732);
nor U4844 (N_4844,N_4743,N_4701);
xnor U4845 (N_4845,N_4694,N_4671);
or U4846 (N_4846,N_4680,N_4603);
and U4847 (N_4847,N_4511,N_4584);
or U4848 (N_4848,N_4621,N_4658);
nand U4849 (N_4849,N_4667,N_4620);
xnor U4850 (N_4850,N_4507,N_4588);
and U4851 (N_4851,N_4539,N_4731);
or U4852 (N_4852,N_4592,N_4578);
xnor U4853 (N_4853,N_4549,N_4574);
nor U4854 (N_4854,N_4700,N_4533);
nor U4855 (N_4855,N_4686,N_4605);
xnor U4856 (N_4856,N_4536,N_4593);
nor U4857 (N_4857,N_4705,N_4624);
xnor U4858 (N_4858,N_4641,N_4506);
nor U4859 (N_4859,N_4684,N_4560);
xor U4860 (N_4860,N_4640,N_4625);
nand U4861 (N_4861,N_4581,N_4662);
or U4862 (N_4862,N_4742,N_4652);
nand U4863 (N_4863,N_4516,N_4598);
nor U4864 (N_4864,N_4734,N_4610);
nor U4865 (N_4865,N_4561,N_4654);
and U4866 (N_4866,N_4594,N_4661);
and U4867 (N_4867,N_4542,N_4553);
or U4868 (N_4868,N_4660,N_4569);
and U4869 (N_4869,N_4647,N_4630);
nand U4870 (N_4870,N_4548,N_4725);
nand U4871 (N_4871,N_4522,N_4669);
or U4872 (N_4872,N_4510,N_4697);
and U4873 (N_4873,N_4699,N_4618);
or U4874 (N_4874,N_4563,N_4649);
and U4875 (N_4875,N_4528,N_4618);
or U4876 (N_4876,N_4713,N_4517);
nor U4877 (N_4877,N_4691,N_4588);
nor U4878 (N_4878,N_4567,N_4725);
nand U4879 (N_4879,N_4693,N_4503);
nor U4880 (N_4880,N_4578,N_4702);
nor U4881 (N_4881,N_4599,N_4578);
or U4882 (N_4882,N_4552,N_4619);
nor U4883 (N_4883,N_4691,N_4514);
xnor U4884 (N_4884,N_4675,N_4612);
or U4885 (N_4885,N_4674,N_4618);
nand U4886 (N_4886,N_4501,N_4624);
nand U4887 (N_4887,N_4608,N_4500);
nand U4888 (N_4888,N_4699,N_4628);
nor U4889 (N_4889,N_4534,N_4684);
nand U4890 (N_4890,N_4623,N_4663);
and U4891 (N_4891,N_4528,N_4594);
or U4892 (N_4892,N_4514,N_4660);
or U4893 (N_4893,N_4605,N_4691);
and U4894 (N_4894,N_4527,N_4699);
nand U4895 (N_4895,N_4698,N_4572);
nand U4896 (N_4896,N_4691,N_4733);
nand U4897 (N_4897,N_4612,N_4702);
nor U4898 (N_4898,N_4547,N_4645);
nand U4899 (N_4899,N_4700,N_4607);
or U4900 (N_4900,N_4741,N_4692);
or U4901 (N_4901,N_4616,N_4555);
nand U4902 (N_4902,N_4522,N_4746);
or U4903 (N_4903,N_4569,N_4500);
and U4904 (N_4904,N_4680,N_4722);
xnor U4905 (N_4905,N_4635,N_4702);
nand U4906 (N_4906,N_4594,N_4653);
nor U4907 (N_4907,N_4546,N_4746);
nor U4908 (N_4908,N_4703,N_4574);
nand U4909 (N_4909,N_4680,N_4706);
or U4910 (N_4910,N_4592,N_4544);
and U4911 (N_4911,N_4621,N_4542);
nor U4912 (N_4912,N_4568,N_4541);
and U4913 (N_4913,N_4693,N_4631);
xnor U4914 (N_4914,N_4620,N_4599);
and U4915 (N_4915,N_4670,N_4631);
nand U4916 (N_4916,N_4514,N_4569);
or U4917 (N_4917,N_4716,N_4508);
nand U4918 (N_4918,N_4744,N_4685);
or U4919 (N_4919,N_4583,N_4659);
nand U4920 (N_4920,N_4527,N_4587);
xor U4921 (N_4921,N_4732,N_4582);
and U4922 (N_4922,N_4527,N_4593);
or U4923 (N_4923,N_4716,N_4660);
and U4924 (N_4924,N_4667,N_4645);
nor U4925 (N_4925,N_4554,N_4650);
nor U4926 (N_4926,N_4506,N_4604);
and U4927 (N_4927,N_4590,N_4742);
nor U4928 (N_4928,N_4501,N_4617);
nor U4929 (N_4929,N_4562,N_4704);
nor U4930 (N_4930,N_4633,N_4505);
or U4931 (N_4931,N_4640,N_4746);
and U4932 (N_4932,N_4644,N_4530);
or U4933 (N_4933,N_4644,N_4689);
nand U4934 (N_4934,N_4502,N_4562);
and U4935 (N_4935,N_4603,N_4674);
and U4936 (N_4936,N_4658,N_4618);
nand U4937 (N_4937,N_4586,N_4569);
xnor U4938 (N_4938,N_4679,N_4728);
nand U4939 (N_4939,N_4682,N_4579);
nand U4940 (N_4940,N_4650,N_4743);
xor U4941 (N_4941,N_4697,N_4747);
and U4942 (N_4942,N_4691,N_4659);
or U4943 (N_4943,N_4737,N_4656);
or U4944 (N_4944,N_4644,N_4557);
nand U4945 (N_4945,N_4675,N_4517);
or U4946 (N_4946,N_4671,N_4670);
xor U4947 (N_4947,N_4517,N_4593);
nor U4948 (N_4948,N_4640,N_4529);
or U4949 (N_4949,N_4521,N_4708);
nor U4950 (N_4950,N_4543,N_4681);
xor U4951 (N_4951,N_4692,N_4506);
nand U4952 (N_4952,N_4562,N_4693);
nand U4953 (N_4953,N_4517,N_4742);
nand U4954 (N_4954,N_4626,N_4659);
and U4955 (N_4955,N_4624,N_4591);
and U4956 (N_4956,N_4706,N_4621);
or U4957 (N_4957,N_4565,N_4518);
and U4958 (N_4958,N_4742,N_4552);
and U4959 (N_4959,N_4634,N_4562);
nor U4960 (N_4960,N_4536,N_4658);
or U4961 (N_4961,N_4700,N_4507);
or U4962 (N_4962,N_4725,N_4731);
or U4963 (N_4963,N_4600,N_4683);
or U4964 (N_4964,N_4558,N_4512);
xnor U4965 (N_4965,N_4641,N_4743);
nor U4966 (N_4966,N_4587,N_4543);
and U4967 (N_4967,N_4686,N_4699);
nand U4968 (N_4968,N_4532,N_4593);
and U4969 (N_4969,N_4629,N_4731);
nand U4970 (N_4970,N_4622,N_4525);
nor U4971 (N_4971,N_4587,N_4610);
xnor U4972 (N_4972,N_4575,N_4652);
or U4973 (N_4973,N_4740,N_4630);
and U4974 (N_4974,N_4522,N_4623);
and U4975 (N_4975,N_4713,N_4685);
and U4976 (N_4976,N_4681,N_4671);
or U4977 (N_4977,N_4547,N_4626);
nor U4978 (N_4978,N_4671,N_4561);
nor U4979 (N_4979,N_4548,N_4550);
or U4980 (N_4980,N_4657,N_4665);
or U4981 (N_4981,N_4685,N_4530);
nand U4982 (N_4982,N_4629,N_4517);
nor U4983 (N_4983,N_4716,N_4605);
nor U4984 (N_4984,N_4711,N_4515);
and U4985 (N_4985,N_4632,N_4589);
xnor U4986 (N_4986,N_4565,N_4721);
nand U4987 (N_4987,N_4582,N_4573);
nor U4988 (N_4988,N_4680,N_4562);
and U4989 (N_4989,N_4738,N_4697);
or U4990 (N_4990,N_4530,N_4637);
xnor U4991 (N_4991,N_4612,N_4516);
nand U4992 (N_4992,N_4714,N_4568);
and U4993 (N_4993,N_4702,N_4506);
nand U4994 (N_4994,N_4558,N_4580);
or U4995 (N_4995,N_4607,N_4615);
nand U4996 (N_4996,N_4589,N_4717);
or U4997 (N_4997,N_4634,N_4500);
nor U4998 (N_4998,N_4597,N_4596);
xor U4999 (N_4999,N_4551,N_4696);
or U5000 (N_5000,N_4881,N_4750);
nand U5001 (N_5001,N_4890,N_4979);
and U5002 (N_5002,N_4771,N_4836);
nand U5003 (N_5003,N_4989,N_4948);
nand U5004 (N_5004,N_4752,N_4903);
or U5005 (N_5005,N_4849,N_4869);
and U5006 (N_5006,N_4764,N_4974);
nor U5007 (N_5007,N_4780,N_4787);
nand U5008 (N_5008,N_4972,N_4843);
or U5009 (N_5009,N_4969,N_4908);
nor U5010 (N_5010,N_4861,N_4916);
xnor U5011 (N_5011,N_4818,N_4924);
and U5012 (N_5012,N_4839,N_4844);
or U5013 (N_5013,N_4954,N_4958);
nor U5014 (N_5014,N_4788,N_4939);
nand U5015 (N_5015,N_4860,N_4819);
or U5016 (N_5016,N_4810,N_4877);
nor U5017 (N_5017,N_4963,N_4929);
nor U5018 (N_5018,N_4811,N_4902);
nor U5019 (N_5019,N_4817,N_4895);
nor U5020 (N_5020,N_4837,N_4891);
or U5021 (N_5021,N_4892,N_4915);
or U5022 (N_5022,N_4883,N_4893);
nor U5023 (N_5023,N_4997,N_4921);
or U5024 (N_5024,N_4941,N_4982);
or U5025 (N_5025,N_4857,N_4832);
and U5026 (N_5026,N_4953,N_4812);
nor U5027 (N_5027,N_4770,N_4785);
and U5028 (N_5028,N_4964,N_4826);
xor U5029 (N_5029,N_4774,N_4793);
or U5030 (N_5030,N_4835,N_4907);
or U5031 (N_5031,N_4971,N_4962);
nand U5032 (N_5032,N_4957,N_4886);
nand U5033 (N_5033,N_4876,N_4808);
nand U5034 (N_5034,N_4760,N_4938);
or U5035 (N_5035,N_4758,N_4859);
and U5036 (N_5036,N_4807,N_4914);
or U5037 (N_5037,N_4961,N_4782);
or U5038 (N_5038,N_4933,N_4983);
nand U5039 (N_5039,N_4755,N_4910);
nor U5040 (N_5040,N_4875,N_4970);
or U5041 (N_5041,N_4827,N_4845);
nor U5042 (N_5042,N_4896,N_4772);
nand U5043 (N_5043,N_4798,N_4757);
and U5044 (N_5044,N_4888,N_4887);
or U5045 (N_5045,N_4976,N_4816);
nand U5046 (N_5046,N_4978,N_4911);
nor U5047 (N_5047,N_4791,N_4765);
nor U5048 (N_5048,N_4966,N_4841);
nor U5049 (N_5049,N_4851,N_4922);
nor U5050 (N_5050,N_4980,N_4850);
and U5051 (N_5051,N_4942,N_4863);
and U5052 (N_5052,N_4824,N_4873);
nand U5053 (N_5053,N_4799,N_4786);
nor U5054 (N_5054,N_4838,N_4777);
and U5055 (N_5055,N_4947,N_4898);
nand U5056 (N_5056,N_4952,N_4813);
xnor U5057 (N_5057,N_4862,N_4889);
and U5058 (N_5058,N_4936,N_4790);
nor U5059 (N_5059,N_4856,N_4965);
and U5060 (N_5060,N_4829,N_4759);
nor U5061 (N_5061,N_4783,N_4925);
xor U5062 (N_5062,N_4918,N_4993);
or U5063 (N_5063,N_4998,N_4804);
or U5064 (N_5064,N_4882,N_4801);
nor U5065 (N_5065,N_4854,N_4814);
xnor U5066 (N_5066,N_4761,N_4830);
xor U5067 (N_5067,N_4754,N_4930);
nand U5068 (N_5068,N_4934,N_4919);
nand U5069 (N_5069,N_4773,N_4950);
nor U5070 (N_5070,N_4840,N_4913);
and U5071 (N_5071,N_4951,N_4956);
or U5072 (N_5072,N_4937,N_4864);
nor U5073 (N_5073,N_4946,N_4763);
nand U5074 (N_5074,N_4795,N_4995);
nor U5075 (N_5075,N_4868,N_4825);
or U5076 (N_5076,N_4821,N_4943);
nor U5077 (N_5077,N_4996,N_4940);
or U5078 (N_5078,N_4977,N_4847);
xor U5079 (N_5079,N_4884,N_4762);
and U5080 (N_5080,N_4784,N_4809);
or U5081 (N_5081,N_4944,N_4778);
nand U5082 (N_5082,N_4990,N_4899);
or U5083 (N_5083,N_4945,N_4949);
xor U5084 (N_5084,N_4988,N_4794);
xor U5085 (N_5085,N_4855,N_4905);
nor U5086 (N_5086,N_4828,N_4792);
nand U5087 (N_5087,N_4960,N_4986);
or U5088 (N_5088,N_4833,N_4897);
nor U5089 (N_5089,N_4879,N_4789);
nor U5090 (N_5090,N_4858,N_4806);
xor U5091 (N_5091,N_4834,N_4871);
or U5092 (N_5092,N_4823,N_4959);
nand U5093 (N_5093,N_4797,N_4932);
nand U5094 (N_5094,N_4776,N_4955);
and U5095 (N_5095,N_4878,N_4874);
and U5096 (N_5096,N_4867,N_4923);
and U5097 (N_5097,N_4842,N_4853);
nor U5098 (N_5098,N_4901,N_4900);
nand U5099 (N_5099,N_4767,N_4894);
or U5100 (N_5100,N_4865,N_4831);
and U5101 (N_5101,N_4815,N_4775);
nor U5102 (N_5102,N_4751,N_4909);
xor U5103 (N_5103,N_4846,N_4968);
nand U5104 (N_5104,N_4880,N_4927);
and U5105 (N_5105,N_4753,N_4768);
nor U5106 (N_5106,N_4992,N_4999);
and U5107 (N_5107,N_4928,N_4852);
or U5108 (N_5108,N_4866,N_4904);
or U5109 (N_5109,N_4872,N_4984);
or U5110 (N_5110,N_4870,N_4805);
and U5111 (N_5111,N_4987,N_4931);
nor U5112 (N_5112,N_4779,N_4822);
nor U5113 (N_5113,N_4985,N_4800);
and U5114 (N_5114,N_4973,N_4967);
xor U5115 (N_5115,N_4991,N_4796);
nand U5116 (N_5116,N_4802,N_4975);
nor U5117 (N_5117,N_4917,N_4803);
and U5118 (N_5118,N_4848,N_4920);
nand U5119 (N_5119,N_4994,N_4781);
or U5120 (N_5120,N_4912,N_4935);
and U5121 (N_5121,N_4769,N_4756);
nor U5122 (N_5122,N_4885,N_4906);
nand U5123 (N_5123,N_4820,N_4926);
nand U5124 (N_5124,N_4766,N_4981);
nor U5125 (N_5125,N_4759,N_4839);
nand U5126 (N_5126,N_4993,N_4806);
or U5127 (N_5127,N_4774,N_4871);
xor U5128 (N_5128,N_4804,N_4942);
nand U5129 (N_5129,N_4790,N_4755);
and U5130 (N_5130,N_4977,N_4841);
or U5131 (N_5131,N_4857,N_4967);
nand U5132 (N_5132,N_4884,N_4857);
nand U5133 (N_5133,N_4838,N_4815);
nor U5134 (N_5134,N_4830,N_4933);
nor U5135 (N_5135,N_4833,N_4791);
xnor U5136 (N_5136,N_4787,N_4842);
xor U5137 (N_5137,N_4880,N_4888);
nor U5138 (N_5138,N_4815,N_4796);
nand U5139 (N_5139,N_4756,N_4941);
and U5140 (N_5140,N_4830,N_4798);
nand U5141 (N_5141,N_4973,N_4974);
nor U5142 (N_5142,N_4774,N_4984);
nand U5143 (N_5143,N_4881,N_4992);
nor U5144 (N_5144,N_4781,N_4799);
and U5145 (N_5145,N_4780,N_4757);
or U5146 (N_5146,N_4782,N_4983);
nor U5147 (N_5147,N_4819,N_4993);
nand U5148 (N_5148,N_4977,N_4894);
or U5149 (N_5149,N_4807,N_4915);
and U5150 (N_5150,N_4841,N_4789);
nor U5151 (N_5151,N_4909,N_4949);
nor U5152 (N_5152,N_4986,N_4894);
and U5153 (N_5153,N_4902,N_4850);
xnor U5154 (N_5154,N_4773,N_4947);
or U5155 (N_5155,N_4982,N_4980);
and U5156 (N_5156,N_4883,N_4996);
nand U5157 (N_5157,N_4878,N_4823);
nand U5158 (N_5158,N_4753,N_4932);
or U5159 (N_5159,N_4790,N_4771);
xor U5160 (N_5160,N_4875,N_4906);
xor U5161 (N_5161,N_4962,N_4912);
or U5162 (N_5162,N_4815,N_4800);
and U5163 (N_5163,N_4922,N_4771);
nand U5164 (N_5164,N_4957,N_4816);
and U5165 (N_5165,N_4855,N_4913);
nand U5166 (N_5166,N_4842,N_4991);
nor U5167 (N_5167,N_4810,N_4921);
and U5168 (N_5168,N_4762,N_4905);
nand U5169 (N_5169,N_4770,N_4769);
nand U5170 (N_5170,N_4961,N_4866);
or U5171 (N_5171,N_4891,N_4964);
nand U5172 (N_5172,N_4843,N_4800);
or U5173 (N_5173,N_4922,N_4778);
xor U5174 (N_5174,N_4915,N_4987);
or U5175 (N_5175,N_4963,N_4882);
nand U5176 (N_5176,N_4993,N_4915);
and U5177 (N_5177,N_4900,N_4799);
nand U5178 (N_5178,N_4862,N_4851);
or U5179 (N_5179,N_4754,N_4769);
and U5180 (N_5180,N_4794,N_4889);
or U5181 (N_5181,N_4955,N_4786);
nand U5182 (N_5182,N_4754,N_4942);
nor U5183 (N_5183,N_4813,N_4778);
nor U5184 (N_5184,N_4918,N_4760);
nor U5185 (N_5185,N_4996,N_4924);
or U5186 (N_5186,N_4898,N_4915);
nand U5187 (N_5187,N_4837,N_4751);
and U5188 (N_5188,N_4919,N_4790);
nor U5189 (N_5189,N_4794,N_4853);
and U5190 (N_5190,N_4918,N_4823);
or U5191 (N_5191,N_4854,N_4760);
or U5192 (N_5192,N_4793,N_4861);
nor U5193 (N_5193,N_4774,N_4801);
xnor U5194 (N_5194,N_4768,N_4964);
xnor U5195 (N_5195,N_4815,N_4914);
or U5196 (N_5196,N_4788,N_4913);
or U5197 (N_5197,N_4849,N_4958);
or U5198 (N_5198,N_4806,N_4898);
xnor U5199 (N_5199,N_4760,N_4992);
xor U5200 (N_5200,N_4852,N_4942);
and U5201 (N_5201,N_4853,N_4960);
nand U5202 (N_5202,N_4836,N_4926);
and U5203 (N_5203,N_4792,N_4965);
nor U5204 (N_5204,N_4915,N_4925);
nor U5205 (N_5205,N_4794,N_4954);
or U5206 (N_5206,N_4942,N_4877);
nor U5207 (N_5207,N_4986,N_4878);
and U5208 (N_5208,N_4766,N_4777);
and U5209 (N_5209,N_4890,N_4895);
and U5210 (N_5210,N_4827,N_4951);
and U5211 (N_5211,N_4952,N_4782);
and U5212 (N_5212,N_4868,N_4766);
nor U5213 (N_5213,N_4976,N_4814);
and U5214 (N_5214,N_4831,N_4963);
nand U5215 (N_5215,N_4800,N_4916);
and U5216 (N_5216,N_4948,N_4955);
or U5217 (N_5217,N_4817,N_4969);
nand U5218 (N_5218,N_4907,N_4957);
and U5219 (N_5219,N_4905,N_4967);
and U5220 (N_5220,N_4790,N_4897);
nand U5221 (N_5221,N_4760,N_4768);
nor U5222 (N_5222,N_4777,N_4767);
nand U5223 (N_5223,N_4907,N_4906);
and U5224 (N_5224,N_4792,N_4812);
or U5225 (N_5225,N_4807,N_4833);
nand U5226 (N_5226,N_4844,N_4948);
nand U5227 (N_5227,N_4992,N_4931);
and U5228 (N_5228,N_4998,N_4960);
or U5229 (N_5229,N_4756,N_4789);
nand U5230 (N_5230,N_4989,N_4956);
and U5231 (N_5231,N_4889,N_4972);
xor U5232 (N_5232,N_4771,N_4841);
or U5233 (N_5233,N_4805,N_4950);
nor U5234 (N_5234,N_4830,N_4760);
and U5235 (N_5235,N_4902,N_4896);
and U5236 (N_5236,N_4998,N_4924);
nand U5237 (N_5237,N_4820,N_4919);
nor U5238 (N_5238,N_4855,N_4850);
and U5239 (N_5239,N_4930,N_4938);
nand U5240 (N_5240,N_4846,N_4937);
nor U5241 (N_5241,N_4853,N_4940);
or U5242 (N_5242,N_4863,N_4792);
nand U5243 (N_5243,N_4946,N_4963);
nand U5244 (N_5244,N_4837,N_4927);
nand U5245 (N_5245,N_4821,N_4925);
xor U5246 (N_5246,N_4810,N_4933);
nor U5247 (N_5247,N_4841,N_4832);
or U5248 (N_5248,N_4775,N_4969);
or U5249 (N_5249,N_4989,N_4857);
and U5250 (N_5250,N_5151,N_5237);
nor U5251 (N_5251,N_5062,N_5161);
or U5252 (N_5252,N_5186,N_5032);
and U5253 (N_5253,N_5189,N_5039);
nand U5254 (N_5254,N_5029,N_5022);
nor U5255 (N_5255,N_5056,N_5191);
nor U5256 (N_5256,N_5068,N_5152);
xnor U5257 (N_5257,N_5118,N_5156);
and U5258 (N_5258,N_5199,N_5141);
nand U5259 (N_5259,N_5247,N_5236);
xor U5260 (N_5260,N_5130,N_5091);
nand U5261 (N_5261,N_5105,N_5088);
or U5262 (N_5262,N_5217,N_5017);
and U5263 (N_5263,N_5226,N_5147);
or U5264 (N_5264,N_5241,N_5221);
or U5265 (N_5265,N_5165,N_5008);
nand U5266 (N_5266,N_5051,N_5041);
or U5267 (N_5267,N_5204,N_5229);
nor U5268 (N_5268,N_5044,N_5111);
nand U5269 (N_5269,N_5164,N_5033);
nand U5270 (N_5270,N_5005,N_5149);
and U5271 (N_5271,N_5097,N_5206);
and U5272 (N_5272,N_5213,N_5163);
and U5273 (N_5273,N_5090,N_5081);
nand U5274 (N_5274,N_5173,N_5170);
xnor U5275 (N_5275,N_5037,N_5135);
nor U5276 (N_5276,N_5181,N_5215);
and U5277 (N_5277,N_5086,N_5107);
and U5278 (N_5278,N_5218,N_5210);
or U5279 (N_5279,N_5203,N_5225);
and U5280 (N_5280,N_5087,N_5198);
nand U5281 (N_5281,N_5004,N_5042);
nor U5282 (N_5282,N_5119,N_5166);
nand U5283 (N_5283,N_5243,N_5072);
and U5284 (N_5284,N_5220,N_5169);
or U5285 (N_5285,N_5002,N_5125);
nand U5286 (N_5286,N_5023,N_5099);
and U5287 (N_5287,N_5054,N_5155);
nor U5288 (N_5288,N_5193,N_5244);
or U5289 (N_5289,N_5240,N_5036);
nor U5290 (N_5290,N_5232,N_5234);
and U5291 (N_5291,N_5142,N_5224);
and U5292 (N_5292,N_5123,N_5074);
xor U5293 (N_5293,N_5235,N_5230);
and U5294 (N_5294,N_5050,N_5188);
nor U5295 (N_5295,N_5172,N_5223);
nand U5296 (N_5296,N_5026,N_5195);
nand U5297 (N_5297,N_5208,N_5146);
xor U5298 (N_5298,N_5115,N_5200);
xnor U5299 (N_5299,N_5011,N_5015);
or U5300 (N_5300,N_5192,N_5053);
and U5301 (N_5301,N_5132,N_5187);
nor U5302 (N_5302,N_5079,N_5185);
xnor U5303 (N_5303,N_5176,N_5231);
and U5304 (N_5304,N_5083,N_5177);
nand U5305 (N_5305,N_5073,N_5212);
nand U5306 (N_5306,N_5158,N_5038);
and U5307 (N_5307,N_5043,N_5064);
nand U5308 (N_5308,N_5127,N_5171);
and U5309 (N_5309,N_5096,N_5067);
nand U5310 (N_5310,N_5092,N_5209);
or U5311 (N_5311,N_5065,N_5108);
nand U5312 (N_5312,N_5194,N_5012);
nor U5313 (N_5313,N_5030,N_5028);
nand U5314 (N_5314,N_5024,N_5070);
xor U5315 (N_5315,N_5134,N_5157);
or U5316 (N_5316,N_5202,N_5001);
nor U5317 (N_5317,N_5093,N_5106);
or U5318 (N_5318,N_5128,N_5129);
nor U5319 (N_5319,N_5003,N_5143);
nor U5320 (N_5320,N_5000,N_5239);
or U5321 (N_5321,N_5047,N_5197);
and U5322 (N_5322,N_5245,N_5178);
nand U5323 (N_5323,N_5190,N_5084);
nor U5324 (N_5324,N_5183,N_5075);
nor U5325 (N_5325,N_5205,N_5122);
nor U5326 (N_5326,N_5154,N_5094);
or U5327 (N_5327,N_5078,N_5100);
or U5328 (N_5328,N_5114,N_5150);
or U5329 (N_5329,N_5139,N_5219);
or U5330 (N_5330,N_5137,N_5216);
nor U5331 (N_5331,N_5184,N_5248);
or U5332 (N_5332,N_5104,N_5233);
nor U5333 (N_5333,N_5201,N_5082);
nand U5334 (N_5334,N_5034,N_5174);
xor U5335 (N_5335,N_5168,N_5080);
or U5336 (N_5336,N_5116,N_5016);
and U5337 (N_5337,N_5018,N_5089);
nand U5338 (N_5338,N_5101,N_5025);
nand U5339 (N_5339,N_5035,N_5162);
nand U5340 (N_5340,N_5175,N_5066);
xor U5341 (N_5341,N_5031,N_5058);
and U5342 (N_5342,N_5242,N_5246);
and U5343 (N_5343,N_5238,N_5059);
xnor U5344 (N_5344,N_5121,N_5144);
nor U5345 (N_5345,N_5019,N_5049);
nand U5346 (N_5346,N_5048,N_5120);
nand U5347 (N_5347,N_5140,N_5027);
or U5348 (N_5348,N_5124,N_5110);
nor U5349 (N_5349,N_5211,N_5249);
or U5350 (N_5350,N_5045,N_5222);
nor U5351 (N_5351,N_5117,N_5040);
or U5352 (N_5352,N_5102,N_5160);
or U5353 (N_5353,N_5006,N_5007);
nand U5354 (N_5354,N_5076,N_5061);
xor U5355 (N_5355,N_5167,N_5126);
or U5356 (N_5356,N_5046,N_5052);
or U5357 (N_5357,N_5098,N_5060);
and U5358 (N_5358,N_5133,N_5013);
nand U5359 (N_5359,N_5227,N_5112);
nor U5360 (N_5360,N_5077,N_5057);
nand U5361 (N_5361,N_5085,N_5138);
nor U5362 (N_5362,N_5095,N_5207);
or U5363 (N_5363,N_5009,N_5063);
and U5364 (N_5364,N_5214,N_5180);
nand U5365 (N_5365,N_5020,N_5148);
or U5366 (N_5366,N_5014,N_5109);
and U5367 (N_5367,N_5228,N_5153);
nor U5368 (N_5368,N_5131,N_5136);
or U5369 (N_5369,N_5055,N_5159);
or U5370 (N_5370,N_5145,N_5196);
xor U5371 (N_5371,N_5069,N_5113);
and U5372 (N_5372,N_5021,N_5179);
nor U5373 (N_5373,N_5182,N_5071);
nand U5374 (N_5374,N_5103,N_5010);
nand U5375 (N_5375,N_5080,N_5041);
nor U5376 (N_5376,N_5211,N_5174);
nor U5377 (N_5377,N_5053,N_5148);
or U5378 (N_5378,N_5032,N_5057);
nor U5379 (N_5379,N_5245,N_5200);
and U5380 (N_5380,N_5125,N_5107);
nand U5381 (N_5381,N_5161,N_5159);
and U5382 (N_5382,N_5067,N_5072);
and U5383 (N_5383,N_5128,N_5135);
nor U5384 (N_5384,N_5212,N_5024);
nor U5385 (N_5385,N_5247,N_5058);
or U5386 (N_5386,N_5208,N_5055);
nand U5387 (N_5387,N_5234,N_5039);
nand U5388 (N_5388,N_5055,N_5181);
nand U5389 (N_5389,N_5020,N_5167);
nand U5390 (N_5390,N_5223,N_5120);
nor U5391 (N_5391,N_5158,N_5196);
and U5392 (N_5392,N_5179,N_5090);
xnor U5393 (N_5393,N_5057,N_5112);
nor U5394 (N_5394,N_5247,N_5099);
and U5395 (N_5395,N_5043,N_5179);
nor U5396 (N_5396,N_5020,N_5108);
nor U5397 (N_5397,N_5137,N_5174);
and U5398 (N_5398,N_5187,N_5084);
nand U5399 (N_5399,N_5090,N_5000);
and U5400 (N_5400,N_5141,N_5213);
nand U5401 (N_5401,N_5026,N_5036);
nor U5402 (N_5402,N_5089,N_5091);
nand U5403 (N_5403,N_5007,N_5029);
and U5404 (N_5404,N_5082,N_5181);
and U5405 (N_5405,N_5175,N_5070);
and U5406 (N_5406,N_5003,N_5002);
or U5407 (N_5407,N_5162,N_5181);
or U5408 (N_5408,N_5137,N_5078);
xor U5409 (N_5409,N_5185,N_5138);
and U5410 (N_5410,N_5246,N_5148);
xnor U5411 (N_5411,N_5055,N_5147);
nor U5412 (N_5412,N_5238,N_5034);
nand U5413 (N_5413,N_5249,N_5241);
nor U5414 (N_5414,N_5106,N_5136);
nor U5415 (N_5415,N_5032,N_5101);
nor U5416 (N_5416,N_5208,N_5071);
or U5417 (N_5417,N_5177,N_5093);
nand U5418 (N_5418,N_5015,N_5207);
or U5419 (N_5419,N_5057,N_5200);
or U5420 (N_5420,N_5042,N_5154);
xor U5421 (N_5421,N_5095,N_5042);
nor U5422 (N_5422,N_5194,N_5212);
nor U5423 (N_5423,N_5210,N_5054);
and U5424 (N_5424,N_5224,N_5051);
and U5425 (N_5425,N_5219,N_5132);
nand U5426 (N_5426,N_5241,N_5218);
nor U5427 (N_5427,N_5112,N_5166);
and U5428 (N_5428,N_5110,N_5134);
nor U5429 (N_5429,N_5181,N_5099);
or U5430 (N_5430,N_5106,N_5014);
nand U5431 (N_5431,N_5162,N_5114);
or U5432 (N_5432,N_5234,N_5062);
and U5433 (N_5433,N_5115,N_5094);
nand U5434 (N_5434,N_5110,N_5009);
nor U5435 (N_5435,N_5238,N_5036);
nor U5436 (N_5436,N_5129,N_5212);
xnor U5437 (N_5437,N_5213,N_5190);
and U5438 (N_5438,N_5060,N_5072);
nor U5439 (N_5439,N_5152,N_5058);
or U5440 (N_5440,N_5145,N_5173);
nand U5441 (N_5441,N_5002,N_5018);
nor U5442 (N_5442,N_5017,N_5236);
nand U5443 (N_5443,N_5123,N_5041);
nor U5444 (N_5444,N_5047,N_5120);
nor U5445 (N_5445,N_5152,N_5208);
xor U5446 (N_5446,N_5085,N_5245);
xor U5447 (N_5447,N_5023,N_5019);
nor U5448 (N_5448,N_5142,N_5229);
or U5449 (N_5449,N_5045,N_5249);
nor U5450 (N_5450,N_5044,N_5113);
nand U5451 (N_5451,N_5085,N_5009);
xor U5452 (N_5452,N_5108,N_5218);
or U5453 (N_5453,N_5137,N_5130);
and U5454 (N_5454,N_5219,N_5231);
nor U5455 (N_5455,N_5138,N_5165);
xnor U5456 (N_5456,N_5188,N_5231);
xnor U5457 (N_5457,N_5001,N_5221);
nor U5458 (N_5458,N_5209,N_5203);
nand U5459 (N_5459,N_5092,N_5075);
or U5460 (N_5460,N_5186,N_5063);
nand U5461 (N_5461,N_5099,N_5210);
nor U5462 (N_5462,N_5212,N_5135);
and U5463 (N_5463,N_5008,N_5227);
nand U5464 (N_5464,N_5097,N_5015);
xor U5465 (N_5465,N_5103,N_5179);
or U5466 (N_5466,N_5112,N_5245);
nor U5467 (N_5467,N_5076,N_5223);
or U5468 (N_5468,N_5012,N_5199);
nor U5469 (N_5469,N_5149,N_5015);
and U5470 (N_5470,N_5029,N_5091);
or U5471 (N_5471,N_5093,N_5111);
and U5472 (N_5472,N_5217,N_5052);
and U5473 (N_5473,N_5163,N_5053);
nor U5474 (N_5474,N_5175,N_5009);
or U5475 (N_5475,N_5105,N_5185);
nand U5476 (N_5476,N_5119,N_5225);
and U5477 (N_5477,N_5042,N_5204);
and U5478 (N_5478,N_5116,N_5047);
and U5479 (N_5479,N_5131,N_5043);
and U5480 (N_5480,N_5133,N_5088);
nand U5481 (N_5481,N_5037,N_5011);
and U5482 (N_5482,N_5041,N_5164);
and U5483 (N_5483,N_5082,N_5038);
and U5484 (N_5484,N_5243,N_5042);
and U5485 (N_5485,N_5163,N_5049);
nand U5486 (N_5486,N_5231,N_5002);
and U5487 (N_5487,N_5098,N_5053);
and U5488 (N_5488,N_5145,N_5143);
nor U5489 (N_5489,N_5075,N_5027);
and U5490 (N_5490,N_5143,N_5047);
nor U5491 (N_5491,N_5010,N_5210);
and U5492 (N_5492,N_5136,N_5166);
xor U5493 (N_5493,N_5061,N_5099);
xor U5494 (N_5494,N_5188,N_5198);
or U5495 (N_5495,N_5048,N_5093);
nor U5496 (N_5496,N_5038,N_5060);
nor U5497 (N_5497,N_5159,N_5074);
nand U5498 (N_5498,N_5100,N_5106);
and U5499 (N_5499,N_5212,N_5001);
nor U5500 (N_5500,N_5286,N_5411);
nand U5501 (N_5501,N_5291,N_5339);
nand U5502 (N_5502,N_5433,N_5284);
and U5503 (N_5503,N_5299,N_5491);
nor U5504 (N_5504,N_5274,N_5407);
nand U5505 (N_5505,N_5409,N_5383);
nand U5506 (N_5506,N_5413,N_5363);
xnor U5507 (N_5507,N_5495,N_5289);
or U5508 (N_5508,N_5482,N_5329);
or U5509 (N_5509,N_5387,N_5323);
nand U5510 (N_5510,N_5271,N_5451);
nor U5511 (N_5511,N_5468,N_5312);
or U5512 (N_5512,N_5301,N_5268);
nand U5513 (N_5513,N_5483,N_5358);
nand U5514 (N_5514,N_5444,N_5362);
and U5515 (N_5515,N_5379,N_5479);
or U5516 (N_5516,N_5399,N_5382);
nand U5517 (N_5517,N_5280,N_5288);
nor U5518 (N_5518,N_5488,N_5348);
and U5519 (N_5519,N_5275,N_5425);
nor U5520 (N_5520,N_5309,N_5297);
nor U5521 (N_5521,N_5269,N_5380);
xor U5522 (N_5522,N_5422,N_5262);
xor U5523 (N_5523,N_5276,N_5345);
xor U5524 (N_5524,N_5469,N_5313);
nor U5525 (N_5525,N_5321,N_5304);
nor U5526 (N_5526,N_5449,N_5394);
or U5527 (N_5527,N_5277,N_5418);
and U5528 (N_5528,N_5455,N_5253);
or U5529 (N_5529,N_5320,N_5443);
and U5530 (N_5530,N_5252,N_5498);
nand U5531 (N_5531,N_5270,N_5251);
nand U5532 (N_5532,N_5279,N_5282);
xor U5533 (N_5533,N_5424,N_5298);
and U5534 (N_5534,N_5361,N_5373);
or U5535 (N_5535,N_5486,N_5341);
nor U5536 (N_5536,N_5344,N_5333);
xor U5537 (N_5537,N_5300,N_5406);
and U5538 (N_5538,N_5336,N_5342);
nor U5539 (N_5539,N_5368,N_5448);
nand U5540 (N_5540,N_5366,N_5352);
nand U5541 (N_5541,N_5293,N_5319);
nand U5542 (N_5542,N_5435,N_5462);
nor U5543 (N_5543,N_5476,N_5439);
nor U5544 (N_5544,N_5317,N_5471);
or U5545 (N_5545,N_5428,N_5485);
or U5546 (N_5546,N_5472,N_5408);
xnor U5547 (N_5547,N_5350,N_5351);
or U5548 (N_5548,N_5402,N_5267);
and U5549 (N_5549,N_5461,N_5403);
xnor U5550 (N_5550,N_5359,N_5384);
or U5551 (N_5551,N_5258,N_5427);
and U5552 (N_5552,N_5255,N_5392);
nor U5553 (N_5553,N_5493,N_5453);
and U5554 (N_5554,N_5434,N_5378);
nor U5555 (N_5555,N_5315,N_5330);
or U5556 (N_5556,N_5480,N_5396);
or U5557 (N_5557,N_5490,N_5260);
and U5558 (N_5558,N_5395,N_5305);
or U5559 (N_5559,N_5326,N_5347);
and U5560 (N_5560,N_5302,N_5343);
nor U5561 (N_5561,N_5474,N_5393);
and U5562 (N_5562,N_5404,N_5442);
and U5563 (N_5563,N_5325,N_5283);
nor U5564 (N_5564,N_5446,N_5464);
nand U5565 (N_5565,N_5445,N_5257);
nor U5566 (N_5566,N_5412,N_5308);
nand U5567 (N_5567,N_5332,N_5459);
nand U5568 (N_5568,N_5294,N_5487);
and U5569 (N_5569,N_5385,N_5458);
nor U5570 (N_5570,N_5381,N_5431);
nand U5571 (N_5571,N_5386,N_5401);
xor U5572 (N_5572,N_5365,N_5263);
nand U5573 (N_5573,N_5254,N_5338);
nand U5574 (N_5574,N_5314,N_5290);
nand U5575 (N_5575,N_5481,N_5375);
or U5576 (N_5576,N_5272,N_5460);
or U5577 (N_5577,N_5410,N_5318);
nor U5578 (N_5578,N_5429,N_5419);
and U5579 (N_5579,N_5369,N_5389);
or U5580 (N_5580,N_5287,N_5273);
nor U5581 (N_5581,N_5440,N_5374);
nor U5582 (N_5582,N_5261,N_5296);
and U5583 (N_5583,N_5370,N_5414);
and U5584 (N_5584,N_5398,N_5447);
or U5585 (N_5585,N_5295,N_5281);
nor U5586 (N_5586,N_5466,N_5372);
nand U5587 (N_5587,N_5457,N_5349);
or U5588 (N_5588,N_5292,N_5285);
nor U5589 (N_5589,N_5250,N_5420);
nor U5590 (N_5590,N_5452,N_5477);
xnor U5591 (N_5591,N_5327,N_5494);
nand U5592 (N_5592,N_5377,N_5278);
nand U5593 (N_5593,N_5416,N_5467);
or U5594 (N_5594,N_5353,N_5334);
nor U5595 (N_5595,N_5324,N_5367);
nor U5596 (N_5596,N_5311,N_5423);
and U5597 (N_5597,N_5355,N_5478);
or U5598 (N_5598,N_5454,N_5316);
nor U5599 (N_5599,N_5357,N_5475);
nand U5600 (N_5600,N_5328,N_5388);
or U5601 (N_5601,N_5415,N_5256);
and U5602 (N_5602,N_5356,N_5266);
and U5603 (N_5603,N_5354,N_5376);
and U5604 (N_5604,N_5489,N_5322);
and U5605 (N_5605,N_5400,N_5346);
nor U5606 (N_5606,N_5436,N_5397);
and U5607 (N_5607,N_5360,N_5496);
or U5608 (N_5608,N_5310,N_5426);
nor U5609 (N_5609,N_5259,N_5438);
nand U5610 (N_5610,N_5391,N_5337);
or U5611 (N_5611,N_5390,N_5437);
or U5612 (N_5612,N_5497,N_5441);
and U5613 (N_5613,N_5465,N_5432);
nand U5614 (N_5614,N_5417,N_5303);
nor U5615 (N_5615,N_5499,N_5450);
or U5616 (N_5616,N_5340,N_5307);
or U5617 (N_5617,N_5470,N_5492);
nor U5618 (N_5618,N_5405,N_5364);
and U5619 (N_5619,N_5463,N_5306);
xor U5620 (N_5620,N_5331,N_5456);
nand U5621 (N_5621,N_5264,N_5265);
or U5622 (N_5622,N_5484,N_5421);
nand U5623 (N_5623,N_5371,N_5335);
and U5624 (N_5624,N_5473,N_5430);
nor U5625 (N_5625,N_5325,N_5444);
nor U5626 (N_5626,N_5455,N_5298);
or U5627 (N_5627,N_5390,N_5482);
and U5628 (N_5628,N_5360,N_5315);
or U5629 (N_5629,N_5345,N_5403);
nor U5630 (N_5630,N_5258,N_5483);
nand U5631 (N_5631,N_5361,N_5379);
nand U5632 (N_5632,N_5305,N_5465);
nor U5633 (N_5633,N_5413,N_5335);
and U5634 (N_5634,N_5368,N_5387);
and U5635 (N_5635,N_5438,N_5387);
or U5636 (N_5636,N_5392,N_5468);
nor U5637 (N_5637,N_5280,N_5369);
nand U5638 (N_5638,N_5274,N_5372);
or U5639 (N_5639,N_5419,N_5396);
and U5640 (N_5640,N_5491,N_5350);
nor U5641 (N_5641,N_5460,N_5370);
and U5642 (N_5642,N_5467,N_5254);
nor U5643 (N_5643,N_5252,N_5358);
nand U5644 (N_5644,N_5457,N_5465);
or U5645 (N_5645,N_5324,N_5348);
nand U5646 (N_5646,N_5422,N_5322);
nand U5647 (N_5647,N_5481,N_5335);
or U5648 (N_5648,N_5478,N_5298);
nand U5649 (N_5649,N_5256,N_5323);
or U5650 (N_5650,N_5302,N_5476);
and U5651 (N_5651,N_5339,N_5477);
or U5652 (N_5652,N_5292,N_5340);
or U5653 (N_5653,N_5438,N_5314);
nand U5654 (N_5654,N_5484,N_5379);
nor U5655 (N_5655,N_5306,N_5279);
nand U5656 (N_5656,N_5366,N_5444);
xor U5657 (N_5657,N_5430,N_5437);
nand U5658 (N_5658,N_5362,N_5385);
and U5659 (N_5659,N_5440,N_5456);
nand U5660 (N_5660,N_5373,N_5473);
and U5661 (N_5661,N_5338,N_5333);
and U5662 (N_5662,N_5493,N_5315);
nand U5663 (N_5663,N_5450,N_5482);
and U5664 (N_5664,N_5326,N_5404);
and U5665 (N_5665,N_5436,N_5360);
and U5666 (N_5666,N_5370,N_5305);
and U5667 (N_5667,N_5355,N_5264);
nor U5668 (N_5668,N_5335,N_5432);
and U5669 (N_5669,N_5460,N_5320);
or U5670 (N_5670,N_5257,N_5408);
nand U5671 (N_5671,N_5486,N_5315);
and U5672 (N_5672,N_5301,N_5257);
or U5673 (N_5673,N_5368,N_5296);
nand U5674 (N_5674,N_5424,N_5409);
or U5675 (N_5675,N_5365,N_5358);
nand U5676 (N_5676,N_5326,N_5292);
xor U5677 (N_5677,N_5383,N_5284);
and U5678 (N_5678,N_5448,N_5311);
and U5679 (N_5679,N_5370,N_5375);
or U5680 (N_5680,N_5251,N_5322);
or U5681 (N_5681,N_5298,N_5456);
nor U5682 (N_5682,N_5377,N_5281);
nand U5683 (N_5683,N_5465,N_5255);
or U5684 (N_5684,N_5468,N_5495);
or U5685 (N_5685,N_5447,N_5377);
and U5686 (N_5686,N_5377,N_5356);
nand U5687 (N_5687,N_5385,N_5412);
nand U5688 (N_5688,N_5382,N_5444);
and U5689 (N_5689,N_5378,N_5424);
and U5690 (N_5690,N_5418,N_5473);
nand U5691 (N_5691,N_5289,N_5323);
nand U5692 (N_5692,N_5434,N_5383);
nor U5693 (N_5693,N_5283,N_5342);
nor U5694 (N_5694,N_5391,N_5268);
or U5695 (N_5695,N_5268,N_5396);
nand U5696 (N_5696,N_5413,N_5250);
nor U5697 (N_5697,N_5308,N_5402);
nand U5698 (N_5698,N_5497,N_5262);
nor U5699 (N_5699,N_5307,N_5403);
and U5700 (N_5700,N_5313,N_5272);
and U5701 (N_5701,N_5368,N_5438);
nand U5702 (N_5702,N_5463,N_5257);
or U5703 (N_5703,N_5493,N_5434);
xor U5704 (N_5704,N_5284,N_5411);
nor U5705 (N_5705,N_5339,N_5306);
xor U5706 (N_5706,N_5342,N_5330);
and U5707 (N_5707,N_5255,N_5268);
and U5708 (N_5708,N_5257,N_5405);
or U5709 (N_5709,N_5395,N_5260);
nor U5710 (N_5710,N_5458,N_5441);
or U5711 (N_5711,N_5482,N_5468);
nor U5712 (N_5712,N_5301,N_5391);
xor U5713 (N_5713,N_5311,N_5373);
nor U5714 (N_5714,N_5282,N_5342);
nand U5715 (N_5715,N_5262,N_5414);
and U5716 (N_5716,N_5266,N_5289);
or U5717 (N_5717,N_5254,N_5288);
xor U5718 (N_5718,N_5327,N_5318);
nor U5719 (N_5719,N_5354,N_5390);
nor U5720 (N_5720,N_5449,N_5359);
nor U5721 (N_5721,N_5417,N_5270);
and U5722 (N_5722,N_5461,N_5451);
nor U5723 (N_5723,N_5306,N_5423);
or U5724 (N_5724,N_5291,N_5255);
nor U5725 (N_5725,N_5302,N_5378);
and U5726 (N_5726,N_5291,N_5344);
nor U5727 (N_5727,N_5437,N_5323);
xnor U5728 (N_5728,N_5368,N_5373);
or U5729 (N_5729,N_5487,N_5479);
nand U5730 (N_5730,N_5395,N_5348);
and U5731 (N_5731,N_5313,N_5494);
and U5732 (N_5732,N_5468,N_5333);
nand U5733 (N_5733,N_5327,N_5362);
and U5734 (N_5734,N_5465,N_5397);
nor U5735 (N_5735,N_5347,N_5337);
nand U5736 (N_5736,N_5310,N_5293);
nand U5737 (N_5737,N_5465,N_5293);
nand U5738 (N_5738,N_5491,N_5304);
nor U5739 (N_5739,N_5472,N_5450);
and U5740 (N_5740,N_5438,N_5455);
or U5741 (N_5741,N_5300,N_5455);
and U5742 (N_5742,N_5311,N_5261);
nor U5743 (N_5743,N_5337,N_5461);
or U5744 (N_5744,N_5459,N_5393);
and U5745 (N_5745,N_5459,N_5391);
xor U5746 (N_5746,N_5493,N_5422);
nor U5747 (N_5747,N_5300,N_5257);
nand U5748 (N_5748,N_5297,N_5264);
or U5749 (N_5749,N_5302,N_5276);
or U5750 (N_5750,N_5563,N_5736);
xnor U5751 (N_5751,N_5562,N_5611);
and U5752 (N_5752,N_5645,N_5732);
and U5753 (N_5753,N_5612,N_5729);
nor U5754 (N_5754,N_5692,N_5578);
nor U5755 (N_5755,N_5727,N_5748);
nor U5756 (N_5756,N_5657,N_5740);
nand U5757 (N_5757,N_5716,N_5577);
xnor U5758 (N_5758,N_5631,N_5518);
nand U5759 (N_5759,N_5633,N_5704);
or U5760 (N_5760,N_5569,N_5618);
nand U5761 (N_5761,N_5521,N_5658);
nor U5762 (N_5762,N_5583,N_5630);
and U5763 (N_5763,N_5509,N_5543);
or U5764 (N_5764,N_5636,N_5683);
nor U5765 (N_5765,N_5580,N_5667);
or U5766 (N_5766,N_5643,N_5553);
and U5767 (N_5767,N_5574,N_5546);
nand U5768 (N_5768,N_5539,N_5620);
or U5769 (N_5769,N_5561,N_5534);
and U5770 (N_5770,N_5549,N_5605);
and U5771 (N_5771,N_5724,N_5695);
nand U5772 (N_5772,N_5529,N_5743);
nand U5773 (N_5773,N_5511,N_5533);
or U5774 (N_5774,N_5671,N_5586);
or U5775 (N_5775,N_5500,N_5689);
or U5776 (N_5776,N_5600,N_5668);
and U5777 (N_5777,N_5610,N_5514);
xor U5778 (N_5778,N_5531,N_5523);
and U5779 (N_5779,N_5641,N_5593);
and U5780 (N_5780,N_5623,N_5552);
nor U5781 (N_5781,N_5520,N_5647);
nor U5782 (N_5782,N_5747,N_5682);
xor U5783 (N_5783,N_5651,N_5628);
and U5784 (N_5784,N_5648,N_5614);
and U5785 (N_5785,N_5607,N_5745);
nor U5786 (N_5786,N_5718,N_5678);
nor U5787 (N_5787,N_5652,N_5591);
nor U5788 (N_5788,N_5693,N_5536);
and U5789 (N_5789,N_5597,N_5505);
and U5790 (N_5790,N_5715,N_5649);
xor U5791 (N_5791,N_5710,N_5741);
nand U5792 (N_5792,N_5542,N_5502);
nor U5793 (N_5793,N_5720,N_5655);
xnor U5794 (N_5794,N_5585,N_5588);
or U5795 (N_5795,N_5621,N_5515);
nand U5796 (N_5796,N_5669,N_5616);
or U5797 (N_5797,N_5653,N_5592);
nand U5798 (N_5798,N_5598,N_5584);
nand U5799 (N_5799,N_5556,N_5567);
and U5800 (N_5800,N_5506,N_5661);
or U5801 (N_5801,N_5595,N_5730);
nor U5802 (N_5802,N_5731,N_5708);
nand U5803 (N_5803,N_5733,N_5650);
xor U5804 (N_5804,N_5530,N_5609);
xor U5805 (N_5805,N_5702,N_5656);
or U5806 (N_5806,N_5679,N_5613);
and U5807 (N_5807,N_5575,N_5725);
or U5808 (N_5808,N_5703,N_5709);
nand U5809 (N_5809,N_5507,N_5604);
or U5810 (N_5810,N_5566,N_5576);
or U5811 (N_5811,N_5599,N_5596);
and U5812 (N_5812,N_5670,N_5626);
nor U5813 (N_5813,N_5617,N_5508);
xnor U5814 (N_5814,N_5560,N_5603);
xor U5815 (N_5815,N_5699,N_5590);
and U5816 (N_5816,N_5545,N_5581);
nor U5817 (N_5817,N_5517,N_5522);
nor U5818 (N_5818,N_5512,N_5606);
nor U5819 (N_5819,N_5712,N_5686);
or U5820 (N_5820,N_5548,N_5537);
nor U5821 (N_5821,N_5632,N_5619);
or U5822 (N_5822,N_5675,N_5642);
nand U5823 (N_5823,N_5737,N_5742);
nor U5824 (N_5824,N_5734,N_5677);
nor U5825 (N_5825,N_5582,N_5565);
nand U5826 (N_5826,N_5663,N_5544);
nand U5827 (N_5827,N_5691,N_5503);
nor U5828 (N_5828,N_5510,N_5570);
and U5829 (N_5829,N_5714,N_5594);
and U5830 (N_5830,N_5538,N_5551);
nand U5831 (N_5831,N_5541,N_5639);
xor U5832 (N_5832,N_5684,N_5719);
or U5833 (N_5833,N_5717,N_5625);
or U5834 (N_5834,N_5571,N_5662);
nand U5835 (N_5835,N_5501,N_5527);
nand U5836 (N_5836,N_5681,N_5634);
or U5837 (N_5837,N_5696,N_5558);
and U5838 (N_5838,N_5680,N_5713);
or U5839 (N_5839,N_5674,N_5555);
nor U5840 (N_5840,N_5685,N_5723);
and U5841 (N_5841,N_5572,N_5644);
and U5842 (N_5842,N_5673,N_5697);
xor U5843 (N_5843,N_5654,N_5705);
nor U5844 (N_5844,N_5640,N_5627);
xnor U5845 (N_5845,N_5706,N_5624);
nand U5846 (N_5846,N_5629,N_5528);
or U5847 (N_5847,N_5519,N_5722);
or U5848 (N_5848,N_5660,N_5749);
or U5849 (N_5849,N_5687,N_5557);
nor U5850 (N_5850,N_5676,N_5587);
and U5851 (N_5851,N_5707,N_5602);
nand U5852 (N_5852,N_5700,N_5622);
or U5853 (N_5853,N_5659,N_5526);
and U5854 (N_5854,N_5688,N_5711);
nand U5855 (N_5855,N_5638,N_5564);
or U5856 (N_5856,N_5664,N_5694);
nor U5857 (N_5857,N_5579,N_5568);
or U5858 (N_5858,N_5601,N_5735);
and U5859 (N_5859,N_5608,N_5666);
nand U5860 (N_5860,N_5525,N_5744);
nor U5861 (N_5861,N_5535,N_5646);
or U5862 (N_5862,N_5746,N_5524);
and U5863 (N_5863,N_5554,N_5589);
or U5864 (N_5864,N_5532,N_5738);
and U5865 (N_5865,N_5637,N_5739);
nand U5866 (N_5866,N_5690,N_5573);
xnor U5867 (N_5867,N_5513,N_5672);
nand U5868 (N_5868,N_5635,N_5547);
or U5869 (N_5869,N_5701,N_5726);
nor U5870 (N_5870,N_5698,N_5665);
nor U5871 (N_5871,N_5728,N_5504);
or U5872 (N_5872,N_5516,N_5559);
or U5873 (N_5873,N_5550,N_5721);
or U5874 (N_5874,N_5540,N_5615);
or U5875 (N_5875,N_5663,N_5670);
or U5876 (N_5876,N_5565,N_5711);
or U5877 (N_5877,N_5705,N_5639);
nor U5878 (N_5878,N_5582,N_5626);
nor U5879 (N_5879,N_5561,N_5538);
xor U5880 (N_5880,N_5547,N_5641);
nand U5881 (N_5881,N_5745,N_5704);
nor U5882 (N_5882,N_5684,N_5516);
xnor U5883 (N_5883,N_5642,N_5514);
xnor U5884 (N_5884,N_5694,N_5630);
nand U5885 (N_5885,N_5681,N_5528);
or U5886 (N_5886,N_5543,N_5691);
nor U5887 (N_5887,N_5737,N_5600);
nor U5888 (N_5888,N_5582,N_5648);
nor U5889 (N_5889,N_5508,N_5652);
or U5890 (N_5890,N_5709,N_5717);
xor U5891 (N_5891,N_5726,N_5513);
or U5892 (N_5892,N_5643,N_5518);
and U5893 (N_5893,N_5562,N_5525);
nor U5894 (N_5894,N_5724,N_5738);
xnor U5895 (N_5895,N_5662,N_5668);
nor U5896 (N_5896,N_5730,N_5582);
and U5897 (N_5897,N_5578,N_5520);
and U5898 (N_5898,N_5558,N_5595);
xnor U5899 (N_5899,N_5533,N_5664);
nand U5900 (N_5900,N_5743,N_5722);
and U5901 (N_5901,N_5632,N_5615);
nand U5902 (N_5902,N_5530,N_5722);
or U5903 (N_5903,N_5694,N_5628);
xnor U5904 (N_5904,N_5545,N_5583);
and U5905 (N_5905,N_5526,N_5697);
and U5906 (N_5906,N_5742,N_5745);
or U5907 (N_5907,N_5619,N_5689);
or U5908 (N_5908,N_5635,N_5650);
nor U5909 (N_5909,N_5511,N_5570);
nand U5910 (N_5910,N_5597,N_5705);
and U5911 (N_5911,N_5643,N_5634);
nand U5912 (N_5912,N_5635,N_5685);
nand U5913 (N_5913,N_5544,N_5741);
nand U5914 (N_5914,N_5589,N_5636);
nor U5915 (N_5915,N_5587,N_5687);
xnor U5916 (N_5916,N_5512,N_5580);
nand U5917 (N_5917,N_5568,N_5663);
nor U5918 (N_5918,N_5711,N_5619);
nor U5919 (N_5919,N_5635,N_5617);
and U5920 (N_5920,N_5593,N_5537);
xnor U5921 (N_5921,N_5515,N_5644);
or U5922 (N_5922,N_5719,N_5718);
or U5923 (N_5923,N_5742,N_5565);
and U5924 (N_5924,N_5546,N_5519);
xor U5925 (N_5925,N_5739,N_5709);
or U5926 (N_5926,N_5622,N_5690);
nor U5927 (N_5927,N_5687,N_5501);
and U5928 (N_5928,N_5740,N_5599);
nor U5929 (N_5929,N_5579,N_5727);
and U5930 (N_5930,N_5515,N_5617);
nor U5931 (N_5931,N_5684,N_5728);
and U5932 (N_5932,N_5701,N_5628);
nand U5933 (N_5933,N_5504,N_5645);
nor U5934 (N_5934,N_5657,N_5589);
nor U5935 (N_5935,N_5702,N_5591);
xnor U5936 (N_5936,N_5565,N_5637);
and U5937 (N_5937,N_5722,N_5699);
and U5938 (N_5938,N_5707,N_5620);
and U5939 (N_5939,N_5590,N_5584);
nand U5940 (N_5940,N_5735,N_5655);
nor U5941 (N_5941,N_5553,N_5586);
nand U5942 (N_5942,N_5742,N_5544);
or U5943 (N_5943,N_5734,N_5714);
or U5944 (N_5944,N_5541,N_5706);
nor U5945 (N_5945,N_5572,N_5530);
or U5946 (N_5946,N_5589,N_5693);
nor U5947 (N_5947,N_5729,N_5736);
and U5948 (N_5948,N_5527,N_5579);
nor U5949 (N_5949,N_5664,N_5702);
and U5950 (N_5950,N_5565,N_5691);
and U5951 (N_5951,N_5542,N_5519);
and U5952 (N_5952,N_5570,N_5514);
or U5953 (N_5953,N_5699,N_5546);
nor U5954 (N_5954,N_5693,N_5738);
and U5955 (N_5955,N_5600,N_5745);
xnor U5956 (N_5956,N_5735,N_5626);
or U5957 (N_5957,N_5689,N_5519);
nand U5958 (N_5958,N_5584,N_5706);
nand U5959 (N_5959,N_5516,N_5653);
nand U5960 (N_5960,N_5569,N_5719);
nor U5961 (N_5961,N_5532,N_5700);
nor U5962 (N_5962,N_5503,N_5711);
nand U5963 (N_5963,N_5693,N_5506);
and U5964 (N_5964,N_5524,N_5561);
and U5965 (N_5965,N_5529,N_5500);
or U5966 (N_5966,N_5634,N_5546);
nand U5967 (N_5967,N_5503,N_5593);
or U5968 (N_5968,N_5568,N_5542);
and U5969 (N_5969,N_5697,N_5737);
nor U5970 (N_5970,N_5586,N_5648);
nand U5971 (N_5971,N_5695,N_5565);
nor U5972 (N_5972,N_5591,N_5632);
nor U5973 (N_5973,N_5733,N_5712);
or U5974 (N_5974,N_5622,N_5736);
or U5975 (N_5975,N_5692,N_5667);
nand U5976 (N_5976,N_5693,N_5510);
and U5977 (N_5977,N_5716,N_5706);
and U5978 (N_5978,N_5684,N_5617);
nor U5979 (N_5979,N_5527,N_5630);
nand U5980 (N_5980,N_5555,N_5614);
and U5981 (N_5981,N_5588,N_5538);
xnor U5982 (N_5982,N_5544,N_5537);
and U5983 (N_5983,N_5645,N_5536);
nor U5984 (N_5984,N_5608,N_5697);
xor U5985 (N_5985,N_5515,N_5597);
nor U5986 (N_5986,N_5686,N_5513);
and U5987 (N_5987,N_5588,N_5656);
nand U5988 (N_5988,N_5519,N_5511);
or U5989 (N_5989,N_5694,N_5710);
nor U5990 (N_5990,N_5513,N_5541);
or U5991 (N_5991,N_5706,N_5649);
or U5992 (N_5992,N_5645,N_5510);
or U5993 (N_5993,N_5703,N_5645);
nand U5994 (N_5994,N_5535,N_5508);
nand U5995 (N_5995,N_5602,N_5694);
nand U5996 (N_5996,N_5680,N_5674);
nor U5997 (N_5997,N_5500,N_5597);
nor U5998 (N_5998,N_5536,N_5597);
nor U5999 (N_5999,N_5584,N_5521);
or U6000 (N_6000,N_5991,N_5838);
nor U6001 (N_6001,N_5810,N_5818);
or U6002 (N_6002,N_5859,N_5948);
or U6003 (N_6003,N_5915,N_5825);
nor U6004 (N_6004,N_5980,N_5949);
nand U6005 (N_6005,N_5773,N_5911);
nor U6006 (N_6006,N_5887,N_5833);
nand U6007 (N_6007,N_5937,N_5976);
or U6008 (N_6008,N_5794,N_5871);
nand U6009 (N_6009,N_5854,N_5930);
xor U6010 (N_6010,N_5858,N_5908);
nor U6011 (N_6011,N_5777,N_5924);
or U6012 (N_6012,N_5954,N_5775);
nand U6013 (N_6013,N_5923,N_5888);
and U6014 (N_6014,N_5761,N_5837);
and U6015 (N_6015,N_5857,N_5804);
nand U6016 (N_6016,N_5769,N_5856);
nor U6017 (N_6017,N_5996,N_5814);
and U6018 (N_6018,N_5989,N_5831);
and U6019 (N_6019,N_5965,N_5907);
or U6020 (N_6020,N_5817,N_5929);
and U6021 (N_6021,N_5821,N_5840);
and U6022 (N_6022,N_5780,N_5984);
nand U6023 (N_6023,N_5851,N_5999);
and U6024 (N_6024,N_5884,N_5849);
or U6025 (N_6025,N_5865,N_5863);
or U6026 (N_6026,N_5811,N_5905);
or U6027 (N_6027,N_5771,N_5787);
or U6028 (N_6028,N_5920,N_5809);
and U6029 (N_6029,N_5791,N_5862);
and U6030 (N_6030,N_5826,N_5874);
xnor U6031 (N_6031,N_5927,N_5952);
or U6032 (N_6032,N_5970,N_5968);
nor U6033 (N_6033,N_5881,N_5788);
nor U6034 (N_6034,N_5990,N_5926);
nand U6035 (N_6035,N_5898,N_5979);
nand U6036 (N_6036,N_5909,N_5992);
or U6037 (N_6037,N_5767,N_5805);
nor U6038 (N_6038,N_5830,N_5764);
and U6039 (N_6039,N_5969,N_5935);
nor U6040 (N_6040,N_5896,N_5768);
or U6041 (N_6041,N_5934,N_5974);
and U6042 (N_6042,N_5950,N_5963);
nor U6043 (N_6043,N_5770,N_5766);
and U6044 (N_6044,N_5759,N_5755);
or U6045 (N_6045,N_5835,N_5997);
nor U6046 (N_6046,N_5802,N_5828);
or U6047 (N_6047,N_5993,N_5815);
and U6048 (N_6048,N_5894,N_5943);
and U6049 (N_6049,N_5936,N_5783);
nor U6050 (N_6050,N_5793,N_5891);
nand U6051 (N_6051,N_5883,N_5803);
or U6052 (N_6052,N_5786,N_5986);
and U6053 (N_6053,N_5752,N_5841);
nand U6054 (N_6054,N_5827,N_5760);
nor U6055 (N_6055,N_5903,N_5978);
nor U6056 (N_6056,N_5901,N_5796);
nor U6057 (N_6057,N_5751,N_5875);
nand U6058 (N_6058,N_5848,N_5958);
or U6059 (N_6059,N_5754,N_5942);
or U6060 (N_6060,N_5800,N_5843);
nor U6061 (N_6061,N_5906,N_5774);
nor U6062 (N_6062,N_5872,N_5779);
or U6063 (N_6063,N_5945,N_5910);
nor U6064 (N_6064,N_5762,N_5822);
and U6065 (N_6065,N_5799,N_5756);
nor U6066 (N_6066,N_5944,N_5964);
nor U6067 (N_6067,N_5880,N_5866);
nand U6068 (N_6068,N_5765,N_5876);
nor U6069 (N_6069,N_5868,N_5961);
and U6070 (N_6070,N_5941,N_5782);
nand U6071 (N_6071,N_5852,N_5878);
nand U6072 (N_6072,N_5988,N_5890);
or U6073 (N_6073,N_5959,N_5972);
or U6074 (N_6074,N_5850,N_5922);
and U6075 (N_6075,N_5873,N_5940);
nor U6076 (N_6076,N_5860,N_5844);
xnor U6077 (N_6077,N_5933,N_5960);
nand U6078 (N_6078,N_5886,N_5892);
xnor U6079 (N_6079,N_5953,N_5987);
or U6080 (N_6080,N_5776,N_5807);
nand U6081 (N_6081,N_5785,N_5897);
xor U6082 (N_6082,N_5913,N_5946);
or U6083 (N_6083,N_5846,N_5947);
or U6084 (N_6084,N_5895,N_5784);
or U6085 (N_6085,N_5882,N_5870);
nand U6086 (N_6086,N_5967,N_5845);
nand U6087 (N_6087,N_5889,N_5763);
nand U6088 (N_6088,N_5998,N_5981);
nor U6089 (N_6089,N_5877,N_5994);
and U6090 (N_6090,N_5932,N_5829);
and U6091 (N_6091,N_5962,N_5772);
xnor U6092 (N_6092,N_5983,N_5753);
nand U6093 (N_6093,N_5973,N_5995);
nor U6094 (N_6094,N_5834,N_5869);
or U6095 (N_6095,N_5975,N_5956);
nor U6096 (N_6096,N_5931,N_5966);
nand U6097 (N_6097,N_5798,N_5939);
nor U6098 (N_6098,N_5912,N_5916);
or U6099 (N_6099,N_5904,N_5938);
nor U6100 (N_6100,N_5847,N_5982);
and U6101 (N_6101,N_5977,N_5855);
nand U6102 (N_6102,N_5806,N_5816);
and U6103 (N_6103,N_5861,N_5914);
nor U6104 (N_6104,N_5864,N_5808);
nor U6105 (N_6105,N_5928,N_5917);
and U6106 (N_6106,N_5839,N_5902);
xnor U6107 (N_6107,N_5820,N_5879);
or U6108 (N_6108,N_5797,N_5842);
and U6109 (N_6109,N_5885,N_5758);
xor U6110 (N_6110,N_5893,N_5750);
or U6111 (N_6111,N_5853,N_5819);
nand U6112 (N_6112,N_5795,N_5823);
nand U6113 (N_6113,N_5812,N_5900);
xor U6114 (N_6114,N_5778,N_5925);
nand U6115 (N_6115,N_5899,N_5832);
nor U6116 (N_6116,N_5781,N_5813);
nor U6117 (N_6117,N_5918,N_5955);
nor U6118 (N_6118,N_5971,N_5919);
nor U6119 (N_6119,N_5957,N_5985);
or U6120 (N_6120,N_5790,N_5824);
nor U6121 (N_6121,N_5951,N_5792);
or U6122 (N_6122,N_5921,N_5789);
or U6123 (N_6123,N_5801,N_5757);
and U6124 (N_6124,N_5867,N_5836);
and U6125 (N_6125,N_5921,N_5991);
or U6126 (N_6126,N_5756,N_5814);
nor U6127 (N_6127,N_5881,N_5802);
and U6128 (N_6128,N_5910,N_5751);
or U6129 (N_6129,N_5777,N_5821);
nand U6130 (N_6130,N_5774,N_5956);
or U6131 (N_6131,N_5767,N_5830);
and U6132 (N_6132,N_5789,N_5893);
nand U6133 (N_6133,N_5935,N_5782);
nand U6134 (N_6134,N_5880,N_5955);
and U6135 (N_6135,N_5910,N_5923);
or U6136 (N_6136,N_5859,N_5825);
nand U6137 (N_6137,N_5829,N_5963);
nand U6138 (N_6138,N_5751,N_5880);
or U6139 (N_6139,N_5811,N_5805);
xnor U6140 (N_6140,N_5818,N_5907);
xnor U6141 (N_6141,N_5872,N_5764);
nor U6142 (N_6142,N_5843,N_5982);
nand U6143 (N_6143,N_5767,N_5915);
nand U6144 (N_6144,N_5942,N_5775);
nor U6145 (N_6145,N_5822,N_5984);
nor U6146 (N_6146,N_5767,N_5936);
and U6147 (N_6147,N_5848,N_5996);
nor U6148 (N_6148,N_5962,N_5845);
and U6149 (N_6149,N_5822,N_5910);
nor U6150 (N_6150,N_5894,N_5963);
nor U6151 (N_6151,N_5962,N_5931);
or U6152 (N_6152,N_5971,N_5939);
nor U6153 (N_6153,N_5867,N_5965);
and U6154 (N_6154,N_5838,N_5784);
or U6155 (N_6155,N_5769,N_5862);
nor U6156 (N_6156,N_5763,N_5794);
nor U6157 (N_6157,N_5957,N_5766);
nor U6158 (N_6158,N_5797,N_5878);
or U6159 (N_6159,N_5955,N_5850);
nor U6160 (N_6160,N_5976,N_5964);
nor U6161 (N_6161,N_5837,N_5929);
xor U6162 (N_6162,N_5768,N_5933);
nor U6163 (N_6163,N_5831,N_5923);
nor U6164 (N_6164,N_5807,N_5841);
and U6165 (N_6165,N_5816,N_5912);
nand U6166 (N_6166,N_5994,N_5992);
nand U6167 (N_6167,N_5874,N_5986);
or U6168 (N_6168,N_5752,N_5825);
nor U6169 (N_6169,N_5794,N_5996);
and U6170 (N_6170,N_5764,N_5787);
or U6171 (N_6171,N_5782,N_5875);
nand U6172 (N_6172,N_5854,N_5827);
nand U6173 (N_6173,N_5841,N_5877);
nand U6174 (N_6174,N_5901,N_5853);
nand U6175 (N_6175,N_5783,N_5803);
nand U6176 (N_6176,N_5792,N_5966);
xor U6177 (N_6177,N_5838,N_5759);
nand U6178 (N_6178,N_5909,N_5954);
and U6179 (N_6179,N_5823,N_5951);
and U6180 (N_6180,N_5760,N_5763);
or U6181 (N_6181,N_5790,N_5992);
nand U6182 (N_6182,N_5865,N_5873);
nor U6183 (N_6183,N_5830,N_5848);
nand U6184 (N_6184,N_5989,N_5770);
nor U6185 (N_6185,N_5983,N_5945);
nor U6186 (N_6186,N_5978,N_5967);
and U6187 (N_6187,N_5825,N_5804);
nand U6188 (N_6188,N_5996,N_5770);
or U6189 (N_6189,N_5762,N_5955);
xor U6190 (N_6190,N_5921,N_5784);
or U6191 (N_6191,N_5828,N_5830);
nand U6192 (N_6192,N_5921,N_5838);
and U6193 (N_6193,N_5911,N_5830);
and U6194 (N_6194,N_5805,N_5945);
and U6195 (N_6195,N_5777,N_5802);
nor U6196 (N_6196,N_5824,N_5834);
and U6197 (N_6197,N_5966,N_5923);
or U6198 (N_6198,N_5930,N_5830);
nand U6199 (N_6199,N_5934,N_5770);
nand U6200 (N_6200,N_5862,N_5843);
nand U6201 (N_6201,N_5844,N_5871);
nor U6202 (N_6202,N_5964,N_5856);
xor U6203 (N_6203,N_5899,N_5915);
or U6204 (N_6204,N_5867,N_5931);
or U6205 (N_6205,N_5842,N_5939);
and U6206 (N_6206,N_5800,N_5771);
nand U6207 (N_6207,N_5938,N_5917);
nor U6208 (N_6208,N_5872,N_5833);
nand U6209 (N_6209,N_5927,N_5993);
and U6210 (N_6210,N_5840,N_5892);
nor U6211 (N_6211,N_5834,N_5773);
or U6212 (N_6212,N_5883,N_5805);
and U6213 (N_6213,N_5754,N_5988);
nand U6214 (N_6214,N_5970,N_5831);
and U6215 (N_6215,N_5900,N_5868);
nor U6216 (N_6216,N_5935,N_5871);
nor U6217 (N_6217,N_5973,N_5915);
and U6218 (N_6218,N_5888,N_5861);
or U6219 (N_6219,N_5883,N_5919);
nor U6220 (N_6220,N_5777,N_5805);
nand U6221 (N_6221,N_5818,N_5951);
xor U6222 (N_6222,N_5865,N_5768);
nand U6223 (N_6223,N_5799,N_5848);
nand U6224 (N_6224,N_5914,N_5834);
nand U6225 (N_6225,N_5904,N_5912);
and U6226 (N_6226,N_5773,N_5878);
nand U6227 (N_6227,N_5817,N_5936);
xnor U6228 (N_6228,N_5995,N_5921);
nand U6229 (N_6229,N_5914,N_5991);
nor U6230 (N_6230,N_5957,N_5800);
or U6231 (N_6231,N_5820,N_5988);
or U6232 (N_6232,N_5799,N_5827);
nand U6233 (N_6233,N_5958,N_5875);
nor U6234 (N_6234,N_5803,N_5824);
nand U6235 (N_6235,N_5756,N_5924);
nand U6236 (N_6236,N_5875,N_5932);
nor U6237 (N_6237,N_5786,N_5842);
nor U6238 (N_6238,N_5785,N_5910);
nor U6239 (N_6239,N_5844,N_5964);
nand U6240 (N_6240,N_5803,N_5896);
and U6241 (N_6241,N_5914,N_5898);
nor U6242 (N_6242,N_5853,N_5953);
nand U6243 (N_6243,N_5961,N_5824);
or U6244 (N_6244,N_5989,N_5913);
or U6245 (N_6245,N_5782,N_5849);
and U6246 (N_6246,N_5975,N_5943);
and U6247 (N_6247,N_5814,N_5853);
or U6248 (N_6248,N_5876,N_5979);
and U6249 (N_6249,N_5829,N_5855);
and U6250 (N_6250,N_6029,N_6014);
nor U6251 (N_6251,N_6080,N_6131);
or U6252 (N_6252,N_6206,N_6141);
and U6253 (N_6253,N_6050,N_6061);
and U6254 (N_6254,N_6181,N_6073);
nor U6255 (N_6255,N_6126,N_6017);
nand U6256 (N_6256,N_6169,N_6196);
or U6257 (N_6257,N_6113,N_6128);
xnor U6258 (N_6258,N_6164,N_6214);
nand U6259 (N_6259,N_6026,N_6237);
and U6260 (N_6260,N_6154,N_6204);
nor U6261 (N_6261,N_6203,N_6124);
and U6262 (N_6262,N_6163,N_6143);
nor U6263 (N_6263,N_6059,N_6069);
xor U6264 (N_6264,N_6234,N_6092);
nor U6265 (N_6265,N_6081,N_6127);
and U6266 (N_6266,N_6117,N_6135);
and U6267 (N_6267,N_6082,N_6111);
nand U6268 (N_6268,N_6040,N_6220);
or U6269 (N_6269,N_6183,N_6245);
nor U6270 (N_6270,N_6200,N_6098);
and U6271 (N_6271,N_6149,N_6132);
nand U6272 (N_6272,N_6019,N_6074);
and U6273 (N_6273,N_6032,N_6167);
xor U6274 (N_6274,N_6025,N_6108);
and U6275 (N_6275,N_6170,N_6065);
nor U6276 (N_6276,N_6036,N_6104);
and U6277 (N_6277,N_6052,N_6191);
and U6278 (N_6278,N_6148,N_6001);
or U6279 (N_6279,N_6178,N_6186);
and U6280 (N_6280,N_6102,N_6229);
nor U6281 (N_6281,N_6125,N_6142);
nor U6282 (N_6282,N_6194,N_6071);
nor U6283 (N_6283,N_6209,N_6168);
or U6284 (N_6284,N_6175,N_6248);
xor U6285 (N_6285,N_6227,N_6153);
xnor U6286 (N_6286,N_6095,N_6078);
nand U6287 (N_6287,N_6043,N_6010);
and U6288 (N_6288,N_6156,N_6101);
and U6289 (N_6289,N_6249,N_6039);
or U6290 (N_6290,N_6027,N_6097);
nand U6291 (N_6291,N_6212,N_6116);
xnor U6292 (N_6292,N_6075,N_6244);
nand U6293 (N_6293,N_6179,N_6042);
nor U6294 (N_6294,N_6151,N_6201);
nor U6295 (N_6295,N_6195,N_6031);
nand U6296 (N_6296,N_6083,N_6238);
and U6297 (N_6297,N_6005,N_6112);
nand U6298 (N_6298,N_6165,N_6003);
nand U6299 (N_6299,N_6033,N_6011);
nand U6300 (N_6300,N_6147,N_6016);
nand U6301 (N_6301,N_6187,N_6085);
or U6302 (N_6302,N_6066,N_6138);
nand U6303 (N_6303,N_6241,N_6225);
nor U6304 (N_6304,N_6094,N_6051);
xnor U6305 (N_6305,N_6224,N_6103);
and U6306 (N_6306,N_6119,N_6202);
and U6307 (N_6307,N_6217,N_6106);
nand U6308 (N_6308,N_6107,N_6110);
nand U6309 (N_6309,N_6053,N_6122);
nand U6310 (N_6310,N_6062,N_6037);
nor U6311 (N_6311,N_6063,N_6197);
xor U6312 (N_6312,N_6172,N_6159);
or U6313 (N_6313,N_6022,N_6076);
nand U6314 (N_6314,N_6171,N_6048);
xnor U6315 (N_6315,N_6176,N_6049);
or U6316 (N_6316,N_6034,N_6079);
nand U6317 (N_6317,N_6060,N_6155);
and U6318 (N_6318,N_6058,N_6247);
and U6319 (N_6319,N_6038,N_6089);
nor U6320 (N_6320,N_6077,N_6223);
and U6321 (N_6321,N_6246,N_6002);
and U6322 (N_6322,N_6045,N_6231);
xnor U6323 (N_6323,N_6193,N_6158);
nand U6324 (N_6324,N_6152,N_6160);
nand U6325 (N_6325,N_6177,N_6232);
or U6326 (N_6326,N_6230,N_6161);
or U6327 (N_6327,N_6144,N_6012);
or U6328 (N_6328,N_6054,N_6235);
nand U6329 (N_6329,N_6105,N_6030);
and U6330 (N_6330,N_6180,N_6162);
nand U6331 (N_6331,N_6024,N_6174);
and U6332 (N_6332,N_6188,N_6136);
xor U6333 (N_6333,N_6004,N_6211);
or U6334 (N_6334,N_6219,N_6129);
nand U6335 (N_6335,N_6087,N_6057);
or U6336 (N_6336,N_6046,N_6222);
or U6337 (N_6337,N_6064,N_6086);
or U6338 (N_6338,N_6173,N_6099);
nand U6339 (N_6339,N_6134,N_6166);
nand U6340 (N_6340,N_6150,N_6013);
nand U6341 (N_6341,N_6228,N_6157);
and U6342 (N_6342,N_6198,N_6121);
nor U6343 (N_6343,N_6139,N_6130);
nor U6344 (N_6344,N_6006,N_6044);
nand U6345 (N_6345,N_6226,N_6239);
nand U6346 (N_6346,N_6015,N_6115);
nor U6347 (N_6347,N_6123,N_6182);
or U6348 (N_6348,N_6096,N_6120);
nor U6349 (N_6349,N_6047,N_6137);
nor U6350 (N_6350,N_6190,N_6100);
nor U6351 (N_6351,N_6146,N_6207);
and U6352 (N_6352,N_6213,N_6242);
nand U6353 (N_6353,N_6091,N_6199);
or U6354 (N_6354,N_6072,N_6210);
xor U6355 (N_6355,N_6218,N_6090);
or U6356 (N_6356,N_6185,N_6068);
xnor U6357 (N_6357,N_6093,N_6215);
and U6358 (N_6358,N_6133,N_6020);
or U6359 (N_6359,N_6055,N_6084);
nor U6360 (N_6360,N_6221,N_6118);
and U6361 (N_6361,N_6041,N_6000);
nand U6362 (N_6362,N_6009,N_6067);
nand U6363 (N_6363,N_6184,N_6140);
and U6364 (N_6364,N_6243,N_6145);
nor U6365 (N_6365,N_6008,N_6240);
and U6366 (N_6366,N_6018,N_6021);
xnor U6367 (N_6367,N_6088,N_6192);
or U6368 (N_6368,N_6208,N_6007);
xor U6369 (N_6369,N_6109,N_6056);
nor U6370 (N_6370,N_6189,N_6236);
or U6371 (N_6371,N_6070,N_6028);
nor U6372 (N_6372,N_6216,N_6205);
or U6373 (N_6373,N_6114,N_6233);
nor U6374 (N_6374,N_6035,N_6023);
and U6375 (N_6375,N_6026,N_6094);
or U6376 (N_6376,N_6201,N_6027);
or U6377 (N_6377,N_6055,N_6067);
or U6378 (N_6378,N_6053,N_6163);
and U6379 (N_6379,N_6034,N_6170);
xnor U6380 (N_6380,N_6220,N_6191);
and U6381 (N_6381,N_6141,N_6136);
nor U6382 (N_6382,N_6224,N_6090);
nand U6383 (N_6383,N_6191,N_6038);
xor U6384 (N_6384,N_6115,N_6176);
nor U6385 (N_6385,N_6050,N_6073);
and U6386 (N_6386,N_6050,N_6144);
nor U6387 (N_6387,N_6159,N_6163);
or U6388 (N_6388,N_6091,N_6057);
xor U6389 (N_6389,N_6055,N_6157);
nand U6390 (N_6390,N_6144,N_6020);
or U6391 (N_6391,N_6146,N_6201);
or U6392 (N_6392,N_6188,N_6063);
and U6393 (N_6393,N_6009,N_6231);
or U6394 (N_6394,N_6021,N_6077);
and U6395 (N_6395,N_6228,N_6184);
and U6396 (N_6396,N_6066,N_6027);
and U6397 (N_6397,N_6096,N_6067);
and U6398 (N_6398,N_6233,N_6159);
nor U6399 (N_6399,N_6160,N_6225);
and U6400 (N_6400,N_6164,N_6165);
and U6401 (N_6401,N_6249,N_6206);
xor U6402 (N_6402,N_6154,N_6147);
and U6403 (N_6403,N_6208,N_6186);
nor U6404 (N_6404,N_6214,N_6014);
nor U6405 (N_6405,N_6093,N_6103);
nand U6406 (N_6406,N_6093,N_6186);
nand U6407 (N_6407,N_6229,N_6162);
and U6408 (N_6408,N_6083,N_6048);
and U6409 (N_6409,N_6083,N_6065);
xnor U6410 (N_6410,N_6187,N_6172);
or U6411 (N_6411,N_6231,N_6142);
and U6412 (N_6412,N_6126,N_6117);
and U6413 (N_6413,N_6036,N_6035);
and U6414 (N_6414,N_6031,N_6179);
nor U6415 (N_6415,N_6030,N_6118);
and U6416 (N_6416,N_6123,N_6154);
xnor U6417 (N_6417,N_6194,N_6135);
or U6418 (N_6418,N_6136,N_6101);
and U6419 (N_6419,N_6003,N_6237);
nor U6420 (N_6420,N_6164,N_6040);
nor U6421 (N_6421,N_6099,N_6221);
and U6422 (N_6422,N_6042,N_6209);
or U6423 (N_6423,N_6160,N_6033);
or U6424 (N_6424,N_6140,N_6101);
and U6425 (N_6425,N_6196,N_6150);
nand U6426 (N_6426,N_6003,N_6214);
nand U6427 (N_6427,N_6041,N_6190);
nor U6428 (N_6428,N_6117,N_6249);
xor U6429 (N_6429,N_6135,N_6088);
and U6430 (N_6430,N_6111,N_6180);
and U6431 (N_6431,N_6068,N_6077);
nor U6432 (N_6432,N_6037,N_6234);
nand U6433 (N_6433,N_6188,N_6088);
nor U6434 (N_6434,N_6216,N_6062);
or U6435 (N_6435,N_6035,N_6096);
and U6436 (N_6436,N_6055,N_6166);
and U6437 (N_6437,N_6078,N_6007);
and U6438 (N_6438,N_6062,N_6228);
nand U6439 (N_6439,N_6129,N_6011);
xor U6440 (N_6440,N_6098,N_6027);
nand U6441 (N_6441,N_6221,N_6207);
or U6442 (N_6442,N_6220,N_6024);
nor U6443 (N_6443,N_6084,N_6044);
and U6444 (N_6444,N_6145,N_6002);
nor U6445 (N_6445,N_6109,N_6187);
or U6446 (N_6446,N_6211,N_6171);
or U6447 (N_6447,N_6090,N_6247);
and U6448 (N_6448,N_6118,N_6119);
nand U6449 (N_6449,N_6046,N_6193);
nor U6450 (N_6450,N_6192,N_6090);
or U6451 (N_6451,N_6234,N_6182);
nand U6452 (N_6452,N_6152,N_6215);
and U6453 (N_6453,N_6216,N_6247);
nand U6454 (N_6454,N_6156,N_6224);
or U6455 (N_6455,N_6082,N_6041);
or U6456 (N_6456,N_6085,N_6157);
nor U6457 (N_6457,N_6119,N_6219);
nand U6458 (N_6458,N_6188,N_6124);
xor U6459 (N_6459,N_6153,N_6031);
xor U6460 (N_6460,N_6136,N_6191);
or U6461 (N_6461,N_6201,N_6148);
or U6462 (N_6462,N_6112,N_6052);
nand U6463 (N_6463,N_6156,N_6084);
nor U6464 (N_6464,N_6147,N_6139);
nor U6465 (N_6465,N_6074,N_6061);
and U6466 (N_6466,N_6061,N_6112);
nor U6467 (N_6467,N_6044,N_6086);
xor U6468 (N_6468,N_6164,N_6043);
nor U6469 (N_6469,N_6137,N_6075);
nor U6470 (N_6470,N_6151,N_6004);
or U6471 (N_6471,N_6212,N_6026);
nor U6472 (N_6472,N_6226,N_6171);
or U6473 (N_6473,N_6182,N_6118);
nor U6474 (N_6474,N_6027,N_6110);
or U6475 (N_6475,N_6022,N_6122);
and U6476 (N_6476,N_6053,N_6146);
and U6477 (N_6477,N_6026,N_6201);
and U6478 (N_6478,N_6033,N_6233);
and U6479 (N_6479,N_6087,N_6109);
or U6480 (N_6480,N_6197,N_6028);
nand U6481 (N_6481,N_6239,N_6032);
nor U6482 (N_6482,N_6181,N_6173);
xnor U6483 (N_6483,N_6032,N_6011);
nor U6484 (N_6484,N_6073,N_6112);
nand U6485 (N_6485,N_6135,N_6147);
and U6486 (N_6486,N_6058,N_6006);
nor U6487 (N_6487,N_6117,N_6012);
or U6488 (N_6488,N_6150,N_6123);
nor U6489 (N_6489,N_6244,N_6030);
nand U6490 (N_6490,N_6056,N_6012);
nor U6491 (N_6491,N_6023,N_6021);
nand U6492 (N_6492,N_6102,N_6083);
or U6493 (N_6493,N_6196,N_6014);
nand U6494 (N_6494,N_6231,N_6111);
and U6495 (N_6495,N_6043,N_6183);
or U6496 (N_6496,N_6017,N_6045);
and U6497 (N_6497,N_6162,N_6066);
and U6498 (N_6498,N_6213,N_6065);
nand U6499 (N_6499,N_6052,N_6126);
or U6500 (N_6500,N_6266,N_6265);
nand U6501 (N_6501,N_6494,N_6328);
or U6502 (N_6502,N_6286,N_6453);
nand U6503 (N_6503,N_6379,N_6438);
or U6504 (N_6504,N_6425,N_6430);
nor U6505 (N_6505,N_6389,N_6352);
and U6506 (N_6506,N_6427,N_6419);
and U6507 (N_6507,N_6472,N_6468);
nor U6508 (N_6508,N_6480,N_6481);
or U6509 (N_6509,N_6339,N_6340);
nand U6510 (N_6510,N_6489,N_6254);
nand U6511 (N_6511,N_6457,N_6487);
xor U6512 (N_6512,N_6293,N_6261);
nor U6513 (N_6513,N_6308,N_6269);
and U6514 (N_6514,N_6448,N_6406);
and U6515 (N_6515,N_6292,N_6374);
and U6516 (N_6516,N_6315,N_6385);
xnor U6517 (N_6517,N_6280,N_6417);
nand U6518 (N_6518,N_6362,N_6262);
and U6519 (N_6519,N_6402,N_6257);
nor U6520 (N_6520,N_6264,N_6253);
or U6521 (N_6521,N_6287,N_6310);
xnor U6522 (N_6522,N_6459,N_6356);
or U6523 (N_6523,N_6268,N_6482);
or U6524 (N_6524,N_6333,N_6358);
or U6525 (N_6525,N_6329,N_6445);
or U6526 (N_6526,N_6289,N_6450);
nor U6527 (N_6527,N_6386,N_6346);
nand U6528 (N_6528,N_6475,N_6439);
nor U6529 (N_6529,N_6449,N_6336);
xnor U6530 (N_6530,N_6321,N_6442);
xor U6531 (N_6531,N_6258,N_6277);
or U6532 (N_6532,N_6460,N_6357);
nor U6533 (N_6533,N_6461,N_6276);
and U6534 (N_6534,N_6484,N_6377);
nand U6535 (N_6535,N_6278,N_6476);
nand U6536 (N_6536,N_6365,N_6473);
nor U6537 (N_6537,N_6413,N_6361);
nand U6538 (N_6538,N_6320,N_6426);
and U6539 (N_6539,N_6465,N_6313);
nor U6540 (N_6540,N_6334,N_6327);
xnor U6541 (N_6541,N_6429,N_6309);
or U6542 (N_6542,N_6302,N_6479);
or U6543 (N_6543,N_6466,N_6314);
nor U6544 (N_6544,N_6298,N_6434);
or U6545 (N_6545,N_6397,N_6267);
and U6546 (N_6546,N_6441,N_6422);
nand U6547 (N_6547,N_6281,N_6279);
nand U6548 (N_6548,N_6393,N_6364);
nand U6549 (N_6549,N_6355,N_6300);
nand U6550 (N_6550,N_6395,N_6363);
and U6551 (N_6551,N_6478,N_6458);
nand U6552 (N_6552,N_6431,N_6295);
or U6553 (N_6553,N_6491,N_6440);
or U6554 (N_6554,N_6303,N_6291);
or U6555 (N_6555,N_6285,N_6403);
nor U6556 (N_6556,N_6273,N_6326);
or U6557 (N_6557,N_6490,N_6260);
and U6558 (N_6558,N_6366,N_6477);
nor U6559 (N_6559,N_6433,N_6437);
nor U6560 (N_6560,N_6367,N_6250);
and U6561 (N_6561,N_6414,N_6432);
nor U6562 (N_6562,N_6497,N_6387);
or U6563 (N_6563,N_6488,N_6469);
and U6564 (N_6564,N_6288,N_6330);
xor U6565 (N_6565,N_6446,N_6272);
nand U6566 (N_6566,N_6408,N_6350);
or U6567 (N_6567,N_6255,N_6375);
nand U6568 (N_6568,N_6382,N_6470);
nor U6569 (N_6569,N_6380,N_6451);
nor U6570 (N_6570,N_6462,N_6322);
nand U6571 (N_6571,N_6370,N_6349);
and U6572 (N_6572,N_6405,N_6492);
or U6573 (N_6573,N_6259,N_6332);
nand U6574 (N_6574,N_6398,N_6344);
and U6575 (N_6575,N_6455,N_6400);
or U6576 (N_6576,N_6467,N_6353);
nor U6577 (N_6577,N_6368,N_6407);
nor U6578 (N_6578,N_6369,N_6474);
or U6579 (N_6579,N_6456,N_6390);
nand U6580 (N_6580,N_6428,N_6270);
nor U6581 (N_6581,N_6415,N_6495);
or U6582 (N_6582,N_6274,N_6294);
and U6583 (N_6583,N_6323,N_6391);
nand U6584 (N_6584,N_6401,N_6411);
nand U6585 (N_6585,N_6435,N_6372);
nand U6586 (N_6586,N_6483,N_6307);
nor U6587 (N_6587,N_6409,N_6452);
and U6588 (N_6588,N_6373,N_6486);
or U6589 (N_6589,N_6394,N_6283);
and U6590 (N_6590,N_6423,N_6347);
and U6591 (N_6591,N_6454,N_6381);
or U6592 (N_6592,N_6444,N_6399);
nor U6593 (N_6593,N_6421,N_6324);
nor U6594 (N_6594,N_6263,N_6348);
or U6595 (N_6595,N_6360,N_6338);
nand U6596 (N_6596,N_6284,N_6376);
nand U6597 (N_6597,N_6384,N_6341);
or U6598 (N_6598,N_6464,N_6251);
nand U6599 (N_6599,N_6316,N_6256);
or U6600 (N_6600,N_6335,N_6297);
xnor U6601 (N_6601,N_6290,N_6304);
nor U6602 (N_6602,N_6371,N_6359);
or U6603 (N_6603,N_6337,N_6404);
nor U6604 (N_6604,N_6319,N_6392);
nor U6605 (N_6605,N_6443,N_6299);
nor U6606 (N_6606,N_6396,N_6282);
xnor U6607 (N_6607,N_6418,N_6447);
nand U6608 (N_6608,N_6252,N_6424);
nor U6609 (N_6609,N_6416,N_6351);
and U6610 (N_6610,N_6345,N_6463);
nand U6611 (N_6611,N_6343,N_6498);
and U6612 (N_6612,N_6378,N_6410);
nor U6613 (N_6613,N_6325,N_6296);
nand U6614 (N_6614,N_6354,N_6485);
nor U6615 (N_6615,N_6420,N_6342);
and U6616 (N_6616,N_6312,N_6301);
or U6617 (N_6617,N_6499,N_6436);
nand U6618 (N_6618,N_6331,N_6496);
nand U6619 (N_6619,N_6271,N_6318);
or U6620 (N_6620,N_6317,N_6471);
nand U6621 (N_6621,N_6412,N_6388);
and U6622 (N_6622,N_6305,N_6383);
nand U6623 (N_6623,N_6275,N_6311);
nor U6624 (N_6624,N_6306,N_6493);
or U6625 (N_6625,N_6351,N_6281);
or U6626 (N_6626,N_6303,N_6321);
nand U6627 (N_6627,N_6405,N_6309);
or U6628 (N_6628,N_6363,N_6378);
nor U6629 (N_6629,N_6361,N_6468);
or U6630 (N_6630,N_6361,N_6387);
nand U6631 (N_6631,N_6336,N_6290);
nor U6632 (N_6632,N_6361,N_6363);
nor U6633 (N_6633,N_6472,N_6250);
nand U6634 (N_6634,N_6449,N_6275);
xor U6635 (N_6635,N_6290,N_6414);
or U6636 (N_6636,N_6462,N_6385);
and U6637 (N_6637,N_6385,N_6425);
nor U6638 (N_6638,N_6344,N_6427);
xnor U6639 (N_6639,N_6347,N_6270);
xor U6640 (N_6640,N_6499,N_6331);
or U6641 (N_6641,N_6440,N_6341);
xor U6642 (N_6642,N_6291,N_6322);
xnor U6643 (N_6643,N_6474,N_6392);
and U6644 (N_6644,N_6482,N_6393);
nor U6645 (N_6645,N_6294,N_6411);
nand U6646 (N_6646,N_6392,N_6252);
nor U6647 (N_6647,N_6452,N_6278);
nand U6648 (N_6648,N_6407,N_6452);
and U6649 (N_6649,N_6317,N_6414);
nor U6650 (N_6650,N_6401,N_6422);
or U6651 (N_6651,N_6264,N_6477);
xnor U6652 (N_6652,N_6424,N_6461);
nand U6653 (N_6653,N_6380,N_6350);
and U6654 (N_6654,N_6299,N_6414);
or U6655 (N_6655,N_6431,N_6488);
nor U6656 (N_6656,N_6306,N_6495);
nand U6657 (N_6657,N_6487,N_6368);
nand U6658 (N_6658,N_6272,N_6496);
nand U6659 (N_6659,N_6263,N_6435);
and U6660 (N_6660,N_6306,N_6423);
or U6661 (N_6661,N_6427,N_6365);
or U6662 (N_6662,N_6334,N_6315);
or U6663 (N_6663,N_6432,N_6337);
and U6664 (N_6664,N_6377,N_6307);
xor U6665 (N_6665,N_6313,N_6373);
or U6666 (N_6666,N_6305,N_6493);
nand U6667 (N_6667,N_6286,N_6442);
xor U6668 (N_6668,N_6341,N_6488);
and U6669 (N_6669,N_6495,N_6471);
and U6670 (N_6670,N_6312,N_6267);
nand U6671 (N_6671,N_6309,N_6384);
nand U6672 (N_6672,N_6395,N_6364);
nand U6673 (N_6673,N_6404,N_6269);
nor U6674 (N_6674,N_6454,N_6256);
or U6675 (N_6675,N_6256,N_6433);
nand U6676 (N_6676,N_6489,N_6261);
nor U6677 (N_6677,N_6392,N_6450);
nor U6678 (N_6678,N_6314,N_6441);
and U6679 (N_6679,N_6293,N_6262);
and U6680 (N_6680,N_6365,N_6471);
and U6681 (N_6681,N_6347,N_6398);
and U6682 (N_6682,N_6289,N_6302);
and U6683 (N_6683,N_6415,N_6428);
or U6684 (N_6684,N_6383,N_6409);
or U6685 (N_6685,N_6402,N_6401);
and U6686 (N_6686,N_6270,N_6388);
nand U6687 (N_6687,N_6319,N_6451);
xor U6688 (N_6688,N_6274,N_6493);
nor U6689 (N_6689,N_6484,N_6417);
xor U6690 (N_6690,N_6337,N_6495);
or U6691 (N_6691,N_6417,N_6378);
and U6692 (N_6692,N_6490,N_6409);
or U6693 (N_6693,N_6491,N_6438);
or U6694 (N_6694,N_6489,N_6378);
nand U6695 (N_6695,N_6310,N_6305);
nor U6696 (N_6696,N_6342,N_6446);
nand U6697 (N_6697,N_6289,N_6272);
nor U6698 (N_6698,N_6321,N_6390);
and U6699 (N_6699,N_6261,N_6307);
xor U6700 (N_6700,N_6254,N_6345);
nor U6701 (N_6701,N_6262,N_6445);
nor U6702 (N_6702,N_6396,N_6422);
nor U6703 (N_6703,N_6303,N_6476);
and U6704 (N_6704,N_6472,N_6397);
nand U6705 (N_6705,N_6410,N_6296);
and U6706 (N_6706,N_6402,N_6497);
or U6707 (N_6707,N_6453,N_6325);
xnor U6708 (N_6708,N_6414,N_6391);
nand U6709 (N_6709,N_6422,N_6361);
nor U6710 (N_6710,N_6390,N_6404);
or U6711 (N_6711,N_6302,N_6396);
xnor U6712 (N_6712,N_6489,N_6333);
nand U6713 (N_6713,N_6263,N_6424);
nand U6714 (N_6714,N_6356,N_6319);
or U6715 (N_6715,N_6283,N_6365);
nor U6716 (N_6716,N_6344,N_6411);
and U6717 (N_6717,N_6312,N_6302);
nor U6718 (N_6718,N_6468,N_6380);
nand U6719 (N_6719,N_6464,N_6286);
nand U6720 (N_6720,N_6425,N_6289);
nor U6721 (N_6721,N_6256,N_6425);
xnor U6722 (N_6722,N_6487,N_6431);
nand U6723 (N_6723,N_6371,N_6313);
or U6724 (N_6724,N_6492,N_6379);
nand U6725 (N_6725,N_6405,N_6260);
nand U6726 (N_6726,N_6442,N_6384);
or U6727 (N_6727,N_6487,N_6325);
nor U6728 (N_6728,N_6410,N_6438);
or U6729 (N_6729,N_6447,N_6398);
and U6730 (N_6730,N_6318,N_6385);
nand U6731 (N_6731,N_6481,N_6390);
xor U6732 (N_6732,N_6284,N_6259);
and U6733 (N_6733,N_6283,N_6357);
xnor U6734 (N_6734,N_6322,N_6481);
xnor U6735 (N_6735,N_6262,N_6469);
and U6736 (N_6736,N_6389,N_6357);
nand U6737 (N_6737,N_6254,N_6359);
xor U6738 (N_6738,N_6344,N_6261);
or U6739 (N_6739,N_6272,N_6455);
nor U6740 (N_6740,N_6388,N_6481);
nand U6741 (N_6741,N_6284,N_6455);
nand U6742 (N_6742,N_6455,N_6363);
and U6743 (N_6743,N_6471,N_6330);
nand U6744 (N_6744,N_6439,N_6345);
or U6745 (N_6745,N_6371,N_6348);
nor U6746 (N_6746,N_6482,N_6433);
xnor U6747 (N_6747,N_6335,N_6444);
or U6748 (N_6748,N_6498,N_6486);
xor U6749 (N_6749,N_6283,N_6345);
and U6750 (N_6750,N_6590,N_6722);
or U6751 (N_6751,N_6716,N_6516);
or U6752 (N_6752,N_6669,N_6537);
nand U6753 (N_6753,N_6707,N_6515);
or U6754 (N_6754,N_6552,N_6731);
or U6755 (N_6755,N_6622,N_6583);
or U6756 (N_6756,N_6738,N_6723);
nor U6757 (N_6757,N_6545,N_6571);
and U6758 (N_6758,N_6619,N_6673);
nor U6759 (N_6759,N_6608,N_6713);
and U6760 (N_6760,N_6726,N_6648);
nor U6761 (N_6761,N_6565,N_6542);
nand U6762 (N_6762,N_6572,N_6748);
or U6763 (N_6763,N_6640,N_6609);
nand U6764 (N_6764,N_6543,N_6501);
nor U6765 (N_6765,N_6574,N_6714);
nor U6766 (N_6766,N_6536,N_6626);
and U6767 (N_6767,N_6560,N_6715);
nand U6768 (N_6768,N_6682,N_6503);
nand U6769 (N_6769,N_6656,N_6676);
and U6770 (N_6770,N_6539,N_6602);
nor U6771 (N_6771,N_6595,N_6576);
xnor U6772 (N_6772,N_6693,N_6559);
and U6773 (N_6773,N_6548,N_6521);
xor U6774 (N_6774,N_6564,N_6652);
nand U6775 (N_6775,N_6677,N_6613);
and U6776 (N_6776,N_6687,N_6581);
and U6777 (N_6777,N_6724,N_6621);
xnor U6778 (N_6778,N_6528,N_6554);
nor U6779 (N_6779,N_6584,N_6502);
and U6780 (N_6780,N_6585,N_6627);
and U6781 (N_6781,N_6728,N_6566);
nand U6782 (N_6782,N_6667,N_6629);
nand U6783 (N_6783,N_6586,N_6601);
or U6784 (N_6784,N_6558,N_6591);
or U6785 (N_6785,N_6665,N_6527);
nand U6786 (N_6786,N_6674,N_6596);
nand U6787 (N_6787,N_6678,N_6697);
xor U6788 (N_6788,N_6611,N_6700);
nor U6789 (N_6789,N_6645,N_6523);
nor U6790 (N_6790,N_6742,N_6637);
xor U6791 (N_6791,N_6568,N_6681);
and U6792 (N_6792,N_6685,N_6666);
nor U6793 (N_6793,N_6517,N_6524);
nand U6794 (N_6794,N_6617,N_6510);
or U6795 (N_6795,N_6746,N_6598);
nand U6796 (N_6796,N_6535,N_6634);
and U6797 (N_6797,N_6551,N_6671);
xnor U6798 (N_6798,N_6507,N_6506);
nor U6799 (N_6799,N_6557,N_6698);
and U6800 (N_6800,N_6588,N_6610);
and U6801 (N_6801,N_6513,N_6623);
and U6802 (N_6802,N_6725,N_6604);
or U6803 (N_6803,N_6544,N_6691);
and U6804 (N_6804,N_6658,N_6555);
nand U6805 (N_6805,N_6597,N_6683);
nand U6806 (N_6806,N_6546,N_6540);
nand U6807 (N_6807,N_6508,N_6525);
nand U6808 (N_6808,N_6662,N_6628);
and U6809 (N_6809,N_6547,N_6708);
or U6810 (N_6810,N_6643,N_6538);
nand U6811 (N_6811,N_6589,N_6570);
and U6812 (N_6812,N_6733,N_6680);
or U6813 (N_6813,N_6718,N_6519);
nor U6814 (N_6814,N_6741,N_6573);
xor U6815 (N_6815,N_6630,N_6654);
and U6816 (N_6816,N_6605,N_6672);
nor U6817 (N_6817,N_6730,N_6679);
nand U6818 (N_6818,N_6534,N_6531);
xnor U6819 (N_6819,N_6655,N_6749);
xnor U6820 (N_6820,N_6578,N_6704);
nor U6821 (N_6821,N_6661,N_6744);
nand U6822 (N_6822,N_6633,N_6532);
nor U6823 (N_6823,N_6505,N_6651);
or U6824 (N_6824,N_6603,N_6659);
and U6825 (N_6825,N_6694,N_6689);
or U6826 (N_6826,N_6699,N_6561);
and U6827 (N_6827,N_6549,N_6649);
and U6828 (N_6828,N_6739,N_6735);
nor U6829 (N_6829,N_6717,N_6706);
and U6830 (N_6830,N_6695,N_6530);
nand U6831 (N_6831,N_6727,N_6575);
and U6832 (N_6832,N_6563,N_6712);
nand U6833 (N_6833,N_6703,N_6675);
or U6834 (N_6834,N_6599,N_6612);
and U6835 (N_6835,N_6593,N_6580);
nand U6836 (N_6836,N_6684,N_6529);
xnor U6837 (N_6837,N_6721,N_6668);
xor U6838 (N_6838,N_6664,N_6512);
nand U6839 (N_6839,N_6556,N_6614);
nand U6840 (N_6840,N_6592,N_6638);
nor U6841 (N_6841,N_6729,N_6747);
xor U6842 (N_6842,N_6607,N_6639);
or U6843 (N_6843,N_6702,N_6579);
or U6844 (N_6844,N_6690,N_6606);
and U6845 (N_6845,N_6709,N_6616);
and U6846 (N_6846,N_6647,N_6657);
or U6847 (N_6847,N_6500,N_6569);
nand U6848 (N_6848,N_6541,N_6520);
xnor U6849 (N_6849,N_6511,N_6526);
xnor U6850 (N_6850,N_6736,N_6653);
nor U6851 (N_6851,N_6562,N_6688);
nor U6852 (N_6852,N_6663,N_6686);
xor U6853 (N_6853,N_6650,N_6644);
and U6854 (N_6854,N_6600,N_6745);
nor U6855 (N_6855,N_6620,N_6631);
or U6856 (N_6856,N_6641,N_6618);
and U6857 (N_6857,N_6553,N_6670);
nor U6858 (N_6858,N_6533,N_6518);
or U6859 (N_6859,N_6625,N_6737);
and U6860 (N_6860,N_6636,N_6740);
or U6861 (N_6861,N_6509,N_6567);
nor U6862 (N_6862,N_6632,N_6642);
and U6863 (N_6863,N_6624,N_6504);
nand U6864 (N_6864,N_6577,N_6732);
nor U6865 (N_6865,N_6705,N_6582);
or U6866 (N_6866,N_6720,N_6660);
and U6867 (N_6867,N_6711,N_6646);
and U6868 (N_6868,N_6635,N_6719);
or U6869 (N_6869,N_6701,N_6594);
or U6870 (N_6870,N_6696,N_6615);
and U6871 (N_6871,N_6522,N_6550);
or U6872 (N_6872,N_6710,N_6514);
nand U6873 (N_6873,N_6692,N_6743);
and U6874 (N_6874,N_6734,N_6587);
nand U6875 (N_6875,N_6595,N_6608);
and U6876 (N_6876,N_6541,N_6608);
nor U6877 (N_6877,N_6645,N_6702);
nand U6878 (N_6878,N_6585,N_6742);
nand U6879 (N_6879,N_6705,N_6532);
nor U6880 (N_6880,N_6507,N_6525);
or U6881 (N_6881,N_6667,N_6584);
or U6882 (N_6882,N_6502,N_6524);
nand U6883 (N_6883,N_6603,N_6718);
nand U6884 (N_6884,N_6608,N_6656);
or U6885 (N_6885,N_6522,N_6505);
nand U6886 (N_6886,N_6684,N_6704);
or U6887 (N_6887,N_6684,N_6589);
nor U6888 (N_6888,N_6599,N_6647);
nand U6889 (N_6889,N_6602,N_6670);
and U6890 (N_6890,N_6542,N_6561);
nor U6891 (N_6891,N_6511,N_6624);
and U6892 (N_6892,N_6641,N_6545);
nand U6893 (N_6893,N_6612,N_6580);
and U6894 (N_6894,N_6539,N_6509);
nand U6895 (N_6895,N_6702,N_6666);
nor U6896 (N_6896,N_6683,N_6550);
nor U6897 (N_6897,N_6597,N_6533);
and U6898 (N_6898,N_6563,N_6717);
and U6899 (N_6899,N_6727,N_6723);
nand U6900 (N_6900,N_6633,N_6687);
nor U6901 (N_6901,N_6596,N_6523);
nor U6902 (N_6902,N_6744,N_6533);
or U6903 (N_6903,N_6551,N_6582);
or U6904 (N_6904,N_6739,N_6605);
nor U6905 (N_6905,N_6511,N_6684);
or U6906 (N_6906,N_6678,N_6718);
nand U6907 (N_6907,N_6510,N_6585);
nor U6908 (N_6908,N_6555,N_6606);
and U6909 (N_6909,N_6583,N_6564);
and U6910 (N_6910,N_6607,N_6709);
xnor U6911 (N_6911,N_6558,N_6655);
nor U6912 (N_6912,N_6515,N_6577);
and U6913 (N_6913,N_6637,N_6650);
nor U6914 (N_6914,N_6579,N_6629);
nand U6915 (N_6915,N_6631,N_6650);
nand U6916 (N_6916,N_6534,N_6650);
nor U6917 (N_6917,N_6718,N_6692);
nor U6918 (N_6918,N_6748,N_6566);
nand U6919 (N_6919,N_6746,N_6556);
or U6920 (N_6920,N_6617,N_6572);
xor U6921 (N_6921,N_6663,N_6635);
and U6922 (N_6922,N_6636,N_6724);
nor U6923 (N_6923,N_6694,N_6546);
and U6924 (N_6924,N_6658,N_6548);
and U6925 (N_6925,N_6559,N_6725);
and U6926 (N_6926,N_6508,N_6649);
nor U6927 (N_6927,N_6710,N_6622);
xnor U6928 (N_6928,N_6730,N_6545);
xnor U6929 (N_6929,N_6585,N_6507);
and U6930 (N_6930,N_6658,N_6603);
nor U6931 (N_6931,N_6583,N_6705);
and U6932 (N_6932,N_6716,N_6727);
nor U6933 (N_6933,N_6689,N_6603);
or U6934 (N_6934,N_6526,N_6635);
nand U6935 (N_6935,N_6664,N_6542);
or U6936 (N_6936,N_6706,N_6687);
and U6937 (N_6937,N_6665,N_6736);
nand U6938 (N_6938,N_6615,N_6682);
or U6939 (N_6939,N_6584,N_6511);
nor U6940 (N_6940,N_6555,N_6743);
nor U6941 (N_6941,N_6647,N_6574);
nor U6942 (N_6942,N_6687,N_6664);
nor U6943 (N_6943,N_6632,N_6652);
nor U6944 (N_6944,N_6728,N_6652);
nor U6945 (N_6945,N_6695,N_6668);
nand U6946 (N_6946,N_6573,N_6528);
nor U6947 (N_6947,N_6525,N_6638);
or U6948 (N_6948,N_6721,N_6506);
nor U6949 (N_6949,N_6595,N_6529);
nand U6950 (N_6950,N_6576,N_6653);
nor U6951 (N_6951,N_6605,N_6721);
nand U6952 (N_6952,N_6507,N_6677);
nor U6953 (N_6953,N_6645,N_6516);
or U6954 (N_6954,N_6695,N_6561);
or U6955 (N_6955,N_6562,N_6708);
and U6956 (N_6956,N_6635,N_6647);
nor U6957 (N_6957,N_6610,N_6692);
or U6958 (N_6958,N_6511,N_6569);
or U6959 (N_6959,N_6704,N_6623);
or U6960 (N_6960,N_6709,N_6706);
xor U6961 (N_6961,N_6651,N_6504);
nor U6962 (N_6962,N_6654,N_6666);
xor U6963 (N_6963,N_6616,N_6507);
and U6964 (N_6964,N_6547,N_6565);
xnor U6965 (N_6965,N_6728,N_6655);
or U6966 (N_6966,N_6601,N_6719);
or U6967 (N_6967,N_6677,N_6610);
nand U6968 (N_6968,N_6693,N_6698);
nor U6969 (N_6969,N_6637,N_6633);
xor U6970 (N_6970,N_6555,N_6711);
and U6971 (N_6971,N_6690,N_6666);
nor U6972 (N_6972,N_6650,N_6636);
nor U6973 (N_6973,N_6607,N_6525);
or U6974 (N_6974,N_6506,N_6596);
or U6975 (N_6975,N_6532,N_6589);
or U6976 (N_6976,N_6504,N_6502);
xor U6977 (N_6977,N_6521,N_6723);
and U6978 (N_6978,N_6699,N_6570);
and U6979 (N_6979,N_6530,N_6709);
nand U6980 (N_6980,N_6571,N_6661);
nor U6981 (N_6981,N_6577,N_6704);
nor U6982 (N_6982,N_6546,N_6590);
nor U6983 (N_6983,N_6686,N_6650);
or U6984 (N_6984,N_6644,N_6652);
xnor U6985 (N_6985,N_6523,N_6525);
nor U6986 (N_6986,N_6641,N_6605);
xor U6987 (N_6987,N_6712,N_6591);
nor U6988 (N_6988,N_6738,N_6695);
xor U6989 (N_6989,N_6612,N_6571);
nor U6990 (N_6990,N_6562,N_6722);
nand U6991 (N_6991,N_6735,N_6610);
xnor U6992 (N_6992,N_6646,N_6599);
and U6993 (N_6993,N_6686,N_6533);
and U6994 (N_6994,N_6720,N_6653);
xor U6995 (N_6995,N_6569,N_6549);
nand U6996 (N_6996,N_6545,N_6729);
nand U6997 (N_6997,N_6698,N_6602);
and U6998 (N_6998,N_6540,N_6642);
and U6999 (N_6999,N_6530,N_6572);
nor U7000 (N_7000,N_6760,N_6833);
nor U7001 (N_7001,N_6981,N_6912);
nand U7002 (N_7002,N_6944,N_6996);
or U7003 (N_7003,N_6942,N_6913);
nand U7004 (N_7004,N_6823,N_6804);
nand U7005 (N_7005,N_6754,N_6995);
nand U7006 (N_7006,N_6851,N_6794);
nor U7007 (N_7007,N_6819,N_6908);
and U7008 (N_7008,N_6963,N_6884);
nor U7009 (N_7009,N_6974,N_6796);
nor U7010 (N_7010,N_6892,N_6930);
or U7011 (N_7011,N_6795,N_6836);
or U7012 (N_7012,N_6898,N_6977);
nand U7013 (N_7013,N_6813,N_6776);
or U7014 (N_7014,N_6972,N_6949);
and U7015 (N_7015,N_6903,N_6784);
or U7016 (N_7016,N_6957,N_6755);
and U7017 (N_7017,N_6826,N_6992);
or U7018 (N_7018,N_6774,N_6879);
or U7019 (N_7019,N_6976,N_6937);
and U7020 (N_7020,N_6779,N_6855);
nor U7021 (N_7021,N_6853,N_6948);
nand U7022 (N_7022,N_6990,N_6874);
nand U7023 (N_7023,N_6939,N_6919);
and U7024 (N_7024,N_6759,N_6814);
and U7025 (N_7025,N_6964,N_6991);
and U7026 (N_7026,N_6928,N_6886);
or U7027 (N_7027,N_6809,N_6959);
or U7028 (N_7028,N_6778,N_6883);
or U7029 (N_7029,N_6858,N_6854);
nor U7030 (N_7030,N_6877,N_6800);
nand U7031 (N_7031,N_6914,N_6897);
nand U7032 (N_7032,N_6911,N_6832);
nand U7033 (N_7033,N_6811,N_6862);
nand U7034 (N_7034,N_6835,N_6988);
nand U7035 (N_7035,N_6772,N_6915);
nor U7036 (N_7036,N_6820,N_6786);
nand U7037 (N_7037,N_6994,N_6758);
or U7038 (N_7038,N_6844,N_6878);
nor U7039 (N_7039,N_6818,N_6801);
and U7040 (N_7040,N_6876,N_6916);
or U7041 (N_7041,N_6782,N_6805);
nand U7042 (N_7042,N_6770,N_6921);
and U7043 (N_7043,N_6783,N_6923);
or U7044 (N_7044,N_6831,N_6924);
and U7045 (N_7045,N_6768,N_6803);
or U7046 (N_7046,N_6899,N_6837);
nand U7047 (N_7047,N_6986,N_6927);
or U7048 (N_7048,N_6989,N_6943);
xnor U7049 (N_7049,N_6781,N_6817);
nor U7050 (N_7050,N_6840,N_6935);
nand U7051 (N_7051,N_6895,N_6864);
nor U7052 (N_7052,N_6936,N_6905);
nor U7053 (N_7053,N_6790,N_6773);
and U7054 (N_7054,N_6802,N_6792);
nor U7055 (N_7055,N_6910,N_6764);
or U7056 (N_7056,N_6769,N_6860);
nand U7057 (N_7057,N_6904,N_6845);
or U7058 (N_7058,N_6987,N_6843);
and U7059 (N_7059,N_6893,N_6785);
nand U7060 (N_7060,N_6940,N_6969);
xor U7061 (N_7061,N_6932,N_6982);
or U7062 (N_7062,N_6975,N_6979);
or U7063 (N_7063,N_6907,N_6882);
or U7064 (N_7064,N_6920,N_6955);
and U7065 (N_7065,N_6791,N_6967);
nand U7066 (N_7066,N_6896,N_6894);
nand U7067 (N_7067,N_6841,N_6946);
nand U7068 (N_7068,N_6767,N_6880);
xor U7069 (N_7069,N_6887,N_6797);
nand U7070 (N_7070,N_6889,N_6900);
or U7071 (N_7071,N_6978,N_6868);
and U7072 (N_7072,N_6909,N_6829);
nor U7073 (N_7073,N_6875,N_6947);
xor U7074 (N_7074,N_6771,N_6857);
or U7075 (N_7075,N_6765,N_6961);
nand U7076 (N_7076,N_6827,N_6922);
and U7077 (N_7077,N_6917,N_6952);
nand U7078 (N_7078,N_6980,N_6762);
xor U7079 (N_7079,N_6834,N_6869);
or U7080 (N_7080,N_6787,N_6867);
xor U7081 (N_7081,N_6956,N_6888);
nor U7082 (N_7082,N_6863,N_6881);
nand U7083 (N_7083,N_6958,N_6777);
nand U7084 (N_7084,N_6852,N_6788);
nand U7085 (N_7085,N_6850,N_6918);
xnor U7086 (N_7086,N_6873,N_6752);
nand U7087 (N_7087,N_6871,N_6756);
nand U7088 (N_7088,N_6842,N_6971);
or U7089 (N_7089,N_6859,N_6954);
nand U7090 (N_7090,N_6866,N_6934);
nand U7091 (N_7091,N_6780,N_6941);
nor U7092 (N_7092,N_6966,N_6806);
xnor U7093 (N_7093,N_6938,N_6789);
or U7094 (N_7094,N_6865,N_6973);
nor U7095 (N_7095,N_6951,N_6950);
xnor U7096 (N_7096,N_6847,N_6825);
nor U7097 (N_7097,N_6838,N_6931);
nand U7098 (N_7098,N_6998,N_6984);
and U7099 (N_7099,N_6906,N_6968);
and U7100 (N_7100,N_6807,N_6815);
nand U7101 (N_7101,N_6985,N_6751);
nand U7102 (N_7102,N_6810,N_6999);
and U7103 (N_7103,N_6945,N_6799);
xnor U7104 (N_7104,N_6953,N_6824);
and U7105 (N_7105,N_6808,N_6793);
nor U7106 (N_7106,N_6856,N_6816);
nand U7107 (N_7107,N_6970,N_6872);
xor U7108 (N_7108,N_6828,N_6870);
nand U7109 (N_7109,N_6925,N_6926);
xor U7110 (N_7110,N_6885,N_6902);
and U7111 (N_7111,N_6753,N_6812);
xor U7112 (N_7112,N_6822,N_6962);
nand U7113 (N_7113,N_6890,N_6750);
and U7114 (N_7114,N_6775,N_6761);
nor U7115 (N_7115,N_6821,N_6763);
or U7116 (N_7116,N_6798,N_6929);
and U7117 (N_7117,N_6849,N_6848);
xor U7118 (N_7118,N_6839,N_6901);
nand U7119 (N_7119,N_6993,N_6846);
nor U7120 (N_7120,N_6983,N_6965);
nand U7121 (N_7121,N_6766,N_6830);
nand U7122 (N_7122,N_6891,N_6960);
nor U7123 (N_7123,N_6997,N_6933);
nand U7124 (N_7124,N_6757,N_6861);
nor U7125 (N_7125,N_6912,N_6892);
or U7126 (N_7126,N_6866,N_6993);
nor U7127 (N_7127,N_6831,N_6952);
nor U7128 (N_7128,N_6983,N_6802);
xnor U7129 (N_7129,N_6761,N_6931);
nand U7130 (N_7130,N_6924,N_6929);
xor U7131 (N_7131,N_6864,N_6828);
and U7132 (N_7132,N_6769,N_6829);
xnor U7133 (N_7133,N_6765,N_6885);
nor U7134 (N_7134,N_6839,N_6775);
nand U7135 (N_7135,N_6767,N_6985);
nand U7136 (N_7136,N_6905,N_6982);
nand U7137 (N_7137,N_6877,N_6894);
nand U7138 (N_7138,N_6881,N_6899);
nand U7139 (N_7139,N_6819,N_6831);
nand U7140 (N_7140,N_6880,N_6799);
or U7141 (N_7141,N_6925,N_6833);
and U7142 (N_7142,N_6908,N_6778);
or U7143 (N_7143,N_6839,N_6885);
xor U7144 (N_7144,N_6845,N_6873);
nor U7145 (N_7145,N_6941,N_6821);
or U7146 (N_7146,N_6860,N_6886);
nor U7147 (N_7147,N_6789,N_6835);
nand U7148 (N_7148,N_6757,N_6811);
and U7149 (N_7149,N_6916,N_6773);
nor U7150 (N_7150,N_6921,N_6842);
or U7151 (N_7151,N_6767,N_6996);
nor U7152 (N_7152,N_6862,N_6773);
nor U7153 (N_7153,N_6851,N_6843);
nor U7154 (N_7154,N_6780,N_6861);
or U7155 (N_7155,N_6887,N_6809);
nand U7156 (N_7156,N_6782,N_6845);
nand U7157 (N_7157,N_6774,N_6767);
xnor U7158 (N_7158,N_6755,N_6971);
or U7159 (N_7159,N_6903,N_6972);
nand U7160 (N_7160,N_6790,N_6891);
or U7161 (N_7161,N_6890,N_6922);
or U7162 (N_7162,N_6990,N_6802);
and U7163 (N_7163,N_6899,N_6796);
nor U7164 (N_7164,N_6915,N_6753);
nand U7165 (N_7165,N_6833,N_6851);
nor U7166 (N_7166,N_6954,N_6780);
nand U7167 (N_7167,N_6996,N_6751);
and U7168 (N_7168,N_6966,N_6849);
nor U7169 (N_7169,N_6807,N_6774);
and U7170 (N_7170,N_6972,N_6881);
or U7171 (N_7171,N_6821,N_6987);
nand U7172 (N_7172,N_6847,N_6790);
nor U7173 (N_7173,N_6859,N_6801);
nor U7174 (N_7174,N_6964,N_6843);
and U7175 (N_7175,N_6930,N_6970);
nor U7176 (N_7176,N_6825,N_6793);
or U7177 (N_7177,N_6926,N_6836);
or U7178 (N_7178,N_6914,N_6899);
or U7179 (N_7179,N_6833,N_6864);
and U7180 (N_7180,N_6974,N_6817);
nand U7181 (N_7181,N_6960,N_6941);
and U7182 (N_7182,N_6974,N_6908);
nor U7183 (N_7183,N_6855,N_6762);
nor U7184 (N_7184,N_6804,N_6788);
nor U7185 (N_7185,N_6942,N_6902);
or U7186 (N_7186,N_6974,N_6978);
nor U7187 (N_7187,N_6844,N_6876);
and U7188 (N_7188,N_6957,N_6807);
or U7189 (N_7189,N_6916,N_6923);
xnor U7190 (N_7190,N_6971,N_6787);
and U7191 (N_7191,N_6911,N_6995);
or U7192 (N_7192,N_6986,N_6962);
or U7193 (N_7193,N_6951,N_6815);
or U7194 (N_7194,N_6997,N_6801);
nor U7195 (N_7195,N_6828,N_6987);
nand U7196 (N_7196,N_6802,N_6957);
nor U7197 (N_7197,N_6840,N_6777);
xor U7198 (N_7198,N_6791,N_6814);
nand U7199 (N_7199,N_6767,N_6998);
nand U7200 (N_7200,N_6821,N_6925);
nand U7201 (N_7201,N_6854,N_6860);
and U7202 (N_7202,N_6984,N_6764);
and U7203 (N_7203,N_6924,N_6766);
nand U7204 (N_7204,N_6759,N_6950);
nor U7205 (N_7205,N_6953,N_6994);
nand U7206 (N_7206,N_6968,N_6957);
nand U7207 (N_7207,N_6958,N_6841);
or U7208 (N_7208,N_6925,N_6921);
nor U7209 (N_7209,N_6987,N_6950);
nor U7210 (N_7210,N_6812,N_6954);
or U7211 (N_7211,N_6857,N_6788);
nor U7212 (N_7212,N_6884,N_6928);
or U7213 (N_7213,N_6799,N_6946);
nand U7214 (N_7214,N_6877,N_6757);
xor U7215 (N_7215,N_6894,N_6850);
xnor U7216 (N_7216,N_6919,N_6915);
nor U7217 (N_7217,N_6775,N_6923);
nand U7218 (N_7218,N_6932,N_6759);
nor U7219 (N_7219,N_6963,N_6799);
and U7220 (N_7220,N_6918,N_6944);
nand U7221 (N_7221,N_6991,N_6916);
xnor U7222 (N_7222,N_6981,N_6868);
nand U7223 (N_7223,N_6817,N_6970);
nand U7224 (N_7224,N_6948,N_6802);
nor U7225 (N_7225,N_6980,N_6848);
nand U7226 (N_7226,N_6864,N_6974);
nand U7227 (N_7227,N_6980,N_6973);
nand U7228 (N_7228,N_6881,N_6838);
or U7229 (N_7229,N_6990,N_6757);
xor U7230 (N_7230,N_6873,N_6773);
and U7231 (N_7231,N_6838,N_6801);
nand U7232 (N_7232,N_6972,N_6940);
nand U7233 (N_7233,N_6936,N_6842);
xnor U7234 (N_7234,N_6899,N_6811);
nor U7235 (N_7235,N_6877,N_6770);
nor U7236 (N_7236,N_6975,N_6985);
nand U7237 (N_7237,N_6769,N_6777);
nor U7238 (N_7238,N_6805,N_6982);
or U7239 (N_7239,N_6947,N_6996);
nor U7240 (N_7240,N_6956,N_6755);
and U7241 (N_7241,N_6800,N_6882);
and U7242 (N_7242,N_6947,N_6894);
or U7243 (N_7243,N_6781,N_6819);
nand U7244 (N_7244,N_6988,N_6883);
nor U7245 (N_7245,N_6840,N_6870);
or U7246 (N_7246,N_6915,N_6888);
and U7247 (N_7247,N_6934,N_6754);
nand U7248 (N_7248,N_6934,N_6823);
and U7249 (N_7249,N_6827,N_6876);
or U7250 (N_7250,N_7121,N_7127);
and U7251 (N_7251,N_7122,N_7247);
nor U7252 (N_7252,N_7153,N_7069);
nand U7253 (N_7253,N_7146,N_7043);
and U7254 (N_7254,N_7210,N_7107);
or U7255 (N_7255,N_7054,N_7185);
nand U7256 (N_7256,N_7162,N_7033);
xnor U7257 (N_7257,N_7198,N_7021);
nand U7258 (N_7258,N_7228,N_7155);
nor U7259 (N_7259,N_7201,N_7110);
or U7260 (N_7260,N_7194,N_7204);
and U7261 (N_7261,N_7189,N_7163);
or U7262 (N_7262,N_7231,N_7184);
xnor U7263 (N_7263,N_7216,N_7106);
or U7264 (N_7264,N_7142,N_7148);
nor U7265 (N_7265,N_7093,N_7056);
xor U7266 (N_7266,N_7232,N_7109);
nor U7267 (N_7267,N_7028,N_7085);
and U7268 (N_7268,N_7213,N_7044);
xor U7269 (N_7269,N_7188,N_7175);
or U7270 (N_7270,N_7136,N_7246);
nand U7271 (N_7271,N_7117,N_7138);
nor U7272 (N_7272,N_7015,N_7080);
or U7273 (N_7273,N_7062,N_7099);
or U7274 (N_7274,N_7087,N_7186);
or U7275 (N_7275,N_7012,N_7149);
and U7276 (N_7276,N_7089,N_7004);
nor U7277 (N_7277,N_7063,N_7249);
nor U7278 (N_7278,N_7157,N_7225);
and U7279 (N_7279,N_7208,N_7196);
and U7280 (N_7280,N_7123,N_7164);
and U7281 (N_7281,N_7035,N_7061);
nor U7282 (N_7282,N_7088,N_7202);
or U7283 (N_7283,N_7240,N_7038);
or U7284 (N_7284,N_7078,N_7008);
and U7285 (N_7285,N_7179,N_7167);
nand U7286 (N_7286,N_7158,N_7124);
xor U7287 (N_7287,N_7095,N_7177);
nor U7288 (N_7288,N_7100,N_7129);
and U7289 (N_7289,N_7126,N_7145);
or U7290 (N_7290,N_7092,N_7226);
xnor U7291 (N_7291,N_7079,N_7005);
nand U7292 (N_7292,N_7140,N_7016);
and U7293 (N_7293,N_7013,N_7019);
or U7294 (N_7294,N_7108,N_7031);
xor U7295 (N_7295,N_7200,N_7191);
nor U7296 (N_7296,N_7036,N_7034);
xor U7297 (N_7297,N_7101,N_7139);
or U7298 (N_7298,N_7055,N_7152);
and U7299 (N_7299,N_7030,N_7025);
or U7300 (N_7300,N_7193,N_7075);
nor U7301 (N_7301,N_7159,N_7022);
nand U7302 (N_7302,N_7026,N_7071);
and U7303 (N_7303,N_7183,N_7230);
and U7304 (N_7304,N_7072,N_7245);
or U7305 (N_7305,N_7074,N_7002);
xor U7306 (N_7306,N_7141,N_7220);
and U7307 (N_7307,N_7115,N_7132);
or U7308 (N_7308,N_7073,N_7187);
and U7309 (N_7309,N_7144,N_7170);
nand U7310 (N_7310,N_7130,N_7120);
and U7311 (N_7311,N_7046,N_7192);
nand U7312 (N_7312,N_7243,N_7116);
nor U7313 (N_7313,N_7211,N_7176);
and U7314 (N_7314,N_7090,N_7011);
and U7315 (N_7315,N_7212,N_7098);
nor U7316 (N_7316,N_7190,N_7165);
or U7317 (N_7317,N_7241,N_7009);
nor U7318 (N_7318,N_7135,N_7239);
nand U7319 (N_7319,N_7023,N_7242);
nand U7320 (N_7320,N_7218,N_7222);
and U7321 (N_7321,N_7058,N_7219);
nand U7322 (N_7322,N_7045,N_7007);
nor U7323 (N_7323,N_7244,N_7137);
nor U7324 (N_7324,N_7097,N_7224);
nor U7325 (N_7325,N_7040,N_7248);
and U7326 (N_7326,N_7174,N_7166);
nor U7327 (N_7327,N_7229,N_7018);
or U7328 (N_7328,N_7215,N_7143);
and U7329 (N_7329,N_7182,N_7236);
and U7330 (N_7330,N_7048,N_7037);
nor U7331 (N_7331,N_7205,N_7029);
or U7332 (N_7332,N_7066,N_7003);
and U7333 (N_7333,N_7150,N_7214);
nor U7334 (N_7334,N_7027,N_7209);
or U7335 (N_7335,N_7151,N_7169);
and U7336 (N_7336,N_7105,N_7227);
nor U7337 (N_7337,N_7047,N_7119);
or U7338 (N_7338,N_7094,N_7081);
nor U7339 (N_7339,N_7118,N_7104);
or U7340 (N_7340,N_7207,N_7147);
or U7341 (N_7341,N_7237,N_7076);
and U7342 (N_7342,N_7235,N_7180);
and U7343 (N_7343,N_7133,N_7065);
or U7344 (N_7344,N_7051,N_7134);
and U7345 (N_7345,N_7161,N_7064);
and U7346 (N_7346,N_7096,N_7041);
nor U7347 (N_7347,N_7050,N_7203);
nor U7348 (N_7348,N_7173,N_7156);
nor U7349 (N_7349,N_7086,N_7032);
and U7350 (N_7350,N_7057,N_7060);
nor U7351 (N_7351,N_7111,N_7112);
and U7352 (N_7352,N_7217,N_7131);
nor U7353 (N_7353,N_7125,N_7067);
and U7354 (N_7354,N_7042,N_7223);
nor U7355 (N_7355,N_7020,N_7197);
and U7356 (N_7356,N_7001,N_7181);
nand U7357 (N_7357,N_7059,N_7221);
nand U7358 (N_7358,N_7154,N_7000);
and U7359 (N_7359,N_7128,N_7178);
nor U7360 (N_7360,N_7091,N_7206);
or U7361 (N_7361,N_7171,N_7113);
xor U7362 (N_7362,N_7070,N_7172);
nor U7363 (N_7363,N_7052,N_7082);
nor U7364 (N_7364,N_7068,N_7010);
and U7365 (N_7365,N_7006,N_7053);
nand U7366 (N_7366,N_7234,N_7168);
and U7367 (N_7367,N_7083,N_7017);
nand U7368 (N_7368,N_7077,N_7084);
nor U7369 (N_7369,N_7114,N_7102);
or U7370 (N_7370,N_7049,N_7014);
and U7371 (N_7371,N_7233,N_7024);
or U7372 (N_7372,N_7103,N_7160);
or U7373 (N_7373,N_7238,N_7195);
or U7374 (N_7374,N_7199,N_7039);
or U7375 (N_7375,N_7194,N_7245);
nor U7376 (N_7376,N_7080,N_7132);
nand U7377 (N_7377,N_7037,N_7230);
nand U7378 (N_7378,N_7002,N_7182);
or U7379 (N_7379,N_7031,N_7016);
and U7380 (N_7380,N_7004,N_7056);
or U7381 (N_7381,N_7181,N_7007);
and U7382 (N_7382,N_7053,N_7214);
nor U7383 (N_7383,N_7148,N_7242);
or U7384 (N_7384,N_7050,N_7169);
nand U7385 (N_7385,N_7165,N_7052);
and U7386 (N_7386,N_7206,N_7010);
nor U7387 (N_7387,N_7111,N_7048);
nor U7388 (N_7388,N_7069,N_7080);
or U7389 (N_7389,N_7240,N_7148);
or U7390 (N_7390,N_7004,N_7005);
xor U7391 (N_7391,N_7093,N_7190);
and U7392 (N_7392,N_7213,N_7241);
nand U7393 (N_7393,N_7018,N_7162);
or U7394 (N_7394,N_7146,N_7114);
nand U7395 (N_7395,N_7049,N_7057);
nor U7396 (N_7396,N_7137,N_7172);
nor U7397 (N_7397,N_7114,N_7068);
nor U7398 (N_7398,N_7236,N_7231);
nand U7399 (N_7399,N_7025,N_7165);
or U7400 (N_7400,N_7221,N_7218);
nand U7401 (N_7401,N_7123,N_7097);
and U7402 (N_7402,N_7039,N_7108);
or U7403 (N_7403,N_7141,N_7097);
xnor U7404 (N_7404,N_7115,N_7107);
or U7405 (N_7405,N_7025,N_7135);
and U7406 (N_7406,N_7013,N_7008);
and U7407 (N_7407,N_7224,N_7103);
or U7408 (N_7408,N_7061,N_7199);
nand U7409 (N_7409,N_7144,N_7048);
nor U7410 (N_7410,N_7065,N_7195);
xnor U7411 (N_7411,N_7170,N_7240);
nand U7412 (N_7412,N_7140,N_7097);
nand U7413 (N_7413,N_7156,N_7123);
nor U7414 (N_7414,N_7124,N_7090);
xor U7415 (N_7415,N_7195,N_7077);
and U7416 (N_7416,N_7195,N_7040);
nor U7417 (N_7417,N_7017,N_7146);
nand U7418 (N_7418,N_7096,N_7036);
nor U7419 (N_7419,N_7159,N_7029);
nand U7420 (N_7420,N_7164,N_7150);
and U7421 (N_7421,N_7129,N_7000);
or U7422 (N_7422,N_7061,N_7106);
nor U7423 (N_7423,N_7005,N_7225);
nor U7424 (N_7424,N_7195,N_7172);
or U7425 (N_7425,N_7213,N_7134);
and U7426 (N_7426,N_7105,N_7072);
nor U7427 (N_7427,N_7171,N_7045);
or U7428 (N_7428,N_7159,N_7180);
nor U7429 (N_7429,N_7027,N_7173);
nor U7430 (N_7430,N_7133,N_7189);
nor U7431 (N_7431,N_7231,N_7160);
or U7432 (N_7432,N_7237,N_7055);
nand U7433 (N_7433,N_7131,N_7138);
nand U7434 (N_7434,N_7227,N_7186);
nand U7435 (N_7435,N_7200,N_7177);
and U7436 (N_7436,N_7193,N_7114);
or U7437 (N_7437,N_7138,N_7042);
and U7438 (N_7438,N_7162,N_7234);
nor U7439 (N_7439,N_7122,N_7213);
xnor U7440 (N_7440,N_7235,N_7199);
and U7441 (N_7441,N_7013,N_7109);
and U7442 (N_7442,N_7163,N_7110);
nor U7443 (N_7443,N_7003,N_7074);
or U7444 (N_7444,N_7240,N_7154);
or U7445 (N_7445,N_7214,N_7088);
nand U7446 (N_7446,N_7195,N_7088);
and U7447 (N_7447,N_7016,N_7060);
nand U7448 (N_7448,N_7220,N_7138);
nand U7449 (N_7449,N_7228,N_7139);
xnor U7450 (N_7450,N_7059,N_7186);
nand U7451 (N_7451,N_7158,N_7034);
nand U7452 (N_7452,N_7118,N_7019);
nand U7453 (N_7453,N_7122,N_7161);
xnor U7454 (N_7454,N_7037,N_7184);
or U7455 (N_7455,N_7203,N_7037);
nand U7456 (N_7456,N_7146,N_7095);
xnor U7457 (N_7457,N_7169,N_7000);
and U7458 (N_7458,N_7145,N_7024);
and U7459 (N_7459,N_7212,N_7244);
xor U7460 (N_7460,N_7231,N_7176);
and U7461 (N_7461,N_7221,N_7210);
or U7462 (N_7462,N_7169,N_7121);
nor U7463 (N_7463,N_7107,N_7041);
nand U7464 (N_7464,N_7036,N_7094);
nor U7465 (N_7465,N_7113,N_7105);
and U7466 (N_7466,N_7238,N_7151);
nand U7467 (N_7467,N_7046,N_7215);
and U7468 (N_7468,N_7050,N_7047);
xnor U7469 (N_7469,N_7215,N_7091);
or U7470 (N_7470,N_7101,N_7041);
nor U7471 (N_7471,N_7056,N_7196);
or U7472 (N_7472,N_7244,N_7124);
and U7473 (N_7473,N_7139,N_7102);
or U7474 (N_7474,N_7136,N_7111);
and U7475 (N_7475,N_7037,N_7136);
nand U7476 (N_7476,N_7117,N_7108);
nand U7477 (N_7477,N_7200,N_7163);
or U7478 (N_7478,N_7237,N_7222);
and U7479 (N_7479,N_7006,N_7114);
nand U7480 (N_7480,N_7079,N_7235);
or U7481 (N_7481,N_7248,N_7073);
nor U7482 (N_7482,N_7117,N_7097);
nor U7483 (N_7483,N_7173,N_7154);
and U7484 (N_7484,N_7160,N_7038);
and U7485 (N_7485,N_7182,N_7007);
nand U7486 (N_7486,N_7230,N_7180);
or U7487 (N_7487,N_7233,N_7244);
and U7488 (N_7488,N_7041,N_7156);
nor U7489 (N_7489,N_7076,N_7052);
nand U7490 (N_7490,N_7242,N_7008);
and U7491 (N_7491,N_7172,N_7136);
and U7492 (N_7492,N_7195,N_7203);
nand U7493 (N_7493,N_7092,N_7210);
nand U7494 (N_7494,N_7167,N_7096);
or U7495 (N_7495,N_7239,N_7103);
and U7496 (N_7496,N_7190,N_7216);
and U7497 (N_7497,N_7092,N_7236);
nor U7498 (N_7498,N_7038,N_7084);
nor U7499 (N_7499,N_7192,N_7244);
or U7500 (N_7500,N_7367,N_7318);
nand U7501 (N_7501,N_7440,N_7323);
nand U7502 (N_7502,N_7411,N_7392);
nand U7503 (N_7503,N_7355,N_7405);
nand U7504 (N_7504,N_7291,N_7398);
nand U7505 (N_7505,N_7287,N_7264);
and U7506 (N_7506,N_7369,N_7317);
and U7507 (N_7507,N_7455,N_7370);
nor U7508 (N_7508,N_7390,N_7424);
nand U7509 (N_7509,N_7302,N_7478);
nor U7510 (N_7510,N_7319,N_7456);
xnor U7511 (N_7511,N_7400,N_7431);
and U7512 (N_7512,N_7450,N_7298);
nor U7513 (N_7513,N_7338,N_7251);
or U7514 (N_7514,N_7384,N_7352);
and U7515 (N_7515,N_7458,N_7362);
and U7516 (N_7516,N_7290,N_7259);
nor U7517 (N_7517,N_7375,N_7328);
xor U7518 (N_7518,N_7413,N_7437);
or U7519 (N_7519,N_7383,N_7409);
nand U7520 (N_7520,N_7356,N_7320);
or U7521 (N_7521,N_7479,N_7301);
or U7522 (N_7522,N_7434,N_7447);
nor U7523 (N_7523,N_7368,N_7307);
or U7524 (N_7524,N_7308,N_7486);
or U7525 (N_7525,N_7295,N_7410);
or U7526 (N_7526,N_7316,N_7267);
and U7527 (N_7527,N_7359,N_7294);
or U7528 (N_7528,N_7348,N_7252);
or U7529 (N_7529,N_7467,N_7423);
nor U7530 (N_7530,N_7349,N_7436);
nor U7531 (N_7531,N_7379,N_7474);
and U7532 (N_7532,N_7339,N_7380);
nor U7533 (N_7533,N_7443,N_7363);
nand U7534 (N_7534,N_7448,N_7310);
nor U7535 (N_7535,N_7300,N_7357);
and U7536 (N_7536,N_7293,N_7490);
and U7537 (N_7537,N_7334,N_7417);
or U7538 (N_7538,N_7358,N_7376);
xnor U7539 (N_7539,N_7461,N_7336);
and U7540 (N_7540,N_7432,N_7489);
and U7541 (N_7541,N_7261,N_7445);
nor U7542 (N_7542,N_7484,N_7406);
xnor U7543 (N_7543,N_7466,N_7414);
xor U7544 (N_7544,N_7347,N_7321);
nand U7545 (N_7545,N_7374,N_7385);
and U7546 (N_7546,N_7340,N_7396);
and U7547 (N_7547,N_7271,N_7332);
and U7548 (N_7548,N_7262,N_7421);
nor U7549 (N_7549,N_7491,N_7419);
nor U7550 (N_7550,N_7258,N_7361);
nor U7551 (N_7551,N_7255,N_7331);
nor U7552 (N_7552,N_7329,N_7283);
or U7553 (N_7553,N_7274,N_7281);
xor U7554 (N_7554,N_7488,N_7464);
xor U7555 (N_7555,N_7366,N_7454);
and U7556 (N_7556,N_7364,N_7256);
nand U7557 (N_7557,N_7312,N_7265);
nor U7558 (N_7558,N_7471,N_7402);
nor U7559 (N_7559,N_7460,N_7343);
nand U7560 (N_7560,N_7278,N_7275);
nor U7561 (N_7561,N_7354,N_7285);
xnor U7562 (N_7562,N_7430,N_7288);
and U7563 (N_7563,N_7482,N_7304);
nand U7564 (N_7564,N_7395,N_7418);
nand U7565 (N_7565,N_7389,N_7483);
or U7566 (N_7566,N_7260,N_7372);
xnor U7567 (N_7567,N_7407,N_7403);
nor U7568 (N_7568,N_7333,N_7435);
or U7569 (N_7569,N_7327,N_7477);
or U7570 (N_7570,N_7404,N_7266);
nor U7571 (N_7571,N_7254,N_7401);
nand U7572 (N_7572,N_7344,N_7444);
or U7573 (N_7573,N_7463,N_7387);
and U7574 (N_7574,N_7276,N_7351);
and U7575 (N_7575,N_7468,N_7373);
nor U7576 (N_7576,N_7330,N_7426);
or U7577 (N_7577,N_7438,N_7498);
and U7578 (N_7578,N_7439,N_7470);
nor U7579 (N_7579,N_7277,N_7415);
or U7580 (N_7580,N_7420,N_7469);
nor U7581 (N_7581,N_7280,N_7350);
nor U7582 (N_7582,N_7270,N_7388);
and U7583 (N_7583,N_7397,N_7416);
nor U7584 (N_7584,N_7353,N_7263);
and U7585 (N_7585,N_7465,N_7472);
and U7586 (N_7586,N_7282,N_7313);
nand U7587 (N_7587,N_7272,N_7335);
nor U7588 (N_7588,N_7441,N_7314);
and U7589 (N_7589,N_7322,N_7299);
or U7590 (N_7590,N_7306,N_7378);
nor U7591 (N_7591,N_7428,N_7408);
or U7592 (N_7592,N_7365,N_7433);
nand U7593 (N_7593,N_7371,N_7481);
or U7594 (N_7594,N_7485,N_7442);
nor U7595 (N_7595,N_7315,N_7412);
xnor U7596 (N_7596,N_7494,N_7475);
or U7597 (N_7597,N_7279,N_7446);
nor U7598 (N_7598,N_7382,N_7493);
nor U7599 (N_7599,N_7296,N_7268);
nor U7600 (N_7600,N_7393,N_7451);
and U7601 (N_7601,N_7346,N_7326);
and U7602 (N_7602,N_7425,N_7253);
and U7603 (N_7603,N_7324,N_7286);
and U7604 (N_7604,N_7462,N_7297);
nor U7605 (N_7605,N_7309,N_7305);
nand U7606 (N_7606,N_7257,N_7399);
and U7607 (N_7607,N_7311,N_7386);
or U7608 (N_7608,N_7492,N_7452);
and U7609 (N_7609,N_7495,N_7427);
nand U7610 (N_7610,N_7480,N_7497);
and U7611 (N_7611,N_7269,N_7457);
or U7612 (N_7612,N_7325,N_7342);
and U7613 (N_7613,N_7487,N_7292);
nand U7614 (N_7614,N_7476,N_7422);
or U7615 (N_7615,N_7496,N_7337);
nor U7616 (N_7616,N_7453,N_7429);
or U7617 (N_7617,N_7381,N_7360);
and U7618 (N_7618,N_7303,N_7289);
and U7619 (N_7619,N_7377,N_7449);
or U7620 (N_7620,N_7459,N_7391);
nor U7621 (N_7621,N_7273,N_7394);
or U7622 (N_7622,N_7345,N_7499);
xor U7623 (N_7623,N_7250,N_7284);
or U7624 (N_7624,N_7473,N_7341);
and U7625 (N_7625,N_7277,N_7398);
and U7626 (N_7626,N_7333,N_7281);
nor U7627 (N_7627,N_7331,N_7292);
nand U7628 (N_7628,N_7279,N_7367);
xor U7629 (N_7629,N_7492,N_7299);
and U7630 (N_7630,N_7348,N_7459);
or U7631 (N_7631,N_7433,N_7291);
or U7632 (N_7632,N_7311,N_7447);
and U7633 (N_7633,N_7442,N_7492);
and U7634 (N_7634,N_7490,N_7302);
and U7635 (N_7635,N_7287,N_7495);
nor U7636 (N_7636,N_7462,N_7374);
and U7637 (N_7637,N_7410,N_7286);
or U7638 (N_7638,N_7363,N_7331);
nand U7639 (N_7639,N_7358,N_7372);
and U7640 (N_7640,N_7366,N_7461);
nor U7641 (N_7641,N_7283,N_7311);
and U7642 (N_7642,N_7327,N_7318);
nand U7643 (N_7643,N_7419,N_7353);
or U7644 (N_7644,N_7490,N_7489);
nand U7645 (N_7645,N_7304,N_7299);
nand U7646 (N_7646,N_7369,N_7485);
nand U7647 (N_7647,N_7428,N_7309);
nand U7648 (N_7648,N_7455,N_7486);
or U7649 (N_7649,N_7251,N_7455);
nand U7650 (N_7650,N_7406,N_7326);
nor U7651 (N_7651,N_7492,N_7450);
nor U7652 (N_7652,N_7485,N_7359);
or U7653 (N_7653,N_7476,N_7365);
nand U7654 (N_7654,N_7343,N_7326);
nor U7655 (N_7655,N_7499,N_7413);
and U7656 (N_7656,N_7298,N_7406);
nand U7657 (N_7657,N_7430,N_7387);
nand U7658 (N_7658,N_7271,N_7280);
or U7659 (N_7659,N_7253,N_7307);
or U7660 (N_7660,N_7479,N_7260);
or U7661 (N_7661,N_7391,N_7290);
xor U7662 (N_7662,N_7457,N_7353);
xnor U7663 (N_7663,N_7253,N_7340);
and U7664 (N_7664,N_7361,N_7492);
xnor U7665 (N_7665,N_7258,N_7362);
nor U7666 (N_7666,N_7360,N_7358);
and U7667 (N_7667,N_7269,N_7268);
or U7668 (N_7668,N_7326,N_7294);
nor U7669 (N_7669,N_7260,N_7388);
nand U7670 (N_7670,N_7418,N_7391);
and U7671 (N_7671,N_7404,N_7333);
nor U7672 (N_7672,N_7490,N_7423);
or U7673 (N_7673,N_7323,N_7448);
or U7674 (N_7674,N_7274,N_7331);
nand U7675 (N_7675,N_7414,N_7385);
xor U7676 (N_7676,N_7324,N_7451);
or U7677 (N_7677,N_7488,N_7484);
and U7678 (N_7678,N_7326,N_7447);
or U7679 (N_7679,N_7343,N_7463);
nor U7680 (N_7680,N_7372,N_7489);
xor U7681 (N_7681,N_7330,N_7403);
or U7682 (N_7682,N_7331,N_7451);
nand U7683 (N_7683,N_7277,N_7433);
and U7684 (N_7684,N_7491,N_7321);
nand U7685 (N_7685,N_7431,N_7303);
nand U7686 (N_7686,N_7492,N_7317);
nor U7687 (N_7687,N_7371,N_7292);
nand U7688 (N_7688,N_7388,N_7486);
and U7689 (N_7689,N_7294,N_7348);
nand U7690 (N_7690,N_7440,N_7331);
nand U7691 (N_7691,N_7288,N_7378);
and U7692 (N_7692,N_7254,N_7434);
nor U7693 (N_7693,N_7326,N_7254);
nor U7694 (N_7694,N_7301,N_7379);
nor U7695 (N_7695,N_7324,N_7275);
or U7696 (N_7696,N_7437,N_7340);
or U7697 (N_7697,N_7497,N_7368);
nand U7698 (N_7698,N_7339,N_7424);
xnor U7699 (N_7699,N_7394,N_7386);
nand U7700 (N_7700,N_7396,N_7261);
or U7701 (N_7701,N_7450,N_7306);
nor U7702 (N_7702,N_7292,N_7339);
and U7703 (N_7703,N_7435,N_7481);
nor U7704 (N_7704,N_7361,N_7311);
and U7705 (N_7705,N_7409,N_7493);
and U7706 (N_7706,N_7289,N_7333);
nor U7707 (N_7707,N_7472,N_7382);
nor U7708 (N_7708,N_7453,N_7487);
and U7709 (N_7709,N_7333,N_7464);
nand U7710 (N_7710,N_7440,N_7264);
nor U7711 (N_7711,N_7431,N_7386);
or U7712 (N_7712,N_7320,N_7313);
nor U7713 (N_7713,N_7376,N_7317);
nor U7714 (N_7714,N_7330,N_7274);
nand U7715 (N_7715,N_7494,N_7420);
nor U7716 (N_7716,N_7352,N_7457);
nand U7717 (N_7717,N_7328,N_7393);
nand U7718 (N_7718,N_7456,N_7372);
nor U7719 (N_7719,N_7484,N_7380);
nor U7720 (N_7720,N_7472,N_7257);
xor U7721 (N_7721,N_7253,N_7282);
nor U7722 (N_7722,N_7316,N_7320);
nor U7723 (N_7723,N_7272,N_7440);
nand U7724 (N_7724,N_7252,N_7370);
nand U7725 (N_7725,N_7405,N_7270);
or U7726 (N_7726,N_7336,N_7309);
nand U7727 (N_7727,N_7410,N_7255);
nor U7728 (N_7728,N_7291,N_7416);
nand U7729 (N_7729,N_7474,N_7445);
nand U7730 (N_7730,N_7254,N_7330);
nor U7731 (N_7731,N_7474,N_7264);
or U7732 (N_7732,N_7342,N_7367);
and U7733 (N_7733,N_7437,N_7463);
or U7734 (N_7734,N_7293,N_7343);
nor U7735 (N_7735,N_7414,N_7422);
xnor U7736 (N_7736,N_7280,N_7348);
and U7737 (N_7737,N_7497,N_7326);
or U7738 (N_7738,N_7359,N_7282);
nand U7739 (N_7739,N_7410,N_7395);
or U7740 (N_7740,N_7479,N_7251);
nor U7741 (N_7741,N_7299,N_7300);
nand U7742 (N_7742,N_7429,N_7336);
nand U7743 (N_7743,N_7372,N_7252);
or U7744 (N_7744,N_7453,N_7376);
and U7745 (N_7745,N_7484,N_7267);
xnor U7746 (N_7746,N_7299,N_7384);
and U7747 (N_7747,N_7486,N_7302);
or U7748 (N_7748,N_7359,N_7273);
nand U7749 (N_7749,N_7326,N_7441);
nand U7750 (N_7750,N_7624,N_7708);
or U7751 (N_7751,N_7566,N_7688);
nand U7752 (N_7752,N_7580,N_7568);
nand U7753 (N_7753,N_7735,N_7594);
nor U7754 (N_7754,N_7672,N_7631);
nand U7755 (N_7755,N_7715,N_7733);
nand U7756 (N_7756,N_7542,N_7643);
or U7757 (N_7757,N_7510,N_7610);
or U7758 (N_7758,N_7554,N_7506);
and U7759 (N_7759,N_7587,N_7679);
xnor U7760 (N_7760,N_7501,N_7584);
or U7761 (N_7761,N_7727,N_7555);
nor U7762 (N_7762,N_7619,N_7695);
xnor U7763 (N_7763,N_7623,N_7627);
nor U7764 (N_7764,N_7591,N_7700);
xnor U7765 (N_7765,N_7660,N_7536);
and U7766 (N_7766,N_7678,N_7663);
and U7767 (N_7767,N_7730,N_7535);
xnor U7768 (N_7768,N_7504,N_7702);
and U7769 (N_7769,N_7686,N_7551);
and U7770 (N_7770,N_7714,N_7519);
or U7771 (N_7771,N_7692,N_7737);
and U7772 (N_7772,N_7509,N_7633);
and U7773 (N_7773,N_7515,N_7603);
nor U7774 (N_7774,N_7673,N_7719);
or U7775 (N_7775,N_7560,N_7683);
nand U7776 (N_7776,N_7634,N_7701);
nor U7777 (N_7777,N_7729,N_7725);
or U7778 (N_7778,N_7629,N_7693);
or U7779 (N_7779,N_7606,N_7516);
nand U7780 (N_7780,N_7508,N_7647);
and U7781 (N_7781,N_7649,N_7710);
nand U7782 (N_7782,N_7637,N_7636);
xnor U7783 (N_7783,N_7675,N_7538);
xnor U7784 (N_7784,N_7747,N_7617);
or U7785 (N_7785,N_7639,N_7746);
or U7786 (N_7786,N_7680,N_7572);
nor U7787 (N_7787,N_7593,N_7529);
or U7788 (N_7788,N_7709,N_7685);
and U7789 (N_7789,N_7728,N_7583);
and U7790 (N_7790,N_7706,N_7615);
nor U7791 (N_7791,N_7716,N_7711);
nor U7792 (N_7792,N_7502,N_7597);
or U7793 (N_7793,N_7612,N_7520);
xor U7794 (N_7794,N_7723,N_7704);
and U7795 (N_7795,N_7736,N_7565);
or U7796 (N_7796,N_7689,N_7563);
or U7797 (N_7797,N_7534,N_7684);
or U7798 (N_7798,N_7674,N_7595);
nor U7799 (N_7799,N_7577,N_7544);
or U7800 (N_7800,N_7525,N_7605);
and U7801 (N_7801,N_7697,N_7666);
xnor U7802 (N_7802,N_7540,N_7552);
nor U7803 (N_7803,N_7651,N_7656);
or U7804 (N_7804,N_7654,N_7588);
and U7805 (N_7805,N_7665,N_7528);
or U7806 (N_7806,N_7599,N_7550);
nand U7807 (N_7807,N_7734,N_7500);
nand U7808 (N_7808,N_7713,N_7640);
nor U7809 (N_7809,N_7720,N_7531);
and U7810 (N_7810,N_7726,N_7748);
and U7811 (N_7811,N_7628,N_7642);
and U7812 (N_7812,N_7682,N_7614);
and U7813 (N_7813,N_7658,N_7703);
or U7814 (N_7814,N_7626,N_7621);
nor U7815 (N_7815,N_7546,N_7681);
nand U7816 (N_7816,N_7718,N_7569);
nor U7817 (N_7817,N_7611,N_7741);
nor U7818 (N_7818,N_7575,N_7644);
or U7819 (N_7819,N_7590,N_7645);
or U7820 (N_7820,N_7514,N_7596);
or U7821 (N_7821,N_7592,N_7669);
nand U7822 (N_7822,N_7705,N_7690);
xnor U7823 (N_7823,N_7582,N_7671);
or U7824 (N_7824,N_7625,N_7613);
and U7825 (N_7825,N_7607,N_7668);
nand U7826 (N_7826,N_7574,N_7586);
and U7827 (N_7827,N_7537,N_7521);
or U7828 (N_7828,N_7602,N_7707);
nor U7829 (N_7829,N_7653,N_7561);
nand U7830 (N_7830,N_7739,N_7717);
and U7831 (N_7831,N_7567,N_7632);
nor U7832 (N_7832,N_7712,N_7664);
nand U7833 (N_7833,N_7573,N_7532);
or U7834 (N_7834,N_7698,N_7524);
and U7835 (N_7835,N_7559,N_7539);
xor U7836 (N_7836,N_7526,N_7740);
nor U7837 (N_7837,N_7601,N_7696);
nor U7838 (N_7838,N_7609,N_7676);
and U7839 (N_7839,N_7608,N_7533);
or U7840 (N_7840,N_7570,N_7722);
or U7841 (N_7841,N_7511,N_7579);
or U7842 (N_7842,N_7505,N_7677);
and U7843 (N_7843,N_7512,N_7589);
or U7844 (N_7844,N_7523,N_7557);
nand U7845 (N_7845,N_7522,N_7742);
nand U7846 (N_7846,N_7691,N_7721);
nand U7847 (N_7847,N_7507,N_7630);
nand U7848 (N_7848,N_7738,N_7518);
or U7849 (N_7849,N_7659,N_7745);
xor U7850 (N_7850,N_7641,N_7662);
xnor U7851 (N_7851,N_7517,N_7556);
nand U7852 (N_7852,N_7558,N_7600);
nand U7853 (N_7853,N_7650,N_7646);
xnor U7854 (N_7854,N_7553,N_7667);
or U7855 (N_7855,N_7622,N_7530);
nor U7856 (N_7856,N_7571,N_7699);
or U7857 (N_7857,N_7657,N_7616);
nand U7858 (N_7858,N_7604,N_7513);
and U7859 (N_7859,N_7749,N_7576);
nand U7860 (N_7860,N_7620,N_7694);
nor U7861 (N_7861,N_7562,N_7547);
and U7862 (N_7862,N_7541,N_7578);
or U7863 (N_7863,N_7648,N_7731);
nand U7864 (N_7864,N_7549,N_7548);
or U7865 (N_7865,N_7545,N_7655);
nand U7866 (N_7866,N_7687,N_7652);
or U7867 (N_7867,N_7743,N_7732);
nand U7868 (N_7868,N_7635,N_7598);
and U7869 (N_7869,N_7527,N_7503);
nor U7870 (N_7870,N_7564,N_7661);
xor U7871 (N_7871,N_7581,N_7670);
nor U7872 (N_7872,N_7638,N_7543);
or U7873 (N_7873,N_7744,N_7585);
nor U7874 (N_7874,N_7618,N_7724);
or U7875 (N_7875,N_7617,N_7525);
nand U7876 (N_7876,N_7643,N_7510);
nor U7877 (N_7877,N_7665,N_7696);
nand U7878 (N_7878,N_7644,N_7648);
and U7879 (N_7879,N_7665,N_7722);
and U7880 (N_7880,N_7700,N_7633);
nor U7881 (N_7881,N_7747,N_7746);
nand U7882 (N_7882,N_7529,N_7657);
and U7883 (N_7883,N_7500,N_7745);
and U7884 (N_7884,N_7719,N_7630);
nand U7885 (N_7885,N_7666,N_7626);
nor U7886 (N_7886,N_7665,N_7545);
nor U7887 (N_7887,N_7632,N_7718);
nor U7888 (N_7888,N_7631,N_7696);
nor U7889 (N_7889,N_7533,N_7731);
nor U7890 (N_7890,N_7518,N_7732);
and U7891 (N_7891,N_7709,N_7546);
nor U7892 (N_7892,N_7646,N_7670);
xor U7893 (N_7893,N_7655,N_7611);
and U7894 (N_7894,N_7654,N_7719);
and U7895 (N_7895,N_7629,N_7700);
xnor U7896 (N_7896,N_7615,N_7593);
and U7897 (N_7897,N_7626,N_7615);
and U7898 (N_7898,N_7680,N_7593);
and U7899 (N_7899,N_7620,N_7680);
nand U7900 (N_7900,N_7564,N_7722);
and U7901 (N_7901,N_7657,N_7587);
xor U7902 (N_7902,N_7637,N_7635);
and U7903 (N_7903,N_7676,N_7608);
nand U7904 (N_7904,N_7616,N_7549);
nand U7905 (N_7905,N_7605,N_7695);
nand U7906 (N_7906,N_7622,N_7510);
nor U7907 (N_7907,N_7572,N_7731);
xnor U7908 (N_7908,N_7613,N_7703);
or U7909 (N_7909,N_7678,N_7509);
nor U7910 (N_7910,N_7557,N_7708);
nor U7911 (N_7911,N_7648,N_7561);
nand U7912 (N_7912,N_7520,N_7699);
nand U7913 (N_7913,N_7574,N_7709);
and U7914 (N_7914,N_7683,N_7689);
nand U7915 (N_7915,N_7571,N_7666);
or U7916 (N_7916,N_7690,N_7501);
xnor U7917 (N_7917,N_7743,N_7618);
nor U7918 (N_7918,N_7531,N_7643);
xnor U7919 (N_7919,N_7643,N_7602);
nor U7920 (N_7920,N_7688,N_7551);
nand U7921 (N_7921,N_7701,N_7738);
xor U7922 (N_7922,N_7657,N_7605);
nor U7923 (N_7923,N_7722,N_7641);
xnor U7924 (N_7924,N_7618,N_7644);
and U7925 (N_7925,N_7633,N_7681);
and U7926 (N_7926,N_7530,N_7630);
nand U7927 (N_7927,N_7569,N_7610);
nand U7928 (N_7928,N_7648,N_7527);
xor U7929 (N_7929,N_7598,N_7608);
nor U7930 (N_7930,N_7742,N_7568);
and U7931 (N_7931,N_7630,N_7563);
and U7932 (N_7932,N_7664,N_7697);
nor U7933 (N_7933,N_7659,N_7671);
or U7934 (N_7934,N_7723,N_7733);
nand U7935 (N_7935,N_7701,N_7691);
xor U7936 (N_7936,N_7567,N_7688);
or U7937 (N_7937,N_7672,N_7675);
nor U7938 (N_7938,N_7654,N_7601);
or U7939 (N_7939,N_7554,N_7626);
nand U7940 (N_7940,N_7537,N_7544);
and U7941 (N_7941,N_7584,N_7510);
nand U7942 (N_7942,N_7665,N_7590);
nor U7943 (N_7943,N_7607,N_7748);
nand U7944 (N_7944,N_7584,N_7574);
or U7945 (N_7945,N_7552,N_7558);
nor U7946 (N_7946,N_7502,N_7713);
or U7947 (N_7947,N_7556,N_7672);
and U7948 (N_7948,N_7525,N_7503);
or U7949 (N_7949,N_7620,N_7558);
or U7950 (N_7950,N_7558,N_7574);
nor U7951 (N_7951,N_7739,N_7672);
or U7952 (N_7952,N_7712,N_7584);
and U7953 (N_7953,N_7516,N_7687);
and U7954 (N_7954,N_7673,N_7683);
and U7955 (N_7955,N_7597,N_7551);
or U7956 (N_7956,N_7727,N_7730);
nand U7957 (N_7957,N_7528,N_7706);
nand U7958 (N_7958,N_7672,N_7735);
xor U7959 (N_7959,N_7534,N_7703);
nor U7960 (N_7960,N_7519,N_7646);
xnor U7961 (N_7961,N_7716,N_7565);
nor U7962 (N_7962,N_7574,N_7671);
nand U7963 (N_7963,N_7607,N_7617);
or U7964 (N_7964,N_7691,N_7730);
and U7965 (N_7965,N_7670,N_7744);
nand U7966 (N_7966,N_7717,N_7592);
and U7967 (N_7967,N_7563,N_7514);
nor U7968 (N_7968,N_7547,N_7720);
xnor U7969 (N_7969,N_7728,N_7722);
nor U7970 (N_7970,N_7713,N_7506);
or U7971 (N_7971,N_7510,N_7526);
nor U7972 (N_7972,N_7626,N_7623);
nand U7973 (N_7973,N_7624,N_7669);
nand U7974 (N_7974,N_7645,N_7510);
nor U7975 (N_7975,N_7624,N_7553);
and U7976 (N_7976,N_7718,N_7558);
and U7977 (N_7977,N_7742,N_7720);
nor U7978 (N_7978,N_7748,N_7502);
nor U7979 (N_7979,N_7588,N_7500);
nand U7980 (N_7980,N_7636,N_7525);
xor U7981 (N_7981,N_7550,N_7741);
nor U7982 (N_7982,N_7573,N_7602);
and U7983 (N_7983,N_7567,N_7507);
or U7984 (N_7984,N_7689,N_7719);
and U7985 (N_7985,N_7603,N_7597);
nor U7986 (N_7986,N_7747,N_7642);
and U7987 (N_7987,N_7616,N_7518);
nand U7988 (N_7988,N_7657,N_7577);
nand U7989 (N_7989,N_7746,N_7569);
xnor U7990 (N_7990,N_7667,N_7585);
and U7991 (N_7991,N_7662,N_7575);
and U7992 (N_7992,N_7571,N_7722);
nor U7993 (N_7993,N_7650,N_7679);
or U7994 (N_7994,N_7680,N_7678);
xor U7995 (N_7995,N_7717,N_7516);
or U7996 (N_7996,N_7702,N_7637);
nand U7997 (N_7997,N_7657,N_7735);
or U7998 (N_7998,N_7566,N_7706);
or U7999 (N_7999,N_7702,N_7554);
nand U8000 (N_8000,N_7839,N_7957);
and U8001 (N_8001,N_7928,N_7791);
nor U8002 (N_8002,N_7809,N_7794);
xor U8003 (N_8003,N_7847,N_7857);
nand U8004 (N_8004,N_7862,N_7906);
nor U8005 (N_8005,N_7821,N_7764);
nand U8006 (N_8006,N_7878,N_7796);
or U8007 (N_8007,N_7785,N_7851);
nand U8008 (N_8008,N_7881,N_7844);
nor U8009 (N_8009,N_7867,N_7769);
or U8010 (N_8010,N_7978,N_7982);
and U8011 (N_8011,N_7830,N_7900);
and U8012 (N_8012,N_7907,N_7870);
nand U8013 (N_8013,N_7858,N_7916);
xnor U8014 (N_8014,N_7751,N_7920);
and U8015 (N_8015,N_7866,N_7997);
xor U8016 (N_8016,N_7893,N_7902);
or U8017 (N_8017,N_7974,N_7938);
xor U8018 (N_8018,N_7989,N_7832);
nor U8019 (N_8019,N_7776,N_7868);
nand U8020 (N_8020,N_7942,N_7967);
and U8021 (N_8021,N_7812,N_7973);
nor U8022 (N_8022,N_7763,N_7879);
nand U8023 (N_8023,N_7940,N_7865);
nor U8024 (N_8024,N_7772,N_7784);
nand U8025 (N_8025,N_7898,N_7930);
nand U8026 (N_8026,N_7932,N_7886);
and U8027 (N_8027,N_7759,N_7952);
nor U8028 (N_8028,N_7833,N_7810);
and U8029 (N_8029,N_7922,N_7929);
and U8030 (N_8030,N_7990,N_7753);
or U8031 (N_8031,N_7792,N_7890);
nand U8032 (N_8032,N_7768,N_7816);
nand U8033 (N_8033,N_7853,N_7789);
nand U8034 (N_8034,N_7939,N_7991);
nor U8035 (N_8035,N_7934,N_7927);
and U8036 (N_8036,N_7935,N_7959);
nand U8037 (N_8037,N_7971,N_7852);
and U8038 (N_8038,N_7774,N_7885);
and U8039 (N_8039,N_7909,N_7761);
and U8040 (N_8040,N_7854,N_7958);
nand U8041 (N_8041,N_7883,N_7856);
or U8042 (N_8042,N_7754,N_7950);
nor U8043 (N_8043,N_7861,N_7814);
and U8044 (N_8044,N_7871,N_7976);
and U8045 (N_8045,N_7756,N_7966);
nand U8046 (N_8046,N_7889,N_7855);
and U8047 (N_8047,N_7829,N_7919);
nand U8048 (N_8048,N_7828,N_7985);
nor U8049 (N_8049,N_7823,N_7888);
or U8050 (N_8050,N_7846,N_7797);
nor U8051 (N_8051,N_7820,N_7944);
or U8052 (N_8052,N_7790,N_7918);
nand U8053 (N_8053,N_7903,N_7795);
and U8054 (N_8054,N_7804,N_7943);
or U8055 (N_8055,N_7936,N_7838);
or U8056 (N_8056,N_7988,N_7801);
and U8057 (N_8057,N_7783,N_7896);
or U8058 (N_8058,N_7782,N_7987);
and U8059 (N_8059,N_7945,N_7937);
and U8060 (N_8060,N_7755,N_7806);
and U8061 (N_8061,N_7824,N_7762);
nor U8062 (N_8062,N_7779,N_7891);
or U8063 (N_8063,N_7897,N_7908);
or U8064 (N_8064,N_7970,N_7981);
or U8065 (N_8065,N_7895,N_7775);
nand U8066 (N_8066,N_7825,N_7994);
or U8067 (N_8067,N_7771,N_7901);
or U8068 (N_8068,N_7880,N_7758);
and U8069 (N_8069,N_7941,N_7805);
or U8070 (N_8070,N_7904,N_7849);
nand U8071 (N_8071,N_7983,N_7815);
nor U8072 (N_8072,N_7822,N_7864);
nand U8073 (N_8073,N_7946,N_7803);
or U8074 (N_8074,N_7962,N_7837);
nand U8075 (N_8075,N_7875,N_7882);
xnor U8076 (N_8076,N_7786,N_7874);
nand U8077 (N_8077,N_7819,N_7811);
or U8078 (N_8078,N_7826,N_7793);
or U8079 (N_8079,N_7817,N_7905);
or U8080 (N_8080,N_7915,N_7788);
nor U8081 (N_8081,N_7965,N_7841);
or U8082 (N_8082,N_7910,N_7876);
xnor U8083 (N_8083,N_7813,N_7963);
or U8084 (N_8084,N_7781,N_7912);
and U8085 (N_8085,N_7859,N_7750);
xnor U8086 (N_8086,N_7827,N_7873);
and U8087 (N_8087,N_7848,N_7926);
nor U8088 (N_8088,N_7760,N_7887);
and U8089 (N_8089,N_7787,N_7773);
or U8090 (N_8090,N_7960,N_7992);
nand U8091 (N_8091,N_7770,N_7984);
and U8092 (N_8092,N_7986,N_7850);
nor U8093 (N_8093,N_7835,N_7951);
or U8094 (N_8094,N_7947,N_7969);
and U8095 (N_8095,N_7802,N_7899);
xor U8096 (N_8096,N_7818,N_7765);
nor U8097 (N_8097,N_7860,N_7993);
and U8098 (N_8098,N_7757,N_7834);
and U8099 (N_8099,N_7869,N_7955);
and U8100 (N_8100,N_7914,N_7799);
nor U8101 (N_8101,N_7842,N_7949);
and U8102 (N_8102,N_7933,N_7923);
nor U8103 (N_8103,N_7980,N_7931);
or U8104 (N_8104,N_7863,N_7766);
and U8105 (N_8105,N_7998,N_7975);
nand U8106 (N_8106,N_7948,N_7892);
or U8107 (N_8107,N_7954,N_7843);
xor U8108 (N_8108,N_7831,N_7961);
and U8109 (N_8109,N_7798,N_7964);
nor U8110 (N_8110,N_7925,N_7872);
nor U8111 (N_8111,N_7808,N_7972);
xnor U8112 (N_8112,N_7894,N_7996);
and U8113 (N_8113,N_7956,N_7752);
nor U8114 (N_8114,N_7845,N_7877);
nand U8115 (N_8115,N_7924,N_7800);
nor U8116 (N_8116,N_7995,N_7840);
or U8117 (N_8117,N_7968,N_7921);
nand U8118 (N_8118,N_7979,N_7999);
and U8119 (N_8119,N_7767,N_7977);
and U8120 (N_8120,N_7780,N_7807);
or U8121 (N_8121,N_7917,N_7911);
nor U8122 (N_8122,N_7884,N_7836);
nor U8123 (N_8123,N_7953,N_7777);
nor U8124 (N_8124,N_7913,N_7778);
nand U8125 (N_8125,N_7952,N_7967);
nor U8126 (N_8126,N_7983,N_7917);
and U8127 (N_8127,N_7912,N_7981);
nor U8128 (N_8128,N_7909,N_7927);
and U8129 (N_8129,N_7761,N_7809);
nor U8130 (N_8130,N_7873,N_7962);
nand U8131 (N_8131,N_7978,N_7993);
and U8132 (N_8132,N_7753,N_7798);
nor U8133 (N_8133,N_7862,N_7785);
and U8134 (N_8134,N_7860,N_7985);
or U8135 (N_8135,N_7986,N_7836);
nand U8136 (N_8136,N_7923,N_7884);
nor U8137 (N_8137,N_7894,N_7946);
and U8138 (N_8138,N_7842,N_7957);
or U8139 (N_8139,N_7928,N_7869);
nand U8140 (N_8140,N_7972,N_7950);
or U8141 (N_8141,N_7809,N_7814);
nor U8142 (N_8142,N_7981,N_7774);
nand U8143 (N_8143,N_7853,N_7870);
and U8144 (N_8144,N_7761,N_7988);
or U8145 (N_8145,N_7831,N_7956);
or U8146 (N_8146,N_7782,N_7920);
xnor U8147 (N_8147,N_7846,N_7989);
nor U8148 (N_8148,N_7948,N_7846);
and U8149 (N_8149,N_7977,N_7946);
nor U8150 (N_8150,N_7929,N_7788);
nor U8151 (N_8151,N_7765,N_7756);
nor U8152 (N_8152,N_7827,N_7984);
or U8153 (N_8153,N_7751,N_7966);
and U8154 (N_8154,N_7804,N_7789);
or U8155 (N_8155,N_7963,N_7782);
or U8156 (N_8156,N_7943,N_7996);
or U8157 (N_8157,N_7946,N_7929);
nand U8158 (N_8158,N_7818,N_7886);
nor U8159 (N_8159,N_7896,N_7820);
nand U8160 (N_8160,N_7770,N_7819);
and U8161 (N_8161,N_7866,N_7956);
xor U8162 (N_8162,N_7971,N_7908);
nor U8163 (N_8163,N_7812,N_7952);
nor U8164 (N_8164,N_7781,N_7850);
xor U8165 (N_8165,N_7855,N_7802);
nand U8166 (N_8166,N_7931,N_7863);
and U8167 (N_8167,N_7929,N_7801);
nor U8168 (N_8168,N_7841,N_7825);
nor U8169 (N_8169,N_7775,N_7938);
and U8170 (N_8170,N_7859,N_7795);
nor U8171 (N_8171,N_7834,N_7817);
and U8172 (N_8172,N_7804,N_7959);
xnor U8173 (N_8173,N_7833,N_7782);
or U8174 (N_8174,N_7815,N_7820);
or U8175 (N_8175,N_7823,N_7957);
or U8176 (N_8176,N_7880,N_7975);
nand U8177 (N_8177,N_7940,N_7772);
or U8178 (N_8178,N_7894,N_7950);
or U8179 (N_8179,N_7857,N_7770);
and U8180 (N_8180,N_7923,N_7988);
nor U8181 (N_8181,N_7888,N_7852);
and U8182 (N_8182,N_7799,N_7942);
nand U8183 (N_8183,N_7922,N_7914);
nor U8184 (N_8184,N_7763,N_7784);
nor U8185 (N_8185,N_7861,N_7862);
or U8186 (N_8186,N_7791,N_7936);
and U8187 (N_8187,N_7966,N_7763);
nor U8188 (N_8188,N_7980,N_7799);
or U8189 (N_8189,N_7759,N_7769);
nor U8190 (N_8190,N_7800,N_7825);
or U8191 (N_8191,N_7820,N_7810);
and U8192 (N_8192,N_7859,N_7804);
or U8193 (N_8193,N_7925,N_7906);
or U8194 (N_8194,N_7909,N_7977);
nor U8195 (N_8195,N_7769,N_7809);
nand U8196 (N_8196,N_7776,N_7881);
nand U8197 (N_8197,N_7894,N_7881);
or U8198 (N_8198,N_7808,N_7769);
and U8199 (N_8199,N_7890,N_7958);
nand U8200 (N_8200,N_7844,N_7836);
nand U8201 (N_8201,N_7779,N_7769);
or U8202 (N_8202,N_7898,N_7944);
nand U8203 (N_8203,N_7979,N_7862);
nor U8204 (N_8204,N_7860,N_7859);
xor U8205 (N_8205,N_7887,N_7952);
nand U8206 (N_8206,N_7870,N_7862);
nor U8207 (N_8207,N_7868,N_7790);
or U8208 (N_8208,N_7808,N_7871);
xor U8209 (N_8209,N_7987,N_7856);
nand U8210 (N_8210,N_7854,N_7756);
nor U8211 (N_8211,N_7922,N_7949);
or U8212 (N_8212,N_7835,N_7781);
nand U8213 (N_8213,N_7989,N_7825);
or U8214 (N_8214,N_7860,N_7963);
nor U8215 (N_8215,N_7985,N_7923);
and U8216 (N_8216,N_7830,N_7848);
or U8217 (N_8217,N_7967,N_7868);
and U8218 (N_8218,N_7842,N_7931);
or U8219 (N_8219,N_7909,N_7771);
nand U8220 (N_8220,N_7817,N_7822);
or U8221 (N_8221,N_7779,N_7873);
nand U8222 (N_8222,N_7974,N_7904);
nor U8223 (N_8223,N_7861,N_7984);
and U8224 (N_8224,N_7819,N_7891);
or U8225 (N_8225,N_7992,N_7930);
nand U8226 (N_8226,N_7979,N_7798);
xor U8227 (N_8227,N_7831,N_7812);
or U8228 (N_8228,N_7816,N_7887);
xor U8229 (N_8229,N_7983,N_7999);
nor U8230 (N_8230,N_7773,N_7906);
or U8231 (N_8231,N_7929,N_7995);
xor U8232 (N_8232,N_7769,N_7822);
and U8233 (N_8233,N_7963,N_7755);
nand U8234 (N_8234,N_7962,N_7858);
nand U8235 (N_8235,N_7843,N_7824);
nor U8236 (N_8236,N_7876,N_7977);
xnor U8237 (N_8237,N_7979,N_7759);
nor U8238 (N_8238,N_7789,N_7866);
nand U8239 (N_8239,N_7868,N_7833);
nor U8240 (N_8240,N_7956,N_7809);
or U8241 (N_8241,N_7994,N_7919);
and U8242 (N_8242,N_7841,N_7816);
or U8243 (N_8243,N_7772,N_7833);
and U8244 (N_8244,N_7752,N_7806);
or U8245 (N_8245,N_7768,N_7864);
or U8246 (N_8246,N_7915,N_7892);
xor U8247 (N_8247,N_7949,N_7770);
or U8248 (N_8248,N_7980,N_7779);
nand U8249 (N_8249,N_7954,N_7859);
or U8250 (N_8250,N_8037,N_8174);
nand U8251 (N_8251,N_8054,N_8212);
or U8252 (N_8252,N_8147,N_8193);
or U8253 (N_8253,N_8041,N_8146);
and U8254 (N_8254,N_8009,N_8097);
or U8255 (N_8255,N_8157,N_8005);
or U8256 (N_8256,N_8040,N_8078);
nand U8257 (N_8257,N_8124,N_8044);
nor U8258 (N_8258,N_8154,N_8080);
nand U8259 (N_8259,N_8083,N_8108);
nor U8260 (N_8260,N_8087,N_8191);
and U8261 (N_8261,N_8067,N_8069);
and U8262 (N_8262,N_8033,N_8053);
and U8263 (N_8263,N_8002,N_8035);
nor U8264 (N_8264,N_8222,N_8130);
nor U8265 (N_8265,N_8221,N_8144);
xnor U8266 (N_8266,N_8224,N_8110);
nor U8267 (N_8267,N_8086,N_8123);
or U8268 (N_8268,N_8202,N_8122);
or U8269 (N_8269,N_8249,N_8014);
or U8270 (N_8270,N_8045,N_8017);
nand U8271 (N_8271,N_8062,N_8029);
nor U8272 (N_8272,N_8127,N_8020);
and U8273 (N_8273,N_8190,N_8197);
nand U8274 (N_8274,N_8194,N_8102);
or U8275 (N_8275,N_8021,N_8074);
nor U8276 (N_8276,N_8213,N_8139);
nor U8277 (N_8277,N_8056,N_8138);
nand U8278 (N_8278,N_8117,N_8200);
nor U8279 (N_8279,N_8066,N_8039);
nand U8280 (N_8280,N_8211,N_8125);
xnor U8281 (N_8281,N_8246,N_8186);
nor U8282 (N_8282,N_8244,N_8068);
xnor U8283 (N_8283,N_8132,N_8073);
nor U8284 (N_8284,N_8134,N_8077);
and U8285 (N_8285,N_8092,N_8170);
or U8286 (N_8286,N_8131,N_8145);
or U8287 (N_8287,N_8004,N_8115);
nand U8288 (N_8288,N_8236,N_8024);
nor U8289 (N_8289,N_8046,N_8215);
or U8290 (N_8290,N_8217,N_8176);
and U8291 (N_8291,N_8049,N_8149);
xnor U8292 (N_8292,N_8114,N_8103);
nand U8293 (N_8293,N_8047,N_8223);
or U8294 (N_8294,N_8084,N_8000);
nor U8295 (N_8295,N_8019,N_8173);
and U8296 (N_8296,N_8133,N_8248);
nand U8297 (N_8297,N_8048,N_8022);
nand U8298 (N_8298,N_8185,N_8028);
or U8299 (N_8299,N_8226,N_8175);
nor U8300 (N_8300,N_8161,N_8172);
or U8301 (N_8301,N_8129,N_8093);
and U8302 (N_8302,N_8201,N_8106);
and U8303 (N_8303,N_8234,N_8027);
or U8304 (N_8304,N_8198,N_8012);
nand U8305 (N_8305,N_8071,N_8099);
or U8306 (N_8306,N_8150,N_8142);
and U8307 (N_8307,N_8178,N_8109);
xor U8308 (N_8308,N_8003,N_8043);
or U8309 (N_8309,N_8206,N_8113);
xor U8310 (N_8310,N_8079,N_8239);
xnor U8311 (N_8311,N_8195,N_8081);
nand U8312 (N_8312,N_8082,N_8156);
nand U8313 (N_8313,N_8231,N_8038);
nor U8314 (N_8314,N_8025,N_8160);
or U8315 (N_8315,N_8180,N_8183);
and U8316 (N_8316,N_8192,N_8100);
nor U8317 (N_8317,N_8036,N_8060);
nand U8318 (N_8318,N_8001,N_8107);
nand U8319 (N_8319,N_8241,N_8119);
and U8320 (N_8320,N_8118,N_8076);
or U8321 (N_8321,N_8013,N_8187);
xor U8322 (N_8322,N_8225,N_8207);
or U8323 (N_8323,N_8152,N_8089);
nor U8324 (N_8324,N_8143,N_8075);
nand U8325 (N_8325,N_8164,N_8232);
xor U8326 (N_8326,N_8235,N_8171);
or U8327 (N_8327,N_8210,N_8196);
or U8328 (N_8328,N_8016,N_8059);
nor U8329 (N_8329,N_8011,N_8165);
nor U8330 (N_8330,N_8141,N_8010);
and U8331 (N_8331,N_8018,N_8237);
nor U8332 (N_8332,N_8051,N_8026);
and U8333 (N_8333,N_8101,N_8179);
nand U8334 (N_8334,N_8162,N_8209);
nand U8335 (N_8335,N_8218,N_8163);
or U8336 (N_8336,N_8182,N_8243);
nor U8337 (N_8337,N_8065,N_8058);
nand U8338 (N_8338,N_8184,N_8168);
nand U8339 (N_8339,N_8121,N_8216);
nor U8340 (N_8340,N_8096,N_8055);
nand U8341 (N_8341,N_8155,N_8167);
and U8342 (N_8342,N_8135,N_8030);
xor U8343 (N_8343,N_8085,N_8137);
or U8344 (N_8344,N_8188,N_8032);
and U8345 (N_8345,N_8151,N_8088);
or U8346 (N_8346,N_8240,N_8219);
xor U8347 (N_8347,N_8064,N_8189);
nand U8348 (N_8348,N_8238,N_8204);
nand U8349 (N_8349,N_8140,N_8159);
or U8350 (N_8350,N_8090,N_8111);
nand U8351 (N_8351,N_8242,N_8112);
nand U8352 (N_8352,N_8247,N_8072);
and U8353 (N_8353,N_8128,N_8148);
and U8354 (N_8354,N_8008,N_8034);
or U8355 (N_8355,N_8042,N_8061);
and U8356 (N_8356,N_8057,N_8166);
or U8357 (N_8357,N_8105,N_8052);
or U8358 (N_8358,N_8098,N_8208);
or U8359 (N_8359,N_8126,N_8214);
nand U8360 (N_8360,N_8094,N_8050);
nor U8361 (N_8361,N_8199,N_8181);
nand U8362 (N_8362,N_8136,N_8177);
and U8363 (N_8363,N_8203,N_8233);
xor U8364 (N_8364,N_8007,N_8104);
nor U8365 (N_8365,N_8153,N_8169);
nor U8366 (N_8366,N_8228,N_8227);
nor U8367 (N_8367,N_8229,N_8205);
nand U8368 (N_8368,N_8023,N_8158);
or U8369 (N_8369,N_8230,N_8120);
nand U8370 (N_8370,N_8063,N_8031);
and U8371 (N_8371,N_8015,N_8116);
nand U8372 (N_8372,N_8091,N_8220);
nor U8373 (N_8373,N_8095,N_8006);
or U8374 (N_8374,N_8070,N_8245);
nor U8375 (N_8375,N_8240,N_8064);
or U8376 (N_8376,N_8228,N_8233);
nor U8377 (N_8377,N_8134,N_8026);
nor U8378 (N_8378,N_8201,N_8119);
and U8379 (N_8379,N_8113,N_8005);
nor U8380 (N_8380,N_8110,N_8121);
xnor U8381 (N_8381,N_8055,N_8051);
nor U8382 (N_8382,N_8195,N_8168);
or U8383 (N_8383,N_8102,N_8108);
nand U8384 (N_8384,N_8130,N_8136);
nand U8385 (N_8385,N_8111,N_8198);
nand U8386 (N_8386,N_8151,N_8133);
nor U8387 (N_8387,N_8220,N_8236);
or U8388 (N_8388,N_8093,N_8133);
xor U8389 (N_8389,N_8164,N_8145);
nand U8390 (N_8390,N_8074,N_8184);
and U8391 (N_8391,N_8136,N_8040);
nor U8392 (N_8392,N_8182,N_8003);
nand U8393 (N_8393,N_8197,N_8021);
xor U8394 (N_8394,N_8216,N_8207);
nand U8395 (N_8395,N_8112,N_8187);
nor U8396 (N_8396,N_8030,N_8194);
nand U8397 (N_8397,N_8160,N_8063);
xnor U8398 (N_8398,N_8209,N_8241);
or U8399 (N_8399,N_8078,N_8099);
nand U8400 (N_8400,N_8114,N_8208);
nor U8401 (N_8401,N_8037,N_8164);
and U8402 (N_8402,N_8220,N_8149);
nand U8403 (N_8403,N_8247,N_8141);
or U8404 (N_8404,N_8194,N_8237);
nor U8405 (N_8405,N_8189,N_8090);
and U8406 (N_8406,N_8024,N_8015);
nor U8407 (N_8407,N_8053,N_8125);
nand U8408 (N_8408,N_8235,N_8173);
xnor U8409 (N_8409,N_8062,N_8076);
xor U8410 (N_8410,N_8013,N_8045);
and U8411 (N_8411,N_8016,N_8100);
and U8412 (N_8412,N_8209,N_8221);
or U8413 (N_8413,N_8208,N_8076);
nand U8414 (N_8414,N_8237,N_8015);
nand U8415 (N_8415,N_8139,N_8202);
nand U8416 (N_8416,N_8164,N_8110);
and U8417 (N_8417,N_8176,N_8055);
nand U8418 (N_8418,N_8223,N_8119);
or U8419 (N_8419,N_8073,N_8097);
xor U8420 (N_8420,N_8109,N_8005);
xnor U8421 (N_8421,N_8032,N_8143);
nand U8422 (N_8422,N_8171,N_8008);
nand U8423 (N_8423,N_8165,N_8126);
or U8424 (N_8424,N_8243,N_8177);
and U8425 (N_8425,N_8044,N_8003);
nand U8426 (N_8426,N_8146,N_8119);
or U8427 (N_8427,N_8072,N_8191);
and U8428 (N_8428,N_8066,N_8038);
and U8429 (N_8429,N_8123,N_8035);
xnor U8430 (N_8430,N_8044,N_8038);
and U8431 (N_8431,N_8115,N_8104);
or U8432 (N_8432,N_8220,N_8057);
or U8433 (N_8433,N_8179,N_8016);
and U8434 (N_8434,N_8212,N_8060);
nand U8435 (N_8435,N_8128,N_8077);
xor U8436 (N_8436,N_8227,N_8128);
and U8437 (N_8437,N_8239,N_8002);
and U8438 (N_8438,N_8020,N_8185);
nand U8439 (N_8439,N_8172,N_8156);
nand U8440 (N_8440,N_8105,N_8058);
and U8441 (N_8441,N_8118,N_8129);
nand U8442 (N_8442,N_8219,N_8200);
nand U8443 (N_8443,N_8011,N_8019);
nor U8444 (N_8444,N_8000,N_8043);
nand U8445 (N_8445,N_8195,N_8179);
and U8446 (N_8446,N_8137,N_8198);
or U8447 (N_8447,N_8128,N_8197);
nand U8448 (N_8448,N_8167,N_8010);
or U8449 (N_8449,N_8112,N_8164);
and U8450 (N_8450,N_8055,N_8031);
nand U8451 (N_8451,N_8146,N_8078);
nand U8452 (N_8452,N_8237,N_8125);
xor U8453 (N_8453,N_8099,N_8140);
nand U8454 (N_8454,N_8114,N_8051);
or U8455 (N_8455,N_8190,N_8039);
and U8456 (N_8456,N_8175,N_8140);
nand U8457 (N_8457,N_8198,N_8031);
or U8458 (N_8458,N_8192,N_8058);
nor U8459 (N_8459,N_8195,N_8028);
nand U8460 (N_8460,N_8214,N_8116);
nand U8461 (N_8461,N_8054,N_8060);
or U8462 (N_8462,N_8182,N_8029);
xor U8463 (N_8463,N_8001,N_8243);
nand U8464 (N_8464,N_8118,N_8035);
nor U8465 (N_8465,N_8159,N_8025);
and U8466 (N_8466,N_8202,N_8031);
and U8467 (N_8467,N_8211,N_8077);
nand U8468 (N_8468,N_8125,N_8035);
nand U8469 (N_8469,N_8140,N_8106);
nor U8470 (N_8470,N_8080,N_8204);
xnor U8471 (N_8471,N_8060,N_8113);
or U8472 (N_8472,N_8048,N_8208);
and U8473 (N_8473,N_8102,N_8041);
or U8474 (N_8474,N_8030,N_8191);
and U8475 (N_8475,N_8019,N_8098);
nand U8476 (N_8476,N_8154,N_8023);
nor U8477 (N_8477,N_8065,N_8113);
xnor U8478 (N_8478,N_8155,N_8228);
and U8479 (N_8479,N_8106,N_8128);
nor U8480 (N_8480,N_8226,N_8141);
xnor U8481 (N_8481,N_8010,N_8096);
nor U8482 (N_8482,N_8064,N_8053);
or U8483 (N_8483,N_8021,N_8232);
xnor U8484 (N_8484,N_8048,N_8124);
nor U8485 (N_8485,N_8144,N_8207);
nor U8486 (N_8486,N_8085,N_8247);
and U8487 (N_8487,N_8033,N_8176);
nor U8488 (N_8488,N_8228,N_8186);
and U8489 (N_8489,N_8095,N_8226);
nand U8490 (N_8490,N_8017,N_8225);
and U8491 (N_8491,N_8199,N_8164);
or U8492 (N_8492,N_8184,N_8169);
xor U8493 (N_8493,N_8162,N_8165);
nor U8494 (N_8494,N_8147,N_8116);
nand U8495 (N_8495,N_8186,N_8180);
nor U8496 (N_8496,N_8097,N_8103);
nand U8497 (N_8497,N_8009,N_8192);
or U8498 (N_8498,N_8050,N_8246);
or U8499 (N_8499,N_8019,N_8042);
nor U8500 (N_8500,N_8489,N_8447);
and U8501 (N_8501,N_8479,N_8385);
or U8502 (N_8502,N_8336,N_8356);
or U8503 (N_8503,N_8254,N_8457);
and U8504 (N_8504,N_8446,N_8308);
nor U8505 (N_8505,N_8473,N_8392);
nor U8506 (N_8506,N_8430,N_8289);
or U8507 (N_8507,N_8375,N_8397);
and U8508 (N_8508,N_8335,N_8478);
and U8509 (N_8509,N_8416,N_8418);
nor U8510 (N_8510,N_8257,N_8406);
nor U8511 (N_8511,N_8367,N_8334);
and U8512 (N_8512,N_8456,N_8444);
or U8513 (N_8513,N_8287,N_8340);
or U8514 (N_8514,N_8424,N_8328);
and U8515 (N_8515,N_8346,N_8267);
and U8516 (N_8516,N_8330,N_8383);
nor U8517 (N_8517,N_8404,N_8290);
or U8518 (N_8518,N_8339,N_8445);
and U8519 (N_8519,N_8304,N_8415);
nor U8520 (N_8520,N_8437,N_8459);
nor U8521 (N_8521,N_8380,N_8493);
and U8522 (N_8522,N_8355,N_8357);
and U8523 (N_8523,N_8495,N_8372);
and U8524 (N_8524,N_8293,N_8402);
nand U8525 (N_8525,N_8496,N_8352);
nor U8526 (N_8526,N_8365,N_8343);
or U8527 (N_8527,N_8266,N_8443);
nand U8528 (N_8528,N_8256,N_8481);
xor U8529 (N_8529,N_8422,N_8258);
or U8530 (N_8530,N_8310,N_8411);
nor U8531 (N_8531,N_8265,N_8262);
nand U8532 (N_8532,N_8313,N_8429);
and U8533 (N_8533,N_8431,N_8299);
nand U8534 (N_8534,N_8464,N_8400);
nor U8535 (N_8535,N_8272,N_8433);
and U8536 (N_8536,N_8461,N_8469);
nor U8537 (N_8537,N_8408,N_8268);
or U8538 (N_8538,N_8485,N_8490);
or U8539 (N_8539,N_8323,N_8337);
and U8540 (N_8540,N_8407,N_8295);
and U8541 (N_8541,N_8492,N_8455);
nor U8542 (N_8542,N_8499,N_8453);
nand U8543 (N_8543,N_8381,N_8345);
and U8544 (N_8544,N_8307,N_8333);
and U8545 (N_8545,N_8428,N_8488);
nor U8546 (N_8546,N_8494,N_8432);
nor U8547 (N_8547,N_8306,N_8399);
nand U8548 (N_8548,N_8250,N_8466);
nor U8549 (N_8549,N_8382,N_8409);
nand U8550 (N_8550,N_8378,N_8401);
nor U8551 (N_8551,N_8362,N_8302);
and U8552 (N_8552,N_8264,N_8449);
nor U8553 (N_8553,N_8315,N_8348);
nand U8554 (N_8554,N_8482,N_8377);
nand U8555 (N_8555,N_8303,N_8475);
nand U8556 (N_8556,N_8270,N_8309);
and U8557 (N_8557,N_8439,N_8369);
nor U8558 (N_8558,N_8423,N_8320);
nand U8559 (N_8559,N_8373,N_8451);
xor U8560 (N_8560,N_8281,N_8284);
nand U8561 (N_8561,N_8487,N_8327);
nand U8562 (N_8562,N_8413,N_8465);
and U8563 (N_8563,N_8458,N_8288);
nor U8564 (N_8564,N_8435,N_8279);
and U8565 (N_8565,N_8316,N_8374);
or U8566 (N_8566,N_8338,N_8462);
or U8567 (N_8567,N_8344,N_8298);
or U8568 (N_8568,N_8483,N_8441);
or U8569 (N_8569,N_8442,N_8470);
or U8570 (N_8570,N_8468,N_8325);
and U8571 (N_8571,N_8305,N_8364);
and U8572 (N_8572,N_8476,N_8283);
nand U8573 (N_8573,N_8387,N_8434);
nand U8574 (N_8574,N_8271,N_8472);
nor U8575 (N_8575,N_8324,N_8454);
nor U8576 (N_8576,N_8425,N_8252);
nor U8577 (N_8577,N_8396,N_8426);
or U8578 (N_8578,N_8276,N_8351);
xor U8579 (N_8579,N_8341,N_8253);
and U8580 (N_8580,N_8359,N_8436);
nor U8581 (N_8581,N_8391,N_8301);
nand U8582 (N_8582,N_8312,N_8342);
xor U8583 (N_8583,N_8286,N_8412);
nor U8584 (N_8584,N_8414,N_8354);
nand U8585 (N_8585,N_8390,N_8350);
and U8586 (N_8586,N_8393,N_8370);
or U8587 (N_8587,N_8389,N_8353);
or U8588 (N_8588,N_8319,N_8280);
or U8589 (N_8589,N_8388,N_8277);
nand U8590 (N_8590,N_8300,N_8450);
nor U8591 (N_8591,N_8405,N_8296);
and U8592 (N_8592,N_8384,N_8349);
nand U8593 (N_8593,N_8297,N_8474);
nand U8594 (N_8594,N_8421,N_8419);
or U8595 (N_8595,N_8486,N_8467);
xnor U8596 (N_8596,N_8285,N_8332);
and U8597 (N_8597,N_8395,N_8292);
nor U8598 (N_8598,N_8260,N_8318);
or U8599 (N_8599,N_8278,N_8347);
or U8600 (N_8600,N_8361,N_8282);
and U8601 (N_8601,N_8366,N_8314);
nor U8602 (N_8602,N_8477,N_8321);
nand U8603 (N_8603,N_8452,N_8491);
nor U8604 (N_8604,N_8484,N_8471);
nor U8605 (N_8605,N_8294,N_8386);
nand U8606 (N_8606,N_8420,N_8261);
and U8607 (N_8607,N_8440,N_8438);
nand U8608 (N_8608,N_8360,N_8274);
nor U8609 (N_8609,N_8329,N_8498);
and U8610 (N_8610,N_8463,N_8427);
and U8611 (N_8611,N_8368,N_8273);
nand U8612 (N_8612,N_8251,N_8379);
nand U8613 (N_8613,N_8269,N_8371);
and U8614 (N_8614,N_8417,N_8322);
nor U8615 (N_8615,N_8259,N_8326);
nor U8616 (N_8616,N_8363,N_8358);
or U8617 (N_8617,N_8291,N_8376);
or U8618 (N_8618,N_8255,N_8410);
nor U8619 (N_8619,N_8394,N_8317);
and U8620 (N_8620,N_8480,N_8263);
nor U8621 (N_8621,N_8403,N_8448);
nor U8622 (N_8622,N_8460,N_8398);
and U8623 (N_8623,N_8311,N_8331);
nor U8624 (N_8624,N_8497,N_8275);
nand U8625 (N_8625,N_8483,N_8469);
and U8626 (N_8626,N_8410,N_8451);
or U8627 (N_8627,N_8445,N_8470);
or U8628 (N_8628,N_8455,N_8316);
nor U8629 (N_8629,N_8480,N_8448);
or U8630 (N_8630,N_8424,N_8472);
nand U8631 (N_8631,N_8269,N_8499);
and U8632 (N_8632,N_8364,N_8315);
or U8633 (N_8633,N_8272,N_8256);
or U8634 (N_8634,N_8333,N_8342);
nand U8635 (N_8635,N_8418,N_8488);
nand U8636 (N_8636,N_8344,N_8470);
and U8637 (N_8637,N_8438,N_8454);
nand U8638 (N_8638,N_8483,N_8254);
xnor U8639 (N_8639,N_8430,N_8358);
xor U8640 (N_8640,N_8287,N_8279);
or U8641 (N_8641,N_8361,N_8489);
or U8642 (N_8642,N_8467,N_8414);
or U8643 (N_8643,N_8380,N_8346);
nor U8644 (N_8644,N_8325,N_8465);
nor U8645 (N_8645,N_8370,N_8268);
or U8646 (N_8646,N_8492,N_8401);
and U8647 (N_8647,N_8448,N_8356);
nor U8648 (N_8648,N_8253,N_8455);
or U8649 (N_8649,N_8386,N_8486);
nand U8650 (N_8650,N_8441,N_8314);
or U8651 (N_8651,N_8423,N_8482);
nand U8652 (N_8652,N_8252,N_8354);
nor U8653 (N_8653,N_8338,N_8467);
or U8654 (N_8654,N_8322,N_8403);
and U8655 (N_8655,N_8477,N_8406);
nor U8656 (N_8656,N_8389,N_8359);
nand U8657 (N_8657,N_8292,N_8324);
and U8658 (N_8658,N_8282,N_8436);
xor U8659 (N_8659,N_8494,N_8306);
xor U8660 (N_8660,N_8414,N_8350);
nor U8661 (N_8661,N_8298,N_8435);
nand U8662 (N_8662,N_8493,N_8401);
nand U8663 (N_8663,N_8383,N_8375);
nand U8664 (N_8664,N_8298,N_8277);
xnor U8665 (N_8665,N_8259,N_8254);
and U8666 (N_8666,N_8478,N_8355);
nand U8667 (N_8667,N_8279,N_8292);
nand U8668 (N_8668,N_8391,N_8407);
and U8669 (N_8669,N_8423,N_8384);
and U8670 (N_8670,N_8492,N_8357);
xor U8671 (N_8671,N_8336,N_8394);
or U8672 (N_8672,N_8352,N_8255);
nand U8673 (N_8673,N_8353,N_8437);
nand U8674 (N_8674,N_8273,N_8404);
or U8675 (N_8675,N_8483,N_8485);
nand U8676 (N_8676,N_8418,N_8450);
xor U8677 (N_8677,N_8334,N_8417);
and U8678 (N_8678,N_8259,N_8332);
or U8679 (N_8679,N_8277,N_8372);
or U8680 (N_8680,N_8398,N_8435);
or U8681 (N_8681,N_8430,N_8311);
or U8682 (N_8682,N_8431,N_8365);
or U8683 (N_8683,N_8322,N_8425);
or U8684 (N_8684,N_8447,N_8390);
nor U8685 (N_8685,N_8412,N_8425);
or U8686 (N_8686,N_8436,N_8270);
nor U8687 (N_8687,N_8429,N_8307);
nor U8688 (N_8688,N_8471,N_8470);
nor U8689 (N_8689,N_8351,N_8361);
nand U8690 (N_8690,N_8358,N_8292);
xor U8691 (N_8691,N_8332,N_8382);
xor U8692 (N_8692,N_8367,N_8311);
or U8693 (N_8693,N_8356,N_8449);
or U8694 (N_8694,N_8265,N_8302);
and U8695 (N_8695,N_8496,N_8499);
and U8696 (N_8696,N_8341,N_8261);
nand U8697 (N_8697,N_8465,N_8341);
nand U8698 (N_8698,N_8350,N_8478);
and U8699 (N_8699,N_8480,N_8256);
xnor U8700 (N_8700,N_8397,N_8321);
nor U8701 (N_8701,N_8385,N_8301);
nand U8702 (N_8702,N_8299,N_8368);
and U8703 (N_8703,N_8302,N_8254);
nor U8704 (N_8704,N_8447,N_8292);
and U8705 (N_8705,N_8363,N_8392);
nand U8706 (N_8706,N_8345,N_8293);
nor U8707 (N_8707,N_8312,N_8395);
or U8708 (N_8708,N_8457,N_8352);
nand U8709 (N_8709,N_8407,N_8322);
xnor U8710 (N_8710,N_8271,N_8322);
nor U8711 (N_8711,N_8353,N_8311);
nor U8712 (N_8712,N_8486,N_8287);
and U8713 (N_8713,N_8420,N_8267);
xor U8714 (N_8714,N_8390,N_8333);
nand U8715 (N_8715,N_8258,N_8468);
nor U8716 (N_8716,N_8261,N_8475);
or U8717 (N_8717,N_8327,N_8359);
nand U8718 (N_8718,N_8357,N_8474);
nand U8719 (N_8719,N_8291,N_8269);
or U8720 (N_8720,N_8299,N_8388);
or U8721 (N_8721,N_8490,N_8398);
nor U8722 (N_8722,N_8304,N_8395);
or U8723 (N_8723,N_8362,N_8338);
nor U8724 (N_8724,N_8492,N_8459);
or U8725 (N_8725,N_8275,N_8286);
or U8726 (N_8726,N_8488,N_8379);
nor U8727 (N_8727,N_8321,N_8414);
nand U8728 (N_8728,N_8273,N_8385);
nor U8729 (N_8729,N_8253,N_8394);
or U8730 (N_8730,N_8378,N_8315);
or U8731 (N_8731,N_8477,N_8428);
nor U8732 (N_8732,N_8442,N_8257);
and U8733 (N_8733,N_8363,N_8495);
xor U8734 (N_8734,N_8361,N_8497);
nor U8735 (N_8735,N_8419,N_8264);
nand U8736 (N_8736,N_8358,N_8471);
or U8737 (N_8737,N_8351,N_8480);
and U8738 (N_8738,N_8319,N_8465);
and U8739 (N_8739,N_8348,N_8460);
and U8740 (N_8740,N_8309,N_8396);
nor U8741 (N_8741,N_8255,N_8346);
and U8742 (N_8742,N_8344,N_8370);
and U8743 (N_8743,N_8418,N_8497);
nor U8744 (N_8744,N_8289,N_8426);
nand U8745 (N_8745,N_8496,N_8384);
or U8746 (N_8746,N_8487,N_8291);
and U8747 (N_8747,N_8334,N_8298);
nor U8748 (N_8748,N_8358,N_8420);
xor U8749 (N_8749,N_8311,N_8321);
and U8750 (N_8750,N_8728,N_8589);
xnor U8751 (N_8751,N_8542,N_8659);
nor U8752 (N_8752,N_8572,N_8606);
nor U8753 (N_8753,N_8534,N_8617);
and U8754 (N_8754,N_8510,N_8502);
or U8755 (N_8755,N_8550,N_8641);
and U8756 (N_8756,N_8601,N_8532);
nand U8757 (N_8757,N_8573,N_8503);
nand U8758 (N_8758,N_8707,N_8729);
or U8759 (N_8759,N_8675,N_8539);
or U8760 (N_8760,N_8545,N_8747);
and U8761 (N_8761,N_8664,N_8613);
nand U8762 (N_8762,N_8555,N_8543);
and U8763 (N_8763,N_8714,N_8533);
or U8764 (N_8764,N_8538,N_8552);
nand U8765 (N_8765,N_8528,N_8662);
and U8766 (N_8766,N_8665,N_8612);
nand U8767 (N_8767,N_8748,N_8574);
xnor U8768 (N_8768,N_8576,N_8727);
nor U8769 (N_8769,N_8703,N_8632);
or U8770 (N_8770,N_8704,N_8581);
nor U8771 (N_8771,N_8577,N_8663);
nor U8772 (N_8772,N_8607,N_8715);
or U8773 (N_8773,N_8518,N_8609);
and U8774 (N_8774,N_8520,N_8526);
nand U8775 (N_8775,N_8745,N_8620);
nand U8776 (N_8776,N_8652,N_8513);
and U8777 (N_8777,N_8621,N_8599);
and U8778 (N_8778,N_8509,N_8567);
and U8779 (N_8779,N_8692,N_8683);
or U8780 (N_8780,N_8564,N_8674);
or U8781 (N_8781,N_8725,N_8682);
nand U8782 (N_8782,N_8535,N_8708);
nand U8783 (N_8783,N_8690,N_8597);
xor U8784 (N_8784,N_8684,N_8546);
nor U8785 (N_8785,N_8596,N_8541);
or U8786 (N_8786,N_8643,N_8590);
nand U8787 (N_8787,N_8669,N_8501);
nand U8788 (N_8788,N_8701,N_8516);
and U8789 (N_8789,N_8673,N_8580);
or U8790 (N_8790,N_8644,N_8651);
and U8791 (N_8791,N_8689,N_8647);
nand U8792 (N_8792,N_8626,N_8640);
or U8793 (N_8793,N_8578,N_8676);
or U8794 (N_8794,N_8653,N_8511);
nand U8795 (N_8795,N_8508,N_8547);
or U8796 (N_8796,N_8672,N_8570);
nand U8797 (N_8797,N_8549,N_8721);
and U8798 (N_8798,N_8575,N_8744);
or U8799 (N_8799,N_8554,N_8595);
xnor U8800 (N_8800,N_8681,N_8678);
nand U8801 (N_8801,N_8749,N_8566);
nor U8802 (N_8802,N_8529,N_8565);
or U8803 (N_8803,N_8537,N_8639);
nand U8804 (N_8804,N_8583,N_8646);
and U8805 (N_8805,N_8695,N_8624);
nand U8806 (N_8806,N_8666,N_8702);
and U8807 (N_8807,N_8638,N_8521);
and U8808 (N_8808,N_8585,N_8522);
or U8809 (N_8809,N_8615,N_8584);
or U8810 (N_8810,N_8658,N_8634);
and U8811 (N_8811,N_8507,N_8723);
nor U8812 (N_8812,N_8616,N_8515);
nand U8813 (N_8813,N_8593,N_8604);
nand U8814 (N_8814,N_8712,N_8530);
nor U8815 (N_8815,N_8568,N_8504);
or U8816 (N_8816,N_8586,N_8711);
nand U8817 (N_8817,N_8741,N_8654);
nand U8818 (N_8818,N_8591,N_8614);
nor U8819 (N_8819,N_8694,N_8734);
xnor U8820 (N_8820,N_8735,N_8619);
xor U8821 (N_8821,N_8661,N_8719);
xnor U8822 (N_8822,N_8602,N_8710);
nor U8823 (N_8823,N_8540,N_8740);
nand U8824 (N_8824,N_8582,N_8699);
nor U8825 (N_8825,N_8667,N_8720);
nand U8826 (N_8826,N_8563,N_8743);
and U8827 (N_8827,N_8608,N_8730);
xor U8828 (N_8828,N_8649,N_8600);
xor U8829 (N_8829,N_8677,N_8746);
or U8830 (N_8830,N_8500,N_8642);
or U8831 (N_8831,N_8645,N_8679);
xnor U8832 (N_8832,N_8569,N_8519);
or U8833 (N_8833,N_8685,N_8724);
nand U8834 (N_8834,N_8698,N_8603);
and U8835 (N_8835,N_8622,N_8737);
nand U8836 (N_8836,N_8717,N_8731);
nor U8837 (N_8837,N_8742,N_8705);
or U8838 (N_8838,N_8637,N_8630);
xnor U8839 (N_8839,N_8610,N_8631);
and U8840 (N_8840,N_8633,N_8571);
or U8841 (N_8841,N_8732,N_8700);
and U8842 (N_8842,N_8693,N_8579);
xnor U8843 (N_8843,N_8588,N_8514);
nand U8844 (N_8844,N_8709,N_8660);
and U8845 (N_8845,N_8636,N_8655);
and U8846 (N_8846,N_8536,N_8611);
xor U8847 (N_8847,N_8629,N_8505);
or U8848 (N_8848,N_8512,N_8562);
and U8849 (N_8849,N_8718,N_8592);
xnor U8850 (N_8850,N_8524,N_8713);
nand U8851 (N_8851,N_8648,N_8671);
and U8852 (N_8852,N_8650,N_8517);
or U8853 (N_8853,N_8527,N_8697);
or U8854 (N_8854,N_8551,N_8668);
and U8855 (N_8855,N_8739,N_8680);
nand U8856 (N_8856,N_8687,N_8587);
or U8857 (N_8857,N_8553,N_8598);
and U8858 (N_8858,N_8531,N_8696);
and U8859 (N_8859,N_8544,N_8722);
and U8860 (N_8860,N_8618,N_8560);
and U8861 (N_8861,N_8605,N_8594);
and U8862 (N_8862,N_8628,N_8635);
and U8863 (N_8863,N_8716,N_8726);
nand U8864 (N_8864,N_8733,N_8548);
nor U8865 (N_8865,N_8738,N_8623);
nor U8866 (N_8866,N_8561,N_8523);
nand U8867 (N_8867,N_8625,N_8736);
or U8868 (N_8868,N_8558,N_8691);
or U8869 (N_8869,N_8656,N_8506);
nor U8870 (N_8870,N_8557,N_8657);
nor U8871 (N_8871,N_8525,N_8556);
and U8872 (N_8872,N_8559,N_8706);
nor U8873 (N_8873,N_8627,N_8686);
and U8874 (N_8874,N_8670,N_8688);
or U8875 (N_8875,N_8512,N_8574);
nand U8876 (N_8876,N_8722,N_8676);
and U8877 (N_8877,N_8616,N_8635);
nor U8878 (N_8878,N_8632,N_8604);
nor U8879 (N_8879,N_8521,N_8574);
nand U8880 (N_8880,N_8628,N_8639);
and U8881 (N_8881,N_8609,N_8595);
nor U8882 (N_8882,N_8560,N_8574);
or U8883 (N_8883,N_8599,N_8530);
and U8884 (N_8884,N_8740,N_8621);
or U8885 (N_8885,N_8534,N_8694);
xnor U8886 (N_8886,N_8520,N_8523);
nor U8887 (N_8887,N_8715,N_8666);
or U8888 (N_8888,N_8549,N_8672);
and U8889 (N_8889,N_8559,N_8733);
and U8890 (N_8890,N_8615,N_8511);
nand U8891 (N_8891,N_8688,N_8517);
or U8892 (N_8892,N_8660,N_8580);
or U8893 (N_8893,N_8532,N_8724);
xor U8894 (N_8894,N_8700,N_8567);
or U8895 (N_8895,N_8690,N_8566);
and U8896 (N_8896,N_8613,N_8693);
and U8897 (N_8897,N_8720,N_8544);
or U8898 (N_8898,N_8684,N_8518);
or U8899 (N_8899,N_8672,N_8685);
nand U8900 (N_8900,N_8575,N_8740);
or U8901 (N_8901,N_8544,N_8599);
or U8902 (N_8902,N_8505,N_8613);
nor U8903 (N_8903,N_8598,N_8676);
nor U8904 (N_8904,N_8721,N_8556);
xor U8905 (N_8905,N_8609,N_8526);
and U8906 (N_8906,N_8660,N_8516);
xor U8907 (N_8907,N_8573,N_8535);
xor U8908 (N_8908,N_8549,N_8722);
nor U8909 (N_8909,N_8686,N_8518);
nor U8910 (N_8910,N_8748,N_8704);
or U8911 (N_8911,N_8682,N_8579);
xnor U8912 (N_8912,N_8582,N_8604);
nor U8913 (N_8913,N_8624,N_8664);
nor U8914 (N_8914,N_8699,N_8511);
and U8915 (N_8915,N_8687,N_8717);
or U8916 (N_8916,N_8514,N_8562);
or U8917 (N_8917,N_8727,N_8639);
and U8918 (N_8918,N_8645,N_8575);
or U8919 (N_8919,N_8705,N_8736);
or U8920 (N_8920,N_8506,N_8617);
or U8921 (N_8921,N_8695,N_8566);
or U8922 (N_8922,N_8568,N_8613);
nor U8923 (N_8923,N_8647,N_8509);
or U8924 (N_8924,N_8536,N_8659);
or U8925 (N_8925,N_8540,N_8560);
and U8926 (N_8926,N_8539,N_8565);
or U8927 (N_8927,N_8685,N_8625);
or U8928 (N_8928,N_8634,N_8717);
nor U8929 (N_8929,N_8680,N_8692);
or U8930 (N_8930,N_8676,N_8631);
nand U8931 (N_8931,N_8695,N_8510);
and U8932 (N_8932,N_8567,N_8562);
xor U8933 (N_8933,N_8743,N_8649);
nor U8934 (N_8934,N_8524,N_8522);
nand U8935 (N_8935,N_8528,N_8610);
or U8936 (N_8936,N_8695,N_8674);
and U8937 (N_8937,N_8559,N_8676);
nor U8938 (N_8938,N_8511,N_8625);
nor U8939 (N_8939,N_8572,N_8711);
and U8940 (N_8940,N_8548,N_8723);
xnor U8941 (N_8941,N_8689,N_8579);
nor U8942 (N_8942,N_8516,N_8537);
nand U8943 (N_8943,N_8732,N_8606);
xor U8944 (N_8944,N_8595,N_8598);
nor U8945 (N_8945,N_8690,N_8729);
and U8946 (N_8946,N_8646,N_8544);
and U8947 (N_8947,N_8590,N_8511);
nand U8948 (N_8948,N_8731,N_8700);
nand U8949 (N_8949,N_8560,N_8676);
nand U8950 (N_8950,N_8501,N_8667);
xor U8951 (N_8951,N_8726,N_8681);
nand U8952 (N_8952,N_8675,N_8746);
nor U8953 (N_8953,N_8572,N_8696);
nand U8954 (N_8954,N_8728,N_8577);
nor U8955 (N_8955,N_8624,N_8515);
or U8956 (N_8956,N_8614,N_8711);
nand U8957 (N_8957,N_8724,N_8636);
and U8958 (N_8958,N_8571,N_8606);
nor U8959 (N_8959,N_8593,N_8587);
or U8960 (N_8960,N_8567,N_8593);
or U8961 (N_8961,N_8709,N_8687);
nand U8962 (N_8962,N_8515,N_8744);
nand U8963 (N_8963,N_8658,N_8682);
nor U8964 (N_8964,N_8703,N_8609);
or U8965 (N_8965,N_8574,N_8581);
xnor U8966 (N_8966,N_8559,N_8688);
nor U8967 (N_8967,N_8652,N_8624);
nand U8968 (N_8968,N_8632,N_8658);
nor U8969 (N_8969,N_8553,N_8534);
xor U8970 (N_8970,N_8596,N_8560);
nand U8971 (N_8971,N_8614,N_8559);
and U8972 (N_8972,N_8718,N_8571);
nand U8973 (N_8973,N_8719,N_8678);
nand U8974 (N_8974,N_8675,N_8613);
and U8975 (N_8975,N_8589,N_8662);
or U8976 (N_8976,N_8668,N_8534);
xor U8977 (N_8977,N_8572,N_8513);
nand U8978 (N_8978,N_8552,N_8723);
or U8979 (N_8979,N_8568,N_8692);
or U8980 (N_8980,N_8542,N_8666);
nand U8981 (N_8981,N_8691,N_8584);
nand U8982 (N_8982,N_8581,N_8691);
nand U8983 (N_8983,N_8741,N_8608);
nand U8984 (N_8984,N_8521,N_8547);
and U8985 (N_8985,N_8654,N_8664);
nand U8986 (N_8986,N_8551,N_8517);
nand U8987 (N_8987,N_8650,N_8550);
xnor U8988 (N_8988,N_8694,N_8591);
nor U8989 (N_8989,N_8583,N_8735);
nand U8990 (N_8990,N_8729,N_8689);
and U8991 (N_8991,N_8703,N_8659);
nor U8992 (N_8992,N_8686,N_8521);
nand U8993 (N_8993,N_8628,N_8659);
nand U8994 (N_8994,N_8709,N_8671);
nor U8995 (N_8995,N_8660,N_8612);
nand U8996 (N_8996,N_8516,N_8655);
and U8997 (N_8997,N_8598,N_8735);
nand U8998 (N_8998,N_8572,N_8553);
nor U8999 (N_8999,N_8501,N_8747);
and U9000 (N_9000,N_8882,N_8926);
nor U9001 (N_9001,N_8862,N_8764);
nor U9002 (N_9002,N_8788,N_8911);
nand U9003 (N_9003,N_8786,N_8797);
and U9004 (N_9004,N_8816,N_8991);
nand U9005 (N_9005,N_8768,N_8906);
or U9006 (N_9006,N_8978,N_8879);
or U9007 (N_9007,N_8957,N_8893);
or U9008 (N_9008,N_8888,N_8806);
or U9009 (N_9009,N_8783,N_8887);
or U9010 (N_9010,N_8897,N_8808);
or U9011 (N_9011,N_8946,N_8892);
and U9012 (N_9012,N_8932,N_8803);
nor U9013 (N_9013,N_8880,N_8940);
or U9014 (N_9014,N_8799,N_8853);
or U9015 (N_9015,N_8979,N_8918);
xor U9016 (N_9016,N_8999,N_8779);
or U9017 (N_9017,N_8908,N_8765);
and U9018 (N_9018,N_8876,N_8949);
nor U9019 (N_9019,N_8867,N_8998);
or U9020 (N_9020,N_8935,N_8873);
nor U9021 (N_9021,N_8841,N_8915);
or U9022 (N_9022,N_8755,N_8798);
and U9023 (N_9023,N_8973,N_8762);
or U9024 (N_9024,N_8829,N_8849);
nor U9025 (N_9025,N_8937,N_8759);
or U9026 (N_9026,N_8811,N_8854);
and U9027 (N_9027,N_8848,N_8913);
or U9028 (N_9028,N_8965,N_8992);
or U9029 (N_9029,N_8758,N_8775);
nand U9030 (N_9030,N_8845,N_8948);
nand U9031 (N_9031,N_8967,N_8781);
or U9032 (N_9032,N_8802,N_8776);
nand U9033 (N_9033,N_8969,N_8984);
nand U9034 (N_9034,N_8910,N_8761);
nand U9035 (N_9035,N_8941,N_8903);
xor U9036 (N_9036,N_8832,N_8934);
or U9037 (N_9037,N_8981,N_8960);
nor U9038 (N_9038,N_8931,N_8977);
and U9039 (N_9039,N_8942,N_8846);
nor U9040 (N_9040,N_8835,N_8902);
and U9041 (N_9041,N_8975,N_8817);
nand U9042 (N_9042,N_8820,N_8877);
nor U9043 (N_9043,N_8985,N_8919);
nand U9044 (N_9044,N_8883,N_8958);
nand U9045 (N_9045,N_8971,N_8885);
nor U9046 (N_9046,N_8815,N_8800);
and U9047 (N_9047,N_8968,N_8970);
or U9048 (N_9048,N_8870,N_8990);
nand U9049 (N_9049,N_8756,N_8881);
nand U9050 (N_9050,N_8872,N_8807);
nand U9051 (N_9051,N_8914,N_8860);
nand U9052 (N_9052,N_8976,N_8950);
and U9053 (N_9053,N_8834,N_8777);
nand U9054 (N_9054,N_8947,N_8994);
or U9055 (N_9055,N_8851,N_8789);
and U9056 (N_9056,N_8982,N_8901);
and U9057 (N_9057,N_8943,N_8997);
nand U9058 (N_9058,N_8858,N_8920);
nand U9059 (N_9059,N_8900,N_8836);
and U9060 (N_9060,N_8780,N_8813);
nor U9061 (N_9061,N_8961,N_8766);
or U9062 (N_9062,N_8884,N_8929);
nor U9063 (N_9063,N_8890,N_8927);
and U9064 (N_9064,N_8814,N_8855);
or U9065 (N_9065,N_8784,N_8963);
nor U9066 (N_9066,N_8822,N_8857);
or U9067 (N_9067,N_8837,N_8778);
nor U9068 (N_9068,N_8819,N_8863);
nor U9069 (N_9069,N_8757,N_8933);
and U9070 (N_9070,N_8763,N_8894);
nor U9071 (N_9071,N_8945,N_8878);
xnor U9072 (N_9072,N_8905,N_8773);
and U9073 (N_9073,N_8767,N_8869);
or U9074 (N_9074,N_8787,N_8843);
nand U9075 (N_9075,N_8791,N_8987);
nor U9076 (N_9076,N_8750,N_8962);
or U9077 (N_9077,N_8801,N_8922);
nand U9078 (N_9078,N_8966,N_8923);
xor U9079 (N_9079,N_8793,N_8988);
or U9080 (N_9080,N_8753,N_8907);
or U9081 (N_9081,N_8833,N_8859);
nand U9082 (N_9082,N_8871,N_8864);
xor U9083 (N_9083,N_8842,N_8930);
nand U9084 (N_9084,N_8754,N_8794);
and U9085 (N_9085,N_8792,N_8782);
nand U9086 (N_9086,N_8856,N_8956);
nor U9087 (N_9087,N_8917,N_8840);
or U9088 (N_9088,N_8861,N_8895);
nor U9089 (N_9089,N_8760,N_8986);
nor U9090 (N_9090,N_8838,N_8874);
nand U9091 (N_9091,N_8824,N_8959);
nand U9092 (N_9092,N_8810,N_8850);
nor U9093 (N_9093,N_8974,N_8996);
nand U9094 (N_9094,N_8852,N_8912);
and U9095 (N_9095,N_8774,N_8939);
or U9096 (N_9096,N_8951,N_8827);
or U9097 (N_9097,N_8790,N_8989);
or U9098 (N_9098,N_8771,N_8889);
xor U9099 (N_9099,N_8875,N_8818);
and U9100 (N_9100,N_8954,N_8795);
nor U9101 (N_9101,N_8830,N_8886);
and U9102 (N_9102,N_8936,N_8839);
and U9103 (N_9103,N_8825,N_8891);
or U9104 (N_9104,N_8925,N_8921);
or U9105 (N_9105,N_8924,N_8831);
and U9106 (N_9106,N_8823,N_8983);
nor U9107 (N_9107,N_8866,N_8898);
nor U9108 (N_9108,N_8972,N_8896);
nor U9109 (N_9109,N_8955,N_8769);
nor U9110 (N_9110,N_8944,N_8909);
and U9111 (N_9111,N_8938,N_8928);
and U9112 (N_9112,N_8916,N_8796);
and U9113 (N_9113,N_8953,N_8904);
and U9114 (N_9114,N_8821,N_8770);
or U9115 (N_9115,N_8952,N_8847);
nor U9116 (N_9116,N_8993,N_8804);
nor U9117 (N_9117,N_8980,N_8899);
nand U9118 (N_9118,N_8812,N_8785);
and U9119 (N_9119,N_8964,N_8772);
nand U9120 (N_9120,N_8868,N_8805);
and U9121 (N_9121,N_8995,N_8828);
and U9122 (N_9122,N_8826,N_8752);
or U9123 (N_9123,N_8809,N_8751);
nor U9124 (N_9124,N_8844,N_8865);
and U9125 (N_9125,N_8815,N_8982);
and U9126 (N_9126,N_8947,N_8797);
or U9127 (N_9127,N_8833,N_8967);
nor U9128 (N_9128,N_8889,N_8762);
nand U9129 (N_9129,N_8915,N_8866);
nor U9130 (N_9130,N_8914,N_8979);
nand U9131 (N_9131,N_8848,N_8987);
xor U9132 (N_9132,N_8817,N_8762);
or U9133 (N_9133,N_8872,N_8829);
nor U9134 (N_9134,N_8898,N_8852);
or U9135 (N_9135,N_8857,N_8826);
xor U9136 (N_9136,N_8767,N_8896);
or U9137 (N_9137,N_8791,N_8814);
nor U9138 (N_9138,N_8893,N_8785);
and U9139 (N_9139,N_8902,N_8855);
and U9140 (N_9140,N_8761,N_8819);
or U9141 (N_9141,N_8817,N_8802);
or U9142 (N_9142,N_8918,N_8889);
and U9143 (N_9143,N_8907,N_8794);
nand U9144 (N_9144,N_8945,N_8754);
and U9145 (N_9145,N_8923,N_8989);
nand U9146 (N_9146,N_8897,N_8826);
nand U9147 (N_9147,N_8987,N_8766);
or U9148 (N_9148,N_8819,N_8827);
or U9149 (N_9149,N_8901,N_8923);
nand U9150 (N_9150,N_8759,N_8774);
nor U9151 (N_9151,N_8948,N_8968);
and U9152 (N_9152,N_8987,N_8820);
nor U9153 (N_9153,N_8878,N_8983);
nand U9154 (N_9154,N_8798,N_8914);
and U9155 (N_9155,N_8822,N_8769);
or U9156 (N_9156,N_8794,N_8886);
nor U9157 (N_9157,N_8790,N_8969);
xor U9158 (N_9158,N_8856,N_8929);
xor U9159 (N_9159,N_8790,N_8776);
nor U9160 (N_9160,N_8924,N_8921);
nand U9161 (N_9161,N_8797,N_8983);
nor U9162 (N_9162,N_8996,N_8804);
and U9163 (N_9163,N_8795,N_8761);
or U9164 (N_9164,N_8773,N_8783);
nand U9165 (N_9165,N_8946,N_8873);
nand U9166 (N_9166,N_8763,N_8755);
xnor U9167 (N_9167,N_8977,N_8767);
or U9168 (N_9168,N_8922,N_8873);
and U9169 (N_9169,N_8767,N_8910);
or U9170 (N_9170,N_8982,N_8804);
and U9171 (N_9171,N_8944,N_8953);
and U9172 (N_9172,N_8961,N_8814);
nor U9173 (N_9173,N_8774,N_8905);
and U9174 (N_9174,N_8864,N_8999);
nand U9175 (N_9175,N_8877,N_8910);
nor U9176 (N_9176,N_8966,N_8784);
nor U9177 (N_9177,N_8845,N_8764);
nor U9178 (N_9178,N_8789,N_8938);
nor U9179 (N_9179,N_8776,N_8966);
and U9180 (N_9180,N_8954,N_8799);
nor U9181 (N_9181,N_8782,N_8837);
nand U9182 (N_9182,N_8917,N_8969);
nand U9183 (N_9183,N_8794,N_8818);
or U9184 (N_9184,N_8967,N_8925);
nand U9185 (N_9185,N_8871,N_8771);
or U9186 (N_9186,N_8944,N_8813);
or U9187 (N_9187,N_8969,N_8934);
nand U9188 (N_9188,N_8932,N_8848);
or U9189 (N_9189,N_8891,N_8805);
or U9190 (N_9190,N_8947,N_8823);
or U9191 (N_9191,N_8922,N_8913);
nor U9192 (N_9192,N_8970,N_8791);
or U9193 (N_9193,N_8755,N_8905);
or U9194 (N_9194,N_8882,N_8776);
and U9195 (N_9195,N_8872,N_8990);
nor U9196 (N_9196,N_8955,N_8993);
nor U9197 (N_9197,N_8800,N_8927);
or U9198 (N_9198,N_8767,N_8828);
nor U9199 (N_9199,N_8896,N_8887);
nor U9200 (N_9200,N_8786,N_8917);
or U9201 (N_9201,N_8914,N_8955);
xor U9202 (N_9202,N_8988,N_8944);
nand U9203 (N_9203,N_8818,N_8979);
nand U9204 (N_9204,N_8877,N_8925);
nand U9205 (N_9205,N_8812,N_8909);
and U9206 (N_9206,N_8909,N_8793);
nand U9207 (N_9207,N_8775,N_8986);
or U9208 (N_9208,N_8789,N_8927);
and U9209 (N_9209,N_8766,N_8863);
xor U9210 (N_9210,N_8923,N_8956);
nand U9211 (N_9211,N_8954,N_8925);
or U9212 (N_9212,N_8897,N_8964);
nor U9213 (N_9213,N_8833,N_8916);
and U9214 (N_9214,N_8909,N_8946);
and U9215 (N_9215,N_8800,N_8921);
xnor U9216 (N_9216,N_8798,N_8856);
xnor U9217 (N_9217,N_8819,N_8766);
nand U9218 (N_9218,N_8832,N_8846);
nor U9219 (N_9219,N_8815,N_8775);
and U9220 (N_9220,N_8855,N_8907);
nand U9221 (N_9221,N_8786,N_8772);
nand U9222 (N_9222,N_8780,N_8897);
or U9223 (N_9223,N_8972,N_8784);
xor U9224 (N_9224,N_8990,N_8987);
nor U9225 (N_9225,N_8937,N_8754);
nor U9226 (N_9226,N_8955,N_8808);
xor U9227 (N_9227,N_8805,N_8869);
xnor U9228 (N_9228,N_8850,N_8811);
or U9229 (N_9229,N_8858,N_8967);
nand U9230 (N_9230,N_8882,N_8851);
and U9231 (N_9231,N_8953,N_8799);
nor U9232 (N_9232,N_8788,N_8888);
nor U9233 (N_9233,N_8825,N_8982);
nor U9234 (N_9234,N_8823,N_8871);
nor U9235 (N_9235,N_8995,N_8886);
or U9236 (N_9236,N_8776,N_8890);
nand U9237 (N_9237,N_8874,N_8787);
and U9238 (N_9238,N_8829,N_8864);
and U9239 (N_9239,N_8856,N_8881);
nor U9240 (N_9240,N_8954,N_8872);
nand U9241 (N_9241,N_8842,N_8992);
nor U9242 (N_9242,N_8871,N_8867);
or U9243 (N_9243,N_8927,N_8980);
nand U9244 (N_9244,N_8899,N_8818);
or U9245 (N_9245,N_8914,N_8977);
nor U9246 (N_9246,N_8939,N_8841);
or U9247 (N_9247,N_8911,N_8913);
xnor U9248 (N_9248,N_8847,N_8964);
nor U9249 (N_9249,N_8869,N_8876);
or U9250 (N_9250,N_9192,N_9019);
and U9251 (N_9251,N_9138,N_9221);
or U9252 (N_9252,N_9238,N_9112);
nand U9253 (N_9253,N_9126,N_9193);
and U9254 (N_9254,N_9158,N_9081);
nand U9255 (N_9255,N_9218,N_9045);
or U9256 (N_9256,N_9249,N_9055);
nand U9257 (N_9257,N_9016,N_9197);
nor U9258 (N_9258,N_9135,N_9005);
nand U9259 (N_9259,N_9109,N_9181);
nor U9260 (N_9260,N_9242,N_9151);
nor U9261 (N_9261,N_9006,N_9104);
or U9262 (N_9262,N_9134,N_9056);
nor U9263 (N_9263,N_9233,N_9062);
nand U9264 (N_9264,N_9153,N_9133);
nor U9265 (N_9265,N_9227,N_9030);
nor U9266 (N_9266,N_9003,N_9129);
nor U9267 (N_9267,N_9149,N_9049);
nand U9268 (N_9268,N_9243,N_9127);
or U9269 (N_9269,N_9080,N_9219);
nand U9270 (N_9270,N_9156,N_9119);
and U9271 (N_9271,N_9234,N_9107);
nor U9272 (N_9272,N_9189,N_9008);
and U9273 (N_9273,N_9177,N_9165);
or U9274 (N_9274,N_9090,N_9122);
and U9275 (N_9275,N_9145,N_9222);
nand U9276 (N_9276,N_9076,N_9067);
and U9277 (N_9277,N_9196,N_9247);
xor U9278 (N_9278,N_9236,N_9210);
nand U9279 (N_9279,N_9182,N_9185);
or U9280 (N_9280,N_9211,N_9052);
nand U9281 (N_9281,N_9002,N_9229);
and U9282 (N_9282,N_9170,N_9139);
or U9283 (N_9283,N_9072,N_9029);
nor U9284 (N_9284,N_9143,N_9036);
and U9285 (N_9285,N_9168,N_9136);
or U9286 (N_9286,N_9075,N_9140);
xnor U9287 (N_9287,N_9022,N_9183);
nand U9288 (N_9288,N_9161,N_9026);
nand U9289 (N_9289,N_9191,N_9204);
or U9290 (N_9290,N_9059,N_9050);
and U9291 (N_9291,N_9113,N_9132);
nor U9292 (N_9292,N_9128,N_9144);
nor U9293 (N_9293,N_9244,N_9024);
and U9294 (N_9294,N_9190,N_9154);
nor U9295 (N_9295,N_9028,N_9150);
or U9296 (N_9296,N_9043,N_9093);
and U9297 (N_9297,N_9035,N_9065);
or U9298 (N_9298,N_9096,N_9082);
xor U9299 (N_9299,N_9091,N_9098);
or U9300 (N_9300,N_9087,N_9245);
nor U9301 (N_9301,N_9173,N_9180);
xnor U9302 (N_9302,N_9051,N_9004);
or U9303 (N_9303,N_9225,N_9032);
nand U9304 (N_9304,N_9202,N_9012);
nor U9305 (N_9305,N_9097,N_9027);
xnor U9306 (N_9306,N_9231,N_9176);
and U9307 (N_9307,N_9048,N_9105);
xor U9308 (N_9308,N_9103,N_9201);
or U9309 (N_9309,N_9046,N_9009);
or U9310 (N_9310,N_9007,N_9246);
and U9311 (N_9311,N_9169,N_9131);
nor U9312 (N_9312,N_9092,N_9198);
nand U9313 (N_9313,N_9042,N_9146);
and U9314 (N_9314,N_9040,N_9175);
and U9315 (N_9315,N_9141,N_9205);
or U9316 (N_9316,N_9148,N_9017);
nand U9317 (N_9317,N_9239,N_9157);
nand U9318 (N_9318,N_9118,N_9155);
nand U9319 (N_9319,N_9071,N_9213);
and U9320 (N_9320,N_9166,N_9115);
or U9321 (N_9321,N_9014,N_9088);
or U9322 (N_9322,N_9130,N_9047);
nor U9323 (N_9323,N_9164,N_9240);
or U9324 (N_9324,N_9174,N_9171);
and U9325 (N_9325,N_9203,N_9064);
and U9326 (N_9326,N_9108,N_9207);
nand U9327 (N_9327,N_9111,N_9089);
nand U9328 (N_9328,N_9068,N_9167);
nand U9329 (N_9329,N_9085,N_9011);
nor U9330 (N_9330,N_9025,N_9106);
and U9331 (N_9331,N_9208,N_9015);
nor U9332 (N_9332,N_9124,N_9001);
nand U9333 (N_9333,N_9194,N_9101);
or U9334 (N_9334,N_9241,N_9023);
nand U9335 (N_9335,N_9121,N_9228);
or U9336 (N_9336,N_9053,N_9230);
nor U9337 (N_9337,N_9078,N_9074);
or U9338 (N_9338,N_9215,N_9084);
or U9339 (N_9339,N_9069,N_9248);
nor U9340 (N_9340,N_9010,N_9125);
or U9341 (N_9341,N_9066,N_9123);
or U9342 (N_9342,N_9034,N_9120);
or U9343 (N_9343,N_9061,N_9060);
nand U9344 (N_9344,N_9083,N_9058);
or U9345 (N_9345,N_9044,N_9147);
or U9346 (N_9346,N_9209,N_9226);
xor U9347 (N_9347,N_9162,N_9033);
and U9348 (N_9348,N_9079,N_9013);
nor U9349 (N_9349,N_9195,N_9159);
xor U9350 (N_9350,N_9172,N_9224);
nand U9351 (N_9351,N_9094,N_9160);
nor U9352 (N_9352,N_9152,N_9200);
or U9353 (N_9353,N_9163,N_9038);
and U9354 (N_9354,N_9178,N_9095);
and U9355 (N_9355,N_9188,N_9018);
and U9356 (N_9356,N_9186,N_9031);
or U9357 (N_9357,N_9137,N_9114);
nand U9358 (N_9358,N_9217,N_9020);
and U9359 (N_9359,N_9086,N_9179);
or U9360 (N_9360,N_9214,N_9077);
nor U9361 (N_9361,N_9212,N_9057);
nand U9362 (N_9362,N_9021,N_9073);
and U9363 (N_9363,N_9102,N_9184);
or U9364 (N_9364,N_9063,N_9206);
and U9365 (N_9365,N_9235,N_9000);
and U9366 (N_9366,N_9223,N_9070);
xor U9367 (N_9367,N_9110,N_9232);
and U9368 (N_9368,N_9187,N_9199);
xor U9369 (N_9369,N_9117,N_9099);
xnor U9370 (N_9370,N_9039,N_9100);
or U9371 (N_9371,N_9116,N_9054);
nand U9372 (N_9372,N_9237,N_9037);
nand U9373 (N_9373,N_9220,N_9216);
or U9374 (N_9374,N_9041,N_9142);
xnor U9375 (N_9375,N_9142,N_9046);
nand U9376 (N_9376,N_9051,N_9077);
and U9377 (N_9377,N_9230,N_9003);
and U9378 (N_9378,N_9191,N_9223);
and U9379 (N_9379,N_9217,N_9154);
or U9380 (N_9380,N_9224,N_9188);
or U9381 (N_9381,N_9016,N_9186);
xor U9382 (N_9382,N_9216,N_9013);
or U9383 (N_9383,N_9126,N_9163);
nor U9384 (N_9384,N_9178,N_9114);
and U9385 (N_9385,N_9167,N_9218);
nor U9386 (N_9386,N_9158,N_9146);
nand U9387 (N_9387,N_9196,N_9098);
or U9388 (N_9388,N_9219,N_9051);
nor U9389 (N_9389,N_9227,N_9096);
nand U9390 (N_9390,N_9126,N_9037);
nor U9391 (N_9391,N_9007,N_9185);
and U9392 (N_9392,N_9089,N_9185);
nor U9393 (N_9393,N_9166,N_9033);
or U9394 (N_9394,N_9138,N_9225);
nand U9395 (N_9395,N_9196,N_9242);
or U9396 (N_9396,N_9232,N_9210);
nor U9397 (N_9397,N_9152,N_9057);
nor U9398 (N_9398,N_9211,N_9010);
nand U9399 (N_9399,N_9134,N_9159);
nand U9400 (N_9400,N_9080,N_9023);
and U9401 (N_9401,N_9010,N_9100);
nand U9402 (N_9402,N_9000,N_9192);
and U9403 (N_9403,N_9108,N_9233);
nand U9404 (N_9404,N_9189,N_9073);
xor U9405 (N_9405,N_9014,N_9169);
or U9406 (N_9406,N_9158,N_9187);
nand U9407 (N_9407,N_9121,N_9041);
and U9408 (N_9408,N_9192,N_9023);
and U9409 (N_9409,N_9074,N_9115);
or U9410 (N_9410,N_9049,N_9208);
or U9411 (N_9411,N_9182,N_9096);
nand U9412 (N_9412,N_9055,N_9056);
or U9413 (N_9413,N_9146,N_9105);
nor U9414 (N_9414,N_9195,N_9249);
and U9415 (N_9415,N_9149,N_9071);
or U9416 (N_9416,N_9093,N_9117);
nand U9417 (N_9417,N_9134,N_9141);
nand U9418 (N_9418,N_9149,N_9219);
or U9419 (N_9419,N_9176,N_9047);
or U9420 (N_9420,N_9110,N_9107);
and U9421 (N_9421,N_9198,N_9117);
nor U9422 (N_9422,N_9022,N_9185);
and U9423 (N_9423,N_9220,N_9147);
and U9424 (N_9424,N_9115,N_9022);
and U9425 (N_9425,N_9003,N_9088);
nand U9426 (N_9426,N_9248,N_9087);
or U9427 (N_9427,N_9108,N_9100);
or U9428 (N_9428,N_9004,N_9102);
and U9429 (N_9429,N_9189,N_9089);
or U9430 (N_9430,N_9129,N_9038);
or U9431 (N_9431,N_9188,N_9001);
or U9432 (N_9432,N_9010,N_9044);
or U9433 (N_9433,N_9139,N_9001);
nor U9434 (N_9434,N_9172,N_9014);
xor U9435 (N_9435,N_9099,N_9055);
nor U9436 (N_9436,N_9148,N_9225);
nor U9437 (N_9437,N_9179,N_9234);
nor U9438 (N_9438,N_9020,N_9113);
nand U9439 (N_9439,N_9145,N_9242);
nand U9440 (N_9440,N_9098,N_9028);
nor U9441 (N_9441,N_9135,N_9020);
nor U9442 (N_9442,N_9049,N_9038);
and U9443 (N_9443,N_9030,N_9097);
nand U9444 (N_9444,N_9132,N_9168);
and U9445 (N_9445,N_9002,N_9108);
nor U9446 (N_9446,N_9040,N_9064);
xnor U9447 (N_9447,N_9148,N_9096);
nand U9448 (N_9448,N_9203,N_9105);
and U9449 (N_9449,N_9088,N_9209);
and U9450 (N_9450,N_9174,N_9050);
nand U9451 (N_9451,N_9245,N_9061);
nand U9452 (N_9452,N_9017,N_9166);
nand U9453 (N_9453,N_9207,N_9163);
nor U9454 (N_9454,N_9194,N_9009);
nand U9455 (N_9455,N_9089,N_9165);
and U9456 (N_9456,N_9233,N_9186);
nor U9457 (N_9457,N_9021,N_9120);
and U9458 (N_9458,N_9224,N_9122);
and U9459 (N_9459,N_9003,N_9241);
nand U9460 (N_9460,N_9045,N_9223);
or U9461 (N_9461,N_9182,N_9141);
nand U9462 (N_9462,N_9121,N_9243);
nor U9463 (N_9463,N_9108,N_9141);
nand U9464 (N_9464,N_9178,N_9228);
nand U9465 (N_9465,N_9138,N_9122);
nand U9466 (N_9466,N_9081,N_9127);
nand U9467 (N_9467,N_9083,N_9190);
nor U9468 (N_9468,N_9248,N_9064);
or U9469 (N_9469,N_9202,N_9007);
or U9470 (N_9470,N_9099,N_9035);
nand U9471 (N_9471,N_9033,N_9199);
xnor U9472 (N_9472,N_9243,N_9134);
or U9473 (N_9473,N_9052,N_9088);
nand U9474 (N_9474,N_9061,N_9031);
and U9475 (N_9475,N_9061,N_9095);
nor U9476 (N_9476,N_9128,N_9071);
or U9477 (N_9477,N_9021,N_9105);
and U9478 (N_9478,N_9182,N_9202);
nor U9479 (N_9479,N_9167,N_9217);
and U9480 (N_9480,N_9032,N_9159);
nand U9481 (N_9481,N_9098,N_9156);
nand U9482 (N_9482,N_9180,N_9016);
nor U9483 (N_9483,N_9123,N_9181);
nand U9484 (N_9484,N_9046,N_9041);
xor U9485 (N_9485,N_9176,N_9010);
and U9486 (N_9486,N_9184,N_9089);
nor U9487 (N_9487,N_9039,N_9085);
nand U9488 (N_9488,N_9230,N_9126);
and U9489 (N_9489,N_9024,N_9004);
nand U9490 (N_9490,N_9220,N_9187);
nor U9491 (N_9491,N_9039,N_9078);
xor U9492 (N_9492,N_9085,N_9022);
nor U9493 (N_9493,N_9081,N_9223);
nand U9494 (N_9494,N_9194,N_9124);
nor U9495 (N_9495,N_9134,N_9165);
nor U9496 (N_9496,N_9136,N_9231);
nor U9497 (N_9497,N_9095,N_9234);
nor U9498 (N_9498,N_9233,N_9092);
nor U9499 (N_9499,N_9020,N_9163);
nand U9500 (N_9500,N_9426,N_9331);
nand U9501 (N_9501,N_9414,N_9418);
or U9502 (N_9502,N_9473,N_9321);
or U9503 (N_9503,N_9481,N_9398);
nor U9504 (N_9504,N_9416,N_9468);
or U9505 (N_9505,N_9439,N_9265);
nand U9506 (N_9506,N_9374,N_9392);
nand U9507 (N_9507,N_9289,N_9371);
or U9508 (N_9508,N_9404,N_9269);
or U9509 (N_9509,N_9447,N_9272);
or U9510 (N_9510,N_9420,N_9460);
and U9511 (N_9511,N_9488,N_9299);
nand U9512 (N_9512,N_9471,N_9415);
nor U9513 (N_9513,N_9252,N_9406);
and U9514 (N_9514,N_9432,N_9445);
nand U9515 (N_9515,N_9405,N_9430);
and U9516 (N_9516,N_9437,N_9485);
nand U9517 (N_9517,N_9452,N_9345);
and U9518 (N_9518,N_9465,N_9346);
or U9519 (N_9519,N_9308,N_9311);
and U9520 (N_9520,N_9334,N_9441);
nor U9521 (N_9521,N_9467,N_9276);
nand U9522 (N_9522,N_9306,N_9261);
or U9523 (N_9523,N_9274,N_9360);
nand U9524 (N_9524,N_9435,N_9352);
nand U9525 (N_9525,N_9494,N_9425);
nand U9526 (N_9526,N_9409,N_9444);
nor U9527 (N_9527,N_9264,N_9387);
and U9528 (N_9528,N_9347,N_9429);
or U9529 (N_9529,N_9332,N_9277);
nand U9530 (N_9530,N_9377,N_9314);
xor U9531 (N_9531,N_9292,N_9280);
nor U9532 (N_9532,N_9367,N_9458);
and U9533 (N_9533,N_9260,N_9421);
and U9534 (N_9534,N_9351,N_9333);
and U9535 (N_9535,N_9325,N_9339);
xnor U9536 (N_9536,N_9318,N_9324);
nor U9537 (N_9537,N_9251,N_9283);
xnor U9538 (N_9538,N_9390,N_9375);
nor U9539 (N_9539,N_9407,N_9461);
nor U9540 (N_9540,N_9436,N_9419);
xnor U9541 (N_9541,N_9479,N_9486);
or U9542 (N_9542,N_9446,N_9361);
nand U9543 (N_9543,N_9357,N_9356);
and U9544 (N_9544,N_9271,N_9381);
or U9545 (N_9545,N_9344,N_9255);
and U9546 (N_9546,N_9484,N_9493);
nand U9547 (N_9547,N_9294,N_9329);
nor U9548 (N_9548,N_9362,N_9455);
nor U9549 (N_9549,N_9433,N_9456);
nor U9550 (N_9550,N_9376,N_9466);
nor U9551 (N_9551,N_9319,N_9423);
and U9552 (N_9552,N_9463,N_9499);
nand U9553 (N_9553,N_9474,N_9364);
or U9554 (N_9554,N_9335,N_9395);
or U9555 (N_9555,N_9396,N_9478);
nand U9556 (N_9556,N_9453,N_9301);
nand U9557 (N_9557,N_9316,N_9326);
nor U9558 (N_9558,N_9350,N_9354);
xor U9559 (N_9559,N_9498,N_9353);
or U9560 (N_9560,N_9393,N_9412);
and U9561 (N_9561,N_9476,N_9257);
xnor U9562 (N_9562,N_9328,N_9338);
nor U9563 (N_9563,N_9259,N_9400);
nand U9564 (N_9564,N_9372,N_9262);
and U9565 (N_9565,N_9451,N_9477);
and U9566 (N_9566,N_9285,N_9293);
or U9567 (N_9567,N_9380,N_9317);
nor U9568 (N_9568,N_9492,N_9284);
and U9569 (N_9569,N_9497,N_9442);
or U9570 (N_9570,N_9300,N_9263);
nand U9571 (N_9571,N_9279,N_9327);
and U9572 (N_9572,N_9403,N_9287);
and U9573 (N_9573,N_9417,N_9449);
xnor U9574 (N_9574,N_9295,N_9408);
and U9575 (N_9575,N_9266,N_9388);
nand U9576 (N_9576,N_9323,N_9472);
and U9577 (N_9577,N_9469,N_9315);
nor U9578 (N_9578,N_9342,N_9495);
and U9579 (N_9579,N_9373,N_9428);
xnor U9580 (N_9580,N_9491,N_9424);
nand U9581 (N_9581,N_9278,N_9330);
nor U9582 (N_9582,N_9394,N_9379);
nand U9583 (N_9583,N_9298,N_9378);
nor U9584 (N_9584,N_9440,N_9302);
nand U9585 (N_9585,N_9487,N_9427);
and U9586 (N_9586,N_9343,N_9312);
xnor U9587 (N_9587,N_9363,N_9391);
nand U9588 (N_9588,N_9422,N_9399);
and U9589 (N_9589,N_9434,N_9454);
nand U9590 (N_9590,N_9496,N_9267);
nand U9591 (N_9591,N_9349,N_9475);
nand U9592 (N_9592,N_9483,N_9450);
nor U9593 (N_9593,N_9309,N_9366);
nand U9594 (N_9594,N_9386,N_9305);
nor U9595 (N_9595,N_9480,N_9438);
nor U9596 (N_9596,N_9322,N_9402);
nor U9597 (N_9597,N_9355,N_9448);
or U9598 (N_9598,N_9250,N_9290);
nor U9599 (N_9599,N_9389,N_9268);
nor U9600 (N_9600,N_9273,N_9358);
nor U9601 (N_9601,N_9359,N_9482);
nand U9602 (N_9602,N_9270,N_9384);
nor U9603 (N_9603,N_9443,N_9303);
and U9604 (N_9604,N_9313,N_9457);
or U9605 (N_9605,N_9336,N_9459);
and U9606 (N_9606,N_9282,N_9431);
and U9607 (N_9607,N_9286,N_9411);
nor U9608 (N_9608,N_9410,N_9348);
xnor U9609 (N_9609,N_9291,N_9470);
and U9610 (N_9610,N_9275,N_9307);
or U9611 (N_9611,N_9365,N_9304);
nand U9612 (N_9612,N_9320,N_9490);
nor U9613 (N_9613,N_9489,N_9340);
and U9614 (N_9614,N_9341,N_9296);
nand U9615 (N_9615,N_9413,N_9337);
or U9616 (N_9616,N_9256,N_9385);
nor U9617 (N_9617,N_9288,N_9382);
nand U9618 (N_9618,N_9253,N_9281);
nor U9619 (N_9619,N_9383,N_9368);
or U9620 (N_9620,N_9401,N_9462);
xnor U9621 (N_9621,N_9370,N_9369);
or U9622 (N_9622,N_9397,N_9310);
nor U9623 (N_9623,N_9297,N_9464);
and U9624 (N_9624,N_9254,N_9258);
or U9625 (N_9625,N_9464,N_9438);
nor U9626 (N_9626,N_9303,N_9272);
nor U9627 (N_9627,N_9305,N_9451);
nand U9628 (N_9628,N_9383,N_9355);
and U9629 (N_9629,N_9449,N_9404);
and U9630 (N_9630,N_9487,N_9342);
nor U9631 (N_9631,N_9495,N_9391);
nand U9632 (N_9632,N_9293,N_9473);
or U9633 (N_9633,N_9300,N_9409);
or U9634 (N_9634,N_9486,N_9449);
and U9635 (N_9635,N_9315,N_9456);
and U9636 (N_9636,N_9408,N_9352);
nand U9637 (N_9637,N_9465,N_9488);
xor U9638 (N_9638,N_9297,N_9257);
nand U9639 (N_9639,N_9385,N_9265);
or U9640 (N_9640,N_9329,N_9477);
or U9641 (N_9641,N_9431,N_9409);
nand U9642 (N_9642,N_9390,N_9458);
nor U9643 (N_9643,N_9412,N_9407);
or U9644 (N_9644,N_9316,N_9413);
nor U9645 (N_9645,N_9251,N_9415);
or U9646 (N_9646,N_9424,N_9253);
nand U9647 (N_9647,N_9352,N_9338);
and U9648 (N_9648,N_9454,N_9420);
nand U9649 (N_9649,N_9460,N_9287);
nand U9650 (N_9650,N_9315,N_9379);
or U9651 (N_9651,N_9322,N_9347);
and U9652 (N_9652,N_9281,N_9364);
xnor U9653 (N_9653,N_9277,N_9335);
and U9654 (N_9654,N_9346,N_9476);
and U9655 (N_9655,N_9334,N_9461);
and U9656 (N_9656,N_9290,N_9377);
xor U9657 (N_9657,N_9391,N_9484);
or U9658 (N_9658,N_9491,N_9382);
nor U9659 (N_9659,N_9428,N_9266);
nand U9660 (N_9660,N_9451,N_9452);
or U9661 (N_9661,N_9346,N_9354);
xor U9662 (N_9662,N_9462,N_9396);
nor U9663 (N_9663,N_9290,N_9358);
and U9664 (N_9664,N_9435,N_9254);
xor U9665 (N_9665,N_9492,N_9314);
nor U9666 (N_9666,N_9344,N_9254);
or U9667 (N_9667,N_9351,N_9466);
and U9668 (N_9668,N_9409,N_9363);
or U9669 (N_9669,N_9286,N_9376);
and U9670 (N_9670,N_9279,N_9325);
nand U9671 (N_9671,N_9434,N_9492);
xnor U9672 (N_9672,N_9271,N_9396);
xor U9673 (N_9673,N_9451,N_9273);
nor U9674 (N_9674,N_9382,N_9485);
nor U9675 (N_9675,N_9286,N_9258);
and U9676 (N_9676,N_9292,N_9427);
and U9677 (N_9677,N_9494,N_9344);
nand U9678 (N_9678,N_9298,N_9426);
and U9679 (N_9679,N_9281,N_9266);
and U9680 (N_9680,N_9354,N_9455);
nor U9681 (N_9681,N_9344,N_9273);
and U9682 (N_9682,N_9473,N_9251);
xor U9683 (N_9683,N_9495,N_9251);
xnor U9684 (N_9684,N_9306,N_9319);
nor U9685 (N_9685,N_9385,N_9481);
or U9686 (N_9686,N_9456,N_9311);
nand U9687 (N_9687,N_9465,N_9338);
or U9688 (N_9688,N_9437,N_9321);
and U9689 (N_9689,N_9358,N_9373);
nor U9690 (N_9690,N_9410,N_9265);
nand U9691 (N_9691,N_9264,N_9327);
and U9692 (N_9692,N_9383,N_9344);
or U9693 (N_9693,N_9338,N_9385);
nand U9694 (N_9694,N_9404,N_9458);
and U9695 (N_9695,N_9398,N_9382);
or U9696 (N_9696,N_9282,N_9419);
nand U9697 (N_9697,N_9497,N_9316);
and U9698 (N_9698,N_9317,N_9379);
or U9699 (N_9699,N_9438,N_9313);
nand U9700 (N_9700,N_9354,N_9311);
nand U9701 (N_9701,N_9324,N_9337);
or U9702 (N_9702,N_9370,N_9330);
and U9703 (N_9703,N_9289,N_9377);
or U9704 (N_9704,N_9467,N_9359);
nand U9705 (N_9705,N_9255,N_9293);
and U9706 (N_9706,N_9279,N_9487);
nand U9707 (N_9707,N_9327,N_9310);
nor U9708 (N_9708,N_9360,N_9282);
nand U9709 (N_9709,N_9340,N_9315);
nand U9710 (N_9710,N_9392,N_9334);
and U9711 (N_9711,N_9337,N_9433);
nor U9712 (N_9712,N_9429,N_9427);
or U9713 (N_9713,N_9491,N_9326);
nand U9714 (N_9714,N_9380,N_9458);
and U9715 (N_9715,N_9296,N_9362);
or U9716 (N_9716,N_9370,N_9486);
or U9717 (N_9717,N_9272,N_9327);
and U9718 (N_9718,N_9357,N_9301);
and U9719 (N_9719,N_9487,N_9470);
or U9720 (N_9720,N_9274,N_9353);
and U9721 (N_9721,N_9263,N_9304);
or U9722 (N_9722,N_9444,N_9448);
or U9723 (N_9723,N_9465,N_9495);
nor U9724 (N_9724,N_9311,N_9465);
and U9725 (N_9725,N_9342,N_9397);
nor U9726 (N_9726,N_9466,N_9305);
xor U9727 (N_9727,N_9359,N_9415);
nand U9728 (N_9728,N_9380,N_9346);
nand U9729 (N_9729,N_9465,N_9460);
xor U9730 (N_9730,N_9461,N_9272);
or U9731 (N_9731,N_9452,N_9393);
nor U9732 (N_9732,N_9376,N_9258);
nor U9733 (N_9733,N_9325,N_9323);
nand U9734 (N_9734,N_9482,N_9253);
nor U9735 (N_9735,N_9372,N_9378);
nor U9736 (N_9736,N_9385,N_9480);
xor U9737 (N_9737,N_9250,N_9382);
and U9738 (N_9738,N_9390,N_9294);
or U9739 (N_9739,N_9252,N_9487);
nor U9740 (N_9740,N_9393,N_9489);
nor U9741 (N_9741,N_9470,N_9377);
nor U9742 (N_9742,N_9332,N_9401);
nand U9743 (N_9743,N_9284,N_9381);
nand U9744 (N_9744,N_9345,N_9446);
or U9745 (N_9745,N_9259,N_9288);
nor U9746 (N_9746,N_9270,N_9276);
and U9747 (N_9747,N_9321,N_9287);
or U9748 (N_9748,N_9402,N_9474);
xor U9749 (N_9749,N_9371,N_9332);
or U9750 (N_9750,N_9538,N_9589);
and U9751 (N_9751,N_9742,N_9708);
nand U9752 (N_9752,N_9710,N_9671);
nor U9753 (N_9753,N_9718,N_9681);
nand U9754 (N_9754,N_9517,N_9669);
and U9755 (N_9755,N_9536,N_9609);
nand U9756 (N_9756,N_9667,N_9737);
nor U9757 (N_9757,N_9626,N_9726);
xor U9758 (N_9758,N_9747,N_9534);
xor U9759 (N_9759,N_9709,N_9744);
nand U9760 (N_9760,N_9503,N_9688);
or U9761 (N_9761,N_9665,N_9720);
nor U9762 (N_9762,N_9684,N_9706);
nand U9763 (N_9763,N_9539,N_9585);
or U9764 (N_9764,N_9593,N_9734);
nand U9765 (N_9765,N_9532,N_9739);
or U9766 (N_9766,N_9654,N_9575);
or U9767 (N_9767,N_9557,N_9535);
and U9768 (N_9768,N_9602,N_9551);
and U9769 (N_9769,N_9633,N_9732);
or U9770 (N_9770,N_9572,N_9554);
nor U9771 (N_9771,N_9679,N_9675);
and U9772 (N_9772,N_9660,N_9701);
xnor U9773 (N_9773,N_9564,N_9603);
xor U9774 (N_9774,N_9627,N_9630);
xnor U9775 (N_9775,N_9512,N_9556);
nor U9776 (N_9776,N_9748,N_9550);
and U9777 (N_9777,N_9592,N_9662);
or U9778 (N_9778,N_9590,N_9659);
or U9779 (N_9779,N_9598,N_9735);
nor U9780 (N_9780,N_9670,N_9501);
nor U9781 (N_9781,N_9656,N_9693);
and U9782 (N_9782,N_9509,N_9635);
or U9783 (N_9783,N_9601,N_9652);
and U9784 (N_9784,N_9518,N_9611);
or U9785 (N_9785,N_9634,N_9588);
xnor U9786 (N_9786,N_9727,N_9678);
or U9787 (N_9787,N_9606,N_9698);
nor U9788 (N_9788,N_9699,N_9730);
and U9789 (N_9789,N_9731,N_9719);
nor U9790 (N_9790,N_9521,N_9607);
nor U9791 (N_9791,N_9676,N_9610);
nor U9792 (N_9792,N_9631,N_9714);
and U9793 (N_9793,N_9566,N_9568);
nor U9794 (N_9794,N_9527,N_9617);
nor U9795 (N_9795,N_9653,N_9571);
or U9796 (N_9796,N_9620,N_9577);
nor U9797 (N_9797,N_9646,N_9658);
and U9798 (N_9798,N_9600,N_9516);
and U9799 (N_9799,N_9548,N_9650);
or U9800 (N_9800,N_9599,N_9622);
or U9801 (N_9801,N_9692,N_9725);
xor U9802 (N_9802,N_9687,N_9682);
nor U9803 (N_9803,N_9613,N_9543);
xnor U9804 (N_9804,N_9594,N_9623);
or U9805 (N_9805,N_9580,N_9639);
and U9806 (N_9806,N_9636,N_9632);
nor U9807 (N_9807,N_9723,N_9537);
nor U9808 (N_9808,N_9582,N_9513);
and U9809 (N_9809,N_9570,N_9530);
or U9810 (N_9810,N_9717,N_9666);
nor U9811 (N_9811,N_9545,N_9638);
nor U9812 (N_9812,N_9612,N_9691);
or U9813 (N_9813,N_9621,N_9547);
nor U9814 (N_9814,N_9668,N_9649);
nand U9815 (N_9815,N_9629,N_9578);
or U9816 (N_9816,N_9746,N_9664);
nand U9817 (N_9817,N_9529,N_9643);
or U9818 (N_9818,N_9561,N_9586);
nand U9819 (N_9819,N_9741,N_9522);
nand U9820 (N_9820,N_9506,N_9644);
nor U9821 (N_9821,N_9648,N_9655);
xnor U9822 (N_9822,N_9715,N_9724);
and U9823 (N_9823,N_9624,N_9673);
or U9824 (N_9824,N_9702,N_9683);
nor U9825 (N_9825,N_9637,N_9553);
and U9826 (N_9826,N_9642,N_9713);
and U9827 (N_9827,N_9510,N_9689);
nor U9828 (N_9828,N_9700,N_9514);
or U9829 (N_9829,N_9595,N_9661);
xnor U9830 (N_9830,N_9574,N_9605);
nand U9831 (N_9831,N_9525,N_9552);
or U9832 (N_9832,N_9641,N_9576);
or U9833 (N_9833,N_9696,N_9504);
and U9834 (N_9834,N_9657,N_9618);
and U9835 (N_9835,N_9721,N_9560);
nor U9836 (N_9836,N_9562,N_9729);
nand U9837 (N_9837,N_9559,N_9672);
or U9838 (N_9838,N_9502,N_9549);
or U9839 (N_9839,N_9523,N_9695);
and U9840 (N_9840,N_9533,N_9645);
or U9841 (N_9841,N_9680,N_9528);
or U9842 (N_9842,N_9567,N_9728);
nor U9843 (N_9843,N_9583,N_9500);
or U9844 (N_9844,N_9531,N_9604);
xnor U9845 (N_9845,N_9722,N_9540);
and U9846 (N_9846,N_9555,N_9738);
nor U9847 (N_9847,N_9743,N_9524);
or U9848 (N_9848,N_9565,N_9515);
and U9849 (N_9849,N_9694,N_9685);
and U9850 (N_9850,N_9558,N_9614);
nor U9851 (N_9851,N_9597,N_9686);
nor U9852 (N_9852,N_9640,N_9511);
or U9853 (N_9853,N_9697,N_9542);
nor U9854 (N_9854,N_9584,N_9508);
nor U9855 (N_9855,N_9573,N_9505);
nor U9856 (N_9856,N_9581,N_9569);
xor U9857 (N_9857,N_9704,N_9712);
or U9858 (N_9858,N_9716,N_9663);
xor U9859 (N_9859,N_9651,N_9608);
xnor U9860 (N_9860,N_9711,N_9690);
and U9861 (N_9861,N_9740,N_9587);
or U9862 (N_9862,N_9703,N_9507);
or U9863 (N_9863,N_9677,N_9736);
nand U9864 (N_9864,N_9563,N_9625);
nand U9865 (N_9865,N_9674,N_9616);
nand U9866 (N_9866,N_9544,N_9749);
xor U9867 (N_9867,N_9619,N_9628);
nor U9868 (N_9868,N_9707,N_9526);
and U9869 (N_9869,N_9591,N_9519);
nand U9870 (N_9870,N_9615,N_9520);
and U9871 (N_9871,N_9579,N_9596);
xnor U9872 (N_9872,N_9546,N_9745);
or U9873 (N_9873,N_9705,N_9541);
and U9874 (N_9874,N_9733,N_9647);
xor U9875 (N_9875,N_9653,N_9516);
xnor U9876 (N_9876,N_9524,N_9646);
or U9877 (N_9877,N_9658,N_9681);
or U9878 (N_9878,N_9534,N_9549);
nand U9879 (N_9879,N_9710,N_9688);
and U9880 (N_9880,N_9515,N_9664);
xnor U9881 (N_9881,N_9596,N_9532);
nor U9882 (N_9882,N_9600,N_9586);
or U9883 (N_9883,N_9671,N_9608);
nand U9884 (N_9884,N_9620,N_9508);
xnor U9885 (N_9885,N_9606,N_9604);
or U9886 (N_9886,N_9614,N_9747);
and U9887 (N_9887,N_9740,N_9549);
nor U9888 (N_9888,N_9679,N_9597);
and U9889 (N_9889,N_9669,N_9520);
nor U9890 (N_9890,N_9717,N_9619);
xnor U9891 (N_9891,N_9513,N_9628);
or U9892 (N_9892,N_9642,N_9595);
or U9893 (N_9893,N_9662,N_9653);
and U9894 (N_9894,N_9512,N_9703);
or U9895 (N_9895,N_9609,N_9719);
nor U9896 (N_9896,N_9600,N_9501);
nand U9897 (N_9897,N_9621,N_9539);
nand U9898 (N_9898,N_9522,N_9596);
or U9899 (N_9899,N_9531,N_9610);
or U9900 (N_9900,N_9731,N_9744);
nand U9901 (N_9901,N_9589,N_9582);
nor U9902 (N_9902,N_9547,N_9738);
nand U9903 (N_9903,N_9593,N_9696);
nor U9904 (N_9904,N_9739,N_9582);
and U9905 (N_9905,N_9695,N_9680);
nand U9906 (N_9906,N_9656,N_9517);
and U9907 (N_9907,N_9595,N_9669);
or U9908 (N_9908,N_9736,N_9523);
or U9909 (N_9909,N_9648,N_9603);
nand U9910 (N_9910,N_9589,N_9668);
nand U9911 (N_9911,N_9714,N_9742);
or U9912 (N_9912,N_9591,N_9564);
and U9913 (N_9913,N_9706,N_9675);
nor U9914 (N_9914,N_9527,N_9745);
and U9915 (N_9915,N_9711,N_9649);
and U9916 (N_9916,N_9679,N_9656);
nand U9917 (N_9917,N_9617,N_9565);
or U9918 (N_9918,N_9640,N_9540);
or U9919 (N_9919,N_9628,N_9722);
nor U9920 (N_9920,N_9586,N_9631);
or U9921 (N_9921,N_9595,N_9503);
xnor U9922 (N_9922,N_9576,N_9563);
or U9923 (N_9923,N_9703,N_9521);
and U9924 (N_9924,N_9600,N_9575);
nand U9925 (N_9925,N_9543,N_9572);
or U9926 (N_9926,N_9579,N_9638);
nor U9927 (N_9927,N_9536,N_9641);
nor U9928 (N_9928,N_9642,N_9677);
xnor U9929 (N_9929,N_9737,N_9609);
nand U9930 (N_9930,N_9574,N_9666);
and U9931 (N_9931,N_9724,N_9509);
or U9932 (N_9932,N_9507,N_9558);
or U9933 (N_9933,N_9632,N_9547);
and U9934 (N_9934,N_9748,N_9613);
xnor U9935 (N_9935,N_9569,N_9553);
nor U9936 (N_9936,N_9685,N_9547);
xnor U9937 (N_9937,N_9638,N_9608);
nor U9938 (N_9938,N_9682,N_9737);
nand U9939 (N_9939,N_9583,N_9593);
and U9940 (N_9940,N_9622,N_9619);
and U9941 (N_9941,N_9516,N_9627);
nand U9942 (N_9942,N_9600,N_9504);
nor U9943 (N_9943,N_9637,N_9570);
or U9944 (N_9944,N_9626,N_9542);
or U9945 (N_9945,N_9554,N_9734);
or U9946 (N_9946,N_9522,N_9617);
or U9947 (N_9947,N_9611,N_9598);
or U9948 (N_9948,N_9517,N_9641);
xor U9949 (N_9949,N_9656,N_9717);
and U9950 (N_9950,N_9568,N_9720);
nand U9951 (N_9951,N_9596,N_9666);
or U9952 (N_9952,N_9579,N_9744);
and U9953 (N_9953,N_9621,N_9531);
nand U9954 (N_9954,N_9638,N_9627);
and U9955 (N_9955,N_9594,N_9653);
nand U9956 (N_9956,N_9653,N_9720);
xnor U9957 (N_9957,N_9691,N_9510);
nor U9958 (N_9958,N_9579,N_9601);
nor U9959 (N_9959,N_9515,N_9749);
or U9960 (N_9960,N_9600,N_9724);
nand U9961 (N_9961,N_9551,N_9730);
and U9962 (N_9962,N_9648,N_9548);
nand U9963 (N_9963,N_9728,N_9671);
nand U9964 (N_9964,N_9512,N_9670);
nand U9965 (N_9965,N_9594,N_9573);
xor U9966 (N_9966,N_9558,N_9657);
nor U9967 (N_9967,N_9684,N_9593);
or U9968 (N_9968,N_9550,N_9665);
xor U9969 (N_9969,N_9603,N_9672);
nor U9970 (N_9970,N_9670,N_9735);
or U9971 (N_9971,N_9567,N_9509);
nand U9972 (N_9972,N_9524,N_9747);
nor U9973 (N_9973,N_9707,N_9656);
nand U9974 (N_9974,N_9610,N_9577);
and U9975 (N_9975,N_9749,N_9624);
nand U9976 (N_9976,N_9516,N_9605);
or U9977 (N_9977,N_9501,N_9689);
nor U9978 (N_9978,N_9619,N_9680);
or U9979 (N_9979,N_9612,N_9709);
and U9980 (N_9980,N_9564,N_9565);
or U9981 (N_9981,N_9632,N_9652);
xor U9982 (N_9982,N_9586,N_9590);
nand U9983 (N_9983,N_9519,N_9523);
or U9984 (N_9984,N_9565,N_9534);
and U9985 (N_9985,N_9697,N_9677);
or U9986 (N_9986,N_9608,N_9544);
or U9987 (N_9987,N_9611,N_9615);
and U9988 (N_9988,N_9739,N_9536);
and U9989 (N_9989,N_9727,N_9502);
nor U9990 (N_9990,N_9742,N_9561);
nand U9991 (N_9991,N_9559,N_9646);
or U9992 (N_9992,N_9512,N_9638);
and U9993 (N_9993,N_9730,N_9705);
nor U9994 (N_9994,N_9542,N_9722);
nor U9995 (N_9995,N_9525,N_9700);
nor U9996 (N_9996,N_9704,N_9530);
xnor U9997 (N_9997,N_9522,N_9533);
nor U9998 (N_9998,N_9538,N_9556);
nand U9999 (N_9999,N_9563,N_9633);
nand U10000 (N_10000,N_9860,N_9907);
nor U10001 (N_10001,N_9855,N_9998);
nor U10002 (N_10002,N_9778,N_9839);
nand U10003 (N_10003,N_9838,N_9758);
nor U10004 (N_10004,N_9824,N_9903);
nor U10005 (N_10005,N_9912,N_9785);
nor U10006 (N_10006,N_9917,N_9941);
or U10007 (N_10007,N_9762,N_9757);
or U10008 (N_10008,N_9773,N_9786);
nor U10009 (N_10009,N_9890,N_9856);
nor U10010 (N_10010,N_9799,N_9957);
and U10011 (N_10011,N_9982,N_9805);
or U10012 (N_10012,N_9835,N_9764);
nand U10013 (N_10013,N_9961,N_9885);
or U10014 (N_10014,N_9775,N_9916);
xnor U10015 (N_10015,N_9965,N_9974);
or U10016 (N_10016,N_9829,N_9783);
nand U10017 (N_10017,N_9940,N_9767);
nand U10018 (N_10018,N_9892,N_9989);
nor U10019 (N_10019,N_9877,N_9910);
nand U10020 (N_10020,N_9928,N_9949);
or U10021 (N_10021,N_9858,N_9886);
nor U10022 (N_10022,N_9825,N_9809);
or U10023 (N_10023,N_9819,N_9863);
and U10024 (N_10024,N_9776,N_9875);
or U10025 (N_10025,N_9792,N_9942);
or U10026 (N_10026,N_9761,N_9960);
or U10027 (N_10027,N_9955,N_9993);
or U10028 (N_10028,N_9843,N_9755);
and U10029 (N_10029,N_9795,N_9823);
nor U10030 (N_10030,N_9876,N_9953);
or U10031 (N_10031,N_9954,N_9756);
nand U10032 (N_10032,N_9872,N_9899);
xnor U10033 (N_10033,N_9870,N_9862);
nor U10034 (N_10034,N_9898,N_9931);
nand U10035 (N_10035,N_9883,N_9781);
or U10036 (N_10036,N_9996,N_9750);
and U10037 (N_10037,N_9936,N_9920);
and U10038 (N_10038,N_9911,N_9826);
nand U10039 (N_10039,N_9810,N_9811);
or U10040 (N_10040,N_9933,N_9895);
xnor U10041 (N_10041,N_9844,N_9999);
nor U10042 (N_10042,N_9754,N_9913);
nor U10043 (N_10043,N_9906,N_9978);
nor U10044 (N_10044,N_9927,N_9925);
nand U10045 (N_10045,N_9963,N_9812);
or U10046 (N_10046,N_9929,N_9793);
or U10047 (N_10047,N_9969,N_9976);
or U10048 (N_10048,N_9851,N_9852);
or U10049 (N_10049,N_9766,N_9820);
nor U10050 (N_10050,N_9956,N_9796);
nand U10051 (N_10051,N_9808,N_9787);
or U10052 (N_10052,N_9948,N_9791);
and U10053 (N_10053,N_9814,N_9822);
or U10054 (N_10054,N_9962,N_9831);
or U10055 (N_10055,N_9945,N_9944);
nand U10056 (N_10056,N_9951,N_9901);
nand U10057 (N_10057,N_9794,N_9866);
and U10058 (N_10058,N_9857,N_9818);
nand U10059 (N_10059,N_9935,N_9986);
and U10060 (N_10060,N_9842,N_9841);
nor U10061 (N_10061,N_9865,N_9804);
and U10062 (N_10062,N_9830,N_9943);
nand U10063 (N_10063,N_9815,N_9952);
or U10064 (N_10064,N_9926,N_9834);
xor U10065 (N_10065,N_9840,N_9788);
and U10066 (N_10066,N_9873,N_9801);
xor U10067 (N_10067,N_9970,N_9971);
xor U10068 (N_10068,N_9868,N_9897);
and U10069 (N_10069,N_9915,N_9784);
nand U10070 (N_10070,N_9871,N_9988);
and U10071 (N_10071,N_9759,N_9847);
or U10072 (N_10072,N_9854,N_9807);
nor U10073 (N_10073,N_9924,N_9769);
xnor U10074 (N_10074,N_9753,N_9896);
and U10075 (N_10075,N_9777,N_9760);
nor U10076 (N_10076,N_9900,N_9946);
or U10077 (N_10077,N_9779,N_9832);
nand U10078 (N_10078,N_9763,N_9816);
nand U10079 (N_10079,N_9751,N_9914);
or U10080 (N_10080,N_9893,N_9967);
xor U10081 (N_10081,N_9836,N_9889);
nor U10082 (N_10082,N_9797,N_9765);
and U10083 (N_10083,N_9947,N_9798);
nand U10084 (N_10084,N_9806,N_9950);
and U10085 (N_10085,N_9992,N_9845);
and U10086 (N_10086,N_9849,N_9828);
nand U10087 (N_10087,N_9983,N_9780);
nand U10088 (N_10088,N_9772,N_9770);
nor U10089 (N_10089,N_9921,N_9939);
nand U10090 (N_10090,N_9874,N_9994);
nand U10091 (N_10091,N_9867,N_9904);
xnor U10092 (N_10092,N_9966,N_9972);
or U10093 (N_10093,N_9959,N_9881);
xor U10094 (N_10094,N_9908,N_9833);
xnor U10095 (N_10095,N_9923,N_9869);
nor U10096 (N_10096,N_9932,N_9752);
nand U10097 (N_10097,N_9888,N_9850);
and U10098 (N_10098,N_9958,N_9853);
nand U10099 (N_10099,N_9977,N_9837);
nor U10100 (N_10100,N_9846,N_9817);
nor U10101 (N_10101,N_9979,N_9902);
and U10102 (N_10102,N_9848,N_9894);
xor U10103 (N_10103,N_9864,N_9973);
nor U10104 (N_10104,N_9782,N_9938);
or U10105 (N_10105,N_9802,N_9882);
or U10106 (N_10106,N_9919,N_9821);
or U10107 (N_10107,N_9887,N_9937);
xor U10108 (N_10108,N_9774,N_9909);
or U10109 (N_10109,N_9922,N_9980);
nand U10110 (N_10110,N_9985,N_9878);
xnor U10111 (N_10111,N_9991,N_9803);
nand U10112 (N_10112,N_9984,N_9918);
nor U10113 (N_10113,N_9879,N_9905);
and U10114 (N_10114,N_9891,N_9997);
nor U10115 (N_10115,N_9990,N_9771);
or U10116 (N_10116,N_9827,N_9995);
nand U10117 (N_10117,N_9859,N_9968);
nand U10118 (N_10118,N_9884,N_9934);
nor U10119 (N_10119,N_9880,N_9987);
nor U10120 (N_10120,N_9964,N_9789);
nand U10121 (N_10121,N_9930,N_9861);
or U10122 (N_10122,N_9790,N_9768);
or U10123 (N_10123,N_9800,N_9975);
or U10124 (N_10124,N_9981,N_9813);
nand U10125 (N_10125,N_9990,N_9943);
nand U10126 (N_10126,N_9882,N_9914);
nor U10127 (N_10127,N_9903,N_9889);
or U10128 (N_10128,N_9795,N_9923);
and U10129 (N_10129,N_9830,N_9840);
nand U10130 (N_10130,N_9985,N_9875);
or U10131 (N_10131,N_9842,N_9972);
or U10132 (N_10132,N_9992,N_9976);
nand U10133 (N_10133,N_9926,N_9998);
and U10134 (N_10134,N_9825,N_9969);
nor U10135 (N_10135,N_9927,N_9833);
nand U10136 (N_10136,N_9946,N_9809);
xnor U10137 (N_10137,N_9852,N_9780);
or U10138 (N_10138,N_9852,N_9831);
nand U10139 (N_10139,N_9890,N_9815);
nor U10140 (N_10140,N_9829,N_9754);
and U10141 (N_10141,N_9980,N_9986);
nand U10142 (N_10142,N_9924,N_9992);
nand U10143 (N_10143,N_9970,N_9812);
nand U10144 (N_10144,N_9986,N_9852);
and U10145 (N_10145,N_9857,N_9977);
or U10146 (N_10146,N_9776,N_9945);
nand U10147 (N_10147,N_9904,N_9772);
or U10148 (N_10148,N_9901,N_9851);
or U10149 (N_10149,N_9893,N_9841);
or U10150 (N_10150,N_9757,N_9828);
nor U10151 (N_10151,N_9995,N_9779);
nor U10152 (N_10152,N_9779,N_9943);
or U10153 (N_10153,N_9921,N_9923);
nor U10154 (N_10154,N_9891,N_9906);
or U10155 (N_10155,N_9826,N_9772);
and U10156 (N_10156,N_9958,N_9801);
and U10157 (N_10157,N_9774,N_9819);
and U10158 (N_10158,N_9967,N_9918);
nand U10159 (N_10159,N_9847,N_9793);
xor U10160 (N_10160,N_9762,N_9921);
nand U10161 (N_10161,N_9916,N_9802);
xnor U10162 (N_10162,N_9762,N_9760);
and U10163 (N_10163,N_9902,N_9944);
or U10164 (N_10164,N_9838,N_9817);
or U10165 (N_10165,N_9835,N_9937);
nor U10166 (N_10166,N_9839,N_9861);
nand U10167 (N_10167,N_9842,N_9961);
and U10168 (N_10168,N_9976,N_9919);
or U10169 (N_10169,N_9931,N_9963);
nor U10170 (N_10170,N_9763,N_9832);
and U10171 (N_10171,N_9957,N_9877);
nor U10172 (N_10172,N_9971,N_9966);
xor U10173 (N_10173,N_9891,N_9850);
nor U10174 (N_10174,N_9879,N_9847);
nor U10175 (N_10175,N_9995,N_9828);
and U10176 (N_10176,N_9837,N_9774);
xor U10177 (N_10177,N_9830,N_9843);
nand U10178 (N_10178,N_9919,N_9925);
and U10179 (N_10179,N_9949,N_9841);
nand U10180 (N_10180,N_9950,N_9792);
and U10181 (N_10181,N_9964,N_9940);
and U10182 (N_10182,N_9825,N_9898);
nor U10183 (N_10183,N_9827,N_9886);
and U10184 (N_10184,N_9977,N_9785);
or U10185 (N_10185,N_9955,N_9991);
nor U10186 (N_10186,N_9874,N_9817);
or U10187 (N_10187,N_9924,N_9904);
nand U10188 (N_10188,N_9897,N_9752);
and U10189 (N_10189,N_9900,N_9750);
or U10190 (N_10190,N_9980,N_9814);
and U10191 (N_10191,N_9992,N_9850);
nor U10192 (N_10192,N_9767,N_9869);
and U10193 (N_10193,N_9924,N_9972);
and U10194 (N_10194,N_9811,N_9769);
and U10195 (N_10195,N_9945,N_9913);
xor U10196 (N_10196,N_9978,N_9781);
or U10197 (N_10197,N_9876,N_9989);
xnor U10198 (N_10198,N_9976,N_9857);
nand U10199 (N_10199,N_9821,N_9995);
or U10200 (N_10200,N_9820,N_9856);
and U10201 (N_10201,N_9853,N_9770);
and U10202 (N_10202,N_9792,N_9952);
and U10203 (N_10203,N_9999,N_9877);
or U10204 (N_10204,N_9804,N_9896);
nand U10205 (N_10205,N_9829,N_9868);
or U10206 (N_10206,N_9984,N_9977);
and U10207 (N_10207,N_9934,N_9978);
or U10208 (N_10208,N_9818,N_9778);
and U10209 (N_10209,N_9892,N_9854);
xnor U10210 (N_10210,N_9775,N_9760);
and U10211 (N_10211,N_9979,N_9967);
and U10212 (N_10212,N_9922,N_9998);
and U10213 (N_10213,N_9823,N_9784);
and U10214 (N_10214,N_9813,N_9933);
nor U10215 (N_10215,N_9789,N_9890);
and U10216 (N_10216,N_9977,N_9835);
and U10217 (N_10217,N_9833,N_9752);
and U10218 (N_10218,N_9912,N_9824);
xnor U10219 (N_10219,N_9994,N_9963);
or U10220 (N_10220,N_9942,N_9913);
nand U10221 (N_10221,N_9906,N_9756);
or U10222 (N_10222,N_9757,N_9830);
nor U10223 (N_10223,N_9996,N_9990);
or U10224 (N_10224,N_9833,N_9858);
and U10225 (N_10225,N_9847,N_9968);
or U10226 (N_10226,N_9997,N_9983);
nand U10227 (N_10227,N_9952,N_9974);
and U10228 (N_10228,N_9952,N_9992);
nand U10229 (N_10229,N_9875,N_9954);
nor U10230 (N_10230,N_9932,N_9827);
nand U10231 (N_10231,N_9935,N_9888);
xnor U10232 (N_10232,N_9754,N_9932);
nand U10233 (N_10233,N_9829,N_9875);
nand U10234 (N_10234,N_9763,N_9833);
nor U10235 (N_10235,N_9833,N_9926);
and U10236 (N_10236,N_9805,N_9910);
nand U10237 (N_10237,N_9944,N_9877);
or U10238 (N_10238,N_9955,N_9977);
nand U10239 (N_10239,N_9945,N_9880);
and U10240 (N_10240,N_9863,N_9772);
and U10241 (N_10241,N_9932,N_9895);
and U10242 (N_10242,N_9893,N_9935);
and U10243 (N_10243,N_9789,N_9946);
nor U10244 (N_10244,N_9808,N_9976);
xnor U10245 (N_10245,N_9784,N_9793);
nor U10246 (N_10246,N_9984,N_9904);
nand U10247 (N_10247,N_9938,N_9796);
nor U10248 (N_10248,N_9798,N_9890);
nor U10249 (N_10249,N_9800,N_9801);
nand U10250 (N_10250,N_10081,N_10195);
nor U10251 (N_10251,N_10221,N_10149);
nor U10252 (N_10252,N_10125,N_10175);
or U10253 (N_10253,N_10211,N_10121);
and U10254 (N_10254,N_10040,N_10181);
and U10255 (N_10255,N_10031,N_10100);
and U10256 (N_10256,N_10109,N_10237);
nor U10257 (N_10257,N_10154,N_10024);
nand U10258 (N_10258,N_10080,N_10161);
nand U10259 (N_10259,N_10135,N_10172);
nor U10260 (N_10260,N_10069,N_10225);
nor U10261 (N_10261,N_10131,N_10168);
nor U10262 (N_10262,N_10037,N_10174);
nand U10263 (N_10263,N_10076,N_10010);
nor U10264 (N_10264,N_10228,N_10022);
or U10265 (N_10265,N_10042,N_10112);
and U10266 (N_10266,N_10227,N_10045);
and U10267 (N_10267,N_10170,N_10056);
nor U10268 (N_10268,N_10219,N_10019);
and U10269 (N_10269,N_10026,N_10214);
or U10270 (N_10270,N_10075,N_10184);
nand U10271 (N_10271,N_10060,N_10111);
nor U10272 (N_10272,N_10063,N_10070);
nor U10273 (N_10273,N_10000,N_10122);
nor U10274 (N_10274,N_10030,N_10004);
nor U10275 (N_10275,N_10114,N_10164);
xor U10276 (N_10276,N_10151,N_10067);
or U10277 (N_10277,N_10082,N_10048);
or U10278 (N_10278,N_10012,N_10206);
and U10279 (N_10279,N_10126,N_10029);
xor U10280 (N_10280,N_10091,N_10025);
xor U10281 (N_10281,N_10079,N_10187);
and U10282 (N_10282,N_10016,N_10053);
nand U10283 (N_10283,N_10192,N_10057);
and U10284 (N_10284,N_10208,N_10018);
or U10285 (N_10285,N_10118,N_10007);
nand U10286 (N_10286,N_10136,N_10215);
and U10287 (N_10287,N_10110,N_10226);
nor U10288 (N_10288,N_10173,N_10236);
xor U10289 (N_10289,N_10142,N_10143);
nor U10290 (N_10290,N_10054,N_10137);
or U10291 (N_10291,N_10127,N_10191);
and U10292 (N_10292,N_10145,N_10116);
and U10293 (N_10293,N_10133,N_10178);
and U10294 (N_10294,N_10249,N_10093);
xnor U10295 (N_10295,N_10005,N_10113);
and U10296 (N_10296,N_10052,N_10244);
and U10297 (N_10297,N_10139,N_10073);
nor U10298 (N_10298,N_10217,N_10130);
or U10299 (N_10299,N_10240,N_10182);
xnor U10300 (N_10300,N_10158,N_10115);
nand U10301 (N_10301,N_10027,N_10190);
and U10302 (N_10302,N_10020,N_10062);
nor U10303 (N_10303,N_10059,N_10041);
or U10304 (N_10304,N_10085,N_10205);
nand U10305 (N_10305,N_10224,N_10159);
or U10306 (N_10306,N_10032,N_10223);
nand U10307 (N_10307,N_10209,N_10165);
and U10308 (N_10308,N_10084,N_10071);
nand U10309 (N_10309,N_10108,N_10101);
nor U10310 (N_10310,N_10144,N_10064);
nor U10311 (N_10311,N_10105,N_10138);
nor U10312 (N_10312,N_10028,N_10203);
nand U10313 (N_10313,N_10207,N_10183);
or U10314 (N_10314,N_10167,N_10086);
or U10315 (N_10315,N_10166,N_10176);
or U10316 (N_10316,N_10128,N_10120);
or U10317 (N_10317,N_10096,N_10050);
and U10318 (N_10318,N_10169,N_10047);
and U10319 (N_10319,N_10193,N_10021);
and U10320 (N_10320,N_10134,N_10160);
nor U10321 (N_10321,N_10017,N_10186);
nor U10322 (N_10322,N_10231,N_10095);
xor U10323 (N_10323,N_10238,N_10148);
or U10324 (N_10324,N_10243,N_10204);
nor U10325 (N_10325,N_10212,N_10008);
nor U10326 (N_10326,N_10147,N_10092);
or U10327 (N_10327,N_10034,N_10180);
or U10328 (N_10328,N_10083,N_10094);
nand U10329 (N_10329,N_10124,N_10119);
and U10330 (N_10330,N_10163,N_10155);
nor U10331 (N_10331,N_10216,N_10104);
xor U10332 (N_10332,N_10189,N_10242);
nand U10333 (N_10333,N_10055,N_10234);
xnor U10334 (N_10334,N_10046,N_10199);
nor U10335 (N_10335,N_10014,N_10089);
nand U10336 (N_10336,N_10011,N_10198);
and U10337 (N_10337,N_10157,N_10090);
and U10338 (N_10338,N_10107,N_10013);
and U10339 (N_10339,N_10074,N_10194);
nand U10340 (N_10340,N_10015,N_10220);
or U10341 (N_10341,N_10132,N_10202);
nand U10342 (N_10342,N_10150,N_10245);
nor U10343 (N_10343,N_10171,N_10117);
nor U10344 (N_10344,N_10088,N_10087);
xor U10345 (N_10345,N_10066,N_10077);
and U10346 (N_10346,N_10072,N_10156);
or U10347 (N_10347,N_10247,N_10248);
nor U10348 (N_10348,N_10210,N_10185);
or U10349 (N_10349,N_10196,N_10246);
nor U10350 (N_10350,N_10241,N_10043);
and U10351 (N_10351,N_10222,N_10001);
nor U10352 (N_10352,N_10065,N_10035);
nand U10353 (N_10353,N_10232,N_10036);
xnor U10354 (N_10354,N_10068,N_10099);
xor U10355 (N_10355,N_10051,N_10200);
xor U10356 (N_10356,N_10103,N_10003);
nor U10357 (N_10357,N_10038,N_10213);
and U10358 (N_10358,N_10146,N_10098);
nand U10359 (N_10359,N_10230,N_10006);
nand U10360 (N_10360,N_10097,N_10140);
or U10361 (N_10361,N_10039,N_10188);
nand U10362 (N_10362,N_10078,N_10179);
nor U10363 (N_10363,N_10233,N_10229);
nand U10364 (N_10364,N_10033,N_10239);
xor U10365 (N_10365,N_10106,N_10044);
and U10366 (N_10366,N_10061,N_10218);
and U10367 (N_10367,N_10177,N_10197);
and U10368 (N_10368,N_10123,N_10049);
nand U10369 (N_10369,N_10102,N_10002);
or U10370 (N_10370,N_10162,N_10023);
nand U10371 (N_10371,N_10235,N_10201);
nor U10372 (N_10372,N_10141,N_10009);
or U10373 (N_10373,N_10152,N_10058);
xor U10374 (N_10374,N_10129,N_10153);
nand U10375 (N_10375,N_10234,N_10174);
and U10376 (N_10376,N_10086,N_10030);
nor U10377 (N_10377,N_10104,N_10220);
and U10378 (N_10378,N_10242,N_10088);
nor U10379 (N_10379,N_10060,N_10047);
nor U10380 (N_10380,N_10070,N_10186);
nor U10381 (N_10381,N_10021,N_10096);
nor U10382 (N_10382,N_10013,N_10248);
and U10383 (N_10383,N_10023,N_10201);
or U10384 (N_10384,N_10133,N_10206);
xnor U10385 (N_10385,N_10235,N_10239);
and U10386 (N_10386,N_10201,N_10236);
nand U10387 (N_10387,N_10050,N_10042);
xor U10388 (N_10388,N_10075,N_10120);
xnor U10389 (N_10389,N_10207,N_10157);
and U10390 (N_10390,N_10221,N_10116);
and U10391 (N_10391,N_10050,N_10106);
and U10392 (N_10392,N_10222,N_10179);
and U10393 (N_10393,N_10099,N_10119);
nand U10394 (N_10394,N_10099,N_10206);
or U10395 (N_10395,N_10168,N_10033);
and U10396 (N_10396,N_10047,N_10137);
or U10397 (N_10397,N_10005,N_10225);
or U10398 (N_10398,N_10037,N_10076);
nand U10399 (N_10399,N_10236,N_10013);
nor U10400 (N_10400,N_10057,N_10206);
nor U10401 (N_10401,N_10230,N_10018);
xor U10402 (N_10402,N_10069,N_10009);
nor U10403 (N_10403,N_10138,N_10033);
nor U10404 (N_10404,N_10239,N_10149);
and U10405 (N_10405,N_10028,N_10181);
and U10406 (N_10406,N_10058,N_10142);
or U10407 (N_10407,N_10134,N_10204);
and U10408 (N_10408,N_10113,N_10053);
or U10409 (N_10409,N_10244,N_10225);
nand U10410 (N_10410,N_10088,N_10009);
xor U10411 (N_10411,N_10162,N_10018);
xor U10412 (N_10412,N_10081,N_10157);
or U10413 (N_10413,N_10053,N_10128);
and U10414 (N_10414,N_10147,N_10242);
nand U10415 (N_10415,N_10101,N_10059);
nor U10416 (N_10416,N_10059,N_10159);
nor U10417 (N_10417,N_10046,N_10035);
nor U10418 (N_10418,N_10181,N_10053);
nor U10419 (N_10419,N_10101,N_10203);
nand U10420 (N_10420,N_10078,N_10175);
and U10421 (N_10421,N_10241,N_10107);
or U10422 (N_10422,N_10161,N_10134);
nor U10423 (N_10423,N_10011,N_10102);
and U10424 (N_10424,N_10199,N_10187);
nand U10425 (N_10425,N_10170,N_10098);
or U10426 (N_10426,N_10047,N_10088);
xnor U10427 (N_10427,N_10088,N_10016);
nor U10428 (N_10428,N_10059,N_10177);
or U10429 (N_10429,N_10158,N_10162);
nor U10430 (N_10430,N_10203,N_10143);
nand U10431 (N_10431,N_10099,N_10091);
nand U10432 (N_10432,N_10082,N_10019);
xnor U10433 (N_10433,N_10000,N_10138);
nand U10434 (N_10434,N_10050,N_10047);
nand U10435 (N_10435,N_10085,N_10042);
and U10436 (N_10436,N_10042,N_10196);
or U10437 (N_10437,N_10204,N_10159);
nand U10438 (N_10438,N_10215,N_10101);
nor U10439 (N_10439,N_10091,N_10046);
nor U10440 (N_10440,N_10246,N_10233);
and U10441 (N_10441,N_10183,N_10121);
and U10442 (N_10442,N_10095,N_10215);
nand U10443 (N_10443,N_10155,N_10141);
nand U10444 (N_10444,N_10123,N_10223);
xnor U10445 (N_10445,N_10197,N_10101);
xnor U10446 (N_10446,N_10016,N_10246);
nand U10447 (N_10447,N_10182,N_10110);
nor U10448 (N_10448,N_10016,N_10002);
xnor U10449 (N_10449,N_10043,N_10085);
or U10450 (N_10450,N_10142,N_10190);
or U10451 (N_10451,N_10063,N_10116);
nand U10452 (N_10452,N_10126,N_10148);
nor U10453 (N_10453,N_10085,N_10124);
and U10454 (N_10454,N_10216,N_10060);
nor U10455 (N_10455,N_10158,N_10119);
and U10456 (N_10456,N_10247,N_10148);
or U10457 (N_10457,N_10035,N_10153);
or U10458 (N_10458,N_10164,N_10001);
or U10459 (N_10459,N_10123,N_10182);
nand U10460 (N_10460,N_10157,N_10209);
nand U10461 (N_10461,N_10004,N_10108);
or U10462 (N_10462,N_10003,N_10153);
xnor U10463 (N_10463,N_10172,N_10108);
nor U10464 (N_10464,N_10105,N_10052);
nor U10465 (N_10465,N_10085,N_10123);
and U10466 (N_10466,N_10192,N_10203);
nor U10467 (N_10467,N_10105,N_10102);
and U10468 (N_10468,N_10214,N_10046);
or U10469 (N_10469,N_10150,N_10000);
nor U10470 (N_10470,N_10055,N_10184);
and U10471 (N_10471,N_10017,N_10079);
or U10472 (N_10472,N_10238,N_10059);
nand U10473 (N_10473,N_10208,N_10165);
or U10474 (N_10474,N_10106,N_10230);
nand U10475 (N_10475,N_10125,N_10200);
or U10476 (N_10476,N_10248,N_10141);
nor U10477 (N_10477,N_10121,N_10177);
nand U10478 (N_10478,N_10176,N_10203);
and U10479 (N_10479,N_10017,N_10138);
xor U10480 (N_10480,N_10075,N_10245);
nor U10481 (N_10481,N_10029,N_10059);
or U10482 (N_10482,N_10089,N_10114);
or U10483 (N_10483,N_10029,N_10171);
xnor U10484 (N_10484,N_10056,N_10124);
nand U10485 (N_10485,N_10214,N_10131);
or U10486 (N_10486,N_10245,N_10163);
nand U10487 (N_10487,N_10007,N_10200);
nand U10488 (N_10488,N_10092,N_10174);
nor U10489 (N_10489,N_10034,N_10227);
nor U10490 (N_10490,N_10070,N_10058);
xor U10491 (N_10491,N_10148,N_10176);
nand U10492 (N_10492,N_10070,N_10156);
nor U10493 (N_10493,N_10024,N_10029);
or U10494 (N_10494,N_10157,N_10037);
nor U10495 (N_10495,N_10119,N_10073);
nand U10496 (N_10496,N_10034,N_10098);
nor U10497 (N_10497,N_10042,N_10015);
or U10498 (N_10498,N_10112,N_10146);
nor U10499 (N_10499,N_10099,N_10201);
or U10500 (N_10500,N_10460,N_10475);
or U10501 (N_10501,N_10273,N_10416);
and U10502 (N_10502,N_10427,N_10397);
nand U10503 (N_10503,N_10330,N_10333);
nand U10504 (N_10504,N_10408,N_10282);
and U10505 (N_10505,N_10342,N_10453);
or U10506 (N_10506,N_10386,N_10417);
nor U10507 (N_10507,N_10355,N_10472);
nor U10508 (N_10508,N_10369,N_10296);
nor U10509 (N_10509,N_10451,N_10395);
or U10510 (N_10510,N_10498,N_10341);
or U10511 (N_10511,N_10365,N_10492);
xnor U10512 (N_10512,N_10388,N_10400);
or U10513 (N_10513,N_10274,N_10410);
or U10514 (N_10514,N_10253,N_10478);
or U10515 (N_10515,N_10422,N_10294);
and U10516 (N_10516,N_10412,N_10316);
or U10517 (N_10517,N_10448,N_10463);
and U10518 (N_10518,N_10315,N_10279);
or U10519 (N_10519,N_10260,N_10298);
or U10520 (N_10520,N_10252,N_10285);
and U10521 (N_10521,N_10444,N_10483);
nor U10522 (N_10522,N_10339,N_10396);
and U10523 (N_10523,N_10467,N_10382);
and U10524 (N_10524,N_10356,N_10265);
nand U10525 (N_10525,N_10357,N_10368);
nor U10526 (N_10526,N_10323,N_10367);
xor U10527 (N_10527,N_10270,N_10462);
xnor U10528 (N_10528,N_10403,N_10343);
and U10529 (N_10529,N_10301,N_10495);
and U10530 (N_10530,N_10360,N_10289);
xor U10531 (N_10531,N_10377,N_10267);
or U10532 (N_10532,N_10476,N_10250);
nand U10533 (N_10533,N_10307,N_10327);
nand U10534 (N_10534,N_10373,N_10364);
nand U10535 (N_10535,N_10271,N_10349);
nand U10536 (N_10536,N_10457,N_10329);
nand U10537 (N_10537,N_10306,N_10455);
and U10538 (N_10538,N_10474,N_10291);
nand U10539 (N_10539,N_10350,N_10280);
and U10540 (N_10540,N_10263,N_10389);
and U10541 (N_10541,N_10458,N_10432);
nand U10542 (N_10542,N_10303,N_10425);
or U10543 (N_10543,N_10299,N_10284);
or U10544 (N_10544,N_10486,N_10380);
nor U10545 (N_10545,N_10259,N_10487);
xnor U10546 (N_10546,N_10496,N_10465);
nor U10547 (N_10547,N_10480,N_10374);
nor U10548 (N_10548,N_10446,N_10429);
or U10549 (N_10549,N_10351,N_10287);
or U10550 (N_10550,N_10399,N_10288);
nor U10551 (N_10551,N_10261,N_10344);
or U10552 (N_10552,N_10449,N_10461);
nand U10553 (N_10553,N_10489,N_10309);
or U10554 (N_10554,N_10346,N_10312);
nand U10555 (N_10555,N_10450,N_10391);
nor U10556 (N_10556,N_10477,N_10407);
and U10557 (N_10557,N_10484,N_10393);
nor U10558 (N_10558,N_10311,N_10482);
nand U10559 (N_10559,N_10286,N_10268);
xnor U10560 (N_10560,N_10387,N_10297);
or U10561 (N_10561,N_10332,N_10276);
xor U10562 (N_10562,N_10293,N_10283);
or U10563 (N_10563,N_10378,N_10469);
xor U10564 (N_10564,N_10302,N_10485);
nor U10565 (N_10565,N_10292,N_10321);
xnor U10566 (N_10566,N_10468,N_10402);
nor U10567 (N_10567,N_10363,N_10390);
nor U10568 (N_10568,N_10337,N_10418);
or U10569 (N_10569,N_10318,N_10305);
or U10570 (N_10570,N_10392,N_10358);
nor U10571 (N_10571,N_10452,N_10423);
nor U10572 (N_10572,N_10257,N_10421);
and U10573 (N_10573,N_10479,N_10488);
and U10574 (N_10574,N_10414,N_10493);
nand U10575 (N_10575,N_10359,N_10319);
xor U10576 (N_10576,N_10385,N_10471);
or U10577 (N_10577,N_10258,N_10320);
nand U10578 (N_10578,N_10456,N_10300);
nor U10579 (N_10579,N_10499,N_10445);
or U10580 (N_10580,N_10381,N_10256);
nor U10581 (N_10581,N_10266,N_10361);
xor U10582 (N_10582,N_10347,N_10411);
nand U10583 (N_10583,N_10371,N_10372);
and U10584 (N_10584,N_10470,N_10466);
or U10585 (N_10585,N_10310,N_10376);
and U10586 (N_10586,N_10272,N_10314);
nand U10587 (N_10587,N_10322,N_10437);
or U10588 (N_10588,N_10324,N_10398);
or U10589 (N_10589,N_10345,N_10336);
or U10590 (N_10590,N_10325,N_10290);
and U10591 (N_10591,N_10459,N_10281);
xor U10592 (N_10592,N_10447,N_10304);
nor U10593 (N_10593,N_10255,N_10328);
and U10594 (N_10594,N_10419,N_10383);
nand U10595 (N_10595,N_10438,N_10335);
or U10596 (N_10596,N_10431,N_10370);
or U10597 (N_10597,N_10443,N_10454);
nor U10598 (N_10598,N_10494,N_10420);
nor U10599 (N_10599,N_10442,N_10491);
and U10600 (N_10600,N_10441,N_10326);
or U10601 (N_10601,N_10426,N_10317);
nand U10602 (N_10602,N_10436,N_10308);
nor U10603 (N_10603,N_10490,N_10424);
nor U10604 (N_10604,N_10439,N_10352);
and U10605 (N_10605,N_10404,N_10278);
xor U10606 (N_10606,N_10481,N_10375);
or U10607 (N_10607,N_10262,N_10277);
or U10608 (N_10608,N_10430,N_10251);
and U10609 (N_10609,N_10415,N_10295);
nand U10610 (N_10610,N_10428,N_10433);
nand U10611 (N_10611,N_10379,N_10353);
or U10612 (N_10612,N_10334,N_10331);
nand U10613 (N_10613,N_10354,N_10406);
or U10614 (N_10614,N_10264,N_10384);
nor U10615 (N_10615,N_10440,N_10405);
xor U10616 (N_10616,N_10313,N_10435);
xor U10617 (N_10617,N_10409,N_10340);
or U10618 (N_10618,N_10464,N_10338);
nor U10619 (N_10619,N_10366,N_10394);
and U10620 (N_10620,N_10401,N_10473);
nor U10621 (N_10621,N_10275,N_10497);
nand U10622 (N_10622,N_10413,N_10269);
or U10623 (N_10623,N_10434,N_10254);
and U10624 (N_10624,N_10348,N_10362);
and U10625 (N_10625,N_10329,N_10288);
or U10626 (N_10626,N_10361,N_10468);
nand U10627 (N_10627,N_10445,N_10335);
or U10628 (N_10628,N_10438,N_10280);
or U10629 (N_10629,N_10424,N_10471);
or U10630 (N_10630,N_10473,N_10355);
nand U10631 (N_10631,N_10262,N_10400);
and U10632 (N_10632,N_10488,N_10440);
nand U10633 (N_10633,N_10394,N_10261);
xnor U10634 (N_10634,N_10309,N_10284);
or U10635 (N_10635,N_10461,N_10318);
nor U10636 (N_10636,N_10275,N_10400);
nor U10637 (N_10637,N_10375,N_10406);
or U10638 (N_10638,N_10291,N_10330);
and U10639 (N_10639,N_10309,N_10304);
and U10640 (N_10640,N_10378,N_10465);
and U10641 (N_10641,N_10265,N_10413);
nand U10642 (N_10642,N_10309,N_10312);
nor U10643 (N_10643,N_10443,N_10344);
or U10644 (N_10644,N_10286,N_10294);
nor U10645 (N_10645,N_10259,N_10382);
nor U10646 (N_10646,N_10331,N_10349);
nor U10647 (N_10647,N_10325,N_10439);
nand U10648 (N_10648,N_10323,N_10314);
and U10649 (N_10649,N_10355,N_10346);
nor U10650 (N_10650,N_10452,N_10451);
and U10651 (N_10651,N_10271,N_10381);
nand U10652 (N_10652,N_10285,N_10454);
nor U10653 (N_10653,N_10437,N_10436);
nor U10654 (N_10654,N_10383,N_10276);
or U10655 (N_10655,N_10481,N_10401);
nand U10656 (N_10656,N_10333,N_10441);
or U10657 (N_10657,N_10456,N_10353);
and U10658 (N_10658,N_10438,N_10383);
xnor U10659 (N_10659,N_10386,N_10403);
nand U10660 (N_10660,N_10487,N_10352);
nor U10661 (N_10661,N_10320,N_10425);
or U10662 (N_10662,N_10342,N_10312);
or U10663 (N_10663,N_10412,N_10298);
nand U10664 (N_10664,N_10402,N_10276);
or U10665 (N_10665,N_10335,N_10430);
or U10666 (N_10666,N_10265,N_10289);
or U10667 (N_10667,N_10407,N_10386);
xor U10668 (N_10668,N_10479,N_10324);
or U10669 (N_10669,N_10354,N_10264);
nor U10670 (N_10670,N_10316,N_10371);
xnor U10671 (N_10671,N_10298,N_10382);
or U10672 (N_10672,N_10340,N_10270);
nand U10673 (N_10673,N_10477,N_10474);
nand U10674 (N_10674,N_10278,N_10334);
nor U10675 (N_10675,N_10346,N_10422);
or U10676 (N_10676,N_10486,N_10286);
or U10677 (N_10677,N_10364,N_10393);
or U10678 (N_10678,N_10436,N_10378);
nor U10679 (N_10679,N_10308,N_10310);
and U10680 (N_10680,N_10343,N_10479);
nand U10681 (N_10681,N_10446,N_10357);
and U10682 (N_10682,N_10261,N_10469);
or U10683 (N_10683,N_10356,N_10328);
and U10684 (N_10684,N_10360,N_10464);
and U10685 (N_10685,N_10271,N_10384);
and U10686 (N_10686,N_10271,N_10279);
nand U10687 (N_10687,N_10291,N_10449);
nand U10688 (N_10688,N_10281,N_10401);
nand U10689 (N_10689,N_10443,N_10416);
or U10690 (N_10690,N_10427,N_10368);
nand U10691 (N_10691,N_10442,N_10260);
or U10692 (N_10692,N_10332,N_10489);
or U10693 (N_10693,N_10411,N_10271);
nor U10694 (N_10694,N_10251,N_10426);
and U10695 (N_10695,N_10434,N_10377);
or U10696 (N_10696,N_10277,N_10358);
nor U10697 (N_10697,N_10435,N_10330);
and U10698 (N_10698,N_10404,N_10322);
and U10699 (N_10699,N_10438,N_10319);
and U10700 (N_10700,N_10383,N_10285);
nand U10701 (N_10701,N_10432,N_10402);
nand U10702 (N_10702,N_10390,N_10340);
or U10703 (N_10703,N_10394,N_10433);
nor U10704 (N_10704,N_10440,N_10295);
nand U10705 (N_10705,N_10258,N_10483);
nor U10706 (N_10706,N_10357,N_10252);
and U10707 (N_10707,N_10424,N_10383);
nor U10708 (N_10708,N_10446,N_10397);
xor U10709 (N_10709,N_10428,N_10364);
xnor U10710 (N_10710,N_10306,N_10347);
nand U10711 (N_10711,N_10292,N_10397);
nand U10712 (N_10712,N_10384,N_10466);
nor U10713 (N_10713,N_10311,N_10347);
xor U10714 (N_10714,N_10306,N_10370);
or U10715 (N_10715,N_10342,N_10439);
xnor U10716 (N_10716,N_10404,N_10317);
nor U10717 (N_10717,N_10499,N_10261);
or U10718 (N_10718,N_10485,N_10451);
or U10719 (N_10719,N_10267,N_10310);
and U10720 (N_10720,N_10482,N_10285);
and U10721 (N_10721,N_10291,N_10423);
and U10722 (N_10722,N_10301,N_10456);
nor U10723 (N_10723,N_10431,N_10373);
xor U10724 (N_10724,N_10393,N_10441);
nor U10725 (N_10725,N_10407,N_10400);
nor U10726 (N_10726,N_10258,N_10383);
or U10727 (N_10727,N_10364,N_10398);
or U10728 (N_10728,N_10337,N_10441);
nor U10729 (N_10729,N_10362,N_10307);
nor U10730 (N_10730,N_10418,N_10341);
nand U10731 (N_10731,N_10377,N_10455);
and U10732 (N_10732,N_10427,N_10280);
or U10733 (N_10733,N_10279,N_10394);
or U10734 (N_10734,N_10449,N_10414);
xor U10735 (N_10735,N_10275,N_10262);
nand U10736 (N_10736,N_10430,N_10305);
nand U10737 (N_10737,N_10417,N_10352);
and U10738 (N_10738,N_10488,N_10366);
xor U10739 (N_10739,N_10413,N_10261);
xnor U10740 (N_10740,N_10396,N_10329);
and U10741 (N_10741,N_10398,N_10322);
xor U10742 (N_10742,N_10417,N_10489);
nor U10743 (N_10743,N_10260,N_10305);
or U10744 (N_10744,N_10313,N_10492);
nand U10745 (N_10745,N_10305,N_10263);
nor U10746 (N_10746,N_10255,N_10374);
nor U10747 (N_10747,N_10274,N_10292);
or U10748 (N_10748,N_10444,N_10486);
xnor U10749 (N_10749,N_10287,N_10482);
nor U10750 (N_10750,N_10560,N_10570);
and U10751 (N_10751,N_10533,N_10547);
or U10752 (N_10752,N_10580,N_10718);
and U10753 (N_10753,N_10563,N_10701);
nand U10754 (N_10754,N_10623,N_10586);
nand U10755 (N_10755,N_10579,N_10581);
nand U10756 (N_10756,N_10531,N_10519);
and U10757 (N_10757,N_10738,N_10639);
nand U10758 (N_10758,N_10610,N_10642);
and U10759 (N_10759,N_10558,N_10515);
and U10760 (N_10760,N_10674,N_10611);
nand U10761 (N_10761,N_10554,N_10732);
nand U10762 (N_10762,N_10552,N_10575);
nand U10763 (N_10763,N_10544,N_10595);
and U10764 (N_10764,N_10619,N_10746);
or U10765 (N_10765,N_10528,N_10647);
nor U10766 (N_10766,N_10548,N_10524);
or U10767 (N_10767,N_10521,N_10724);
and U10768 (N_10768,N_10561,N_10540);
and U10769 (N_10769,N_10697,N_10733);
nor U10770 (N_10770,N_10512,N_10657);
and U10771 (N_10771,N_10664,N_10542);
nand U10772 (N_10772,N_10720,N_10740);
and U10773 (N_10773,N_10567,N_10603);
or U10774 (N_10774,N_10641,N_10582);
xor U10775 (N_10775,N_10666,N_10680);
nand U10776 (N_10776,N_10510,N_10714);
and U10777 (N_10777,N_10506,N_10559);
or U10778 (N_10778,N_10630,N_10659);
nor U10779 (N_10779,N_10646,N_10537);
and U10780 (N_10780,N_10728,N_10648);
and U10781 (N_10781,N_10652,N_10503);
and U10782 (N_10782,N_10587,N_10594);
nor U10783 (N_10783,N_10622,N_10711);
nor U10784 (N_10784,N_10520,N_10694);
and U10785 (N_10785,N_10629,N_10545);
nand U10786 (N_10786,N_10699,N_10716);
xnor U10787 (N_10787,N_10655,N_10574);
or U10788 (N_10788,N_10583,N_10693);
and U10789 (N_10789,N_10654,N_10690);
nor U10790 (N_10790,N_10549,N_10634);
or U10791 (N_10791,N_10597,N_10590);
xnor U10792 (N_10792,N_10627,N_10565);
nand U10793 (N_10793,N_10509,N_10741);
nand U10794 (N_10794,N_10593,N_10553);
or U10795 (N_10795,N_10538,N_10721);
or U10796 (N_10796,N_10650,N_10612);
and U10797 (N_10797,N_10566,N_10600);
xor U10798 (N_10798,N_10617,N_10747);
nand U10799 (N_10799,N_10722,N_10700);
xor U10800 (N_10800,N_10526,N_10516);
or U10801 (N_10801,N_10576,N_10673);
or U10802 (N_10802,N_10698,N_10504);
nand U10803 (N_10803,N_10692,N_10651);
nor U10804 (N_10804,N_10691,N_10726);
nor U10805 (N_10805,N_10735,N_10679);
nand U10806 (N_10806,N_10685,N_10705);
nand U10807 (N_10807,N_10522,N_10669);
and U10808 (N_10808,N_10745,N_10517);
nor U10809 (N_10809,N_10631,N_10686);
and U10810 (N_10810,N_10620,N_10536);
xor U10811 (N_10811,N_10681,N_10696);
and U10812 (N_10812,N_10736,N_10523);
nor U10813 (N_10813,N_10557,N_10719);
or U10814 (N_10814,N_10638,N_10500);
and U10815 (N_10815,N_10505,N_10507);
nor U10816 (N_10816,N_10602,N_10532);
and U10817 (N_10817,N_10573,N_10713);
nor U10818 (N_10818,N_10739,N_10535);
xnor U10819 (N_10819,N_10596,N_10725);
nor U10820 (N_10820,N_10584,N_10618);
nor U10821 (N_10821,N_10742,N_10605);
nor U10822 (N_10822,N_10637,N_10682);
nand U10823 (N_10823,N_10710,N_10550);
nor U10824 (N_10824,N_10723,N_10562);
xnor U10825 (N_10825,N_10684,N_10615);
nor U10826 (N_10826,N_10683,N_10546);
xor U10827 (N_10827,N_10644,N_10670);
and U10828 (N_10828,N_10555,N_10525);
nand U10829 (N_10829,N_10585,N_10571);
or U10830 (N_10830,N_10606,N_10708);
nor U10831 (N_10831,N_10727,N_10621);
and U10832 (N_10832,N_10633,N_10660);
and U10833 (N_10833,N_10530,N_10592);
nor U10834 (N_10834,N_10743,N_10663);
nor U10835 (N_10835,N_10707,N_10508);
or U10836 (N_10836,N_10599,N_10501);
or U10837 (N_10837,N_10632,N_10695);
nand U10838 (N_10838,N_10712,N_10613);
or U10839 (N_10839,N_10709,N_10676);
and U10840 (N_10840,N_10703,N_10628);
or U10841 (N_10841,N_10578,N_10672);
and U10842 (N_10842,N_10518,N_10729);
and U10843 (N_10843,N_10737,N_10706);
nor U10844 (N_10844,N_10588,N_10744);
or U10845 (N_10845,N_10529,N_10608);
or U10846 (N_10846,N_10704,N_10730);
and U10847 (N_10847,N_10625,N_10715);
or U10848 (N_10848,N_10572,N_10717);
and U10849 (N_10849,N_10748,N_10636);
nand U10850 (N_10850,N_10662,N_10564);
nand U10851 (N_10851,N_10607,N_10689);
nand U10852 (N_10852,N_10624,N_10502);
nor U10853 (N_10853,N_10658,N_10577);
or U10854 (N_10854,N_10635,N_10687);
or U10855 (N_10855,N_10551,N_10661);
xnor U10856 (N_10856,N_10527,N_10626);
nor U10857 (N_10857,N_10667,N_10749);
and U10858 (N_10858,N_10734,N_10569);
nor U10859 (N_10859,N_10556,N_10671);
or U10860 (N_10860,N_10616,N_10653);
and U10861 (N_10861,N_10702,N_10543);
xor U10862 (N_10862,N_10589,N_10640);
nand U10863 (N_10863,N_10668,N_10539);
and U10864 (N_10864,N_10614,N_10645);
or U10865 (N_10865,N_10678,N_10541);
nor U10866 (N_10866,N_10731,N_10675);
nor U10867 (N_10867,N_10568,N_10609);
or U10868 (N_10868,N_10604,N_10534);
and U10869 (N_10869,N_10591,N_10688);
nor U10870 (N_10870,N_10513,N_10601);
nand U10871 (N_10871,N_10598,N_10649);
and U10872 (N_10872,N_10643,N_10514);
nor U10873 (N_10873,N_10677,N_10656);
and U10874 (N_10874,N_10511,N_10665);
nand U10875 (N_10875,N_10644,N_10626);
nor U10876 (N_10876,N_10681,N_10652);
nor U10877 (N_10877,N_10532,N_10636);
nor U10878 (N_10878,N_10662,N_10529);
or U10879 (N_10879,N_10503,N_10628);
nor U10880 (N_10880,N_10561,N_10589);
nand U10881 (N_10881,N_10615,N_10679);
nand U10882 (N_10882,N_10716,N_10679);
or U10883 (N_10883,N_10665,N_10731);
xnor U10884 (N_10884,N_10725,N_10677);
nand U10885 (N_10885,N_10573,N_10602);
nor U10886 (N_10886,N_10529,N_10729);
nor U10887 (N_10887,N_10519,N_10593);
nor U10888 (N_10888,N_10559,N_10677);
nor U10889 (N_10889,N_10542,N_10585);
nand U10890 (N_10890,N_10549,N_10593);
or U10891 (N_10891,N_10582,N_10563);
or U10892 (N_10892,N_10591,N_10606);
or U10893 (N_10893,N_10509,N_10705);
and U10894 (N_10894,N_10559,N_10613);
nor U10895 (N_10895,N_10642,N_10584);
or U10896 (N_10896,N_10569,N_10749);
and U10897 (N_10897,N_10552,N_10507);
or U10898 (N_10898,N_10700,N_10601);
nor U10899 (N_10899,N_10749,N_10733);
or U10900 (N_10900,N_10546,N_10555);
and U10901 (N_10901,N_10614,N_10602);
nor U10902 (N_10902,N_10637,N_10664);
xor U10903 (N_10903,N_10657,N_10606);
nand U10904 (N_10904,N_10600,N_10636);
nor U10905 (N_10905,N_10587,N_10565);
nand U10906 (N_10906,N_10701,N_10689);
nor U10907 (N_10907,N_10698,N_10579);
or U10908 (N_10908,N_10726,N_10738);
nand U10909 (N_10909,N_10592,N_10656);
nand U10910 (N_10910,N_10735,N_10602);
xor U10911 (N_10911,N_10630,N_10679);
nor U10912 (N_10912,N_10631,N_10585);
nand U10913 (N_10913,N_10521,N_10503);
or U10914 (N_10914,N_10710,N_10603);
xor U10915 (N_10915,N_10508,N_10661);
xor U10916 (N_10916,N_10651,N_10740);
xor U10917 (N_10917,N_10597,N_10739);
or U10918 (N_10918,N_10622,N_10709);
nand U10919 (N_10919,N_10548,N_10525);
or U10920 (N_10920,N_10718,N_10614);
nor U10921 (N_10921,N_10711,N_10651);
xor U10922 (N_10922,N_10620,N_10700);
or U10923 (N_10923,N_10528,N_10505);
nor U10924 (N_10924,N_10682,N_10524);
nor U10925 (N_10925,N_10527,N_10590);
and U10926 (N_10926,N_10520,N_10718);
nand U10927 (N_10927,N_10506,N_10739);
nor U10928 (N_10928,N_10624,N_10581);
and U10929 (N_10929,N_10634,N_10678);
nor U10930 (N_10930,N_10544,N_10531);
nor U10931 (N_10931,N_10613,N_10664);
and U10932 (N_10932,N_10515,N_10532);
nand U10933 (N_10933,N_10677,N_10577);
nand U10934 (N_10934,N_10722,N_10627);
nand U10935 (N_10935,N_10581,N_10700);
nor U10936 (N_10936,N_10604,N_10560);
nand U10937 (N_10937,N_10591,N_10728);
nand U10938 (N_10938,N_10739,N_10595);
nor U10939 (N_10939,N_10716,N_10678);
nor U10940 (N_10940,N_10694,N_10571);
nand U10941 (N_10941,N_10557,N_10555);
nor U10942 (N_10942,N_10713,N_10575);
or U10943 (N_10943,N_10672,N_10511);
nor U10944 (N_10944,N_10749,N_10524);
or U10945 (N_10945,N_10726,N_10522);
nor U10946 (N_10946,N_10734,N_10713);
or U10947 (N_10947,N_10665,N_10622);
nand U10948 (N_10948,N_10566,N_10601);
xor U10949 (N_10949,N_10716,N_10645);
and U10950 (N_10950,N_10565,N_10559);
nand U10951 (N_10951,N_10612,N_10640);
nor U10952 (N_10952,N_10523,N_10508);
and U10953 (N_10953,N_10729,N_10697);
and U10954 (N_10954,N_10626,N_10628);
nand U10955 (N_10955,N_10501,N_10678);
nand U10956 (N_10956,N_10620,N_10709);
xor U10957 (N_10957,N_10609,N_10708);
and U10958 (N_10958,N_10525,N_10542);
nor U10959 (N_10959,N_10659,N_10599);
nand U10960 (N_10960,N_10736,N_10553);
nand U10961 (N_10961,N_10546,N_10509);
nor U10962 (N_10962,N_10545,N_10503);
nand U10963 (N_10963,N_10572,N_10728);
or U10964 (N_10964,N_10547,N_10544);
or U10965 (N_10965,N_10690,N_10682);
nand U10966 (N_10966,N_10561,N_10584);
and U10967 (N_10967,N_10713,N_10721);
nor U10968 (N_10968,N_10711,N_10598);
nor U10969 (N_10969,N_10667,N_10743);
or U10970 (N_10970,N_10657,N_10724);
nand U10971 (N_10971,N_10725,N_10745);
and U10972 (N_10972,N_10731,N_10576);
and U10973 (N_10973,N_10554,N_10612);
nor U10974 (N_10974,N_10561,N_10709);
or U10975 (N_10975,N_10749,N_10589);
nand U10976 (N_10976,N_10618,N_10635);
nor U10977 (N_10977,N_10699,N_10557);
nor U10978 (N_10978,N_10508,N_10620);
and U10979 (N_10979,N_10720,N_10690);
nand U10980 (N_10980,N_10702,N_10684);
nand U10981 (N_10981,N_10717,N_10592);
and U10982 (N_10982,N_10594,N_10560);
or U10983 (N_10983,N_10582,N_10748);
nor U10984 (N_10984,N_10676,N_10749);
or U10985 (N_10985,N_10691,N_10583);
xor U10986 (N_10986,N_10632,N_10533);
nand U10987 (N_10987,N_10631,N_10637);
and U10988 (N_10988,N_10694,N_10594);
or U10989 (N_10989,N_10542,N_10622);
and U10990 (N_10990,N_10510,N_10608);
xor U10991 (N_10991,N_10592,N_10744);
nand U10992 (N_10992,N_10526,N_10596);
or U10993 (N_10993,N_10570,N_10572);
nand U10994 (N_10994,N_10640,N_10577);
nor U10995 (N_10995,N_10636,N_10631);
nor U10996 (N_10996,N_10504,N_10683);
or U10997 (N_10997,N_10728,N_10743);
xor U10998 (N_10998,N_10508,N_10524);
and U10999 (N_10999,N_10617,N_10739);
nor U11000 (N_11000,N_10835,N_10774);
or U11001 (N_11001,N_10897,N_10798);
or U11002 (N_11002,N_10904,N_10843);
or U11003 (N_11003,N_10971,N_10969);
or U11004 (N_11004,N_10828,N_10803);
nor U11005 (N_11005,N_10787,N_10766);
nor U11006 (N_11006,N_10918,N_10764);
and U11007 (N_11007,N_10826,N_10955);
nand U11008 (N_11008,N_10895,N_10915);
nor U11009 (N_11009,N_10963,N_10861);
and U11010 (N_11010,N_10898,N_10778);
and U11011 (N_11011,N_10813,N_10867);
nor U11012 (N_11012,N_10773,N_10775);
and U11013 (N_11013,N_10769,N_10820);
nand U11014 (N_11014,N_10792,N_10929);
nor U11015 (N_11015,N_10967,N_10854);
or U11016 (N_11016,N_10964,N_10873);
or U11017 (N_11017,N_10819,N_10836);
nor U11018 (N_11018,N_10887,N_10882);
nand U11019 (N_11019,N_10881,N_10831);
nor U11020 (N_11020,N_10868,N_10757);
and U11021 (N_11021,N_10864,N_10900);
and U11022 (N_11022,N_10811,N_10932);
and U11023 (N_11023,N_10771,N_10890);
or U11024 (N_11024,N_10908,N_10834);
and U11025 (N_11025,N_10847,N_10916);
and U11026 (N_11026,N_10888,N_10917);
nand U11027 (N_11027,N_10911,N_10752);
or U11028 (N_11028,N_10842,N_10875);
nand U11029 (N_11029,N_10833,N_10782);
nor U11030 (N_11030,N_10808,N_10982);
or U11031 (N_11031,N_10956,N_10869);
and U11032 (N_11032,N_10844,N_10777);
or U11033 (N_11033,N_10905,N_10876);
and U11034 (N_11034,N_10935,N_10958);
nand U11035 (N_11035,N_10993,N_10800);
nor U11036 (N_11036,N_10959,N_10952);
and U11037 (N_11037,N_10756,N_10913);
and U11038 (N_11038,N_10906,N_10884);
xnor U11039 (N_11039,N_10767,N_10762);
xor U11040 (N_11040,N_10822,N_10791);
and U11041 (N_11041,N_10794,N_10957);
nand U11042 (N_11042,N_10933,N_10992);
or U11043 (N_11043,N_10863,N_10815);
nand U11044 (N_11044,N_10780,N_10907);
or U11045 (N_11045,N_10807,N_10901);
and U11046 (N_11046,N_10758,N_10928);
nand U11047 (N_11047,N_10997,N_10987);
nor U11048 (N_11048,N_10983,N_10856);
xnor U11049 (N_11049,N_10921,N_10995);
nor U11050 (N_11050,N_10806,N_10781);
nand U11051 (N_11051,N_10853,N_10872);
and U11052 (N_11052,N_10804,N_10974);
nand U11053 (N_11053,N_10972,N_10991);
and U11054 (N_11054,N_10981,N_10893);
nor U11055 (N_11055,N_10919,N_10862);
and U11056 (N_11056,N_10858,N_10903);
or U11057 (N_11057,N_10846,N_10943);
nand U11058 (N_11058,N_10816,N_10988);
or U11059 (N_11059,N_10899,N_10772);
nor U11060 (N_11060,N_10986,N_10962);
and U11061 (N_11061,N_10896,N_10785);
or U11062 (N_11062,N_10754,N_10937);
nor U11063 (N_11063,N_10924,N_10954);
nor U11064 (N_11064,N_10985,N_10759);
nor U11065 (N_11065,N_10852,N_10824);
nand U11066 (N_11066,N_10947,N_10878);
nand U11067 (N_11067,N_10855,N_10930);
or U11068 (N_11068,N_10920,N_10946);
or U11069 (N_11069,N_10953,N_10970);
or U11070 (N_11070,N_10949,N_10849);
and U11071 (N_11071,N_10980,N_10830);
or U11072 (N_11072,N_10945,N_10998);
nor U11073 (N_11073,N_10802,N_10796);
nor U11074 (N_11074,N_10942,N_10829);
xnor U11075 (N_11075,N_10977,N_10851);
nand U11076 (N_11076,N_10838,N_10776);
nand U11077 (N_11077,N_10886,N_10750);
nor U11078 (N_11078,N_10821,N_10944);
nor U11079 (N_11079,N_10818,N_10883);
nor U11080 (N_11080,N_10765,N_10927);
nand U11081 (N_11081,N_10914,N_10976);
and U11082 (N_11082,N_10910,N_10793);
xor U11083 (N_11083,N_10812,N_10809);
xor U11084 (N_11084,N_10832,N_10926);
or U11085 (N_11085,N_10984,N_10999);
nand U11086 (N_11086,N_10751,N_10790);
and U11087 (N_11087,N_10845,N_10990);
and U11088 (N_11088,N_10870,N_10841);
nand U11089 (N_11089,N_10940,N_10891);
nor U11090 (N_11090,N_10857,N_10966);
nand U11091 (N_11091,N_10892,N_10784);
nor U11092 (N_11092,N_10755,N_10837);
or U11093 (N_11093,N_10931,N_10839);
or U11094 (N_11094,N_10894,N_10939);
and U11095 (N_11095,N_10817,N_10961);
nand U11096 (N_11096,N_10871,N_10960);
or U11097 (N_11097,N_10951,N_10760);
or U11098 (N_11098,N_10934,N_10797);
nor U11099 (N_11099,N_10768,N_10779);
nor U11100 (N_11100,N_10877,N_10975);
nor U11101 (N_11101,N_10789,N_10799);
nor U11102 (N_11102,N_10860,N_10979);
nor U11103 (N_11103,N_10761,N_10825);
and U11104 (N_11104,N_10936,N_10938);
or U11105 (N_11105,N_10885,N_10879);
or U11106 (N_11106,N_10859,N_10770);
or U11107 (N_11107,N_10965,N_10989);
or U11108 (N_11108,N_10923,N_10948);
and U11109 (N_11109,N_10788,N_10810);
or U11110 (N_11110,N_10840,N_10848);
or U11111 (N_11111,N_10786,N_10889);
nand U11112 (N_11112,N_10973,N_10994);
or U11113 (N_11113,N_10941,N_10783);
nand U11114 (N_11114,N_10805,N_10880);
xor U11115 (N_11115,N_10823,N_10866);
nor U11116 (N_11116,N_10968,N_10950);
nand U11117 (N_11117,N_10801,N_10763);
and U11118 (N_11118,N_10827,N_10922);
nand U11119 (N_11119,N_10850,N_10902);
or U11120 (N_11120,N_10978,N_10753);
nand U11121 (N_11121,N_10925,N_10912);
and U11122 (N_11122,N_10996,N_10814);
or U11123 (N_11123,N_10795,N_10909);
nor U11124 (N_11124,N_10874,N_10865);
and U11125 (N_11125,N_10757,N_10876);
or U11126 (N_11126,N_10994,N_10887);
nor U11127 (N_11127,N_10846,N_10888);
nor U11128 (N_11128,N_10974,N_10931);
and U11129 (N_11129,N_10820,N_10886);
or U11130 (N_11130,N_10799,N_10897);
and U11131 (N_11131,N_10827,N_10840);
nand U11132 (N_11132,N_10758,N_10856);
xnor U11133 (N_11133,N_10905,N_10942);
nand U11134 (N_11134,N_10756,N_10892);
or U11135 (N_11135,N_10961,N_10758);
or U11136 (N_11136,N_10901,N_10782);
nand U11137 (N_11137,N_10922,N_10866);
nor U11138 (N_11138,N_10800,N_10791);
and U11139 (N_11139,N_10772,N_10914);
or U11140 (N_11140,N_10808,N_10965);
nand U11141 (N_11141,N_10907,N_10998);
nand U11142 (N_11142,N_10785,N_10979);
nand U11143 (N_11143,N_10929,N_10968);
and U11144 (N_11144,N_10877,N_10949);
and U11145 (N_11145,N_10901,N_10960);
and U11146 (N_11146,N_10893,N_10807);
nor U11147 (N_11147,N_10957,N_10972);
and U11148 (N_11148,N_10993,N_10919);
xnor U11149 (N_11149,N_10955,N_10805);
and U11150 (N_11150,N_10755,N_10855);
and U11151 (N_11151,N_10827,N_10886);
or U11152 (N_11152,N_10770,N_10785);
and U11153 (N_11153,N_10829,N_10821);
nor U11154 (N_11154,N_10786,N_10831);
xor U11155 (N_11155,N_10968,N_10935);
xor U11156 (N_11156,N_10910,N_10964);
nand U11157 (N_11157,N_10991,N_10852);
nand U11158 (N_11158,N_10774,N_10884);
nor U11159 (N_11159,N_10927,N_10878);
or U11160 (N_11160,N_10944,N_10894);
nand U11161 (N_11161,N_10966,N_10780);
nand U11162 (N_11162,N_10860,N_10750);
and U11163 (N_11163,N_10870,N_10863);
and U11164 (N_11164,N_10762,N_10761);
nand U11165 (N_11165,N_10979,N_10977);
xor U11166 (N_11166,N_10934,N_10909);
and U11167 (N_11167,N_10955,N_10834);
nand U11168 (N_11168,N_10938,N_10898);
nor U11169 (N_11169,N_10874,N_10843);
nand U11170 (N_11170,N_10872,N_10847);
nand U11171 (N_11171,N_10900,N_10887);
or U11172 (N_11172,N_10760,N_10941);
nor U11173 (N_11173,N_10893,N_10849);
and U11174 (N_11174,N_10879,N_10844);
and U11175 (N_11175,N_10972,N_10925);
or U11176 (N_11176,N_10969,N_10986);
and U11177 (N_11177,N_10765,N_10897);
nand U11178 (N_11178,N_10756,N_10781);
nand U11179 (N_11179,N_10781,N_10784);
and U11180 (N_11180,N_10758,N_10814);
and U11181 (N_11181,N_10779,N_10832);
nor U11182 (N_11182,N_10794,N_10844);
xor U11183 (N_11183,N_10849,N_10999);
nand U11184 (N_11184,N_10802,N_10819);
and U11185 (N_11185,N_10906,N_10890);
nor U11186 (N_11186,N_10778,N_10856);
and U11187 (N_11187,N_10848,N_10761);
nand U11188 (N_11188,N_10817,N_10969);
and U11189 (N_11189,N_10967,N_10836);
and U11190 (N_11190,N_10843,N_10842);
nor U11191 (N_11191,N_10811,N_10850);
or U11192 (N_11192,N_10922,N_10913);
nor U11193 (N_11193,N_10834,N_10968);
nor U11194 (N_11194,N_10996,N_10780);
nand U11195 (N_11195,N_10792,N_10750);
and U11196 (N_11196,N_10991,N_10950);
nor U11197 (N_11197,N_10836,N_10954);
nand U11198 (N_11198,N_10975,N_10758);
or U11199 (N_11199,N_10753,N_10781);
nand U11200 (N_11200,N_10898,N_10989);
or U11201 (N_11201,N_10804,N_10873);
or U11202 (N_11202,N_10779,N_10965);
or U11203 (N_11203,N_10760,N_10807);
and U11204 (N_11204,N_10936,N_10977);
and U11205 (N_11205,N_10970,N_10800);
nor U11206 (N_11206,N_10929,N_10899);
nand U11207 (N_11207,N_10880,N_10988);
and U11208 (N_11208,N_10819,N_10849);
nand U11209 (N_11209,N_10866,N_10790);
xnor U11210 (N_11210,N_10751,N_10762);
xor U11211 (N_11211,N_10839,N_10895);
or U11212 (N_11212,N_10776,N_10768);
nand U11213 (N_11213,N_10942,N_10830);
or U11214 (N_11214,N_10799,N_10752);
or U11215 (N_11215,N_10869,N_10788);
and U11216 (N_11216,N_10852,N_10856);
and U11217 (N_11217,N_10998,N_10986);
nor U11218 (N_11218,N_10976,N_10959);
nand U11219 (N_11219,N_10826,N_10768);
or U11220 (N_11220,N_10945,N_10777);
nand U11221 (N_11221,N_10931,N_10778);
and U11222 (N_11222,N_10983,N_10895);
nor U11223 (N_11223,N_10794,N_10837);
nor U11224 (N_11224,N_10973,N_10888);
nor U11225 (N_11225,N_10996,N_10906);
and U11226 (N_11226,N_10903,N_10864);
nor U11227 (N_11227,N_10976,N_10783);
nor U11228 (N_11228,N_10830,N_10796);
and U11229 (N_11229,N_10761,N_10921);
nand U11230 (N_11230,N_10766,N_10896);
nor U11231 (N_11231,N_10912,N_10932);
xor U11232 (N_11232,N_10871,N_10792);
and U11233 (N_11233,N_10943,N_10772);
nor U11234 (N_11234,N_10968,N_10998);
xnor U11235 (N_11235,N_10921,N_10868);
and U11236 (N_11236,N_10929,N_10844);
or U11237 (N_11237,N_10956,N_10789);
or U11238 (N_11238,N_10786,N_10973);
nor U11239 (N_11239,N_10752,N_10963);
xnor U11240 (N_11240,N_10971,N_10810);
or U11241 (N_11241,N_10872,N_10989);
or U11242 (N_11242,N_10964,N_10871);
nor U11243 (N_11243,N_10953,N_10980);
xor U11244 (N_11244,N_10955,N_10818);
and U11245 (N_11245,N_10889,N_10894);
nand U11246 (N_11246,N_10963,N_10927);
nor U11247 (N_11247,N_10825,N_10983);
nand U11248 (N_11248,N_10915,N_10937);
nand U11249 (N_11249,N_10785,N_10823);
and U11250 (N_11250,N_11196,N_11003);
nor U11251 (N_11251,N_11051,N_11249);
and U11252 (N_11252,N_11229,N_11123);
xnor U11253 (N_11253,N_11060,N_11248);
and U11254 (N_11254,N_11234,N_11041);
nand U11255 (N_11255,N_11243,N_11087);
or U11256 (N_11256,N_11077,N_11108);
nor U11257 (N_11257,N_11138,N_11109);
and U11258 (N_11258,N_11068,N_11223);
and U11259 (N_11259,N_11105,N_11094);
or U11260 (N_11260,N_11128,N_11129);
nor U11261 (N_11261,N_11042,N_11029);
nor U11262 (N_11262,N_11066,N_11119);
or U11263 (N_11263,N_11165,N_11074);
and U11264 (N_11264,N_11048,N_11011);
nor U11265 (N_11265,N_11148,N_11175);
or U11266 (N_11266,N_11132,N_11233);
or U11267 (N_11267,N_11019,N_11155);
nand U11268 (N_11268,N_11047,N_11080);
xor U11269 (N_11269,N_11036,N_11215);
xor U11270 (N_11270,N_11247,N_11143);
and U11271 (N_11271,N_11067,N_11001);
and U11272 (N_11272,N_11224,N_11020);
xnor U11273 (N_11273,N_11059,N_11065);
or U11274 (N_11274,N_11056,N_11179);
or U11275 (N_11275,N_11151,N_11133);
and U11276 (N_11276,N_11070,N_11016);
or U11277 (N_11277,N_11153,N_11122);
nor U11278 (N_11278,N_11012,N_11021);
and U11279 (N_11279,N_11236,N_11171);
nand U11280 (N_11280,N_11189,N_11045);
nor U11281 (N_11281,N_11213,N_11192);
and U11282 (N_11282,N_11219,N_11194);
nor U11283 (N_11283,N_11208,N_11046);
and U11284 (N_11284,N_11174,N_11025);
xnor U11285 (N_11285,N_11071,N_11052);
nand U11286 (N_11286,N_11135,N_11217);
nand U11287 (N_11287,N_11100,N_11187);
nor U11288 (N_11288,N_11050,N_11076);
and U11289 (N_11289,N_11164,N_11026);
nand U11290 (N_11290,N_11203,N_11034);
or U11291 (N_11291,N_11211,N_11005);
nand U11292 (N_11292,N_11043,N_11134);
and U11293 (N_11293,N_11140,N_11239);
nor U11294 (N_11294,N_11181,N_11144);
nand U11295 (N_11295,N_11141,N_11009);
nand U11296 (N_11296,N_11010,N_11082);
nor U11297 (N_11297,N_11202,N_11245);
nand U11298 (N_11298,N_11062,N_11168);
or U11299 (N_11299,N_11089,N_11201);
nor U11300 (N_11300,N_11107,N_11205);
and U11301 (N_11301,N_11156,N_11055);
and U11302 (N_11302,N_11013,N_11083);
and U11303 (N_11303,N_11182,N_11014);
nand U11304 (N_11304,N_11147,N_11235);
nand U11305 (N_11305,N_11091,N_11081);
nand U11306 (N_11306,N_11183,N_11112);
or U11307 (N_11307,N_11125,N_11212);
nand U11308 (N_11308,N_11096,N_11173);
nor U11309 (N_11309,N_11024,N_11238);
or U11310 (N_11310,N_11064,N_11007);
and U11311 (N_11311,N_11149,N_11127);
nand U11312 (N_11312,N_11113,N_11210);
xnor U11313 (N_11313,N_11162,N_11220);
xor U11314 (N_11314,N_11161,N_11184);
or U11315 (N_11315,N_11037,N_11090);
nand U11316 (N_11316,N_11028,N_11114);
or U11317 (N_11317,N_11057,N_11242);
xor U11318 (N_11318,N_11004,N_11118);
or U11319 (N_11319,N_11126,N_11111);
nor U11320 (N_11320,N_11098,N_11102);
xnor U11321 (N_11321,N_11008,N_11216);
and U11322 (N_11322,N_11237,N_11244);
nand U11323 (N_11323,N_11150,N_11241);
or U11324 (N_11324,N_11157,N_11185);
nor U11325 (N_11325,N_11204,N_11000);
or U11326 (N_11326,N_11172,N_11200);
xnor U11327 (N_11327,N_11103,N_11191);
and U11328 (N_11328,N_11033,N_11088);
nor U11329 (N_11329,N_11221,N_11079);
xor U11330 (N_11330,N_11228,N_11222);
xnor U11331 (N_11331,N_11032,N_11058);
or U11332 (N_11332,N_11137,N_11152);
nand U11333 (N_11333,N_11063,N_11085);
nand U11334 (N_11334,N_11193,N_11017);
xnor U11335 (N_11335,N_11110,N_11044);
and U11336 (N_11336,N_11023,N_11231);
nor U11337 (N_11337,N_11053,N_11073);
nand U11338 (N_11338,N_11158,N_11084);
and U11339 (N_11339,N_11131,N_11031);
nor U11340 (N_11340,N_11095,N_11054);
or U11341 (N_11341,N_11145,N_11142);
nor U11342 (N_11342,N_11022,N_11092);
xor U11343 (N_11343,N_11186,N_11136);
nand U11344 (N_11344,N_11195,N_11104);
nor U11345 (N_11345,N_11072,N_11206);
nor U11346 (N_11346,N_11099,N_11188);
nor U11347 (N_11347,N_11207,N_11086);
nor U11348 (N_11348,N_11078,N_11115);
nor U11349 (N_11349,N_11146,N_11121);
xnor U11350 (N_11350,N_11075,N_11209);
or U11351 (N_11351,N_11169,N_11199);
and U11352 (N_11352,N_11176,N_11097);
and U11353 (N_11353,N_11240,N_11035);
and U11354 (N_11354,N_11178,N_11160);
nor U11355 (N_11355,N_11232,N_11166);
or U11356 (N_11356,N_11139,N_11226);
or U11357 (N_11357,N_11177,N_11198);
nor U11358 (N_11358,N_11163,N_11230);
nor U11359 (N_11359,N_11039,N_11018);
xor U11360 (N_11360,N_11061,N_11101);
and U11361 (N_11361,N_11225,N_11027);
nand U11362 (N_11362,N_11038,N_11117);
and U11363 (N_11363,N_11116,N_11170);
or U11364 (N_11364,N_11006,N_11106);
xnor U11365 (N_11365,N_11124,N_11214);
xor U11366 (N_11366,N_11069,N_11197);
nor U11367 (N_11367,N_11167,N_11049);
nand U11368 (N_11368,N_11159,N_11218);
nand U11369 (N_11369,N_11227,N_11120);
nand U11370 (N_11370,N_11030,N_11002);
and U11371 (N_11371,N_11040,N_11154);
nand U11372 (N_11372,N_11246,N_11190);
nor U11373 (N_11373,N_11130,N_11015);
and U11374 (N_11374,N_11180,N_11093);
and U11375 (N_11375,N_11013,N_11018);
xor U11376 (N_11376,N_11096,N_11222);
or U11377 (N_11377,N_11006,N_11169);
or U11378 (N_11378,N_11053,N_11249);
nor U11379 (N_11379,N_11010,N_11095);
xnor U11380 (N_11380,N_11173,N_11054);
nor U11381 (N_11381,N_11160,N_11173);
nand U11382 (N_11382,N_11213,N_11011);
nor U11383 (N_11383,N_11200,N_11189);
nor U11384 (N_11384,N_11218,N_11053);
nor U11385 (N_11385,N_11025,N_11016);
xor U11386 (N_11386,N_11044,N_11204);
and U11387 (N_11387,N_11132,N_11244);
xnor U11388 (N_11388,N_11095,N_11062);
xor U11389 (N_11389,N_11208,N_11232);
nor U11390 (N_11390,N_11100,N_11193);
nor U11391 (N_11391,N_11175,N_11095);
or U11392 (N_11392,N_11244,N_11161);
and U11393 (N_11393,N_11237,N_11151);
nor U11394 (N_11394,N_11061,N_11007);
nor U11395 (N_11395,N_11248,N_11005);
nor U11396 (N_11396,N_11023,N_11041);
xor U11397 (N_11397,N_11182,N_11238);
or U11398 (N_11398,N_11077,N_11097);
and U11399 (N_11399,N_11072,N_11052);
nand U11400 (N_11400,N_11117,N_11154);
and U11401 (N_11401,N_11004,N_11207);
and U11402 (N_11402,N_11024,N_11152);
or U11403 (N_11403,N_11211,N_11043);
nor U11404 (N_11404,N_11232,N_11117);
or U11405 (N_11405,N_11095,N_11161);
and U11406 (N_11406,N_11088,N_11124);
nor U11407 (N_11407,N_11224,N_11002);
or U11408 (N_11408,N_11121,N_11249);
or U11409 (N_11409,N_11095,N_11101);
or U11410 (N_11410,N_11070,N_11166);
nand U11411 (N_11411,N_11035,N_11091);
or U11412 (N_11412,N_11197,N_11136);
nand U11413 (N_11413,N_11061,N_11051);
nor U11414 (N_11414,N_11079,N_11145);
nand U11415 (N_11415,N_11120,N_11050);
nand U11416 (N_11416,N_11131,N_11065);
nand U11417 (N_11417,N_11187,N_11103);
and U11418 (N_11418,N_11037,N_11117);
or U11419 (N_11419,N_11132,N_11217);
nand U11420 (N_11420,N_11200,N_11019);
nand U11421 (N_11421,N_11006,N_11124);
or U11422 (N_11422,N_11010,N_11168);
nand U11423 (N_11423,N_11026,N_11065);
nand U11424 (N_11424,N_11102,N_11219);
nor U11425 (N_11425,N_11119,N_11166);
and U11426 (N_11426,N_11166,N_11197);
and U11427 (N_11427,N_11141,N_11027);
and U11428 (N_11428,N_11128,N_11088);
nand U11429 (N_11429,N_11052,N_11138);
and U11430 (N_11430,N_11153,N_11093);
or U11431 (N_11431,N_11199,N_11099);
nor U11432 (N_11432,N_11045,N_11081);
and U11433 (N_11433,N_11247,N_11075);
nor U11434 (N_11434,N_11213,N_11194);
and U11435 (N_11435,N_11176,N_11078);
or U11436 (N_11436,N_11016,N_11108);
or U11437 (N_11437,N_11234,N_11017);
and U11438 (N_11438,N_11022,N_11053);
nor U11439 (N_11439,N_11174,N_11044);
xor U11440 (N_11440,N_11159,N_11115);
nand U11441 (N_11441,N_11233,N_11106);
nor U11442 (N_11442,N_11124,N_11130);
and U11443 (N_11443,N_11237,N_11009);
nor U11444 (N_11444,N_11070,N_11064);
and U11445 (N_11445,N_11091,N_11075);
nor U11446 (N_11446,N_11172,N_11142);
and U11447 (N_11447,N_11091,N_11167);
or U11448 (N_11448,N_11190,N_11152);
nand U11449 (N_11449,N_11022,N_11018);
or U11450 (N_11450,N_11169,N_11237);
and U11451 (N_11451,N_11235,N_11038);
nand U11452 (N_11452,N_11127,N_11007);
or U11453 (N_11453,N_11146,N_11163);
and U11454 (N_11454,N_11028,N_11122);
and U11455 (N_11455,N_11074,N_11225);
and U11456 (N_11456,N_11103,N_11243);
or U11457 (N_11457,N_11009,N_11226);
nor U11458 (N_11458,N_11174,N_11169);
or U11459 (N_11459,N_11088,N_11096);
xor U11460 (N_11460,N_11246,N_11238);
or U11461 (N_11461,N_11205,N_11092);
or U11462 (N_11462,N_11028,N_11226);
or U11463 (N_11463,N_11211,N_11210);
or U11464 (N_11464,N_11126,N_11142);
xnor U11465 (N_11465,N_11011,N_11168);
or U11466 (N_11466,N_11215,N_11002);
nor U11467 (N_11467,N_11073,N_11088);
nor U11468 (N_11468,N_11141,N_11056);
or U11469 (N_11469,N_11044,N_11079);
or U11470 (N_11470,N_11126,N_11081);
or U11471 (N_11471,N_11108,N_11167);
nor U11472 (N_11472,N_11015,N_11071);
or U11473 (N_11473,N_11029,N_11226);
nor U11474 (N_11474,N_11075,N_11016);
nand U11475 (N_11475,N_11100,N_11077);
xnor U11476 (N_11476,N_11186,N_11153);
or U11477 (N_11477,N_11201,N_11046);
xor U11478 (N_11478,N_11180,N_11035);
nand U11479 (N_11479,N_11111,N_11206);
or U11480 (N_11480,N_11151,N_11192);
or U11481 (N_11481,N_11024,N_11164);
and U11482 (N_11482,N_11118,N_11149);
nor U11483 (N_11483,N_11153,N_11034);
nand U11484 (N_11484,N_11243,N_11062);
nor U11485 (N_11485,N_11013,N_11107);
or U11486 (N_11486,N_11187,N_11088);
nor U11487 (N_11487,N_11206,N_11229);
or U11488 (N_11488,N_11247,N_11079);
nand U11489 (N_11489,N_11207,N_11144);
nor U11490 (N_11490,N_11140,N_11117);
or U11491 (N_11491,N_11028,N_11218);
and U11492 (N_11492,N_11163,N_11187);
nand U11493 (N_11493,N_11103,N_11156);
nand U11494 (N_11494,N_11059,N_11137);
or U11495 (N_11495,N_11171,N_11046);
nand U11496 (N_11496,N_11213,N_11035);
nor U11497 (N_11497,N_11110,N_11135);
or U11498 (N_11498,N_11063,N_11228);
and U11499 (N_11499,N_11067,N_11194);
nand U11500 (N_11500,N_11445,N_11327);
nor U11501 (N_11501,N_11304,N_11387);
nor U11502 (N_11502,N_11410,N_11282);
nand U11503 (N_11503,N_11310,N_11415);
and U11504 (N_11504,N_11260,N_11442);
and U11505 (N_11505,N_11276,N_11389);
nand U11506 (N_11506,N_11396,N_11308);
or U11507 (N_11507,N_11429,N_11272);
nor U11508 (N_11508,N_11340,N_11256);
nor U11509 (N_11509,N_11373,N_11388);
nor U11510 (N_11510,N_11288,N_11400);
nand U11511 (N_11511,N_11265,N_11252);
nor U11512 (N_11512,N_11314,N_11458);
or U11513 (N_11513,N_11324,N_11376);
nand U11514 (N_11514,N_11253,N_11379);
nor U11515 (N_11515,N_11422,N_11286);
nand U11516 (N_11516,N_11451,N_11417);
xnor U11517 (N_11517,N_11386,N_11341);
or U11518 (N_11518,N_11457,N_11478);
nor U11519 (N_11519,N_11266,N_11473);
nor U11520 (N_11520,N_11366,N_11362);
nor U11521 (N_11521,N_11274,N_11433);
or U11522 (N_11522,N_11295,N_11330);
nand U11523 (N_11523,N_11438,N_11497);
nor U11524 (N_11524,N_11254,N_11323);
or U11525 (N_11525,N_11350,N_11412);
nor U11526 (N_11526,N_11358,N_11494);
or U11527 (N_11527,N_11405,N_11292);
or U11528 (N_11528,N_11461,N_11313);
nand U11529 (N_11529,N_11480,N_11434);
nand U11530 (N_11530,N_11481,N_11432);
nor U11531 (N_11531,N_11264,N_11296);
nand U11532 (N_11532,N_11431,N_11482);
nor U11533 (N_11533,N_11468,N_11331);
and U11534 (N_11534,N_11407,N_11294);
nand U11535 (N_11535,N_11290,N_11428);
or U11536 (N_11536,N_11479,N_11498);
xnor U11537 (N_11537,N_11333,N_11332);
nand U11538 (N_11538,N_11357,N_11441);
or U11539 (N_11539,N_11287,N_11409);
nand U11540 (N_11540,N_11278,N_11289);
nor U11541 (N_11541,N_11477,N_11488);
xnor U11542 (N_11542,N_11349,N_11370);
and U11543 (N_11543,N_11444,N_11420);
or U11544 (N_11544,N_11413,N_11305);
and U11545 (N_11545,N_11427,N_11462);
or U11546 (N_11546,N_11275,N_11382);
and U11547 (N_11547,N_11401,N_11408);
or U11548 (N_11548,N_11476,N_11414);
or U11549 (N_11549,N_11336,N_11467);
and U11550 (N_11550,N_11423,N_11365);
nor U11551 (N_11551,N_11418,N_11353);
and U11552 (N_11552,N_11262,N_11369);
or U11553 (N_11553,N_11377,N_11250);
or U11554 (N_11554,N_11281,N_11368);
and U11555 (N_11555,N_11328,N_11380);
and U11556 (N_11556,N_11465,N_11348);
or U11557 (N_11557,N_11321,N_11391);
xor U11558 (N_11558,N_11483,N_11364);
or U11559 (N_11559,N_11449,N_11251);
and U11560 (N_11560,N_11472,N_11440);
nand U11561 (N_11561,N_11454,N_11471);
and U11562 (N_11562,N_11456,N_11463);
nor U11563 (N_11563,N_11485,N_11335);
nand U11564 (N_11564,N_11312,N_11325);
or U11565 (N_11565,N_11398,N_11383);
and U11566 (N_11566,N_11402,N_11273);
nand U11567 (N_11567,N_11326,N_11351);
or U11568 (N_11568,N_11371,N_11303);
and U11569 (N_11569,N_11342,N_11355);
and U11570 (N_11570,N_11270,N_11437);
and U11571 (N_11571,N_11404,N_11311);
nand U11572 (N_11572,N_11384,N_11318);
nor U11573 (N_11573,N_11393,N_11363);
xor U11574 (N_11574,N_11285,N_11315);
nor U11575 (N_11575,N_11334,N_11446);
and U11576 (N_11576,N_11470,N_11347);
nor U11577 (N_11577,N_11421,N_11359);
nor U11578 (N_11578,N_11424,N_11487);
and U11579 (N_11579,N_11302,N_11263);
nand U11580 (N_11580,N_11392,N_11399);
nand U11581 (N_11581,N_11416,N_11474);
and U11582 (N_11582,N_11490,N_11435);
or U11583 (N_11583,N_11259,N_11492);
nor U11584 (N_11584,N_11269,N_11352);
xnor U11585 (N_11585,N_11280,N_11301);
or U11586 (N_11586,N_11299,N_11374);
or U11587 (N_11587,N_11447,N_11367);
xor U11588 (N_11588,N_11452,N_11279);
and U11589 (N_11589,N_11258,N_11453);
and U11590 (N_11590,N_11450,N_11339);
nand U11591 (N_11591,N_11356,N_11493);
nand U11592 (N_11592,N_11425,N_11329);
nand U11593 (N_11593,N_11344,N_11277);
and U11594 (N_11594,N_11464,N_11489);
or U11595 (N_11595,N_11390,N_11496);
or U11596 (N_11596,N_11411,N_11257);
or U11597 (N_11597,N_11439,N_11338);
nand U11598 (N_11598,N_11406,N_11309);
or U11599 (N_11599,N_11475,N_11316);
nand U11600 (N_11600,N_11271,N_11378);
and U11601 (N_11601,N_11306,N_11322);
or U11602 (N_11602,N_11486,N_11298);
nand U11603 (N_11603,N_11343,N_11419);
and U11604 (N_11604,N_11495,N_11261);
and U11605 (N_11605,N_11372,N_11268);
xnor U11606 (N_11606,N_11443,N_11267);
or U11607 (N_11607,N_11300,N_11346);
nor U11608 (N_11608,N_11337,N_11491);
nand U11609 (N_11609,N_11381,N_11283);
xnor U11610 (N_11610,N_11361,N_11395);
nor U11611 (N_11611,N_11255,N_11307);
nand U11612 (N_11612,N_11499,N_11459);
xnor U11613 (N_11613,N_11385,N_11345);
nor U11614 (N_11614,N_11466,N_11360);
nor U11615 (N_11615,N_11291,N_11469);
or U11616 (N_11616,N_11354,N_11484);
or U11617 (N_11617,N_11436,N_11455);
nand U11618 (N_11618,N_11448,N_11317);
and U11619 (N_11619,N_11297,N_11426);
and U11620 (N_11620,N_11430,N_11403);
nand U11621 (N_11621,N_11320,N_11375);
nand U11622 (N_11622,N_11319,N_11394);
or U11623 (N_11623,N_11284,N_11460);
nand U11624 (N_11624,N_11397,N_11293);
nor U11625 (N_11625,N_11323,N_11334);
and U11626 (N_11626,N_11336,N_11448);
xnor U11627 (N_11627,N_11287,N_11411);
or U11628 (N_11628,N_11388,N_11307);
and U11629 (N_11629,N_11306,N_11258);
nand U11630 (N_11630,N_11371,N_11343);
nand U11631 (N_11631,N_11486,N_11301);
nand U11632 (N_11632,N_11476,N_11490);
nand U11633 (N_11633,N_11322,N_11315);
and U11634 (N_11634,N_11274,N_11422);
nor U11635 (N_11635,N_11410,N_11340);
and U11636 (N_11636,N_11314,N_11486);
and U11637 (N_11637,N_11437,N_11367);
and U11638 (N_11638,N_11486,N_11395);
nor U11639 (N_11639,N_11361,N_11365);
and U11640 (N_11640,N_11253,N_11366);
xnor U11641 (N_11641,N_11455,N_11345);
xor U11642 (N_11642,N_11262,N_11405);
nand U11643 (N_11643,N_11367,N_11456);
nand U11644 (N_11644,N_11434,N_11419);
or U11645 (N_11645,N_11399,N_11262);
nor U11646 (N_11646,N_11479,N_11390);
nor U11647 (N_11647,N_11251,N_11253);
and U11648 (N_11648,N_11253,N_11304);
nand U11649 (N_11649,N_11303,N_11412);
xor U11650 (N_11650,N_11268,N_11287);
xnor U11651 (N_11651,N_11295,N_11344);
xnor U11652 (N_11652,N_11291,N_11394);
nand U11653 (N_11653,N_11425,N_11309);
or U11654 (N_11654,N_11492,N_11289);
nor U11655 (N_11655,N_11307,N_11276);
nand U11656 (N_11656,N_11373,N_11484);
xnor U11657 (N_11657,N_11263,N_11448);
xor U11658 (N_11658,N_11256,N_11319);
nor U11659 (N_11659,N_11275,N_11251);
or U11660 (N_11660,N_11349,N_11352);
nand U11661 (N_11661,N_11335,N_11326);
xnor U11662 (N_11662,N_11350,N_11438);
nand U11663 (N_11663,N_11471,N_11421);
or U11664 (N_11664,N_11340,N_11420);
or U11665 (N_11665,N_11377,N_11302);
or U11666 (N_11666,N_11253,N_11387);
or U11667 (N_11667,N_11272,N_11252);
xnor U11668 (N_11668,N_11420,N_11455);
and U11669 (N_11669,N_11350,N_11483);
xor U11670 (N_11670,N_11433,N_11364);
or U11671 (N_11671,N_11496,N_11336);
nor U11672 (N_11672,N_11466,N_11401);
and U11673 (N_11673,N_11408,N_11375);
nor U11674 (N_11674,N_11320,N_11417);
nand U11675 (N_11675,N_11390,N_11363);
and U11676 (N_11676,N_11416,N_11396);
nand U11677 (N_11677,N_11373,N_11347);
and U11678 (N_11678,N_11268,N_11432);
xor U11679 (N_11679,N_11345,N_11257);
and U11680 (N_11680,N_11290,N_11274);
xnor U11681 (N_11681,N_11444,N_11429);
or U11682 (N_11682,N_11350,N_11470);
and U11683 (N_11683,N_11312,N_11251);
nor U11684 (N_11684,N_11272,N_11473);
nor U11685 (N_11685,N_11336,N_11418);
and U11686 (N_11686,N_11267,N_11357);
nor U11687 (N_11687,N_11347,N_11422);
nand U11688 (N_11688,N_11483,N_11424);
or U11689 (N_11689,N_11450,N_11371);
nand U11690 (N_11690,N_11286,N_11335);
and U11691 (N_11691,N_11455,N_11400);
xnor U11692 (N_11692,N_11401,N_11428);
nor U11693 (N_11693,N_11473,N_11330);
and U11694 (N_11694,N_11372,N_11330);
nor U11695 (N_11695,N_11398,N_11333);
nor U11696 (N_11696,N_11356,N_11440);
or U11697 (N_11697,N_11308,N_11397);
nor U11698 (N_11698,N_11394,N_11276);
nor U11699 (N_11699,N_11460,N_11391);
nor U11700 (N_11700,N_11335,N_11266);
or U11701 (N_11701,N_11412,N_11405);
and U11702 (N_11702,N_11423,N_11447);
or U11703 (N_11703,N_11487,N_11430);
or U11704 (N_11704,N_11278,N_11298);
or U11705 (N_11705,N_11295,N_11419);
and U11706 (N_11706,N_11319,N_11367);
nand U11707 (N_11707,N_11456,N_11341);
or U11708 (N_11708,N_11480,N_11423);
nor U11709 (N_11709,N_11487,N_11476);
nand U11710 (N_11710,N_11468,N_11362);
nand U11711 (N_11711,N_11339,N_11348);
nor U11712 (N_11712,N_11447,N_11468);
nand U11713 (N_11713,N_11389,N_11440);
and U11714 (N_11714,N_11459,N_11273);
nand U11715 (N_11715,N_11294,N_11455);
or U11716 (N_11716,N_11366,N_11495);
nand U11717 (N_11717,N_11428,N_11268);
xnor U11718 (N_11718,N_11498,N_11432);
xnor U11719 (N_11719,N_11499,N_11259);
and U11720 (N_11720,N_11293,N_11352);
nor U11721 (N_11721,N_11408,N_11299);
or U11722 (N_11722,N_11456,N_11350);
or U11723 (N_11723,N_11314,N_11464);
nand U11724 (N_11724,N_11389,N_11272);
and U11725 (N_11725,N_11470,N_11403);
or U11726 (N_11726,N_11421,N_11483);
nand U11727 (N_11727,N_11427,N_11423);
or U11728 (N_11728,N_11475,N_11297);
and U11729 (N_11729,N_11473,N_11491);
nand U11730 (N_11730,N_11273,N_11494);
nand U11731 (N_11731,N_11340,N_11489);
nor U11732 (N_11732,N_11270,N_11325);
xnor U11733 (N_11733,N_11438,N_11370);
or U11734 (N_11734,N_11418,N_11470);
nand U11735 (N_11735,N_11364,N_11294);
nand U11736 (N_11736,N_11363,N_11414);
nor U11737 (N_11737,N_11498,N_11340);
nor U11738 (N_11738,N_11254,N_11318);
or U11739 (N_11739,N_11399,N_11309);
and U11740 (N_11740,N_11285,N_11292);
xnor U11741 (N_11741,N_11435,N_11426);
nand U11742 (N_11742,N_11477,N_11384);
nor U11743 (N_11743,N_11445,N_11452);
nor U11744 (N_11744,N_11301,N_11319);
nand U11745 (N_11745,N_11382,N_11324);
and U11746 (N_11746,N_11257,N_11404);
nor U11747 (N_11747,N_11324,N_11283);
nand U11748 (N_11748,N_11325,N_11267);
or U11749 (N_11749,N_11444,N_11474);
xnor U11750 (N_11750,N_11561,N_11552);
or U11751 (N_11751,N_11513,N_11709);
nor U11752 (N_11752,N_11586,N_11651);
nand U11753 (N_11753,N_11705,N_11596);
nor U11754 (N_11754,N_11643,N_11687);
nand U11755 (N_11755,N_11637,N_11531);
or U11756 (N_11756,N_11517,N_11731);
and U11757 (N_11757,N_11623,N_11524);
and U11758 (N_11758,N_11663,N_11676);
nand U11759 (N_11759,N_11630,N_11656);
nor U11760 (N_11760,N_11591,N_11512);
nand U11761 (N_11761,N_11657,N_11523);
and U11762 (N_11762,N_11723,N_11600);
or U11763 (N_11763,N_11617,N_11627);
nor U11764 (N_11764,N_11710,N_11638);
or U11765 (N_11765,N_11572,N_11641);
or U11766 (N_11766,N_11511,N_11587);
or U11767 (N_11767,N_11539,N_11615);
nand U11768 (N_11768,N_11554,N_11717);
nand U11769 (N_11769,N_11607,N_11648);
or U11770 (N_11770,N_11509,N_11741);
and U11771 (N_11771,N_11556,N_11721);
or U11772 (N_11772,N_11722,N_11635);
or U11773 (N_11773,N_11730,N_11749);
nand U11774 (N_11774,N_11739,N_11745);
or U11775 (N_11775,N_11661,N_11677);
or U11776 (N_11776,N_11646,N_11619);
nand U11777 (N_11777,N_11604,N_11550);
or U11778 (N_11778,N_11534,N_11580);
nor U11779 (N_11779,N_11589,N_11634);
or U11780 (N_11780,N_11636,N_11503);
or U11781 (N_11781,N_11658,N_11695);
nand U11782 (N_11782,N_11538,N_11598);
and U11783 (N_11783,N_11674,N_11558);
nand U11784 (N_11784,N_11546,N_11733);
and U11785 (N_11785,N_11563,N_11685);
nand U11786 (N_11786,N_11704,N_11715);
nand U11787 (N_11787,N_11675,N_11662);
and U11788 (N_11788,N_11545,N_11644);
xnor U11789 (N_11789,N_11747,N_11738);
nand U11790 (N_11790,N_11574,N_11640);
nand U11791 (N_11791,N_11616,N_11667);
nor U11792 (N_11792,N_11566,N_11567);
nor U11793 (N_11793,N_11713,N_11577);
nor U11794 (N_11794,N_11548,N_11726);
and U11795 (N_11795,N_11532,N_11578);
and U11796 (N_11796,N_11740,N_11610);
nand U11797 (N_11797,N_11633,N_11520);
nand U11798 (N_11798,N_11691,N_11543);
xor U11799 (N_11799,N_11576,N_11670);
nand U11800 (N_11800,N_11564,N_11729);
and U11801 (N_11801,N_11519,N_11699);
or U11802 (N_11802,N_11725,N_11526);
xnor U11803 (N_11803,N_11582,N_11609);
nor U11804 (N_11804,N_11506,N_11716);
nor U11805 (N_11805,N_11621,N_11605);
or U11806 (N_11806,N_11693,N_11712);
nand U11807 (N_11807,N_11614,N_11736);
xor U11808 (N_11808,N_11711,N_11655);
xor U11809 (N_11809,N_11501,N_11690);
nor U11810 (N_11810,N_11683,N_11706);
nand U11811 (N_11811,N_11568,N_11748);
or U11812 (N_11812,N_11629,N_11560);
nand U11813 (N_11813,N_11537,N_11642);
nand U11814 (N_11814,N_11626,N_11708);
or U11815 (N_11815,N_11652,N_11562);
and U11816 (N_11816,N_11625,N_11530);
nor U11817 (N_11817,N_11664,N_11624);
and U11818 (N_11818,N_11601,N_11592);
or U11819 (N_11819,N_11732,N_11536);
and U11820 (N_11820,N_11698,N_11692);
nand U11821 (N_11821,N_11659,N_11593);
and U11822 (N_11822,N_11514,N_11516);
or U11823 (N_11823,N_11744,N_11602);
and U11824 (N_11824,N_11533,N_11718);
nand U11825 (N_11825,N_11703,N_11719);
or U11826 (N_11826,N_11666,N_11724);
nor U11827 (N_11827,N_11702,N_11594);
or U11828 (N_11828,N_11660,N_11544);
nor U11829 (N_11829,N_11599,N_11689);
xor U11830 (N_11830,N_11620,N_11518);
xnor U11831 (N_11831,N_11701,N_11547);
nor U11832 (N_11832,N_11672,N_11588);
xor U11833 (N_11833,N_11682,N_11579);
or U11834 (N_11834,N_11590,N_11707);
nand U11835 (N_11835,N_11505,N_11597);
nand U11836 (N_11836,N_11565,N_11528);
xor U11837 (N_11837,N_11510,N_11611);
nand U11838 (N_11838,N_11671,N_11569);
nand U11839 (N_11839,N_11535,N_11612);
nor U11840 (N_11840,N_11504,N_11649);
nand U11841 (N_11841,N_11618,N_11581);
nand U11842 (N_11842,N_11606,N_11684);
or U11843 (N_11843,N_11502,N_11631);
nand U11844 (N_11844,N_11727,N_11622);
or U11845 (N_11845,N_11608,N_11720);
nor U11846 (N_11846,N_11541,N_11737);
or U11847 (N_11847,N_11522,N_11678);
nand U11848 (N_11848,N_11645,N_11696);
and U11849 (N_11849,N_11653,N_11585);
nor U11850 (N_11850,N_11673,N_11654);
and U11851 (N_11851,N_11575,N_11680);
and U11852 (N_11852,N_11603,N_11500);
and U11853 (N_11853,N_11714,N_11694);
nand U11854 (N_11854,N_11743,N_11742);
nor U11855 (N_11855,N_11735,N_11686);
or U11856 (N_11856,N_11542,N_11688);
or U11857 (N_11857,N_11555,N_11697);
nor U11858 (N_11858,N_11647,N_11632);
nand U11859 (N_11859,N_11507,N_11628);
nor U11860 (N_11860,N_11728,N_11521);
nand U11861 (N_11861,N_11573,N_11527);
xnor U11862 (N_11862,N_11650,N_11529);
nor U11863 (N_11863,N_11613,N_11570);
nand U11864 (N_11864,N_11583,N_11559);
and U11865 (N_11865,N_11681,N_11557);
or U11866 (N_11866,N_11679,N_11700);
nor U11867 (N_11867,N_11668,N_11746);
nor U11868 (N_11868,N_11525,N_11571);
and U11869 (N_11869,N_11669,N_11595);
or U11870 (N_11870,N_11584,N_11549);
and U11871 (N_11871,N_11551,N_11515);
nand U11872 (N_11872,N_11734,N_11508);
nor U11873 (N_11873,N_11665,N_11553);
or U11874 (N_11874,N_11639,N_11540);
nand U11875 (N_11875,N_11629,N_11740);
nand U11876 (N_11876,N_11652,N_11599);
or U11877 (N_11877,N_11644,N_11581);
and U11878 (N_11878,N_11565,N_11550);
xor U11879 (N_11879,N_11620,N_11567);
nand U11880 (N_11880,N_11554,N_11606);
and U11881 (N_11881,N_11562,N_11511);
xor U11882 (N_11882,N_11559,N_11644);
or U11883 (N_11883,N_11749,N_11503);
or U11884 (N_11884,N_11514,N_11628);
or U11885 (N_11885,N_11638,N_11596);
and U11886 (N_11886,N_11616,N_11517);
nand U11887 (N_11887,N_11526,N_11631);
or U11888 (N_11888,N_11650,N_11640);
or U11889 (N_11889,N_11702,N_11649);
and U11890 (N_11890,N_11667,N_11562);
nand U11891 (N_11891,N_11540,N_11709);
and U11892 (N_11892,N_11621,N_11666);
nand U11893 (N_11893,N_11720,N_11655);
nor U11894 (N_11894,N_11644,N_11518);
nand U11895 (N_11895,N_11702,N_11664);
or U11896 (N_11896,N_11658,N_11516);
and U11897 (N_11897,N_11643,N_11708);
nor U11898 (N_11898,N_11693,N_11563);
and U11899 (N_11899,N_11508,N_11729);
or U11900 (N_11900,N_11714,N_11534);
or U11901 (N_11901,N_11522,N_11719);
nand U11902 (N_11902,N_11591,N_11618);
and U11903 (N_11903,N_11628,N_11544);
nor U11904 (N_11904,N_11735,N_11688);
and U11905 (N_11905,N_11614,N_11710);
and U11906 (N_11906,N_11715,N_11514);
or U11907 (N_11907,N_11514,N_11567);
and U11908 (N_11908,N_11622,N_11747);
and U11909 (N_11909,N_11671,N_11550);
or U11910 (N_11910,N_11636,N_11540);
nor U11911 (N_11911,N_11681,N_11619);
and U11912 (N_11912,N_11511,N_11745);
nand U11913 (N_11913,N_11705,N_11626);
nand U11914 (N_11914,N_11668,N_11678);
nand U11915 (N_11915,N_11683,N_11556);
and U11916 (N_11916,N_11543,N_11698);
xnor U11917 (N_11917,N_11637,N_11736);
nor U11918 (N_11918,N_11733,N_11603);
nand U11919 (N_11919,N_11645,N_11692);
nor U11920 (N_11920,N_11574,N_11634);
nand U11921 (N_11921,N_11702,N_11718);
nand U11922 (N_11922,N_11658,N_11630);
nand U11923 (N_11923,N_11652,N_11530);
nor U11924 (N_11924,N_11706,N_11673);
and U11925 (N_11925,N_11681,N_11533);
nand U11926 (N_11926,N_11590,N_11738);
nor U11927 (N_11927,N_11523,N_11743);
nor U11928 (N_11928,N_11685,N_11611);
or U11929 (N_11929,N_11743,N_11635);
and U11930 (N_11930,N_11524,N_11604);
xnor U11931 (N_11931,N_11736,N_11525);
and U11932 (N_11932,N_11638,N_11601);
nand U11933 (N_11933,N_11658,N_11701);
nor U11934 (N_11934,N_11513,N_11740);
nor U11935 (N_11935,N_11629,N_11666);
or U11936 (N_11936,N_11743,N_11717);
xnor U11937 (N_11937,N_11604,N_11722);
or U11938 (N_11938,N_11607,N_11576);
nor U11939 (N_11939,N_11633,N_11652);
or U11940 (N_11940,N_11589,N_11641);
nor U11941 (N_11941,N_11730,N_11511);
or U11942 (N_11942,N_11602,N_11503);
nand U11943 (N_11943,N_11670,N_11514);
xor U11944 (N_11944,N_11548,N_11582);
and U11945 (N_11945,N_11502,N_11664);
nor U11946 (N_11946,N_11567,N_11578);
and U11947 (N_11947,N_11747,N_11581);
or U11948 (N_11948,N_11563,N_11605);
and U11949 (N_11949,N_11603,N_11638);
nor U11950 (N_11950,N_11508,N_11596);
and U11951 (N_11951,N_11618,N_11617);
or U11952 (N_11952,N_11741,N_11723);
or U11953 (N_11953,N_11533,N_11629);
nand U11954 (N_11954,N_11605,N_11713);
and U11955 (N_11955,N_11705,N_11512);
or U11956 (N_11956,N_11684,N_11711);
nand U11957 (N_11957,N_11714,N_11536);
nand U11958 (N_11958,N_11714,N_11652);
and U11959 (N_11959,N_11520,N_11731);
or U11960 (N_11960,N_11579,N_11710);
xnor U11961 (N_11961,N_11597,N_11677);
or U11962 (N_11962,N_11699,N_11560);
nand U11963 (N_11963,N_11683,N_11733);
or U11964 (N_11964,N_11692,N_11583);
xnor U11965 (N_11965,N_11568,N_11650);
nand U11966 (N_11966,N_11516,N_11602);
nand U11967 (N_11967,N_11574,N_11501);
nor U11968 (N_11968,N_11712,N_11690);
nor U11969 (N_11969,N_11639,N_11502);
or U11970 (N_11970,N_11734,N_11501);
and U11971 (N_11971,N_11545,N_11717);
nor U11972 (N_11972,N_11557,N_11549);
or U11973 (N_11973,N_11722,N_11698);
nand U11974 (N_11974,N_11747,N_11563);
nand U11975 (N_11975,N_11599,N_11510);
nand U11976 (N_11976,N_11666,N_11718);
nand U11977 (N_11977,N_11523,N_11534);
nor U11978 (N_11978,N_11634,N_11562);
nand U11979 (N_11979,N_11703,N_11745);
nand U11980 (N_11980,N_11597,N_11707);
and U11981 (N_11981,N_11666,N_11593);
nand U11982 (N_11982,N_11575,N_11648);
xor U11983 (N_11983,N_11702,N_11535);
or U11984 (N_11984,N_11521,N_11645);
or U11985 (N_11985,N_11655,N_11723);
xnor U11986 (N_11986,N_11503,N_11661);
and U11987 (N_11987,N_11682,N_11552);
nor U11988 (N_11988,N_11718,N_11538);
nand U11989 (N_11989,N_11726,N_11574);
nor U11990 (N_11990,N_11619,N_11536);
nand U11991 (N_11991,N_11683,N_11597);
nand U11992 (N_11992,N_11651,N_11551);
and U11993 (N_11993,N_11571,N_11685);
and U11994 (N_11994,N_11649,N_11610);
nor U11995 (N_11995,N_11661,N_11539);
nand U11996 (N_11996,N_11656,N_11565);
nor U11997 (N_11997,N_11637,N_11617);
and U11998 (N_11998,N_11508,N_11695);
nor U11999 (N_11999,N_11714,N_11543);
nand U12000 (N_12000,N_11884,N_11771);
and U12001 (N_12001,N_11756,N_11916);
or U12002 (N_12002,N_11997,N_11868);
xor U12003 (N_12003,N_11977,N_11948);
nand U12004 (N_12004,N_11768,N_11945);
and U12005 (N_12005,N_11811,N_11949);
nor U12006 (N_12006,N_11967,N_11984);
and U12007 (N_12007,N_11780,N_11930);
and U12008 (N_12008,N_11969,N_11975);
nand U12009 (N_12009,N_11786,N_11833);
and U12010 (N_12010,N_11989,N_11912);
nor U12011 (N_12011,N_11792,N_11750);
xor U12012 (N_12012,N_11751,N_11787);
or U12013 (N_12013,N_11800,N_11812);
and U12014 (N_12014,N_11767,N_11951);
nand U12015 (N_12015,N_11866,N_11932);
nor U12016 (N_12016,N_11842,N_11878);
or U12017 (N_12017,N_11801,N_11791);
and U12018 (N_12018,N_11760,N_11858);
or U12019 (N_12019,N_11821,N_11924);
or U12020 (N_12020,N_11936,N_11946);
or U12021 (N_12021,N_11860,N_11753);
nand U12022 (N_12022,N_11877,N_11772);
xor U12023 (N_12023,N_11976,N_11900);
and U12024 (N_12024,N_11938,N_11937);
xor U12025 (N_12025,N_11859,N_11993);
or U12026 (N_12026,N_11826,N_11835);
and U12027 (N_12027,N_11939,N_11857);
nor U12028 (N_12028,N_11973,N_11817);
xnor U12029 (N_12029,N_11910,N_11864);
and U12030 (N_12030,N_11942,N_11820);
nand U12031 (N_12031,N_11844,N_11954);
and U12032 (N_12032,N_11790,N_11809);
and U12033 (N_12033,N_11763,N_11961);
nand U12034 (N_12034,N_11779,N_11956);
or U12035 (N_12035,N_11959,N_11778);
and U12036 (N_12036,N_11869,N_11853);
nor U12037 (N_12037,N_11836,N_11974);
and U12038 (N_12038,N_11970,N_11873);
and U12039 (N_12039,N_11906,N_11996);
nand U12040 (N_12040,N_11931,N_11901);
nor U12041 (N_12041,N_11886,N_11825);
or U12042 (N_12042,N_11807,N_11773);
and U12043 (N_12043,N_11905,N_11913);
xor U12044 (N_12044,N_11843,N_11830);
nand U12045 (N_12045,N_11828,N_11834);
and U12046 (N_12046,N_11920,N_11950);
or U12047 (N_12047,N_11991,N_11761);
nor U12048 (N_12048,N_11758,N_11865);
nor U12049 (N_12049,N_11781,N_11965);
or U12050 (N_12050,N_11889,N_11867);
nand U12051 (N_12051,N_11789,N_11802);
nand U12052 (N_12052,N_11831,N_11794);
or U12053 (N_12053,N_11861,N_11907);
or U12054 (N_12054,N_11943,N_11847);
nand U12055 (N_12055,N_11770,N_11926);
nand U12056 (N_12056,N_11851,N_11927);
nand U12057 (N_12057,N_11933,N_11882);
or U12058 (N_12058,N_11755,N_11776);
or U12059 (N_12059,N_11875,N_11962);
xnor U12060 (N_12060,N_11966,N_11968);
nor U12061 (N_12061,N_11915,N_11850);
nand U12062 (N_12062,N_11971,N_11764);
or U12063 (N_12063,N_11885,N_11898);
nand U12064 (N_12064,N_11797,N_11978);
nand U12065 (N_12065,N_11862,N_11964);
nor U12066 (N_12066,N_11827,N_11793);
nand U12067 (N_12067,N_11982,N_11934);
xor U12068 (N_12068,N_11899,N_11958);
nor U12069 (N_12069,N_11904,N_11838);
nand U12070 (N_12070,N_11888,N_11928);
or U12071 (N_12071,N_11863,N_11871);
and U12072 (N_12072,N_11784,N_11788);
and U12073 (N_12073,N_11908,N_11849);
or U12074 (N_12074,N_11994,N_11941);
nand U12075 (N_12075,N_11796,N_11894);
nand U12076 (N_12076,N_11981,N_11872);
nand U12077 (N_12077,N_11909,N_11810);
nor U12078 (N_12078,N_11819,N_11983);
and U12079 (N_12079,N_11952,N_11947);
nor U12080 (N_12080,N_11798,N_11953);
nor U12081 (N_12081,N_11769,N_11917);
nor U12082 (N_12082,N_11895,N_11757);
nor U12083 (N_12083,N_11785,N_11783);
and U12084 (N_12084,N_11852,N_11766);
or U12085 (N_12085,N_11824,N_11923);
and U12086 (N_12086,N_11804,N_11919);
nor U12087 (N_12087,N_11822,N_11918);
and U12088 (N_12088,N_11874,N_11903);
and U12089 (N_12089,N_11955,N_11808);
nand U12090 (N_12090,N_11775,N_11896);
nand U12091 (N_12091,N_11841,N_11979);
nor U12092 (N_12092,N_11914,N_11985);
nor U12093 (N_12093,N_11774,N_11972);
nor U12094 (N_12094,N_11876,N_11883);
nand U12095 (N_12095,N_11799,N_11944);
nor U12096 (N_12096,N_11856,N_11890);
or U12097 (N_12097,N_11752,N_11832);
nor U12098 (N_12098,N_11987,N_11814);
nand U12099 (N_12099,N_11887,N_11777);
or U12100 (N_12100,N_11829,N_11922);
nand U12101 (N_12101,N_11870,N_11840);
nand U12102 (N_12102,N_11782,N_11960);
nand U12103 (N_12103,N_11759,N_11765);
nand U12104 (N_12104,N_11988,N_11813);
xor U12105 (N_12105,N_11839,N_11806);
or U12106 (N_12106,N_11921,N_11940);
and U12107 (N_12107,N_11880,N_11911);
and U12108 (N_12108,N_11855,N_11805);
or U12109 (N_12109,N_11881,N_11957);
xnor U12110 (N_12110,N_11999,N_11963);
and U12111 (N_12111,N_11897,N_11845);
and U12112 (N_12112,N_11995,N_11879);
and U12113 (N_12113,N_11986,N_11990);
and U12114 (N_12114,N_11935,N_11893);
and U12115 (N_12115,N_11980,N_11992);
or U12116 (N_12116,N_11818,N_11846);
nand U12117 (N_12117,N_11892,N_11891);
and U12118 (N_12118,N_11815,N_11925);
and U12119 (N_12119,N_11837,N_11803);
and U12120 (N_12120,N_11998,N_11854);
nor U12121 (N_12121,N_11929,N_11902);
nand U12122 (N_12122,N_11762,N_11754);
and U12123 (N_12123,N_11823,N_11795);
nand U12124 (N_12124,N_11848,N_11816);
nor U12125 (N_12125,N_11781,N_11774);
nand U12126 (N_12126,N_11918,N_11843);
xor U12127 (N_12127,N_11812,N_11883);
nand U12128 (N_12128,N_11911,N_11868);
nand U12129 (N_12129,N_11804,N_11952);
or U12130 (N_12130,N_11975,N_11844);
nor U12131 (N_12131,N_11954,N_11795);
and U12132 (N_12132,N_11757,N_11893);
or U12133 (N_12133,N_11928,N_11963);
and U12134 (N_12134,N_11987,N_11843);
xor U12135 (N_12135,N_11770,N_11767);
nor U12136 (N_12136,N_11862,N_11786);
nand U12137 (N_12137,N_11835,N_11900);
nand U12138 (N_12138,N_11835,N_11987);
nor U12139 (N_12139,N_11774,N_11763);
or U12140 (N_12140,N_11908,N_11918);
nand U12141 (N_12141,N_11900,N_11762);
nor U12142 (N_12142,N_11830,N_11841);
and U12143 (N_12143,N_11819,N_11875);
and U12144 (N_12144,N_11872,N_11766);
nor U12145 (N_12145,N_11871,N_11908);
and U12146 (N_12146,N_11780,N_11909);
nand U12147 (N_12147,N_11782,N_11918);
nand U12148 (N_12148,N_11962,N_11933);
nand U12149 (N_12149,N_11991,N_11786);
nand U12150 (N_12150,N_11769,N_11972);
or U12151 (N_12151,N_11789,N_11856);
nand U12152 (N_12152,N_11754,N_11857);
nor U12153 (N_12153,N_11818,N_11888);
or U12154 (N_12154,N_11814,N_11931);
nand U12155 (N_12155,N_11830,N_11804);
nand U12156 (N_12156,N_11949,N_11931);
and U12157 (N_12157,N_11794,N_11905);
and U12158 (N_12158,N_11884,N_11945);
xor U12159 (N_12159,N_11753,N_11971);
nand U12160 (N_12160,N_11841,N_11995);
nor U12161 (N_12161,N_11896,N_11892);
nand U12162 (N_12162,N_11799,N_11950);
nand U12163 (N_12163,N_11919,N_11836);
nor U12164 (N_12164,N_11759,N_11826);
xor U12165 (N_12165,N_11800,N_11903);
and U12166 (N_12166,N_11840,N_11999);
or U12167 (N_12167,N_11846,N_11750);
or U12168 (N_12168,N_11997,N_11950);
xor U12169 (N_12169,N_11840,N_11751);
and U12170 (N_12170,N_11889,N_11781);
or U12171 (N_12171,N_11858,N_11857);
or U12172 (N_12172,N_11965,N_11942);
and U12173 (N_12173,N_11880,N_11927);
xor U12174 (N_12174,N_11908,N_11772);
nor U12175 (N_12175,N_11810,N_11900);
nor U12176 (N_12176,N_11999,N_11826);
nor U12177 (N_12177,N_11763,N_11867);
and U12178 (N_12178,N_11846,N_11987);
nand U12179 (N_12179,N_11805,N_11970);
nor U12180 (N_12180,N_11882,N_11892);
xnor U12181 (N_12181,N_11954,N_11949);
nor U12182 (N_12182,N_11766,N_11974);
and U12183 (N_12183,N_11837,N_11879);
xor U12184 (N_12184,N_11803,N_11985);
nand U12185 (N_12185,N_11766,N_11826);
nor U12186 (N_12186,N_11976,N_11856);
or U12187 (N_12187,N_11769,N_11961);
and U12188 (N_12188,N_11783,N_11756);
xnor U12189 (N_12189,N_11769,N_11934);
and U12190 (N_12190,N_11796,N_11962);
nand U12191 (N_12191,N_11770,N_11857);
or U12192 (N_12192,N_11959,N_11888);
and U12193 (N_12193,N_11861,N_11853);
or U12194 (N_12194,N_11853,N_11960);
nand U12195 (N_12195,N_11775,N_11947);
nand U12196 (N_12196,N_11918,N_11933);
nand U12197 (N_12197,N_11910,N_11901);
nor U12198 (N_12198,N_11766,N_11751);
xor U12199 (N_12199,N_11893,N_11794);
xor U12200 (N_12200,N_11959,N_11919);
nor U12201 (N_12201,N_11768,N_11824);
nor U12202 (N_12202,N_11867,N_11795);
or U12203 (N_12203,N_11931,N_11921);
nand U12204 (N_12204,N_11823,N_11953);
and U12205 (N_12205,N_11967,N_11896);
nor U12206 (N_12206,N_11886,N_11828);
and U12207 (N_12207,N_11826,N_11872);
and U12208 (N_12208,N_11958,N_11876);
nor U12209 (N_12209,N_11907,N_11880);
and U12210 (N_12210,N_11796,N_11918);
nand U12211 (N_12211,N_11907,N_11771);
and U12212 (N_12212,N_11847,N_11776);
and U12213 (N_12213,N_11763,N_11846);
or U12214 (N_12214,N_11797,N_11794);
nor U12215 (N_12215,N_11953,N_11785);
or U12216 (N_12216,N_11944,N_11798);
nand U12217 (N_12217,N_11918,N_11926);
nand U12218 (N_12218,N_11921,N_11972);
nand U12219 (N_12219,N_11999,N_11778);
xnor U12220 (N_12220,N_11774,N_11890);
nand U12221 (N_12221,N_11993,N_11783);
and U12222 (N_12222,N_11834,N_11776);
nor U12223 (N_12223,N_11775,N_11872);
xor U12224 (N_12224,N_11817,N_11968);
and U12225 (N_12225,N_11859,N_11971);
and U12226 (N_12226,N_11796,N_11878);
and U12227 (N_12227,N_11798,N_11763);
or U12228 (N_12228,N_11939,N_11935);
nor U12229 (N_12229,N_11914,N_11816);
and U12230 (N_12230,N_11870,N_11930);
or U12231 (N_12231,N_11768,N_11859);
nor U12232 (N_12232,N_11941,N_11915);
nor U12233 (N_12233,N_11764,N_11849);
and U12234 (N_12234,N_11907,N_11900);
or U12235 (N_12235,N_11768,N_11909);
nand U12236 (N_12236,N_11920,N_11972);
and U12237 (N_12237,N_11976,N_11926);
nor U12238 (N_12238,N_11873,N_11770);
xnor U12239 (N_12239,N_11843,N_11792);
xnor U12240 (N_12240,N_11997,N_11858);
or U12241 (N_12241,N_11942,N_11824);
xor U12242 (N_12242,N_11857,N_11913);
nor U12243 (N_12243,N_11845,N_11949);
nor U12244 (N_12244,N_11903,N_11795);
or U12245 (N_12245,N_11868,N_11772);
nor U12246 (N_12246,N_11803,N_11943);
and U12247 (N_12247,N_11846,N_11942);
or U12248 (N_12248,N_11935,N_11950);
and U12249 (N_12249,N_11779,N_11933);
and U12250 (N_12250,N_12226,N_12087);
or U12251 (N_12251,N_12149,N_12208);
nand U12252 (N_12252,N_12134,N_12094);
and U12253 (N_12253,N_12012,N_12186);
nor U12254 (N_12254,N_12187,N_12133);
or U12255 (N_12255,N_12170,N_12054);
or U12256 (N_12256,N_12061,N_12140);
xor U12257 (N_12257,N_12021,N_12029);
or U12258 (N_12258,N_12037,N_12048);
or U12259 (N_12259,N_12102,N_12229);
nor U12260 (N_12260,N_12042,N_12193);
nor U12261 (N_12261,N_12212,N_12028);
and U12262 (N_12262,N_12230,N_12143);
nand U12263 (N_12263,N_12014,N_12181);
nor U12264 (N_12264,N_12023,N_12137);
nand U12265 (N_12265,N_12110,N_12169);
nor U12266 (N_12266,N_12041,N_12103);
and U12267 (N_12267,N_12113,N_12010);
or U12268 (N_12268,N_12058,N_12067);
and U12269 (N_12269,N_12111,N_12013);
and U12270 (N_12270,N_12056,N_12178);
nand U12271 (N_12271,N_12172,N_12232);
or U12272 (N_12272,N_12018,N_12130);
nor U12273 (N_12273,N_12147,N_12151);
xnor U12274 (N_12274,N_12096,N_12183);
nor U12275 (N_12275,N_12034,N_12148);
and U12276 (N_12276,N_12166,N_12224);
or U12277 (N_12277,N_12157,N_12233);
or U12278 (N_12278,N_12081,N_12194);
nor U12279 (N_12279,N_12083,N_12039);
xnor U12280 (N_12280,N_12091,N_12249);
and U12281 (N_12281,N_12045,N_12216);
and U12282 (N_12282,N_12240,N_12248);
nor U12283 (N_12283,N_12180,N_12150);
or U12284 (N_12284,N_12132,N_12182);
nor U12285 (N_12285,N_12162,N_12128);
nand U12286 (N_12286,N_12158,N_12079);
nand U12287 (N_12287,N_12218,N_12235);
nand U12288 (N_12288,N_12173,N_12024);
nor U12289 (N_12289,N_12084,N_12247);
or U12290 (N_12290,N_12106,N_12074);
or U12291 (N_12291,N_12122,N_12097);
and U12292 (N_12292,N_12154,N_12228);
nor U12293 (N_12293,N_12125,N_12060);
or U12294 (N_12294,N_12209,N_12201);
or U12295 (N_12295,N_12070,N_12167);
nor U12296 (N_12296,N_12105,N_12065);
or U12297 (N_12297,N_12114,N_12118);
nand U12298 (N_12298,N_12221,N_12119);
nand U12299 (N_12299,N_12030,N_12197);
nor U12300 (N_12300,N_12007,N_12190);
nand U12301 (N_12301,N_12146,N_12196);
and U12302 (N_12302,N_12124,N_12062);
nand U12303 (N_12303,N_12211,N_12077);
nor U12304 (N_12304,N_12176,N_12005);
nor U12305 (N_12305,N_12243,N_12055);
or U12306 (N_12306,N_12052,N_12003);
xnor U12307 (N_12307,N_12101,N_12078);
and U12308 (N_12308,N_12053,N_12080);
and U12309 (N_12309,N_12036,N_12239);
nor U12310 (N_12310,N_12164,N_12126);
and U12311 (N_12311,N_12185,N_12090);
nand U12312 (N_12312,N_12108,N_12051);
nor U12313 (N_12313,N_12203,N_12234);
xor U12314 (N_12314,N_12099,N_12059);
nor U12315 (N_12315,N_12104,N_12214);
nor U12316 (N_12316,N_12191,N_12050);
nand U12317 (N_12317,N_12092,N_12189);
and U12318 (N_12318,N_12107,N_12109);
or U12319 (N_12319,N_12076,N_12044);
or U12320 (N_12320,N_12188,N_12011);
and U12321 (N_12321,N_12142,N_12217);
nor U12322 (N_12322,N_12004,N_12156);
and U12323 (N_12323,N_12222,N_12066);
nand U12324 (N_12324,N_12015,N_12174);
or U12325 (N_12325,N_12038,N_12095);
nand U12326 (N_12326,N_12071,N_12144);
or U12327 (N_12327,N_12121,N_12026);
nand U12328 (N_12328,N_12075,N_12245);
or U12329 (N_12329,N_12246,N_12027);
nor U12330 (N_12330,N_12152,N_12159);
and U12331 (N_12331,N_12072,N_12000);
nor U12332 (N_12332,N_12223,N_12006);
nand U12333 (N_12333,N_12184,N_12195);
or U12334 (N_12334,N_12225,N_12117);
or U12335 (N_12335,N_12236,N_12213);
nand U12336 (N_12336,N_12177,N_12093);
nand U12337 (N_12337,N_12206,N_12215);
and U12338 (N_12338,N_12068,N_12116);
nand U12339 (N_12339,N_12033,N_12161);
xor U12340 (N_12340,N_12237,N_12231);
nor U12341 (N_12341,N_12022,N_12017);
nand U12342 (N_12342,N_12088,N_12002);
nand U12343 (N_12343,N_12069,N_12085);
nor U12344 (N_12344,N_12057,N_12242);
or U12345 (N_12345,N_12160,N_12032);
nand U12346 (N_12346,N_12238,N_12227);
or U12347 (N_12347,N_12123,N_12192);
or U12348 (N_12348,N_12171,N_12244);
nor U12349 (N_12349,N_12199,N_12219);
nand U12350 (N_12350,N_12112,N_12127);
nor U12351 (N_12351,N_12009,N_12016);
or U12352 (N_12352,N_12141,N_12086);
or U12353 (N_12353,N_12198,N_12100);
nand U12354 (N_12354,N_12210,N_12008);
or U12355 (N_12355,N_12179,N_12063);
or U12356 (N_12356,N_12200,N_12064);
and U12357 (N_12357,N_12241,N_12139);
nand U12358 (N_12358,N_12165,N_12073);
and U12359 (N_12359,N_12046,N_12020);
nand U12360 (N_12360,N_12082,N_12129);
nor U12361 (N_12361,N_12089,N_12145);
and U12362 (N_12362,N_12019,N_12120);
nand U12363 (N_12363,N_12049,N_12202);
xor U12364 (N_12364,N_12204,N_12205);
nor U12365 (N_12365,N_12115,N_12163);
nand U12366 (N_12366,N_12001,N_12035);
or U12367 (N_12367,N_12207,N_12098);
nand U12368 (N_12368,N_12025,N_12153);
nor U12369 (N_12369,N_12040,N_12043);
or U12370 (N_12370,N_12155,N_12131);
and U12371 (N_12371,N_12136,N_12135);
or U12372 (N_12372,N_12220,N_12047);
or U12373 (N_12373,N_12168,N_12138);
nor U12374 (N_12374,N_12175,N_12031);
and U12375 (N_12375,N_12184,N_12236);
and U12376 (N_12376,N_12235,N_12015);
nor U12377 (N_12377,N_12243,N_12186);
or U12378 (N_12378,N_12166,N_12156);
nand U12379 (N_12379,N_12164,N_12070);
xor U12380 (N_12380,N_12091,N_12152);
nand U12381 (N_12381,N_12021,N_12014);
nand U12382 (N_12382,N_12037,N_12222);
or U12383 (N_12383,N_12166,N_12054);
nor U12384 (N_12384,N_12011,N_12224);
nand U12385 (N_12385,N_12198,N_12152);
and U12386 (N_12386,N_12213,N_12163);
or U12387 (N_12387,N_12129,N_12164);
xor U12388 (N_12388,N_12040,N_12104);
nand U12389 (N_12389,N_12100,N_12043);
xnor U12390 (N_12390,N_12084,N_12004);
or U12391 (N_12391,N_12237,N_12000);
or U12392 (N_12392,N_12197,N_12228);
or U12393 (N_12393,N_12085,N_12070);
xor U12394 (N_12394,N_12242,N_12072);
nor U12395 (N_12395,N_12037,N_12024);
and U12396 (N_12396,N_12147,N_12246);
nor U12397 (N_12397,N_12220,N_12081);
nor U12398 (N_12398,N_12193,N_12040);
nor U12399 (N_12399,N_12007,N_12113);
or U12400 (N_12400,N_12184,N_12055);
nand U12401 (N_12401,N_12027,N_12210);
or U12402 (N_12402,N_12078,N_12164);
nand U12403 (N_12403,N_12139,N_12238);
nor U12404 (N_12404,N_12064,N_12087);
and U12405 (N_12405,N_12157,N_12190);
nor U12406 (N_12406,N_12240,N_12215);
xor U12407 (N_12407,N_12164,N_12106);
nor U12408 (N_12408,N_12151,N_12024);
nand U12409 (N_12409,N_12052,N_12226);
nand U12410 (N_12410,N_12232,N_12040);
xnor U12411 (N_12411,N_12150,N_12028);
nor U12412 (N_12412,N_12029,N_12201);
nand U12413 (N_12413,N_12049,N_12248);
nand U12414 (N_12414,N_12038,N_12119);
nor U12415 (N_12415,N_12028,N_12072);
or U12416 (N_12416,N_12011,N_12220);
and U12417 (N_12417,N_12123,N_12007);
or U12418 (N_12418,N_12005,N_12194);
nor U12419 (N_12419,N_12082,N_12145);
nand U12420 (N_12420,N_12054,N_12012);
nand U12421 (N_12421,N_12090,N_12220);
xnor U12422 (N_12422,N_12209,N_12113);
nand U12423 (N_12423,N_12119,N_12032);
nand U12424 (N_12424,N_12142,N_12013);
nor U12425 (N_12425,N_12137,N_12025);
and U12426 (N_12426,N_12153,N_12189);
nor U12427 (N_12427,N_12078,N_12162);
or U12428 (N_12428,N_12136,N_12224);
or U12429 (N_12429,N_12113,N_12085);
nand U12430 (N_12430,N_12157,N_12057);
nand U12431 (N_12431,N_12027,N_12143);
and U12432 (N_12432,N_12083,N_12187);
nor U12433 (N_12433,N_12000,N_12030);
nand U12434 (N_12434,N_12102,N_12073);
nand U12435 (N_12435,N_12056,N_12092);
or U12436 (N_12436,N_12180,N_12116);
xnor U12437 (N_12437,N_12044,N_12103);
or U12438 (N_12438,N_12067,N_12078);
nor U12439 (N_12439,N_12044,N_12167);
and U12440 (N_12440,N_12205,N_12075);
xor U12441 (N_12441,N_12232,N_12012);
and U12442 (N_12442,N_12173,N_12151);
nor U12443 (N_12443,N_12026,N_12061);
and U12444 (N_12444,N_12051,N_12094);
nand U12445 (N_12445,N_12239,N_12070);
or U12446 (N_12446,N_12188,N_12043);
nand U12447 (N_12447,N_12218,N_12201);
and U12448 (N_12448,N_12178,N_12123);
and U12449 (N_12449,N_12218,N_12049);
nor U12450 (N_12450,N_12168,N_12122);
and U12451 (N_12451,N_12066,N_12096);
or U12452 (N_12452,N_12008,N_12127);
nor U12453 (N_12453,N_12163,N_12185);
nand U12454 (N_12454,N_12114,N_12175);
xnor U12455 (N_12455,N_12199,N_12038);
xor U12456 (N_12456,N_12185,N_12006);
xor U12457 (N_12457,N_12161,N_12225);
nand U12458 (N_12458,N_12125,N_12062);
nand U12459 (N_12459,N_12223,N_12217);
or U12460 (N_12460,N_12076,N_12060);
or U12461 (N_12461,N_12224,N_12179);
or U12462 (N_12462,N_12189,N_12012);
nand U12463 (N_12463,N_12150,N_12162);
xnor U12464 (N_12464,N_12060,N_12179);
and U12465 (N_12465,N_12085,N_12104);
and U12466 (N_12466,N_12101,N_12241);
nand U12467 (N_12467,N_12154,N_12225);
or U12468 (N_12468,N_12059,N_12216);
or U12469 (N_12469,N_12146,N_12176);
nor U12470 (N_12470,N_12211,N_12054);
and U12471 (N_12471,N_12061,N_12106);
nor U12472 (N_12472,N_12008,N_12194);
nand U12473 (N_12473,N_12194,N_12099);
nand U12474 (N_12474,N_12247,N_12004);
nand U12475 (N_12475,N_12176,N_12042);
nor U12476 (N_12476,N_12242,N_12156);
nor U12477 (N_12477,N_12249,N_12226);
nor U12478 (N_12478,N_12128,N_12084);
and U12479 (N_12479,N_12105,N_12100);
xor U12480 (N_12480,N_12118,N_12212);
nand U12481 (N_12481,N_12090,N_12155);
and U12482 (N_12482,N_12037,N_12025);
xnor U12483 (N_12483,N_12008,N_12161);
and U12484 (N_12484,N_12230,N_12211);
or U12485 (N_12485,N_12227,N_12217);
or U12486 (N_12486,N_12156,N_12216);
or U12487 (N_12487,N_12116,N_12207);
nor U12488 (N_12488,N_12241,N_12039);
nor U12489 (N_12489,N_12212,N_12195);
nor U12490 (N_12490,N_12123,N_12013);
xor U12491 (N_12491,N_12200,N_12245);
and U12492 (N_12492,N_12240,N_12143);
or U12493 (N_12493,N_12238,N_12010);
xnor U12494 (N_12494,N_12101,N_12194);
xor U12495 (N_12495,N_12129,N_12099);
nand U12496 (N_12496,N_12087,N_12212);
or U12497 (N_12497,N_12052,N_12099);
nand U12498 (N_12498,N_12107,N_12158);
nor U12499 (N_12499,N_12078,N_12188);
or U12500 (N_12500,N_12397,N_12271);
nand U12501 (N_12501,N_12401,N_12451);
nor U12502 (N_12502,N_12419,N_12368);
nor U12503 (N_12503,N_12478,N_12370);
or U12504 (N_12504,N_12369,N_12492);
nand U12505 (N_12505,N_12471,N_12295);
xor U12506 (N_12506,N_12319,N_12278);
xnor U12507 (N_12507,N_12480,N_12377);
or U12508 (N_12508,N_12406,N_12498);
nand U12509 (N_12509,N_12350,N_12389);
and U12510 (N_12510,N_12321,N_12291);
and U12511 (N_12511,N_12349,N_12265);
and U12512 (N_12512,N_12495,N_12470);
nor U12513 (N_12513,N_12435,N_12279);
or U12514 (N_12514,N_12491,N_12310);
nor U12515 (N_12515,N_12384,N_12475);
and U12516 (N_12516,N_12477,N_12381);
xnor U12517 (N_12517,N_12443,N_12302);
nor U12518 (N_12518,N_12269,N_12315);
nor U12519 (N_12519,N_12432,N_12476);
nor U12520 (N_12520,N_12380,N_12410);
nand U12521 (N_12521,N_12494,N_12374);
nand U12522 (N_12522,N_12454,N_12296);
nand U12523 (N_12523,N_12450,N_12353);
and U12524 (N_12524,N_12379,N_12462);
xnor U12525 (N_12525,N_12479,N_12273);
nor U12526 (N_12526,N_12425,N_12362);
nor U12527 (N_12527,N_12441,N_12412);
nand U12528 (N_12528,N_12482,N_12489);
nor U12529 (N_12529,N_12324,N_12403);
or U12530 (N_12530,N_12264,N_12300);
or U12531 (N_12531,N_12343,N_12294);
nand U12532 (N_12532,N_12405,N_12335);
or U12533 (N_12533,N_12298,N_12260);
nand U12534 (N_12534,N_12290,N_12305);
nand U12535 (N_12535,N_12372,N_12272);
nor U12536 (N_12536,N_12408,N_12304);
nand U12537 (N_12537,N_12391,N_12430);
and U12538 (N_12538,N_12359,N_12440);
nand U12539 (N_12539,N_12329,N_12276);
and U12540 (N_12540,N_12460,N_12325);
xor U12541 (N_12541,N_12448,N_12442);
or U12542 (N_12542,N_12337,N_12268);
or U12543 (N_12543,N_12348,N_12254);
nand U12544 (N_12544,N_12438,N_12292);
and U12545 (N_12545,N_12250,N_12434);
nand U12546 (N_12546,N_12277,N_12318);
nor U12547 (N_12547,N_12474,N_12280);
nor U12548 (N_12548,N_12499,N_12385);
nor U12549 (N_12549,N_12483,N_12469);
nand U12550 (N_12550,N_12358,N_12309);
and U12551 (N_12551,N_12285,N_12449);
or U12552 (N_12552,N_12466,N_12399);
nor U12553 (N_12553,N_12259,N_12418);
nor U12554 (N_12554,N_12320,N_12312);
or U12555 (N_12555,N_12365,N_12283);
and U12556 (N_12556,N_12398,N_12452);
nor U12557 (N_12557,N_12252,N_12458);
or U12558 (N_12558,N_12331,N_12444);
xnor U12559 (N_12559,N_12496,N_12356);
and U12560 (N_12560,N_12352,N_12354);
or U12561 (N_12561,N_12407,N_12263);
or U12562 (N_12562,N_12427,N_12393);
and U12563 (N_12563,N_12313,N_12428);
xor U12564 (N_12564,N_12334,N_12357);
and U12565 (N_12565,N_12484,N_12333);
nor U12566 (N_12566,N_12308,N_12409);
nor U12567 (N_12567,N_12416,N_12388);
or U12568 (N_12568,N_12346,N_12338);
or U12569 (N_12569,N_12340,N_12275);
xnor U12570 (N_12570,N_12465,N_12424);
or U12571 (N_12571,N_12431,N_12378);
nand U12572 (N_12572,N_12323,N_12421);
or U12573 (N_12573,N_12404,N_12303);
or U12574 (N_12574,N_12293,N_12307);
xor U12575 (N_12575,N_12341,N_12464);
nor U12576 (N_12576,N_12355,N_12387);
nor U12577 (N_12577,N_12426,N_12473);
and U12578 (N_12578,N_12488,N_12327);
and U12579 (N_12579,N_12455,N_12375);
xor U12580 (N_12580,N_12422,N_12395);
or U12581 (N_12581,N_12345,N_12363);
nor U12582 (N_12582,N_12456,N_12306);
nand U12583 (N_12583,N_12386,N_12415);
or U12584 (N_12584,N_12314,N_12461);
or U12585 (N_12585,N_12344,N_12330);
and U12586 (N_12586,N_12366,N_12383);
or U12587 (N_12587,N_12487,N_12485);
or U12588 (N_12588,N_12282,N_12286);
and U12589 (N_12589,N_12394,N_12360);
nand U12590 (N_12590,N_12367,N_12402);
nand U12591 (N_12591,N_12347,N_12453);
and U12592 (N_12592,N_12270,N_12437);
xor U12593 (N_12593,N_12262,N_12467);
or U12594 (N_12594,N_12253,N_12447);
or U12595 (N_12595,N_12301,N_12486);
or U12596 (N_12596,N_12289,N_12261);
nor U12597 (N_12597,N_12342,N_12255);
nand U12598 (N_12598,N_12463,N_12468);
and U12599 (N_12599,N_12413,N_12351);
xnor U12600 (N_12600,N_12392,N_12256);
or U12601 (N_12601,N_12439,N_12481);
nand U12602 (N_12602,N_12288,N_12361);
or U12603 (N_12603,N_12257,N_12400);
nor U12604 (N_12604,N_12336,N_12251);
nand U12605 (N_12605,N_12445,N_12339);
nor U12606 (N_12606,N_12472,N_12316);
xor U12607 (N_12607,N_12322,N_12382);
or U12608 (N_12608,N_12417,N_12390);
and U12609 (N_12609,N_12274,N_12436);
or U12610 (N_12610,N_12311,N_12411);
xnor U12611 (N_12611,N_12299,N_12429);
or U12612 (N_12612,N_12376,N_12446);
or U12613 (N_12613,N_12457,N_12493);
xor U12614 (N_12614,N_12414,N_12332);
nor U12615 (N_12615,N_12297,N_12287);
and U12616 (N_12616,N_12364,N_12459);
nand U12617 (N_12617,N_12490,N_12266);
or U12618 (N_12618,N_12420,N_12267);
nor U12619 (N_12619,N_12326,N_12396);
xor U12620 (N_12620,N_12258,N_12373);
nand U12621 (N_12621,N_12328,N_12497);
or U12622 (N_12622,N_12433,N_12284);
nor U12623 (N_12623,N_12371,N_12281);
or U12624 (N_12624,N_12317,N_12423);
nor U12625 (N_12625,N_12372,N_12466);
xnor U12626 (N_12626,N_12333,N_12325);
nand U12627 (N_12627,N_12405,N_12265);
nor U12628 (N_12628,N_12491,N_12489);
or U12629 (N_12629,N_12438,N_12268);
nand U12630 (N_12630,N_12373,N_12378);
or U12631 (N_12631,N_12255,N_12467);
and U12632 (N_12632,N_12430,N_12334);
nor U12633 (N_12633,N_12379,N_12442);
nand U12634 (N_12634,N_12399,N_12378);
and U12635 (N_12635,N_12493,N_12388);
and U12636 (N_12636,N_12411,N_12255);
and U12637 (N_12637,N_12309,N_12446);
nor U12638 (N_12638,N_12492,N_12253);
nor U12639 (N_12639,N_12392,N_12305);
nand U12640 (N_12640,N_12390,N_12275);
and U12641 (N_12641,N_12317,N_12447);
xnor U12642 (N_12642,N_12404,N_12417);
and U12643 (N_12643,N_12351,N_12288);
nand U12644 (N_12644,N_12444,N_12440);
nor U12645 (N_12645,N_12254,N_12293);
and U12646 (N_12646,N_12268,N_12260);
xnor U12647 (N_12647,N_12428,N_12329);
xor U12648 (N_12648,N_12398,N_12348);
or U12649 (N_12649,N_12377,N_12407);
or U12650 (N_12650,N_12318,N_12479);
nand U12651 (N_12651,N_12485,N_12423);
and U12652 (N_12652,N_12323,N_12274);
and U12653 (N_12653,N_12389,N_12306);
or U12654 (N_12654,N_12367,N_12263);
or U12655 (N_12655,N_12384,N_12333);
nor U12656 (N_12656,N_12491,N_12321);
nand U12657 (N_12657,N_12495,N_12478);
xor U12658 (N_12658,N_12403,N_12259);
xor U12659 (N_12659,N_12417,N_12487);
nand U12660 (N_12660,N_12400,N_12441);
or U12661 (N_12661,N_12498,N_12395);
nand U12662 (N_12662,N_12322,N_12324);
nand U12663 (N_12663,N_12365,N_12378);
nand U12664 (N_12664,N_12264,N_12413);
nand U12665 (N_12665,N_12438,N_12270);
or U12666 (N_12666,N_12337,N_12438);
nor U12667 (N_12667,N_12258,N_12321);
nand U12668 (N_12668,N_12424,N_12338);
and U12669 (N_12669,N_12383,N_12388);
and U12670 (N_12670,N_12465,N_12484);
nor U12671 (N_12671,N_12482,N_12344);
and U12672 (N_12672,N_12455,N_12370);
and U12673 (N_12673,N_12414,N_12469);
nor U12674 (N_12674,N_12388,N_12483);
and U12675 (N_12675,N_12417,N_12313);
or U12676 (N_12676,N_12439,N_12264);
nand U12677 (N_12677,N_12439,N_12318);
and U12678 (N_12678,N_12357,N_12305);
or U12679 (N_12679,N_12266,N_12484);
nor U12680 (N_12680,N_12371,N_12324);
or U12681 (N_12681,N_12431,N_12410);
nand U12682 (N_12682,N_12364,N_12341);
nor U12683 (N_12683,N_12432,N_12300);
or U12684 (N_12684,N_12288,N_12437);
or U12685 (N_12685,N_12463,N_12420);
and U12686 (N_12686,N_12258,N_12485);
and U12687 (N_12687,N_12285,N_12484);
or U12688 (N_12688,N_12439,N_12443);
or U12689 (N_12689,N_12381,N_12405);
nand U12690 (N_12690,N_12330,N_12476);
nand U12691 (N_12691,N_12400,N_12446);
or U12692 (N_12692,N_12384,N_12395);
nand U12693 (N_12693,N_12407,N_12286);
and U12694 (N_12694,N_12424,N_12440);
nor U12695 (N_12695,N_12387,N_12268);
nor U12696 (N_12696,N_12271,N_12333);
and U12697 (N_12697,N_12334,N_12394);
nand U12698 (N_12698,N_12438,N_12267);
and U12699 (N_12699,N_12411,N_12327);
nor U12700 (N_12700,N_12353,N_12418);
xnor U12701 (N_12701,N_12251,N_12328);
and U12702 (N_12702,N_12269,N_12360);
nor U12703 (N_12703,N_12411,N_12368);
nand U12704 (N_12704,N_12365,N_12272);
nand U12705 (N_12705,N_12381,N_12280);
xnor U12706 (N_12706,N_12477,N_12446);
or U12707 (N_12707,N_12413,N_12476);
xor U12708 (N_12708,N_12375,N_12402);
nand U12709 (N_12709,N_12278,N_12492);
nand U12710 (N_12710,N_12448,N_12435);
or U12711 (N_12711,N_12336,N_12408);
or U12712 (N_12712,N_12431,N_12327);
and U12713 (N_12713,N_12453,N_12394);
nand U12714 (N_12714,N_12475,N_12297);
and U12715 (N_12715,N_12376,N_12346);
xnor U12716 (N_12716,N_12284,N_12473);
and U12717 (N_12717,N_12389,N_12291);
nor U12718 (N_12718,N_12471,N_12273);
nand U12719 (N_12719,N_12499,N_12432);
nor U12720 (N_12720,N_12364,N_12296);
or U12721 (N_12721,N_12374,N_12499);
or U12722 (N_12722,N_12431,N_12445);
and U12723 (N_12723,N_12284,N_12271);
or U12724 (N_12724,N_12314,N_12469);
nand U12725 (N_12725,N_12475,N_12274);
or U12726 (N_12726,N_12350,N_12497);
nor U12727 (N_12727,N_12402,N_12252);
or U12728 (N_12728,N_12364,N_12424);
and U12729 (N_12729,N_12325,N_12269);
or U12730 (N_12730,N_12365,N_12296);
nand U12731 (N_12731,N_12278,N_12461);
and U12732 (N_12732,N_12412,N_12310);
or U12733 (N_12733,N_12470,N_12371);
nor U12734 (N_12734,N_12362,N_12409);
and U12735 (N_12735,N_12392,N_12261);
nand U12736 (N_12736,N_12453,N_12419);
or U12737 (N_12737,N_12365,N_12315);
nand U12738 (N_12738,N_12351,N_12273);
nor U12739 (N_12739,N_12255,N_12397);
nand U12740 (N_12740,N_12485,N_12425);
nor U12741 (N_12741,N_12494,N_12413);
nor U12742 (N_12742,N_12358,N_12442);
nor U12743 (N_12743,N_12492,N_12365);
or U12744 (N_12744,N_12274,N_12383);
xnor U12745 (N_12745,N_12467,N_12474);
xor U12746 (N_12746,N_12424,N_12370);
or U12747 (N_12747,N_12276,N_12368);
or U12748 (N_12748,N_12493,N_12272);
xnor U12749 (N_12749,N_12388,N_12264);
nand U12750 (N_12750,N_12702,N_12712);
or U12751 (N_12751,N_12603,N_12620);
xor U12752 (N_12752,N_12565,N_12654);
nor U12753 (N_12753,N_12531,N_12608);
and U12754 (N_12754,N_12672,N_12635);
nor U12755 (N_12755,N_12539,N_12749);
nor U12756 (N_12756,N_12516,N_12515);
or U12757 (N_12757,N_12541,N_12545);
xnor U12758 (N_12758,N_12696,N_12551);
nor U12759 (N_12759,N_12505,N_12562);
nand U12760 (N_12760,N_12630,N_12560);
and U12761 (N_12761,N_12552,N_12631);
nor U12762 (N_12762,N_12665,N_12546);
or U12763 (N_12763,N_12746,N_12523);
and U12764 (N_12764,N_12729,N_12659);
nor U12765 (N_12765,N_12563,N_12590);
or U12766 (N_12766,N_12673,N_12599);
and U12767 (N_12767,N_12597,N_12613);
nor U12768 (N_12768,N_12667,N_12503);
and U12769 (N_12769,N_12549,N_12610);
nand U12770 (N_12770,N_12506,N_12695);
and U12771 (N_12771,N_12533,N_12732);
or U12772 (N_12772,N_12596,N_12534);
nor U12773 (N_12773,N_12527,N_12553);
or U12774 (N_12774,N_12726,N_12711);
or U12775 (N_12775,N_12583,N_12688);
and U12776 (N_12776,N_12598,N_12669);
nand U12777 (N_12777,N_12522,N_12571);
nor U12778 (N_12778,N_12594,N_12718);
and U12779 (N_12779,N_12528,N_12614);
or U12780 (N_12780,N_12623,N_12679);
and U12781 (N_12781,N_12537,N_12676);
nand U12782 (N_12782,N_12683,N_12576);
nor U12783 (N_12783,N_12525,N_12550);
and U12784 (N_12784,N_12710,N_12668);
nand U12785 (N_12785,N_12543,N_12713);
nor U12786 (N_12786,N_12578,N_12649);
nand U12787 (N_12787,N_12540,N_12733);
or U12788 (N_12788,N_12555,N_12740);
and U12789 (N_12789,N_12684,N_12514);
or U12790 (N_12790,N_12737,N_12618);
nand U12791 (N_12791,N_12606,N_12512);
xor U12792 (N_12792,N_12530,N_12617);
and U12793 (N_12793,N_12619,N_12724);
xnor U12794 (N_12794,N_12697,N_12723);
or U12795 (N_12795,N_12587,N_12642);
or U12796 (N_12796,N_12532,N_12508);
and U12797 (N_12797,N_12526,N_12575);
nand U12798 (N_12798,N_12709,N_12693);
and U12799 (N_12799,N_12557,N_12666);
nor U12800 (N_12800,N_12636,N_12502);
nor U12801 (N_12801,N_12558,N_12577);
nand U12802 (N_12802,N_12687,N_12564);
xnor U12803 (N_12803,N_12645,N_12580);
xor U12804 (N_12804,N_12612,N_12632);
nor U12805 (N_12805,N_12520,N_12664);
nand U12806 (N_12806,N_12556,N_12727);
or U12807 (N_12807,N_12529,N_12691);
nand U12808 (N_12808,N_12653,N_12699);
nor U12809 (N_12809,N_12521,N_12700);
and U12810 (N_12810,N_12627,N_12601);
nor U12811 (N_12811,N_12567,N_12588);
and U12812 (N_12812,N_12542,N_12638);
nor U12813 (N_12813,N_12743,N_12714);
nor U12814 (N_12814,N_12655,N_12643);
xnor U12815 (N_12815,N_12509,N_12573);
nand U12816 (N_12816,N_12500,N_12742);
xnor U12817 (N_12817,N_12731,N_12650);
or U12818 (N_12818,N_12559,N_12744);
nor U12819 (N_12819,N_12621,N_12730);
nand U12820 (N_12820,N_12615,N_12535);
or U12821 (N_12821,N_12652,N_12547);
nor U12822 (N_12822,N_12611,N_12517);
or U12823 (N_12823,N_12504,N_12678);
and U12824 (N_12824,N_12640,N_12704);
or U12825 (N_12825,N_12706,N_12569);
or U12826 (N_12826,N_12663,N_12717);
nor U12827 (N_12827,N_12689,N_12698);
nor U12828 (N_12828,N_12637,N_12670);
or U12829 (N_12829,N_12589,N_12658);
or U12830 (N_12830,N_12662,N_12507);
nand U12831 (N_12831,N_12736,N_12681);
and U12832 (N_12832,N_12707,N_12511);
and U12833 (N_12833,N_12604,N_12656);
nand U12834 (N_12834,N_12701,N_12519);
nor U12835 (N_12835,N_12671,N_12641);
and U12836 (N_12836,N_12660,N_12719);
nor U12837 (N_12837,N_12579,N_12566);
nor U12838 (N_12838,N_12720,N_12685);
and U12839 (N_12839,N_12651,N_12748);
nor U12840 (N_12840,N_12657,N_12626);
xor U12841 (N_12841,N_12739,N_12647);
and U12842 (N_12842,N_12682,N_12694);
nor U12843 (N_12843,N_12524,N_12734);
nor U12844 (N_12844,N_12536,N_12554);
nand U12845 (N_12845,N_12633,N_12741);
and U12846 (N_12846,N_12570,N_12747);
xor U12847 (N_12847,N_12593,N_12501);
nand U12848 (N_12848,N_12634,N_12722);
nor U12849 (N_12849,N_12605,N_12624);
nor U12850 (N_12850,N_12690,N_12703);
nor U12851 (N_12851,N_12677,N_12648);
or U12852 (N_12852,N_12622,N_12538);
nand U12853 (N_12853,N_12629,N_12628);
or U12854 (N_12854,N_12745,N_12600);
xnor U12855 (N_12855,N_12721,N_12510);
nand U12856 (N_12856,N_12602,N_12574);
or U12857 (N_12857,N_12513,N_12616);
nor U12858 (N_12858,N_12708,N_12609);
or U12859 (N_12859,N_12625,N_12728);
nand U12860 (N_12860,N_12738,N_12572);
nand U12861 (N_12861,N_12561,N_12715);
and U12862 (N_12862,N_12585,N_12548);
or U12863 (N_12863,N_12675,N_12646);
xnor U12864 (N_12864,N_12725,N_12584);
xor U12865 (N_12865,N_12661,N_12568);
and U12866 (N_12866,N_12716,N_12582);
or U12867 (N_12867,N_12581,N_12518);
nand U12868 (N_12868,N_12591,N_12674);
and U12869 (N_12869,N_12644,N_12680);
and U12870 (N_12870,N_12692,N_12735);
or U12871 (N_12871,N_12705,N_12607);
nand U12872 (N_12872,N_12595,N_12586);
or U12873 (N_12873,N_12544,N_12592);
nand U12874 (N_12874,N_12686,N_12639);
xor U12875 (N_12875,N_12648,N_12697);
nand U12876 (N_12876,N_12684,N_12596);
and U12877 (N_12877,N_12736,N_12711);
xor U12878 (N_12878,N_12564,N_12523);
or U12879 (N_12879,N_12692,N_12526);
nor U12880 (N_12880,N_12610,N_12623);
nand U12881 (N_12881,N_12548,N_12703);
nand U12882 (N_12882,N_12746,N_12510);
or U12883 (N_12883,N_12728,N_12569);
nand U12884 (N_12884,N_12528,N_12650);
and U12885 (N_12885,N_12656,N_12595);
nand U12886 (N_12886,N_12640,N_12699);
or U12887 (N_12887,N_12594,N_12539);
nor U12888 (N_12888,N_12718,N_12727);
nand U12889 (N_12889,N_12736,N_12695);
and U12890 (N_12890,N_12637,N_12623);
or U12891 (N_12891,N_12601,N_12708);
nand U12892 (N_12892,N_12715,N_12725);
or U12893 (N_12893,N_12692,N_12748);
or U12894 (N_12894,N_12597,N_12737);
and U12895 (N_12895,N_12741,N_12716);
and U12896 (N_12896,N_12585,N_12747);
and U12897 (N_12897,N_12543,N_12573);
or U12898 (N_12898,N_12516,N_12507);
or U12899 (N_12899,N_12554,N_12706);
nand U12900 (N_12900,N_12507,N_12619);
and U12901 (N_12901,N_12543,N_12535);
nor U12902 (N_12902,N_12590,N_12730);
or U12903 (N_12903,N_12515,N_12535);
or U12904 (N_12904,N_12743,N_12703);
and U12905 (N_12905,N_12585,N_12666);
and U12906 (N_12906,N_12668,N_12650);
nand U12907 (N_12907,N_12556,N_12566);
or U12908 (N_12908,N_12684,N_12573);
or U12909 (N_12909,N_12542,N_12696);
and U12910 (N_12910,N_12635,N_12603);
nor U12911 (N_12911,N_12670,N_12672);
xnor U12912 (N_12912,N_12626,N_12505);
nand U12913 (N_12913,N_12674,N_12613);
nand U12914 (N_12914,N_12556,N_12568);
or U12915 (N_12915,N_12520,N_12648);
nand U12916 (N_12916,N_12645,N_12551);
nand U12917 (N_12917,N_12513,N_12528);
and U12918 (N_12918,N_12655,N_12590);
nor U12919 (N_12919,N_12698,N_12547);
nor U12920 (N_12920,N_12519,N_12523);
xor U12921 (N_12921,N_12634,N_12545);
nor U12922 (N_12922,N_12717,N_12733);
nand U12923 (N_12923,N_12694,N_12555);
and U12924 (N_12924,N_12613,N_12527);
nand U12925 (N_12925,N_12627,N_12619);
nor U12926 (N_12926,N_12700,N_12628);
nand U12927 (N_12927,N_12579,N_12530);
or U12928 (N_12928,N_12534,N_12727);
or U12929 (N_12929,N_12583,N_12669);
and U12930 (N_12930,N_12697,N_12556);
nand U12931 (N_12931,N_12662,N_12567);
or U12932 (N_12932,N_12574,N_12616);
or U12933 (N_12933,N_12530,N_12534);
nand U12934 (N_12934,N_12629,N_12603);
nand U12935 (N_12935,N_12573,N_12695);
nand U12936 (N_12936,N_12625,N_12553);
and U12937 (N_12937,N_12613,N_12549);
and U12938 (N_12938,N_12707,N_12690);
nor U12939 (N_12939,N_12662,N_12623);
and U12940 (N_12940,N_12705,N_12541);
and U12941 (N_12941,N_12703,N_12567);
nor U12942 (N_12942,N_12702,N_12532);
and U12943 (N_12943,N_12500,N_12637);
and U12944 (N_12944,N_12653,N_12686);
nand U12945 (N_12945,N_12646,N_12729);
or U12946 (N_12946,N_12749,N_12643);
and U12947 (N_12947,N_12502,N_12730);
and U12948 (N_12948,N_12617,N_12611);
or U12949 (N_12949,N_12626,N_12526);
nor U12950 (N_12950,N_12645,N_12656);
nand U12951 (N_12951,N_12683,N_12550);
and U12952 (N_12952,N_12686,N_12665);
or U12953 (N_12953,N_12591,N_12647);
nor U12954 (N_12954,N_12724,N_12670);
nor U12955 (N_12955,N_12699,N_12726);
or U12956 (N_12956,N_12695,N_12521);
nor U12957 (N_12957,N_12654,N_12641);
or U12958 (N_12958,N_12638,N_12709);
and U12959 (N_12959,N_12633,N_12703);
and U12960 (N_12960,N_12522,N_12593);
and U12961 (N_12961,N_12713,N_12709);
and U12962 (N_12962,N_12743,N_12646);
nor U12963 (N_12963,N_12718,N_12630);
or U12964 (N_12964,N_12638,N_12677);
nor U12965 (N_12965,N_12520,N_12654);
nand U12966 (N_12966,N_12580,N_12713);
nor U12967 (N_12967,N_12702,N_12689);
and U12968 (N_12968,N_12633,N_12748);
and U12969 (N_12969,N_12645,N_12567);
nor U12970 (N_12970,N_12727,N_12504);
xor U12971 (N_12971,N_12741,N_12603);
or U12972 (N_12972,N_12573,N_12620);
nand U12973 (N_12973,N_12583,N_12515);
nor U12974 (N_12974,N_12710,N_12566);
and U12975 (N_12975,N_12534,N_12712);
nand U12976 (N_12976,N_12580,N_12641);
nand U12977 (N_12977,N_12691,N_12732);
and U12978 (N_12978,N_12610,N_12733);
or U12979 (N_12979,N_12567,N_12535);
or U12980 (N_12980,N_12616,N_12520);
nand U12981 (N_12981,N_12679,N_12597);
nor U12982 (N_12982,N_12658,N_12599);
nand U12983 (N_12983,N_12620,N_12680);
nand U12984 (N_12984,N_12698,N_12637);
nand U12985 (N_12985,N_12726,N_12706);
or U12986 (N_12986,N_12542,N_12518);
xnor U12987 (N_12987,N_12522,N_12616);
nor U12988 (N_12988,N_12676,N_12645);
and U12989 (N_12989,N_12714,N_12689);
nor U12990 (N_12990,N_12746,N_12708);
or U12991 (N_12991,N_12505,N_12580);
nor U12992 (N_12992,N_12530,N_12737);
or U12993 (N_12993,N_12663,N_12649);
nor U12994 (N_12994,N_12653,N_12664);
or U12995 (N_12995,N_12634,N_12532);
xor U12996 (N_12996,N_12519,N_12527);
or U12997 (N_12997,N_12740,N_12566);
nand U12998 (N_12998,N_12725,N_12701);
or U12999 (N_12999,N_12602,N_12511);
nor U13000 (N_13000,N_12783,N_12851);
or U13001 (N_13001,N_12994,N_12806);
nor U13002 (N_13002,N_12912,N_12856);
and U13003 (N_13003,N_12770,N_12928);
and U13004 (N_13004,N_12914,N_12801);
nor U13005 (N_13005,N_12891,N_12820);
and U13006 (N_13006,N_12924,N_12976);
or U13007 (N_13007,N_12958,N_12870);
nand U13008 (N_13008,N_12903,N_12967);
and U13009 (N_13009,N_12835,N_12800);
xor U13010 (N_13010,N_12962,N_12769);
or U13011 (N_13011,N_12969,N_12937);
nor U13012 (N_13012,N_12838,N_12947);
nor U13013 (N_13013,N_12951,N_12916);
or U13014 (N_13014,N_12885,N_12817);
nand U13015 (N_13015,N_12865,N_12883);
nor U13016 (N_13016,N_12946,N_12918);
or U13017 (N_13017,N_12857,N_12753);
and U13018 (N_13018,N_12797,N_12847);
or U13019 (N_13019,N_12935,N_12989);
nand U13020 (N_13020,N_12982,N_12970);
or U13021 (N_13021,N_12786,N_12861);
and U13022 (N_13022,N_12874,N_12775);
nor U13023 (N_13023,N_12878,N_12884);
nand U13024 (N_13024,N_12944,N_12984);
nand U13025 (N_13025,N_12790,N_12936);
nor U13026 (N_13026,N_12755,N_12866);
or U13027 (N_13027,N_12767,N_12909);
and U13028 (N_13028,N_12754,N_12873);
nor U13029 (N_13029,N_12888,N_12986);
nor U13030 (N_13030,N_12802,N_12807);
or U13031 (N_13031,N_12834,N_12899);
xnor U13032 (N_13032,N_12990,N_12798);
or U13033 (N_13033,N_12752,N_12824);
or U13034 (N_13034,N_12751,N_12893);
or U13035 (N_13035,N_12814,N_12862);
nor U13036 (N_13036,N_12995,N_12975);
and U13037 (N_13037,N_12945,N_12942);
or U13038 (N_13038,N_12904,N_12964);
xor U13039 (N_13039,N_12882,N_12842);
and U13040 (N_13040,N_12950,N_12913);
xor U13041 (N_13041,N_12941,N_12987);
and U13042 (N_13042,N_12860,N_12889);
nor U13043 (N_13043,N_12940,N_12934);
and U13044 (N_13044,N_12818,N_12845);
nor U13045 (N_13045,N_12892,N_12826);
nand U13046 (N_13046,N_12762,N_12796);
nand U13047 (N_13047,N_12778,N_12821);
and U13048 (N_13048,N_12991,N_12863);
nand U13049 (N_13049,N_12988,N_12760);
and U13050 (N_13050,N_12898,N_12864);
nand U13051 (N_13051,N_12768,N_12774);
or U13052 (N_13052,N_12811,N_12779);
nand U13053 (N_13053,N_12812,N_12894);
nand U13054 (N_13054,N_12854,N_12922);
or U13055 (N_13055,N_12792,N_12771);
nor U13056 (N_13056,N_12780,N_12999);
and U13057 (N_13057,N_12756,N_12897);
or U13058 (N_13058,N_12939,N_12895);
xnor U13059 (N_13059,N_12773,N_12795);
or U13060 (N_13060,N_12846,N_12997);
nand U13061 (N_13061,N_12829,N_12876);
or U13062 (N_13062,N_12996,N_12849);
or U13063 (N_13063,N_12993,N_12759);
nand U13064 (N_13064,N_12973,N_12850);
and U13065 (N_13065,N_12900,N_12948);
nor U13066 (N_13066,N_12877,N_12839);
and U13067 (N_13067,N_12929,N_12926);
nor U13068 (N_13068,N_12750,N_12852);
nand U13069 (N_13069,N_12831,N_12979);
nor U13070 (N_13070,N_12772,N_12933);
and U13071 (N_13071,N_12886,N_12963);
nand U13072 (N_13072,N_12954,N_12917);
nand U13073 (N_13073,N_12765,N_12853);
or U13074 (N_13074,N_12804,N_12789);
or U13075 (N_13075,N_12887,N_12784);
nor U13076 (N_13076,N_12881,N_12932);
or U13077 (N_13077,N_12761,N_12957);
nand U13078 (N_13078,N_12825,N_12906);
nor U13079 (N_13079,N_12896,N_12844);
nand U13080 (N_13080,N_12799,N_12978);
or U13081 (N_13081,N_12920,N_12827);
nand U13082 (N_13082,N_12943,N_12902);
or U13083 (N_13083,N_12901,N_12828);
or U13084 (N_13084,N_12983,N_12974);
xnor U13085 (N_13085,N_12910,N_12869);
and U13086 (N_13086,N_12848,N_12757);
and U13087 (N_13087,N_12766,N_12810);
nor U13088 (N_13088,N_12822,N_12785);
or U13089 (N_13089,N_12980,N_12794);
nor U13090 (N_13090,N_12938,N_12890);
nor U13091 (N_13091,N_12919,N_12777);
nand U13092 (N_13092,N_12808,N_12809);
and U13093 (N_13093,N_12966,N_12868);
nor U13094 (N_13094,N_12992,N_12764);
or U13095 (N_13095,N_12927,N_12781);
nand U13096 (N_13096,N_12787,N_12915);
xnor U13097 (N_13097,N_12833,N_12921);
or U13098 (N_13098,N_12972,N_12953);
nor U13099 (N_13099,N_12859,N_12841);
or U13100 (N_13100,N_12837,N_12758);
and U13101 (N_13101,N_12855,N_12843);
nor U13102 (N_13102,N_12880,N_12830);
nand U13103 (N_13103,N_12952,N_12965);
nor U13104 (N_13104,N_12875,N_12840);
and U13105 (N_13105,N_12836,N_12908);
nand U13106 (N_13106,N_12949,N_12905);
and U13107 (N_13107,N_12763,N_12931);
nand U13108 (N_13108,N_12793,N_12985);
or U13109 (N_13109,N_12871,N_12791);
or U13110 (N_13110,N_12930,N_12907);
nand U13111 (N_13111,N_12776,N_12925);
nor U13112 (N_13112,N_12832,N_12872);
and U13113 (N_13113,N_12813,N_12819);
or U13114 (N_13114,N_12805,N_12960);
nor U13115 (N_13115,N_12959,N_12867);
nand U13116 (N_13116,N_12971,N_12816);
and U13117 (N_13117,N_12956,N_12911);
nand U13118 (N_13118,N_12955,N_12961);
nor U13119 (N_13119,N_12879,N_12788);
or U13120 (N_13120,N_12858,N_12782);
nand U13121 (N_13121,N_12968,N_12923);
nand U13122 (N_13122,N_12998,N_12981);
nor U13123 (N_13123,N_12815,N_12823);
nor U13124 (N_13124,N_12803,N_12977);
nand U13125 (N_13125,N_12793,N_12916);
nor U13126 (N_13126,N_12919,N_12766);
nor U13127 (N_13127,N_12840,N_12900);
nand U13128 (N_13128,N_12771,N_12855);
xor U13129 (N_13129,N_12794,N_12771);
nor U13130 (N_13130,N_12806,N_12851);
or U13131 (N_13131,N_12945,N_12838);
and U13132 (N_13132,N_12948,N_12997);
nor U13133 (N_13133,N_12858,N_12996);
nor U13134 (N_13134,N_12761,N_12861);
nor U13135 (N_13135,N_12981,N_12791);
and U13136 (N_13136,N_12835,N_12777);
nor U13137 (N_13137,N_12954,N_12770);
and U13138 (N_13138,N_12820,N_12987);
and U13139 (N_13139,N_12790,N_12978);
xnor U13140 (N_13140,N_12781,N_12864);
xnor U13141 (N_13141,N_12771,N_12804);
xor U13142 (N_13142,N_12847,N_12854);
and U13143 (N_13143,N_12936,N_12911);
or U13144 (N_13144,N_12773,N_12946);
nor U13145 (N_13145,N_12752,N_12784);
and U13146 (N_13146,N_12784,N_12941);
or U13147 (N_13147,N_12939,N_12965);
or U13148 (N_13148,N_12897,N_12871);
and U13149 (N_13149,N_12771,N_12936);
nor U13150 (N_13150,N_12949,N_12898);
nand U13151 (N_13151,N_12887,N_12836);
nand U13152 (N_13152,N_12996,N_12795);
nand U13153 (N_13153,N_12830,N_12789);
nand U13154 (N_13154,N_12937,N_12897);
or U13155 (N_13155,N_12793,N_12903);
xnor U13156 (N_13156,N_12999,N_12968);
and U13157 (N_13157,N_12833,N_12895);
and U13158 (N_13158,N_12913,N_12795);
and U13159 (N_13159,N_12758,N_12793);
and U13160 (N_13160,N_12750,N_12763);
and U13161 (N_13161,N_12841,N_12984);
nand U13162 (N_13162,N_12804,N_12919);
or U13163 (N_13163,N_12832,N_12996);
nor U13164 (N_13164,N_12878,N_12940);
nor U13165 (N_13165,N_12797,N_12801);
nor U13166 (N_13166,N_12931,N_12797);
xnor U13167 (N_13167,N_12852,N_12824);
nor U13168 (N_13168,N_12795,N_12919);
nor U13169 (N_13169,N_12897,N_12913);
nand U13170 (N_13170,N_12776,N_12790);
xor U13171 (N_13171,N_12839,N_12851);
nor U13172 (N_13172,N_12932,N_12968);
nor U13173 (N_13173,N_12945,N_12903);
nor U13174 (N_13174,N_12765,N_12824);
nor U13175 (N_13175,N_12832,N_12917);
or U13176 (N_13176,N_12752,N_12843);
or U13177 (N_13177,N_12759,N_12773);
xor U13178 (N_13178,N_12974,N_12917);
and U13179 (N_13179,N_12929,N_12863);
nor U13180 (N_13180,N_12790,N_12799);
or U13181 (N_13181,N_12804,N_12828);
and U13182 (N_13182,N_12979,N_12922);
or U13183 (N_13183,N_12821,N_12960);
nor U13184 (N_13184,N_12946,N_12835);
nor U13185 (N_13185,N_12850,N_12911);
nor U13186 (N_13186,N_12928,N_12752);
nor U13187 (N_13187,N_12835,N_12795);
nor U13188 (N_13188,N_12779,N_12957);
and U13189 (N_13189,N_12781,N_12976);
nand U13190 (N_13190,N_12804,N_12930);
nand U13191 (N_13191,N_12891,N_12768);
or U13192 (N_13192,N_12828,N_12834);
or U13193 (N_13193,N_12840,N_12775);
nor U13194 (N_13194,N_12947,N_12852);
or U13195 (N_13195,N_12861,N_12766);
nand U13196 (N_13196,N_12832,N_12767);
nor U13197 (N_13197,N_12806,N_12877);
and U13198 (N_13198,N_12771,N_12832);
xnor U13199 (N_13199,N_12764,N_12774);
nand U13200 (N_13200,N_12828,N_12816);
and U13201 (N_13201,N_12838,N_12998);
or U13202 (N_13202,N_12908,N_12778);
nand U13203 (N_13203,N_12769,N_12994);
and U13204 (N_13204,N_12938,N_12897);
and U13205 (N_13205,N_12823,N_12938);
xor U13206 (N_13206,N_12984,N_12779);
nand U13207 (N_13207,N_12958,N_12757);
xor U13208 (N_13208,N_12859,N_12852);
nand U13209 (N_13209,N_12995,N_12842);
nor U13210 (N_13210,N_12789,N_12984);
nand U13211 (N_13211,N_12874,N_12778);
nand U13212 (N_13212,N_12804,N_12941);
and U13213 (N_13213,N_12855,N_12834);
nor U13214 (N_13214,N_12834,N_12762);
nand U13215 (N_13215,N_12829,N_12982);
nor U13216 (N_13216,N_12825,N_12885);
and U13217 (N_13217,N_12774,N_12754);
xnor U13218 (N_13218,N_12907,N_12756);
and U13219 (N_13219,N_12943,N_12929);
and U13220 (N_13220,N_12859,N_12803);
and U13221 (N_13221,N_12974,N_12763);
and U13222 (N_13222,N_12978,N_12988);
or U13223 (N_13223,N_12878,N_12854);
nand U13224 (N_13224,N_12822,N_12808);
nor U13225 (N_13225,N_12941,N_12771);
nand U13226 (N_13226,N_12935,N_12797);
and U13227 (N_13227,N_12888,N_12926);
and U13228 (N_13228,N_12808,N_12862);
and U13229 (N_13229,N_12949,N_12809);
or U13230 (N_13230,N_12891,N_12812);
nand U13231 (N_13231,N_12929,N_12854);
and U13232 (N_13232,N_12771,N_12992);
nor U13233 (N_13233,N_12830,N_12915);
xor U13234 (N_13234,N_12895,N_12899);
or U13235 (N_13235,N_12909,N_12819);
and U13236 (N_13236,N_12987,N_12957);
and U13237 (N_13237,N_12868,N_12804);
nand U13238 (N_13238,N_12862,N_12763);
or U13239 (N_13239,N_12914,N_12854);
or U13240 (N_13240,N_12800,N_12810);
nor U13241 (N_13241,N_12865,N_12836);
or U13242 (N_13242,N_12840,N_12827);
nand U13243 (N_13243,N_12767,N_12838);
and U13244 (N_13244,N_12905,N_12833);
nor U13245 (N_13245,N_12965,N_12784);
nor U13246 (N_13246,N_12920,N_12919);
and U13247 (N_13247,N_12874,N_12836);
or U13248 (N_13248,N_12857,N_12916);
nand U13249 (N_13249,N_12802,N_12822);
or U13250 (N_13250,N_13065,N_13244);
xor U13251 (N_13251,N_13175,N_13114);
nor U13252 (N_13252,N_13106,N_13185);
and U13253 (N_13253,N_13205,N_13157);
and U13254 (N_13254,N_13060,N_13131);
or U13255 (N_13255,N_13159,N_13195);
and U13256 (N_13256,N_13110,N_13230);
and U13257 (N_13257,N_13162,N_13071);
or U13258 (N_13258,N_13059,N_13011);
nand U13259 (N_13259,N_13103,N_13246);
or U13260 (N_13260,N_13031,N_13228);
or U13261 (N_13261,N_13191,N_13168);
xnor U13262 (N_13262,N_13098,N_13123);
nand U13263 (N_13263,N_13221,N_13188);
nor U13264 (N_13264,N_13143,N_13164);
or U13265 (N_13265,N_13112,N_13196);
nor U13266 (N_13266,N_13202,N_13058);
nor U13267 (N_13267,N_13139,N_13227);
nand U13268 (N_13268,N_13086,N_13117);
nand U13269 (N_13269,N_13160,N_13122);
nor U13270 (N_13270,N_13240,N_13197);
and U13271 (N_13271,N_13001,N_13033);
or U13272 (N_13272,N_13237,N_13146);
or U13273 (N_13273,N_13163,N_13049);
and U13274 (N_13274,N_13004,N_13152);
and U13275 (N_13275,N_13018,N_13245);
and U13276 (N_13276,N_13064,N_13095);
nor U13277 (N_13277,N_13238,N_13116);
or U13278 (N_13278,N_13153,N_13189);
nand U13279 (N_13279,N_13040,N_13073);
or U13280 (N_13280,N_13102,N_13134);
xor U13281 (N_13281,N_13050,N_13150);
xor U13282 (N_13282,N_13120,N_13124);
nor U13283 (N_13283,N_13019,N_13027);
nand U13284 (N_13284,N_13022,N_13192);
and U13285 (N_13285,N_13078,N_13200);
and U13286 (N_13286,N_13198,N_13066);
nor U13287 (N_13287,N_13101,N_13247);
xor U13288 (N_13288,N_13068,N_13155);
and U13289 (N_13289,N_13046,N_13145);
and U13290 (N_13290,N_13051,N_13125);
or U13291 (N_13291,N_13056,N_13016);
nand U13292 (N_13292,N_13069,N_13231);
and U13293 (N_13293,N_13020,N_13063);
nand U13294 (N_13294,N_13072,N_13184);
nor U13295 (N_13295,N_13029,N_13061);
nand U13296 (N_13296,N_13190,N_13206);
nand U13297 (N_13297,N_13218,N_13142);
nor U13298 (N_13298,N_13234,N_13107);
nand U13299 (N_13299,N_13109,N_13130);
nand U13300 (N_13300,N_13235,N_13092);
xnor U13301 (N_13301,N_13126,N_13085);
xor U13302 (N_13302,N_13242,N_13104);
nor U13303 (N_13303,N_13222,N_13147);
and U13304 (N_13304,N_13167,N_13075);
and U13305 (N_13305,N_13089,N_13201);
nand U13306 (N_13306,N_13249,N_13013);
or U13307 (N_13307,N_13127,N_13052);
nor U13308 (N_13308,N_13096,N_13165);
nor U13309 (N_13309,N_13180,N_13177);
nand U13310 (N_13310,N_13079,N_13045);
or U13311 (N_13311,N_13121,N_13181);
nand U13312 (N_13312,N_13156,N_13225);
nand U13313 (N_13313,N_13178,N_13008);
or U13314 (N_13314,N_13236,N_13111);
nor U13315 (N_13315,N_13183,N_13014);
nor U13316 (N_13316,N_13074,N_13173);
and U13317 (N_13317,N_13039,N_13132);
or U13318 (N_13318,N_13009,N_13118);
nor U13319 (N_13319,N_13047,N_13161);
or U13320 (N_13320,N_13084,N_13158);
and U13321 (N_13321,N_13044,N_13091);
xor U13322 (N_13322,N_13224,N_13149);
and U13323 (N_13323,N_13024,N_13210);
or U13324 (N_13324,N_13119,N_13172);
nor U13325 (N_13325,N_13010,N_13216);
nand U13326 (N_13326,N_13076,N_13229);
and U13327 (N_13327,N_13169,N_13128);
or U13328 (N_13328,N_13211,N_13193);
or U13329 (N_13329,N_13048,N_13219);
and U13330 (N_13330,N_13232,N_13088);
nand U13331 (N_13331,N_13062,N_13166);
and U13332 (N_13332,N_13017,N_13041);
nand U13333 (N_13333,N_13209,N_13151);
xor U13334 (N_13334,N_13241,N_13093);
nor U13335 (N_13335,N_13203,N_13057);
nor U13336 (N_13336,N_13021,N_13115);
nor U13337 (N_13337,N_13182,N_13037);
and U13338 (N_13338,N_13032,N_13034);
or U13339 (N_13339,N_13215,N_13030);
nor U13340 (N_13340,N_13187,N_13179);
nand U13341 (N_13341,N_13204,N_13105);
or U13342 (N_13342,N_13070,N_13080);
nor U13343 (N_13343,N_13067,N_13137);
nor U13344 (N_13344,N_13006,N_13136);
nor U13345 (N_13345,N_13000,N_13199);
nand U13346 (N_13346,N_13170,N_13007);
and U13347 (N_13347,N_13043,N_13082);
nand U13348 (N_13348,N_13243,N_13171);
nand U13349 (N_13349,N_13217,N_13081);
or U13350 (N_13350,N_13023,N_13015);
nor U13351 (N_13351,N_13208,N_13077);
nor U13352 (N_13352,N_13002,N_13053);
nand U13353 (N_13353,N_13012,N_13113);
nand U13354 (N_13354,N_13226,N_13129);
or U13355 (N_13355,N_13055,N_13099);
and U13356 (N_13356,N_13138,N_13026);
or U13357 (N_13357,N_13028,N_13108);
or U13358 (N_13358,N_13005,N_13094);
nand U13359 (N_13359,N_13220,N_13154);
or U13360 (N_13360,N_13144,N_13042);
and U13361 (N_13361,N_13223,N_13133);
nand U13362 (N_13362,N_13207,N_13176);
and U13363 (N_13363,N_13003,N_13194);
nor U13364 (N_13364,N_13097,N_13038);
nand U13365 (N_13365,N_13174,N_13100);
nor U13366 (N_13366,N_13036,N_13148);
nand U13367 (N_13367,N_13233,N_13213);
nor U13368 (N_13368,N_13135,N_13186);
xnor U13369 (N_13369,N_13141,N_13025);
or U13370 (N_13370,N_13214,N_13212);
nor U13371 (N_13371,N_13087,N_13140);
or U13372 (N_13372,N_13248,N_13090);
nor U13373 (N_13373,N_13083,N_13239);
and U13374 (N_13374,N_13035,N_13054);
xnor U13375 (N_13375,N_13221,N_13083);
nand U13376 (N_13376,N_13027,N_13080);
xnor U13377 (N_13377,N_13116,N_13095);
or U13378 (N_13378,N_13006,N_13070);
xor U13379 (N_13379,N_13221,N_13187);
or U13380 (N_13380,N_13028,N_13115);
or U13381 (N_13381,N_13182,N_13120);
or U13382 (N_13382,N_13217,N_13115);
and U13383 (N_13383,N_13109,N_13035);
xor U13384 (N_13384,N_13056,N_13012);
and U13385 (N_13385,N_13065,N_13139);
nor U13386 (N_13386,N_13210,N_13079);
or U13387 (N_13387,N_13226,N_13132);
nor U13388 (N_13388,N_13033,N_13046);
or U13389 (N_13389,N_13114,N_13038);
and U13390 (N_13390,N_13184,N_13070);
nand U13391 (N_13391,N_13177,N_13195);
xnor U13392 (N_13392,N_13089,N_13149);
nor U13393 (N_13393,N_13104,N_13238);
or U13394 (N_13394,N_13213,N_13201);
nand U13395 (N_13395,N_13010,N_13032);
nor U13396 (N_13396,N_13163,N_13069);
nor U13397 (N_13397,N_13036,N_13243);
xnor U13398 (N_13398,N_13204,N_13197);
or U13399 (N_13399,N_13066,N_13234);
nand U13400 (N_13400,N_13133,N_13048);
and U13401 (N_13401,N_13006,N_13022);
and U13402 (N_13402,N_13108,N_13007);
or U13403 (N_13403,N_13110,N_13098);
nor U13404 (N_13404,N_13153,N_13194);
nand U13405 (N_13405,N_13041,N_13169);
and U13406 (N_13406,N_13146,N_13162);
nor U13407 (N_13407,N_13177,N_13085);
and U13408 (N_13408,N_13103,N_13121);
nor U13409 (N_13409,N_13185,N_13013);
and U13410 (N_13410,N_13185,N_13146);
or U13411 (N_13411,N_13140,N_13149);
and U13412 (N_13412,N_13218,N_13160);
or U13413 (N_13413,N_13173,N_13051);
nor U13414 (N_13414,N_13062,N_13044);
nor U13415 (N_13415,N_13202,N_13124);
nand U13416 (N_13416,N_13232,N_13136);
or U13417 (N_13417,N_13206,N_13127);
nand U13418 (N_13418,N_13117,N_13120);
and U13419 (N_13419,N_13199,N_13178);
or U13420 (N_13420,N_13105,N_13089);
and U13421 (N_13421,N_13057,N_13080);
nand U13422 (N_13422,N_13039,N_13122);
nand U13423 (N_13423,N_13093,N_13103);
nor U13424 (N_13424,N_13096,N_13234);
nor U13425 (N_13425,N_13127,N_13227);
nor U13426 (N_13426,N_13147,N_13001);
nand U13427 (N_13427,N_13075,N_13202);
xor U13428 (N_13428,N_13194,N_13057);
nand U13429 (N_13429,N_13199,N_13208);
nor U13430 (N_13430,N_13237,N_13221);
or U13431 (N_13431,N_13238,N_13181);
nand U13432 (N_13432,N_13120,N_13155);
or U13433 (N_13433,N_13015,N_13077);
nor U13434 (N_13434,N_13088,N_13155);
and U13435 (N_13435,N_13041,N_13230);
and U13436 (N_13436,N_13075,N_13039);
and U13437 (N_13437,N_13246,N_13059);
nand U13438 (N_13438,N_13204,N_13235);
and U13439 (N_13439,N_13141,N_13106);
nand U13440 (N_13440,N_13147,N_13137);
and U13441 (N_13441,N_13153,N_13057);
and U13442 (N_13442,N_13071,N_13021);
nand U13443 (N_13443,N_13241,N_13182);
or U13444 (N_13444,N_13073,N_13213);
nand U13445 (N_13445,N_13096,N_13015);
and U13446 (N_13446,N_13043,N_13126);
or U13447 (N_13447,N_13070,N_13124);
and U13448 (N_13448,N_13085,N_13139);
nor U13449 (N_13449,N_13148,N_13100);
and U13450 (N_13450,N_13179,N_13185);
nor U13451 (N_13451,N_13189,N_13178);
xnor U13452 (N_13452,N_13156,N_13240);
nor U13453 (N_13453,N_13083,N_13203);
nand U13454 (N_13454,N_13218,N_13176);
nor U13455 (N_13455,N_13126,N_13016);
nor U13456 (N_13456,N_13142,N_13147);
and U13457 (N_13457,N_13036,N_13108);
nand U13458 (N_13458,N_13174,N_13064);
xor U13459 (N_13459,N_13239,N_13039);
nor U13460 (N_13460,N_13053,N_13236);
nor U13461 (N_13461,N_13130,N_13131);
or U13462 (N_13462,N_13002,N_13150);
xnor U13463 (N_13463,N_13233,N_13025);
xor U13464 (N_13464,N_13170,N_13213);
or U13465 (N_13465,N_13010,N_13113);
nand U13466 (N_13466,N_13024,N_13019);
and U13467 (N_13467,N_13069,N_13219);
nor U13468 (N_13468,N_13062,N_13211);
and U13469 (N_13469,N_13110,N_13122);
nor U13470 (N_13470,N_13180,N_13200);
or U13471 (N_13471,N_13144,N_13218);
or U13472 (N_13472,N_13086,N_13177);
and U13473 (N_13473,N_13007,N_13189);
nand U13474 (N_13474,N_13136,N_13191);
nor U13475 (N_13475,N_13068,N_13146);
nor U13476 (N_13476,N_13137,N_13240);
nand U13477 (N_13477,N_13200,N_13043);
xnor U13478 (N_13478,N_13213,N_13091);
nand U13479 (N_13479,N_13238,N_13172);
nand U13480 (N_13480,N_13105,N_13227);
nor U13481 (N_13481,N_13123,N_13023);
xor U13482 (N_13482,N_13139,N_13110);
nor U13483 (N_13483,N_13138,N_13151);
and U13484 (N_13484,N_13233,N_13003);
xor U13485 (N_13485,N_13199,N_13227);
and U13486 (N_13486,N_13007,N_13155);
nand U13487 (N_13487,N_13055,N_13147);
and U13488 (N_13488,N_13059,N_13097);
and U13489 (N_13489,N_13026,N_13016);
xor U13490 (N_13490,N_13030,N_13137);
or U13491 (N_13491,N_13193,N_13201);
nand U13492 (N_13492,N_13053,N_13216);
or U13493 (N_13493,N_13147,N_13070);
nor U13494 (N_13494,N_13041,N_13167);
and U13495 (N_13495,N_13206,N_13105);
nand U13496 (N_13496,N_13100,N_13241);
nor U13497 (N_13497,N_13148,N_13212);
or U13498 (N_13498,N_13044,N_13050);
nand U13499 (N_13499,N_13236,N_13005);
or U13500 (N_13500,N_13311,N_13465);
nand U13501 (N_13501,N_13369,N_13476);
nor U13502 (N_13502,N_13336,N_13497);
nor U13503 (N_13503,N_13484,N_13331);
nor U13504 (N_13504,N_13393,N_13401);
nor U13505 (N_13505,N_13489,N_13410);
and U13506 (N_13506,N_13304,N_13335);
nand U13507 (N_13507,N_13288,N_13388);
and U13508 (N_13508,N_13409,N_13290);
and U13509 (N_13509,N_13265,N_13271);
or U13510 (N_13510,N_13360,N_13491);
xnor U13511 (N_13511,N_13306,N_13418);
and U13512 (N_13512,N_13408,N_13332);
nand U13513 (N_13513,N_13439,N_13452);
nor U13514 (N_13514,N_13350,N_13414);
xor U13515 (N_13515,N_13253,N_13425);
and U13516 (N_13516,N_13457,N_13260);
and U13517 (N_13517,N_13250,N_13405);
nor U13518 (N_13518,N_13477,N_13321);
or U13519 (N_13519,N_13356,N_13424);
nand U13520 (N_13520,N_13313,N_13376);
or U13521 (N_13521,N_13381,N_13257);
xnor U13522 (N_13522,N_13458,N_13494);
or U13523 (N_13523,N_13454,N_13286);
and U13524 (N_13524,N_13415,N_13363);
and U13525 (N_13525,N_13298,N_13374);
and U13526 (N_13526,N_13398,N_13432);
and U13527 (N_13527,N_13428,N_13462);
xor U13528 (N_13528,N_13366,N_13268);
and U13529 (N_13529,N_13362,N_13277);
and U13530 (N_13530,N_13389,N_13478);
nand U13531 (N_13531,N_13481,N_13404);
or U13532 (N_13532,N_13364,N_13365);
xor U13533 (N_13533,N_13334,N_13443);
and U13534 (N_13534,N_13254,N_13479);
or U13535 (N_13535,N_13347,N_13296);
and U13536 (N_13536,N_13352,N_13324);
nor U13537 (N_13537,N_13303,N_13498);
nand U13538 (N_13538,N_13323,N_13377);
and U13539 (N_13539,N_13270,N_13278);
or U13540 (N_13540,N_13289,N_13480);
and U13541 (N_13541,N_13444,N_13280);
and U13542 (N_13542,N_13293,N_13499);
or U13543 (N_13543,N_13252,N_13421);
or U13544 (N_13544,N_13433,N_13463);
nor U13545 (N_13545,N_13281,N_13383);
nor U13546 (N_13546,N_13263,N_13272);
nand U13547 (N_13547,N_13372,N_13367);
or U13548 (N_13548,N_13468,N_13385);
nand U13549 (N_13549,N_13403,N_13422);
and U13550 (N_13550,N_13450,N_13420);
nand U13551 (N_13551,N_13431,N_13305);
nand U13552 (N_13552,N_13451,N_13449);
or U13553 (N_13553,N_13387,N_13346);
or U13554 (N_13554,N_13283,N_13308);
xnor U13555 (N_13555,N_13442,N_13392);
nor U13556 (N_13556,N_13291,N_13474);
or U13557 (N_13557,N_13416,N_13292);
or U13558 (N_13558,N_13391,N_13340);
or U13559 (N_13559,N_13373,N_13471);
and U13560 (N_13560,N_13485,N_13475);
and U13561 (N_13561,N_13371,N_13267);
nand U13562 (N_13562,N_13456,N_13294);
xnor U13563 (N_13563,N_13353,N_13368);
nand U13564 (N_13564,N_13255,N_13328);
nor U13565 (N_13565,N_13406,N_13466);
nand U13566 (N_13566,N_13329,N_13397);
xor U13567 (N_13567,N_13488,N_13486);
and U13568 (N_13568,N_13354,N_13445);
nor U13569 (N_13569,N_13297,N_13417);
nand U13570 (N_13570,N_13258,N_13345);
or U13571 (N_13571,N_13279,N_13349);
nor U13572 (N_13572,N_13423,N_13317);
or U13573 (N_13573,N_13419,N_13438);
and U13574 (N_13574,N_13256,N_13310);
or U13575 (N_13575,N_13327,N_13251);
nand U13576 (N_13576,N_13487,N_13436);
and U13577 (N_13577,N_13446,N_13435);
nor U13578 (N_13578,N_13273,N_13276);
xor U13579 (N_13579,N_13390,N_13427);
nor U13580 (N_13580,N_13312,N_13274);
nor U13581 (N_13581,N_13300,N_13453);
and U13582 (N_13582,N_13259,N_13315);
or U13583 (N_13583,N_13299,N_13316);
nor U13584 (N_13584,N_13266,N_13430);
nand U13585 (N_13585,N_13341,N_13295);
or U13586 (N_13586,N_13412,N_13429);
and U13587 (N_13587,N_13492,N_13382);
and U13588 (N_13588,N_13496,N_13459);
nor U13589 (N_13589,N_13396,N_13322);
and U13590 (N_13590,N_13284,N_13482);
and U13591 (N_13591,N_13455,N_13394);
or U13592 (N_13592,N_13490,N_13287);
xnor U13593 (N_13593,N_13302,N_13344);
or U13594 (N_13594,N_13309,N_13307);
nor U13595 (N_13595,N_13264,N_13441);
or U13596 (N_13596,N_13275,N_13469);
xnor U13597 (N_13597,N_13342,N_13285);
nor U13598 (N_13598,N_13282,N_13337);
xnor U13599 (N_13599,N_13378,N_13318);
nand U13600 (N_13600,N_13361,N_13357);
or U13601 (N_13601,N_13437,N_13262);
nand U13602 (N_13602,N_13325,N_13330);
nand U13603 (N_13603,N_13269,N_13339);
and U13604 (N_13604,N_13375,N_13380);
or U13605 (N_13605,N_13402,N_13395);
nor U13606 (N_13606,N_13470,N_13434);
and U13607 (N_13607,N_13413,N_13355);
nor U13608 (N_13608,N_13379,N_13461);
and U13609 (N_13609,N_13464,N_13261);
nand U13610 (N_13610,N_13333,N_13343);
nor U13611 (N_13611,N_13472,N_13460);
nor U13612 (N_13612,N_13358,N_13301);
xor U13613 (N_13613,N_13351,N_13386);
and U13614 (N_13614,N_13384,N_13399);
nor U13615 (N_13615,N_13448,N_13407);
and U13616 (N_13616,N_13338,N_13447);
nand U13617 (N_13617,N_13483,N_13314);
and U13618 (N_13618,N_13493,N_13440);
and U13619 (N_13619,N_13348,N_13473);
nor U13620 (N_13620,N_13359,N_13495);
nand U13621 (N_13621,N_13370,N_13326);
xnor U13622 (N_13622,N_13319,N_13426);
or U13623 (N_13623,N_13467,N_13400);
nand U13624 (N_13624,N_13411,N_13320);
and U13625 (N_13625,N_13308,N_13497);
nor U13626 (N_13626,N_13295,N_13314);
nand U13627 (N_13627,N_13392,N_13378);
or U13628 (N_13628,N_13342,N_13331);
or U13629 (N_13629,N_13263,N_13425);
nand U13630 (N_13630,N_13302,N_13398);
nor U13631 (N_13631,N_13253,N_13381);
nor U13632 (N_13632,N_13293,N_13262);
or U13633 (N_13633,N_13322,N_13300);
or U13634 (N_13634,N_13349,N_13495);
or U13635 (N_13635,N_13419,N_13341);
nor U13636 (N_13636,N_13442,N_13271);
or U13637 (N_13637,N_13271,N_13474);
nand U13638 (N_13638,N_13455,N_13347);
xnor U13639 (N_13639,N_13285,N_13369);
or U13640 (N_13640,N_13496,N_13451);
and U13641 (N_13641,N_13286,N_13323);
nand U13642 (N_13642,N_13317,N_13498);
xor U13643 (N_13643,N_13413,N_13313);
nor U13644 (N_13644,N_13290,N_13273);
nand U13645 (N_13645,N_13374,N_13329);
nand U13646 (N_13646,N_13496,N_13443);
and U13647 (N_13647,N_13358,N_13304);
xnor U13648 (N_13648,N_13330,N_13283);
nor U13649 (N_13649,N_13334,N_13264);
and U13650 (N_13650,N_13386,N_13442);
and U13651 (N_13651,N_13487,N_13291);
nand U13652 (N_13652,N_13275,N_13497);
and U13653 (N_13653,N_13449,N_13287);
nand U13654 (N_13654,N_13495,N_13257);
and U13655 (N_13655,N_13485,N_13447);
or U13656 (N_13656,N_13439,N_13263);
or U13657 (N_13657,N_13309,N_13378);
and U13658 (N_13658,N_13381,N_13447);
and U13659 (N_13659,N_13370,N_13420);
or U13660 (N_13660,N_13323,N_13345);
or U13661 (N_13661,N_13367,N_13466);
and U13662 (N_13662,N_13389,N_13432);
nand U13663 (N_13663,N_13391,N_13343);
nor U13664 (N_13664,N_13252,N_13264);
nand U13665 (N_13665,N_13376,N_13356);
nand U13666 (N_13666,N_13289,N_13285);
and U13667 (N_13667,N_13378,N_13450);
and U13668 (N_13668,N_13359,N_13278);
xnor U13669 (N_13669,N_13399,N_13347);
or U13670 (N_13670,N_13441,N_13356);
xor U13671 (N_13671,N_13368,N_13255);
or U13672 (N_13672,N_13389,N_13281);
nor U13673 (N_13673,N_13469,N_13450);
or U13674 (N_13674,N_13283,N_13294);
xor U13675 (N_13675,N_13452,N_13376);
or U13676 (N_13676,N_13316,N_13497);
or U13677 (N_13677,N_13315,N_13474);
or U13678 (N_13678,N_13455,N_13415);
and U13679 (N_13679,N_13462,N_13251);
or U13680 (N_13680,N_13264,N_13339);
xor U13681 (N_13681,N_13434,N_13356);
and U13682 (N_13682,N_13265,N_13439);
nor U13683 (N_13683,N_13273,N_13319);
nor U13684 (N_13684,N_13272,N_13460);
nor U13685 (N_13685,N_13480,N_13397);
or U13686 (N_13686,N_13364,N_13336);
nand U13687 (N_13687,N_13329,N_13424);
or U13688 (N_13688,N_13438,N_13493);
or U13689 (N_13689,N_13345,N_13336);
and U13690 (N_13690,N_13470,N_13339);
nand U13691 (N_13691,N_13491,N_13264);
or U13692 (N_13692,N_13296,N_13448);
and U13693 (N_13693,N_13374,N_13438);
or U13694 (N_13694,N_13476,N_13459);
nand U13695 (N_13695,N_13296,N_13315);
or U13696 (N_13696,N_13301,N_13334);
and U13697 (N_13697,N_13300,N_13347);
or U13698 (N_13698,N_13453,N_13371);
nor U13699 (N_13699,N_13443,N_13478);
or U13700 (N_13700,N_13321,N_13423);
nand U13701 (N_13701,N_13335,N_13281);
nor U13702 (N_13702,N_13335,N_13302);
nor U13703 (N_13703,N_13324,N_13319);
or U13704 (N_13704,N_13426,N_13254);
or U13705 (N_13705,N_13422,N_13261);
and U13706 (N_13706,N_13490,N_13462);
nand U13707 (N_13707,N_13272,N_13368);
nor U13708 (N_13708,N_13394,N_13372);
or U13709 (N_13709,N_13261,N_13406);
or U13710 (N_13710,N_13490,N_13318);
nor U13711 (N_13711,N_13357,N_13399);
xnor U13712 (N_13712,N_13405,N_13449);
nor U13713 (N_13713,N_13479,N_13333);
or U13714 (N_13714,N_13384,N_13493);
or U13715 (N_13715,N_13307,N_13490);
or U13716 (N_13716,N_13328,N_13296);
or U13717 (N_13717,N_13348,N_13486);
and U13718 (N_13718,N_13312,N_13479);
nand U13719 (N_13719,N_13369,N_13493);
nand U13720 (N_13720,N_13342,N_13470);
or U13721 (N_13721,N_13431,N_13373);
nand U13722 (N_13722,N_13470,N_13453);
and U13723 (N_13723,N_13318,N_13344);
xor U13724 (N_13724,N_13250,N_13387);
nand U13725 (N_13725,N_13453,N_13414);
nor U13726 (N_13726,N_13307,N_13491);
or U13727 (N_13727,N_13377,N_13303);
or U13728 (N_13728,N_13350,N_13391);
nand U13729 (N_13729,N_13387,N_13287);
nand U13730 (N_13730,N_13429,N_13326);
nor U13731 (N_13731,N_13307,N_13419);
nor U13732 (N_13732,N_13298,N_13268);
or U13733 (N_13733,N_13277,N_13343);
nor U13734 (N_13734,N_13274,N_13478);
xnor U13735 (N_13735,N_13372,N_13381);
nor U13736 (N_13736,N_13328,N_13410);
nand U13737 (N_13737,N_13336,N_13365);
or U13738 (N_13738,N_13487,N_13351);
nor U13739 (N_13739,N_13477,N_13462);
nor U13740 (N_13740,N_13331,N_13470);
or U13741 (N_13741,N_13437,N_13469);
or U13742 (N_13742,N_13449,N_13482);
and U13743 (N_13743,N_13491,N_13467);
xnor U13744 (N_13744,N_13279,N_13483);
nor U13745 (N_13745,N_13368,N_13454);
nor U13746 (N_13746,N_13489,N_13351);
nand U13747 (N_13747,N_13313,N_13361);
nor U13748 (N_13748,N_13414,N_13346);
and U13749 (N_13749,N_13270,N_13348);
nand U13750 (N_13750,N_13704,N_13652);
or U13751 (N_13751,N_13733,N_13570);
xor U13752 (N_13752,N_13666,N_13727);
or U13753 (N_13753,N_13639,N_13675);
and U13754 (N_13754,N_13636,N_13577);
or U13755 (N_13755,N_13564,N_13695);
and U13756 (N_13756,N_13690,N_13615);
nor U13757 (N_13757,N_13614,N_13606);
nor U13758 (N_13758,N_13519,N_13559);
nor U13759 (N_13759,N_13589,N_13629);
or U13760 (N_13760,N_13503,N_13693);
or U13761 (N_13761,N_13571,N_13644);
nand U13762 (N_13762,N_13598,N_13719);
xor U13763 (N_13763,N_13726,N_13696);
and U13764 (N_13764,N_13676,N_13712);
and U13765 (N_13765,N_13720,N_13545);
or U13766 (N_13766,N_13707,N_13534);
and U13767 (N_13767,N_13584,N_13647);
nand U13768 (N_13768,N_13583,N_13731);
and U13769 (N_13769,N_13670,N_13531);
nor U13770 (N_13770,N_13607,N_13723);
nor U13771 (N_13771,N_13658,N_13625);
nand U13772 (N_13772,N_13743,N_13595);
nor U13773 (N_13773,N_13588,N_13590);
and U13774 (N_13774,N_13669,N_13725);
nand U13775 (N_13775,N_13691,N_13515);
and U13776 (N_13776,N_13527,N_13558);
or U13777 (N_13777,N_13543,N_13643);
and U13778 (N_13778,N_13701,N_13742);
nor U13779 (N_13779,N_13721,N_13679);
nor U13780 (N_13780,N_13506,N_13568);
and U13781 (N_13781,N_13600,N_13610);
and U13782 (N_13782,N_13623,N_13664);
xnor U13783 (N_13783,N_13548,N_13594);
xor U13784 (N_13784,N_13737,N_13672);
nand U13785 (N_13785,N_13605,N_13582);
and U13786 (N_13786,N_13668,N_13619);
nand U13787 (N_13787,N_13654,N_13523);
nand U13788 (N_13788,N_13551,N_13550);
nor U13789 (N_13789,N_13706,N_13536);
nand U13790 (N_13790,N_13716,N_13710);
or U13791 (N_13791,N_13509,N_13674);
nor U13792 (N_13792,N_13673,N_13626);
nor U13793 (N_13793,N_13732,N_13524);
and U13794 (N_13794,N_13697,N_13662);
xnor U13795 (N_13795,N_13546,N_13596);
and U13796 (N_13796,N_13717,N_13741);
nor U13797 (N_13797,N_13572,N_13659);
and U13798 (N_13798,N_13702,N_13665);
nand U13799 (N_13799,N_13580,N_13628);
or U13800 (N_13800,N_13698,N_13516);
and U13801 (N_13801,N_13530,N_13533);
nor U13802 (N_13802,N_13542,N_13620);
nor U13803 (N_13803,N_13526,N_13556);
nor U13804 (N_13804,N_13535,N_13729);
nand U13805 (N_13805,N_13681,N_13554);
nor U13806 (N_13806,N_13512,N_13624);
nand U13807 (N_13807,N_13529,N_13688);
or U13808 (N_13808,N_13603,N_13569);
or U13809 (N_13809,N_13648,N_13663);
and U13810 (N_13810,N_13678,N_13514);
and U13811 (N_13811,N_13660,N_13521);
or U13812 (N_13812,N_13646,N_13601);
or U13813 (N_13813,N_13632,N_13645);
or U13814 (N_13814,N_13748,N_13642);
nand U13815 (N_13815,N_13520,N_13700);
nor U13816 (N_13816,N_13560,N_13627);
nand U13817 (N_13817,N_13508,N_13692);
or U13818 (N_13818,N_13730,N_13581);
xor U13819 (N_13819,N_13597,N_13504);
and U13820 (N_13820,N_13685,N_13734);
nand U13821 (N_13821,N_13630,N_13576);
nand U13822 (N_13822,N_13746,N_13735);
xnor U13823 (N_13823,N_13714,N_13507);
or U13824 (N_13824,N_13565,N_13552);
and U13825 (N_13825,N_13612,N_13653);
nand U13826 (N_13826,N_13609,N_13703);
or U13827 (N_13827,N_13640,N_13682);
or U13828 (N_13828,N_13745,N_13722);
or U13829 (N_13829,N_13689,N_13709);
nand U13830 (N_13830,N_13541,N_13562);
or U13831 (N_13831,N_13593,N_13537);
nor U13832 (N_13832,N_13747,N_13728);
nand U13833 (N_13833,N_13736,N_13749);
xnor U13834 (N_13834,N_13621,N_13538);
or U13835 (N_13835,N_13680,N_13511);
nand U13836 (N_13836,N_13586,N_13656);
nand U13837 (N_13837,N_13738,N_13677);
xor U13838 (N_13838,N_13574,N_13641);
nor U13839 (N_13839,N_13505,N_13599);
nand U13840 (N_13840,N_13638,N_13502);
xor U13841 (N_13841,N_13667,N_13585);
and U13842 (N_13842,N_13715,N_13522);
nor U13843 (N_13843,N_13724,N_13602);
nand U13844 (N_13844,N_13687,N_13683);
nand U13845 (N_13845,N_13718,N_13557);
nor U13846 (N_13846,N_13711,N_13547);
nor U13847 (N_13847,N_13563,N_13561);
or U13848 (N_13848,N_13573,N_13579);
or U13849 (N_13849,N_13532,N_13528);
nor U13850 (N_13850,N_13555,N_13513);
or U13851 (N_13851,N_13618,N_13635);
and U13852 (N_13852,N_13671,N_13604);
xor U13853 (N_13853,N_13631,N_13661);
nand U13854 (N_13854,N_13501,N_13739);
xnor U13855 (N_13855,N_13611,N_13651);
xnor U13856 (N_13856,N_13740,N_13622);
and U13857 (N_13857,N_13517,N_13566);
xor U13858 (N_13858,N_13713,N_13578);
or U13859 (N_13859,N_13634,N_13657);
nor U13860 (N_13860,N_13694,N_13544);
and U13861 (N_13861,N_13616,N_13613);
xnor U13862 (N_13862,N_13549,N_13518);
nand U13863 (N_13863,N_13684,N_13539);
nand U13864 (N_13864,N_13591,N_13699);
or U13865 (N_13865,N_13744,N_13540);
and U13866 (N_13866,N_13650,N_13655);
xor U13867 (N_13867,N_13510,N_13567);
nor U13868 (N_13868,N_13592,N_13587);
nor U13869 (N_13869,N_13649,N_13608);
nor U13870 (N_13870,N_13705,N_13553);
xor U13871 (N_13871,N_13500,N_13575);
nor U13872 (N_13872,N_13708,N_13637);
nand U13873 (N_13873,N_13525,N_13686);
nand U13874 (N_13874,N_13633,N_13617);
and U13875 (N_13875,N_13651,N_13743);
nand U13876 (N_13876,N_13551,N_13679);
nor U13877 (N_13877,N_13595,N_13736);
or U13878 (N_13878,N_13506,N_13702);
nand U13879 (N_13879,N_13702,N_13658);
nor U13880 (N_13880,N_13633,N_13647);
and U13881 (N_13881,N_13642,N_13719);
nor U13882 (N_13882,N_13580,N_13636);
and U13883 (N_13883,N_13552,N_13606);
nand U13884 (N_13884,N_13666,N_13717);
or U13885 (N_13885,N_13584,N_13615);
nor U13886 (N_13886,N_13631,N_13550);
xnor U13887 (N_13887,N_13677,N_13604);
xor U13888 (N_13888,N_13566,N_13706);
nor U13889 (N_13889,N_13549,N_13603);
nor U13890 (N_13890,N_13746,N_13633);
nand U13891 (N_13891,N_13710,N_13741);
or U13892 (N_13892,N_13516,N_13651);
nor U13893 (N_13893,N_13655,N_13644);
nor U13894 (N_13894,N_13634,N_13692);
nor U13895 (N_13895,N_13534,N_13619);
and U13896 (N_13896,N_13733,N_13742);
or U13897 (N_13897,N_13606,N_13549);
or U13898 (N_13898,N_13738,N_13586);
nand U13899 (N_13899,N_13611,N_13653);
nand U13900 (N_13900,N_13516,N_13676);
or U13901 (N_13901,N_13612,N_13644);
nand U13902 (N_13902,N_13631,N_13584);
nand U13903 (N_13903,N_13643,N_13578);
nor U13904 (N_13904,N_13729,N_13680);
and U13905 (N_13905,N_13701,N_13627);
nand U13906 (N_13906,N_13704,N_13540);
xnor U13907 (N_13907,N_13679,N_13643);
and U13908 (N_13908,N_13565,N_13705);
and U13909 (N_13909,N_13728,N_13605);
nor U13910 (N_13910,N_13585,N_13563);
xor U13911 (N_13911,N_13542,N_13666);
and U13912 (N_13912,N_13659,N_13635);
xor U13913 (N_13913,N_13731,N_13645);
nand U13914 (N_13914,N_13564,N_13579);
nor U13915 (N_13915,N_13716,N_13542);
and U13916 (N_13916,N_13743,N_13663);
nor U13917 (N_13917,N_13616,N_13528);
and U13918 (N_13918,N_13641,N_13640);
and U13919 (N_13919,N_13662,N_13552);
and U13920 (N_13920,N_13532,N_13740);
nor U13921 (N_13921,N_13692,N_13646);
or U13922 (N_13922,N_13660,N_13619);
nor U13923 (N_13923,N_13675,N_13536);
nand U13924 (N_13924,N_13648,N_13650);
xnor U13925 (N_13925,N_13624,N_13605);
and U13926 (N_13926,N_13551,N_13669);
and U13927 (N_13927,N_13519,N_13625);
nor U13928 (N_13928,N_13677,N_13691);
xnor U13929 (N_13929,N_13698,N_13749);
nor U13930 (N_13930,N_13646,N_13662);
xor U13931 (N_13931,N_13649,N_13653);
nand U13932 (N_13932,N_13676,N_13605);
nand U13933 (N_13933,N_13615,N_13694);
nor U13934 (N_13934,N_13676,N_13571);
xnor U13935 (N_13935,N_13671,N_13503);
nand U13936 (N_13936,N_13728,N_13681);
nand U13937 (N_13937,N_13697,N_13610);
or U13938 (N_13938,N_13701,N_13656);
nor U13939 (N_13939,N_13632,N_13508);
nand U13940 (N_13940,N_13638,N_13579);
and U13941 (N_13941,N_13507,N_13556);
and U13942 (N_13942,N_13505,N_13636);
nand U13943 (N_13943,N_13731,N_13685);
and U13944 (N_13944,N_13614,N_13547);
and U13945 (N_13945,N_13516,N_13662);
nand U13946 (N_13946,N_13740,N_13563);
and U13947 (N_13947,N_13637,N_13660);
or U13948 (N_13948,N_13501,N_13627);
or U13949 (N_13949,N_13690,N_13653);
nand U13950 (N_13950,N_13648,N_13609);
nand U13951 (N_13951,N_13605,N_13682);
and U13952 (N_13952,N_13654,N_13600);
or U13953 (N_13953,N_13577,N_13523);
and U13954 (N_13954,N_13588,N_13748);
nand U13955 (N_13955,N_13649,N_13579);
nand U13956 (N_13956,N_13629,N_13655);
or U13957 (N_13957,N_13538,N_13567);
nand U13958 (N_13958,N_13545,N_13561);
and U13959 (N_13959,N_13543,N_13528);
nor U13960 (N_13960,N_13631,N_13510);
and U13961 (N_13961,N_13528,N_13603);
nor U13962 (N_13962,N_13711,N_13610);
nand U13963 (N_13963,N_13669,N_13538);
or U13964 (N_13964,N_13600,N_13691);
xnor U13965 (N_13965,N_13609,N_13647);
or U13966 (N_13966,N_13591,N_13694);
and U13967 (N_13967,N_13613,N_13505);
nor U13968 (N_13968,N_13541,N_13718);
nor U13969 (N_13969,N_13518,N_13695);
and U13970 (N_13970,N_13723,N_13502);
nor U13971 (N_13971,N_13730,N_13678);
nand U13972 (N_13972,N_13559,N_13631);
and U13973 (N_13973,N_13596,N_13695);
xor U13974 (N_13974,N_13635,N_13693);
and U13975 (N_13975,N_13528,N_13732);
or U13976 (N_13976,N_13726,N_13578);
or U13977 (N_13977,N_13674,N_13681);
nand U13978 (N_13978,N_13554,N_13744);
or U13979 (N_13979,N_13508,N_13573);
nand U13980 (N_13980,N_13686,N_13733);
or U13981 (N_13981,N_13689,N_13719);
xnor U13982 (N_13982,N_13555,N_13607);
and U13983 (N_13983,N_13710,N_13717);
xor U13984 (N_13984,N_13611,N_13691);
or U13985 (N_13985,N_13646,N_13548);
or U13986 (N_13986,N_13668,N_13565);
nand U13987 (N_13987,N_13680,N_13507);
or U13988 (N_13988,N_13712,N_13610);
or U13989 (N_13989,N_13590,N_13744);
or U13990 (N_13990,N_13713,N_13580);
and U13991 (N_13991,N_13596,N_13563);
nor U13992 (N_13992,N_13737,N_13522);
nor U13993 (N_13993,N_13675,N_13703);
or U13994 (N_13994,N_13725,N_13502);
nor U13995 (N_13995,N_13601,N_13561);
nand U13996 (N_13996,N_13548,N_13629);
and U13997 (N_13997,N_13615,N_13565);
xor U13998 (N_13998,N_13542,N_13623);
and U13999 (N_13999,N_13742,N_13559);
nand U14000 (N_14000,N_13999,N_13963);
nand U14001 (N_14001,N_13959,N_13898);
nand U14002 (N_14002,N_13965,N_13975);
nor U14003 (N_14003,N_13945,N_13765);
and U14004 (N_14004,N_13946,N_13978);
nand U14005 (N_14005,N_13914,N_13873);
nand U14006 (N_14006,N_13922,N_13821);
nand U14007 (N_14007,N_13795,N_13984);
or U14008 (N_14008,N_13957,N_13920);
and U14009 (N_14009,N_13871,N_13993);
or U14010 (N_14010,N_13777,N_13900);
nand U14011 (N_14011,N_13919,N_13915);
nor U14012 (N_14012,N_13980,N_13880);
or U14013 (N_14013,N_13787,N_13952);
nand U14014 (N_14014,N_13867,N_13961);
nand U14015 (N_14015,N_13889,N_13947);
or U14016 (N_14016,N_13790,N_13771);
and U14017 (N_14017,N_13837,N_13971);
or U14018 (N_14018,N_13904,N_13996);
nor U14019 (N_14019,N_13859,N_13995);
and U14020 (N_14020,N_13877,N_13903);
xnor U14021 (N_14021,N_13912,N_13878);
nand U14022 (N_14022,N_13936,N_13908);
xnor U14023 (N_14023,N_13809,N_13778);
and U14024 (N_14024,N_13933,N_13817);
nand U14025 (N_14025,N_13813,N_13940);
and U14026 (N_14026,N_13949,N_13766);
or U14027 (N_14027,N_13774,N_13960);
nand U14028 (N_14028,N_13828,N_13966);
nor U14029 (N_14029,N_13868,N_13769);
nand U14030 (N_14030,N_13927,N_13930);
nand U14031 (N_14031,N_13982,N_13841);
or U14032 (N_14032,N_13845,N_13954);
nand U14033 (N_14033,N_13779,N_13754);
or U14034 (N_14034,N_13901,N_13872);
nand U14035 (N_14035,N_13796,N_13881);
and U14036 (N_14036,N_13836,N_13921);
xnor U14037 (N_14037,N_13770,N_13789);
nor U14038 (N_14038,N_13998,N_13833);
or U14039 (N_14039,N_13792,N_13929);
nor U14040 (N_14040,N_13994,N_13839);
and U14041 (N_14041,N_13838,N_13879);
nand U14042 (N_14042,N_13857,N_13970);
nor U14043 (N_14043,N_13955,N_13764);
nand U14044 (N_14044,N_13870,N_13938);
or U14045 (N_14045,N_13884,N_13798);
and U14046 (N_14046,N_13799,N_13866);
xnor U14047 (N_14047,N_13926,N_13829);
or U14048 (N_14048,N_13784,N_13823);
nor U14049 (N_14049,N_13953,N_13899);
or U14050 (N_14050,N_13834,N_13827);
nand U14051 (N_14051,N_13830,N_13756);
xor U14052 (N_14052,N_13819,N_13917);
xnor U14053 (N_14053,N_13810,N_13925);
and U14054 (N_14054,N_13928,N_13939);
or U14055 (N_14055,N_13761,N_13869);
and U14056 (N_14056,N_13846,N_13876);
nor U14057 (N_14057,N_13956,N_13805);
nor U14058 (N_14058,N_13976,N_13825);
nand U14059 (N_14059,N_13986,N_13785);
or U14060 (N_14060,N_13814,N_13797);
and U14061 (N_14061,N_13931,N_13840);
and U14062 (N_14062,N_13985,N_13818);
nor U14063 (N_14063,N_13832,N_13969);
nand U14064 (N_14064,N_13782,N_13944);
and U14065 (N_14065,N_13831,N_13895);
or U14066 (N_14066,N_13786,N_13794);
and U14067 (N_14067,N_13972,N_13842);
or U14068 (N_14068,N_13806,N_13775);
nand U14069 (N_14069,N_13891,N_13916);
nand U14070 (N_14070,N_13791,N_13804);
or U14071 (N_14071,N_13820,N_13850);
nand U14072 (N_14072,N_13835,N_13997);
or U14073 (N_14073,N_13896,N_13865);
or U14074 (N_14074,N_13948,N_13853);
or U14075 (N_14075,N_13801,N_13780);
or U14076 (N_14076,N_13907,N_13934);
and U14077 (N_14077,N_13852,N_13849);
or U14078 (N_14078,N_13812,N_13860);
nor U14079 (N_14079,N_13824,N_13958);
and U14080 (N_14080,N_13760,N_13894);
nor U14081 (N_14081,N_13882,N_13807);
or U14082 (N_14082,N_13858,N_13808);
nand U14083 (N_14083,N_13755,N_13815);
nand U14084 (N_14084,N_13773,N_13855);
or U14085 (N_14085,N_13793,N_13757);
and U14086 (N_14086,N_13967,N_13803);
nor U14087 (N_14087,N_13935,N_13883);
and U14088 (N_14088,N_13950,N_13800);
nand U14089 (N_14089,N_13826,N_13979);
nor U14090 (N_14090,N_13816,N_13753);
or U14091 (N_14091,N_13943,N_13888);
nand U14092 (N_14092,N_13759,N_13863);
xor U14093 (N_14093,N_13856,N_13981);
nor U14094 (N_14094,N_13767,N_13968);
nand U14095 (N_14095,N_13751,N_13851);
nand U14096 (N_14096,N_13750,N_13758);
nor U14097 (N_14097,N_13974,N_13862);
nand U14098 (N_14098,N_13892,N_13875);
and U14099 (N_14099,N_13991,N_13977);
and U14100 (N_14100,N_13923,N_13848);
nand U14101 (N_14101,N_13890,N_13781);
nor U14102 (N_14102,N_13788,N_13918);
or U14103 (N_14103,N_13990,N_13763);
and U14104 (N_14104,N_13905,N_13886);
and U14105 (N_14105,N_13989,N_13893);
nand U14106 (N_14106,N_13902,N_13874);
nor U14107 (N_14107,N_13861,N_13962);
xnor U14108 (N_14108,N_13897,N_13941);
and U14109 (N_14109,N_13924,N_13776);
or U14110 (N_14110,N_13887,N_13762);
or U14111 (N_14111,N_13911,N_13772);
or U14112 (N_14112,N_13847,N_13854);
nor U14113 (N_14113,N_13987,N_13864);
nand U14114 (N_14114,N_13906,N_13983);
nand U14115 (N_14115,N_13783,N_13811);
or U14116 (N_14116,N_13843,N_13822);
nor U14117 (N_14117,N_13802,N_13910);
nor U14118 (N_14118,N_13913,N_13885);
nand U14119 (N_14119,N_13937,N_13992);
nor U14120 (N_14120,N_13973,N_13768);
nand U14121 (N_14121,N_13988,N_13964);
and U14122 (N_14122,N_13951,N_13942);
or U14123 (N_14123,N_13844,N_13752);
and U14124 (N_14124,N_13932,N_13909);
nand U14125 (N_14125,N_13947,N_13877);
and U14126 (N_14126,N_13931,N_13921);
nor U14127 (N_14127,N_13947,N_13890);
nand U14128 (N_14128,N_13911,N_13811);
xnor U14129 (N_14129,N_13837,N_13910);
nor U14130 (N_14130,N_13804,N_13829);
and U14131 (N_14131,N_13839,N_13798);
and U14132 (N_14132,N_13993,N_13963);
and U14133 (N_14133,N_13833,N_13873);
or U14134 (N_14134,N_13764,N_13896);
or U14135 (N_14135,N_13932,N_13872);
and U14136 (N_14136,N_13882,N_13948);
and U14137 (N_14137,N_13871,N_13890);
nor U14138 (N_14138,N_13865,N_13755);
or U14139 (N_14139,N_13759,N_13778);
or U14140 (N_14140,N_13948,N_13918);
nand U14141 (N_14141,N_13760,N_13897);
or U14142 (N_14142,N_13997,N_13977);
nand U14143 (N_14143,N_13939,N_13816);
or U14144 (N_14144,N_13884,N_13834);
xnor U14145 (N_14145,N_13796,N_13830);
nand U14146 (N_14146,N_13889,N_13922);
nor U14147 (N_14147,N_13959,N_13962);
xor U14148 (N_14148,N_13755,N_13903);
and U14149 (N_14149,N_13958,N_13861);
nand U14150 (N_14150,N_13769,N_13938);
xor U14151 (N_14151,N_13784,N_13753);
and U14152 (N_14152,N_13761,N_13853);
nor U14153 (N_14153,N_13851,N_13983);
xnor U14154 (N_14154,N_13982,N_13761);
or U14155 (N_14155,N_13964,N_13843);
nand U14156 (N_14156,N_13898,N_13893);
and U14157 (N_14157,N_13833,N_13926);
and U14158 (N_14158,N_13963,N_13878);
nand U14159 (N_14159,N_13825,N_13922);
and U14160 (N_14160,N_13761,N_13827);
and U14161 (N_14161,N_13780,N_13900);
or U14162 (N_14162,N_13994,N_13984);
and U14163 (N_14163,N_13939,N_13967);
or U14164 (N_14164,N_13982,N_13837);
or U14165 (N_14165,N_13892,N_13832);
and U14166 (N_14166,N_13810,N_13990);
and U14167 (N_14167,N_13806,N_13825);
nand U14168 (N_14168,N_13944,N_13791);
or U14169 (N_14169,N_13905,N_13917);
nor U14170 (N_14170,N_13858,N_13769);
and U14171 (N_14171,N_13925,N_13885);
or U14172 (N_14172,N_13861,N_13922);
and U14173 (N_14173,N_13832,N_13866);
xnor U14174 (N_14174,N_13857,N_13895);
and U14175 (N_14175,N_13891,N_13859);
nand U14176 (N_14176,N_13998,N_13822);
nor U14177 (N_14177,N_13753,N_13991);
nor U14178 (N_14178,N_13839,N_13902);
nor U14179 (N_14179,N_13901,N_13755);
or U14180 (N_14180,N_13839,N_13880);
xor U14181 (N_14181,N_13871,N_13824);
nand U14182 (N_14182,N_13856,N_13945);
and U14183 (N_14183,N_13794,N_13827);
and U14184 (N_14184,N_13964,N_13855);
or U14185 (N_14185,N_13873,N_13776);
and U14186 (N_14186,N_13985,N_13942);
or U14187 (N_14187,N_13770,N_13758);
and U14188 (N_14188,N_13958,N_13911);
nand U14189 (N_14189,N_13792,N_13882);
xnor U14190 (N_14190,N_13777,N_13869);
and U14191 (N_14191,N_13871,N_13813);
or U14192 (N_14192,N_13766,N_13936);
xnor U14193 (N_14193,N_13901,N_13871);
and U14194 (N_14194,N_13954,N_13767);
xor U14195 (N_14195,N_13892,N_13837);
nor U14196 (N_14196,N_13801,N_13895);
nor U14197 (N_14197,N_13839,N_13780);
nand U14198 (N_14198,N_13945,N_13850);
and U14199 (N_14199,N_13921,N_13794);
and U14200 (N_14200,N_13888,N_13904);
nand U14201 (N_14201,N_13864,N_13847);
and U14202 (N_14202,N_13978,N_13800);
or U14203 (N_14203,N_13866,N_13761);
or U14204 (N_14204,N_13944,N_13922);
or U14205 (N_14205,N_13896,N_13824);
nor U14206 (N_14206,N_13764,N_13915);
or U14207 (N_14207,N_13816,N_13833);
nand U14208 (N_14208,N_13838,N_13803);
nand U14209 (N_14209,N_13909,N_13800);
nand U14210 (N_14210,N_13903,N_13953);
and U14211 (N_14211,N_13767,N_13875);
and U14212 (N_14212,N_13774,N_13989);
nor U14213 (N_14213,N_13794,N_13760);
nand U14214 (N_14214,N_13806,N_13803);
nand U14215 (N_14215,N_13987,N_13870);
and U14216 (N_14216,N_13885,N_13837);
nand U14217 (N_14217,N_13769,N_13985);
nor U14218 (N_14218,N_13811,N_13980);
nor U14219 (N_14219,N_13820,N_13782);
xnor U14220 (N_14220,N_13810,N_13849);
or U14221 (N_14221,N_13932,N_13777);
and U14222 (N_14222,N_13754,N_13891);
or U14223 (N_14223,N_13988,N_13768);
nor U14224 (N_14224,N_13897,N_13908);
nand U14225 (N_14225,N_13905,N_13803);
nand U14226 (N_14226,N_13779,N_13845);
nand U14227 (N_14227,N_13978,N_13890);
nor U14228 (N_14228,N_13989,N_13807);
nor U14229 (N_14229,N_13953,N_13873);
and U14230 (N_14230,N_13775,N_13963);
nand U14231 (N_14231,N_13985,N_13792);
nor U14232 (N_14232,N_13956,N_13936);
nor U14233 (N_14233,N_13897,N_13961);
xor U14234 (N_14234,N_13994,N_13821);
nand U14235 (N_14235,N_13866,N_13865);
nor U14236 (N_14236,N_13827,N_13777);
or U14237 (N_14237,N_13985,N_13805);
or U14238 (N_14238,N_13870,N_13965);
nand U14239 (N_14239,N_13824,N_13964);
or U14240 (N_14240,N_13917,N_13953);
and U14241 (N_14241,N_13857,N_13903);
and U14242 (N_14242,N_13925,N_13984);
or U14243 (N_14243,N_13934,N_13799);
or U14244 (N_14244,N_13942,N_13871);
or U14245 (N_14245,N_13838,N_13866);
and U14246 (N_14246,N_13910,N_13971);
xnor U14247 (N_14247,N_13858,N_13953);
or U14248 (N_14248,N_13880,N_13904);
or U14249 (N_14249,N_13961,N_13892);
nand U14250 (N_14250,N_14014,N_14103);
and U14251 (N_14251,N_14046,N_14033);
xnor U14252 (N_14252,N_14110,N_14232);
or U14253 (N_14253,N_14093,N_14116);
and U14254 (N_14254,N_14109,N_14023);
nand U14255 (N_14255,N_14215,N_14170);
or U14256 (N_14256,N_14231,N_14101);
or U14257 (N_14257,N_14107,N_14187);
and U14258 (N_14258,N_14088,N_14239);
or U14259 (N_14259,N_14063,N_14171);
xnor U14260 (N_14260,N_14245,N_14080);
nor U14261 (N_14261,N_14055,N_14237);
and U14262 (N_14262,N_14203,N_14135);
nand U14263 (N_14263,N_14013,N_14005);
or U14264 (N_14264,N_14126,N_14027);
xor U14265 (N_14265,N_14053,N_14037);
nor U14266 (N_14266,N_14190,N_14102);
and U14267 (N_14267,N_14029,N_14106);
and U14268 (N_14268,N_14087,N_14158);
or U14269 (N_14269,N_14057,N_14092);
nor U14270 (N_14270,N_14097,N_14207);
and U14271 (N_14271,N_14168,N_14175);
and U14272 (N_14272,N_14185,N_14218);
nor U14273 (N_14273,N_14129,N_14241);
nand U14274 (N_14274,N_14018,N_14176);
nand U14275 (N_14275,N_14236,N_14000);
nand U14276 (N_14276,N_14211,N_14049);
nor U14277 (N_14277,N_14073,N_14162);
nor U14278 (N_14278,N_14165,N_14076);
nor U14279 (N_14279,N_14065,N_14086);
nor U14280 (N_14280,N_14172,N_14052);
nand U14281 (N_14281,N_14007,N_14206);
xnor U14282 (N_14282,N_14193,N_14167);
nor U14283 (N_14283,N_14161,N_14138);
nand U14284 (N_14284,N_14079,N_14201);
nor U14285 (N_14285,N_14121,N_14113);
and U14286 (N_14286,N_14226,N_14091);
nand U14287 (N_14287,N_14142,N_14177);
nor U14288 (N_14288,N_14212,N_14009);
or U14289 (N_14289,N_14143,N_14140);
xnor U14290 (N_14290,N_14216,N_14024);
or U14291 (N_14291,N_14221,N_14081);
xnor U14292 (N_14292,N_14146,N_14108);
or U14293 (N_14293,N_14134,N_14072);
xor U14294 (N_14294,N_14032,N_14133);
xor U14295 (N_14295,N_14038,N_14050);
nor U14296 (N_14296,N_14095,N_14249);
nand U14297 (N_14297,N_14229,N_14243);
or U14298 (N_14298,N_14208,N_14213);
or U14299 (N_14299,N_14217,N_14045);
nand U14300 (N_14300,N_14137,N_14228);
and U14301 (N_14301,N_14220,N_14227);
or U14302 (N_14302,N_14136,N_14042);
xnor U14303 (N_14303,N_14010,N_14112);
or U14304 (N_14304,N_14044,N_14059);
nor U14305 (N_14305,N_14130,N_14094);
or U14306 (N_14306,N_14145,N_14122);
and U14307 (N_14307,N_14131,N_14002);
and U14308 (N_14308,N_14124,N_14128);
nor U14309 (N_14309,N_14144,N_14036);
xnor U14310 (N_14310,N_14153,N_14152);
nand U14311 (N_14311,N_14222,N_14047);
nand U14312 (N_14312,N_14031,N_14118);
xnor U14313 (N_14313,N_14008,N_14233);
nand U14314 (N_14314,N_14068,N_14111);
xor U14315 (N_14315,N_14077,N_14182);
nor U14316 (N_14316,N_14085,N_14021);
or U14317 (N_14317,N_14214,N_14141);
nor U14318 (N_14318,N_14240,N_14067);
nor U14319 (N_14319,N_14058,N_14139);
and U14320 (N_14320,N_14003,N_14051);
and U14321 (N_14321,N_14192,N_14189);
xnor U14322 (N_14322,N_14011,N_14040);
nand U14323 (N_14323,N_14075,N_14069);
and U14324 (N_14324,N_14154,N_14209);
and U14325 (N_14325,N_14039,N_14159);
nand U14326 (N_14326,N_14205,N_14117);
nor U14327 (N_14327,N_14166,N_14001);
nor U14328 (N_14328,N_14004,N_14078);
xor U14329 (N_14329,N_14225,N_14160);
or U14330 (N_14330,N_14123,N_14188);
nand U14331 (N_14331,N_14071,N_14016);
or U14332 (N_14332,N_14163,N_14178);
nor U14333 (N_14333,N_14084,N_14025);
nor U14334 (N_14334,N_14061,N_14096);
or U14335 (N_14335,N_14242,N_14089);
and U14336 (N_14336,N_14043,N_14235);
nand U14337 (N_14337,N_14019,N_14132);
nor U14338 (N_14338,N_14186,N_14064);
nor U14339 (N_14339,N_14164,N_14082);
nor U14340 (N_14340,N_14173,N_14184);
nor U14341 (N_14341,N_14174,N_14198);
nand U14342 (N_14342,N_14098,N_14197);
nor U14343 (N_14343,N_14017,N_14156);
and U14344 (N_14344,N_14028,N_14114);
nand U14345 (N_14345,N_14247,N_14204);
and U14346 (N_14346,N_14148,N_14169);
xnor U14347 (N_14347,N_14248,N_14191);
nand U14348 (N_14348,N_14151,N_14066);
or U14349 (N_14349,N_14070,N_14194);
or U14350 (N_14350,N_14041,N_14034);
nand U14351 (N_14351,N_14115,N_14012);
nand U14352 (N_14352,N_14224,N_14099);
nor U14353 (N_14353,N_14149,N_14244);
xnor U14354 (N_14354,N_14210,N_14090);
nand U14355 (N_14355,N_14127,N_14030);
nor U14356 (N_14356,N_14155,N_14074);
nor U14357 (N_14357,N_14181,N_14195);
or U14358 (N_14358,N_14147,N_14100);
xor U14359 (N_14359,N_14035,N_14119);
nor U14360 (N_14360,N_14060,N_14157);
nand U14361 (N_14361,N_14150,N_14202);
or U14362 (N_14362,N_14083,N_14022);
nor U14363 (N_14363,N_14026,N_14199);
and U14364 (N_14364,N_14200,N_14015);
nand U14365 (N_14365,N_14120,N_14006);
and U14366 (N_14366,N_14125,N_14219);
or U14367 (N_14367,N_14246,N_14180);
or U14368 (N_14368,N_14054,N_14056);
nor U14369 (N_14369,N_14223,N_14020);
or U14370 (N_14370,N_14183,N_14062);
nor U14371 (N_14371,N_14234,N_14048);
nand U14372 (N_14372,N_14179,N_14105);
or U14373 (N_14373,N_14238,N_14104);
nand U14374 (N_14374,N_14196,N_14230);
xor U14375 (N_14375,N_14211,N_14085);
nor U14376 (N_14376,N_14025,N_14114);
nor U14377 (N_14377,N_14215,N_14050);
nand U14378 (N_14378,N_14240,N_14071);
nor U14379 (N_14379,N_14097,N_14035);
nor U14380 (N_14380,N_14001,N_14176);
nand U14381 (N_14381,N_14081,N_14181);
or U14382 (N_14382,N_14139,N_14194);
nand U14383 (N_14383,N_14194,N_14247);
nor U14384 (N_14384,N_14088,N_14211);
and U14385 (N_14385,N_14099,N_14080);
nor U14386 (N_14386,N_14024,N_14152);
xor U14387 (N_14387,N_14100,N_14006);
nand U14388 (N_14388,N_14106,N_14103);
xor U14389 (N_14389,N_14103,N_14240);
nor U14390 (N_14390,N_14186,N_14154);
and U14391 (N_14391,N_14011,N_14065);
nor U14392 (N_14392,N_14190,N_14227);
or U14393 (N_14393,N_14165,N_14193);
or U14394 (N_14394,N_14134,N_14145);
and U14395 (N_14395,N_14224,N_14067);
and U14396 (N_14396,N_14164,N_14180);
or U14397 (N_14397,N_14181,N_14064);
nor U14398 (N_14398,N_14045,N_14133);
nor U14399 (N_14399,N_14006,N_14001);
and U14400 (N_14400,N_14224,N_14037);
and U14401 (N_14401,N_14140,N_14009);
nand U14402 (N_14402,N_14029,N_14112);
xor U14403 (N_14403,N_14093,N_14038);
xor U14404 (N_14404,N_14153,N_14218);
and U14405 (N_14405,N_14246,N_14174);
and U14406 (N_14406,N_14034,N_14086);
nor U14407 (N_14407,N_14121,N_14008);
nand U14408 (N_14408,N_14041,N_14232);
nor U14409 (N_14409,N_14139,N_14192);
nand U14410 (N_14410,N_14051,N_14081);
nand U14411 (N_14411,N_14181,N_14089);
or U14412 (N_14412,N_14019,N_14134);
nand U14413 (N_14413,N_14035,N_14062);
or U14414 (N_14414,N_14158,N_14231);
nor U14415 (N_14415,N_14059,N_14247);
and U14416 (N_14416,N_14166,N_14227);
nand U14417 (N_14417,N_14152,N_14247);
xor U14418 (N_14418,N_14068,N_14066);
nor U14419 (N_14419,N_14107,N_14191);
xor U14420 (N_14420,N_14027,N_14030);
nand U14421 (N_14421,N_14004,N_14073);
and U14422 (N_14422,N_14176,N_14130);
nand U14423 (N_14423,N_14102,N_14188);
or U14424 (N_14424,N_14109,N_14083);
or U14425 (N_14425,N_14107,N_14124);
and U14426 (N_14426,N_14209,N_14027);
and U14427 (N_14427,N_14101,N_14155);
and U14428 (N_14428,N_14221,N_14158);
or U14429 (N_14429,N_14244,N_14119);
nand U14430 (N_14430,N_14009,N_14048);
nand U14431 (N_14431,N_14060,N_14208);
nand U14432 (N_14432,N_14152,N_14043);
xnor U14433 (N_14433,N_14056,N_14006);
nor U14434 (N_14434,N_14078,N_14145);
xor U14435 (N_14435,N_14054,N_14088);
or U14436 (N_14436,N_14218,N_14213);
nor U14437 (N_14437,N_14055,N_14048);
xnor U14438 (N_14438,N_14030,N_14209);
and U14439 (N_14439,N_14004,N_14076);
nand U14440 (N_14440,N_14210,N_14104);
and U14441 (N_14441,N_14240,N_14045);
and U14442 (N_14442,N_14249,N_14199);
nand U14443 (N_14443,N_14039,N_14205);
or U14444 (N_14444,N_14132,N_14174);
nor U14445 (N_14445,N_14131,N_14180);
xor U14446 (N_14446,N_14022,N_14066);
and U14447 (N_14447,N_14127,N_14178);
xor U14448 (N_14448,N_14089,N_14171);
nand U14449 (N_14449,N_14230,N_14180);
and U14450 (N_14450,N_14227,N_14085);
nor U14451 (N_14451,N_14044,N_14144);
or U14452 (N_14452,N_14100,N_14215);
and U14453 (N_14453,N_14188,N_14077);
or U14454 (N_14454,N_14027,N_14160);
nand U14455 (N_14455,N_14192,N_14025);
nand U14456 (N_14456,N_14013,N_14016);
nand U14457 (N_14457,N_14131,N_14019);
or U14458 (N_14458,N_14141,N_14020);
nand U14459 (N_14459,N_14184,N_14248);
nand U14460 (N_14460,N_14009,N_14206);
and U14461 (N_14461,N_14236,N_14039);
nand U14462 (N_14462,N_14118,N_14068);
nor U14463 (N_14463,N_14082,N_14052);
and U14464 (N_14464,N_14185,N_14007);
nand U14465 (N_14465,N_14054,N_14162);
and U14466 (N_14466,N_14037,N_14025);
or U14467 (N_14467,N_14156,N_14063);
nor U14468 (N_14468,N_14138,N_14036);
and U14469 (N_14469,N_14075,N_14182);
or U14470 (N_14470,N_14236,N_14201);
xnor U14471 (N_14471,N_14124,N_14038);
xor U14472 (N_14472,N_14217,N_14076);
nand U14473 (N_14473,N_14211,N_14097);
xnor U14474 (N_14474,N_14210,N_14163);
or U14475 (N_14475,N_14108,N_14245);
nand U14476 (N_14476,N_14248,N_14124);
or U14477 (N_14477,N_14156,N_14157);
or U14478 (N_14478,N_14145,N_14164);
or U14479 (N_14479,N_14135,N_14191);
nand U14480 (N_14480,N_14067,N_14061);
xor U14481 (N_14481,N_14188,N_14091);
or U14482 (N_14482,N_14247,N_14011);
and U14483 (N_14483,N_14147,N_14085);
nor U14484 (N_14484,N_14069,N_14053);
xor U14485 (N_14485,N_14218,N_14009);
or U14486 (N_14486,N_14230,N_14155);
and U14487 (N_14487,N_14060,N_14222);
and U14488 (N_14488,N_14045,N_14031);
nand U14489 (N_14489,N_14072,N_14080);
nor U14490 (N_14490,N_14164,N_14167);
nor U14491 (N_14491,N_14000,N_14023);
nand U14492 (N_14492,N_14141,N_14132);
and U14493 (N_14493,N_14068,N_14022);
or U14494 (N_14494,N_14038,N_14021);
nand U14495 (N_14495,N_14146,N_14139);
nor U14496 (N_14496,N_14158,N_14134);
or U14497 (N_14497,N_14169,N_14078);
nand U14498 (N_14498,N_14045,N_14156);
nor U14499 (N_14499,N_14066,N_14188);
nand U14500 (N_14500,N_14415,N_14416);
or U14501 (N_14501,N_14449,N_14399);
nor U14502 (N_14502,N_14436,N_14331);
or U14503 (N_14503,N_14406,N_14393);
and U14504 (N_14504,N_14255,N_14271);
nor U14505 (N_14505,N_14361,N_14412);
nand U14506 (N_14506,N_14464,N_14287);
nor U14507 (N_14507,N_14463,N_14297);
or U14508 (N_14508,N_14346,N_14370);
or U14509 (N_14509,N_14476,N_14429);
and U14510 (N_14510,N_14304,N_14282);
nor U14511 (N_14511,N_14278,N_14395);
or U14512 (N_14512,N_14337,N_14270);
nand U14513 (N_14513,N_14440,N_14432);
xnor U14514 (N_14514,N_14260,N_14422);
and U14515 (N_14515,N_14377,N_14456);
nor U14516 (N_14516,N_14286,N_14284);
xor U14517 (N_14517,N_14450,N_14333);
and U14518 (N_14518,N_14491,N_14258);
or U14519 (N_14519,N_14367,N_14434);
or U14520 (N_14520,N_14276,N_14389);
and U14521 (N_14521,N_14413,N_14482);
nand U14522 (N_14522,N_14397,N_14443);
or U14523 (N_14523,N_14497,N_14322);
and U14524 (N_14524,N_14380,N_14439);
and U14525 (N_14525,N_14310,N_14479);
nor U14526 (N_14526,N_14483,N_14314);
and U14527 (N_14527,N_14364,N_14332);
nor U14528 (N_14528,N_14461,N_14343);
nor U14529 (N_14529,N_14308,N_14360);
and U14530 (N_14530,N_14379,N_14452);
and U14531 (N_14531,N_14363,N_14475);
and U14532 (N_14532,N_14285,N_14474);
and U14533 (N_14533,N_14359,N_14495);
nor U14534 (N_14534,N_14394,N_14471);
nor U14535 (N_14535,N_14290,N_14273);
nor U14536 (N_14536,N_14431,N_14354);
or U14537 (N_14537,N_14374,N_14467);
nor U14538 (N_14538,N_14274,N_14468);
and U14539 (N_14539,N_14267,N_14460);
nor U14540 (N_14540,N_14300,N_14388);
nor U14541 (N_14541,N_14466,N_14329);
nand U14542 (N_14542,N_14369,N_14311);
or U14543 (N_14543,N_14384,N_14349);
nor U14544 (N_14544,N_14465,N_14455);
xnor U14545 (N_14545,N_14423,N_14317);
nor U14546 (N_14546,N_14433,N_14376);
nor U14547 (N_14547,N_14302,N_14498);
and U14548 (N_14548,N_14470,N_14437);
nor U14549 (N_14549,N_14404,N_14477);
nand U14550 (N_14550,N_14484,N_14387);
nor U14551 (N_14551,N_14252,N_14303);
nand U14552 (N_14552,N_14417,N_14487);
nor U14553 (N_14553,N_14294,N_14488);
xnor U14554 (N_14554,N_14435,N_14368);
nand U14555 (N_14555,N_14398,N_14373);
or U14556 (N_14556,N_14499,N_14313);
nor U14557 (N_14557,N_14338,N_14350);
nand U14558 (N_14558,N_14307,N_14353);
nand U14559 (N_14559,N_14279,N_14426);
and U14560 (N_14560,N_14462,N_14478);
or U14561 (N_14561,N_14288,N_14485);
xor U14562 (N_14562,N_14289,N_14262);
nand U14563 (N_14563,N_14472,N_14266);
and U14564 (N_14564,N_14486,N_14447);
nor U14565 (N_14565,N_14281,N_14489);
xor U14566 (N_14566,N_14493,N_14299);
nand U14567 (N_14567,N_14425,N_14321);
nand U14568 (N_14568,N_14257,N_14328);
or U14569 (N_14569,N_14371,N_14298);
and U14570 (N_14570,N_14254,N_14330);
or U14571 (N_14571,N_14480,N_14438);
or U14572 (N_14572,N_14420,N_14362);
or U14573 (N_14573,N_14419,N_14277);
nand U14574 (N_14574,N_14272,N_14347);
nand U14575 (N_14575,N_14342,N_14283);
nand U14576 (N_14576,N_14441,N_14268);
and U14577 (N_14577,N_14275,N_14336);
nand U14578 (N_14578,N_14265,N_14339);
nand U14579 (N_14579,N_14424,N_14319);
nor U14580 (N_14580,N_14459,N_14293);
and U14581 (N_14581,N_14357,N_14340);
and U14582 (N_14582,N_14358,N_14325);
or U14583 (N_14583,N_14291,N_14391);
or U14584 (N_14584,N_14344,N_14295);
and U14585 (N_14585,N_14372,N_14334);
nand U14586 (N_14586,N_14315,N_14356);
nand U14587 (N_14587,N_14296,N_14251);
nand U14588 (N_14588,N_14400,N_14263);
nor U14589 (N_14589,N_14401,N_14316);
or U14590 (N_14590,N_14309,N_14366);
or U14591 (N_14591,N_14445,N_14469);
and U14592 (N_14592,N_14341,N_14454);
and U14593 (N_14593,N_14355,N_14410);
nand U14594 (N_14594,N_14261,N_14259);
nand U14595 (N_14595,N_14408,N_14378);
and U14596 (N_14596,N_14327,N_14442);
or U14597 (N_14597,N_14335,N_14292);
nor U14598 (N_14598,N_14256,N_14326);
xor U14599 (N_14599,N_14418,N_14444);
or U14600 (N_14600,N_14407,N_14305);
or U14601 (N_14601,N_14481,N_14375);
and U14602 (N_14602,N_14494,N_14280);
and U14603 (N_14603,N_14414,N_14385);
and U14604 (N_14604,N_14386,N_14352);
nor U14605 (N_14605,N_14383,N_14411);
nand U14606 (N_14606,N_14451,N_14320);
or U14607 (N_14607,N_14306,N_14402);
or U14608 (N_14608,N_14382,N_14490);
nand U14609 (N_14609,N_14427,N_14448);
nor U14610 (N_14610,N_14409,N_14381);
nand U14611 (N_14611,N_14348,N_14473);
nand U14612 (N_14612,N_14324,N_14446);
and U14613 (N_14613,N_14492,N_14269);
nand U14614 (N_14614,N_14405,N_14421);
nand U14615 (N_14615,N_14250,N_14390);
and U14616 (N_14616,N_14396,N_14496);
nand U14617 (N_14617,N_14312,N_14253);
and U14618 (N_14618,N_14428,N_14403);
and U14619 (N_14619,N_14392,N_14458);
and U14620 (N_14620,N_14457,N_14323);
or U14621 (N_14621,N_14264,N_14345);
xnor U14622 (N_14622,N_14301,N_14318);
or U14623 (N_14623,N_14453,N_14430);
or U14624 (N_14624,N_14351,N_14365);
and U14625 (N_14625,N_14281,N_14448);
nor U14626 (N_14626,N_14273,N_14433);
or U14627 (N_14627,N_14298,N_14425);
or U14628 (N_14628,N_14494,N_14468);
and U14629 (N_14629,N_14434,N_14337);
nor U14630 (N_14630,N_14308,N_14407);
nand U14631 (N_14631,N_14356,N_14428);
and U14632 (N_14632,N_14356,N_14286);
or U14633 (N_14633,N_14393,N_14294);
or U14634 (N_14634,N_14497,N_14333);
nand U14635 (N_14635,N_14329,N_14367);
xnor U14636 (N_14636,N_14431,N_14366);
or U14637 (N_14637,N_14426,N_14351);
or U14638 (N_14638,N_14277,N_14326);
or U14639 (N_14639,N_14274,N_14353);
nand U14640 (N_14640,N_14497,N_14318);
or U14641 (N_14641,N_14263,N_14478);
nand U14642 (N_14642,N_14456,N_14277);
or U14643 (N_14643,N_14457,N_14308);
xor U14644 (N_14644,N_14344,N_14440);
or U14645 (N_14645,N_14292,N_14422);
nor U14646 (N_14646,N_14351,N_14282);
and U14647 (N_14647,N_14327,N_14305);
and U14648 (N_14648,N_14429,N_14457);
nand U14649 (N_14649,N_14386,N_14369);
and U14650 (N_14650,N_14458,N_14376);
nor U14651 (N_14651,N_14425,N_14452);
and U14652 (N_14652,N_14453,N_14412);
and U14653 (N_14653,N_14385,N_14450);
or U14654 (N_14654,N_14282,N_14349);
nor U14655 (N_14655,N_14464,N_14392);
nand U14656 (N_14656,N_14407,N_14454);
or U14657 (N_14657,N_14268,N_14472);
nand U14658 (N_14658,N_14350,N_14358);
and U14659 (N_14659,N_14316,N_14430);
and U14660 (N_14660,N_14418,N_14427);
nand U14661 (N_14661,N_14382,N_14453);
nand U14662 (N_14662,N_14257,N_14437);
or U14663 (N_14663,N_14404,N_14439);
nor U14664 (N_14664,N_14271,N_14387);
or U14665 (N_14665,N_14416,N_14287);
nor U14666 (N_14666,N_14483,N_14430);
or U14667 (N_14667,N_14325,N_14266);
nand U14668 (N_14668,N_14261,N_14423);
and U14669 (N_14669,N_14478,N_14313);
or U14670 (N_14670,N_14267,N_14272);
and U14671 (N_14671,N_14407,N_14351);
nand U14672 (N_14672,N_14382,N_14297);
xor U14673 (N_14673,N_14431,N_14443);
and U14674 (N_14674,N_14495,N_14405);
or U14675 (N_14675,N_14365,N_14305);
nor U14676 (N_14676,N_14423,N_14441);
nand U14677 (N_14677,N_14490,N_14283);
nand U14678 (N_14678,N_14450,N_14335);
or U14679 (N_14679,N_14357,N_14313);
and U14680 (N_14680,N_14390,N_14373);
and U14681 (N_14681,N_14466,N_14484);
or U14682 (N_14682,N_14405,N_14398);
nor U14683 (N_14683,N_14418,N_14278);
xnor U14684 (N_14684,N_14393,N_14261);
and U14685 (N_14685,N_14351,N_14451);
nand U14686 (N_14686,N_14328,N_14424);
nor U14687 (N_14687,N_14315,N_14300);
or U14688 (N_14688,N_14286,N_14459);
nand U14689 (N_14689,N_14288,N_14272);
and U14690 (N_14690,N_14489,N_14498);
nor U14691 (N_14691,N_14278,N_14388);
and U14692 (N_14692,N_14389,N_14316);
nand U14693 (N_14693,N_14254,N_14275);
and U14694 (N_14694,N_14263,N_14495);
or U14695 (N_14695,N_14305,N_14330);
nor U14696 (N_14696,N_14258,N_14257);
or U14697 (N_14697,N_14326,N_14323);
nand U14698 (N_14698,N_14488,N_14448);
xnor U14699 (N_14699,N_14387,N_14360);
or U14700 (N_14700,N_14409,N_14255);
or U14701 (N_14701,N_14472,N_14425);
or U14702 (N_14702,N_14399,N_14404);
nor U14703 (N_14703,N_14266,N_14282);
or U14704 (N_14704,N_14439,N_14386);
and U14705 (N_14705,N_14317,N_14369);
and U14706 (N_14706,N_14269,N_14473);
nand U14707 (N_14707,N_14408,N_14321);
xor U14708 (N_14708,N_14333,N_14417);
nand U14709 (N_14709,N_14269,N_14491);
xor U14710 (N_14710,N_14341,N_14299);
or U14711 (N_14711,N_14353,N_14269);
and U14712 (N_14712,N_14361,N_14384);
and U14713 (N_14713,N_14317,N_14269);
nand U14714 (N_14714,N_14390,N_14394);
xnor U14715 (N_14715,N_14363,N_14457);
nor U14716 (N_14716,N_14348,N_14354);
nor U14717 (N_14717,N_14287,N_14473);
nor U14718 (N_14718,N_14454,N_14370);
or U14719 (N_14719,N_14411,N_14404);
xnor U14720 (N_14720,N_14283,N_14312);
xnor U14721 (N_14721,N_14476,N_14403);
nand U14722 (N_14722,N_14478,N_14496);
nor U14723 (N_14723,N_14352,N_14380);
nor U14724 (N_14724,N_14494,N_14354);
nand U14725 (N_14725,N_14494,N_14317);
and U14726 (N_14726,N_14325,N_14368);
xor U14727 (N_14727,N_14261,N_14446);
and U14728 (N_14728,N_14395,N_14309);
or U14729 (N_14729,N_14324,N_14376);
nand U14730 (N_14730,N_14384,N_14418);
xor U14731 (N_14731,N_14396,N_14367);
or U14732 (N_14732,N_14459,N_14328);
nor U14733 (N_14733,N_14481,N_14294);
nor U14734 (N_14734,N_14405,N_14377);
or U14735 (N_14735,N_14375,N_14338);
and U14736 (N_14736,N_14279,N_14414);
and U14737 (N_14737,N_14473,N_14311);
and U14738 (N_14738,N_14427,N_14344);
xor U14739 (N_14739,N_14289,N_14427);
xnor U14740 (N_14740,N_14440,N_14381);
and U14741 (N_14741,N_14272,N_14474);
and U14742 (N_14742,N_14339,N_14341);
or U14743 (N_14743,N_14273,N_14398);
nor U14744 (N_14744,N_14306,N_14291);
and U14745 (N_14745,N_14320,N_14294);
nand U14746 (N_14746,N_14266,N_14369);
nand U14747 (N_14747,N_14447,N_14377);
and U14748 (N_14748,N_14477,N_14385);
nand U14749 (N_14749,N_14295,N_14363);
and U14750 (N_14750,N_14585,N_14631);
xnor U14751 (N_14751,N_14726,N_14649);
or U14752 (N_14752,N_14692,N_14674);
or U14753 (N_14753,N_14538,N_14640);
xnor U14754 (N_14754,N_14673,N_14688);
or U14755 (N_14755,N_14614,N_14623);
nand U14756 (N_14756,N_14700,N_14633);
and U14757 (N_14757,N_14509,N_14703);
and U14758 (N_14758,N_14643,N_14507);
and U14759 (N_14759,N_14510,N_14530);
or U14760 (N_14760,N_14722,N_14542);
nand U14761 (N_14761,N_14734,N_14537);
nand U14762 (N_14762,N_14705,N_14588);
or U14763 (N_14763,N_14744,N_14682);
xor U14764 (N_14764,N_14604,N_14583);
xnor U14765 (N_14765,N_14712,N_14600);
and U14766 (N_14766,N_14672,N_14586);
or U14767 (N_14767,N_14724,N_14638);
or U14768 (N_14768,N_14644,N_14717);
nor U14769 (N_14769,N_14540,N_14581);
or U14770 (N_14770,N_14701,N_14660);
nand U14771 (N_14771,N_14580,N_14691);
nor U14772 (N_14772,N_14518,N_14582);
xor U14773 (N_14773,N_14661,N_14730);
and U14774 (N_14774,N_14523,N_14664);
nor U14775 (N_14775,N_14541,N_14591);
and U14776 (N_14776,N_14655,N_14652);
nand U14777 (N_14777,N_14728,N_14749);
nand U14778 (N_14778,N_14519,N_14587);
nor U14779 (N_14779,N_14677,N_14566);
or U14780 (N_14780,N_14647,N_14666);
and U14781 (N_14781,N_14571,N_14511);
or U14782 (N_14782,N_14513,N_14517);
xor U14783 (N_14783,N_14683,N_14619);
or U14784 (N_14784,N_14748,N_14743);
nor U14785 (N_14785,N_14626,N_14694);
or U14786 (N_14786,N_14628,N_14556);
or U14787 (N_14787,N_14684,N_14596);
nand U14788 (N_14788,N_14563,N_14565);
or U14789 (N_14789,N_14716,N_14708);
or U14790 (N_14790,N_14551,N_14552);
nor U14791 (N_14791,N_14697,N_14501);
and U14792 (N_14792,N_14569,N_14528);
or U14793 (N_14793,N_14693,N_14606);
and U14794 (N_14794,N_14520,N_14531);
nor U14795 (N_14795,N_14555,N_14742);
nand U14796 (N_14796,N_14747,N_14533);
and U14797 (N_14797,N_14745,N_14512);
nor U14798 (N_14798,N_14639,N_14738);
or U14799 (N_14799,N_14746,N_14667);
or U14800 (N_14800,N_14613,N_14572);
nor U14801 (N_14801,N_14645,N_14713);
or U14802 (N_14802,N_14579,N_14627);
or U14803 (N_14803,N_14608,N_14634);
nand U14804 (N_14804,N_14632,N_14729);
and U14805 (N_14805,N_14637,N_14603);
nand U14806 (N_14806,N_14567,N_14611);
nor U14807 (N_14807,N_14594,N_14609);
xnor U14808 (N_14808,N_14592,N_14553);
xor U14809 (N_14809,N_14521,N_14699);
xor U14810 (N_14810,N_14605,N_14737);
nor U14811 (N_14811,N_14695,N_14725);
and U14812 (N_14812,N_14736,N_14656);
xor U14813 (N_14813,N_14589,N_14678);
or U14814 (N_14814,N_14715,N_14545);
or U14815 (N_14815,N_14557,N_14687);
or U14816 (N_14816,N_14524,N_14577);
or U14817 (N_14817,N_14584,N_14597);
nand U14818 (N_14818,N_14731,N_14680);
xnor U14819 (N_14819,N_14503,N_14668);
or U14820 (N_14820,N_14617,N_14689);
or U14821 (N_14821,N_14598,N_14685);
xor U14822 (N_14822,N_14669,N_14721);
or U14823 (N_14823,N_14739,N_14532);
nand U14824 (N_14824,N_14535,N_14612);
nor U14825 (N_14825,N_14522,N_14505);
nand U14826 (N_14826,N_14706,N_14558);
or U14827 (N_14827,N_14602,N_14711);
nand U14828 (N_14828,N_14618,N_14727);
and U14829 (N_14829,N_14709,N_14679);
nand U14830 (N_14830,N_14681,N_14526);
xnor U14831 (N_14831,N_14576,N_14620);
and U14832 (N_14832,N_14593,N_14615);
nor U14833 (N_14833,N_14574,N_14527);
nor U14834 (N_14834,N_14675,N_14502);
and U14835 (N_14835,N_14696,N_14568);
nand U14836 (N_14836,N_14686,N_14559);
or U14837 (N_14837,N_14657,N_14590);
xor U14838 (N_14838,N_14514,N_14653);
nor U14839 (N_14839,N_14740,N_14543);
nand U14840 (N_14840,N_14698,N_14508);
or U14841 (N_14841,N_14500,N_14610);
or U14842 (N_14842,N_14525,N_14515);
and U14843 (N_14843,N_14710,N_14735);
nor U14844 (N_14844,N_14646,N_14648);
or U14845 (N_14845,N_14671,N_14570);
nand U14846 (N_14846,N_14539,N_14719);
nor U14847 (N_14847,N_14536,N_14595);
and U14848 (N_14848,N_14670,N_14658);
and U14849 (N_14849,N_14629,N_14676);
nor U14850 (N_14850,N_14650,N_14718);
and U14851 (N_14851,N_14662,N_14732);
nand U14852 (N_14852,N_14636,N_14704);
nor U14853 (N_14853,N_14506,N_14573);
or U14854 (N_14854,N_14654,N_14578);
and U14855 (N_14855,N_14642,N_14575);
or U14856 (N_14856,N_14548,N_14562);
nand U14857 (N_14857,N_14659,N_14564);
and U14858 (N_14858,N_14741,N_14547);
nor U14859 (N_14859,N_14663,N_14720);
nand U14860 (N_14860,N_14630,N_14607);
nand U14861 (N_14861,N_14601,N_14714);
nand U14862 (N_14862,N_14560,N_14561);
nor U14863 (N_14863,N_14622,N_14625);
or U14864 (N_14864,N_14616,N_14504);
and U14865 (N_14865,N_14733,N_14534);
nor U14866 (N_14866,N_14550,N_14651);
and U14867 (N_14867,N_14723,N_14641);
nor U14868 (N_14868,N_14544,N_14516);
and U14869 (N_14869,N_14554,N_14624);
nand U14870 (N_14870,N_14665,N_14702);
and U14871 (N_14871,N_14599,N_14635);
nand U14872 (N_14872,N_14621,N_14529);
nor U14873 (N_14873,N_14707,N_14690);
nor U14874 (N_14874,N_14549,N_14546);
or U14875 (N_14875,N_14744,N_14533);
xnor U14876 (N_14876,N_14594,N_14509);
and U14877 (N_14877,N_14685,N_14595);
and U14878 (N_14878,N_14671,N_14549);
nand U14879 (N_14879,N_14528,N_14640);
nand U14880 (N_14880,N_14513,N_14680);
and U14881 (N_14881,N_14570,N_14596);
and U14882 (N_14882,N_14694,N_14590);
nand U14883 (N_14883,N_14626,N_14585);
or U14884 (N_14884,N_14680,N_14643);
or U14885 (N_14885,N_14554,N_14642);
xnor U14886 (N_14886,N_14692,N_14654);
and U14887 (N_14887,N_14559,N_14595);
and U14888 (N_14888,N_14622,N_14699);
nor U14889 (N_14889,N_14526,N_14699);
and U14890 (N_14890,N_14654,N_14565);
and U14891 (N_14891,N_14748,N_14599);
and U14892 (N_14892,N_14731,N_14538);
nor U14893 (N_14893,N_14652,N_14699);
nor U14894 (N_14894,N_14560,N_14634);
and U14895 (N_14895,N_14605,N_14555);
nor U14896 (N_14896,N_14501,N_14706);
nand U14897 (N_14897,N_14580,N_14551);
and U14898 (N_14898,N_14648,N_14569);
nor U14899 (N_14899,N_14587,N_14535);
xnor U14900 (N_14900,N_14634,N_14621);
and U14901 (N_14901,N_14731,N_14628);
nor U14902 (N_14902,N_14727,N_14695);
and U14903 (N_14903,N_14562,N_14524);
and U14904 (N_14904,N_14628,N_14616);
and U14905 (N_14905,N_14674,N_14615);
xor U14906 (N_14906,N_14624,N_14571);
or U14907 (N_14907,N_14655,N_14527);
nand U14908 (N_14908,N_14581,N_14720);
nand U14909 (N_14909,N_14706,N_14611);
and U14910 (N_14910,N_14741,N_14590);
or U14911 (N_14911,N_14657,N_14529);
nand U14912 (N_14912,N_14651,N_14510);
nor U14913 (N_14913,N_14720,N_14729);
xnor U14914 (N_14914,N_14525,N_14744);
and U14915 (N_14915,N_14593,N_14656);
nand U14916 (N_14916,N_14621,N_14571);
nor U14917 (N_14917,N_14614,N_14709);
xor U14918 (N_14918,N_14736,N_14535);
nor U14919 (N_14919,N_14554,N_14596);
or U14920 (N_14920,N_14662,N_14557);
nand U14921 (N_14921,N_14603,N_14504);
or U14922 (N_14922,N_14548,N_14695);
or U14923 (N_14923,N_14548,N_14541);
or U14924 (N_14924,N_14672,N_14528);
and U14925 (N_14925,N_14541,N_14526);
xnor U14926 (N_14926,N_14539,N_14599);
nor U14927 (N_14927,N_14696,N_14743);
or U14928 (N_14928,N_14684,N_14648);
xor U14929 (N_14929,N_14551,N_14728);
or U14930 (N_14930,N_14562,N_14552);
nand U14931 (N_14931,N_14552,N_14535);
nor U14932 (N_14932,N_14673,N_14576);
and U14933 (N_14933,N_14620,N_14677);
xnor U14934 (N_14934,N_14554,N_14672);
nand U14935 (N_14935,N_14734,N_14619);
nor U14936 (N_14936,N_14522,N_14603);
nand U14937 (N_14937,N_14690,N_14621);
and U14938 (N_14938,N_14617,N_14712);
nand U14939 (N_14939,N_14687,N_14527);
or U14940 (N_14940,N_14554,N_14592);
nand U14941 (N_14941,N_14532,N_14703);
nor U14942 (N_14942,N_14560,N_14715);
nor U14943 (N_14943,N_14513,N_14735);
nor U14944 (N_14944,N_14528,N_14746);
nand U14945 (N_14945,N_14630,N_14726);
nor U14946 (N_14946,N_14625,N_14558);
nand U14947 (N_14947,N_14739,N_14561);
nor U14948 (N_14948,N_14535,N_14550);
nor U14949 (N_14949,N_14676,N_14655);
and U14950 (N_14950,N_14619,N_14685);
nand U14951 (N_14951,N_14576,N_14540);
or U14952 (N_14952,N_14673,N_14635);
and U14953 (N_14953,N_14541,N_14525);
nand U14954 (N_14954,N_14697,N_14603);
nor U14955 (N_14955,N_14715,N_14543);
nor U14956 (N_14956,N_14749,N_14710);
and U14957 (N_14957,N_14675,N_14727);
nor U14958 (N_14958,N_14646,N_14578);
nor U14959 (N_14959,N_14692,N_14737);
nand U14960 (N_14960,N_14700,N_14732);
nor U14961 (N_14961,N_14609,N_14591);
or U14962 (N_14962,N_14727,N_14728);
or U14963 (N_14963,N_14614,N_14619);
or U14964 (N_14964,N_14728,N_14545);
and U14965 (N_14965,N_14698,N_14594);
and U14966 (N_14966,N_14747,N_14716);
nand U14967 (N_14967,N_14544,N_14684);
nor U14968 (N_14968,N_14688,N_14680);
nor U14969 (N_14969,N_14629,N_14624);
xor U14970 (N_14970,N_14746,N_14551);
nor U14971 (N_14971,N_14674,N_14542);
nand U14972 (N_14972,N_14538,N_14744);
and U14973 (N_14973,N_14671,N_14709);
nand U14974 (N_14974,N_14675,N_14668);
nand U14975 (N_14975,N_14736,N_14667);
nand U14976 (N_14976,N_14514,N_14666);
xnor U14977 (N_14977,N_14722,N_14610);
and U14978 (N_14978,N_14701,N_14546);
nor U14979 (N_14979,N_14516,N_14650);
or U14980 (N_14980,N_14567,N_14664);
and U14981 (N_14981,N_14518,N_14666);
and U14982 (N_14982,N_14634,N_14702);
and U14983 (N_14983,N_14649,N_14704);
or U14984 (N_14984,N_14713,N_14571);
or U14985 (N_14985,N_14567,N_14617);
nand U14986 (N_14986,N_14635,N_14748);
xor U14987 (N_14987,N_14691,N_14609);
or U14988 (N_14988,N_14699,N_14597);
and U14989 (N_14989,N_14693,N_14580);
nor U14990 (N_14990,N_14567,N_14686);
and U14991 (N_14991,N_14540,N_14538);
or U14992 (N_14992,N_14685,N_14558);
or U14993 (N_14993,N_14501,N_14728);
and U14994 (N_14994,N_14648,N_14736);
nor U14995 (N_14995,N_14613,N_14657);
and U14996 (N_14996,N_14517,N_14748);
and U14997 (N_14997,N_14609,N_14647);
nor U14998 (N_14998,N_14689,N_14546);
nor U14999 (N_14999,N_14701,N_14667);
or U15000 (N_15000,N_14966,N_14795);
nand U15001 (N_15001,N_14761,N_14931);
or U15002 (N_15002,N_14834,N_14967);
xnor U15003 (N_15003,N_14932,N_14804);
nand U15004 (N_15004,N_14753,N_14918);
nor U15005 (N_15005,N_14896,N_14789);
nor U15006 (N_15006,N_14828,N_14872);
nand U15007 (N_15007,N_14874,N_14940);
nand U15008 (N_15008,N_14776,N_14861);
and U15009 (N_15009,N_14801,N_14954);
and U15010 (N_15010,N_14963,N_14751);
nor U15011 (N_15011,N_14847,N_14781);
and U15012 (N_15012,N_14826,N_14916);
nand U15013 (N_15013,N_14886,N_14901);
nor U15014 (N_15014,N_14927,N_14929);
nand U15015 (N_15015,N_14843,N_14914);
nor U15016 (N_15016,N_14868,N_14875);
nor U15017 (N_15017,N_14835,N_14906);
nand U15018 (N_15018,N_14923,N_14971);
nor U15019 (N_15019,N_14904,N_14827);
and U15020 (N_15020,N_14850,N_14911);
nor U15021 (N_15021,N_14957,N_14993);
nor U15022 (N_15022,N_14976,N_14894);
or U15023 (N_15023,N_14972,N_14889);
xor U15024 (N_15024,N_14917,N_14752);
or U15025 (N_15025,N_14756,N_14785);
nand U15026 (N_15026,N_14829,N_14989);
nand U15027 (N_15027,N_14974,N_14900);
xnor U15028 (N_15028,N_14837,N_14962);
or U15029 (N_15029,N_14750,N_14771);
nor U15030 (N_15030,N_14965,N_14867);
nand U15031 (N_15031,N_14824,N_14964);
xnor U15032 (N_15032,N_14767,N_14882);
xor U15033 (N_15033,N_14952,N_14769);
and U15034 (N_15034,N_14864,N_14758);
nor U15035 (N_15035,N_14833,N_14869);
and U15036 (N_15036,N_14848,N_14890);
or U15037 (N_15037,N_14854,N_14786);
nor U15038 (N_15038,N_14772,N_14936);
nor U15039 (N_15039,N_14788,N_14798);
xnor U15040 (N_15040,N_14888,N_14812);
nand U15041 (N_15041,N_14773,N_14770);
and U15042 (N_15042,N_14898,N_14779);
nand U15043 (N_15043,N_14836,N_14921);
nor U15044 (N_15044,N_14947,N_14846);
nor U15045 (N_15045,N_14938,N_14809);
or U15046 (N_15046,N_14897,N_14825);
and U15047 (N_15047,N_14803,N_14873);
nor U15048 (N_15048,N_14978,N_14794);
or U15049 (N_15049,N_14999,N_14941);
nor U15050 (N_15050,N_14881,N_14939);
nor U15051 (N_15051,N_14946,N_14983);
or U15052 (N_15052,N_14830,N_14977);
and U15053 (N_15053,N_14760,N_14992);
and U15054 (N_15054,N_14968,N_14956);
or U15055 (N_15055,N_14959,N_14997);
and U15056 (N_15056,N_14996,N_14823);
xor U15057 (N_15057,N_14984,N_14793);
nand U15058 (N_15058,N_14818,N_14925);
nor U15059 (N_15059,N_14919,N_14821);
nand U15060 (N_15060,N_14950,N_14951);
nand U15061 (N_15061,N_14844,N_14775);
and U15062 (N_15062,N_14883,N_14885);
and U15063 (N_15063,N_14949,N_14852);
xnor U15064 (N_15064,N_14870,N_14855);
and U15065 (N_15065,N_14928,N_14980);
nor U15066 (N_15066,N_14831,N_14865);
and U15067 (N_15067,N_14853,N_14995);
nor U15068 (N_15068,N_14849,N_14907);
or U15069 (N_15069,N_14944,N_14930);
nand U15070 (N_15070,N_14948,N_14895);
xor U15071 (N_15071,N_14819,N_14981);
nand U15072 (N_15072,N_14856,N_14892);
or U15073 (N_15073,N_14808,N_14934);
nor U15074 (N_15074,N_14859,N_14796);
nand U15075 (N_15075,N_14822,N_14990);
and U15076 (N_15076,N_14858,N_14813);
and U15077 (N_15077,N_14862,N_14961);
xor U15078 (N_15078,N_14778,N_14902);
or U15079 (N_15079,N_14797,N_14942);
nor U15080 (N_15080,N_14887,N_14899);
or U15081 (N_15081,N_14879,N_14933);
or U15082 (N_15082,N_14987,N_14790);
or U15083 (N_15083,N_14816,N_14857);
or U15084 (N_15084,N_14945,N_14991);
nor U15085 (N_15085,N_14800,N_14876);
or U15086 (N_15086,N_14943,N_14810);
and U15087 (N_15087,N_14994,N_14937);
or U15088 (N_15088,N_14893,N_14908);
or U15089 (N_15089,N_14764,N_14910);
and U15090 (N_15090,N_14979,N_14973);
or U15091 (N_15091,N_14969,N_14909);
and U15092 (N_15092,N_14985,N_14960);
xor U15093 (N_15093,N_14860,N_14988);
nand U15094 (N_15094,N_14754,N_14975);
or U15095 (N_15095,N_14851,N_14762);
nand U15096 (N_15096,N_14784,N_14866);
and U15097 (N_15097,N_14871,N_14799);
nor U15098 (N_15098,N_14998,N_14806);
or U15099 (N_15099,N_14926,N_14884);
nor U15100 (N_15100,N_14805,N_14839);
or U15101 (N_15101,N_14755,N_14915);
and U15102 (N_15102,N_14841,N_14891);
nand U15103 (N_15103,N_14768,N_14807);
nand U15104 (N_15104,N_14955,N_14791);
xnor U15105 (N_15105,N_14912,N_14958);
or U15106 (N_15106,N_14863,N_14905);
xnor U15107 (N_15107,N_14832,N_14953);
nor U15108 (N_15108,N_14815,N_14986);
nand U15109 (N_15109,N_14903,N_14935);
nand U15110 (N_15110,N_14757,N_14766);
nor U15111 (N_15111,N_14842,N_14838);
xnor U15112 (N_15112,N_14782,N_14763);
or U15113 (N_15113,N_14814,N_14802);
nand U15114 (N_15114,N_14774,N_14878);
and U15115 (N_15115,N_14982,N_14924);
and U15116 (N_15116,N_14780,N_14845);
nor U15117 (N_15117,N_14765,N_14920);
nor U15118 (N_15118,N_14787,N_14820);
and U15119 (N_15119,N_14840,N_14913);
and U15120 (N_15120,N_14922,N_14817);
xnor U15121 (N_15121,N_14759,N_14811);
nor U15122 (N_15122,N_14880,N_14777);
nand U15123 (N_15123,N_14792,N_14783);
nand U15124 (N_15124,N_14877,N_14970);
nand U15125 (N_15125,N_14941,N_14860);
nor U15126 (N_15126,N_14932,N_14812);
nor U15127 (N_15127,N_14757,N_14962);
nor U15128 (N_15128,N_14878,N_14913);
and U15129 (N_15129,N_14966,N_14963);
or U15130 (N_15130,N_14788,N_14838);
nand U15131 (N_15131,N_14767,N_14885);
or U15132 (N_15132,N_14770,N_14829);
nor U15133 (N_15133,N_14874,N_14965);
and U15134 (N_15134,N_14964,N_14770);
nor U15135 (N_15135,N_14838,N_14850);
nor U15136 (N_15136,N_14763,N_14847);
or U15137 (N_15137,N_14982,N_14974);
and U15138 (N_15138,N_14780,N_14952);
nand U15139 (N_15139,N_14935,N_14808);
nor U15140 (N_15140,N_14776,N_14804);
nand U15141 (N_15141,N_14924,N_14826);
nand U15142 (N_15142,N_14916,N_14806);
or U15143 (N_15143,N_14787,N_14957);
xnor U15144 (N_15144,N_14830,N_14887);
or U15145 (N_15145,N_14931,N_14892);
xor U15146 (N_15146,N_14909,N_14953);
nor U15147 (N_15147,N_14806,N_14953);
nand U15148 (N_15148,N_14992,N_14754);
nand U15149 (N_15149,N_14807,N_14863);
and U15150 (N_15150,N_14972,N_14847);
nor U15151 (N_15151,N_14896,N_14954);
xor U15152 (N_15152,N_14823,N_14817);
nor U15153 (N_15153,N_14876,N_14878);
nor U15154 (N_15154,N_14947,N_14870);
and U15155 (N_15155,N_14980,N_14937);
or U15156 (N_15156,N_14835,N_14757);
nor U15157 (N_15157,N_14904,N_14976);
xnor U15158 (N_15158,N_14956,N_14907);
nor U15159 (N_15159,N_14961,N_14965);
nand U15160 (N_15160,N_14783,N_14776);
nor U15161 (N_15161,N_14906,N_14787);
xor U15162 (N_15162,N_14965,N_14889);
or U15163 (N_15163,N_14778,N_14912);
nor U15164 (N_15164,N_14881,N_14953);
nor U15165 (N_15165,N_14997,N_14822);
and U15166 (N_15166,N_14780,N_14784);
nand U15167 (N_15167,N_14883,N_14850);
xnor U15168 (N_15168,N_14951,N_14892);
nand U15169 (N_15169,N_14998,N_14917);
or U15170 (N_15170,N_14919,N_14850);
and U15171 (N_15171,N_14827,N_14897);
or U15172 (N_15172,N_14760,N_14775);
and U15173 (N_15173,N_14979,N_14778);
or U15174 (N_15174,N_14843,N_14989);
and U15175 (N_15175,N_14968,N_14864);
nand U15176 (N_15176,N_14972,N_14887);
nand U15177 (N_15177,N_14956,N_14878);
nor U15178 (N_15178,N_14886,N_14995);
nor U15179 (N_15179,N_14922,N_14928);
or U15180 (N_15180,N_14871,N_14813);
or U15181 (N_15181,N_14994,N_14815);
and U15182 (N_15182,N_14937,N_14960);
nand U15183 (N_15183,N_14996,N_14855);
and U15184 (N_15184,N_14899,N_14750);
nor U15185 (N_15185,N_14785,N_14767);
and U15186 (N_15186,N_14918,N_14967);
and U15187 (N_15187,N_14837,N_14866);
and U15188 (N_15188,N_14960,N_14842);
or U15189 (N_15189,N_14780,N_14987);
xor U15190 (N_15190,N_14825,N_14785);
nand U15191 (N_15191,N_14886,N_14963);
and U15192 (N_15192,N_14867,N_14960);
and U15193 (N_15193,N_14974,N_14873);
and U15194 (N_15194,N_14868,N_14855);
and U15195 (N_15195,N_14768,N_14879);
nor U15196 (N_15196,N_14890,N_14774);
nor U15197 (N_15197,N_14938,N_14899);
nor U15198 (N_15198,N_14840,N_14771);
nor U15199 (N_15199,N_14917,N_14757);
and U15200 (N_15200,N_14987,N_14852);
nor U15201 (N_15201,N_14819,N_14897);
nand U15202 (N_15202,N_14798,N_14911);
and U15203 (N_15203,N_14934,N_14759);
xnor U15204 (N_15204,N_14909,N_14973);
or U15205 (N_15205,N_14780,N_14800);
nand U15206 (N_15206,N_14910,N_14877);
or U15207 (N_15207,N_14779,N_14946);
nand U15208 (N_15208,N_14934,N_14864);
and U15209 (N_15209,N_14841,N_14884);
nor U15210 (N_15210,N_14900,N_14841);
and U15211 (N_15211,N_14920,N_14948);
and U15212 (N_15212,N_14971,N_14962);
and U15213 (N_15213,N_14767,N_14847);
or U15214 (N_15214,N_14789,N_14930);
or U15215 (N_15215,N_14948,N_14916);
nor U15216 (N_15216,N_14982,N_14847);
and U15217 (N_15217,N_14864,N_14973);
or U15218 (N_15218,N_14753,N_14982);
nand U15219 (N_15219,N_14758,N_14949);
and U15220 (N_15220,N_14866,N_14840);
nor U15221 (N_15221,N_14869,N_14935);
nor U15222 (N_15222,N_14846,N_14798);
xor U15223 (N_15223,N_14750,N_14765);
or U15224 (N_15224,N_14970,N_14793);
and U15225 (N_15225,N_14956,N_14872);
nor U15226 (N_15226,N_14986,N_14936);
nor U15227 (N_15227,N_14977,N_14930);
and U15228 (N_15228,N_14904,N_14886);
xnor U15229 (N_15229,N_14762,N_14870);
and U15230 (N_15230,N_14872,N_14949);
and U15231 (N_15231,N_14763,N_14915);
nor U15232 (N_15232,N_14833,N_14942);
and U15233 (N_15233,N_14755,N_14903);
and U15234 (N_15234,N_14752,N_14847);
or U15235 (N_15235,N_14988,N_14908);
nor U15236 (N_15236,N_14988,N_14750);
nand U15237 (N_15237,N_14898,N_14881);
and U15238 (N_15238,N_14952,N_14781);
and U15239 (N_15239,N_14818,N_14804);
nand U15240 (N_15240,N_14980,N_14950);
nor U15241 (N_15241,N_14757,N_14951);
xnor U15242 (N_15242,N_14753,N_14764);
or U15243 (N_15243,N_14843,N_14826);
or U15244 (N_15244,N_14815,N_14857);
and U15245 (N_15245,N_14803,N_14880);
or U15246 (N_15246,N_14896,N_14860);
nand U15247 (N_15247,N_14819,N_14941);
nor U15248 (N_15248,N_14816,N_14815);
or U15249 (N_15249,N_14971,N_14952);
nand U15250 (N_15250,N_15202,N_15102);
and U15251 (N_15251,N_15244,N_15094);
or U15252 (N_15252,N_15151,N_15084);
nor U15253 (N_15253,N_15081,N_15025);
nand U15254 (N_15254,N_15049,N_15132);
and U15255 (N_15255,N_15221,N_15188);
or U15256 (N_15256,N_15237,N_15184);
or U15257 (N_15257,N_15074,N_15182);
and U15258 (N_15258,N_15110,N_15013);
nand U15259 (N_15259,N_15108,N_15091);
nor U15260 (N_15260,N_15011,N_15208);
or U15261 (N_15261,N_15076,N_15080);
or U15262 (N_15262,N_15028,N_15157);
and U15263 (N_15263,N_15001,N_15064);
and U15264 (N_15264,N_15130,N_15048);
nand U15265 (N_15265,N_15008,N_15159);
and U15266 (N_15266,N_15134,N_15021);
nand U15267 (N_15267,N_15045,N_15195);
or U15268 (N_15268,N_15220,N_15210);
or U15269 (N_15269,N_15227,N_15065);
and U15270 (N_15270,N_15191,N_15027);
nand U15271 (N_15271,N_15103,N_15003);
nand U15272 (N_15272,N_15068,N_15038);
nand U15273 (N_15273,N_15169,N_15053);
or U15274 (N_15274,N_15040,N_15183);
and U15275 (N_15275,N_15109,N_15181);
or U15276 (N_15276,N_15017,N_15160);
nor U15277 (N_15277,N_15128,N_15047);
or U15278 (N_15278,N_15225,N_15033);
and U15279 (N_15279,N_15034,N_15111);
and U15280 (N_15280,N_15187,N_15089);
nor U15281 (N_15281,N_15217,N_15120);
or U15282 (N_15282,N_15072,N_15239);
nand U15283 (N_15283,N_15155,N_15143);
nor U15284 (N_15284,N_15205,N_15164);
nor U15285 (N_15285,N_15119,N_15235);
or U15286 (N_15286,N_15026,N_15144);
or U15287 (N_15287,N_15173,N_15057);
and U15288 (N_15288,N_15106,N_15179);
and U15289 (N_15289,N_15212,N_15036);
nand U15290 (N_15290,N_15168,N_15185);
nand U15291 (N_15291,N_15096,N_15060);
nand U15292 (N_15292,N_15046,N_15122);
or U15293 (N_15293,N_15054,N_15056);
or U15294 (N_15294,N_15207,N_15206);
xnor U15295 (N_15295,N_15009,N_15166);
and U15296 (N_15296,N_15136,N_15113);
or U15297 (N_15297,N_15148,N_15088);
nand U15298 (N_15298,N_15032,N_15000);
and U15299 (N_15299,N_15229,N_15236);
nand U15300 (N_15300,N_15020,N_15247);
nor U15301 (N_15301,N_15012,N_15135);
nand U15302 (N_15302,N_15002,N_15117);
and U15303 (N_15303,N_15177,N_15006);
xor U15304 (N_15304,N_15125,N_15077);
nor U15305 (N_15305,N_15243,N_15142);
and U15306 (N_15306,N_15153,N_15055);
nand U15307 (N_15307,N_15004,N_15052);
nor U15308 (N_15308,N_15198,N_15190);
nor U15309 (N_15309,N_15051,N_15116);
or U15310 (N_15310,N_15124,N_15101);
nor U15311 (N_15311,N_15174,N_15231);
xor U15312 (N_15312,N_15010,N_15211);
nand U15313 (N_15313,N_15133,N_15029);
or U15314 (N_15314,N_15005,N_15215);
nor U15315 (N_15315,N_15121,N_15093);
nor U15316 (N_15316,N_15024,N_15234);
nand U15317 (N_15317,N_15186,N_15150);
and U15318 (N_15318,N_15097,N_15178);
and U15319 (N_15319,N_15085,N_15209);
or U15320 (N_15320,N_15100,N_15249);
nand U15321 (N_15321,N_15015,N_15203);
nand U15322 (N_15322,N_15149,N_15140);
and U15323 (N_15323,N_15030,N_15146);
nor U15324 (N_15324,N_15167,N_15196);
nand U15325 (N_15325,N_15066,N_15067);
or U15326 (N_15326,N_15241,N_15044);
nor U15327 (N_15327,N_15043,N_15158);
nand U15328 (N_15328,N_15083,N_15233);
and U15329 (N_15329,N_15194,N_15090);
and U15330 (N_15330,N_15213,N_15246);
nor U15331 (N_15331,N_15214,N_15063);
or U15332 (N_15332,N_15138,N_15131);
nand U15333 (N_15333,N_15087,N_15098);
nand U15334 (N_15334,N_15023,N_15050);
and U15335 (N_15335,N_15242,N_15156);
nand U15336 (N_15336,N_15031,N_15176);
nand U15337 (N_15337,N_15218,N_15129);
or U15338 (N_15338,N_15042,N_15059);
nor U15339 (N_15339,N_15163,N_15018);
nand U15340 (N_15340,N_15114,N_15171);
and U15341 (N_15341,N_15022,N_15082);
nor U15342 (N_15342,N_15228,N_15137);
nand U15343 (N_15343,N_15180,N_15092);
or U15344 (N_15344,N_15104,N_15014);
nor U15345 (N_15345,N_15071,N_15039);
xor U15346 (N_15346,N_15172,N_15248);
nor U15347 (N_15347,N_15118,N_15161);
nor U15348 (N_15348,N_15070,N_15238);
or U15349 (N_15349,N_15019,N_15086);
nor U15350 (N_15350,N_15170,N_15069);
nor U15351 (N_15351,N_15061,N_15219);
and U15352 (N_15352,N_15105,N_15078);
nor U15353 (N_15353,N_15079,N_15232);
nand U15354 (N_15354,N_15007,N_15037);
nand U15355 (N_15355,N_15123,N_15035);
nor U15356 (N_15356,N_15062,N_15197);
and U15357 (N_15357,N_15165,N_15095);
nand U15358 (N_15358,N_15226,N_15073);
nor U15359 (N_15359,N_15189,N_15200);
or U15360 (N_15360,N_15192,N_15107);
nor U15361 (N_15361,N_15041,N_15141);
nor U15362 (N_15362,N_15115,N_15240);
and U15363 (N_15363,N_15147,N_15216);
and U15364 (N_15364,N_15112,N_15099);
nor U15365 (N_15365,N_15201,N_15199);
nor U15366 (N_15366,N_15152,N_15245);
nor U15367 (N_15367,N_15145,N_15222);
nand U15368 (N_15368,N_15162,N_15224);
nand U15369 (N_15369,N_15016,N_15127);
nor U15370 (N_15370,N_15075,N_15223);
nand U15371 (N_15371,N_15193,N_15139);
nor U15372 (N_15372,N_15154,N_15058);
or U15373 (N_15373,N_15204,N_15230);
nand U15374 (N_15374,N_15126,N_15175);
or U15375 (N_15375,N_15027,N_15032);
or U15376 (N_15376,N_15170,N_15129);
and U15377 (N_15377,N_15187,N_15188);
and U15378 (N_15378,N_15055,N_15190);
or U15379 (N_15379,N_15193,N_15144);
nand U15380 (N_15380,N_15214,N_15108);
nand U15381 (N_15381,N_15123,N_15194);
nand U15382 (N_15382,N_15233,N_15228);
and U15383 (N_15383,N_15136,N_15220);
nand U15384 (N_15384,N_15127,N_15249);
and U15385 (N_15385,N_15048,N_15186);
or U15386 (N_15386,N_15003,N_15051);
and U15387 (N_15387,N_15089,N_15171);
nor U15388 (N_15388,N_15009,N_15035);
or U15389 (N_15389,N_15000,N_15029);
and U15390 (N_15390,N_15174,N_15149);
and U15391 (N_15391,N_15026,N_15038);
or U15392 (N_15392,N_15185,N_15127);
or U15393 (N_15393,N_15193,N_15119);
nand U15394 (N_15394,N_15039,N_15027);
or U15395 (N_15395,N_15090,N_15027);
nand U15396 (N_15396,N_15157,N_15207);
or U15397 (N_15397,N_15063,N_15198);
nand U15398 (N_15398,N_15115,N_15152);
nand U15399 (N_15399,N_15134,N_15216);
or U15400 (N_15400,N_15040,N_15081);
and U15401 (N_15401,N_15064,N_15009);
nand U15402 (N_15402,N_15125,N_15190);
or U15403 (N_15403,N_15210,N_15231);
xor U15404 (N_15404,N_15079,N_15230);
and U15405 (N_15405,N_15209,N_15171);
nor U15406 (N_15406,N_15003,N_15034);
nand U15407 (N_15407,N_15105,N_15150);
nand U15408 (N_15408,N_15131,N_15030);
and U15409 (N_15409,N_15199,N_15045);
or U15410 (N_15410,N_15207,N_15019);
nand U15411 (N_15411,N_15041,N_15122);
nor U15412 (N_15412,N_15151,N_15178);
or U15413 (N_15413,N_15042,N_15234);
nor U15414 (N_15414,N_15024,N_15117);
nand U15415 (N_15415,N_15028,N_15026);
xor U15416 (N_15416,N_15197,N_15038);
and U15417 (N_15417,N_15011,N_15222);
or U15418 (N_15418,N_15002,N_15030);
or U15419 (N_15419,N_15103,N_15237);
nor U15420 (N_15420,N_15152,N_15094);
nand U15421 (N_15421,N_15042,N_15214);
and U15422 (N_15422,N_15084,N_15172);
nand U15423 (N_15423,N_15180,N_15211);
nor U15424 (N_15424,N_15157,N_15237);
or U15425 (N_15425,N_15170,N_15037);
nor U15426 (N_15426,N_15242,N_15084);
and U15427 (N_15427,N_15177,N_15065);
nand U15428 (N_15428,N_15080,N_15210);
or U15429 (N_15429,N_15044,N_15164);
nor U15430 (N_15430,N_15106,N_15124);
nor U15431 (N_15431,N_15084,N_15076);
or U15432 (N_15432,N_15186,N_15198);
nand U15433 (N_15433,N_15145,N_15240);
and U15434 (N_15434,N_15241,N_15068);
and U15435 (N_15435,N_15195,N_15142);
nand U15436 (N_15436,N_15112,N_15226);
nor U15437 (N_15437,N_15244,N_15005);
nand U15438 (N_15438,N_15111,N_15092);
nand U15439 (N_15439,N_15242,N_15206);
or U15440 (N_15440,N_15193,N_15163);
and U15441 (N_15441,N_15217,N_15110);
nand U15442 (N_15442,N_15140,N_15069);
or U15443 (N_15443,N_15141,N_15140);
and U15444 (N_15444,N_15209,N_15219);
nor U15445 (N_15445,N_15091,N_15160);
nor U15446 (N_15446,N_15223,N_15197);
nand U15447 (N_15447,N_15043,N_15020);
nand U15448 (N_15448,N_15006,N_15104);
or U15449 (N_15449,N_15155,N_15107);
and U15450 (N_15450,N_15017,N_15184);
and U15451 (N_15451,N_15060,N_15089);
or U15452 (N_15452,N_15086,N_15221);
and U15453 (N_15453,N_15017,N_15034);
nor U15454 (N_15454,N_15231,N_15092);
or U15455 (N_15455,N_15247,N_15136);
xor U15456 (N_15456,N_15081,N_15149);
and U15457 (N_15457,N_15155,N_15105);
and U15458 (N_15458,N_15115,N_15001);
and U15459 (N_15459,N_15005,N_15174);
xor U15460 (N_15460,N_15015,N_15204);
xor U15461 (N_15461,N_15047,N_15162);
nand U15462 (N_15462,N_15236,N_15080);
nor U15463 (N_15463,N_15105,N_15234);
or U15464 (N_15464,N_15172,N_15045);
and U15465 (N_15465,N_15126,N_15063);
nor U15466 (N_15466,N_15207,N_15078);
or U15467 (N_15467,N_15237,N_15007);
and U15468 (N_15468,N_15028,N_15229);
or U15469 (N_15469,N_15183,N_15238);
and U15470 (N_15470,N_15223,N_15135);
nand U15471 (N_15471,N_15164,N_15220);
nor U15472 (N_15472,N_15209,N_15233);
nand U15473 (N_15473,N_15177,N_15035);
nand U15474 (N_15474,N_15174,N_15111);
nor U15475 (N_15475,N_15057,N_15142);
or U15476 (N_15476,N_15078,N_15165);
and U15477 (N_15477,N_15115,N_15147);
xnor U15478 (N_15478,N_15174,N_15242);
xnor U15479 (N_15479,N_15143,N_15069);
nand U15480 (N_15480,N_15221,N_15176);
nand U15481 (N_15481,N_15075,N_15040);
or U15482 (N_15482,N_15053,N_15244);
and U15483 (N_15483,N_15057,N_15075);
and U15484 (N_15484,N_15159,N_15103);
nor U15485 (N_15485,N_15238,N_15098);
xor U15486 (N_15486,N_15229,N_15240);
or U15487 (N_15487,N_15075,N_15234);
or U15488 (N_15488,N_15041,N_15040);
nor U15489 (N_15489,N_15088,N_15051);
xor U15490 (N_15490,N_15181,N_15199);
nand U15491 (N_15491,N_15107,N_15040);
nor U15492 (N_15492,N_15197,N_15238);
nor U15493 (N_15493,N_15008,N_15070);
nand U15494 (N_15494,N_15125,N_15010);
or U15495 (N_15495,N_15156,N_15021);
and U15496 (N_15496,N_15131,N_15059);
nor U15497 (N_15497,N_15246,N_15040);
and U15498 (N_15498,N_15214,N_15174);
nand U15499 (N_15499,N_15206,N_15094);
or U15500 (N_15500,N_15421,N_15424);
nor U15501 (N_15501,N_15403,N_15297);
xnor U15502 (N_15502,N_15451,N_15367);
or U15503 (N_15503,N_15287,N_15469);
nand U15504 (N_15504,N_15393,N_15271);
and U15505 (N_15505,N_15292,N_15251);
nor U15506 (N_15506,N_15395,N_15428);
nand U15507 (N_15507,N_15337,N_15381);
nor U15508 (N_15508,N_15334,N_15408);
nor U15509 (N_15509,N_15429,N_15448);
xor U15510 (N_15510,N_15455,N_15325);
or U15511 (N_15511,N_15301,N_15311);
nand U15512 (N_15512,N_15371,N_15364);
nand U15513 (N_15513,N_15348,N_15450);
or U15514 (N_15514,N_15291,N_15365);
nand U15515 (N_15515,N_15378,N_15274);
nand U15516 (N_15516,N_15306,N_15336);
and U15517 (N_15517,N_15338,N_15422);
or U15518 (N_15518,N_15404,N_15315);
nand U15519 (N_15519,N_15280,N_15376);
nand U15520 (N_15520,N_15405,N_15265);
nor U15521 (N_15521,N_15307,N_15354);
or U15522 (N_15522,N_15415,N_15452);
and U15523 (N_15523,N_15268,N_15281);
nor U15524 (N_15524,N_15407,N_15355);
and U15525 (N_15525,N_15495,N_15266);
and U15526 (N_15526,N_15313,N_15279);
nor U15527 (N_15527,N_15436,N_15487);
xnor U15528 (N_15528,N_15308,N_15396);
nor U15529 (N_15529,N_15445,N_15253);
nand U15530 (N_15530,N_15300,N_15299);
or U15531 (N_15531,N_15321,N_15277);
and U15532 (N_15532,N_15391,N_15317);
nor U15533 (N_15533,N_15411,N_15482);
nand U15534 (N_15534,N_15400,N_15419);
nor U15535 (N_15535,N_15256,N_15484);
nor U15536 (N_15536,N_15471,N_15432);
nor U15537 (N_15537,N_15352,N_15273);
or U15538 (N_15538,N_15453,N_15394);
xor U15539 (N_15539,N_15302,N_15449);
or U15540 (N_15540,N_15383,N_15476);
and U15541 (N_15541,N_15350,N_15288);
and U15542 (N_15542,N_15462,N_15374);
nor U15543 (N_15543,N_15314,N_15373);
nor U15544 (N_15544,N_15328,N_15435);
nor U15545 (N_15545,N_15434,N_15417);
nor U15546 (N_15546,N_15379,N_15282);
xor U15547 (N_15547,N_15456,N_15298);
nor U15548 (N_15548,N_15349,N_15262);
nor U15549 (N_15549,N_15255,N_15397);
and U15550 (N_15550,N_15473,N_15335);
nand U15551 (N_15551,N_15486,N_15330);
nand U15552 (N_15552,N_15464,N_15252);
nand U15553 (N_15553,N_15346,N_15358);
nand U15554 (N_15554,N_15284,N_15320);
nor U15555 (N_15555,N_15309,N_15363);
nand U15556 (N_15556,N_15490,N_15327);
or U15557 (N_15557,N_15390,N_15384);
and U15558 (N_15558,N_15339,N_15485);
nor U15559 (N_15559,N_15324,N_15410);
nor U15560 (N_15560,N_15446,N_15347);
nand U15561 (N_15561,N_15468,N_15312);
nor U15562 (N_15562,N_15488,N_15254);
nor U15563 (N_15563,N_15305,N_15402);
and U15564 (N_15564,N_15480,N_15294);
and U15565 (N_15565,N_15423,N_15406);
or U15566 (N_15566,N_15275,N_15440);
nand U15567 (N_15567,N_15351,N_15389);
or U15568 (N_15568,N_15409,N_15380);
nor U15569 (N_15569,N_15318,N_15319);
nand U15570 (N_15570,N_15303,N_15283);
and U15571 (N_15571,N_15276,N_15342);
nor U15572 (N_15572,N_15344,N_15343);
and U15573 (N_15573,N_15392,N_15472);
or U15574 (N_15574,N_15420,N_15295);
or U15575 (N_15575,N_15430,N_15426);
nand U15576 (N_15576,N_15413,N_15465);
nand U15577 (N_15577,N_15326,N_15382);
or U15578 (N_15578,N_15250,N_15362);
xnor U15579 (N_15579,N_15447,N_15479);
nor U15580 (N_15580,N_15458,N_15491);
nand U15581 (N_15581,N_15481,N_15401);
nand U15582 (N_15582,N_15498,N_15340);
nand U15583 (N_15583,N_15412,N_15427);
and U15584 (N_15584,N_15457,N_15475);
and U15585 (N_15585,N_15493,N_15441);
or U15586 (N_15586,N_15345,N_15377);
nand U15587 (N_15587,N_15269,N_15454);
nand U15588 (N_15588,N_15296,N_15261);
or U15589 (N_15589,N_15353,N_15375);
and U15590 (N_15590,N_15463,N_15263);
nor U15591 (N_15591,N_15399,N_15386);
or U15592 (N_15592,N_15433,N_15477);
or U15593 (N_15593,N_15304,N_15289);
or U15594 (N_15594,N_15368,N_15425);
nand U15595 (N_15595,N_15461,N_15466);
or U15596 (N_15596,N_15285,N_15489);
and U15597 (N_15597,N_15444,N_15499);
nand U15598 (N_15598,N_15310,N_15478);
nand U15599 (N_15599,N_15439,N_15356);
and U15600 (N_15600,N_15437,N_15372);
and U15601 (N_15601,N_15492,N_15467);
or U15602 (N_15602,N_15385,N_15278);
nor U15603 (N_15603,N_15470,N_15357);
nor U15604 (N_15604,N_15259,N_15360);
nand U15605 (N_15605,N_15323,N_15459);
nand U15606 (N_15606,N_15416,N_15359);
and U15607 (N_15607,N_15497,N_15267);
nand U15608 (N_15608,N_15370,N_15272);
or U15609 (N_15609,N_15290,N_15431);
and U15610 (N_15610,N_15361,N_15366);
nor U15611 (N_15611,N_15443,N_15460);
nor U15612 (N_15612,N_15331,N_15316);
nor U15613 (N_15613,N_15332,N_15496);
or U15614 (N_15614,N_15494,N_15414);
and U15615 (N_15615,N_15438,N_15341);
nor U15616 (N_15616,N_15260,N_15442);
nor U15617 (N_15617,N_15418,N_15388);
xnor U15618 (N_15618,N_15329,N_15333);
or U15619 (N_15619,N_15258,N_15293);
nand U15620 (N_15620,N_15270,N_15322);
and U15621 (N_15621,N_15286,N_15387);
nor U15622 (N_15622,N_15264,N_15474);
nor U15623 (N_15623,N_15369,N_15398);
or U15624 (N_15624,N_15483,N_15257);
or U15625 (N_15625,N_15483,N_15256);
nor U15626 (N_15626,N_15440,N_15259);
xor U15627 (N_15627,N_15389,N_15489);
xor U15628 (N_15628,N_15461,N_15359);
nor U15629 (N_15629,N_15395,N_15295);
nand U15630 (N_15630,N_15335,N_15250);
or U15631 (N_15631,N_15328,N_15477);
or U15632 (N_15632,N_15431,N_15425);
or U15633 (N_15633,N_15339,N_15353);
or U15634 (N_15634,N_15433,N_15465);
nand U15635 (N_15635,N_15451,N_15479);
nor U15636 (N_15636,N_15335,N_15480);
and U15637 (N_15637,N_15461,N_15322);
and U15638 (N_15638,N_15321,N_15447);
nand U15639 (N_15639,N_15477,N_15453);
or U15640 (N_15640,N_15251,N_15315);
nor U15641 (N_15641,N_15454,N_15302);
and U15642 (N_15642,N_15419,N_15312);
and U15643 (N_15643,N_15474,N_15335);
nor U15644 (N_15644,N_15480,N_15483);
nor U15645 (N_15645,N_15310,N_15432);
and U15646 (N_15646,N_15315,N_15363);
nand U15647 (N_15647,N_15449,N_15314);
and U15648 (N_15648,N_15418,N_15373);
nand U15649 (N_15649,N_15382,N_15404);
nand U15650 (N_15650,N_15301,N_15471);
or U15651 (N_15651,N_15390,N_15268);
nor U15652 (N_15652,N_15340,N_15363);
nor U15653 (N_15653,N_15482,N_15260);
or U15654 (N_15654,N_15290,N_15332);
xnor U15655 (N_15655,N_15496,N_15495);
nor U15656 (N_15656,N_15290,N_15272);
or U15657 (N_15657,N_15309,N_15366);
or U15658 (N_15658,N_15415,N_15264);
or U15659 (N_15659,N_15417,N_15333);
or U15660 (N_15660,N_15316,N_15373);
nor U15661 (N_15661,N_15348,N_15432);
nand U15662 (N_15662,N_15326,N_15308);
and U15663 (N_15663,N_15351,N_15458);
and U15664 (N_15664,N_15437,N_15483);
nor U15665 (N_15665,N_15394,N_15402);
xnor U15666 (N_15666,N_15254,N_15283);
xnor U15667 (N_15667,N_15470,N_15302);
nand U15668 (N_15668,N_15339,N_15456);
xor U15669 (N_15669,N_15353,N_15455);
and U15670 (N_15670,N_15474,N_15456);
or U15671 (N_15671,N_15401,N_15405);
or U15672 (N_15672,N_15362,N_15372);
and U15673 (N_15673,N_15411,N_15490);
nor U15674 (N_15674,N_15469,N_15310);
nand U15675 (N_15675,N_15345,N_15490);
nand U15676 (N_15676,N_15399,N_15304);
or U15677 (N_15677,N_15305,N_15411);
and U15678 (N_15678,N_15482,N_15453);
and U15679 (N_15679,N_15428,N_15313);
xor U15680 (N_15680,N_15488,N_15496);
nand U15681 (N_15681,N_15431,N_15300);
and U15682 (N_15682,N_15441,N_15410);
or U15683 (N_15683,N_15307,N_15421);
nand U15684 (N_15684,N_15347,N_15372);
nor U15685 (N_15685,N_15489,N_15322);
nand U15686 (N_15686,N_15432,N_15346);
and U15687 (N_15687,N_15276,N_15314);
nor U15688 (N_15688,N_15326,N_15353);
nand U15689 (N_15689,N_15264,N_15383);
or U15690 (N_15690,N_15454,N_15487);
nor U15691 (N_15691,N_15367,N_15261);
or U15692 (N_15692,N_15457,N_15302);
nor U15693 (N_15693,N_15290,N_15296);
xor U15694 (N_15694,N_15387,N_15270);
or U15695 (N_15695,N_15437,N_15493);
nand U15696 (N_15696,N_15435,N_15260);
and U15697 (N_15697,N_15312,N_15333);
and U15698 (N_15698,N_15343,N_15252);
xor U15699 (N_15699,N_15321,N_15498);
and U15700 (N_15700,N_15479,N_15250);
and U15701 (N_15701,N_15311,N_15445);
nor U15702 (N_15702,N_15497,N_15375);
xor U15703 (N_15703,N_15448,N_15473);
nor U15704 (N_15704,N_15253,N_15386);
or U15705 (N_15705,N_15454,N_15495);
nand U15706 (N_15706,N_15256,N_15281);
nand U15707 (N_15707,N_15275,N_15424);
nor U15708 (N_15708,N_15273,N_15262);
and U15709 (N_15709,N_15414,N_15429);
nand U15710 (N_15710,N_15307,N_15346);
or U15711 (N_15711,N_15411,N_15458);
nor U15712 (N_15712,N_15282,N_15474);
nand U15713 (N_15713,N_15356,N_15486);
and U15714 (N_15714,N_15250,N_15324);
nand U15715 (N_15715,N_15417,N_15436);
nand U15716 (N_15716,N_15302,N_15462);
and U15717 (N_15717,N_15481,N_15495);
xor U15718 (N_15718,N_15442,N_15332);
or U15719 (N_15719,N_15281,N_15422);
and U15720 (N_15720,N_15261,N_15294);
xor U15721 (N_15721,N_15293,N_15434);
nand U15722 (N_15722,N_15474,N_15457);
or U15723 (N_15723,N_15470,N_15473);
or U15724 (N_15724,N_15407,N_15269);
or U15725 (N_15725,N_15327,N_15260);
xor U15726 (N_15726,N_15297,N_15477);
nor U15727 (N_15727,N_15281,N_15430);
or U15728 (N_15728,N_15482,N_15491);
and U15729 (N_15729,N_15278,N_15414);
nand U15730 (N_15730,N_15373,N_15353);
or U15731 (N_15731,N_15457,N_15491);
nor U15732 (N_15732,N_15424,N_15408);
nand U15733 (N_15733,N_15439,N_15303);
or U15734 (N_15734,N_15271,N_15413);
nor U15735 (N_15735,N_15498,N_15376);
nand U15736 (N_15736,N_15485,N_15319);
nand U15737 (N_15737,N_15441,N_15449);
and U15738 (N_15738,N_15295,N_15360);
and U15739 (N_15739,N_15478,N_15464);
nand U15740 (N_15740,N_15457,N_15391);
nor U15741 (N_15741,N_15430,N_15454);
and U15742 (N_15742,N_15410,N_15282);
and U15743 (N_15743,N_15406,N_15486);
nand U15744 (N_15744,N_15485,N_15434);
nor U15745 (N_15745,N_15439,N_15406);
and U15746 (N_15746,N_15329,N_15486);
xor U15747 (N_15747,N_15437,N_15313);
nand U15748 (N_15748,N_15405,N_15439);
and U15749 (N_15749,N_15406,N_15388);
nor U15750 (N_15750,N_15690,N_15614);
and U15751 (N_15751,N_15543,N_15645);
or U15752 (N_15752,N_15596,N_15574);
nand U15753 (N_15753,N_15508,N_15653);
and U15754 (N_15754,N_15749,N_15619);
nor U15755 (N_15755,N_15666,N_15697);
nand U15756 (N_15756,N_15707,N_15718);
and U15757 (N_15757,N_15580,N_15513);
nor U15758 (N_15758,N_15684,N_15665);
or U15759 (N_15759,N_15618,N_15539);
or U15760 (N_15760,N_15724,N_15521);
or U15761 (N_15761,N_15719,N_15652);
or U15762 (N_15762,N_15698,N_15639);
or U15763 (N_15763,N_15609,N_15623);
or U15764 (N_15764,N_15607,N_15629);
nand U15765 (N_15765,N_15627,N_15567);
and U15766 (N_15766,N_15660,N_15691);
or U15767 (N_15767,N_15694,N_15667);
nand U15768 (N_15768,N_15516,N_15727);
nor U15769 (N_15769,N_15664,N_15599);
nand U15770 (N_15770,N_15601,N_15568);
or U15771 (N_15771,N_15566,N_15522);
nor U15772 (N_15772,N_15529,N_15687);
nand U15773 (N_15773,N_15643,N_15569);
and U15774 (N_15774,N_15524,N_15525);
nand U15775 (N_15775,N_15734,N_15702);
nand U15776 (N_15776,N_15725,N_15688);
nor U15777 (N_15777,N_15588,N_15530);
or U15778 (N_15778,N_15547,N_15693);
or U15779 (N_15779,N_15650,N_15642);
and U15780 (N_15780,N_15681,N_15542);
nor U15781 (N_15781,N_15550,N_15748);
xor U15782 (N_15782,N_15502,N_15575);
or U15783 (N_15783,N_15680,N_15590);
and U15784 (N_15784,N_15617,N_15635);
or U15785 (N_15785,N_15597,N_15742);
xor U15786 (N_15786,N_15729,N_15555);
and U15787 (N_15787,N_15556,N_15634);
nor U15788 (N_15788,N_15579,N_15517);
nor U15789 (N_15789,N_15583,N_15740);
and U15790 (N_15790,N_15705,N_15658);
nor U15791 (N_15791,N_15551,N_15535);
nand U15792 (N_15792,N_15577,N_15563);
and U15793 (N_15793,N_15527,N_15509);
and U15794 (N_15794,N_15704,N_15626);
nor U15795 (N_15795,N_15602,N_15651);
nor U15796 (N_15796,N_15578,N_15710);
xor U15797 (N_15797,N_15662,N_15655);
nor U15798 (N_15798,N_15512,N_15659);
and U15799 (N_15799,N_15562,N_15733);
nor U15800 (N_15800,N_15552,N_15739);
nor U15801 (N_15801,N_15743,N_15554);
nand U15802 (N_15802,N_15671,N_15620);
nand U15803 (N_15803,N_15510,N_15615);
nor U15804 (N_15804,N_15696,N_15737);
xnor U15805 (N_15805,N_15637,N_15648);
xnor U15806 (N_15806,N_15631,N_15561);
nand U15807 (N_15807,N_15703,N_15537);
and U15808 (N_15808,N_15582,N_15689);
or U15809 (N_15809,N_15676,N_15553);
and U15810 (N_15810,N_15505,N_15683);
or U15811 (N_15811,N_15685,N_15745);
nor U15812 (N_15812,N_15589,N_15514);
nand U15813 (N_15813,N_15647,N_15721);
or U15814 (N_15814,N_15538,N_15591);
nor U15815 (N_15815,N_15669,N_15560);
xor U15816 (N_15816,N_15515,N_15730);
nor U15817 (N_15817,N_15570,N_15576);
nor U15818 (N_15818,N_15732,N_15564);
or U15819 (N_15819,N_15741,N_15519);
nor U15820 (N_15820,N_15621,N_15507);
and U15821 (N_15821,N_15706,N_15641);
nand U15822 (N_15822,N_15501,N_15565);
or U15823 (N_15823,N_15675,N_15610);
nor U15824 (N_15824,N_15709,N_15544);
nor U15825 (N_15825,N_15678,N_15686);
and U15826 (N_15826,N_15715,N_15711);
nand U15827 (N_15827,N_15649,N_15605);
and U15828 (N_15828,N_15500,N_15644);
and U15829 (N_15829,N_15661,N_15624);
xnor U15830 (N_15830,N_15673,N_15593);
nor U15831 (N_15831,N_15573,N_15726);
or U15832 (N_15832,N_15598,N_15528);
nor U15833 (N_15833,N_15511,N_15677);
xnor U15834 (N_15834,N_15723,N_15746);
nand U15835 (N_15835,N_15592,N_15572);
and U15836 (N_15836,N_15633,N_15587);
or U15837 (N_15837,N_15716,N_15744);
nand U15838 (N_15838,N_15548,N_15594);
and U15839 (N_15839,N_15526,N_15520);
or U15840 (N_15840,N_15714,N_15581);
nand U15841 (N_15841,N_15612,N_15630);
and U15842 (N_15842,N_15540,N_15603);
nand U15843 (N_15843,N_15747,N_15503);
nor U15844 (N_15844,N_15534,N_15692);
and U15845 (N_15845,N_15628,N_15533);
nor U15846 (N_15846,N_15622,N_15695);
nand U15847 (N_15847,N_15504,N_15640);
and U15848 (N_15848,N_15546,N_15604);
xor U15849 (N_15849,N_15549,N_15632);
nor U15850 (N_15850,N_15600,N_15638);
and U15851 (N_15851,N_15506,N_15700);
or U15852 (N_15852,N_15532,N_15646);
nand U15853 (N_15853,N_15682,N_15668);
nand U15854 (N_15854,N_15735,N_15670);
nor U15855 (N_15855,N_15713,N_15679);
nor U15856 (N_15856,N_15731,N_15586);
nor U15857 (N_15857,N_15736,N_15523);
nor U15858 (N_15858,N_15738,N_15571);
nand U15859 (N_15859,N_15595,N_15616);
or U15860 (N_15860,N_15541,N_15654);
or U15861 (N_15861,N_15636,N_15717);
or U15862 (N_15862,N_15531,N_15606);
or U15863 (N_15863,N_15585,N_15625);
nand U15864 (N_15864,N_15558,N_15657);
or U15865 (N_15865,N_15557,N_15613);
nor U15866 (N_15866,N_15518,N_15722);
nor U15867 (N_15867,N_15728,N_15663);
and U15868 (N_15868,N_15536,N_15712);
xnor U15869 (N_15869,N_15559,N_15584);
nor U15870 (N_15870,N_15656,N_15720);
nand U15871 (N_15871,N_15674,N_15608);
and U15872 (N_15872,N_15545,N_15708);
and U15873 (N_15873,N_15611,N_15701);
or U15874 (N_15874,N_15699,N_15672);
and U15875 (N_15875,N_15729,N_15585);
nor U15876 (N_15876,N_15572,N_15659);
or U15877 (N_15877,N_15550,N_15668);
xnor U15878 (N_15878,N_15741,N_15595);
or U15879 (N_15879,N_15693,N_15730);
or U15880 (N_15880,N_15609,N_15612);
and U15881 (N_15881,N_15689,N_15620);
or U15882 (N_15882,N_15575,N_15610);
nor U15883 (N_15883,N_15508,N_15552);
or U15884 (N_15884,N_15508,N_15567);
nand U15885 (N_15885,N_15551,N_15573);
xnor U15886 (N_15886,N_15626,N_15637);
nor U15887 (N_15887,N_15552,N_15599);
nand U15888 (N_15888,N_15541,N_15550);
or U15889 (N_15889,N_15526,N_15655);
nor U15890 (N_15890,N_15657,N_15593);
or U15891 (N_15891,N_15687,N_15564);
nand U15892 (N_15892,N_15708,N_15560);
nor U15893 (N_15893,N_15654,N_15555);
nand U15894 (N_15894,N_15552,N_15547);
and U15895 (N_15895,N_15722,N_15715);
and U15896 (N_15896,N_15619,N_15716);
or U15897 (N_15897,N_15746,N_15534);
xor U15898 (N_15898,N_15621,N_15559);
nor U15899 (N_15899,N_15706,N_15582);
nand U15900 (N_15900,N_15740,N_15504);
xnor U15901 (N_15901,N_15632,N_15749);
or U15902 (N_15902,N_15651,N_15500);
nand U15903 (N_15903,N_15540,N_15574);
nand U15904 (N_15904,N_15627,N_15548);
xnor U15905 (N_15905,N_15723,N_15653);
and U15906 (N_15906,N_15659,N_15733);
nor U15907 (N_15907,N_15738,N_15661);
nor U15908 (N_15908,N_15573,N_15708);
and U15909 (N_15909,N_15698,N_15663);
or U15910 (N_15910,N_15630,N_15672);
and U15911 (N_15911,N_15718,N_15562);
nand U15912 (N_15912,N_15712,N_15647);
xor U15913 (N_15913,N_15603,N_15548);
and U15914 (N_15914,N_15655,N_15530);
and U15915 (N_15915,N_15676,N_15654);
or U15916 (N_15916,N_15651,N_15636);
and U15917 (N_15917,N_15692,N_15726);
or U15918 (N_15918,N_15737,N_15588);
xnor U15919 (N_15919,N_15745,N_15583);
nor U15920 (N_15920,N_15696,N_15545);
or U15921 (N_15921,N_15620,N_15632);
and U15922 (N_15922,N_15500,N_15516);
or U15923 (N_15923,N_15559,N_15684);
nor U15924 (N_15924,N_15520,N_15632);
xnor U15925 (N_15925,N_15699,N_15629);
and U15926 (N_15926,N_15563,N_15696);
nand U15927 (N_15927,N_15512,N_15579);
xor U15928 (N_15928,N_15596,N_15672);
and U15929 (N_15929,N_15603,N_15564);
nand U15930 (N_15930,N_15673,N_15675);
and U15931 (N_15931,N_15504,N_15728);
and U15932 (N_15932,N_15649,N_15515);
or U15933 (N_15933,N_15680,N_15616);
or U15934 (N_15934,N_15597,N_15607);
or U15935 (N_15935,N_15529,N_15680);
or U15936 (N_15936,N_15696,N_15624);
nand U15937 (N_15937,N_15572,N_15679);
nand U15938 (N_15938,N_15596,N_15723);
nor U15939 (N_15939,N_15520,N_15719);
nand U15940 (N_15940,N_15656,N_15675);
nor U15941 (N_15941,N_15650,N_15711);
nor U15942 (N_15942,N_15550,N_15536);
and U15943 (N_15943,N_15606,N_15745);
and U15944 (N_15944,N_15564,N_15517);
and U15945 (N_15945,N_15701,N_15603);
or U15946 (N_15946,N_15639,N_15634);
xnor U15947 (N_15947,N_15710,N_15509);
nor U15948 (N_15948,N_15641,N_15514);
nand U15949 (N_15949,N_15702,N_15731);
nand U15950 (N_15950,N_15657,N_15667);
nand U15951 (N_15951,N_15587,N_15725);
nand U15952 (N_15952,N_15510,N_15732);
and U15953 (N_15953,N_15599,N_15712);
nor U15954 (N_15954,N_15646,N_15517);
xnor U15955 (N_15955,N_15572,N_15660);
nand U15956 (N_15956,N_15666,N_15560);
nand U15957 (N_15957,N_15710,N_15585);
nand U15958 (N_15958,N_15554,N_15539);
nor U15959 (N_15959,N_15562,N_15622);
nor U15960 (N_15960,N_15535,N_15543);
or U15961 (N_15961,N_15542,N_15585);
and U15962 (N_15962,N_15547,N_15702);
nand U15963 (N_15963,N_15507,N_15657);
nand U15964 (N_15964,N_15733,N_15739);
nor U15965 (N_15965,N_15543,N_15594);
or U15966 (N_15966,N_15688,N_15573);
nor U15967 (N_15967,N_15592,N_15589);
xor U15968 (N_15968,N_15697,N_15692);
and U15969 (N_15969,N_15555,N_15738);
and U15970 (N_15970,N_15565,N_15695);
nor U15971 (N_15971,N_15579,N_15572);
nor U15972 (N_15972,N_15526,N_15505);
xor U15973 (N_15973,N_15548,N_15683);
nor U15974 (N_15974,N_15715,N_15602);
nor U15975 (N_15975,N_15508,N_15707);
and U15976 (N_15976,N_15727,N_15715);
nand U15977 (N_15977,N_15519,N_15715);
nor U15978 (N_15978,N_15746,N_15606);
or U15979 (N_15979,N_15602,N_15596);
nand U15980 (N_15980,N_15665,N_15580);
and U15981 (N_15981,N_15609,N_15563);
and U15982 (N_15982,N_15605,N_15630);
nand U15983 (N_15983,N_15746,N_15667);
nor U15984 (N_15984,N_15526,N_15600);
or U15985 (N_15985,N_15657,N_15561);
nand U15986 (N_15986,N_15737,N_15559);
or U15987 (N_15987,N_15572,N_15563);
xor U15988 (N_15988,N_15657,N_15607);
or U15989 (N_15989,N_15569,N_15624);
and U15990 (N_15990,N_15599,N_15742);
nand U15991 (N_15991,N_15615,N_15640);
nor U15992 (N_15992,N_15558,N_15574);
xor U15993 (N_15993,N_15732,N_15651);
or U15994 (N_15994,N_15715,N_15673);
nor U15995 (N_15995,N_15633,N_15735);
nor U15996 (N_15996,N_15724,N_15610);
and U15997 (N_15997,N_15552,N_15646);
nand U15998 (N_15998,N_15648,N_15604);
or U15999 (N_15999,N_15541,N_15658);
nor U16000 (N_16000,N_15768,N_15761);
nor U16001 (N_16001,N_15938,N_15787);
and U16002 (N_16002,N_15861,N_15809);
nor U16003 (N_16003,N_15990,N_15961);
nand U16004 (N_16004,N_15802,N_15808);
nor U16005 (N_16005,N_15998,N_15979);
xnor U16006 (N_16006,N_15828,N_15889);
nand U16007 (N_16007,N_15759,N_15864);
and U16008 (N_16008,N_15976,N_15982);
xnor U16009 (N_16009,N_15912,N_15935);
or U16010 (N_16010,N_15795,N_15902);
nor U16011 (N_16011,N_15874,N_15868);
or U16012 (N_16012,N_15940,N_15806);
nor U16013 (N_16013,N_15904,N_15962);
and U16014 (N_16014,N_15816,N_15996);
nand U16015 (N_16015,N_15790,N_15815);
or U16016 (N_16016,N_15865,N_15754);
nor U16017 (N_16017,N_15972,N_15992);
xnor U16018 (N_16018,N_15769,N_15755);
and U16019 (N_16019,N_15948,N_15870);
or U16020 (N_16020,N_15873,N_15953);
nand U16021 (N_16021,N_15977,N_15974);
nor U16022 (N_16022,N_15975,N_15852);
and U16023 (N_16023,N_15871,N_15872);
nand U16024 (N_16024,N_15867,N_15877);
xor U16025 (N_16025,N_15941,N_15841);
xor U16026 (N_16026,N_15956,N_15993);
nor U16027 (N_16027,N_15763,N_15910);
xor U16028 (N_16028,N_15777,N_15931);
nor U16029 (N_16029,N_15804,N_15882);
and U16030 (N_16030,N_15911,N_15897);
nand U16031 (N_16031,N_15752,N_15876);
nor U16032 (N_16032,N_15893,N_15926);
nand U16033 (N_16033,N_15793,N_15879);
nor U16034 (N_16034,N_15950,N_15837);
nand U16035 (N_16035,N_15934,N_15830);
or U16036 (N_16036,N_15778,N_15963);
nand U16037 (N_16037,N_15878,N_15775);
and U16038 (N_16038,N_15845,N_15818);
nor U16039 (N_16039,N_15805,N_15796);
nor U16040 (N_16040,N_15967,N_15855);
nor U16041 (N_16041,N_15903,N_15987);
nand U16042 (N_16042,N_15829,N_15881);
nand U16043 (N_16043,N_15901,N_15913);
and U16044 (N_16044,N_15801,N_15899);
or U16045 (N_16045,N_15853,N_15789);
or U16046 (N_16046,N_15946,N_15863);
and U16047 (N_16047,N_15764,N_15827);
nor U16048 (N_16048,N_15826,N_15915);
nor U16049 (N_16049,N_15905,N_15997);
nor U16050 (N_16050,N_15986,N_15779);
or U16051 (N_16051,N_15758,N_15887);
nor U16052 (N_16052,N_15896,N_15980);
and U16053 (N_16053,N_15858,N_15782);
or U16054 (N_16054,N_15957,N_15774);
or U16055 (N_16055,N_15952,N_15895);
xnor U16056 (N_16056,N_15866,N_15919);
nand U16057 (N_16057,N_15978,N_15999);
nor U16058 (N_16058,N_15995,N_15890);
nor U16059 (N_16059,N_15844,N_15908);
nand U16060 (N_16060,N_15851,N_15854);
nor U16061 (N_16061,N_15825,N_15760);
nor U16062 (N_16062,N_15925,N_15924);
and U16063 (N_16063,N_15822,N_15862);
xor U16064 (N_16064,N_15847,N_15799);
nor U16065 (N_16065,N_15892,N_15835);
xnor U16066 (N_16066,N_15970,N_15791);
xnor U16067 (N_16067,N_15824,N_15770);
nand U16068 (N_16068,N_15803,N_15918);
and U16069 (N_16069,N_15885,N_15785);
nand U16070 (N_16070,N_15848,N_15914);
or U16071 (N_16071,N_15906,N_15860);
and U16072 (N_16072,N_15772,N_15943);
or U16073 (N_16073,N_15836,N_15766);
and U16074 (N_16074,N_15944,N_15811);
and U16075 (N_16075,N_15928,N_15788);
and U16076 (N_16076,N_15959,N_15831);
nor U16077 (N_16077,N_15888,N_15939);
nand U16078 (N_16078,N_15923,N_15960);
nand U16079 (N_16079,N_15984,N_15771);
nor U16080 (N_16080,N_15821,N_15880);
or U16081 (N_16081,N_15898,N_15762);
nand U16082 (N_16082,N_15842,N_15843);
and U16083 (N_16083,N_15932,N_15966);
or U16084 (N_16084,N_15994,N_15930);
nand U16085 (N_16085,N_15800,N_15832);
nor U16086 (N_16086,N_15951,N_15968);
and U16087 (N_16087,N_15813,N_15786);
xnor U16088 (N_16088,N_15798,N_15814);
nand U16089 (N_16089,N_15794,N_15783);
nand U16090 (N_16090,N_15884,N_15776);
or U16091 (N_16091,N_15920,N_15933);
nand U16092 (N_16092,N_15927,N_15954);
nor U16093 (N_16093,N_15929,N_15989);
or U16094 (N_16094,N_15753,N_15833);
nor U16095 (N_16095,N_15859,N_15857);
nand U16096 (N_16096,N_15947,N_15936);
xor U16097 (N_16097,N_15909,N_15945);
or U16098 (N_16098,N_15869,N_15988);
nand U16099 (N_16099,N_15767,N_15894);
and U16100 (N_16100,N_15991,N_15823);
nor U16101 (N_16101,N_15916,N_15765);
and U16102 (N_16102,N_15875,N_15750);
and U16103 (N_16103,N_15840,N_15757);
nor U16104 (N_16104,N_15942,N_15964);
and U16105 (N_16105,N_15839,N_15751);
nand U16106 (N_16106,N_15838,N_15773);
nand U16107 (N_16107,N_15958,N_15797);
xnor U16108 (N_16108,N_15792,N_15955);
nand U16109 (N_16109,N_15850,N_15781);
nand U16110 (N_16110,N_15812,N_15917);
and U16111 (N_16111,N_15810,N_15985);
or U16112 (N_16112,N_15922,N_15891);
xor U16113 (N_16113,N_15900,N_15907);
nor U16114 (N_16114,N_15780,N_15983);
or U16115 (N_16115,N_15846,N_15973);
nand U16116 (N_16116,N_15756,N_15849);
nor U16117 (N_16117,N_15820,N_15886);
nor U16118 (N_16118,N_15971,N_15807);
nor U16119 (N_16119,N_15921,N_15817);
nand U16120 (N_16120,N_15819,N_15949);
nand U16121 (N_16121,N_15834,N_15965);
nand U16122 (N_16122,N_15969,N_15937);
xor U16123 (N_16123,N_15883,N_15856);
nand U16124 (N_16124,N_15981,N_15784);
nand U16125 (N_16125,N_15863,N_15910);
or U16126 (N_16126,N_15894,N_15992);
and U16127 (N_16127,N_15786,N_15870);
or U16128 (N_16128,N_15993,N_15856);
and U16129 (N_16129,N_15969,N_15894);
nor U16130 (N_16130,N_15876,N_15849);
nor U16131 (N_16131,N_15978,N_15755);
nand U16132 (N_16132,N_15926,N_15936);
nor U16133 (N_16133,N_15947,N_15975);
or U16134 (N_16134,N_15768,N_15927);
nand U16135 (N_16135,N_15899,N_15842);
nand U16136 (N_16136,N_15882,N_15825);
xor U16137 (N_16137,N_15766,N_15824);
nand U16138 (N_16138,N_15988,N_15877);
and U16139 (N_16139,N_15992,N_15853);
nand U16140 (N_16140,N_15854,N_15810);
nand U16141 (N_16141,N_15919,N_15807);
nor U16142 (N_16142,N_15769,N_15902);
xnor U16143 (N_16143,N_15913,N_15950);
xnor U16144 (N_16144,N_15770,N_15811);
xnor U16145 (N_16145,N_15790,N_15816);
or U16146 (N_16146,N_15986,N_15917);
nor U16147 (N_16147,N_15949,N_15838);
or U16148 (N_16148,N_15809,N_15759);
nor U16149 (N_16149,N_15962,N_15804);
nand U16150 (N_16150,N_15987,N_15870);
or U16151 (N_16151,N_15985,N_15792);
nand U16152 (N_16152,N_15943,N_15924);
xnor U16153 (N_16153,N_15927,N_15882);
nand U16154 (N_16154,N_15778,N_15826);
or U16155 (N_16155,N_15757,N_15845);
nand U16156 (N_16156,N_15788,N_15987);
nand U16157 (N_16157,N_15880,N_15851);
nand U16158 (N_16158,N_15840,N_15861);
nand U16159 (N_16159,N_15987,N_15864);
and U16160 (N_16160,N_15963,N_15894);
and U16161 (N_16161,N_15874,N_15755);
nand U16162 (N_16162,N_15916,N_15921);
or U16163 (N_16163,N_15854,N_15954);
nand U16164 (N_16164,N_15874,N_15910);
xor U16165 (N_16165,N_15981,N_15781);
nand U16166 (N_16166,N_15836,N_15774);
nor U16167 (N_16167,N_15999,N_15831);
and U16168 (N_16168,N_15786,N_15820);
or U16169 (N_16169,N_15814,N_15986);
nand U16170 (N_16170,N_15952,N_15967);
or U16171 (N_16171,N_15919,N_15930);
nand U16172 (N_16172,N_15844,N_15772);
or U16173 (N_16173,N_15758,N_15862);
nand U16174 (N_16174,N_15804,N_15988);
or U16175 (N_16175,N_15873,N_15961);
and U16176 (N_16176,N_15930,N_15783);
and U16177 (N_16177,N_15874,N_15919);
and U16178 (N_16178,N_15956,N_15766);
xnor U16179 (N_16179,N_15936,N_15903);
or U16180 (N_16180,N_15901,N_15751);
nor U16181 (N_16181,N_15941,N_15932);
or U16182 (N_16182,N_15874,N_15982);
or U16183 (N_16183,N_15850,N_15753);
or U16184 (N_16184,N_15926,N_15841);
or U16185 (N_16185,N_15844,N_15938);
and U16186 (N_16186,N_15877,N_15967);
xnor U16187 (N_16187,N_15895,N_15773);
nor U16188 (N_16188,N_15877,N_15751);
and U16189 (N_16189,N_15856,N_15771);
or U16190 (N_16190,N_15907,N_15947);
or U16191 (N_16191,N_15876,N_15987);
nand U16192 (N_16192,N_15888,N_15756);
and U16193 (N_16193,N_15843,N_15862);
and U16194 (N_16194,N_15966,N_15845);
nand U16195 (N_16195,N_15810,N_15918);
and U16196 (N_16196,N_15760,N_15886);
xnor U16197 (N_16197,N_15910,N_15995);
or U16198 (N_16198,N_15815,N_15857);
nand U16199 (N_16199,N_15754,N_15930);
nor U16200 (N_16200,N_15988,N_15950);
xor U16201 (N_16201,N_15953,N_15776);
and U16202 (N_16202,N_15826,N_15989);
nor U16203 (N_16203,N_15858,N_15978);
nand U16204 (N_16204,N_15854,N_15751);
nor U16205 (N_16205,N_15923,N_15775);
nand U16206 (N_16206,N_15811,N_15989);
or U16207 (N_16207,N_15896,N_15759);
xor U16208 (N_16208,N_15815,N_15877);
nor U16209 (N_16209,N_15951,N_15949);
nand U16210 (N_16210,N_15981,N_15787);
nor U16211 (N_16211,N_15929,N_15811);
nor U16212 (N_16212,N_15911,N_15853);
and U16213 (N_16213,N_15969,N_15956);
nand U16214 (N_16214,N_15781,N_15831);
nand U16215 (N_16215,N_15952,N_15914);
xnor U16216 (N_16216,N_15966,N_15876);
nand U16217 (N_16217,N_15861,N_15834);
xnor U16218 (N_16218,N_15937,N_15786);
nand U16219 (N_16219,N_15940,N_15825);
and U16220 (N_16220,N_15900,N_15984);
nand U16221 (N_16221,N_15853,N_15850);
and U16222 (N_16222,N_15862,N_15942);
or U16223 (N_16223,N_15762,N_15881);
nor U16224 (N_16224,N_15952,N_15788);
xnor U16225 (N_16225,N_15900,N_15983);
nand U16226 (N_16226,N_15918,N_15900);
nor U16227 (N_16227,N_15803,N_15786);
or U16228 (N_16228,N_15964,N_15883);
nand U16229 (N_16229,N_15821,N_15799);
or U16230 (N_16230,N_15845,N_15751);
or U16231 (N_16231,N_15781,N_15809);
or U16232 (N_16232,N_15914,N_15817);
nand U16233 (N_16233,N_15935,N_15796);
and U16234 (N_16234,N_15984,N_15766);
nand U16235 (N_16235,N_15816,N_15975);
or U16236 (N_16236,N_15951,N_15853);
and U16237 (N_16237,N_15874,N_15977);
or U16238 (N_16238,N_15825,N_15976);
nor U16239 (N_16239,N_15902,N_15825);
nand U16240 (N_16240,N_15885,N_15755);
nand U16241 (N_16241,N_15762,N_15937);
and U16242 (N_16242,N_15843,N_15904);
nand U16243 (N_16243,N_15987,N_15827);
xor U16244 (N_16244,N_15831,N_15859);
nand U16245 (N_16245,N_15961,N_15911);
nor U16246 (N_16246,N_15756,N_15772);
and U16247 (N_16247,N_15782,N_15781);
or U16248 (N_16248,N_15755,N_15867);
nand U16249 (N_16249,N_15927,N_15962);
nor U16250 (N_16250,N_16232,N_16039);
nand U16251 (N_16251,N_16211,N_16041);
nor U16252 (N_16252,N_16019,N_16246);
nor U16253 (N_16253,N_16035,N_16215);
nor U16254 (N_16254,N_16025,N_16114);
nor U16255 (N_16255,N_16173,N_16070);
nor U16256 (N_16256,N_16110,N_16089);
or U16257 (N_16257,N_16013,N_16068);
and U16258 (N_16258,N_16072,N_16037);
and U16259 (N_16259,N_16212,N_16238);
and U16260 (N_16260,N_16117,N_16091);
xor U16261 (N_16261,N_16048,N_16154);
nor U16262 (N_16262,N_16209,N_16051);
xor U16263 (N_16263,N_16180,N_16160);
nand U16264 (N_16264,N_16038,N_16172);
nand U16265 (N_16265,N_16121,N_16189);
nor U16266 (N_16266,N_16171,N_16136);
and U16267 (N_16267,N_16186,N_16129);
nand U16268 (N_16268,N_16236,N_16231);
or U16269 (N_16269,N_16248,N_16020);
and U16270 (N_16270,N_16198,N_16216);
nand U16271 (N_16271,N_16144,N_16204);
and U16272 (N_16272,N_16192,N_16014);
and U16273 (N_16273,N_16179,N_16240);
nor U16274 (N_16274,N_16078,N_16193);
nor U16275 (N_16275,N_16113,N_16063);
nand U16276 (N_16276,N_16067,N_16184);
or U16277 (N_16277,N_16061,N_16194);
xnor U16278 (N_16278,N_16124,N_16066);
and U16279 (N_16279,N_16233,N_16191);
and U16280 (N_16280,N_16178,N_16017);
and U16281 (N_16281,N_16137,N_16128);
and U16282 (N_16282,N_16029,N_16023);
or U16283 (N_16283,N_16073,N_16177);
or U16284 (N_16284,N_16057,N_16226);
and U16285 (N_16285,N_16123,N_16045);
nor U16286 (N_16286,N_16166,N_16127);
and U16287 (N_16287,N_16132,N_16008);
xor U16288 (N_16288,N_16043,N_16203);
nand U16289 (N_16289,N_16021,N_16060);
nor U16290 (N_16290,N_16088,N_16143);
nor U16291 (N_16291,N_16028,N_16097);
nor U16292 (N_16292,N_16222,N_16183);
or U16293 (N_16293,N_16015,N_16100);
and U16294 (N_16294,N_16010,N_16182);
or U16295 (N_16295,N_16138,N_16086);
xnor U16296 (N_16296,N_16170,N_16081);
or U16297 (N_16297,N_16167,N_16082);
nand U16298 (N_16298,N_16053,N_16148);
nand U16299 (N_16299,N_16224,N_16220);
and U16300 (N_16300,N_16245,N_16207);
nand U16301 (N_16301,N_16103,N_16175);
or U16302 (N_16302,N_16056,N_16142);
nor U16303 (N_16303,N_16149,N_16007);
nor U16304 (N_16304,N_16181,N_16087);
and U16305 (N_16305,N_16237,N_16151);
nor U16306 (N_16306,N_16046,N_16225);
nand U16307 (N_16307,N_16164,N_16161);
nor U16308 (N_16308,N_16002,N_16027);
xor U16309 (N_16309,N_16031,N_16093);
and U16310 (N_16310,N_16205,N_16197);
nand U16311 (N_16311,N_16201,N_16147);
nor U16312 (N_16312,N_16247,N_16096);
and U16313 (N_16313,N_16158,N_16241);
nand U16314 (N_16314,N_16016,N_16141);
or U16315 (N_16315,N_16064,N_16140);
and U16316 (N_16316,N_16047,N_16018);
nor U16317 (N_16317,N_16210,N_16139);
and U16318 (N_16318,N_16155,N_16090);
nand U16319 (N_16319,N_16168,N_16187);
nor U16320 (N_16320,N_16012,N_16242);
or U16321 (N_16321,N_16011,N_16026);
or U16322 (N_16322,N_16076,N_16176);
nand U16323 (N_16323,N_16085,N_16101);
nor U16324 (N_16324,N_16145,N_16024);
nor U16325 (N_16325,N_16218,N_16111);
nand U16326 (N_16326,N_16163,N_16115);
nor U16327 (N_16327,N_16069,N_16102);
xor U16328 (N_16328,N_16032,N_16050);
or U16329 (N_16329,N_16243,N_16005);
nor U16330 (N_16330,N_16042,N_16217);
nand U16331 (N_16331,N_16214,N_16099);
xnor U16332 (N_16332,N_16004,N_16157);
nor U16333 (N_16333,N_16062,N_16120);
nand U16334 (N_16334,N_16156,N_16249);
nand U16335 (N_16335,N_16098,N_16077);
or U16336 (N_16336,N_16075,N_16169);
nor U16337 (N_16337,N_16190,N_16119);
nand U16338 (N_16338,N_16234,N_16055);
nand U16339 (N_16339,N_16044,N_16079);
nor U16340 (N_16340,N_16105,N_16221);
nor U16341 (N_16341,N_16083,N_16213);
and U16342 (N_16342,N_16109,N_16125);
or U16343 (N_16343,N_16244,N_16059);
or U16344 (N_16344,N_16159,N_16195);
nand U16345 (N_16345,N_16022,N_16230);
and U16346 (N_16346,N_16092,N_16058);
or U16347 (N_16347,N_16208,N_16219);
or U16348 (N_16348,N_16104,N_16084);
and U16349 (N_16349,N_16131,N_16094);
and U16350 (N_16350,N_16065,N_16223);
nor U16351 (N_16351,N_16074,N_16006);
nand U16352 (N_16352,N_16165,N_16229);
nor U16353 (N_16353,N_16071,N_16054);
or U16354 (N_16354,N_16235,N_16034);
nor U16355 (N_16355,N_16095,N_16116);
and U16356 (N_16356,N_16185,N_16049);
nand U16357 (N_16357,N_16174,N_16152);
nor U16358 (N_16358,N_16135,N_16126);
or U16359 (N_16359,N_16000,N_16001);
nor U16360 (N_16360,N_16108,N_16199);
or U16361 (N_16361,N_16202,N_16112);
nand U16362 (N_16362,N_16153,N_16003);
nor U16363 (N_16363,N_16188,N_16196);
nand U16364 (N_16364,N_16040,N_16107);
or U16365 (N_16365,N_16033,N_16052);
nor U16366 (N_16366,N_16206,N_16134);
nand U16367 (N_16367,N_16106,N_16146);
nor U16368 (N_16368,N_16122,N_16228);
or U16369 (N_16369,N_16036,N_16227);
nor U16370 (N_16370,N_16150,N_16162);
nand U16371 (N_16371,N_16239,N_16080);
and U16372 (N_16372,N_16133,N_16009);
nand U16373 (N_16373,N_16200,N_16118);
xnor U16374 (N_16374,N_16030,N_16130);
nand U16375 (N_16375,N_16123,N_16127);
xor U16376 (N_16376,N_16134,N_16028);
nor U16377 (N_16377,N_16150,N_16202);
nor U16378 (N_16378,N_16205,N_16121);
nand U16379 (N_16379,N_16133,N_16194);
nand U16380 (N_16380,N_16183,N_16139);
nand U16381 (N_16381,N_16043,N_16042);
or U16382 (N_16382,N_16175,N_16006);
nor U16383 (N_16383,N_16179,N_16000);
and U16384 (N_16384,N_16183,N_16227);
and U16385 (N_16385,N_16151,N_16170);
nor U16386 (N_16386,N_16087,N_16224);
nand U16387 (N_16387,N_16198,N_16062);
nor U16388 (N_16388,N_16188,N_16095);
xnor U16389 (N_16389,N_16172,N_16109);
nor U16390 (N_16390,N_16184,N_16032);
and U16391 (N_16391,N_16023,N_16242);
and U16392 (N_16392,N_16060,N_16103);
nand U16393 (N_16393,N_16081,N_16016);
nand U16394 (N_16394,N_16078,N_16071);
or U16395 (N_16395,N_16064,N_16187);
and U16396 (N_16396,N_16234,N_16153);
nor U16397 (N_16397,N_16229,N_16120);
or U16398 (N_16398,N_16131,N_16133);
or U16399 (N_16399,N_16083,N_16155);
nand U16400 (N_16400,N_16100,N_16178);
and U16401 (N_16401,N_16020,N_16173);
and U16402 (N_16402,N_16106,N_16247);
nand U16403 (N_16403,N_16132,N_16151);
nor U16404 (N_16404,N_16018,N_16010);
nand U16405 (N_16405,N_16005,N_16212);
and U16406 (N_16406,N_16132,N_16233);
xnor U16407 (N_16407,N_16065,N_16056);
and U16408 (N_16408,N_16173,N_16117);
nand U16409 (N_16409,N_16082,N_16201);
xor U16410 (N_16410,N_16213,N_16167);
nand U16411 (N_16411,N_16152,N_16020);
nor U16412 (N_16412,N_16118,N_16020);
xor U16413 (N_16413,N_16000,N_16023);
and U16414 (N_16414,N_16142,N_16162);
and U16415 (N_16415,N_16081,N_16213);
xnor U16416 (N_16416,N_16131,N_16150);
nor U16417 (N_16417,N_16154,N_16167);
nand U16418 (N_16418,N_16093,N_16197);
xnor U16419 (N_16419,N_16003,N_16135);
xnor U16420 (N_16420,N_16194,N_16135);
and U16421 (N_16421,N_16235,N_16039);
nand U16422 (N_16422,N_16116,N_16010);
nand U16423 (N_16423,N_16113,N_16006);
xnor U16424 (N_16424,N_16101,N_16089);
or U16425 (N_16425,N_16210,N_16203);
or U16426 (N_16426,N_16006,N_16249);
or U16427 (N_16427,N_16106,N_16026);
nor U16428 (N_16428,N_16191,N_16195);
or U16429 (N_16429,N_16097,N_16199);
nand U16430 (N_16430,N_16154,N_16119);
xnor U16431 (N_16431,N_16035,N_16187);
or U16432 (N_16432,N_16050,N_16174);
nor U16433 (N_16433,N_16104,N_16235);
nand U16434 (N_16434,N_16200,N_16158);
xor U16435 (N_16435,N_16003,N_16198);
nand U16436 (N_16436,N_16227,N_16046);
nand U16437 (N_16437,N_16154,N_16135);
xnor U16438 (N_16438,N_16022,N_16181);
and U16439 (N_16439,N_16247,N_16075);
and U16440 (N_16440,N_16037,N_16141);
xnor U16441 (N_16441,N_16178,N_16018);
nand U16442 (N_16442,N_16242,N_16047);
or U16443 (N_16443,N_16230,N_16109);
or U16444 (N_16444,N_16018,N_16162);
xnor U16445 (N_16445,N_16020,N_16099);
or U16446 (N_16446,N_16056,N_16072);
and U16447 (N_16447,N_16153,N_16112);
xor U16448 (N_16448,N_16153,N_16064);
and U16449 (N_16449,N_16158,N_16056);
nor U16450 (N_16450,N_16100,N_16047);
nor U16451 (N_16451,N_16076,N_16248);
nor U16452 (N_16452,N_16207,N_16248);
or U16453 (N_16453,N_16162,N_16079);
or U16454 (N_16454,N_16086,N_16135);
nand U16455 (N_16455,N_16099,N_16041);
nand U16456 (N_16456,N_16182,N_16157);
xor U16457 (N_16457,N_16187,N_16241);
and U16458 (N_16458,N_16063,N_16067);
or U16459 (N_16459,N_16097,N_16168);
or U16460 (N_16460,N_16082,N_16212);
nor U16461 (N_16461,N_16161,N_16024);
nand U16462 (N_16462,N_16085,N_16182);
nor U16463 (N_16463,N_16178,N_16190);
xnor U16464 (N_16464,N_16207,N_16177);
and U16465 (N_16465,N_16242,N_16111);
nand U16466 (N_16466,N_16118,N_16000);
nor U16467 (N_16467,N_16245,N_16124);
or U16468 (N_16468,N_16196,N_16084);
or U16469 (N_16469,N_16062,N_16100);
nor U16470 (N_16470,N_16083,N_16196);
or U16471 (N_16471,N_16178,N_16036);
or U16472 (N_16472,N_16033,N_16187);
nor U16473 (N_16473,N_16088,N_16125);
or U16474 (N_16474,N_16169,N_16034);
nand U16475 (N_16475,N_16106,N_16214);
or U16476 (N_16476,N_16176,N_16208);
nand U16477 (N_16477,N_16245,N_16017);
nor U16478 (N_16478,N_16052,N_16170);
and U16479 (N_16479,N_16150,N_16058);
nor U16480 (N_16480,N_16233,N_16112);
nand U16481 (N_16481,N_16124,N_16023);
nand U16482 (N_16482,N_16171,N_16158);
and U16483 (N_16483,N_16013,N_16154);
nor U16484 (N_16484,N_16241,N_16156);
nand U16485 (N_16485,N_16064,N_16041);
or U16486 (N_16486,N_16206,N_16223);
or U16487 (N_16487,N_16220,N_16088);
or U16488 (N_16488,N_16126,N_16210);
or U16489 (N_16489,N_16144,N_16200);
xor U16490 (N_16490,N_16164,N_16094);
nor U16491 (N_16491,N_16077,N_16194);
and U16492 (N_16492,N_16175,N_16245);
nor U16493 (N_16493,N_16139,N_16182);
and U16494 (N_16494,N_16061,N_16221);
nand U16495 (N_16495,N_16225,N_16174);
and U16496 (N_16496,N_16095,N_16072);
xor U16497 (N_16497,N_16216,N_16238);
and U16498 (N_16498,N_16112,N_16209);
or U16499 (N_16499,N_16037,N_16015);
nand U16500 (N_16500,N_16303,N_16336);
and U16501 (N_16501,N_16350,N_16255);
nor U16502 (N_16502,N_16429,N_16483);
or U16503 (N_16503,N_16289,N_16369);
and U16504 (N_16504,N_16436,N_16494);
or U16505 (N_16505,N_16444,N_16320);
nor U16506 (N_16506,N_16394,N_16437);
or U16507 (N_16507,N_16312,N_16277);
or U16508 (N_16508,N_16364,N_16391);
nand U16509 (N_16509,N_16270,N_16259);
nor U16510 (N_16510,N_16254,N_16251);
and U16511 (N_16511,N_16304,N_16380);
and U16512 (N_16512,N_16454,N_16296);
and U16513 (N_16513,N_16461,N_16498);
nor U16514 (N_16514,N_16458,N_16333);
or U16515 (N_16515,N_16319,N_16478);
nand U16516 (N_16516,N_16393,N_16323);
nand U16517 (N_16517,N_16311,N_16362);
or U16518 (N_16518,N_16385,N_16479);
xor U16519 (N_16519,N_16432,N_16463);
nand U16520 (N_16520,N_16347,N_16353);
nor U16521 (N_16521,N_16417,N_16400);
nand U16522 (N_16522,N_16337,N_16398);
nor U16523 (N_16523,N_16370,N_16274);
and U16524 (N_16524,N_16467,N_16309);
and U16525 (N_16525,N_16314,N_16407);
nor U16526 (N_16526,N_16420,N_16491);
nand U16527 (N_16527,N_16342,N_16470);
or U16528 (N_16528,N_16443,N_16451);
nand U16529 (N_16529,N_16327,N_16334);
and U16530 (N_16530,N_16381,N_16424);
nor U16531 (N_16531,N_16371,N_16448);
and U16532 (N_16532,N_16452,N_16344);
nor U16533 (N_16533,N_16408,N_16335);
nand U16534 (N_16534,N_16267,N_16495);
xor U16535 (N_16535,N_16261,N_16425);
nand U16536 (N_16536,N_16300,N_16285);
nand U16537 (N_16537,N_16378,N_16410);
nor U16538 (N_16538,N_16477,N_16271);
or U16539 (N_16539,N_16307,N_16315);
nor U16540 (N_16540,N_16288,N_16262);
and U16541 (N_16541,N_16366,N_16442);
nand U16542 (N_16542,N_16357,N_16340);
nand U16543 (N_16543,N_16313,N_16496);
nor U16544 (N_16544,N_16439,N_16283);
nor U16545 (N_16545,N_16422,N_16459);
or U16546 (N_16546,N_16302,N_16490);
nor U16547 (N_16547,N_16409,N_16317);
xnor U16548 (N_16548,N_16310,N_16373);
or U16549 (N_16549,N_16419,N_16338);
nand U16550 (N_16550,N_16469,N_16292);
nor U16551 (N_16551,N_16430,N_16272);
nand U16552 (N_16552,N_16497,N_16301);
nand U16553 (N_16553,N_16428,N_16284);
or U16554 (N_16554,N_16265,N_16395);
and U16555 (N_16555,N_16476,N_16396);
and U16556 (N_16556,N_16368,N_16389);
and U16557 (N_16557,N_16305,N_16298);
xnor U16558 (N_16558,N_16355,N_16471);
xnor U16559 (N_16559,N_16325,N_16457);
nor U16560 (N_16560,N_16482,N_16372);
and U16561 (N_16561,N_16418,N_16299);
nand U16562 (N_16562,N_16433,N_16485);
xnor U16563 (N_16563,N_16308,N_16435);
nor U16564 (N_16564,N_16331,N_16268);
xnor U16565 (N_16565,N_16266,N_16354);
nand U16566 (N_16566,N_16447,N_16499);
nand U16567 (N_16567,N_16421,N_16453);
nor U16568 (N_16568,N_16392,N_16413);
or U16569 (N_16569,N_16423,N_16412);
and U16570 (N_16570,N_16460,N_16363);
nor U16571 (N_16571,N_16466,N_16359);
nand U16572 (N_16572,N_16273,N_16352);
and U16573 (N_16573,N_16358,N_16434);
and U16574 (N_16574,N_16402,N_16322);
nand U16575 (N_16575,N_16411,N_16275);
nand U16576 (N_16576,N_16374,N_16360);
nand U16577 (N_16577,N_16329,N_16427);
or U16578 (N_16578,N_16257,N_16446);
or U16579 (N_16579,N_16328,N_16252);
nand U16580 (N_16580,N_16324,N_16449);
and U16581 (N_16581,N_16339,N_16450);
nand U16582 (N_16582,N_16397,N_16474);
and U16583 (N_16583,N_16464,N_16287);
nand U16584 (N_16584,N_16367,N_16383);
or U16585 (N_16585,N_16440,N_16390);
or U16586 (N_16586,N_16375,N_16330);
or U16587 (N_16587,N_16297,N_16462);
and U16588 (N_16588,N_16404,N_16293);
or U16589 (N_16589,N_16455,N_16486);
or U16590 (N_16590,N_16492,N_16406);
or U16591 (N_16591,N_16441,N_16332);
nand U16592 (N_16592,N_16489,N_16269);
nand U16593 (N_16593,N_16253,N_16351);
nor U16594 (N_16594,N_16260,N_16263);
nand U16595 (N_16595,N_16356,N_16405);
or U16596 (N_16596,N_16286,N_16276);
nand U16597 (N_16597,N_16401,N_16426);
xnor U16598 (N_16598,N_16488,N_16365);
nand U16599 (N_16599,N_16377,N_16388);
and U16600 (N_16600,N_16291,N_16321);
nor U16601 (N_16601,N_16399,N_16493);
nand U16602 (N_16602,N_16487,N_16465);
nor U16603 (N_16603,N_16475,N_16403);
or U16604 (N_16604,N_16258,N_16387);
nor U16605 (N_16605,N_16468,N_16415);
nor U16606 (N_16606,N_16414,N_16326);
or U16607 (N_16607,N_16318,N_16294);
and U16608 (N_16608,N_16438,N_16278);
or U16609 (N_16609,N_16316,N_16345);
xor U16610 (N_16610,N_16376,N_16382);
nand U16611 (N_16611,N_16250,N_16343);
nand U16612 (N_16612,N_16264,N_16456);
nor U16613 (N_16613,N_16282,N_16481);
nand U16614 (N_16614,N_16346,N_16431);
nand U16615 (N_16615,N_16256,N_16280);
or U16616 (N_16616,N_16341,N_16295);
nand U16617 (N_16617,N_16473,N_16484);
nor U16618 (N_16618,N_16379,N_16349);
nor U16619 (N_16619,N_16480,N_16281);
nor U16620 (N_16620,N_16386,N_16416);
xnor U16621 (N_16621,N_16384,N_16348);
and U16622 (N_16622,N_16279,N_16306);
xor U16623 (N_16623,N_16290,N_16445);
and U16624 (N_16624,N_16472,N_16361);
and U16625 (N_16625,N_16328,N_16416);
nor U16626 (N_16626,N_16491,N_16481);
and U16627 (N_16627,N_16489,N_16268);
nand U16628 (N_16628,N_16385,N_16478);
nor U16629 (N_16629,N_16255,N_16285);
and U16630 (N_16630,N_16358,N_16491);
xor U16631 (N_16631,N_16316,N_16335);
xor U16632 (N_16632,N_16380,N_16469);
or U16633 (N_16633,N_16440,N_16250);
nor U16634 (N_16634,N_16461,N_16323);
and U16635 (N_16635,N_16445,N_16256);
and U16636 (N_16636,N_16398,N_16264);
or U16637 (N_16637,N_16280,N_16329);
and U16638 (N_16638,N_16317,N_16418);
nor U16639 (N_16639,N_16274,N_16254);
nor U16640 (N_16640,N_16377,N_16428);
or U16641 (N_16641,N_16318,N_16426);
nor U16642 (N_16642,N_16253,N_16271);
and U16643 (N_16643,N_16319,N_16371);
nand U16644 (N_16644,N_16459,N_16409);
or U16645 (N_16645,N_16299,N_16304);
nand U16646 (N_16646,N_16348,N_16426);
or U16647 (N_16647,N_16428,N_16322);
nand U16648 (N_16648,N_16302,N_16479);
or U16649 (N_16649,N_16350,N_16304);
nor U16650 (N_16650,N_16372,N_16301);
and U16651 (N_16651,N_16396,N_16288);
and U16652 (N_16652,N_16430,N_16448);
nor U16653 (N_16653,N_16347,N_16437);
nor U16654 (N_16654,N_16375,N_16441);
or U16655 (N_16655,N_16291,N_16354);
or U16656 (N_16656,N_16291,N_16477);
or U16657 (N_16657,N_16342,N_16434);
nor U16658 (N_16658,N_16406,N_16421);
nor U16659 (N_16659,N_16331,N_16320);
nand U16660 (N_16660,N_16450,N_16491);
nor U16661 (N_16661,N_16334,N_16378);
nand U16662 (N_16662,N_16286,N_16336);
nand U16663 (N_16663,N_16375,N_16357);
nand U16664 (N_16664,N_16494,N_16373);
or U16665 (N_16665,N_16476,N_16266);
or U16666 (N_16666,N_16482,N_16307);
nor U16667 (N_16667,N_16325,N_16296);
and U16668 (N_16668,N_16450,N_16272);
nor U16669 (N_16669,N_16269,N_16480);
or U16670 (N_16670,N_16489,N_16301);
or U16671 (N_16671,N_16417,N_16496);
nor U16672 (N_16672,N_16417,N_16456);
nand U16673 (N_16673,N_16423,N_16474);
nand U16674 (N_16674,N_16413,N_16486);
nor U16675 (N_16675,N_16363,N_16395);
nand U16676 (N_16676,N_16440,N_16376);
and U16677 (N_16677,N_16340,N_16450);
nand U16678 (N_16678,N_16284,N_16491);
nor U16679 (N_16679,N_16286,N_16250);
nor U16680 (N_16680,N_16423,N_16364);
nor U16681 (N_16681,N_16388,N_16283);
nand U16682 (N_16682,N_16371,N_16351);
or U16683 (N_16683,N_16267,N_16367);
and U16684 (N_16684,N_16397,N_16268);
nand U16685 (N_16685,N_16471,N_16311);
nor U16686 (N_16686,N_16369,N_16290);
xor U16687 (N_16687,N_16347,N_16406);
nand U16688 (N_16688,N_16457,N_16470);
and U16689 (N_16689,N_16354,N_16393);
nor U16690 (N_16690,N_16270,N_16367);
nor U16691 (N_16691,N_16303,N_16389);
and U16692 (N_16692,N_16420,N_16366);
nor U16693 (N_16693,N_16497,N_16289);
or U16694 (N_16694,N_16467,N_16325);
and U16695 (N_16695,N_16258,N_16353);
and U16696 (N_16696,N_16311,N_16450);
nor U16697 (N_16697,N_16340,N_16333);
and U16698 (N_16698,N_16491,N_16374);
and U16699 (N_16699,N_16416,N_16271);
nand U16700 (N_16700,N_16336,N_16419);
nor U16701 (N_16701,N_16499,N_16483);
and U16702 (N_16702,N_16351,N_16470);
nand U16703 (N_16703,N_16332,N_16267);
or U16704 (N_16704,N_16259,N_16257);
or U16705 (N_16705,N_16355,N_16262);
and U16706 (N_16706,N_16311,N_16374);
nand U16707 (N_16707,N_16486,N_16482);
nand U16708 (N_16708,N_16449,N_16488);
and U16709 (N_16709,N_16301,N_16463);
xor U16710 (N_16710,N_16477,N_16318);
and U16711 (N_16711,N_16433,N_16342);
or U16712 (N_16712,N_16375,N_16442);
or U16713 (N_16713,N_16381,N_16380);
and U16714 (N_16714,N_16441,N_16488);
nand U16715 (N_16715,N_16472,N_16363);
nand U16716 (N_16716,N_16361,N_16436);
nor U16717 (N_16717,N_16454,N_16494);
xnor U16718 (N_16718,N_16309,N_16337);
or U16719 (N_16719,N_16271,N_16380);
nand U16720 (N_16720,N_16367,N_16454);
nor U16721 (N_16721,N_16348,N_16290);
or U16722 (N_16722,N_16329,N_16271);
and U16723 (N_16723,N_16338,N_16300);
or U16724 (N_16724,N_16491,N_16381);
or U16725 (N_16725,N_16296,N_16321);
nand U16726 (N_16726,N_16424,N_16416);
xor U16727 (N_16727,N_16482,N_16444);
nand U16728 (N_16728,N_16319,N_16424);
nor U16729 (N_16729,N_16383,N_16462);
or U16730 (N_16730,N_16396,N_16434);
or U16731 (N_16731,N_16295,N_16317);
nor U16732 (N_16732,N_16403,N_16258);
or U16733 (N_16733,N_16300,N_16251);
nand U16734 (N_16734,N_16377,N_16253);
or U16735 (N_16735,N_16333,N_16400);
nand U16736 (N_16736,N_16471,N_16365);
and U16737 (N_16737,N_16374,N_16283);
and U16738 (N_16738,N_16441,N_16381);
nor U16739 (N_16739,N_16296,N_16405);
nor U16740 (N_16740,N_16432,N_16434);
or U16741 (N_16741,N_16410,N_16416);
or U16742 (N_16742,N_16252,N_16383);
nand U16743 (N_16743,N_16461,N_16497);
xnor U16744 (N_16744,N_16332,N_16389);
nand U16745 (N_16745,N_16437,N_16378);
or U16746 (N_16746,N_16487,N_16264);
and U16747 (N_16747,N_16377,N_16305);
xnor U16748 (N_16748,N_16337,N_16325);
and U16749 (N_16749,N_16369,N_16467);
or U16750 (N_16750,N_16615,N_16707);
nand U16751 (N_16751,N_16632,N_16540);
nor U16752 (N_16752,N_16613,N_16538);
or U16753 (N_16753,N_16746,N_16587);
or U16754 (N_16754,N_16590,N_16607);
and U16755 (N_16755,N_16649,N_16554);
nand U16756 (N_16756,N_16627,N_16702);
or U16757 (N_16757,N_16659,N_16548);
and U16758 (N_16758,N_16528,N_16695);
or U16759 (N_16759,N_16550,N_16551);
or U16760 (N_16760,N_16720,N_16749);
nor U16761 (N_16761,N_16565,N_16737);
or U16762 (N_16762,N_16648,N_16501);
and U16763 (N_16763,N_16748,N_16559);
nor U16764 (N_16764,N_16512,N_16709);
nand U16765 (N_16765,N_16608,N_16732);
and U16766 (N_16766,N_16623,N_16686);
nor U16767 (N_16767,N_16500,N_16730);
or U16768 (N_16768,N_16536,N_16561);
or U16769 (N_16769,N_16638,N_16566);
nor U16770 (N_16770,N_16517,N_16696);
nand U16771 (N_16771,N_16634,N_16541);
nor U16772 (N_16772,N_16666,N_16604);
and U16773 (N_16773,N_16745,N_16593);
nand U16774 (N_16774,N_16653,N_16673);
and U16775 (N_16775,N_16739,N_16681);
nor U16776 (N_16776,N_16645,N_16506);
or U16777 (N_16777,N_16513,N_16526);
nor U16778 (N_16778,N_16585,N_16642);
and U16779 (N_16779,N_16625,N_16520);
and U16780 (N_16780,N_16650,N_16669);
or U16781 (N_16781,N_16522,N_16651);
nor U16782 (N_16782,N_16605,N_16719);
or U16783 (N_16783,N_16524,N_16738);
nor U16784 (N_16784,N_16609,N_16602);
or U16785 (N_16785,N_16519,N_16544);
or U16786 (N_16786,N_16597,N_16722);
nand U16787 (N_16787,N_16622,N_16711);
nor U16788 (N_16788,N_16510,N_16578);
nand U16789 (N_16789,N_16654,N_16743);
or U16790 (N_16790,N_16619,N_16674);
nor U16791 (N_16791,N_16714,N_16700);
or U16792 (N_16792,N_16682,N_16708);
or U16793 (N_16793,N_16598,N_16736);
nand U16794 (N_16794,N_16539,N_16533);
or U16795 (N_16795,N_16564,N_16571);
nand U16796 (N_16796,N_16557,N_16701);
and U16797 (N_16797,N_16637,N_16610);
or U16798 (N_16798,N_16592,N_16555);
and U16799 (N_16799,N_16705,N_16588);
or U16800 (N_16800,N_16663,N_16572);
and U16801 (N_16801,N_16710,N_16567);
nor U16802 (N_16802,N_16546,N_16727);
and U16803 (N_16803,N_16694,N_16547);
nand U16804 (N_16804,N_16678,N_16630);
and U16805 (N_16805,N_16715,N_16503);
xor U16806 (N_16806,N_16689,N_16685);
nand U16807 (N_16807,N_16661,N_16516);
or U16808 (N_16808,N_16677,N_16680);
or U16809 (N_16809,N_16635,N_16633);
nand U16810 (N_16810,N_16583,N_16672);
nor U16811 (N_16811,N_16644,N_16570);
or U16812 (N_16812,N_16591,N_16553);
or U16813 (N_16813,N_16576,N_16717);
nand U16814 (N_16814,N_16729,N_16636);
nor U16815 (N_16815,N_16667,N_16640);
nor U16816 (N_16816,N_16693,N_16660);
nand U16817 (N_16817,N_16603,N_16525);
or U16818 (N_16818,N_16740,N_16531);
nor U16819 (N_16819,N_16665,N_16628);
nand U16820 (N_16820,N_16586,N_16684);
nand U16821 (N_16821,N_16574,N_16600);
and U16822 (N_16822,N_16725,N_16699);
nor U16823 (N_16823,N_16620,N_16691);
or U16824 (N_16824,N_16690,N_16545);
nor U16825 (N_16825,N_16573,N_16664);
and U16826 (N_16826,N_16534,N_16502);
nor U16827 (N_16827,N_16558,N_16601);
nor U16828 (N_16828,N_16703,N_16529);
nor U16829 (N_16829,N_16584,N_16569);
nor U16830 (N_16830,N_16514,N_16643);
xnor U16831 (N_16831,N_16560,N_16579);
xor U16832 (N_16832,N_16655,N_16589);
or U16833 (N_16833,N_16543,N_16647);
nor U16834 (N_16834,N_16624,N_16641);
or U16835 (N_16835,N_16713,N_16712);
xor U16836 (N_16836,N_16537,N_16679);
nand U16837 (N_16837,N_16671,N_16568);
nand U16838 (N_16838,N_16532,N_16563);
and U16839 (N_16839,N_16515,N_16611);
nand U16840 (N_16840,N_16616,N_16508);
and U16841 (N_16841,N_16704,N_16658);
nand U16842 (N_16842,N_16698,N_16511);
or U16843 (N_16843,N_16744,N_16724);
nand U16844 (N_16844,N_16580,N_16716);
nor U16845 (N_16845,N_16676,N_16728);
xor U16846 (N_16846,N_16523,N_16646);
and U16847 (N_16847,N_16507,N_16639);
xor U16848 (N_16848,N_16521,N_16656);
or U16849 (N_16849,N_16505,N_16733);
or U16850 (N_16850,N_16683,N_16509);
or U16851 (N_16851,N_16617,N_16629);
and U16852 (N_16852,N_16599,N_16631);
nor U16853 (N_16853,N_16552,N_16535);
nor U16854 (N_16854,N_16612,N_16542);
and U16855 (N_16855,N_16562,N_16596);
nand U16856 (N_16856,N_16626,N_16575);
xnor U16857 (N_16857,N_16581,N_16726);
nand U16858 (N_16858,N_16731,N_16668);
nor U16859 (N_16859,N_16530,N_16556);
or U16860 (N_16860,N_16652,N_16692);
nor U16861 (N_16861,N_16582,N_16577);
nand U16862 (N_16862,N_16747,N_16706);
nand U16863 (N_16863,N_16742,N_16618);
and U16864 (N_16864,N_16527,N_16687);
nand U16865 (N_16865,N_16614,N_16734);
nand U16866 (N_16866,N_16735,N_16504);
xnor U16867 (N_16867,N_16621,N_16594);
nand U16868 (N_16868,N_16721,N_16595);
xnor U16869 (N_16869,N_16518,N_16670);
xor U16870 (N_16870,N_16723,N_16662);
nor U16871 (N_16871,N_16741,N_16697);
or U16872 (N_16872,N_16549,N_16675);
and U16873 (N_16873,N_16718,N_16606);
xor U16874 (N_16874,N_16688,N_16657);
nor U16875 (N_16875,N_16511,N_16650);
nor U16876 (N_16876,N_16651,N_16626);
and U16877 (N_16877,N_16702,N_16531);
nand U16878 (N_16878,N_16548,N_16654);
or U16879 (N_16879,N_16507,N_16733);
and U16880 (N_16880,N_16506,N_16722);
and U16881 (N_16881,N_16680,N_16529);
nand U16882 (N_16882,N_16506,N_16511);
and U16883 (N_16883,N_16525,N_16516);
nor U16884 (N_16884,N_16667,N_16720);
or U16885 (N_16885,N_16547,N_16685);
or U16886 (N_16886,N_16694,N_16731);
and U16887 (N_16887,N_16504,N_16633);
or U16888 (N_16888,N_16674,N_16546);
or U16889 (N_16889,N_16655,N_16553);
nand U16890 (N_16890,N_16715,N_16727);
nor U16891 (N_16891,N_16559,N_16547);
or U16892 (N_16892,N_16520,N_16600);
xor U16893 (N_16893,N_16567,N_16614);
and U16894 (N_16894,N_16702,N_16592);
and U16895 (N_16895,N_16718,N_16705);
nand U16896 (N_16896,N_16676,N_16649);
nor U16897 (N_16897,N_16579,N_16653);
or U16898 (N_16898,N_16570,N_16660);
nand U16899 (N_16899,N_16726,N_16588);
and U16900 (N_16900,N_16618,N_16587);
nand U16901 (N_16901,N_16735,N_16621);
nand U16902 (N_16902,N_16576,N_16515);
nor U16903 (N_16903,N_16624,N_16734);
nor U16904 (N_16904,N_16669,N_16685);
nor U16905 (N_16905,N_16538,N_16690);
or U16906 (N_16906,N_16745,N_16571);
nand U16907 (N_16907,N_16552,N_16532);
nand U16908 (N_16908,N_16740,N_16558);
xor U16909 (N_16909,N_16587,N_16528);
or U16910 (N_16910,N_16681,N_16636);
xor U16911 (N_16911,N_16609,N_16695);
or U16912 (N_16912,N_16548,N_16611);
or U16913 (N_16913,N_16523,N_16662);
nand U16914 (N_16914,N_16534,N_16582);
nor U16915 (N_16915,N_16518,N_16506);
or U16916 (N_16916,N_16528,N_16568);
and U16917 (N_16917,N_16587,N_16743);
nor U16918 (N_16918,N_16702,N_16551);
xor U16919 (N_16919,N_16615,N_16672);
and U16920 (N_16920,N_16561,N_16681);
or U16921 (N_16921,N_16678,N_16655);
and U16922 (N_16922,N_16737,N_16726);
xnor U16923 (N_16923,N_16595,N_16740);
nand U16924 (N_16924,N_16547,N_16633);
nand U16925 (N_16925,N_16522,N_16605);
and U16926 (N_16926,N_16688,N_16604);
nor U16927 (N_16927,N_16658,N_16606);
xor U16928 (N_16928,N_16720,N_16693);
nand U16929 (N_16929,N_16536,N_16553);
nor U16930 (N_16930,N_16523,N_16621);
or U16931 (N_16931,N_16513,N_16609);
and U16932 (N_16932,N_16700,N_16609);
xor U16933 (N_16933,N_16575,N_16609);
nor U16934 (N_16934,N_16588,N_16659);
nand U16935 (N_16935,N_16691,N_16745);
or U16936 (N_16936,N_16537,N_16733);
or U16937 (N_16937,N_16581,N_16576);
nand U16938 (N_16938,N_16663,N_16745);
nand U16939 (N_16939,N_16524,N_16573);
and U16940 (N_16940,N_16519,N_16570);
nor U16941 (N_16941,N_16509,N_16638);
nand U16942 (N_16942,N_16549,N_16699);
nand U16943 (N_16943,N_16602,N_16627);
or U16944 (N_16944,N_16666,N_16590);
nor U16945 (N_16945,N_16707,N_16685);
and U16946 (N_16946,N_16629,N_16642);
or U16947 (N_16947,N_16628,N_16652);
or U16948 (N_16948,N_16668,N_16656);
nor U16949 (N_16949,N_16519,N_16640);
nor U16950 (N_16950,N_16590,N_16697);
and U16951 (N_16951,N_16635,N_16690);
or U16952 (N_16952,N_16699,N_16505);
nand U16953 (N_16953,N_16569,N_16596);
xnor U16954 (N_16954,N_16729,N_16589);
nand U16955 (N_16955,N_16576,N_16742);
nand U16956 (N_16956,N_16558,N_16543);
nor U16957 (N_16957,N_16517,N_16744);
and U16958 (N_16958,N_16557,N_16726);
nor U16959 (N_16959,N_16508,N_16668);
and U16960 (N_16960,N_16541,N_16522);
and U16961 (N_16961,N_16657,N_16650);
nand U16962 (N_16962,N_16646,N_16699);
and U16963 (N_16963,N_16649,N_16736);
and U16964 (N_16964,N_16600,N_16646);
or U16965 (N_16965,N_16577,N_16720);
or U16966 (N_16966,N_16641,N_16672);
and U16967 (N_16967,N_16590,N_16525);
or U16968 (N_16968,N_16687,N_16582);
xnor U16969 (N_16969,N_16598,N_16709);
nor U16970 (N_16970,N_16637,N_16574);
or U16971 (N_16971,N_16500,N_16576);
xor U16972 (N_16972,N_16635,N_16663);
nand U16973 (N_16973,N_16697,N_16676);
nand U16974 (N_16974,N_16671,N_16641);
nand U16975 (N_16975,N_16671,N_16575);
or U16976 (N_16976,N_16714,N_16721);
nand U16977 (N_16977,N_16730,N_16707);
or U16978 (N_16978,N_16708,N_16606);
nand U16979 (N_16979,N_16539,N_16591);
or U16980 (N_16980,N_16606,N_16592);
and U16981 (N_16981,N_16550,N_16618);
xor U16982 (N_16982,N_16728,N_16544);
nor U16983 (N_16983,N_16685,N_16505);
xor U16984 (N_16984,N_16725,N_16726);
or U16985 (N_16985,N_16643,N_16517);
or U16986 (N_16986,N_16533,N_16593);
and U16987 (N_16987,N_16603,N_16660);
and U16988 (N_16988,N_16632,N_16551);
nand U16989 (N_16989,N_16569,N_16739);
nor U16990 (N_16990,N_16593,N_16644);
nor U16991 (N_16991,N_16591,N_16608);
nor U16992 (N_16992,N_16674,N_16574);
and U16993 (N_16993,N_16522,N_16711);
and U16994 (N_16994,N_16634,N_16633);
or U16995 (N_16995,N_16747,N_16546);
or U16996 (N_16996,N_16524,N_16584);
nand U16997 (N_16997,N_16685,N_16571);
nand U16998 (N_16998,N_16598,N_16740);
or U16999 (N_16999,N_16520,N_16603);
or U17000 (N_17000,N_16768,N_16885);
nor U17001 (N_17001,N_16819,N_16873);
and U17002 (N_17002,N_16827,N_16944);
and U17003 (N_17003,N_16894,N_16908);
or U17004 (N_17004,N_16915,N_16783);
xor U17005 (N_17005,N_16960,N_16948);
and U17006 (N_17006,N_16881,N_16792);
nand U17007 (N_17007,N_16921,N_16923);
or U17008 (N_17008,N_16765,N_16866);
and U17009 (N_17009,N_16968,N_16935);
and U17010 (N_17010,N_16858,N_16817);
and U17011 (N_17011,N_16869,N_16839);
or U17012 (N_17012,N_16967,N_16891);
or U17013 (N_17013,N_16876,N_16798);
nor U17014 (N_17014,N_16984,N_16912);
and U17015 (N_17015,N_16970,N_16871);
nand U17016 (N_17016,N_16950,N_16842);
nor U17017 (N_17017,N_16867,N_16974);
or U17018 (N_17018,N_16816,N_16977);
nand U17019 (N_17019,N_16895,N_16851);
or U17020 (N_17020,N_16859,N_16820);
nand U17021 (N_17021,N_16870,N_16802);
or U17022 (N_17022,N_16814,N_16933);
nand U17023 (N_17023,N_16770,N_16840);
nor U17024 (N_17024,N_16972,N_16872);
nand U17025 (N_17025,N_16823,N_16826);
nor U17026 (N_17026,N_16793,N_16898);
nor U17027 (N_17027,N_16796,N_16964);
nor U17028 (N_17028,N_16801,N_16957);
or U17029 (N_17029,N_16848,N_16784);
nor U17030 (N_17030,N_16811,N_16996);
and U17031 (N_17031,N_16892,N_16804);
and U17032 (N_17032,N_16767,N_16924);
nor U17033 (N_17033,N_16779,N_16962);
or U17034 (N_17034,N_16799,N_16937);
xnor U17035 (N_17035,N_16963,N_16751);
and U17036 (N_17036,N_16834,N_16874);
and U17037 (N_17037,N_16807,N_16931);
or U17038 (N_17038,N_16907,N_16754);
nand U17039 (N_17039,N_16810,N_16916);
nor U17040 (N_17040,N_16975,N_16791);
nor U17041 (N_17041,N_16868,N_16945);
nand U17042 (N_17042,N_16759,N_16939);
or U17043 (N_17043,N_16919,N_16828);
or U17044 (N_17044,N_16949,N_16986);
nor U17045 (N_17045,N_16806,N_16978);
nor U17046 (N_17046,N_16786,N_16794);
nor U17047 (N_17047,N_16880,N_16890);
and U17048 (N_17048,N_16928,N_16753);
nor U17049 (N_17049,N_16882,N_16929);
or U17050 (N_17050,N_16847,N_16887);
nor U17051 (N_17051,N_16987,N_16833);
or U17052 (N_17052,N_16903,N_16992);
nor U17053 (N_17053,N_16763,N_16854);
nand U17054 (N_17054,N_16989,N_16954);
and U17055 (N_17055,N_16782,N_16941);
nor U17056 (N_17056,N_16965,N_16750);
and U17057 (N_17057,N_16983,N_16875);
or U17058 (N_17058,N_16829,N_16864);
or U17059 (N_17059,N_16818,N_16886);
or U17060 (N_17060,N_16809,N_16857);
nand U17061 (N_17061,N_16926,N_16862);
or U17062 (N_17062,N_16911,N_16961);
and U17063 (N_17063,N_16925,N_16756);
nand U17064 (N_17064,N_16772,N_16774);
xnor U17065 (N_17065,N_16959,N_16952);
and U17066 (N_17066,N_16805,N_16942);
xnor U17067 (N_17067,N_16976,N_16995);
and U17068 (N_17068,N_16990,N_16943);
or U17069 (N_17069,N_16932,N_16877);
nor U17070 (N_17070,N_16896,N_16918);
and U17071 (N_17071,N_16865,N_16758);
or U17072 (N_17072,N_16988,N_16997);
or U17073 (N_17073,N_16955,N_16914);
or U17074 (N_17074,N_16778,N_16755);
nand U17075 (N_17075,N_16897,N_16789);
xnor U17076 (N_17076,N_16856,N_16910);
nand U17077 (N_17077,N_16993,N_16830);
or U17078 (N_17078,N_16902,N_16860);
and U17079 (N_17079,N_16821,N_16940);
and U17080 (N_17080,N_16913,N_16780);
or U17081 (N_17081,N_16953,N_16863);
xor U17082 (N_17082,N_16788,N_16785);
nor U17083 (N_17083,N_16760,N_16832);
and U17084 (N_17084,N_16951,N_16998);
nand U17085 (N_17085,N_16999,N_16822);
and U17086 (N_17086,N_16781,N_16973);
nand U17087 (N_17087,N_16884,N_16812);
xor U17088 (N_17088,N_16800,N_16837);
xor U17089 (N_17089,N_16917,N_16879);
or U17090 (N_17090,N_16927,N_16938);
and U17091 (N_17091,N_16813,N_16775);
nor U17092 (N_17092,N_16849,N_16769);
nand U17093 (N_17093,N_16991,N_16808);
nand U17094 (N_17094,N_16878,N_16994);
nor U17095 (N_17095,N_16900,N_16803);
nor U17096 (N_17096,N_16776,N_16764);
or U17097 (N_17097,N_16982,N_16852);
or U17098 (N_17098,N_16980,N_16883);
nor U17099 (N_17099,N_16845,N_16752);
and U17100 (N_17100,N_16844,N_16850);
nand U17101 (N_17101,N_16787,N_16985);
and U17102 (N_17102,N_16888,N_16936);
and U17103 (N_17103,N_16843,N_16922);
nor U17104 (N_17104,N_16889,N_16761);
xnor U17105 (N_17105,N_16846,N_16906);
or U17106 (N_17106,N_16904,N_16777);
xor U17107 (N_17107,N_16971,N_16909);
and U17108 (N_17108,N_16946,N_16853);
nor U17109 (N_17109,N_16825,N_16947);
xnor U17110 (N_17110,N_16838,N_16893);
and U17111 (N_17111,N_16815,N_16855);
nor U17112 (N_17112,N_16958,N_16797);
and U17113 (N_17113,N_16979,N_16981);
xnor U17114 (N_17114,N_16771,N_16905);
xor U17115 (N_17115,N_16831,N_16930);
and U17116 (N_17116,N_16795,N_16966);
and U17117 (N_17117,N_16901,N_16824);
or U17118 (N_17118,N_16899,N_16934);
nor U17119 (N_17119,N_16762,N_16766);
nor U17120 (N_17120,N_16920,N_16969);
nand U17121 (N_17121,N_16956,N_16773);
nand U17122 (N_17122,N_16841,N_16757);
and U17123 (N_17123,N_16836,N_16861);
nand U17124 (N_17124,N_16790,N_16835);
or U17125 (N_17125,N_16795,N_16910);
nor U17126 (N_17126,N_16811,N_16842);
or U17127 (N_17127,N_16924,N_16799);
or U17128 (N_17128,N_16944,N_16751);
and U17129 (N_17129,N_16988,N_16956);
nor U17130 (N_17130,N_16840,N_16884);
or U17131 (N_17131,N_16805,N_16857);
and U17132 (N_17132,N_16902,N_16839);
nor U17133 (N_17133,N_16830,N_16843);
or U17134 (N_17134,N_16812,N_16892);
nor U17135 (N_17135,N_16950,N_16911);
and U17136 (N_17136,N_16964,N_16923);
xnor U17137 (N_17137,N_16906,N_16947);
or U17138 (N_17138,N_16996,N_16791);
or U17139 (N_17139,N_16839,N_16965);
nand U17140 (N_17140,N_16792,N_16886);
nor U17141 (N_17141,N_16862,N_16826);
and U17142 (N_17142,N_16921,N_16933);
nand U17143 (N_17143,N_16897,N_16800);
nor U17144 (N_17144,N_16763,N_16880);
nor U17145 (N_17145,N_16900,N_16867);
and U17146 (N_17146,N_16822,N_16851);
nor U17147 (N_17147,N_16765,N_16838);
and U17148 (N_17148,N_16828,N_16819);
nand U17149 (N_17149,N_16978,N_16801);
and U17150 (N_17150,N_16859,N_16850);
or U17151 (N_17151,N_16845,N_16968);
or U17152 (N_17152,N_16923,N_16981);
xnor U17153 (N_17153,N_16783,N_16864);
nor U17154 (N_17154,N_16761,N_16770);
or U17155 (N_17155,N_16789,N_16761);
xor U17156 (N_17156,N_16987,N_16755);
and U17157 (N_17157,N_16882,N_16859);
xor U17158 (N_17158,N_16879,N_16961);
nand U17159 (N_17159,N_16986,N_16997);
nor U17160 (N_17160,N_16985,N_16763);
and U17161 (N_17161,N_16817,N_16762);
and U17162 (N_17162,N_16949,N_16974);
xnor U17163 (N_17163,N_16832,N_16891);
nor U17164 (N_17164,N_16846,N_16936);
or U17165 (N_17165,N_16850,N_16987);
or U17166 (N_17166,N_16895,N_16998);
nand U17167 (N_17167,N_16771,N_16825);
nor U17168 (N_17168,N_16769,N_16897);
xor U17169 (N_17169,N_16945,N_16825);
or U17170 (N_17170,N_16821,N_16773);
xnor U17171 (N_17171,N_16803,N_16937);
nor U17172 (N_17172,N_16835,N_16883);
and U17173 (N_17173,N_16804,N_16750);
nand U17174 (N_17174,N_16852,N_16868);
or U17175 (N_17175,N_16996,N_16817);
nand U17176 (N_17176,N_16965,N_16909);
xor U17177 (N_17177,N_16812,N_16814);
nor U17178 (N_17178,N_16901,N_16962);
nor U17179 (N_17179,N_16848,N_16923);
nand U17180 (N_17180,N_16831,N_16760);
and U17181 (N_17181,N_16883,N_16914);
nor U17182 (N_17182,N_16998,N_16833);
nand U17183 (N_17183,N_16989,N_16792);
xor U17184 (N_17184,N_16936,N_16873);
nand U17185 (N_17185,N_16935,N_16794);
and U17186 (N_17186,N_16775,N_16925);
nand U17187 (N_17187,N_16798,N_16804);
nand U17188 (N_17188,N_16898,N_16910);
and U17189 (N_17189,N_16928,N_16825);
nor U17190 (N_17190,N_16826,N_16827);
nand U17191 (N_17191,N_16981,N_16879);
xor U17192 (N_17192,N_16931,N_16933);
or U17193 (N_17193,N_16992,N_16837);
nand U17194 (N_17194,N_16985,N_16931);
nand U17195 (N_17195,N_16893,N_16787);
nor U17196 (N_17196,N_16946,N_16824);
and U17197 (N_17197,N_16903,N_16891);
xor U17198 (N_17198,N_16969,N_16815);
nand U17199 (N_17199,N_16881,N_16798);
or U17200 (N_17200,N_16807,N_16829);
nand U17201 (N_17201,N_16929,N_16911);
nand U17202 (N_17202,N_16958,N_16953);
xnor U17203 (N_17203,N_16807,N_16996);
or U17204 (N_17204,N_16858,N_16930);
nor U17205 (N_17205,N_16807,N_16806);
nand U17206 (N_17206,N_16830,N_16941);
and U17207 (N_17207,N_16868,N_16816);
or U17208 (N_17208,N_16964,N_16762);
and U17209 (N_17209,N_16985,N_16902);
nand U17210 (N_17210,N_16755,N_16932);
or U17211 (N_17211,N_16813,N_16783);
nand U17212 (N_17212,N_16831,N_16853);
nand U17213 (N_17213,N_16804,N_16885);
or U17214 (N_17214,N_16994,N_16818);
nor U17215 (N_17215,N_16830,N_16809);
and U17216 (N_17216,N_16781,N_16815);
and U17217 (N_17217,N_16791,N_16830);
nor U17218 (N_17218,N_16943,N_16878);
xnor U17219 (N_17219,N_16833,N_16919);
or U17220 (N_17220,N_16850,N_16958);
and U17221 (N_17221,N_16802,N_16760);
and U17222 (N_17222,N_16975,N_16755);
and U17223 (N_17223,N_16826,N_16857);
nor U17224 (N_17224,N_16894,N_16848);
or U17225 (N_17225,N_16791,N_16897);
and U17226 (N_17226,N_16805,N_16990);
or U17227 (N_17227,N_16873,N_16834);
and U17228 (N_17228,N_16849,N_16968);
nand U17229 (N_17229,N_16827,N_16753);
or U17230 (N_17230,N_16943,N_16886);
or U17231 (N_17231,N_16777,N_16857);
or U17232 (N_17232,N_16938,N_16869);
nor U17233 (N_17233,N_16753,N_16792);
nand U17234 (N_17234,N_16986,N_16881);
nand U17235 (N_17235,N_16872,N_16771);
nand U17236 (N_17236,N_16952,N_16894);
or U17237 (N_17237,N_16863,N_16801);
or U17238 (N_17238,N_16868,N_16821);
nor U17239 (N_17239,N_16937,N_16941);
nor U17240 (N_17240,N_16931,N_16767);
nor U17241 (N_17241,N_16780,N_16856);
or U17242 (N_17242,N_16979,N_16770);
nand U17243 (N_17243,N_16776,N_16914);
nor U17244 (N_17244,N_16937,N_16887);
or U17245 (N_17245,N_16798,N_16791);
and U17246 (N_17246,N_16997,N_16822);
and U17247 (N_17247,N_16966,N_16865);
and U17248 (N_17248,N_16904,N_16874);
nor U17249 (N_17249,N_16998,N_16859);
or U17250 (N_17250,N_17209,N_17245);
nand U17251 (N_17251,N_17095,N_17240);
or U17252 (N_17252,N_17087,N_17066);
xor U17253 (N_17253,N_17170,N_17041);
and U17254 (N_17254,N_17004,N_17035);
xnor U17255 (N_17255,N_17136,N_17194);
nor U17256 (N_17256,N_17142,N_17201);
and U17257 (N_17257,N_17239,N_17164);
and U17258 (N_17258,N_17060,N_17156);
nand U17259 (N_17259,N_17071,N_17248);
or U17260 (N_17260,N_17040,N_17028);
or U17261 (N_17261,N_17155,N_17097);
xnor U17262 (N_17262,N_17169,N_17161);
xor U17263 (N_17263,N_17183,N_17079);
xnor U17264 (N_17264,N_17176,N_17019);
and U17265 (N_17265,N_17214,N_17243);
or U17266 (N_17266,N_17069,N_17159);
nand U17267 (N_17267,N_17084,N_17190);
nand U17268 (N_17268,N_17249,N_17027);
nor U17269 (N_17269,N_17160,N_17026);
xor U17270 (N_17270,N_17171,N_17064);
or U17271 (N_17271,N_17120,N_17049);
or U17272 (N_17272,N_17085,N_17198);
and U17273 (N_17273,N_17094,N_17032);
or U17274 (N_17274,N_17061,N_17114);
nor U17275 (N_17275,N_17217,N_17130);
or U17276 (N_17276,N_17074,N_17106);
nor U17277 (N_17277,N_17015,N_17024);
or U17278 (N_17278,N_17222,N_17111);
nor U17279 (N_17279,N_17224,N_17012);
nor U17280 (N_17280,N_17047,N_17175);
nor U17281 (N_17281,N_17033,N_17244);
and U17282 (N_17282,N_17105,N_17018);
nor U17283 (N_17283,N_17002,N_17067);
and U17284 (N_17284,N_17126,N_17133);
nor U17285 (N_17285,N_17090,N_17208);
nor U17286 (N_17286,N_17186,N_17148);
nand U17287 (N_17287,N_17059,N_17116);
nor U17288 (N_17288,N_17213,N_17246);
nand U17289 (N_17289,N_17101,N_17221);
xnor U17290 (N_17290,N_17013,N_17187);
nand U17291 (N_17291,N_17141,N_17073);
xnor U17292 (N_17292,N_17167,N_17216);
nor U17293 (N_17293,N_17045,N_17080);
and U17294 (N_17294,N_17072,N_17006);
and U17295 (N_17295,N_17168,N_17088);
or U17296 (N_17296,N_17078,N_17063);
nand U17297 (N_17297,N_17189,N_17247);
or U17298 (N_17298,N_17099,N_17092);
nor U17299 (N_17299,N_17112,N_17234);
nand U17300 (N_17300,N_17134,N_17154);
and U17301 (N_17301,N_17009,N_17124);
or U17302 (N_17302,N_17083,N_17178);
nand U17303 (N_17303,N_17029,N_17044);
nor U17304 (N_17304,N_17196,N_17150);
and U17305 (N_17305,N_17211,N_17203);
and U17306 (N_17306,N_17065,N_17098);
nand U17307 (N_17307,N_17139,N_17162);
and U17308 (N_17308,N_17200,N_17191);
nor U17309 (N_17309,N_17193,N_17192);
nor U17310 (N_17310,N_17146,N_17145);
and U17311 (N_17311,N_17125,N_17242);
and U17312 (N_17312,N_17058,N_17207);
nor U17313 (N_17313,N_17227,N_17199);
nand U17314 (N_17314,N_17157,N_17118);
nor U17315 (N_17315,N_17212,N_17152);
nor U17316 (N_17316,N_17011,N_17108);
nor U17317 (N_17317,N_17131,N_17100);
nor U17318 (N_17318,N_17054,N_17057);
nand U17319 (N_17319,N_17158,N_17025);
nand U17320 (N_17320,N_17021,N_17218);
and U17321 (N_17321,N_17128,N_17204);
nand U17322 (N_17322,N_17149,N_17091);
and U17323 (N_17323,N_17003,N_17153);
nor U17324 (N_17324,N_17031,N_17023);
nand U17325 (N_17325,N_17001,N_17237);
nor U17326 (N_17326,N_17181,N_17219);
nand U17327 (N_17327,N_17037,N_17038);
nand U17328 (N_17328,N_17143,N_17121);
or U17329 (N_17329,N_17166,N_17119);
xnor U17330 (N_17330,N_17104,N_17020);
and U17331 (N_17331,N_17123,N_17205);
nor U17332 (N_17332,N_17117,N_17053);
or U17333 (N_17333,N_17238,N_17180);
and U17334 (N_17334,N_17228,N_17068);
and U17335 (N_17335,N_17113,N_17036);
nor U17336 (N_17336,N_17102,N_17138);
or U17337 (N_17337,N_17109,N_17232);
and U17338 (N_17338,N_17043,N_17052);
or U17339 (N_17339,N_17165,N_17077);
or U17340 (N_17340,N_17140,N_17127);
nand U17341 (N_17341,N_17179,N_17184);
and U17342 (N_17342,N_17030,N_17223);
and U17343 (N_17343,N_17177,N_17051);
nand U17344 (N_17344,N_17229,N_17235);
nand U17345 (N_17345,N_17225,N_17202);
nand U17346 (N_17346,N_17034,N_17107);
and U17347 (N_17347,N_17005,N_17014);
or U17348 (N_17348,N_17210,N_17086);
and U17349 (N_17349,N_17151,N_17132);
nand U17350 (N_17350,N_17185,N_17215);
nand U17351 (N_17351,N_17050,N_17236);
or U17352 (N_17352,N_17076,N_17096);
or U17353 (N_17353,N_17163,N_17046);
or U17354 (N_17354,N_17137,N_17144);
nor U17355 (N_17355,N_17174,N_17093);
or U17356 (N_17356,N_17182,N_17007);
or U17357 (N_17357,N_17241,N_17220);
nor U17358 (N_17358,N_17075,N_17081);
xnor U17359 (N_17359,N_17055,N_17230);
or U17360 (N_17360,N_17197,N_17056);
or U17361 (N_17361,N_17135,N_17226);
nor U17362 (N_17362,N_17089,N_17129);
nor U17363 (N_17363,N_17070,N_17188);
or U17364 (N_17364,N_17206,N_17022);
nand U17365 (N_17365,N_17042,N_17172);
and U17366 (N_17366,N_17195,N_17233);
or U17367 (N_17367,N_17010,N_17231);
or U17368 (N_17368,N_17082,N_17017);
nand U17369 (N_17369,N_17115,N_17039);
or U17370 (N_17370,N_17048,N_17062);
and U17371 (N_17371,N_17008,N_17103);
xnor U17372 (N_17372,N_17110,N_17016);
or U17373 (N_17373,N_17147,N_17122);
or U17374 (N_17374,N_17000,N_17173);
or U17375 (N_17375,N_17127,N_17083);
nand U17376 (N_17376,N_17243,N_17237);
nand U17377 (N_17377,N_17102,N_17171);
or U17378 (N_17378,N_17131,N_17062);
nand U17379 (N_17379,N_17013,N_17181);
nand U17380 (N_17380,N_17225,N_17109);
nand U17381 (N_17381,N_17020,N_17083);
nand U17382 (N_17382,N_17230,N_17236);
nor U17383 (N_17383,N_17236,N_17200);
and U17384 (N_17384,N_17006,N_17066);
nand U17385 (N_17385,N_17026,N_17097);
xnor U17386 (N_17386,N_17178,N_17096);
and U17387 (N_17387,N_17215,N_17127);
nor U17388 (N_17388,N_17075,N_17169);
nand U17389 (N_17389,N_17154,N_17071);
or U17390 (N_17390,N_17112,N_17183);
xnor U17391 (N_17391,N_17089,N_17224);
nor U17392 (N_17392,N_17134,N_17035);
and U17393 (N_17393,N_17143,N_17142);
nand U17394 (N_17394,N_17172,N_17088);
nand U17395 (N_17395,N_17054,N_17242);
or U17396 (N_17396,N_17149,N_17088);
nor U17397 (N_17397,N_17230,N_17023);
and U17398 (N_17398,N_17234,N_17167);
and U17399 (N_17399,N_17209,N_17130);
nand U17400 (N_17400,N_17165,N_17162);
xor U17401 (N_17401,N_17178,N_17051);
nor U17402 (N_17402,N_17005,N_17104);
and U17403 (N_17403,N_17201,N_17117);
and U17404 (N_17404,N_17119,N_17066);
or U17405 (N_17405,N_17020,N_17141);
or U17406 (N_17406,N_17086,N_17050);
or U17407 (N_17407,N_17077,N_17243);
and U17408 (N_17408,N_17172,N_17092);
nand U17409 (N_17409,N_17215,N_17135);
and U17410 (N_17410,N_17199,N_17047);
nor U17411 (N_17411,N_17122,N_17025);
nand U17412 (N_17412,N_17014,N_17194);
and U17413 (N_17413,N_17056,N_17165);
and U17414 (N_17414,N_17122,N_17242);
or U17415 (N_17415,N_17242,N_17009);
nor U17416 (N_17416,N_17097,N_17015);
nand U17417 (N_17417,N_17195,N_17207);
nand U17418 (N_17418,N_17001,N_17216);
or U17419 (N_17419,N_17189,N_17009);
and U17420 (N_17420,N_17133,N_17121);
nand U17421 (N_17421,N_17022,N_17077);
xor U17422 (N_17422,N_17245,N_17041);
nor U17423 (N_17423,N_17072,N_17145);
or U17424 (N_17424,N_17000,N_17229);
or U17425 (N_17425,N_17101,N_17214);
nand U17426 (N_17426,N_17071,N_17061);
and U17427 (N_17427,N_17146,N_17100);
or U17428 (N_17428,N_17247,N_17238);
or U17429 (N_17429,N_17153,N_17088);
nand U17430 (N_17430,N_17039,N_17225);
nor U17431 (N_17431,N_17060,N_17178);
nand U17432 (N_17432,N_17004,N_17037);
nor U17433 (N_17433,N_17037,N_17147);
or U17434 (N_17434,N_17192,N_17088);
nand U17435 (N_17435,N_17073,N_17135);
nor U17436 (N_17436,N_17097,N_17202);
nor U17437 (N_17437,N_17105,N_17098);
nand U17438 (N_17438,N_17215,N_17110);
xnor U17439 (N_17439,N_17185,N_17234);
nand U17440 (N_17440,N_17016,N_17127);
or U17441 (N_17441,N_17170,N_17248);
and U17442 (N_17442,N_17118,N_17126);
and U17443 (N_17443,N_17011,N_17047);
nand U17444 (N_17444,N_17046,N_17145);
nor U17445 (N_17445,N_17068,N_17056);
xnor U17446 (N_17446,N_17163,N_17215);
or U17447 (N_17447,N_17138,N_17245);
nand U17448 (N_17448,N_17022,N_17158);
or U17449 (N_17449,N_17169,N_17193);
or U17450 (N_17450,N_17224,N_17003);
nor U17451 (N_17451,N_17119,N_17210);
xnor U17452 (N_17452,N_17091,N_17040);
nand U17453 (N_17453,N_17139,N_17014);
nand U17454 (N_17454,N_17002,N_17150);
or U17455 (N_17455,N_17148,N_17110);
nand U17456 (N_17456,N_17212,N_17010);
nor U17457 (N_17457,N_17105,N_17234);
or U17458 (N_17458,N_17158,N_17071);
and U17459 (N_17459,N_17058,N_17204);
or U17460 (N_17460,N_17106,N_17153);
and U17461 (N_17461,N_17212,N_17215);
nand U17462 (N_17462,N_17247,N_17143);
and U17463 (N_17463,N_17001,N_17012);
and U17464 (N_17464,N_17050,N_17204);
or U17465 (N_17465,N_17106,N_17217);
or U17466 (N_17466,N_17030,N_17246);
and U17467 (N_17467,N_17074,N_17164);
nand U17468 (N_17468,N_17006,N_17218);
and U17469 (N_17469,N_17192,N_17163);
or U17470 (N_17470,N_17138,N_17195);
nand U17471 (N_17471,N_17016,N_17067);
and U17472 (N_17472,N_17094,N_17178);
nor U17473 (N_17473,N_17166,N_17078);
and U17474 (N_17474,N_17230,N_17204);
and U17475 (N_17475,N_17088,N_17202);
and U17476 (N_17476,N_17162,N_17185);
or U17477 (N_17477,N_17177,N_17060);
nand U17478 (N_17478,N_17096,N_17125);
nand U17479 (N_17479,N_17153,N_17244);
xnor U17480 (N_17480,N_17136,N_17134);
nand U17481 (N_17481,N_17113,N_17100);
or U17482 (N_17482,N_17022,N_17117);
or U17483 (N_17483,N_17203,N_17190);
nand U17484 (N_17484,N_17089,N_17176);
nor U17485 (N_17485,N_17056,N_17095);
nand U17486 (N_17486,N_17133,N_17017);
nor U17487 (N_17487,N_17145,N_17118);
nor U17488 (N_17488,N_17101,N_17093);
nand U17489 (N_17489,N_17039,N_17220);
and U17490 (N_17490,N_17122,N_17204);
and U17491 (N_17491,N_17196,N_17013);
or U17492 (N_17492,N_17036,N_17051);
and U17493 (N_17493,N_17244,N_17139);
nor U17494 (N_17494,N_17005,N_17188);
and U17495 (N_17495,N_17114,N_17067);
nor U17496 (N_17496,N_17155,N_17126);
nand U17497 (N_17497,N_17153,N_17039);
and U17498 (N_17498,N_17206,N_17010);
or U17499 (N_17499,N_17187,N_17105);
xor U17500 (N_17500,N_17435,N_17377);
nand U17501 (N_17501,N_17489,N_17257);
nor U17502 (N_17502,N_17326,N_17283);
nand U17503 (N_17503,N_17259,N_17334);
and U17504 (N_17504,N_17412,N_17278);
and U17505 (N_17505,N_17411,N_17343);
and U17506 (N_17506,N_17347,N_17492);
nand U17507 (N_17507,N_17498,N_17319);
nand U17508 (N_17508,N_17332,N_17462);
and U17509 (N_17509,N_17469,N_17318);
nor U17510 (N_17510,N_17494,N_17311);
nand U17511 (N_17511,N_17383,N_17300);
nor U17512 (N_17512,N_17262,N_17437);
and U17513 (N_17513,N_17299,N_17488);
or U17514 (N_17514,N_17407,N_17484);
nor U17515 (N_17515,N_17273,N_17364);
or U17516 (N_17516,N_17324,N_17301);
nor U17517 (N_17517,N_17430,N_17298);
nor U17518 (N_17518,N_17452,N_17256);
nor U17519 (N_17519,N_17395,N_17270);
or U17520 (N_17520,N_17281,N_17422);
nor U17521 (N_17521,N_17385,N_17370);
nand U17522 (N_17522,N_17445,N_17432);
and U17523 (N_17523,N_17255,N_17434);
or U17524 (N_17524,N_17316,N_17467);
or U17525 (N_17525,N_17457,N_17483);
or U17526 (N_17526,N_17455,N_17325);
nand U17527 (N_17527,N_17464,N_17312);
and U17528 (N_17528,N_17250,N_17386);
nor U17529 (N_17529,N_17353,N_17289);
or U17530 (N_17530,N_17405,N_17320);
or U17531 (N_17531,N_17305,N_17479);
and U17532 (N_17532,N_17307,N_17267);
nand U17533 (N_17533,N_17251,N_17297);
and U17534 (N_17534,N_17427,N_17482);
nand U17535 (N_17535,N_17431,N_17308);
nor U17536 (N_17536,N_17379,N_17294);
nand U17537 (N_17537,N_17272,N_17443);
nor U17538 (N_17538,N_17436,N_17402);
nor U17539 (N_17539,N_17252,N_17254);
xnor U17540 (N_17540,N_17453,N_17444);
and U17541 (N_17541,N_17306,N_17388);
nand U17542 (N_17542,N_17295,N_17361);
nand U17543 (N_17543,N_17313,N_17333);
or U17544 (N_17544,N_17274,N_17268);
nor U17545 (N_17545,N_17303,N_17440);
xor U17546 (N_17546,N_17354,N_17264);
or U17547 (N_17547,N_17459,N_17485);
xnor U17548 (N_17548,N_17378,N_17328);
xor U17549 (N_17549,N_17366,N_17321);
nand U17550 (N_17550,N_17408,N_17269);
nor U17551 (N_17551,N_17286,N_17428);
nor U17552 (N_17552,N_17403,N_17465);
or U17553 (N_17553,N_17439,N_17429);
and U17554 (N_17554,N_17397,N_17310);
xnor U17555 (N_17555,N_17461,N_17293);
and U17556 (N_17556,N_17367,N_17495);
nor U17557 (N_17557,N_17394,N_17265);
and U17558 (N_17558,N_17373,N_17474);
nor U17559 (N_17559,N_17337,N_17416);
and U17560 (N_17560,N_17491,N_17365);
nor U17561 (N_17561,N_17414,N_17350);
nand U17562 (N_17562,N_17392,N_17415);
nor U17563 (N_17563,N_17384,N_17380);
nor U17564 (N_17564,N_17327,N_17401);
or U17565 (N_17565,N_17263,N_17499);
nand U17566 (N_17566,N_17450,N_17399);
and U17567 (N_17567,N_17477,N_17302);
and U17568 (N_17568,N_17336,N_17331);
nand U17569 (N_17569,N_17476,N_17390);
or U17570 (N_17570,N_17381,N_17340);
and U17571 (N_17571,N_17418,N_17348);
and U17572 (N_17572,N_17292,N_17346);
and U17573 (N_17573,N_17339,N_17473);
xor U17574 (N_17574,N_17447,N_17456);
nand U17575 (N_17575,N_17420,N_17438);
nor U17576 (N_17576,N_17344,N_17351);
nand U17577 (N_17577,N_17478,N_17376);
nand U17578 (N_17578,N_17475,N_17374);
nor U17579 (N_17579,N_17466,N_17362);
nor U17580 (N_17580,N_17486,N_17309);
and U17581 (N_17581,N_17359,N_17451);
nor U17582 (N_17582,N_17279,N_17285);
and U17583 (N_17583,N_17345,N_17442);
nor U17584 (N_17584,N_17425,N_17463);
nand U17585 (N_17585,N_17446,N_17406);
nand U17586 (N_17586,N_17417,N_17448);
or U17587 (N_17587,N_17358,N_17314);
or U17588 (N_17588,N_17369,N_17372);
or U17589 (N_17589,N_17387,N_17282);
and U17590 (N_17590,N_17284,N_17360);
or U17591 (N_17591,N_17410,N_17341);
and U17592 (N_17592,N_17287,N_17441);
nand U17593 (N_17593,N_17330,N_17391);
xnor U17594 (N_17594,N_17490,N_17357);
xnor U17595 (N_17595,N_17496,N_17253);
or U17596 (N_17596,N_17355,N_17389);
or U17597 (N_17597,N_17460,N_17481);
nor U17598 (N_17598,N_17419,N_17413);
and U17599 (N_17599,N_17424,N_17480);
and U17600 (N_17600,N_17315,N_17421);
nand U17601 (N_17601,N_17280,N_17449);
nor U17602 (N_17602,N_17290,N_17471);
xnor U17603 (N_17603,N_17404,N_17396);
nand U17604 (N_17604,N_17393,N_17433);
xnor U17605 (N_17605,N_17382,N_17266);
and U17606 (N_17606,N_17323,N_17296);
and U17607 (N_17607,N_17458,N_17349);
xor U17608 (N_17608,N_17487,N_17423);
nor U17609 (N_17609,N_17375,N_17363);
xnor U17610 (N_17610,N_17258,N_17304);
nor U17611 (N_17611,N_17288,N_17260);
nor U17612 (N_17612,N_17342,N_17398);
or U17613 (N_17613,N_17400,N_17493);
nand U17614 (N_17614,N_17497,N_17356);
nor U17615 (N_17615,N_17472,N_17352);
or U17616 (N_17616,N_17454,N_17371);
nor U17617 (N_17617,N_17317,N_17271);
nor U17618 (N_17618,N_17470,N_17276);
nor U17619 (N_17619,N_17322,N_17277);
and U17620 (N_17620,N_17426,N_17409);
nand U17621 (N_17621,N_17291,N_17468);
nand U17622 (N_17622,N_17275,N_17368);
nand U17623 (N_17623,N_17338,N_17329);
nand U17624 (N_17624,N_17261,N_17335);
and U17625 (N_17625,N_17348,N_17446);
xnor U17626 (N_17626,N_17491,N_17334);
xnor U17627 (N_17627,N_17467,N_17408);
nor U17628 (N_17628,N_17253,N_17405);
and U17629 (N_17629,N_17472,N_17460);
xor U17630 (N_17630,N_17379,N_17404);
nor U17631 (N_17631,N_17293,N_17443);
and U17632 (N_17632,N_17285,N_17405);
nor U17633 (N_17633,N_17375,N_17345);
nor U17634 (N_17634,N_17279,N_17286);
and U17635 (N_17635,N_17450,N_17487);
xnor U17636 (N_17636,N_17280,N_17284);
nor U17637 (N_17637,N_17425,N_17306);
and U17638 (N_17638,N_17258,N_17341);
xnor U17639 (N_17639,N_17280,N_17269);
xnor U17640 (N_17640,N_17350,N_17309);
or U17641 (N_17641,N_17264,N_17344);
nand U17642 (N_17642,N_17475,N_17456);
or U17643 (N_17643,N_17377,N_17428);
and U17644 (N_17644,N_17493,N_17427);
nor U17645 (N_17645,N_17290,N_17497);
nand U17646 (N_17646,N_17368,N_17497);
or U17647 (N_17647,N_17281,N_17453);
or U17648 (N_17648,N_17451,N_17460);
nor U17649 (N_17649,N_17482,N_17365);
and U17650 (N_17650,N_17459,N_17377);
nor U17651 (N_17651,N_17254,N_17286);
or U17652 (N_17652,N_17415,N_17325);
or U17653 (N_17653,N_17463,N_17485);
nor U17654 (N_17654,N_17316,N_17483);
nor U17655 (N_17655,N_17456,N_17304);
or U17656 (N_17656,N_17470,N_17317);
nand U17657 (N_17657,N_17463,N_17395);
or U17658 (N_17658,N_17275,N_17298);
and U17659 (N_17659,N_17474,N_17448);
and U17660 (N_17660,N_17357,N_17452);
and U17661 (N_17661,N_17383,N_17396);
nand U17662 (N_17662,N_17436,N_17256);
or U17663 (N_17663,N_17451,N_17300);
and U17664 (N_17664,N_17475,N_17380);
nand U17665 (N_17665,N_17426,N_17294);
and U17666 (N_17666,N_17324,N_17371);
or U17667 (N_17667,N_17369,N_17392);
or U17668 (N_17668,N_17285,N_17354);
nand U17669 (N_17669,N_17325,N_17406);
nand U17670 (N_17670,N_17258,N_17311);
or U17671 (N_17671,N_17456,N_17350);
nor U17672 (N_17672,N_17482,N_17251);
and U17673 (N_17673,N_17420,N_17351);
or U17674 (N_17674,N_17408,N_17308);
nor U17675 (N_17675,N_17469,N_17417);
and U17676 (N_17676,N_17451,N_17349);
and U17677 (N_17677,N_17473,N_17264);
or U17678 (N_17678,N_17251,N_17320);
or U17679 (N_17679,N_17258,N_17312);
or U17680 (N_17680,N_17260,N_17474);
or U17681 (N_17681,N_17344,N_17314);
xor U17682 (N_17682,N_17466,N_17389);
or U17683 (N_17683,N_17439,N_17344);
and U17684 (N_17684,N_17325,N_17478);
or U17685 (N_17685,N_17414,N_17434);
and U17686 (N_17686,N_17262,N_17422);
nor U17687 (N_17687,N_17466,N_17322);
or U17688 (N_17688,N_17295,N_17469);
nor U17689 (N_17689,N_17396,N_17401);
nand U17690 (N_17690,N_17497,N_17337);
and U17691 (N_17691,N_17474,N_17295);
nor U17692 (N_17692,N_17312,N_17328);
nor U17693 (N_17693,N_17299,N_17458);
nor U17694 (N_17694,N_17317,N_17494);
and U17695 (N_17695,N_17378,N_17344);
xor U17696 (N_17696,N_17421,N_17256);
or U17697 (N_17697,N_17375,N_17301);
nor U17698 (N_17698,N_17418,N_17444);
nand U17699 (N_17699,N_17388,N_17367);
and U17700 (N_17700,N_17468,N_17350);
nor U17701 (N_17701,N_17268,N_17375);
nand U17702 (N_17702,N_17334,N_17264);
or U17703 (N_17703,N_17349,N_17318);
nor U17704 (N_17704,N_17381,N_17416);
nor U17705 (N_17705,N_17378,N_17433);
nand U17706 (N_17706,N_17431,N_17426);
nor U17707 (N_17707,N_17351,N_17284);
and U17708 (N_17708,N_17362,N_17425);
or U17709 (N_17709,N_17487,N_17292);
and U17710 (N_17710,N_17347,N_17294);
nand U17711 (N_17711,N_17433,N_17387);
and U17712 (N_17712,N_17406,N_17411);
nand U17713 (N_17713,N_17362,N_17305);
xor U17714 (N_17714,N_17466,N_17492);
and U17715 (N_17715,N_17257,N_17452);
or U17716 (N_17716,N_17388,N_17456);
nor U17717 (N_17717,N_17348,N_17498);
nor U17718 (N_17718,N_17350,N_17443);
or U17719 (N_17719,N_17480,N_17430);
nor U17720 (N_17720,N_17351,N_17473);
nor U17721 (N_17721,N_17441,N_17377);
and U17722 (N_17722,N_17363,N_17286);
and U17723 (N_17723,N_17441,N_17411);
and U17724 (N_17724,N_17356,N_17377);
nor U17725 (N_17725,N_17251,N_17274);
and U17726 (N_17726,N_17382,N_17356);
nand U17727 (N_17727,N_17275,N_17362);
nor U17728 (N_17728,N_17349,N_17305);
nor U17729 (N_17729,N_17284,N_17429);
or U17730 (N_17730,N_17361,N_17446);
and U17731 (N_17731,N_17441,N_17352);
nand U17732 (N_17732,N_17373,N_17282);
xnor U17733 (N_17733,N_17496,N_17313);
nor U17734 (N_17734,N_17463,N_17259);
xnor U17735 (N_17735,N_17443,N_17307);
or U17736 (N_17736,N_17251,N_17347);
nor U17737 (N_17737,N_17420,N_17484);
or U17738 (N_17738,N_17366,N_17283);
and U17739 (N_17739,N_17307,N_17292);
nor U17740 (N_17740,N_17470,N_17335);
nor U17741 (N_17741,N_17298,N_17270);
nand U17742 (N_17742,N_17450,N_17365);
nor U17743 (N_17743,N_17277,N_17358);
or U17744 (N_17744,N_17326,N_17319);
or U17745 (N_17745,N_17448,N_17487);
or U17746 (N_17746,N_17458,N_17350);
nand U17747 (N_17747,N_17368,N_17411);
nand U17748 (N_17748,N_17387,N_17293);
nor U17749 (N_17749,N_17398,N_17419);
xor U17750 (N_17750,N_17530,N_17503);
and U17751 (N_17751,N_17683,N_17524);
nor U17752 (N_17752,N_17581,N_17596);
xnor U17753 (N_17753,N_17553,N_17686);
and U17754 (N_17754,N_17500,N_17516);
nand U17755 (N_17755,N_17515,N_17710);
and U17756 (N_17756,N_17695,N_17501);
and U17757 (N_17757,N_17592,N_17608);
nor U17758 (N_17758,N_17625,N_17676);
or U17759 (N_17759,N_17694,N_17588);
nor U17760 (N_17760,N_17711,N_17585);
nor U17761 (N_17761,N_17582,N_17525);
and U17762 (N_17762,N_17613,N_17675);
or U17763 (N_17763,N_17743,N_17504);
nor U17764 (N_17764,N_17658,N_17598);
nor U17765 (N_17765,N_17571,N_17745);
nand U17766 (N_17766,N_17519,N_17599);
nor U17767 (N_17767,N_17680,N_17568);
nand U17768 (N_17768,N_17586,N_17632);
nand U17769 (N_17769,N_17721,N_17744);
nand U17770 (N_17770,N_17544,N_17541);
nor U17771 (N_17771,N_17562,N_17591);
nor U17772 (N_17772,N_17555,N_17733);
and U17773 (N_17773,N_17741,N_17656);
nand U17774 (N_17774,N_17737,N_17649);
and U17775 (N_17775,N_17612,N_17674);
or U17776 (N_17776,N_17651,N_17603);
nand U17777 (N_17777,N_17566,N_17734);
nand U17778 (N_17778,N_17652,N_17725);
nor U17779 (N_17779,N_17696,N_17636);
nand U17780 (N_17780,N_17546,N_17663);
and U17781 (N_17781,N_17563,N_17614);
and U17782 (N_17782,N_17653,N_17668);
and U17783 (N_17783,N_17620,N_17729);
nand U17784 (N_17784,N_17719,N_17552);
or U17785 (N_17785,N_17617,N_17749);
nor U17786 (N_17786,N_17679,N_17742);
xnor U17787 (N_17787,N_17600,N_17660);
and U17788 (N_17788,N_17528,N_17706);
xor U17789 (N_17789,N_17505,N_17661);
nand U17790 (N_17790,N_17644,N_17690);
and U17791 (N_17791,N_17681,N_17638);
nor U17792 (N_17792,N_17718,N_17510);
xor U17793 (N_17793,N_17507,N_17622);
nor U17794 (N_17794,N_17590,N_17716);
nand U17795 (N_17795,N_17672,N_17678);
and U17796 (N_17796,N_17704,N_17539);
or U17797 (N_17797,N_17692,N_17574);
or U17798 (N_17798,N_17579,N_17732);
nand U17799 (N_17799,N_17543,N_17626);
nand U17800 (N_17800,N_17748,N_17691);
and U17801 (N_17801,N_17575,N_17534);
and U17802 (N_17802,N_17667,N_17738);
or U17803 (N_17803,N_17594,N_17736);
or U17804 (N_17804,N_17578,N_17561);
and U17805 (N_17805,N_17560,N_17689);
xor U17806 (N_17806,N_17746,N_17595);
nand U17807 (N_17807,N_17610,N_17628);
nor U17808 (N_17808,N_17641,N_17542);
xor U17809 (N_17809,N_17739,N_17597);
and U17810 (N_17810,N_17580,N_17577);
and U17811 (N_17811,N_17526,N_17545);
and U17812 (N_17812,N_17670,N_17708);
nor U17813 (N_17813,N_17556,N_17611);
or U17814 (N_17814,N_17671,N_17509);
xnor U17815 (N_17815,N_17618,N_17720);
nand U17816 (N_17816,N_17634,N_17698);
or U17817 (N_17817,N_17664,N_17687);
xnor U17818 (N_17818,N_17537,N_17707);
or U17819 (N_17819,N_17605,N_17685);
nand U17820 (N_17820,N_17593,N_17547);
nor U17821 (N_17821,N_17647,N_17631);
or U17822 (N_17822,N_17551,N_17558);
and U17823 (N_17823,N_17601,N_17703);
and U17824 (N_17824,N_17548,N_17570);
nor U17825 (N_17825,N_17557,N_17702);
nand U17826 (N_17826,N_17657,N_17604);
nand U17827 (N_17827,N_17639,N_17502);
and U17828 (N_17828,N_17727,N_17701);
or U17829 (N_17829,N_17648,N_17536);
and U17830 (N_17830,N_17717,N_17514);
nor U17831 (N_17831,N_17659,N_17730);
nor U17832 (N_17832,N_17573,N_17511);
nor U17833 (N_17833,N_17728,N_17602);
and U17834 (N_17834,N_17535,N_17682);
and U17835 (N_17835,N_17633,N_17550);
nor U17836 (N_17836,N_17677,N_17508);
nor U17837 (N_17837,N_17584,N_17529);
or U17838 (N_17838,N_17665,N_17623);
nand U17839 (N_17839,N_17627,N_17650);
or U17840 (N_17840,N_17635,N_17666);
or U17841 (N_17841,N_17616,N_17576);
xor U17842 (N_17842,N_17731,N_17589);
or U17843 (N_17843,N_17724,N_17654);
nor U17844 (N_17844,N_17655,N_17523);
and U17845 (N_17845,N_17637,N_17567);
nor U17846 (N_17846,N_17583,N_17747);
and U17847 (N_17847,N_17533,N_17640);
nor U17848 (N_17848,N_17615,N_17700);
xnor U17849 (N_17849,N_17669,N_17532);
and U17850 (N_17850,N_17735,N_17609);
nor U17851 (N_17851,N_17619,N_17606);
nand U17852 (N_17852,N_17624,N_17565);
xnor U17853 (N_17853,N_17642,N_17722);
nand U17854 (N_17854,N_17549,N_17643);
and U17855 (N_17855,N_17629,N_17512);
and U17856 (N_17856,N_17518,N_17527);
or U17857 (N_17857,N_17569,N_17673);
and U17858 (N_17858,N_17705,N_17693);
and U17859 (N_17859,N_17531,N_17699);
or U17860 (N_17860,N_17572,N_17715);
nand U17861 (N_17861,N_17621,N_17538);
nor U17862 (N_17862,N_17712,N_17513);
or U17863 (N_17863,N_17517,N_17564);
and U17864 (N_17864,N_17684,N_17714);
and U17865 (N_17865,N_17662,N_17559);
and U17866 (N_17866,N_17587,N_17521);
and U17867 (N_17867,N_17688,N_17554);
nand U17868 (N_17868,N_17726,N_17506);
nand U17869 (N_17869,N_17522,N_17713);
or U17870 (N_17870,N_17646,N_17607);
nand U17871 (N_17871,N_17723,N_17630);
nand U17872 (N_17872,N_17709,N_17645);
or U17873 (N_17873,N_17540,N_17520);
and U17874 (N_17874,N_17697,N_17740);
or U17875 (N_17875,N_17708,N_17735);
and U17876 (N_17876,N_17670,N_17663);
and U17877 (N_17877,N_17723,N_17737);
nor U17878 (N_17878,N_17707,N_17552);
nor U17879 (N_17879,N_17545,N_17559);
nand U17880 (N_17880,N_17622,N_17637);
and U17881 (N_17881,N_17740,N_17650);
nand U17882 (N_17882,N_17510,N_17659);
nand U17883 (N_17883,N_17615,N_17665);
and U17884 (N_17884,N_17511,N_17637);
or U17885 (N_17885,N_17719,N_17627);
and U17886 (N_17886,N_17540,N_17573);
and U17887 (N_17887,N_17561,N_17734);
or U17888 (N_17888,N_17630,N_17740);
xor U17889 (N_17889,N_17513,N_17724);
and U17890 (N_17890,N_17735,N_17595);
or U17891 (N_17891,N_17588,N_17662);
and U17892 (N_17892,N_17726,N_17537);
or U17893 (N_17893,N_17677,N_17614);
and U17894 (N_17894,N_17547,N_17576);
nand U17895 (N_17895,N_17679,N_17511);
or U17896 (N_17896,N_17528,N_17657);
and U17897 (N_17897,N_17706,N_17598);
and U17898 (N_17898,N_17658,N_17576);
xor U17899 (N_17899,N_17593,N_17528);
nand U17900 (N_17900,N_17586,N_17502);
nand U17901 (N_17901,N_17583,N_17700);
nor U17902 (N_17902,N_17655,N_17576);
nand U17903 (N_17903,N_17638,N_17586);
or U17904 (N_17904,N_17698,N_17582);
nand U17905 (N_17905,N_17525,N_17550);
xnor U17906 (N_17906,N_17669,N_17661);
nand U17907 (N_17907,N_17599,N_17699);
xor U17908 (N_17908,N_17511,N_17576);
or U17909 (N_17909,N_17510,N_17600);
xnor U17910 (N_17910,N_17604,N_17526);
and U17911 (N_17911,N_17579,N_17722);
xnor U17912 (N_17912,N_17717,N_17611);
and U17913 (N_17913,N_17562,N_17604);
nand U17914 (N_17914,N_17655,N_17654);
nand U17915 (N_17915,N_17624,N_17663);
and U17916 (N_17916,N_17507,N_17711);
nor U17917 (N_17917,N_17691,N_17617);
or U17918 (N_17918,N_17549,N_17742);
xor U17919 (N_17919,N_17587,N_17573);
nand U17920 (N_17920,N_17671,N_17674);
nand U17921 (N_17921,N_17561,N_17709);
or U17922 (N_17922,N_17605,N_17649);
and U17923 (N_17923,N_17736,N_17575);
and U17924 (N_17924,N_17728,N_17551);
nor U17925 (N_17925,N_17661,N_17557);
nand U17926 (N_17926,N_17734,N_17708);
nand U17927 (N_17927,N_17656,N_17585);
or U17928 (N_17928,N_17600,N_17628);
nand U17929 (N_17929,N_17732,N_17606);
xor U17930 (N_17930,N_17683,N_17595);
xor U17931 (N_17931,N_17602,N_17650);
xor U17932 (N_17932,N_17513,N_17605);
nor U17933 (N_17933,N_17545,N_17673);
or U17934 (N_17934,N_17677,N_17573);
nor U17935 (N_17935,N_17646,N_17745);
nand U17936 (N_17936,N_17564,N_17635);
nand U17937 (N_17937,N_17683,N_17536);
and U17938 (N_17938,N_17608,N_17653);
and U17939 (N_17939,N_17724,N_17702);
or U17940 (N_17940,N_17511,N_17656);
and U17941 (N_17941,N_17649,N_17540);
nand U17942 (N_17942,N_17628,N_17643);
or U17943 (N_17943,N_17651,N_17561);
xor U17944 (N_17944,N_17728,N_17683);
nor U17945 (N_17945,N_17500,N_17669);
nand U17946 (N_17946,N_17663,N_17687);
or U17947 (N_17947,N_17656,N_17721);
nand U17948 (N_17948,N_17592,N_17719);
nand U17949 (N_17949,N_17540,N_17683);
nor U17950 (N_17950,N_17542,N_17552);
nor U17951 (N_17951,N_17722,N_17531);
nor U17952 (N_17952,N_17697,N_17543);
nor U17953 (N_17953,N_17515,N_17587);
nor U17954 (N_17954,N_17526,N_17580);
xnor U17955 (N_17955,N_17723,N_17681);
or U17956 (N_17956,N_17622,N_17645);
nor U17957 (N_17957,N_17591,N_17692);
nor U17958 (N_17958,N_17519,N_17707);
or U17959 (N_17959,N_17690,N_17585);
xor U17960 (N_17960,N_17630,N_17744);
nand U17961 (N_17961,N_17645,N_17516);
nand U17962 (N_17962,N_17734,N_17635);
and U17963 (N_17963,N_17650,N_17529);
nor U17964 (N_17964,N_17740,N_17666);
and U17965 (N_17965,N_17643,N_17666);
nor U17966 (N_17966,N_17599,N_17726);
xnor U17967 (N_17967,N_17675,N_17704);
or U17968 (N_17968,N_17734,N_17581);
or U17969 (N_17969,N_17719,N_17642);
and U17970 (N_17970,N_17639,N_17749);
or U17971 (N_17971,N_17523,N_17732);
nor U17972 (N_17972,N_17721,N_17545);
nor U17973 (N_17973,N_17520,N_17536);
nor U17974 (N_17974,N_17652,N_17564);
nand U17975 (N_17975,N_17627,N_17607);
or U17976 (N_17976,N_17584,N_17720);
nand U17977 (N_17977,N_17552,N_17680);
xnor U17978 (N_17978,N_17539,N_17746);
and U17979 (N_17979,N_17709,N_17693);
nor U17980 (N_17980,N_17664,N_17667);
nand U17981 (N_17981,N_17619,N_17609);
nor U17982 (N_17982,N_17522,N_17635);
nor U17983 (N_17983,N_17534,N_17661);
nand U17984 (N_17984,N_17740,N_17658);
and U17985 (N_17985,N_17632,N_17685);
or U17986 (N_17986,N_17537,N_17671);
and U17987 (N_17987,N_17693,N_17623);
and U17988 (N_17988,N_17709,N_17570);
nor U17989 (N_17989,N_17613,N_17542);
nor U17990 (N_17990,N_17703,N_17690);
nor U17991 (N_17991,N_17706,N_17664);
xor U17992 (N_17992,N_17616,N_17547);
or U17993 (N_17993,N_17563,N_17679);
nand U17994 (N_17994,N_17582,N_17566);
nor U17995 (N_17995,N_17597,N_17511);
nor U17996 (N_17996,N_17636,N_17624);
nand U17997 (N_17997,N_17614,N_17601);
nand U17998 (N_17998,N_17612,N_17642);
nand U17999 (N_17999,N_17506,N_17736);
or U18000 (N_18000,N_17877,N_17836);
nand U18001 (N_18001,N_17878,N_17982);
or U18002 (N_18002,N_17862,N_17959);
nor U18003 (N_18003,N_17827,N_17778);
nand U18004 (N_18004,N_17930,N_17957);
and U18005 (N_18005,N_17782,N_17979);
and U18006 (N_18006,N_17758,N_17799);
nor U18007 (N_18007,N_17847,N_17820);
nor U18008 (N_18008,N_17876,N_17939);
nand U18009 (N_18009,N_17993,N_17826);
and U18010 (N_18010,N_17938,N_17814);
and U18011 (N_18011,N_17794,N_17991);
nor U18012 (N_18012,N_17984,N_17844);
or U18013 (N_18013,N_17910,N_17797);
nor U18014 (N_18014,N_17976,N_17951);
and U18015 (N_18015,N_17969,N_17856);
or U18016 (N_18016,N_17792,N_17981);
xor U18017 (N_18017,N_17815,N_17953);
or U18018 (N_18018,N_17803,N_17915);
or U18019 (N_18019,N_17858,N_17997);
or U18020 (N_18020,N_17934,N_17839);
nor U18021 (N_18021,N_17865,N_17898);
nor U18022 (N_18022,N_17870,N_17837);
or U18023 (N_18023,N_17774,N_17853);
or U18024 (N_18024,N_17808,N_17777);
nand U18025 (N_18025,N_17932,N_17947);
and U18026 (N_18026,N_17920,N_17955);
or U18027 (N_18027,N_17998,N_17761);
and U18028 (N_18028,N_17764,N_17968);
or U18029 (N_18029,N_17884,N_17956);
and U18030 (N_18030,N_17874,N_17785);
and U18031 (N_18031,N_17929,N_17845);
nand U18032 (N_18032,N_17965,N_17816);
nand U18033 (N_18033,N_17834,N_17952);
or U18034 (N_18034,N_17882,N_17909);
and U18035 (N_18035,N_17750,N_17925);
nand U18036 (N_18036,N_17994,N_17786);
and U18037 (N_18037,N_17989,N_17897);
and U18038 (N_18038,N_17978,N_17887);
xnor U18039 (N_18039,N_17986,N_17935);
nor U18040 (N_18040,N_17917,N_17829);
and U18041 (N_18041,N_17775,N_17755);
nor U18042 (N_18042,N_17894,N_17942);
and U18043 (N_18043,N_17901,N_17893);
and U18044 (N_18044,N_17810,N_17937);
and U18045 (N_18045,N_17851,N_17988);
or U18046 (N_18046,N_17971,N_17788);
nand U18047 (N_18047,N_17944,N_17921);
nor U18048 (N_18048,N_17802,N_17916);
nor U18049 (N_18049,N_17757,N_17871);
nand U18050 (N_18050,N_17756,N_17776);
nand U18051 (N_18051,N_17752,N_17817);
nor U18052 (N_18052,N_17945,N_17821);
xor U18053 (N_18053,N_17967,N_17779);
or U18054 (N_18054,N_17828,N_17783);
and U18055 (N_18055,N_17983,N_17905);
and U18056 (N_18056,N_17970,N_17809);
nor U18057 (N_18057,N_17825,N_17843);
nor U18058 (N_18058,N_17850,N_17823);
nand U18059 (N_18059,N_17769,N_17973);
nor U18060 (N_18060,N_17869,N_17906);
and U18061 (N_18061,N_17966,N_17943);
nor U18062 (N_18062,N_17807,N_17914);
nand U18063 (N_18063,N_17846,N_17805);
and U18064 (N_18064,N_17883,N_17963);
or U18065 (N_18065,N_17762,N_17811);
and U18066 (N_18066,N_17852,N_17949);
nor U18067 (N_18067,N_17872,N_17889);
or U18068 (N_18068,N_17787,N_17855);
and U18069 (N_18069,N_17833,N_17796);
nor U18070 (N_18070,N_17751,N_17767);
nor U18071 (N_18071,N_17912,N_17886);
nand U18072 (N_18072,N_17819,N_17806);
nand U18073 (N_18073,N_17922,N_17899);
or U18074 (N_18074,N_17964,N_17911);
nor U18075 (N_18075,N_17812,N_17908);
nand U18076 (N_18076,N_17880,N_17977);
nand U18077 (N_18077,N_17900,N_17896);
or U18078 (N_18078,N_17924,N_17831);
and U18079 (N_18079,N_17781,N_17798);
nand U18080 (N_18080,N_17926,N_17879);
nor U18081 (N_18081,N_17904,N_17913);
nor U18082 (N_18082,N_17830,N_17974);
and U18083 (N_18083,N_17996,N_17948);
or U18084 (N_18084,N_17760,N_17768);
nor U18085 (N_18085,N_17773,N_17753);
and U18086 (N_18086,N_17946,N_17840);
and U18087 (N_18087,N_17789,N_17958);
nor U18088 (N_18088,N_17867,N_17864);
nand U18089 (N_18089,N_17780,N_17891);
or U18090 (N_18090,N_17972,N_17890);
or U18091 (N_18091,N_17975,N_17868);
nand U18092 (N_18092,N_17784,N_17854);
nand U18093 (N_18093,N_17860,N_17818);
nand U18094 (N_18094,N_17990,N_17822);
nand U18095 (N_18095,N_17927,N_17841);
nand U18096 (N_18096,N_17804,N_17923);
nand U18097 (N_18097,N_17832,N_17875);
xor U18098 (N_18098,N_17903,N_17961);
nor U18099 (N_18099,N_17892,N_17885);
nand U18100 (N_18100,N_17863,N_17772);
nor U18101 (N_18101,N_17962,N_17933);
nor U18102 (N_18102,N_17848,N_17980);
or U18103 (N_18103,N_17861,N_17992);
xor U18104 (N_18104,N_17941,N_17763);
nand U18105 (N_18105,N_17759,N_17881);
or U18106 (N_18106,N_17960,N_17936);
nand U18107 (N_18107,N_17907,N_17813);
nor U18108 (N_18108,N_17928,N_17824);
nor U18109 (N_18109,N_17793,N_17866);
and U18110 (N_18110,N_17835,N_17771);
and U18111 (N_18111,N_17770,N_17791);
nor U18112 (N_18112,N_17838,N_17987);
xnor U18113 (N_18113,N_17754,N_17931);
xnor U18114 (N_18114,N_17918,N_17999);
and U18115 (N_18115,N_17954,N_17800);
nor U18116 (N_18116,N_17849,N_17873);
and U18117 (N_18117,N_17795,N_17950);
or U18118 (N_18118,N_17995,N_17859);
and U18119 (N_18119,N_17801,N_17895);
xnor U18120 (N_18120,N_17985,N_17902);
nand U18121 (N_18121,N_17765,N_17766);
and U18122 (N_18122,N_17888,N_17842);
and U18123 (N_18123,N_17940,N_17790);
nand U18124 (N_18124,N_17857,N_17919);
or U18125 (N_18125,N_17920,N_17857);
and U18126 (N_18126,N_17911,N_17759);
and U18127 (N_18127,N_17946,N_17939);
xnor U18128 (N_18128,N_17847,N_17886);
or U18129 (N_18129,N_17798,N_17765);
nor U18130 (N_18130,N_17831,N_17935);
nand U18131 (N_18131,N_17870,N_17855);
nor U18132 (N_18132,N_17921,N_17784);
or U18133 (N_18133,N_17929,N_17761);
and U18134 (N_18134,N_17775,N_17925);
nand U18135 (N_18135,N_17859,N_17968);
nor U18136 (N_18136,N_17928,N_17979);
and U18137 (N_18137,N_17951,N_17828);
xnor U18138 (N_18138,N_17761,N_17820);
and U18139 (N_18139,N_17933,N_17899);
nand U18140 (N_18140,N_17912,N_17817);
or U18141 (N_18141,N_17795,N_17814);
and U18142 (N_18142,N_17908,N_17779);
nand U18143 (N_18143,N_17918,N_17825);
and U18144 (N_18144,N_17823,N_17941);
xnor U18145 (N_18145,N_17964,N_17931);
or U18146 (N_18146,N_17811,N_17758);
xnor U18147 (N_18147,N_17762,N_17884);
nor U18148 (N_18148,N_17816,N_17777);
or U18149 (N_18149,N_17775,N_17874);
or U18150 (N_18150,N_17836,N_17945);
nand U18151 (N_18151,N_17945,N_17962);
nor U18152 (N_18152,N_17852,N_17932);
or U18153 (N_18153,N_17992,N_17916);
nor U18154 (N_18154,N_17995,N_17872);
nand U18155 (N_18155,N_17847,N_17889);
or U18156 (N_18156,N_17769,N_17791);
or U18157 (N_18157,N_17902,N_17765);
or U18158 (N_18158,N_17882,N_17804);
or U18159 (N_18159,N_17776,N_17920);
xor U18160 (N_18160,N_17812,N_17782);
nand U18161 (N_18161,N_17819,N_17943);
nand U18162 (N_18162,N_17885,N_17979);
nand U18163 (N_18163,N_17964,N_17815);
nand U18164 (N_18164,N_17770,N_17864);
nor U18165 (N_18165,N_17767,N_17958);
xnor U18166 (N_18166,N_17973,N_17886);
nor U18167 (N_18167,N_17904,N_17861);
and U18168 (N_18168,N_17811,N_17886);
nand U18169 (N_18169,N_17842,N_17882);
or U18170 (N_18170,N_17765,N_17975);
xnor U18171 (N_18171,N_17865,N_17988);
or U18172 (N_18172,N_17852,N_17896);
nand U18173 (N_18173,N_17782,N_17923);
and U18174 (N_18174,N_17974,N_17962);
nor U18175 (N_18175,N_17782,N_17992);
or U18176 (N_18176,N_17988,N_17849);
nand U18177 (N_18177,N_17873,N_17977);
xnor U18178 (N_18178,N_17814,N_17940);
nor U18179 (N_18179,N_17786,N_17944);
nand U18180 (N_18180,N_17832,N_17856);
nand U18181 (N_18181,N_17985,N_17862);
nor U18182 (N_18182,N_17807,N_17960);
nand U18183 (N_18183,N_17818,N_17798);
nor U18184 (N_18184,N_17844,N_17854);
nand U18185 (N_18185,N_17934,N_17925);
nor U18186 (N_18186,N_17936,N_17999);
xor U18187 (N_18187,N_17885,N_17837);
xor U18188 (N_18188,N_17893,N_17896);
xor U18189 (N_18189,N_17753,N_17952);
xnor U18190 (N_18190,N_17926,N_17775);
and U18191 (N_18191,N_17752,N_17900);
xor U18192 (N_18192,N_17844,N_17934);
or U18193 (N_18193,N_17935,N_17921);
or U18194 (N_18194,N_17760,N_17967);
or U18195 (N_18195,N_17901,N_17960);
and U18196 (N_18196,N_17936,N_17932);
nor U18197 (N_18197,N_17754,N_17944);
nand U18198 (N_18198,N_17964,N_17778);
or U18199 (N_18199,N_17939,N_17921);
and U18200 (N_18200,N_17974,N_17872);
nor U18201 (N_18201,N_17848,N_17770);
nand U18202 (N_18202,N_17777,N_17925);
nand U18203 (N_18203,N_17989,N_17823);
nor U18204 (N_18204,N_17854,N_17971);
and U18205 (N_18205,N_17975,N_17812);
nor U18206 (N_18206,N_17961,N_17874);
and U18207 (N_18207,N_17832,N_17887);
xnor U18208 (N_18208,N_17772,N_17876);
and U18209 (N_18209,N_17960,N_17974);
nand U18210 (N_18210,N_17903,N_17808);
nand U18211 (N_18211,N_17921,N_17865);
xor U18212 (N_18212,N_17862,N_17753);
or U18213 (N_18213,N_17776,N_17926);
or U18214 (N_18214,N_17972,N_17868);
and U18215 (N_18215,N_17967,N_17933);
nand U18216 (N_18216,N_17873,N_17952);
and U18217 (N_18217,N_17751,N_17827);
nand U18218 (N_18218,N_17985,N_17860);
or U18219 (N_18219,N_17798,N_17903);
nor U18220 (N_18220,N_17888,N_17966);
nor U18221 (N_18221,N_17847,N_17957);
nand U18222 (N_18222,N_17839,N_17771);
nand U18223 (N_18223,N_17788,N_17846);
or U18224 (N_18224,N_17969,N_17841);
nor U18225 (N_18225,N_17943,N_17820);
nor U18226 (N_18226,N_17977,N_17817);
or U18227 (N_18227,N_17937,N_17806);
or U18228 (N_18228,N_17823,N_17867);
and U18229 (N_18229,N_17792,N_17800);
and U18230 (N_18230,N_17871,N_17979);
and U18231 (N_18231,N_17938,N_17997);
xor U18232 (N_18232,N_17937,N_17819);
nor U18233 (N_18233,N_17834,N_17811);
nor U18234 (N_18234,N_17962,N_17821);
nand U18235 (N_18235,N_17976,N_17796);
xor U18236 (N_18236,N_17908,N_17832);
nor U18237 (N_18237,N_17777,N_17776);
and U18238 (N_18238,N_17924,N_17803);
and U18239 (N_18239,N_17781,N_17962);
nand U18240 (N_18240,N_17806,N_17809);
xnor U18241 (N_18241,N_17753,N_17782);
or U18242 (N_18242,N_17962,N_17876);
or U18243 (N_18243,N_17847,N_17875);
nor U18244 (N_18244,N_17960,N_17832);
or U18245 (N_18245,N_17891,N_17957);
nor U18246 (N_18246,N_17814,N_17917);
or U18247 (N_18247,N_17925,N_17832);
or U18248 (N_18248,N_17822,N_17899);
and U18249 (N_18249,N_17890,N_17796);
and U18250 (N_18250,N_18168,N_18004);
and U18251 (N_18251,N_18121,N_18194);
xnor U18252 (N_18252,N_18196,N_18115);
xor U18253 (N_18253,N_18070,N_18128);
xnor U18254 (N_18254,N_18003,N_18110);
xor U18255 (N_18255,N_18246,N_18107);
nand U18256 (N_18256,N_18187,N_18222);
nand U18257 (N_18257,N_18073,N_18149);
nor U18258 (N_18258,N_18211,N_18068);
nand U18259 (N_18259,N_18025,N_18199);
nand U18260 (N_18260,N_18086,N_18219);
nor U18261 (N_18261,N_18208,N_18132);
nor U18262 (N_18262,N_18021,N_18046);
or U18263 (N_18263,N_18190,N_18005);
xnor U18264 (N_18264,N_18215,N_18001);
nor U18265 (N_18265,N_18154,N_18014);
nand U18266 (N_18266,N_18147,N_18201);
or U18267 (N_18267,N_18036,N_18085);
xor U18268 (N_18268,N_18138,N_18205);
xor U18269 (N_18269,N_18016,N_18009);
nand U18270 (N_18270,N_18166,N_18091);
nor U18271 (N_18271,N_18139,N_18209);
or U18272 (N_18272,N_18096,N_18114);
or U18273 (N_18273,N_18071,N_18062);
and U18274 (N_18274,N_18193,N_18051);
nand U18275 (N_18275,N_18028,N_18093);
nor U18276 (N_18276,N_18191,N_18109);
and U18277 (N_18277,N_18133,N_18239);
nand U18278 (N_18278,N_18000,N_18195);
and U18279 (N_18279,N_18017,N_18220);
nor U18280 (N_18280,N_18098,N_18024);
and U18281 (N_18281,N_18235,N_18167);
or U18282 (N_18282,N_18026,N_18238);
and U18283 (N_18283,N_18088,N_18100);
and U18284 (N_18284,N_18069,N_18175);
nand U18285 (N_18285,N_18124,N_18127);
xnor U18286 (N_18286,N_18226,N_18185);
or U18287 (N_18287,N_18148,N_18162);
nor U18288 (N_18288,N_18081,N_18237);
nand U18289 (N_18289,N_18032,N_18053);
and U18290 (N_18290,N_18008,N_18249);
or U18291 (N_18291,N_18236,N_18058);
or U18292 (N_18292,N_18192,N_18160);
or U18293 (N_18293,N_18035,N_18182);
or U18294 (N_18294,N_18243,N_18152);
or U18295 (N_18295,N_18130,N_18184);
xnor U18296 (N_18296,N_18150,N_18179);
or U18297 (N_18297,N_18020,N_18097);
and U18298 (N_18298,N_18012,N_18181);
nor U18299 (N_18299,N_18059,N_18230);
nand U18300 (N_18300,N_18161,N_18045);
or U18301 (N_18301,N_18142,N_18052);
or U18302 (N_18302,N_18146,N_18087);
nand U18303 (N_18303,N_18171,N_18145);
nand U18304 (N_18304,N_18119,N_18228);
and U18305 (N_18305,N_18245,N_18247);
nand U18306 (N_18306,N_18013,N_18105);
or U18307 (N_18307,N_18083,N_18022);
nand U18308 (N_18308,N_18204,N_18177);
or U18309 (N_18309,N_18134,N_18223);
and U18310 (N_18310,N_18011,N_18126);
xnor U18311 (N_18311,N_18188,N_18065);
nor U18312 (N_18312,N_18094,N_18061);
or U18313 (N_18313,N_18057,N_18244);
nand U18314 (N_18314,N_18229,N_18186);
nor U18315 (N_18315,N_18210,N_18200);
and U18316 (N_18316,N_18217,N_18082);
nand U18317 (N_18317,N_18189,N_18066);
and U18318 (N_18318,N_18033,N_18136);
nand U18319 (N_18319,N_18180,N_18216);
nand U18320 (N_18320,N_18163,N_18221);
nor U18321 (N_18321,N_18248,N_18164);
and U18322 (N_18322,N_18241,N_18002);
nand U18323 (N_18323,N_18074,N_18176);
xor U18324 (N_18324,N_18039,N_18027);
nor U18325 (N_18325,N_18231,N_18112);
or U18326 (N_18326,N_18178,N_18144);
or U18327 (N_18327,N_18125,N_18084);
nand U18328 (N_18328,N_18077,N_18198);
nand U18329 (N_18329,N_18055,N_18054);
and U18330 (N_18330,N_18099,N_18117);
nor U18331 (N_18331,N_18072,N_18232);
nor U18332 (N_18332,N_18056,N_18165);
nand U18333 (N_18333,N_18170,N_18102);
xnor U18334 (N_18334,N_18106,N_18218);
nand U18335 (N_18335,N_18183,N_18143);
and U18336 (N_18336,N_18120,N_18037);
nand U18337 (N_18337,N_18048,N_18038);
nand U18338 (N_18338,N_18197,N_18063);
xnor U18339 (N_18339,N_18101,N_18233);
nor U18340 (N_18340,N_18043,N_18019);
nand U18341 (N_18341,N_18047,N_18067);
or U18342 (N_18342,N_18213,N_18123);
nand U18343 (N_18343,N_18122,N_18018);
nand U18344 (N_18344,N_18203,N_18023);
and U18345 (N_18345,N_18156,N_18049);
and U18346 (N_18346,N_18040,N_18075);
and U18347 (N_18347,N_18174,N_18206);
and U18348 (N_18348,N_18140,N_18118);
and U18349 (N_18349,N_18214,N_18030);
and U18350 (N_18350,N_18079,N_18010);
nand U18351 (N_18351,N_18006,N_18064);
or U18352 (N_18352,N_18207,N_18224);
nand U18353 (N_18353,N_18078,N_18092);
nor U18354 (N_18354,N_18007,N_18242);
nand U18355 (N_18355,N_18135,N_18157);
and U18356 (N_18356,N_18015,N_18080);
and U18357 (N_18357,N_18050,N_18113);
or U18358 (N_18358,N_18225,N_18173);
nand U18359 (N_18359,N_18159,N_18169);
and U18360 (N_18360,N_18095,N_18111);
nor U18361 (N_18361,N_18041,N_18108);
nor U18362 (N_18362,N_18090,N_18116);
or U18363 (N_18363,N_18131,N_18137);
nand U18364 (N_18364,N_18042,N_18044);
nand U18365 (N_18365,N_18240,N_18031);
and U18366 (N_18366,N_18060,N_18227);
and U18367 (N_18367,N_18141,N_18153);
nor U18368 (N_18368,N_18104,N_18103);
nand U18369 (N_18369,N_18034,N_18151);
nand U18370 (N_18370,N_18158,N_18212);
or U18371 (N_18371,N_18155,N_18234);
nor U18372 (N_18372,N_18172,N_18129);
nand U18373 (N_18373,N_18089,N_18076);
nand U18374 (N_18374,N_18202,N_18029);
nand U18375 (N_18375,N_18181,N_18183);
or U18376 (N_18376,N_18186,N_18216);
nand U18377 (N_18377,N_18189,N_18039);
nand U18378 (N_18378,N_18209,N_18093);
xor U18379 (N_18379,N_18075,N_18031);
or U18380 (N_18380,N_18119,N_18164);
nor U18381 (N_18381,N_18077,N_18058);
and U18382 (N_18382,N_18195,N_18115);
and U18383 (N_18383,N_18068,N_18107);
or U18384 (N_18384,N_18015,N_18114);
nor U18385 (N_18385,N_18004,N_18237);
nand U18386 (N_18386,N_18072,N_18031);
nor U18387 (N_18387,N_18112,N_18053);
and U18388 (N_18388,N_18187,N_18020);
and U18389 (N_18389,N_18001,N_18032);
and U18390 (N_18390,N_18185,N_18089);
nand U18391 (N_18391,N_18180,N_18241);
and U18392 (N_18392,N_18043,N_18130);
nor U18393 (N_18393,N_18046,N_18127);
nand U18394 (N_18394,N_18230,N_18065);
nor U18395 (N_18395,N_18141,N_18220);
nor U18396 (N_18396,N_18011,N_18170);
nand U18397 (N_18397,N_18237,N_18050);
and U18398 (N_18398,N_18022,N_18053);
and U18399 (N_18399,N_18078,N_18118);
xor U18400 (N_18400,N_18057,N_18190);
and U18401 (N_18401,N_18063,N_18156);
nand U18402 (N_18402,N_18090,N_18224);
and U18403 (N_18403,N_18098,N_18003);
and U18404 (N_18404,N_18114,N_18085);
or U18405 (N_18405,N_18022,N_18166);
nor U18406 (N_18406,N_18106,N_18156);
and U18407 (N_18407,N_18192,N_18162);
and U18408 (N_18408,N_18085,N_18065);
and U18409 (N_18409,N_18130,N_18137);
nand U18410 (N_18410,N_18089,N_18233);
and U18411 (N_18411,N_18094,N_18060);
nor U18412 (N_18412,N_18160,N_18206);
or U18413 (N_18413,N_18164,N_18084);
nand U18414 (N_18414,N_18153,N_18085);
nand U18415 (N_18415,N_18213,N_18031);
and U18416 (N_18416,N_18033,N_18034);
nor U18417 (N_18417,N_18131,N_18148);
or U18418 (N_18418,N_18015,N_18178);
or U18419 (N_18419,N_18077,N_18196);
or U18420 (N_18420,N_18016,N_18109);
and U18421 (N_18421,N_18046,N_18208);
or U18422 (N_18422,N_18225,N_18136);
and U18423 (N_18423,N_18099,N_18148);
or U18424 (N_18424,N_18132,N_18148);
or U18425 (N_18425,N_18141,N_18236);
xnor U18426 (N_18426,N_18090,N_18165);
or U18427 (N_18427,N_18122,N_18052);
nor U18428 (N_18428,N_18075,N_18037);
nand U18429 (N_18429,N_18153,N_18001);
nor U18430 (N_18430,N_18129,N_18121);
nor U18431 (N_18431,N_18154,N_18046);
and U18432 (N_18432,N_18119,N_18005);
or U18433 (N_18433,N_18044,N_18240);
nor U18434 (N_18434,N_18107,N_18030);
and U18435 (N_18435,N_18173,N_18085);
nor U18436 (N_18436,N_18245,N_18249);
nand U18437 (N_18437,N_18152,N_18083);
nor U18438 (N_18438,N_18083,N_18204);
nand U18439 (N_18439,N_18001,N_18131);
nor U18440 (N_18440,N_18166,N_18076);
or U18441 (N_18441,N_18166,N_18070);
xnor U18442 (N_18442,N_18127,N_18166);
or U18443 (N_18443,N_18113,N_18155);
and U18444 (N_18444,N_18215,N_18151);
or U18445 (N_18445,N_18021,N_18207);
or U18446 (N_18446,N_18091,N_18099);
nand U18447 (N_18447,N_18121,N_18055);
nor U18448 (N_18448,N_18181,N_18120);
or U18449 (N_18449,N_18121,N_18021);
or U18450 (N_18450,N_18212,N_18166);
or U18451 (N_18451,N_18242,N_18220);
and U18452 (N_18452,N_18186,N_18050);
nor U18453 (N_18453,N_18023,N_18095);
xor U18454 (N_18454,N_18069,N_18087);
nand U18455 (N_18455,N_18154,N_18030);
or U18456 (N_18456,N_18079,N_18054);
nor U18457 (N_18457,N_18222,N_18181);
and U18458 (N_18458,N_18248,N_18175);
or U18459 (N_18459,N_18171,N_18188);
nand U18460 (N_18460,N_18073,N_18009);
or U18461 (N_18461,N_18159,N_18071);
and U18462 (N_18462,N_18026,N_18234);
xor U18463 (N_18463,N_18120,N_18099);
or U18464 (N_18464,N_18117,N_18061);
and U18465 (N_18465,N_18211,N_18001);
or U18466 (N_18466,N_18046,N_18239);
or U18467 (N_18467,N_18109,N_18212);
or U18468 (N_18468,N_18166,N_18163);
nand U18469 (N_18469,N_18029,N_18187);
and U18470 (N_18470,N_18041,N_18023);
or U18471 (N_18471,N_18189,N_18051);
xnor U18472 (N_18472,N_18108,N_18100);
nor U18473 (N_18473,N_18014,N_18171);
or U18474 (N_18474,N_18188,N_18004);
or U18475 (N_18475,N_18095,N_18078);
and U18476 (N_18476,N_18102,N_18201);
xor U18477 (N_18477,N_18115,N_18131);
nand U18478 (N_18478,N_18063,N_18025);
nand U18479 (N_18479,N_18064,N_18214);
nand U18480 (N_18480,N_18090,N_18048);
or U18481 (N_18481,N_18141,N_18215);
or U18482 (N_18482,N_18200,N_18205);
nor U18483 (N_18483,N_18076,N_18200);
and U18484 (N_18484,N_18070,N_18215);
nor U18485 (N_18485,N_18233,N_18012);
nor U18486 (N_18486,N_18203,N_18043);
and U18487 (N_18487,N_18030,N_18227);
and U18488 (N_18488,N_18199,N_18065);
and U18489 (N_18489,N_18020,N_18088);
nor U18490 (N_18490,N_18084,N_18036);
and U18491 (N_18491,N_18124,N_18107);
nor U18492 (N_18492,N_18129,N_18064);
nor U18493 (N_18493,N_18144,N_18227);
and U18494 (N_18494,N_18214,N_18243);
nor U18495 (N_18495,N_18012,N_18040);
nor U18496 (N_18496,N_18207,N_18095);
nor U18497 (N_18497,N_18068,N_18204);
xor U18498 (N_18498,N_18057,N_18033);
and U18499 (N_18499,N_18052,N_18109);
nand U18500 (N_18500,N_18363,N_18331);
xor U18501 (N_18501,N_18268,N_18291);
nor U18502 (N_18502,N_18356,N_18479);
nand U18503 (N_18503,N_18279,N_18453);
nor U18504 (N_18504,N_18494,N_18354);
nor U18505 (N_18505,N_18409,N_18349);
or U18506 (N_18506,N_18469,N_18317);
nor U18507 (N_18507,N_18498,N_18250);
and U18508 (N_18508,N_18302,N_18486);
or U18509 (N_18509,N_18493,N_18490);
or U18510 (N_18510,N_18315,N_18402);
nand U18511 (N_18511,N_18377,N_18344);
and U18512 (N_18512,N_18254,N_18446);
nor U18513 (N_18513,N_18350,N_18466);
xor U18514 (N_18514,N_18467,N_18316);
xnor U18515 (N_18515,N_18267,N_18388);
nand U18516 (N_18516,N_18259,N_18472);
and U18517 (N_18517,N_18442,N_18357);
and U18518 (N_18518,N_18425,N_18367);
nor U18519 (N_18519,N_18386,N_18487);
nor U18520 (N_18520,N_18297,N_18435);
and U18521 (N_18521,N_18376,N_18491);
nor U18522 (N_18522,N_18318,N_18396);
and U18523 (N_18523,N_18445,N_18395);
or U18524 (N_18524,N_18265,N_18403);
nor U18525 (N_18525,N_18387,N_18275);
nand U18526 (N_18526,N_18366,N_18382);
nand U18527 (N_18527,N_18372,N_18443);
nand U18528 (N_18528,N_18251,N_18390);
or U18529 (N_18529,N_18285,N_18482);
nor U18530 (N_18530,N_18458,N_18408);
and U18531 (N_18531,N_18401,N_18459);
nand U18532 (N_18532,N_18394,N_18295);
or U18533 (N_18533,N_18389,N_18293);
xor U18534 (N_18534,N_18499,N_18457);
nor U18535 (N_18535,N_18264,N_18448);
or U18536 (N_18536,N_18370,N_18436);
and U18537 (N_18537,N_18263,N_18451);
and U18538 (N_18538,N_18447,N_18477);
and U18539 (N_18539,N_18280,N_18368);
and U18540 (N_18540,N_18299,N_18307);
nand U18541 (N_18541,N_18474,N_18450);
or U18542 (N_18542,N_18359,N_18369);
and U18543 (N_18543,N_18497,N_18257);
and U18544 (N_18544,N_18411,N_18489);
nor U18545 (N_18545,N_18320,N_18337);
nor U18546 (N_18546,N_18346,N_18405);
nor U18547 (N_18547,N_18439,N_18314);
or U18548 (N_18548,N_18277,N_18271);
and U18549 (N_18549,N_18471,N_18373);
or U18550 (N_18550,N_18294,N_18261);
nor U18551 (N_18551,N_18272,N_18422);
nor U18552 (N_18552,N_18292,N_18371);
nand U18553 (N_18553,N_18340,N_18381);
xor U18554 (N_18554,N_18461,N_18334);
nor U18555 (N_18555,N_18266,N_18400);
or U18556 (N_18556,N_18426,N_18290);
and U18557 (N_18557,N_18260,N_18470);
nor U18558 (N_18558,N_18270,N_18355);
and U18559 (N_18559,N_18454,N_18282);
nor U18560 (N_18560,N_18319,N_18335);
xnor U18561 (N_18561,N_18361,N_18485);
nand U18562 (N_18562,N_18488,N_18296);
or U18563 (N_18563,N_18385,N_18484);
or U18564 (N_18564,N_18300,N_18305);
or U18565 (N_18565,N_18420,N_18256);
nor U18566 (N_18566,N_18496,N_18347);
nor U18567 (N_18567,N_18364,N_18399);
or U18568 (N_18568,N_18417,N_18276);
xor U18569 (N_18569,N_18495,N_18433);
nor U18570 (N_18570,N_18283,N_18483);
or U18571 (N_18571,N_18413,N_18343);
and U18572 (N_18572,N_18427,N_18342);
and U18573 (N_18573,N_18456,N_18407);
or U18574 (N_18574,N_18353,N_18289);
xnor U18575 (N_18575,N_18406,N_18383);
nor U18576 (N_18576,N_18431,N_18336);
nor U18577 (N_18577,N_18330,N_18262);
nand U18578 (N_18578,N_18460,N_18480);
and U18579 (N_18579,N_18392,N_18324);
nand U18580 (N_18580,N_18288,N_18437);
nor U18581 (N_18581,N_18393,N_18312);
xnor U18582 (N_18582,N_18398,N_18306);
nand U18583 (N_18583,N_18284,N_18452);
or U18584 (N_18584,N_18255,N_18352);
and U18585 (N_18585,N_18360,N_18327);
xor U18586 (N_18586,N_18309,N_18419);
and U18587 (N_18587,N_18468,N_18478);
nand U18588 (N_18588,N_18310,N_18345);
and U18589 (N_18589,N_18323,N_18338);
nor U18590 (N_18590,N_18311,N_18434);
xor U18591 (N_18591,N_18326,N_18412);
or U18592 (N_18592,N_18430,N_18341);
nand U18593 (N_18593,N_18473,N_18463);
nor U18594 (N_18594,N_18333,N_18358);
nor U18595 (N_18595,N_18440,N_18438);
or U18596 (N_18596,N_18252,N_18415);
nor U18597 (N_18597,N_18339,N_18423);
and U18598 (N_18598,N_18432,N_18329);
and U18599 (N_18599,N_18384,N_18322);
or U18600 (N_18600,N_18418,N_18391);
and U18601 (N_18601,N_18428,N_18424);
nor U18602 (N_18602,N_18429,N_18313);
nor U18603 (N_18603,N_18278,N_18380);
or U18604 (N_18604,N_18301,N_18328);
xnor U18605 (N_18605,N_18374,N_18325);
nand U18606 (N_18606,N_18269,N_18379);
nand U18607 (N_18607,N_18375,N_18274);
or U18608 (N_18608,N_18287,N_18397);
nand U18609 (N_18609,N_18281,N_18308);
nand U18610 (N_18610,N_18286,N_18298);
nor U18611 (N_18611,N_18253,N_18378);
and U18612 (N_18612,N_18464,N_18441);
and U18613 (N_18613,N_18304,N_18475);
or U18614 (N_18614,N_18444,N_18365);
nand U18615 (N_18615,N_18414,N_18351);
nand U18616 (N_18616,N_18416,N_18332);
and U18617 (N_18617,N_18465,N_18462);
or U18618 (N_18618,N_18476,N_18273);
nand U18619 (N_18619,N_18449,N_18421);
and U18620 (N_18620,N_18303,N_18404);
xor U18621 (N_18621,N_18258,N_18410);
and U18622 (N_18622,N_18321,N_18455);
nand U18623 (N_18623,N_18492,N_18362);
nand U18624 (N_18624,N_18348,N_18481);
nand U18625 (N_18625,N_18346,N_18468);
or U18626 (N_18626,N_18293,N_18291);
and U18627 (N_18627,N_18496,N_18250);
xor U18628 (N_18628,N_18251,N_18345);
nor U18629 (N_18629,N_18359,N_18256);
nor U18630 (N_18630,N_18274,N_18499);
or U18631 (N_18631,N_18283,N_18353);
nand U18632 (N_18632,N_18369,N_18429);
nor U18633 (N_18633,N_18467,N_18485);
or U18634 (N_18634,N_18401,N_18363);
or U18635 (N_18635,N_18458,N_18378);
xnor U18636 (N_18636,N_18421,N_18433);
and U18637 (N_18637,N_18451,N_18403);
nor U18638 (N_18638,N_18430,N_18317);
or U18639 (N_18639,N_18341,N_18451);
nor U18640 (N_18640,N_18451,N_18356);
nand U18641 (N_18641,N_18266,N_18324);
or U18642 (N_18642,N_18264,N_18361);
and U18643 (N_18643,N_18426,N_18343);
nand U18644 (N_18644,N_18362,N_18450);
xnor U18645 (N_18645,N_18267,N_18404);
xnor U18646 (N_18646,N_18285,N_18255);
xnor U18647 (N_18647,N_18317,N_18439);
and U18648 (N_18648,N_18404,N_18353);
and U18649 (N_18649,N_18317,N_18435);
and U18650 (N_18650,N_18254,N_18337);
and U18651 (N_18651,N_18412,N_18421);
xnor U18652 (N_18652,N_18354,N_18265);
or U18653 (N_18653,N_18385,N_18279);
xor U18654 (N_18654,N_18271,N_18279);
nor U18655 (N_18655,N_18316,N_18411);
xnor U18656 (N_18656,N_18483,N_18300);
or U18657 (N_18657,N_18277,N_18478);
nor U18658 (N_18658,N_18411,N_18394);
nor U18659 (N_18659,N_18459,N_18446);
nand U18660 (N_18660,N_18273,N_18412);
or U18661 (N_18661,N_18422,N_18292);
and U18662 (N_18662,N_18309,N_18473);
nand U18663 (N_18663,N_18368,N_18372);
nand U18664 (N_18664,N_18375,N_18310);
and U18665 (N_18665,N_18298,N_18400);
xor U18666 (N_18666,N_18366,N_18438);
nand U18667 (N_18667,N_18361,N_18328);
nor U18668 (N_18668,N_18396,N_18427);
xor U18669 (N_18669,N_18419,N_18493);
or U18670 (N_18670,N_18433,N_18251);
and U18671 (N_18671,N_18307,N_18258);
or U18672 (N_18672,N_18435,N_18254);
xor U18673 (N_18673,N_18293,N_18440);
and U18674 (N_18674,N_18394,N_18441);
nor U18675 (N_18675,N_18339,N_18428);
and U18676 (N_18676,N_18307,N_18363);
or U18677 (N_18677,N_18461,N_18309);
or U18678 (N_18678,N_18327,N_18470);
nor U18679 (N_18679,N_18337,N_18353);
or U18680 (N_18680,N_18316,N_18297);
nor U18681 (N_18681,N_18396,N_18430);
or U18682 (N_18682,N_18341,N_18478);
nor U18683 (N_18683,N_18433,N_18338);
nand U18684 (N_18684,N_18314,N_18310);
nor U18685 (N_18685,N_18488,N_18427);
nand U18686 (N_18686,N_18377,N_18457);
nand U18687 (N_18687,N_18318,N_18468);
nor U18688 (N_18688,N_18479,N_18471);
and U18689 (N_18689,N_18265,N_18487);
nor U18690 (N_18690,N_18383,N_18497);
nor U18691 (N_18691,N_18433,N_18292);
nor U18692 (N_18692,N_18265,N_18479);
or U18693 (N_18693,N_18490,N_18458);
or U18694 (N_18694,N_18488,N_18476);
or U18695 (N_18695,N_18440,N_18273);
or U18696 (N_18696,N_18395,N_18444);
or U18697 (N_18697,N_18499,N_18407);
and U18698 (N_18698,N_18299,N_18424);
and U18699 (N_18699,N_18443,N_18409);
or U18700 (N_18700,N_18324,N_18435);
nor U18701 (N_18701,N_18391,N_18361);
xor U18702 (N_18702,N_18469,N_18483);
or U18703 (N_18703,N_18386,N_18373);
nand U18704 (N_18704,N_18364,N_18489);
nor U18705 (N_18705,N_18484,N_18374);
nor U18706 (N_18706,N_18388,N_18339);
and U18707 (N_18707,N_18266,N_18298);
nand U18708 (N_18708,N_18499,N_18476);
nand U18709 (N_18709,N_18486,N_18368);
nor U18710 (N_18710,N_18456,N_18290);
nor U18711 (N_18711,N_18282,N_18427);
nand U18712 (N_18712,N_18495,N_18318);
nand U18713 (N_18713,N_18322,N_18362);
or U18714 (N_18714,N_18293,N_18372);
or U18715 (N_18715,N_18298,N_18339);
nor U18716 (N_18716,N_18435,N_18255);
nand U18717 (N_18717,N_18255,N_18289);
nor U18718 (N_18718,N_18478,N_18412);
nor U18719 (N_18719,N_18486,N_18387);
and U18720 (N_18720,N_18325,N_18285);
nor U18721 (N_18721,N_18254,N_18352);
or U18722 (N_18722,N_18347,N_18276);
nand U18723 (N_18723,N_18438,N_18315);
nor U18724 (N_18724,N_18344,N_18396);
xor U18725 (N_18725,N_18446,N_18368);
and U18726 (N_18726,N_18324,N_18385);
and U18727 (N_18727,N_18448,N_18365);
nand U18728 (N_18728,N_18414,N_18261);
nand U18729 (N_18729,N_18324,N_18424);
and U18730 (N_18730,N_18286,N_18350);
nor U18731 (N_18731,N_18389,N_18490);
and U18732 (N_18732,N_18370,N_18266);
nor U18733 (N_18733,N_18299,N_18371);
or U18734 (N_18734,N_18432,N_18277);
nor U18735 (N_18735,N_18487,N_18266);
nor U18736 (N_18736,N_18258,N_18426);
xor U18737 (N_18737,N_18256,N_18375);
or U18738 (N_18738,N_18399,N_18323);
nor U18739 (N_18739,N_18328,N_18456);
and U18740 (N_18740,N_18442,N_18468);
and U18741 (N_18741,N_18356,N_18442);
or U18742 (N_18742,N_18478,N_18421);
and U18743 (N_18743,N_18382,N_18324);
and U18744 (N_18744,N_18425,N_18311);
and U18745 (N_18745,N_18388,N_18357);
and U18746 (N_18746,N_18362,N_18487);
and U18747 (N_18747,N_18323,N_18401);
nor U18748 (N_18748,N_18327,N_18371);
xor U18749 (N_18749,N_18327,N_18454);
and U18750 (N_18750,N_18715,N_18741);
nand U18751 (N_18751,N_18660,N_18706);
nor U18752 (N_18752,N_18724,N_18710);
or U18753 (N_18753,N_18620,N_18596);
or U18754 (N_18754,N_18569,N_18704);
nor U18755 (N_18755,N_18632,N_18636);
nand U18756 (N_18756,N_18644,N_18694);
nor U18757 (N_18757,N_18650,N_18717);
xor U18758 (N_18758,N_18568,N_18647);
or U18759 (N_18759,N_18581,N_18624);
nor U18760 (N_18760,N_18504,N_18690);
nand U18761 (N_18761,N_18517,N_18551);
and U18762 (N_18762,N_18676,N_18668);
xnor U18763 (N_18763,N_18548,N_18610);
nor U18764 (N_18764,N_18574,N_18746);
and U18765 (N_18765,N_18714,N_18728);
or U18766 (N_18766,N_18567,N_18540);
or U18767 (N_18767,N_18508,N_18611);
nor U18768 (N_18768,N_18723,N_18661);
xnor U18769 (N_18769,N_18643,N_18675);
or U18770 (N_18770,N_18555,N_18701);
or U18771 (N_18771,N_18747,N_18580);
nand U18772 (N_18772,N_18594,N_18640);
nor U18773 (N_18773,N_18545,N_18565);
nand U18774 (N_18774,N_18615,N_18516);
nand U18775 (N_18775,N_18633,N_18674);
nand U18776 (N_18776,N_18634,N_18539);
and U18777 (N_18777,N_18659,N_18595);
xnor U18778 (N_18778,N_18607,N_18500);
nor U18779 (N_18779,N_18708,N_18657);
nor U18780 (N_18780,N_18671,N_18656);
or U18781 (N_18781,N_18572,N_18592);
nor U18782 (N_18782,N_18652,N_18679);
xnor U18783 (N_18783,N_18625,N_18550);
and U18784 (N_18784,N_18692,N_18522);
nor U18785 (N_18785,N_18547,N_18685);
and U18786 (N_18786,N_18651,N_18618);
or U18787 (N_18787,N_18556,N_18716);
nand U18788 (N_18788,N_18506,N_18672);
or U18789 (N_18789,N_18510,N_18546);
nand U18790 (N_18790,N_18501,N_18740);
xnor U18791 (N_18791,N_18721,N_18518);
nand U18792 (N_18792,N_18537,N_18609);
or U18793 (N_18793,N_18649,N_18626);
nand U18794 (N_18794,N_18613,N_18505);
and U18795 (N_18795,N_18738,N_18635);
or U18796 (N_18796,N_18532,N_18523);
nand U18797 (N_18797,N_18667,N_18709);
nor U18798 (N_18798,N_18673,N_18515);
nand U18799 (N_18799,N_18733,N_18684);
nand U18800 (N_18800,N_18639,N_18621);
and U18801 (N_18801,N_18564,N_18648);
nor U18802 (N_18802,N_18503,N_18511);
xnor U18803 (N_18803,N_18641,N_18599);
or U18804 (N_18804,N_18662,N_18588);
and U18805 (N_18805,N_18622,N_18585);
nand U18806 (N_18806,N_18554,N_18749);
or U18807 (N_18807,N_18642,N_18552);
or U18808 (N_18808,N_18605,N_18597);
nor U18809 (N_18809,N_18557,N_18521);
nand U18810 (N_18810,N_18587,N_18720);
nor U18811 (N_18811,N_18654,N_18589);
and U18812 (N_18812,N_18570,N_18735);
and U18813 (N_18813,N_18655,N_18602);
nor U18814 (N_18814,N_18616,N_18682);
or U18815 (N_18815,N_18719,N_18743);
xor U18816 (N_18816,N_18584,N_18577);
and U18817 (N_18817,N_18600,N_18653);
nand U18818 (N_18818,N_18691,N_18663);
nand U18819 (N_18819,N_18543,N_18628);
nand U18820 (N_18820,N_18512,N_18737);
and U18821 (N_18821,N_18705,N_18680);
nor U18822 (N_18822,N_18559,N_18617);
nor U18823 (N_18823,N_18700,N_18612);
and U18824 (N_18824,N_18534,N_18645);
nand U18825 (N_18825,N_18703,N_18713);
xor U18826 (N_18826,N_18528,N_18677);
nand U18827 (N_18827,N_18695,N_18542);
nor U18828 (N_18828,N_18718,N_18524);
nor U18829 (N_18829,N_18502,N_18688);
and U18830 (N_18830,N_18711,N_18725);
xor U18831 (N_18831,N_18614,N_18604);
nand U18832 (N_18832,N_18519,N_18726);
xnor U18833 (N_18833,N_18527,N_18686);
and U18834 (N_18834,N_18665,N_18520);
nand U18835 (N_18835,N_18683,N_18514);
nand U18836 (N_18836,N_18729,N_18526);
nand U18837 (N_18837,N_18608,N_18730);
or U18838 (N_18838,N_18707,N_18558);
xnor U18839 (N_18839,N_18638,N_18727);
or U18840 (N_18840,N_18531,N_18541);
nand U18841 (N_18841,N_18593,N_18582);
nand U18842 (N_18842,N_18576,N_18549);
nor U18843 (N_18843,N_18678,N_18731);
or U18844 (N_18844,N_18578,N_18579);
xor U18845 (N_18845,N_18509,N_18533);
xnor U18846 (N_18846,N_18734,N_18560);
and U18847 (N_18847,N_18525,N_18748);
nand U18848 (N_18848,N_18536,N_18669);
nor U18849 (N_18849,N_18631,N_18629);
and U18850 (N_18850,N_18699,N_18736);
nand U18851 (N_18851,N_18666,N_18658);
nor U18852 (N_18852,N_18619,N_18646);
nand U18853 (N_18853,N_18732,N_18689);
or U18854 (N_18854,N_18606,N_18571);
or U18855 (N_18855,N_18681,N_18697);
and U18856 (N_18856,N_18507,N_18553);
and U18857 (N_18857,N_18598,N_18575);
nand U18858 (N_18858,N_18603,N_18573);
or U18859 (N_18859,N_18583,N_18529);
and U18860 (N_18860,N_18693,N_18530);
xor U18861 (N_18861,N_18590,N_18712);
nand U18862 (N_18862,N_18586,N_18601);
xnor U18863 (N_18863,N_18744,N_18563);
or U18864 (N_18864,N_18623,N_18630);
nor U18865 (N_18865,N_18544,N_18742);
and U18866 (N_18866,N_18739,N_18670);
nand U18867 (N_18867,N_18637,N_18745);
and U18868 (N_18868,N_18664,N_18702);
and U18869 (N_18869,N_18561,N_18566);
and U18870 (N_18870,N_18687,N_18538);
or U18871 (N_18871,N_18591,N_18627);
or U18872 (N_18872,N_18562,N_18535);
and U18873 (N_18873,N_18513,N_18698);
and U18874 (N_18874,N_18696,N_18722);
nor U18875 (N_18875,N_18551,N_18655);
or U18876 (N_18876,N_18598,N_18619);
and U18877 (N_18877,N_18525,N_18705);
or U18878 (N_18878,N_18562,N_18602);
nand U18879 (N_18879,N_18689,N_18532);
and U18880 (N_18880,N_18657,N_18696);
nor U18881 (N_18881,N_18646,N_18565);
xor U18882 (N_18882,N_18733,N_18691);
nand U18883 (N_18883,N_18737,N_18618);
nand U18884 (N_18884,N_18575,N_18729);
xor U18885 (N_18885,N_18699,N_18530);
nand U18886 (N_18886,N_18670,N_18708);
nand U18887 (N_18887,N_18647,N_18560);
nand U18888 (N_18888,N_18717,N_18748);
nor U18889 (N_18889,N_18505,N_18661);
nor U18890 (N_18890,N_18714,N_18556);
nor U18891 (N_18891,N_18705,N_18650);
or U18892 (N_18892,N_18568,N_18632);
nand U18893 (N_18893,N_18589,N_18536);
nor U18894 (N_18894,N_18574,N_18623);
or U18895 (N_18895,N_18576,N_18736);
and U18896 (N_18896,N_18650,N_18548);
nor U18897 (N_18897,N_18690,N_18525);
nor U18898 (N_18898,N_18741,N_18534);
and U18899 (N_18899,N_18537,N_18559);
or U18900 (N_18900,N_18643,N_18713);
or U18901 (N_18901,N_18627,N_18553);
or U18902 (N_18902,N_18548,N_18667);
or U18903 (N_18903,N_18513,N_18510);
nor U18904 (N_18904,N_18524,N_18512);
nor U18905 (N_18905,N_18612,N_18692);
or U18906 (N_18906,N_18549,N_18503);
nand U18907 (N_18907,N_18577,N_18511);
or U18908 (N_18908,N_18612,N_18544);
and U18909 (N_18909,N_18587,N_18706);
or U18910 (N_18910,N_18682,N_18643);
nand U18911 (N_18911,N_18516,N_18601);
nand U18912 (N_18912,N_18669,N_18630);
nor U18913 (N_18913,N_18530,N_18687);
and U18914 (N_18914,N_18508,N_18610);
nor U18915 (N_18915,N_18525,N_18731);
and U18916 (N_18916,N_18654,N_18743);
nor U18917 (N_18917,N_18712,N_18560);
or U18918 (N_18918,N_18573,N_18703);
nand U18919 (N_18919,N_18505,N_18527);
and U18920 (N_18920,N_18509,N_18535);
nand U18921 (N_18921,N_18533,N_18536);
nand U18922 (N_18922,N_18723,N_18658);
and U18923 (N_18923,N_18539,N_18628);
and U18924 (N_18924,N_18676,N_18709);
and U18925 (N_18925,N_18615,N_18704);
and U18926 (N_18926,N_18638,N_18677);
and U18927 (N_18927,N_18563,N_18659);
nand U18928 (N_18928,N_18608,N_18726);
nor U18929 (N_18929,N_18733,N_18742);
or U18930 (N_18930,N_18575,N_18749);
nand U18931 (N_18931,N_18721,N_18591);
nand U18932 (N_18932,N_18560,N_18604);
and U18933 (N_18933,N_18531,N_18630);
and U18934 (N_18934,N_18704,N_18617);
or U18935 (N_18935,N_18630,N_18617);
and U18936 (N_18936,N_18698,N_18697);
nor U18937 (N_18937,N_18632,N_18578);
and U18938 (N_18938,N_18547,N_18648);
nor U18939 (N_18939,N_18703,N_18665);
or U18940 (N_18940,N_18600,N_18695);
xor U18941 (N_18941,N_18654,N_18602);
nor U18942 (N_18942,N_18594,N_18688);
and U18943 (N_18943,N_18693,N_18578);
nor U18944 (N_18944,N_18585,N_18558);
nand U18945 (N_18945,N_18716,N_18720);
nor U18946 (N_18946,N_18630,N_18663);
or U18947 (N_18947,N_18597,N_18623);
and U18948 (N_18948,N_18694,N_18527);
xnor U18949 (N_18949,N_18609,N_18668);
nor U18950 (N_18950,N_18640,N_18539);
and U18951 (N_18951,N_18737,N_18579);
and U18952 (N_18952,N_18712,N_18624);
xor U18953 (N_18953,N_18648,N_18722);
nand U18954 (N_18954,N_18712,N_18703);
or U18955 (N_18955,N_18567,N_18506);
or U18956 (N_18956,N_18702,N_18501);
and U18957 (N_18957,N_18724,N_18514);
nand U18958 (N_18958,N_18650,N_18711);
nor U18959 (N_18959,N_18502,N_18692);
and U18960 (N_18960,N_18530,N_18653);
or U18961 (N_18961,N_18540,N_18616);
nor U18962 (N_18962,N_18641,N_18622);
nand U18963 (N_18963,N_18739,N_18715);
and U18964 (N_18964,N_18708,N_18665);
or U18965 (N_18965,N_18637,N_18748);
xor U18966 (N_18966,N_18652,N_18654);
or U18967 (N_18967,N_18698,N_18500);
or U18968 (N_18968,N_18584,N_18651);
or U18969 (N_18969,N_18654,N_18747);
or U18970 (N_18970,N_18741,N_18692);
and U18971 (N_18971,N_18747,N_18676);
nor U18972 (N_18972,N_18712,N_18584);
and U18973 (N_18973,N_18557,N_18744);
or U18974 (N_18974,N_18644,N_18728);
nand U18975 (N_18975,N_18645,N_18529);
and U18976 (N_18976,N_18538,N_18571);
and U18977 (N_18977,N_18723,N_18589);
nand U18978 (N_18978,N_18529,N_18676);
nand U18979 (N_18979,N_18738,N_18545);
or U18980 (N_18980,N_18676,N_18607);
nand U18981 (N_18981,N_18689,N_18525);
nor U18982 (N_18982,N_18705,N_18727);
or U18983 (N_18983,N_18604,N_18629);
nor U18984 (N_18984,N_18594,N_18577);
or U18985 (N_18985,N_18629,N_18630);
nand U18986 (N_18986,N_18625,N_18636);
xor U18987 (N_18987,N_18568,N_18738);
and U18988 (N_18988,N_18654,N_18551);
or U18989 (N_18989,N_18571,N_18618);
nor U18990 (N_18990,N_18630,N_18590);
and U18991 (N_18991,N_18661,N_18589);
and U18992 (N_18992,N_18703,N_18578);
or U18993 (N_18993,N_18593,N_18680);
or U18994 (N_18994,N_18525,N_18577);
nand U18995 (N_18995,N_18535,N_18710);
nor U18996 (N_18996,N_18543,N_18721);
nor U18997 (N_18997,N_18715,N_18682);
and U18998 (N_18998,N_18739,N_18561);
or U18999 (N_18999,N_18599,N_18564);
or U19000 (N_19000,N_18962,N_18837);
and U19001 (N_19001,N_18860,N_18864);
nand U19002 (N_19002,N_18768,N_18957);
nor U19003 (N_19003,N_18903,N_18914);
nand U19004 (N_19004,N_18956,N_18806);
nand U19005 (N_19005,N_18867,N_18835);
xnor U19006 (N_19006,N_18763,N_18881);
or U19007 (N_19007,N_18930,N_18898);
nand U19008 (N_19008,N_18868,N_18983);
or U19009 (N_19009,N_18890,N_18945);
and U19010 (N_19010,N_18911,N_18841);
nand U19011 (N_19011,N_18821,N_18793);
or U19012 (N_19012,N_18838,N_18882);
nor U19013 (N_19013,N_18862,N_18985);
or U19014 (N_19014,N_18847,N_18842);
or U19015 (N_19015,N_18978,N_18873);
nor U19016 (N_19016,N_18980,N_18974);
and U19017 (N_19017,N_18917,N_18807);
or U19018 (N_19018,N_18839,N_18755);
or U19019 (N_19019,N_18822,N_18887);
nand U19020 (N_19020,N_18846,N_18958);
and U19021 (N_19021,N_18815,N_18893);
nor U19022 (N_19022,N_18984,N_18961);
nand U19023 (N_19023,N_18801,N_18830);
nand U19024 (N_19024,N_18943,N_18912);
and U19025 (N_19025,N_18762,N_18900);
nand U19026 (N_19026,N_18992,N_18771);
nand U19027 (N_19027,N_18963,N_18781);
nor U19028 (N_19028,N_18902,N_18858);
and U19029 (N_19029,N_18937,N_18895);
or U19030 (N_19030,N_18897,N_18832);
nor U19031 (N_19031,N_18805,N_18971);
xnor U19032 (N_19032,N_18855,N_18975);
xnor U19033 (N_19033,N_18901,N_18852);
nor U19034 (N_19034,N_18758,N_18828);
xnor U19035 (N_19035,N_18787,N_18936);
nand U19036 (N_19036,N_18986,N_18918);
xnor U19037 (N_19037,N_18996,N_18848);
or U19038 (N_19038,N_18889,N_18764);
and U19039 (N_19039,N_18818,N_18861);
and U19040 (N_19040,N_18891,N_18924);
or U19041 (N_19041,N_18790,N_18761);
and U19042 (N_19042,N_18977,N_18817);
nor U19043 (N_19043,N_18849,N_18976);
nor U19044 (N_19044,N_18944,N_18916);
and U19045 (N_19045,N_18997,N_18925);
and U19046 (N_19046,N_18913,N_18833);
and U19047 (N_19047,N_18788,N_18759);
xnor U19048 (N_19048,N_18797,N_18998);
xor U19049 (N_19049,N_18757,N_18774);
nor U19050 (N_19050,N_18791,N_18987);
nand U19051 (N_19051,N_18922,N_18959);
and U19052 (N_19052,N_18840,N_18967);
nor U19053 (N_19053,N_18792,N_18954);
nand U19054 (N_19054,N_18784,N_18823);
and U19055 (N_19055,N_18753,N_18926);
and U19056 (N_19056,N_18874,N_18777);
xnor U19057 (N_19057,N_18907,N_18814);
or U19058 (N_19058,N_18994,N_18779);
nand U19059 (N_19059,N_18804,N_18851);
and U19060 (N_19060,N_18871,N_18919);
nand U19061 (N_19061,N_18812,N_18942);
or U19062 (N_19062,N_18827,N_18766);
and U19063 (N_19063,N_18915,N_18960);
xor U19064 (N_19064,N_18780,N_18866);
and U19065 (N_19065,N_18775,N_18949);
and U19066 (N_19066,N_18770,N_18968);
or U19067 (N_19067,N_18786,N_18896);
nor U19068 (N_19068,N_18934,N_18773);
nand U19069 (N_19069,N_18908,N_18836);
and U19070 (N_19070,N_18878,N_18798);
and U19071 (N_19071,N_18938,N_18850);
nor U19072 (N_19072,N_18950,N_18865);
nor U19073 (N_19073,N_18880,N_18800);
and U19074 (N_19074,N_18816,N_18795);
nand U19075 (N_19075,N_18776,N_18785);
nor U19076 (N_19076,N_18857,N_18813);
or U19077 (N_19077,N_18988,N_18808);
nand U19078 (N_19078,N_18905,N_18935);
xor U19079 (N_19079,N_18966,N_18810);
nand U19080 (N_19080,N_18826,N_18820);
or U19081 (N_19081,N_18760,N_18991);
xor U19082 (N_19082,N_18769,N_18802);
nor U19083 (N_19083,N_18778,N_18829);
and U19084 (N_19084,N_18927,N_18932);
and U19085 (N_19085,N_18892,N_18794);
and U19086 (N_19086,N_18854,N_18824);
nand U19087 (N_19087,N_18767,N_18969);
or U19088 (N_19088,N_18894,N_18789);
or U19089 (N_19089,N_18904,N_18843);
nor U19090 (N_19090,N_18884,N_18948);
and U19091 (N_19091,N_18990,N_18796);
nand U19092 (N_19092,N_18899,N_18947);
or U19093 (N_19093,N_18886,N_18799);
nand U19094 (N_19094,N_18946,N_18853);
and U19095 (N_19095,N_18982,N_18993);
or U19096 (N_19096,N_18750,N_18970);
or U19097 (N_19097,N_18951,N_18885);
and U19098 (N_19098,N_18856,N_18844);
and U19099 (N_19099,N_18909,N_18964);
nand U19100 (N_19100,N_18923,N_18863);
nand U19101 (N_19101,N_18952,N_18955);
or U19102 (N_19102,N_18933,N_18869);
and U19103 (N_19103,N_18809,N_18831);
and U19104 (N_19104,N_18941,N_18859);
nor U19105 (N_19105,N_18883,N_18877);
nand U19106 (N_19106,N_18876,N_18995);
nand U19107 (N_19107,N_18929,N_18765);
and U19108 (N_19108,N_18965,N_18920);
and U19109 (N_19109,N_18875,N_18756);
xor U19110 (N_19110,N_18953,N_18973);
and U19111 (N_19111,N_18979,N_18888);
and U19112 (N_19112,N_18783,N_18752);
and U19113 (N_19113,N_18921,N_18845);
and U19114 (N_19114,N_18834,N_18906);
or U19115 (N_19115,N_18811,N_18870);
or U19116 (N_19116,N_18910,N_18772);
or U19117 (N_19117,N_18999,N_18782);
or U19118 (N_19118,N_18981,N_18972);
nor U19119 (N_19119,N_18819,N_18939);
nor U19120 (N_19120,N_18989,N_18879);
and U19121 (N_19121,N_18940,N_18754);
nand U19122 (N_19122,N_18931,N_18825);
and U19123 (N_19123,N_18928,N_18751);
or U19124 (N_19124,N_18872,N_18803);
nand U19125 (N_19125,N_18814,N_18846);
and U19126 (N_19126,N_18895,N_18876);
or U19127 (N_19127,N_18787,N_18824);
or U19128 (N_19128,N_18825,N_18764);
and U19129 (N_19129,N_18895,N_18977);
or U19130 (N_19130,N_18968,N_18963);
or U19131 (N_19131,N_18887,N_18844);
xnor U19132 (N_19132,N_18929,N_18805);
nand U19133 (N_19133,N_18934,N_18816);
nand U19134 (N_19134,N_18812,N_18816);
nand U19135 (N_19135,N_18807,N_18866);
nor U19136 (N_19136,N_18837,N_18847);
or U19137 (N_19137,N_18849,N_18867);
nand U19138 (N_19138,N_18940,N_18865);
nor U19139 (N_19139,N_18876,N_18769);
or U19140 (N_19140,N_18974,N_18997);
or U19141 (N_19141,N_18879,N_18845);
or U19142 (N_19142,N_18857,N_18940);
nand U19143 (N_19143,N_18771,N_18764);
or U19144 (N_19144,N_18760,N_18891);
nand U19145 (N_19145,N_18958,N_18971);
and U19146 (N_19146,N_18978,N_18770);
nand U19147 (N_19147,N_18903,N_18980);
nand U19148 (N_19148,N_18779,N_18773);
and U19149 (N_19149,N_18885,N_18961);
or U19150 (N_19150,N_18864,N_18960);
or U19151 (N_19151,N_18824,N_18995);
or U19152 (N_19152,N_18904,N_18811);
nor U19153 (N_19153,N_18923,N_18887);
or U19154 (N_19154,N_18801,N_18775);
or U19155 (N_19155,N_18756,N_18939);
or U19156 (N_19156,N_18987,N_18976);
or U19157 (N_19157,N_18911,N_18880);
nor U19158 (N_19158,N_18832,N_18947);
xor U19159 (N_19159,N_18888,N_18919);
nor U19160 (N_19160,N_18830,N_18937);
nor U19161 (N_19161,N_18861,N_18830);
nor U19162 (N_19162,N_18848,N_18821);
and U19163 (N_19163,N_18912,N_18866);
and U19164 (N_19164,N_18795,N_18857);
and U19165 (N_19165,N_18803,N_18751);
and U19166 (N_19166,N_18766,N_18881);
nand U19167 (N_19167,N_18769,N_18804);
nor U19168 (N_19168,N_18948,N_18964);
or U19169 (N_19169,N_18803,N_18991);
or U19170 (N_19170,N_18864,N_18893);
nand U19171 (N_19171,N_18980,N_18826);
nand U19172 (N_19172,N_18976,N_18959);
nor U19173 (N_19173,N_18891,N_18906);
and U19174 (N_19174,N_18900,N_18985);
nand U19175 (N_19175,N_18771,N_18782);
or U19176 (N_19176,N_18750,N_18751);
or U19177 (N_19177,N_18990,N_18854);
xor U19178 (N_19178,N_18910,N_18996);
or U19179 (N_19179,N_18783,N_18911);
or U19180 (N_19180,N_18854,N_18846);
and U19181 (N_19181,N_18971,N_18930);
nor U19182 (N_19182,N_18834,N_18840);
nand U19183 (N_19183,N_18864,N_18771);
nor U19184 (N_19184,N_18882,N_18868);
or U19185 (N_19185,N_18770,N_18916);
or U19186 (N_19186,N_18800,N_18753);
nand U19187 (N_19187,N_18844,N_18764);
or U19188 (N_19188,N_18976,N_18891);
or U19189 (N_19189,N_18889,N_18897);
nor U19190 (N_19190,N_18838,N_18906);
xor U19191 (N_19191,N_18755,N_18771);
and U19192 (N_19192,N_18802,N_18799);
nor U19193 (N_19193,N_18773,N_18899);
and U19194 (N_19194,N_18805,N_18785);
or U19195 (N_19195,N_18954,N_18883);
nand U19196 (N_19196,N_18860,N_18962);
nor U19197 (N_19197,N_18975,N_18802);
and U19198 (N_19198,N_18862,N_18785);
xnor U19199 (N_19199,N_18987,N_18890);
nand U19200 (N_19200,N_18926,N_18834);
nand U19201 (N_19201,N_18841,N_18854);
and U19202 (N_19202,N_18830,N_18762);
nor U19203 (N_19203,N_18910,N_18964);
nor U19204 (N_19204,N_18975,N_18814);
or U19205 (N_19205,N_18830,N_18921);
and U19206 (N_19206,N_18945,N_18967);
or U19207 (N_19207,N_18916,N_18852);
and U19208 (N_19208,N_18798,N_18773);
nor U19209 (N_19209,N_18873,N_18869);
and U19210 (N_19210,N_18777,N_18828);
and U19211 (N_19211,N_18940,N_18917);
or U19212 (N_19212,N_18771,N_18944);
or U19213 (N_19213,N_18770,N_18778);
nand U19214 (N_19214,N_18979,N_18801);
and U19215 (N_19215,N_18921,N_18970);
and U19216 (N_19216,N_18795,N_18751);
nor U19217 (N_19217,N_18970,N_18763);
nor U19218 (N_19218,N_18959,N_18991);
nand U19219 (N_19219,N_18823,N_18921);
or U19220 (N_19220,N_18857,N_18787);
and U19221 (N_19221,N_18837,N_18956);
xor U19222 (N_19222,N_18975,N_18844);
nor U19223 (N_19223,N_18806,N_18953);
and U19224 (N_19224,N_18955,N_18919);
nand U19225 (N_19225,N_18924,N_18920);
nand U19226 (N_19226,N_18820,N_18825);
or U19227 (N_19227,N_18966,N_18793);
nand U19228 (N_19228,N_18782,N_18817);
nand U19229 (N_19229,N_18846,N_18961);
and U19230 (N_19230,N_18922,N_18931);
nand U19231 (N_19231,N_18909,N_18860);
nor U19232 (N_19232,N_18824,N_18860);
nor U19233 (N_19233,N_18992,N_18922);
nor U19234 (N_19234,N_18973,N_18962);
nand U19235 (N_19235,N_18995,N_18804);
or U19236 (N_19236,N_18827,N_18772);
or U19237 (N_19237,N_18962,N_18854);
nor U19238 (N_19238,N_18952,N_18957);
and U19239 (N_19239,N_18945,N_18782);
or U19240 (N_19240,N_18761,N_18944);
nor U19241 (N_19241,N_18972,N_18827);
nor U19242 (N_19242,N_18854,N_18830);
and U19243 (N_19243,N_18805,N_18813);
or U19244 (N_19244,N_18793,N_18803);
or U19245 (N_19245,N_18865,N_18766);
nand U19246 (N_19246,N_18980,N_18976);
xnor U19247 (N_19247,N_18837,N_18934);
nand U19248 (N_19248,N_18969,N_18945);
or U19249 (N_19249,N_18751,N_18932);
nand U19250 (N_19250,N_19170,N_19158);
nor U19251 (N_19251,N_19069,N_19146);
xnor U19252 (N_19252,N_19238,N_19172);
nor U19253 (N_19253,N_19211,N_19067);
or U19254 (N_19254,N_19034,N_19151);
nand U19255 (N_19255,N_19056,N_19131);
or U19256 (N_19256,N_19096,N_19047);
nand U19257 (N_19257,N_19048,N_19176);
nor U19258 (N_19258,N_19178,N_19104);
or U19259 (N_19259,N_19013,N_19006);
nor U19260 (N_19260,N_19156,N_19198);
and U19261 (N_19261,N_19208,N_19074);
nand U19262 (N_19262,N_19194,N_19025);
nand U19263 (N_19263,N_19183,N_19210);
and U19264 (N_19264,N_19168,N_19177);
and U19265 (N_19265,N_19139,N_19209);
and U19266 (N_19266,N_19097,N_19231);
nand U19267 (N_19267,N_19041,N_19027);
xnor U19268 (N_19268,N_19164,N_19108);
xnor U19269 (N_19269,N_19123,N_19112);
nand U19270 (N_19270,N_19109,N_19053);
nor U19271 (N_19271,N_19125,N_19229);
and U19272 (N_19272,N_19161,N_19024);
or U19273 (N_19273,N_19003,N_19050);
xnor U19274 (N_19274,N_19145,N_19026);
and U19275 (N_19275,N_19187,N_19245);
and U19276 (N_19276,N_19110,N_19102);
and U19277 (N_19277,N_19002,N_19084);
xor U19278 (N_19278,N_19230,N_19153);
xor U19279 (N_19279,N_19023,N_19241);
and U19280 (N_19280,N_19031,N_19220);
and U19281 (N_19281,N_19179,N_19132);
nor U19282 (N_19282,N_19243,N_19080);
nand U19283 (N_19283,N_19160,N_19149);
nand U19284 (N_19284,N_19045,N_19181);
nor U19285 (N_19285,N_19219,N_19009);
and U19286 (N_19286,N_19166,N_19234);
nor U19287 (N_19287,N_19068,N_19094);
nand U19288 (N_19288,N_19205,N_19138);
and U19289 (N_19289,N_19144,N_19193);
or U19290 (N_19290,N_19196,N_19165);
nand U19291 (N_19291,N_19235,N_19036);
and U19292 (N_19292,N_19117,N_19140);
and U19293 (N_19293,N_19182,N_19055);
nor U19294 (N_19294,N_19022,N_19215);
xnor U19295 (N_19295,N_19197,N_19174);
or U19296 (N_19296,N_19044,N_19118);
xnor U19297 (N_19297,N_19103,N_19248);
xnor U19298 (N_19298,N_19119,N_19085);
and U19299 (N_19299,N_19092,N_19099);
or U19300 (N_19300,N_19224,N_19037);
and U19301 (N_19301,N_19116,N_19206);
xnor U19302 (N_19302,N_19163,N_19191);
or U19303 (N_19303,N_19076,N_19126);
or U19304 (N_19304,N_19066,N_19190);
nor U19305 (N_19305,N_19042,N_19061);
nor U19306 (N_19306,N_19054,N_19073);
nand U19307 (N_19307,N_19071,N_19000);
nor U19308 (N_19308,N_19012,N_19011);
or U19309 (N_19309,N_19095,N_19154);
and U19310 (N_19310,N_19184,N_19088);
nand U19311 (N_19311,N_19155,N_19098);
xor U19312 (N_19312,N_19083,N_19033);
and U19313 (N_19313,N_19028,N_19049);
and U19314 (N_19314,N_19030,N_19032);
and U19315 (N_19315,N_19135,N_19005);
nand U19316 (N_19316,N_19058,N_19090);
xor U19317 (N_19317,N_19019,N_19147);
nor U19318 (N_19318,N_19226,N_19100);
and U19319 (N_19319,N_19192,N_19065);
nand U19320 (N_19320,N_19222,N_19015);
nand U19321 (N_19321,N_19203,N_19200);
and U19322 (N_19322,N_19150,N_19249);
nor U19323 (N_19323,N_19244,N_19081);
or U19324 (N_19324,N_19039,N_19010);
nor U19325 (N_19325,N_19225,N_19130);
or U19326 (N_19326,N_19242,N_19101);
or U19327 (N_19327,N_19121,N_19070);
nor U19328 (N_19328,N_19082,N_19223);
nand U19329 (N_19329,N_19029,N_19152);
and U19330 (N_19330,N_19133,N_19207);
nand U19331 (N_19331,N_19228,N_19046);
and U19332 (N_19332,N_19122,N_19239);
nand U19333 (N_19333,N_19077,N_19114);
nand U19334 (N_19334,N_19051,N_19062);
and U19335 (N_19335,N_19201,N_19246);
nor U19336 (N_19336,N_19204,N_19093);
and U19337 (N_19337,N_19004,N_19129);
or U19338 (N_19338,N_19162,N_19087);
nand U19339 (N_19339,N_19064,N_19079);
nand U19340 (N_19340,N_19169,N_19137);
nand U19341 (N_19341,N_19008,N_19141);
or U19342 (N_19342,N_19038,N_19236);
nor U19343 (N_19343,N_19186,N_19035);
xor U19344 (N_19344,N_19159,N_19021);
nand U19345 (N_19345,N_19189,N_19040);
xnor U19346 (N_19346,N_19173,N_19167);
or U19347 (N_19347,N_19227,N_19124);
nand U19348 (N_19348,N_19142,N_19195);
nor U19349 (N_19349,N_19202,N_19217);
and U19350 (N_19350,N_19240,N_19134);
or U19351 (N_19351,N_19001,N_19188);
nand U19352 (N_19352,N_19016,N_19106);
nor U19353 (N_19353,N_19237,N_19214);
and U19354 (N_19354,N_19136,N_19089);
nand U19355 (N_19355,N_19014,N_19143);
nor U19356 (N_19356,N_19247,N_19128);
and U19357 (N_19357,N_19075,N_19111);
xnor U19358 (N_19358,N_19043,N_19180);
nor U19359 (N_19359,N_19020,N_19059);
and U19360 (N_19360,N_19086,N_19199);
nor U19361 (N_19361,N_19221,N_19213);
or U19362 (N_19362,N_19091,N_19171);
and U19363 (N_19363,N_19052,N_19185);
and U19364 (N_19364,N_19120,N_19212);
nand U19365 (N_19365,N_19233,N_19078);
and U19366 (N_19366,N_19218,N_19007);
nor U19367 (N_19367,N_19157,N_19072);
xnor U19368 (N_19368,N_19017,N_19018);
nand U19369 (N_19369,N_19216,N_19115);
nor U19370 (N_19370,N_19105,N_19113);
nand U19371 (N_19371,N_19107,N_19057);
and U19372 (N_19372,N_19060,N_19063);
nor U19373 (N_19373,N_19175,N_19148);
nand U19374 (N_19374,N_19127,N_19232);
and U19375 (N_19375,N_19135,N_19028);
nor U19376 (N_19376,N_19026,N_19078);
nor U19377 (N_19377,N_19091,N_19240);
or U19378 (N_19378,N_19119,N_19014);
nand U19379 (N_19379,N_19067,N_19146);
nor U19380 (N_19380,N_19223,N_19154);
and U19381 (N_19381,N_19196,N_19144);
nand U19382 (N_19382,N_19199,N_19214);
nand U19383 (N_19383,N_19232,N_19064);
xnor U19384 (N_19384,N_19025,N_19044);
nor U19385 (N_19385,N_19142,N_19182);
or U19386 (N_19386,N_19084,N_19211);
nor U19387 (N_19387,N_19076,N_19094);
or U19388 (N_19388,N_19215,N_19180);
and U19389 (N_19389,N_19158,N_19215);
xor U19390 (N_19390,N_19155,N_19047);
and U19391 (N_19391,N_19090,N_19092);
nand U19392 (N_19392,N_19082,N_19081);
and U19393 (N_19393,N_19019,N_19081);
and U19394 (N_19394,N_19002,N_19020);
nand U19395 (N_19395,N_19083,N_19114);
and U19396 (N_19396,N_19051,N_19209);
nand U19397 (N_19397,N_19082,N_19066);
and U19398 (N_19398,N_19226,N_19085);
and U19399 (N_19399,N_19221,N_19147);
nor U19400 (N_19400,N_19157,N_19010);
and U19401 (N_19401,N_19152,N_19067);
and U19402 (N_19402,N_19226,N_19192);
nor U19403 (N_19403,N_19225,N_19144);
or U19404 (N_19404,N_19176,N_19242);
nor U19405 (N_19405,N_19242,N_19245);
and U19406 (N_19406,N_19118,N_19060);
or U19407 (N_19407,N_19054,N_19122);
and U19408 (N_19408,N_19107,N_19023);
nor U19409 (N_19409,N_19035,N_19094);
or U19410 (N_19410,N_19099,N_19037);
or U19411 (N_19411,N_19135,N_19237);
nor U19412 (N_19412,N_19208,N_19121);
xnor U19413 (N_19413,N_19024,N_19105);
or U19414 (N_19414,N_19236,N_19069);
nor U19415 (N_19415,N_19216,N_19136);
or U19416 (N_19416,N_19132,N_19178);
nand U19417 (N_19417,N_19012,N_19150);
nor U19418 (N_19418,N_19079,N_19088);
xor U19419 (N_19419,N_19185,N_19043);
nor U19420 (N_19420,N_19093,N_19000);
and U19421 (N_19421,N_19143,N_19197);
nor U19422 (N_19422,N_19094,N_19182);
nor U19423 (N_19423,N_19069,N_19114);
or U19424 (N_19424,N_19117,N_19031);
and U19425 (N_19425,N_19104,N_19066);
xor U19426 (N_19426,N_19230,N_19045);
or U19427 (N_19427,N_19224,N_19006);
and U19428 (N_19428,N_19108,N_19105);
and U19429 (N_19429,N_19118,N_19095);
or U19430 (N_19430,N_19224,N_19028);
and U19431 (N_19431,N_19208,N_19196);
xor U19432 (N_19432,N_19066,N_19037);
or U19433 (N_19433,N_19034,N_19071);
and U19434 (N_19434,N_19027,N_19020);
and U19435 (N_19435,N_19063,N_19199);
nor U19436 (N_19436,N_19139,N_19185);
and U19437 (N_19437,N_19132,N_19231);
nand U19438 (N_19438,N_19076,N_19144);
nor U19439 (N_19439,N_19162,N_19061);
nor U19440 (N_19440,N_19173,N_19157);
nand U19441 (N_19441,N_19215,N_19021);
nor U19442 (N_19442,N_19147,N_19098);
xnor U19443 (N_19443,N_19153,N_19173);
nand U19444 (N_19444,N_19244,N_19035);
nand U19445 (N_19445,N_19013,N_19192);
or U19446 (N_19446,N_19116,N_19050);
and U19447 (N_19447,N_19070,N_19042);
or U19448 (N_19448,N_19243,N_19099);
xnor U19449 (N_19449,N_19034,N_19087);
nor U19450 (N_19450,N_19239,N_19063);
or U19451 (N_19451,N_19013,N_19128);
or U19452 (N_19452,N_19041,N_19174);
nor U19453 (N_19453,N_19023,N_19199);
xnor U19454 (N_19454,N_19168,N_19042);
and U19455 (N_19455,N_19128,N_19156);
or U19456 (N_19456,N_19201,N_19036);
nor U19457 (N_19457,N_19126,N_19061);
nand U19458 (N_19458,N_19036,N_19011);
nor U19459 (N_19459,N_19211,N_19023);
nand U19460 (N_19460,N_19225,N_19069);
or U19461 (N_19461,N_19136,N_19070);
nand U19462 (N_19462,N_19099,N_19155);
nand U19463 (N_19463,N_19112,N_19168);
nand U19464 (N_19464,N_19130,N_19010);
and U19465 (N_19465,N_19092,N_19103);
nor U19466 (N_19466,N_19121,N_19079);
nor U19467 (N_19467,N_19133,N_19243);
or U19468 (N_19468,N_19144,N_19071);
nand U19469 (N_19469,N_19205,N_19074);
nor U19470 (N_19470,N_19221,N_19012);
or U19471 (N_19471,N_19212,N_19203);
and U19472 (N_19472,N_19230,N_19160);
xnor U19473 (N_19473,N_19020,N_19061);
and U19474 (N_19474,N_19210,N_19160);
or U19475 (N_19475,N_19192,N_19177);
nand U19476 (N_19476,N_19075,N_19137);
nor U19477 (N_19477,N_19124,N_19058);
nand U19478 (N_19478,N_19170,N_19108);
nor U19479 (N_19479,N_19060,N_19033);
or U19480 (N_19480,N_19128,N_19072);
nand U19481 (N_19481,N_19183,N_19019);
or U19482 (N_19482,N_19094,N_19240);
or U19483 (N_19483,N_19150,N_19077);
nand U19484 (N_19484,N_19125,N_19028);
and U19485 (N_19485,N_19031,N_19219);
and U19486 (N_19486,N_19017,N_19138);
and U19487 (N_19487,N_19014,N_19111);
nand U19488 (N_19488,N_19120,N_19042);
and U19489 (N_19489,N_19165,N_19216);
and U19490 (N_19490,N_19039,N_19022);
and U19491 (N_19491,N_19158,N_19085);
or U19492 (N_19492,N_19056,N_19213);
or U19493 (N_19493,N_19126,N_19190);
nand U19494 (N_19494,N_19194,N_19026);
or U19495 (N_19495,N_19085,N_19234);
xor U19496 (N_19496,N_19238,N_19034);
nor U19497 (N_19497,N_19057,N_19092);
nand U19498 (N_19498,N_19101,N_19069);
nand U19499 (N_19499,N_19017,N_19007);
or U19500 (N_19500,N_19474,N_19430);
nor U19501 (N_19501,N_19420,N_19482);
nor U19502 (N_19502,N_19453,N_19466);
nand U19503 (N_19503,N_19313,N_19419);
nand U19504 (N_19504,N_19257,N_19256);
and U19505 (N_19505,N_19417,N_19387);
or U19506 (N_19506,N_19471,N_19371);
nor U19507 (N_19507,N_19410,N_19350);
xnor U19508 (N_19508,N_19403,N_19270);
and U19509 (N_19509,N_19394,N_19438);
nand U19510 (N_19510,N_19253,N_19268);
nand U19511 (N_19511,N_19284,N_19349);
and U19512 (N_19512,N_19289,N_19365);
nand U19513 (N_19513,N_19393,N_19288);
nand U19514 (N_19514,N_19261,N_19279);
or U19515 (N_19515,N_19359,N_19331);
or U19516 (N_19516,N_19367,N_19377);
nand U19517 (N_19517,N_19290,N_19298);
nor U19518 (N_19518,N_19335,N_19328);
xor U19519 (N_19519,N_19469,N_19461);
nor U19520 (N_19520,N_19418,N_19498);
nand U19521 (N_19521,N_19300,N_19472);
or U19522 (N_19522,N_19323,N_19434);
nand U19523 (N_19523,N_19433,N_19250);
and U19524 (N_19524,N_19283,N_19446);
or U19525 (N_19525,N_19338,N_19368);
or U19526 (N_19526,N_19319,N_19330);
xnor U19527 (N_19527,N_19355,N_19413);
xnor U19528 (N_19528,N_19314,N_19342);
nor U19529 (N_19529,N_19439,N_19347);
nand U19530 (N_19530,N_19399,N_19346);
and U19531 (N_19531,N_19448,N_19302);
or U19532 (N_19532,N_19389,N_19460);
nand U19533 (N_19533,N_19405,N_19372);
xnor U19534 (N_19534,N_19479,N_19429);
nand U19535 (N_19535,N_19386,N_19409);
or U19536 (N_19536,N_19485,N_19275);
and U19537 (N_19537,N_19316,N_19476);
nor U19538 (N_19538,N_19340,N_19470);
or U19539 (N_19539,N_19269,N_19447);
nor U19540 (N_19540,N_19325,N_19293);
xnor U19541 (N_19541,N_19396,N_19424);
or U19542 (N_19542,N_19273,N_19352);
nand U19543 (N_19543,N_19265,N_19334);
nor U19544 (N_19544,N_19337,N_19499);
xnor U19545 (N_19545,N_19489,N_19307);
nor U19546 (N_19546,N_19304,N_19407);
nor U19547 (N_19547,N_19291,N_19363);
and U19548 (N_19548,N_19381,N_19455);
xnor U19549 (N_19549,N_19361,N_19408);
and U19550 (N_19550,N_19451,N_19495);
xnor U19551 (N_19551,N_19286,N_19422);
and U19552 (N_19552,N_19467,N_19327);
or U19553 (N_19553,N_19456,N_19440);
and U19554 (N_19554,N_19374,N_19481);
and U19555 (N_19555,N_19390,N_19322);
or U19556 (N_19556,N_19339,N_19445);
xor U19557 (N_19557,N_19303,N_19406);
and U19558 (N_19558,N_19262,N_19294);
nor U19559 (N_19559,N_19383,N_19404);
xnor U19560 (N_19560,N_19492,N_19296);
xor U19561 (N_19561,N_19473,N_19345);
nor U19562 (N_19562,N_19266,N_19358);
nor U19563 (N_19563,N_19332,N_19395);
or U19564 (N_19564,N_19251,N_19295);
and U19565 (N_19565,N_19311,N_19398);
xor U19566 (N_19566,N_19309,N_19380);
nand U19567 (N_19567,N_19397,N_19324);
nand U19568 (N_19568,N_19252,N_19486);
and U19569 (N_19569,N_19321,N_19475);
and U19570 (N_19570,N_19497,N_19435);
nor U19571 (N_19571,N_19391,N_19369);
nand U19572 (N_19572,N_19312,N_19348);
nand U19573 (N_19573,N_19452,N_19400);
nor U19574 (N_19574,N_19494,N_19378);
xnor U19575 (N_19575,N_19259,N_19427);
nand U19576 (N_19576,N_19281,N_19305);
nand U19577 (N_19577,N_19462,N_19276);
or U19578 (N_19578,N_19382,N_19306);
and U19579 (N_19579,N_19336,N_19326);
nand U19580 (N_19580,N_19333,N_19356);
nor U19581 (N_19581,N_19457,N_19272);
xnor U19582 (N_19582,N_19370,N_19432);
nor U19583 (N_19583,N_19488,N_19375);
nor U19584 (N_19584,N_19428,N_19384);
or U19585 (N_19585,N_19354,N_19360);
and U19586 (N_19586,N_19416,N_19301);
nor U19587 (N_19587,N_19425,N_19415);
xor U19588 (N_19588,N_19443,N_19357);
nor U19589 (N_19589,N_19411,N_19401);
and U19590 (N_19590,N_19423,N_19379);
nand U19591 (N_19591,N_19285,N_19491);
and U19592 (N_19592,N_19351,N_19441);
nand U19593 (N_19593,N_19280,N_19437);
and U19594 (N_19594,N_19282,N_19431);
nand U19595 (N_19595,N_19373,N_19264);
nand U19596 (N_19596,N_19483,N_19477);
and U19597 (N_19597,N_19315,N_19388);
xor U19598 (N_19598,N_19436,N_19278);
nor U19599 (N_19599,N_19478,N_19297);
or U19600 (N_19600,N_19287,N_19343);
nor U19601 (N_19601,N_19442,N_19366);
nand U19602 (N_19602,N_19414,N_19317);
and U19603 (N_19603,N_19362,N_19493);
nor U19604 (N_19604,N_19444,N_19459);
and U19605 (N_19605,N_19292,N_19484);
nand U19606 (N_19606,N_19412,N_19465);
or U19607 (N_19607,N_19310,N_19376);
or U19608 (N_19608,N_19490,N_19308);
nor U19609 (N_19609,N_19458,N_19385);
and U19610 (N_19610,N_19464,N_19450);
xor U19611 (N_19611,N_19480,N_19254);
or U19612 (N_19612,N_19463,N_19454);
nor U19613 (N_19613,N_19318,N_19402);
nor U19614 (N_19614,N_19341,N_19260);
and U19615 (N_19615,N_19274,N_19320);
nand U19616 (N_19616,N_19299,N_19258);
nor U19617 (N_19617,N_19267,N_19449);
and U19618 (N_19618,N_19344,N_19329);
nor U19619 (N_19619,N_19392,N_19468);
nand U19620 (N_19620,N_19487,N_19255);
nand U19621 (N_19621,N_19421,N_19364);
xor U19622 (N_19622,N_19426,N_19353);
nor U19623 (N_19623,N_19263,N_19277);
xnor U19624 (N_19624,N_19496,N_19271);
nand U19625 (N_19625,N_19271,N_19414);
and U19626 (N_19626,N_19373,N_19432);
nor U19627 (N_19627,N_19483,N_19365);
or U19628 (N_19628,N_19416,N_19430);
nor U19629 (N_19629,N_19459,N_19331);
nand U19630 (N_19630,N_19394,N_19377);
xnor U19631 (N_19631,N_19320,N_19305);
or U19632 (N_19632,N_19275,N_19419);
nand U19633 (N_19633,N_19431,N_19258);
nand U19634 (N_19634,N_19491,N_19479);
and U19635 (N_19635,N_19268,N_19277);
nor U19636 (N_19636,N_19486,N_19386);
nand U19637 (N_19637,N_19275,N_19386);
and U19638 (N_19638,N_19490,N_19466);
nor U19639 (N_19639,N_19445,N_19387);
and U19640 (N_19640,N_19380,N_19324);
xor U19641 (N_19641,N_19271,N_19476);
nand U19642 (N_19642,N_19478,N_19259);
or U19643 (N_19643,N_19449,N_19400);
or U19644 (N_19644,N_19452,N_19300);
nand U19645 (N_19645,N_19473,N_19361);
and U19646 (N_19646,N_19384,N_19300);
and U19647 (N_19647,N_19250,N_19493);
or U19648 (N_19648,N_19285,N_19348);
and U19649 (N_19649,N_19314,N_19370);
and U19650 (N_19650,N_19449,N_19293);
nand U19651 (N_19651,N_19420,N_19277);
nand U19652 (N_19652,N_19393,N_19451);
nand U19653 (N_19653,N_19391,N_19262);
and U19654 (N_19654,N_19256,N_19378);
nand U19655 (N_19655,N_19443,N_19288);
and U19656 (N_19656,N_19489,N_19435);
nor U19657 (N_19657,N_19412,N_19457);
nor U19658 (N_19658,N_19273,N_19317);
and U19659 (N_19659,N_19453,N_19298);
nor U19660 (N_19660,N_19287,N_19389);
xnor U19661 (N_19661,N_19349,N_19320);
or U19662 (N_19662,N_19317,N_19417);
and U19663 (N_19663,N_19496,N_19423);
or U19664 (N_19664,N_19292,N_19408);
nor U19665 (N_19665,N_19446,N_19459);
or U19666 (N_19666,N_19462,N_19343);
nor U19667 (N_19667,N_19370,N_19469);
or U19668 (N_19668,N_19412,N_19259);
and U19669 (N_19669,N_19261,N_19448);
or U19670 (N_19670,N_19339,N_19315);
and U19671 (N_19671,N_19296,N_19498);
xor U19672 (N_19672,N_19355,N_19332);
or U19673 (N_19673,N_19268,N_19474);
xor U19674 (N_19674,N_19320,N_19250);
and U19675 (N_19675,N_19271,N_19494);
nor U19676 (N_19676,N_19359,N_19493);
or U19677 (N_19677,N_19364,N_19383);
or U19678 (N_19678,N_19364,N_19264);
nor U19679 (N_19679,N_19357,N_19266);
nand U19680 (N_19680,N_19257,N_19315);
nand U19681 (N_19681,N_19376,N_19372);
and U19682 (N_19682,N_19277,N_19313);
and U19683 (N_19683,N_19297,N_19453);
and U19684 (N_19684,N_19460,N_19273);
nand U19685 (N_19685,N_19444,N_19436);
and U19686 (N_19686,N_19309,N_19265);
or U19687 (N_19687,N_19290,N_19453);
or U19688 (N_19688,N_19390,N_19280);
nor U19689 (N_19689,N_19415,N_19390);
or U19690 (N_19690,N_19485,N_19279);
nand U19691 (N_19691,N_19499,N_19470);
nor U19692 (N_19692,N_19418,N_19462);
nand U19693 (N_19693,N_19416,N_19482);
or U19694 (N_19694,N_19390,N_19417);
and U19695 (N_19695,N_19316,N_19264);
and U19696 (N_19696,N_19374,N_19397);
and U19697 (N_19697,N_19333,N_19428);
nor U19698 (N_19698,N_19333,N_19353);
nand U19699 (N_19699,N_19499,N_19422);
and U19700 (N_19700,N_19275,N_19468);
nand U19701 (N_19701,N_19326,N_19269);
nand U19702 (N_19702,N_19439,N_19360);
nand U19703 (N_19703,N_19449,N_19356);
nand U19704 (N_19704,N_19306,N_19362);
or U19705 (N_19705,N_19437,N_19390);
nor U19706 (N_19706,N_19483,N_19468);
xnor U19707 (N_19707,N_19410,N_19407);
or U19708 (N_19708,N_19481,N_19442);
nand U19709 (N_19709,N_19484,N_19333);
and U19710 (N_19710,N_19387,N_19418);
nor U19711 (N_19711,N_19259,N_19305);
nor U19712 (N_19712,N_19443,N_19302);
nor U19713 (N_19713,N_19375,N_19485);
nand U19714 (N_19714,N_19470,N_19440);
nor U19715 (N_19715,N_19492,N_19388);
and U19716 (N_19716,N_19439,N_19383);
and U19717 (N_19717,N_19423,N_19280);
and U19718 (N_19718,N_19397,N_19276);
and U19719 (N_19719,N_19473,N_19451);
and U19720 (N_19720,N_19250,N_19312);
and U19721 (N_19721,N_19273,N_19446);
nor U19722 (N_19722,N_19363,N_19482);
or U19723 (N_19723,N_19266,N_19254);
nor U19724 (N_19724,N_19373,N_19282);
nand U19725 (N_19725,N_19366,N_19341);
nand U19726 (N_19726,N_19429,N_19384);
nand U19727 (N_19727,N_19363,N_19465);
and U19728 (N_19728,N_19357,N_19265);
nor U19729 (N_19729,N_19383,N_19459);
xnor U19730 (N_19730,N_19377,N_19329);
and U19731 (N_19731,N_19375,N_19481);
nand U19732 (N_19732,N_19378,N_19364);
nand U19733 (N_19733,N_19450,N_19397);
and U19734 (N_19734,N_19343,N_19258);
and U19735 (N_19735,N_19381,N_19415);
nand U19736 (N_19736,N_19495,N_19412);
or U19737 (N_19737,N_19476,N_19403);
or U19738 (N_19738,N_19325,N_19364);
xor U19739 (N_19739,N_19464,N_19457);
xnor U19740 (N_19740,N_19426,N_19405);
nand U19741 (N_19741,N_19470,N_19497);
and U19742 (N_19742,N_19353,N_19373);
or U19743 (N_19743,N_19424,N_19356);
and U19744 (N_19744,N_19447,N_19436);
or U19745 (N_19745,N_19392,N_19328);
nand U19746 (N_19746,N_19295,N_19258);
or U19747 (N_19747,N_19324,N_19268);
nand U19748 (N_19748,N_19353,N_19330);
nor U19749 (N_19749,N_19388,N_19442);
or U19750 (N_19750,N_19689,N_19693);
nor U19751 (N_19751,N_19502,N_19621);
nor U19752 (N_19752,N_19730,N_19635);
or U19753 (N_19753,N_19717,N_19666);
nand U19754 (N_19754,N_19654,N_19676);
nand U19755 (N_19755,N_19560,N_19683);
nand U19756 (N_19756,N_19569,N_19627);
nand U19757 (N_19757,N_19741,N_19699);
and U19758 (N_19758,N_19700,N_19634);
nor U19759 (N_19759,N_19570,N_19610);
and U19760 (N_19760,N_19680,N_19644);
or U19761 (N_19761,N_19512,N_19547);
nand U19762 (N_19762,N_19546,N_19723);
or U19763 (N_19763,N_19539,N_19647);
nand U19764 (N_19764,N_19500,N_19590);
and U19765 (N_19765,N_19646,N_19556);
and U19766 (N_19766,N_19516,N_19582);
or U19767 (N_19767,N_19648,N_19624);
xor U19768 (N_19768,N_19507,N_19731);
xor U19769 (N_19769,N_19506,N_19612);
and U19770 (N_19770,N_19725,N_19508);
nor U19771 (N_19771,N_19585,N_19628);
or U19772 (N_19772,N_19598,N_19707);
or U19773 (N_19773,N_19688,N_19637);
and U19774 (N_19774,N_19573,N_19626);
and U19775 (N_19775,N_19538,N_19607);
and U19776 (N_19776,N_19535,N_19521);
nand U19777 (N_19777,N_19663,N_19727);
nand U19778 (N_19778,N_19713,N_19668);
or U19779 (N_19779,N_19739,N_19733);
and U19780 (N_19780,N_19669,N_19740);
nor U19781 (N_19781,N_19597,N_19691);
or U19782 (N_19782,N_19599,N_19682);
and U19783 (N_19783,N_19536,N_19613);
nor U19784 (N_19784,N_19686,N_19608);
and U19785 (N_19785,N_19653,N_19641);
and U19786 (N_19786,N_19665,N_19672);
and U19787 (N_19787,N_19574,N_19636);
nand U19788 (N_19788,N_19711,N_19735);
nand U19789 (N_19789,N_19588,N_19609);
nand U19790 (N_19790,N_19584,N_19677);
or U19791 (N_19791,N_19652,N_19620);
and U19792 (N_19792,N_19530,N_19600);
and U19793 (N_19793,N_19728,N_19593);
nor U19794 (N_19794,N_19695,N_19642);
and U19795 (N_19795,N_19643,N_19625);
and U19796 (N_19796,N_19747,N_19571);
nand U19797 (N_19797,N_19532,N_19640);
xnor U19798 (N_19798,N_19748,N_19659);
nand U19799 (N_19799,N_19687,N_19519);
nand U19800 (N_19800,N_19509,N_19743);
or U19801 (N_19801,N_19709,N_19722);
nand U19802 (N_19802,N_19716,N_19721);
nor U19803 (N_19803,N_19617,N_19726);
and U19804 (N_19804,N_19685,N_19745);
or U19805 (N_19805,N_19697,N_19522);
nand U19806 (N_19806,N_19596,N_19517);
and U19807 (N_19807,N_19515,N_19719);
nor U19808 (N_19808,N_19629,N_19632);
and U19809 (N_19809,N_19631,N_19592);
xnor U19810 (N_19810,N_19575,N_19664);
nor U19811 (N_19811,N_19523,N_19501);
xor U19812 (N_19812,N_19715,N_19553);
and U19813 (N_19813,N_19537,N_19557);
nand U19814 (N_19814,N_19558,N_19542);
or U19815 (N_19815,N_19618,N_19619);
nand U19816 (N_19816,N_19576,N_19744);
or U19817 (N_19817,N_19615,N_19681);
or U19818 (N_19818,N_19565,N_19630);
nor U19819 (N_19819,N_19503,N_19587);
nor U19820 (N_19820,N_19742,N_19572);
nor U19821 (N_19821,N_19712,N_19550);
nand U19822 (N_19822,N_19579,N_19692);
or U19823 (N_19823,N_19533,N_19678);
or U19824 (N_19824,N_19749,N_19606);
nor U19825 (N_19825,N_19710,N_19520);
nor U19826 (N_19826,N_19734,N_19605);
nor U19827 (N_19827,N_19566,N_19594);
and U19828 (N_19828,N_19564,N_19737);
nor U19829 (N_19829,N_19718,N_19581);
and U19830 (N_19830,N_19651,N_19667);
nor U19831 (N_19831,N_19578,N_19544);
xnor U19832 (N_19832,N_19633,N_19614);
and U19833 (N_19833,N_19561,N_19701);
nand U19834 (N_19834,N_19541,N_19696);
nor U19835 (N_19835,N_19673,N_19703);
and U19836 (N_19836,N_19562,N_19555);
xnor U19837 (N_19837,N_19510,N_19661);
nand U19838 (N_19838,N_19655,N_19704);
nor U19839 (N_19839,N_19513,N_19702);
nand U19840 (N_19840,N_19505,N_19720);
nand U19841 (N_19841,N_19738,N_19559);
xnor U19842 (N_19842,N_19658,N_19529);
and U19843 (N_19843,N_19623,N_19604);
or U19844 (N_19844,N_19545,N_19679);
nand U19845 (N_19845,N_19675,N_19694);
and U19846 (N_19846,N_19563,N_19638);
nor U19847 (N_19847,N_19543,N_19583);
and U19848 (N_19848,N_19586,N_19526);
xor U19849 (N_19849,N_19534,N_19746);
nor U19850 (N_19850,N_19705,N_19657);
nand U19851 (N_19851,N_19603,N_19577);
nand U19852 (N_19852,N_19662,N_19548);
nor U19853 (N_19853,N_19554,N_19660);
and U19854 (N_19854,N_19708,N_19567);
nor U19855 (N_19855,N_19616,N_19698);
nand U19856 (N_19856,N_19650,N_19595);
and U19857 (N_19857,N_19580,N_19706);
nand U19858 (N_19858,N_19591,N_19525);
nor U19859 (N_19859,N_19551,N_19674);
nor U19860 (N_19860,N_19602,N_19514);
nand U19861 (N_19861,N_19622,N_19656);
nand U19862 (N_19862,N_19504,N_19732);
nor U19863 (N_19863,N_19528,N_19527);
or U19864 (N_19864,N_19524,N_19645);
or U19865 (N_19865,N_19611,N_19714);
nor U19866 (N_19866,N_19540,N_19736);
nand U19867 (N_19867,N_19568,N_19511);
or U19868 (N_19868,N_19724,N_19601);
nand U19869 (N_19869,N_19552,N_19671);
and U19870 (N_19870,N_19639,N_19684);
or U19871 (N_19871,N_19729,N_19531);
and U19872 (N_19872,N_19690,N_19549);
or U19873 (N_19873,N_19518,N_19649);
or U19874 (N_19874,N_19670,N_19589);
nor U19875 (N_19875,N_19746,N_19543);
nand U19876 (N_19876,N_19507,N_19682);
or U19877 (N_19877,N_19696,N_19617);
nor U19878 (N_19878,N_19739,N_19555);
nand U19879 (N_19879,N_19621,N_19666);
and U19880 (N_19880,N_19707,N_19721);
and U19881 (N_19881,N_19664,N_19704);
nor U19882 (N_19882,N_19635,N_19520);
nor U19883 (N_19883,N_19575,N_19581);
nand U19884 (N_19884,N_19592,N_19709);
nor U19885 (N_19885,N_19519,N_19691);
and U19886 (N_19886,N_19644,N_19568);
or U19887 (N_19887,N_19531,N_19630);
nand U19888 (N_19888,N_19644,N_19668);
nand U19889 (N_19889,N_19620,N_19687);
xnor U19890 (N_19890,N_19693,N_19739);
nand U19891 (N_19891,N_19635,N_19587);
or U19892 (N_19892,N_19602,N_19674);
nor U19893 (N_19893,N_19567,N_19516);
and U19894 (N_19894,N_19702,N_19747);
xor U19895 (N_19895,N_19732,N_19539);
nor U19896 (N_19896,N_19726,N_19618);
and U19897 (N_19897,N_19571,N_19643);
nand U19898 (N_19898,N_19514,N_19576);
nand U19899 (N_19899,N_19747,N_19537);
xor U19900 (N_19900,N_19737,N_19648);
and U19901 (N_19901,N_19706,N_19583);
xnor U19902 (N_19902,N_19505,N_19537);
or U19903 (N_19903,N_19529,N_19669);
nor U19904 (N_19904,N_19692,N_19601);
and U19905 (N_19905,N_19527,N_19731);
or U19906 (N_19906,N_19593,N_19664);
and U19907 (N_19907,N_19634,N_19683);
xor U19908 (N_19908,N_19740,N_19667);
xor U19909 (N_19909,N_19692,N_19539);
nor U19910 (N_19910,N_19728,N_19622);
or U19911 (N_19911,N_19567,N_19715);
or U19912 (N_19912,N_19646,N_19598);
nor U19913 (N_19913,N_19522,N_19704);
or U19914 (N_19914,N_19695,N_19690);
and U19915 (N_19915,N_19605,N_19599);
and U19916 (N_19916,N_19559,N_19581);
or U19917 (N_19917,N_19732,N_19736);
nor U19918 (N_19918,N_19709,N_19683);
nand U19919 (N_19919,N_19704,N_19744);
and U19920 (N_19920,N_19518,N_19745);
nand U19921 (N_19921,N_19691,N_19682);
nor U19922 (N_19922,N_19663,N_19692);
nor U19923 (N_19923,N_19696,N_19592);
xor U19924 (N_19924,N_19632,N_19614);
nand U19925 (N_19925,N_19690,N_19729);
or U19926 (N_19926,N_19553,N_19731);
and U19927 (N_19927,N_19678,N_19727);
and U19928 (N_19928,N_19547,N_19515);
nand U19929 (N_19929,N_19704,N_19585);
or U19930 (N_19930,N_19643,N_19640);
xnor U19931 (N_19931,N_19549,N_19719);
nand U19932 (N_19932,N_19695,N_19613);
and U19933 (N_19933,N_19579,N_19626);
and U19934 (N_19934,N_19611,N_19659);
nand U19935 (N_19935,N_19674,N_19665);
nor U19936 (N_19936,N_19553,N_19706);
or U19937 (N_19937,N_19749,N_19649);
and U19938 (N_19938,N_19510,N_19748);
nor U19939 (N_19939,N_19689,N_19511);
and U19940 (N_19940,N_19670,N_19706);
and U19941 (N_19941,N_19552,N_19731);
nor U19942 (N_19942,N_19604,N_19746);
and U19943 (N_19943,N_19530,N_19646);
or U19944 (N_19944,N_19710,N_19559);
and U19945 (N_19945,N_19535,N_19545);
and U19946 (N_19946,N_19656,N_19731);
and U19947 (N_19947,N_19695,N_19547);
and U19948 (N_19948,N_19637,N_19548);
or U19949 (N_19949,N_19544,N_19678);
or U19950 (N_19950,N_19557,N_19548);
nand U19951 (N_19951,N_19561,N_19557);
or U19952 (N_19952,N_19524,N_19546);
nor U19953 (N_19953,N_19626,N_19593);
nand U19954 (N_19954,N_19598,N_19520);
nand U19955 (N_19955,N_19690,N_19641);
nand U19956 (N_19956,N_19516,N_19630);
and U19957 (N_19957,N_19628,N_19538);
and U19958 (N_19958,N_19647,N_19669);
or U19959 (N_19959,N_19653,N_19520);
nand U19960 (N_19960,N_19668,N_19553);
and U19961 (N_19961,N_19694,N_19656);
xor U19962 (N_19962,N_19578,N_19653);
nand U19963 (N_19963,N_19622,N_19574);
nand U19964 (N_19964,N_19693,N_19681);
nand U19965 (N_19965,N_19619,N_19657);
or U19966 (N_19966,N_19567,N_19500);
nor U19967 (N_19967,N_19735,N_19722);
or U19968 (N_19968,N_19549,N_19568);
nor U19969 (N_19969,N_19744,N_19573);
nand U19970 (N_19970,N_19616,N_19590);
and U19971 (N_19971,N_19618,N_19675);
nand U19972 (N_19972,N_19697,N_19726);
and U19973 (N_19973,N_19730,N_19663);
or U19974 (N_19974,N_19615,N_19662);
nand U19975 (N_19975,N_19602,N_19595);
nand U19976 (N_19976,N_19704,N_19666);
nand U19977 (N_19977,N_19711,N_19659);
and U19978 (N_19978,N_19628,N_19645);
nand U19979 (N_19979,N_19697,N_19685);
or U19980 (N_19980,N_19720,N_19748);
nor U19981 (N_19981,N_19621,N_19699);
and U19982 (N_19982,N_19662,N_19730);
and U19983 (N_19983,N_19581,N_19744);
xor U19984 (N_19984,N_19664,N_19527);
nand U19985 (N_19985,N_19518,N_19719);
xor U19986 (N_19986,N_19665,N_19577);
xnor U19987 (N_19987,N_19643,N_19711);
and U19988 (N_19988,N_19729,N_19508);
nand U19989 (N_19989,N_19684,N_19712);
and U19990 (N_19990,N_19546,N_19517);
nor U19991 (N_19991,N_19504,N_19720);
and U19992 (N_19992,N_19702,N_19698);
nor U19993 (N_19993,N_19723,N_19733);
nand U19994 (N_19994,N_19731,N_19525);
nor U19995 (N_19995,N_19739,N_19543);
nand U19996 (N_19996,N_19525,N_19697);
or U19997 (N_19997,N_19714,N_19712);
or U19998 (N_19998,N_19694,N_19513);
and U19999 (N_19999,N_19703,N_19603);
or UO_0 (O_0,N_19769,N_19874);
xor UO_1 (O_1,N_19973,N_19960);
nor UO_2 (O_2,N_19901,N_19869);
or UO_3 (O_3,N_19799,N_19822);
or UO_4 (O_4,N_19850,N_19770);
or UO_5 (O_5,N_19995,N_19956);
and UO_6 (O_6,N_19875,N_19857);
or UO_7 (O_7,N_19759,N_19972);
nand UO_8 (O_8,N_19929,N_19924);
or UO_9 (O_9,N_19826,N_19785);
nor UO_10 (O_10,N_19800,N_19763);
or UO_11 (O_11,N_19774,N_19779);
xor UO_12 (O_12,N_19928,N_19893);
nand UO_13 (O_13,N_19903,N_19767);
xnor UO_14 (O_14,N_19915,N_19978);
nor UO_15 (O_15,N_19834,N_19912);
nor UO_16 (O_16,N_19852,N_19982);
or UO_17 (O_17,N_19992,N_19753);
or UO_18 (O_18,N_19780,N_19938);
or UO_19 (O_19,N_19983,N_19756);
nor UO_20 (O_20,N_19803,N_19896);
and UO_21 (O_21,N_19889,N_19867);
and UO_22 (O_22,N_19911,N_19768);
nor UO_23 (O_23,N_19825,N_19784);
and UO_24 (O_24,N_19847,N_19815);
or UO_25 (O_25,N_19891,N_19844);
nand UO_26 (O_26,N_19892,N_19921);
nand UO_27 (O_27,N_19955,N_19760);
nand UO_28 (O_28,N_19809,N_19835);
nor UO_29 (O_29,N_19843,N_19794);
nor UO_30 (O_30,N_19860,N_19861);
nor UO_31 (O_31,N_19888,N_19933);
nor UO_32 (O_32,N_19854,N_19899);
and UO_33 (O_33,N_19919,N_19975);
and UO_34 (O_34,N_19864,N_19971);
nor UO_35 (O_35,N_19751,N_19908);
nor UO_36 (O_36,N_19851,N_19841);
nand UO_37 (O_37,N_19793,N_19996);
nor UO_38 (O_38,N_19820,N_19991);
nor UO_39 (O_39,N_19942,N_19909);
nor UO_40 (O_40,N_19918,N_19957);
nand UO_41 (O_41,N_19946,N_19798);
nor UO_42 (O_42,N_19750,N_19900);
xor UO_43 (O_43,N_19872,N_19807);
nand UO_44 (O_44,N_19894,N_19881);
nand UO_45 (O_45,N_19859,N_19849);
or UO_46 (O_46,N_19974,N_19837);
nor UO_47 (O_47,N_19987,N_19878);
and UO_48 (O_48,N_19865,N_19949);
and UO_49 (O_49,N_19808,N_19817);
or UO_50 (O_50,N_19999,N_19968);
and UO_51 (O_51,N_19887,N_19805);
nor UO_52 (O_52,N_19787,N_19922);
and UO_53 (O_53,N_19790,N_19836);
or UO_54 (O_54,N_19950,N_19776);
xnor UO_55 (O_55,N_19804,N_19965);
nor UO_56 (O_56,N_19883,N_19797);
nand UO_57 (O_57,N_19816,N_19970);
and UO_58 (O_58,N_19876,N_19752);
xor UO_59 (O_59,N_19917,N_19882);
nor UO_60 (O_60,N_19827,N_19765);
xnor UO_61 (O_61,N_19904,N_19947);
xor UO_62 (O_62,N_19961,N_19819);
nor UO_63 (O_63,N_19945,N_19940);
nand UO_64 (O_64,N_19831,N_19858);
and UO_65 (O_65,N_19846,N_19979);
nand UO_66 (O_66,N_19840,N_19762);
and UO_67 (O_67,N_19905,N_19885);
or UO_68 (O_68,N_19890,N_19862);
nand UO_69 (O_69,N_19783,N_19997);
or UO_70 (O_70,N_19833,N_19796);
nand UO_71 (O_71,N_19856,N_19907);
or UO_72 (O_72,N_19761,N_19788);
or UO_73 (O_73,N_19944,N_19966);
or UO_74 (O_74,N_19939,N_19772);
nand UO_75 (O_75,N_19895,N_19778);
and UO_76 (O_76,N_19832,N_19792);
nand UO_77 (O_77,N_19980,N_19935);
nand UO_78 (O_78,N_19998,N_19814);
and UO_79 (O_79,N_19927,N_19879);
or UO_80 (O_80,N_19910,N_19838);
or UO_81 (O_81,N_19936,N_19986);
or UO_82 (O_82,N_19818,N_19994);
xnor UO_83 (O_83,N_19871,N_19842);
nor UO_84 (O_84,N_19959,N_19926);
xnor UO_85 (O_85,N_19934,N_19773);
and UO_86 (O_86,N_19810,N_19951);
and UO_87 (O_87,N_19870,N_19764);
nand UO_88 (O_88,N_19988,N_19898);
nor UO_89 (O_89,N_19902,N_19990);
and UO_90 (O_90,N_19954,N_19916);
nor UO_91 (O_91,N_19771,N_19828);
nor UO_92 (O_92,N_19863,N_19967);
nor UO_93 (O_93,N_19877,N_19873);
and UO_94 (O_94,N_19806,N_19932);
nor UO_95 (O_95,N_19839,N_19853);
and UO_96 (O_96,N_19984,N_19913);
nor UO_97 (O_97,N_19845,N_19964);
nor UO_98 (O_98,N_19766,N_19930);
nor UO_99 (O_99,N_19830,N_19981);
and UO_100 (O_100,N_19897,N_19777);
nor UO_101 (O_101,N_19813,N_19989);
or UO_102 (O_102,N_19914,N_19884);
nor UO_103 (O_103,N_19824,N_19985);
and UO_104 (O_104,N_19923,N_19920);
nor UO_105 (O_105,N_19958,N_19906);
nand UO_106 (O_106,N_19812,N_19931);
nand UO_107 (O_107,N_19758,N_19755);
nor UO_108 (O_108,N_19811,N_19782);
nand UO_109 (O_109,N_19855,N_19937);
xnor UO_110 (O_110,N_19848,N_19791);
or UO_111 (O_111,N_19821,N_19823);
nand UO_112 (O_112,N_19943,N_19801);
or UO_113 (O_113,N_19795,N_19953);
nand UO_114 (O_114,N_19829,N_19802);
nor UO_115 (O_115,N_19948,N_19880);
and UO_116 (O_116,N_19886,N_19789);
or UO_117 (O_117,N_19868,N_19866);
nor UO_118 (O_118,N_19977,N_19962);
nand UO_119 (O_119,N_19941,N_19775);
nor UO_120 (O_120,N_19754,N_19952);
and UO_121 (O_121,N_19993,N_19757);
nor UO_122 (O_122,N_19969,N_19963);
nor UO_123 (O_123,N_19781,N_19925);
nor UO_124 (O_124,N_19786,N_19976);
and UO_125 (O_125,N_19767,N_19761);
xnor UO_126 (O_126,N_19960,N_19768);
nand UO_127 (O_127,N_19983,N_19833);
nor UO_128 (O_128,N_19937,N_19818);
nor UO_129 (O_129,N_19933,N_19845);
xor UO_130 (O_130,N_19814,N_19911);
nand UO_131 (O_131,N_19990,N_19837);
nor UO_132 (O_132,N_19964,N_19927);
nor UO_133 (O_133,N_19803,N_19763);
or UO_134 (O_134,N_19801,N_19824);
or UO_135 (O_135,N_19895,N_19795);
or UO_136 (O_136,N_19807,N_19906);
nand UO_137 (O_137,N_19777,N_19846);
or UO_138 (O_138,N_19833,N_19880);
or UO_139 (O_139,N_19793,N_19962);
and UO_140 (O_140,N_19811,N_19927);
nor UO_141 (O_141,N_19946,N_19979);
and UO_142 (O_142,N_19780,N_19913);
nor UO_143 (O_143,N_19833,N_19774);
nand UO_144 (O_144,N_19837,N_19802);
nand UO_145 (O_145,N_19820,N_19892);
and UO_146 (O_146,N_19935,N_19865);
or UO_147 (O_147,N_19923,N_19876);
nor UO_148 (O_148,N_19767,N_19754);
nor UO_149 (O_149,N_19888,N_19974);
nor UO_150 (O_150,N_19804,N_19833);
nor UO_151 (O_151,N_19927,N_19995);
nor UO_152 (O_152,N_19919,N_19777);
or UO_153 (O_153,N_19886,N_19897);
nand UO_154 (O_154,N_19991,N_19842);
nor UO_155 (O_155,N_19874,N_19878);
xor UO_156 (O_156,N_19855,N_19949);
and UO_157 (O_157,N_19871,N_19912);
nor UO_158 (O_158,N_19892,N_19962);
nand UO_159 (O_159,N_19753,N_19879);
and UO_160 (O_160,N_19969,N_19822);
nor UO_161 (O_161,N_19810,N_19845);
nand UO_162 (O_162,N_19817,N_19864);
nor UO_163 (O_163,N_19807,N_19892);
xnor UO_164 (O_164,N_19809,N_19801);
and UO_165 (O_165,N_19881,N_19895);
and UO_166 (O_166,N_19890,N_19891);
and UO_167 (O_167,N_19877,N_19862);
and UO_168 (O_168,N_19978,N_19808);
nor UO_169 (O_169,N_19950,N_19765);
or UO_170 (O_170,N_19864,N_19795);
or UO_171 (O_171,N_19983,N_19755);
xor UO_172 (O_172,N_19751,N_19755);
or UO_173 (O_173,N_19870,N_19946);
or UO_174 (O_174,N_19796,N_19819);
nor UO_175 (O_175,N_19785,N_19860);
nor UO_176 (O_176,N_19791,N_19855);
nand UO_177 (O_177,N_19999,N_19771);
nand UO_178 (O_178,N_19768,N_19886);
and UO_179 (O_179,N_19864,N_19787);
nand UO_180 (O_180,N_19945,N_19853);
or UO_181 (O_181,N_19760,N_19818);
nor UO_182 (O_182,N_19909,N_19844);
or UO_183 (O_183,N_19789,N_19929);
or UO_184 (O_184,N_19840,N_19915);
or UO_185 (O_185,N_19835,N_19932);
nand UO_186 (O_186,N_19807,N_19948);
xnor UO_187 (O_187,N_19943,N_19830);
and UO_188 (O_188,N_19981,N_19937);
nand UO_189 (O_189,N_19930,N_19985);
xnor UO_190 (O_190,N_19837,N_19790);
nor UO_191 (O_191,N_19829,N_19786);
nand UO_192 (O_192,N_19992,N_19799);
nor UO_193 (O_193,N_19840,N_19960);
and UO_194 (O_194,N_19880,N_19797);
xor UO_195 (O_195,N_19811,N_19840);
and UO_196 (O_196,N_19807,N_19805);
and UO_197 (O_197,N_19999,N_19874);
and UO_198 (O_198,N_19903,N_19935);
xnor UO_199 (O_199,N_19892,N_19758);
or UO_200 (O_200,N_19820,N_19778);
and UO_201 (O_201,N_19798,N_19819);
or UO_202 (O_202,N_19753,N_19819);
xnor UO_203 (O_203,N_19848,N_19945);
and UO_204 (O_204,N_19751,N_19964);
or UO_205 (O_205,N_19994,N_19972);
nor UO_206 (O_206,N_19790,N_19877);
or UO_207 (O_207,N_19898,N_19978);
nand UO_208 (O_208,N_19836,N_19969);
or UO_209 (O_209,N_19789,N_19760);
and UO_210 (O_210,N_19779,N_19999);
nor UO_211 (O_211,N_19984,N_19905);
or UO_212 (O_212,N_19875,N_19929);
nor UO_213 (O_213,N_19990,N_19918);
nor UO_214 (O_214,N_19753,N_19871);
nor UO_215 (O_215,N_19759,N_19836);
and UO_216 (O_216,N_19850,N_19840);
or UO_217 (O_217,N_19880,N_19937);
nor UO_218 (O_218,N_19953,N_19870);
nor UO_219 (O_219,N_19864,N_19885);
or UO_220 (O_220,N_19860,N_19938);
xor UO_221 (O_221,N_19939,N_19920);
or UO_222 (O_222,N_19897,N_19856);
and UO_223 (O_223,N_19920,N_19965);
or UO_224 (O_224,N_19983,N_19822);
nand UO_225 (O_225,N_19762,N_19938);
nand UO_226 (O_226,N_19883,N_19785);
nor UO_227 (O_227,N_19901,N_19753);
nand UO_228 (O_228,N_19973,N_19767);
or UO_229 (O_229,N_19975,N_19867);
nand UO_230 (O_230,N_19810,N_19909);
nand UO_231 (O_231,N_19875,N_19802);
nand UO_232 (O_232,N_19767,N_19783);
or UO_233 (O_233,N_19861,N_19952);
and UO_234 (O_234,N_19835,N_19832);
or UO_235 (O_235,N_19981,N_19846);
and UO_236 (O_236,N_19865,N_19802);
nor UO_237 (O_237,N_19957,N_19870);
nand UO_238 (O_238,N_19989,N_19854);
or UO_239 (O_239,N_19935,N_19895);
or UO_240 (O_240,N_19879,N_19790);
xnor UO_241 (O_241,N_19973,N_19999);
and UO_242 (O_242,N_19857,N_19903);
and UO_243 (O_243,N_19930,N_19886);
or UO_244 (O_244,N_19909,N_19895);
nor UO_245 (O_245,N_19821,N_19873);
xnor UO_246 (O_246,N_19922,N_19910);
nand UO_247 (O_247,N_19893,N_19765);
nor UO_248 (O_248,N_19899,N_19793);
xnor UO_249 (O_249,N_19799,N_19872);
or UO_250 (O_250,N_19814,N_19908);
nor UO_251 (O_251,N_19923,N_19973);
and UO_252 (O_252,N_19771,N_19817);
and UO_253 (O_253,N_19825,N_19828);
or UO_254 (O_254,N_19896,N_19906);
nand UO_255 (O_255,N_19750,N_19867);
and UO_256 (O_256,N_19868,N_19826);
nand UO_257 (O_257,N_19875,N_19934);
nand UO_258 (O_258,N_19928,N_19830);
and UO_259 (O_259,N_19867,N_19767);
or UO_260 (O_260,N_19932,N_19779);
nand UO_261 (O_261,N_19918,N_19751);
or UO_262 (O_262,N_19824,N_19898);
nor UO_263 (O_263,N_19974,N_19943);
nand UO_264 (O_264,N_19967,N_19941);
or UO_265 (O_265,N_19852,N_19938);
and UO_266 (O_266,N_19861,N_19934);
nor UO_267 (O_267,N_19837,N_19854);
nand UO_268 (O_268,N_19935,N_19951);
and UO_269 (O_269,N_19874,N_19945);
and UO_270 (O_270,N_19768,N_19983);
nor UO_271 (O_271,N_19803,N_19880);
and UO_272 (O_272,N_19772,N_19881);
nand UO_273 (O_273,N_19771,N_19847);
or UO_274 (O_274,N_19942,N_19952);
nand UO_275 (O_275,N_19902,N_19820);
nand UO_276 (O_276,N_19996,N_19965);
nand UO_277 (O_277,N_19805,N_19992);
or UO_278 (O_278,N_19892,N_19946);
nor UO_279 (O_279,N_19964,N_19941);
or UO_280 (O_280,N_19971,N_19855);
nand UO_281 (O_281,N_19910,N_19980);
and UO_282 (O_282,N_19872,N_19991);
xor UO_283 (O_283,N_19859,N_19836);
and UO_284 (O_284,N_19779,N_19895);
nand UO_285 (O_285,N_19798,N_19862);
nand UO_286 (O_286,N_19759,N_19976);
xnor UO_287 (O_287,N_19839,N_19973);
nor UO_288 (O_288,N_19753,N_19840);
xnor UO_289 (O_289,N_19813,N_19819);
and UO_290 (O_290,N_19852,N_19817);
nand UO_291 (O_291,N_19982,N_19851);
or UO_292 (O_292,N_19921,N_19985);
and UO_293 (O_293,N_19948,N_19793);
or UO_294 (O_294,N_19840,N_19761);
nor UO_295 (O_295,N_19828,N_19754);
and UO_296 (O_296,N_19936,N_19800);
nor UO_297 (O_297,N_19826,N_19977);
and UO_298 (O_298,N_19951,N_19931);
and UO_299 (O_299,N_19772,N_19801);
and UO_300 (O_300,N_19898,N_19765);
xnor UO_301 (O_301,N_19955,N_19954);
and UO_302 (O_302,N_19877,N_19913);
nand UO_303 (O_303,N_19956,N_19952);
or UO_304 (O_304,N_19942,N_19856);
and UO_305 (O_305,N_19819,N_19762);
nor UO_306 (O_306,N_19906,N_19921);
or UO_307 (O_307,N_19911,N_19777);
nand UO_308 (O_308,N_19943,N_19938);
xnor UO_309 (O_309,N_19989,N_19821);
xor UO_310 (O_310,N_19876,N_19773);
nand UO_311 (O_311,N_19871,N_19763);
nor UO_312 (O_312,N_19944,N_19911);
nand UO_313 (O_313,N_19992,N_19796);
nor UO_314 (O_314,N_19862,N_19951);
nor UO_315 (O_315,N_19787,N_19939);
nor UO_316 (O_316,N_19815,N_19995);
xor UO_317 (O_317,N_19883,N_19770);
or UO_318 (O_318,N_19847,N_19793);
xor UO_319 (O_319,N_19919,N_19897);
xor UO_320 (O_320,N_19776,N_19932);
nor UO_321 (O_321,N_19752,N_19842);
nor UO_322 (O_322,N_19989,N_19764);
and UO_323 (O_323,N_19861,N_19852);
nor UO_324 (O_324,N_19752,N_19921);
and UO_325 (O_325,N_19854,N_19931);
or UO_326 (O_326,N_19949,N_19861);
or UO_327 (O_327,N_19915,N_19998);
xor UO_328 (O_328,N_19890,N_19878);
and UO_329 (O_329,N_19853,N_19892);
nand UO_330 (O_330,N_19773,N_19925);
nand UO_331 (O_331,N_19992,N_19984);
or UO_332 (O_332,N_19906,N_19780);
nand UO_333 (O_333,N_19934,N_19818);
nor UO_334 (O_334,N_19990,N_19921);
nor UO_335 (O_335,N_19947,N_19800);
nand UO_336 (O_336,N_19757,N_19901);
nand UO_337 (O_337,N_19880,N_19958);
or UO_338 (O_338,N_19944,N_19887);
and UO_339 (O_339,N_19753,N_19891);
nor UO_340 (O_340,N_19962,N_19939);
and UO_341 (O_341,N_19801,N_19915);
and UO_342 (O_342,N_19776,N_19935);
nand UO_343 (O_343,N_19975,N_19930);
nor UO_344 (O_344,N_19753,N_19866);
and UO_345 (O_345,N_19779,N_19832);
or UO_346 (O_346,N_19901,N_19925);
nand UO_347 (O_347,N_19853,N_19847);
xnor UO_348 (O_348,N_19946,N_19938);
nand UO_349 (O_349,N_19980,N_19832);
nor UO_350 (O_350,N_19936,N_19978);
nor UO_351 (O_351,N_19833,N_19893);
or UO_352 (O_352,N_19991,N_19886);
nand UO_353 (O_353,N_19822,N_19875);
and UO_354 (O_354,N_19956,N_19850);
nand UO_355 (O_355,N_19891,N_19947);
or UO_356 (O_356,N_19925,N_19972);
nand UO_357 (O_357,N_19952,N_19971);
nand UO_358 (O_358,N_19862,N_19815);
and UO_359 (O_359,N_19985,N_19883);
or UO_360 (O_360,N_19968,N_19820);
and UO_361 (O_361,N_19950,N_19918);
or UO_362 (O_362,N_19995,N_19953);
nand UO_363 (O_363,N_19776,N_19910);
nand UO_364 (O_364,N_19959,N_19859);
nor UO_365 (O_365,N_19830,N_19805);
and UO_366 (O_366,N_19799,N_19894);
or UO_367 (O_367,N_19955,N_19776);
or UO_368 (O_368,N_19910,N_19981);
and UO_369 (O_369,N_19753,N_19847);
nand UO_370 (O_370,N_19870,N_19829);
nor UO_371 (O_371,N_19965,N_19993);
nand UO_372 (O_372,N_19997,N_19876);
nand UO_373 (O_373,N_19777,N_19977);
or UO_374 (O_374,N_19821,N_19960);
and UO_375 (O_375,N_19755,N_19994);
nand UO_376 (O_376,N_19796,N_19761);
nor UO_377 (O_377,N_19805,N_19838);
nor UO_378 (O_378,N_19917,N_19953);
and UO_379 (O_379,N_19787,N_19869);
nand UO_380 (O_380,N_19879,N_19758);
nor UO_381 (O_381,N_19946,N_19929);
nand UO_382 (O_382,N_19900,N_19783);
nor UO_383 (O_383,N_19840,N_19869);
and UO_384 (O_384,N_19790,N_19849);
and UO_385 (O_385,N_19894,N_19928);
and UO_386 (O_386,N_19753,N_19993);
or UO_387 (O_387,N_19885,N_19751);
or UO_388 (O_388,N_19887,N_19987);
or UO_389 (O_389,N_19800,N_19814);
and UO_390 (O_390,N_19890,N_19888);
nor UO_391 (O_391,N_19992,N_19770);
xnor UO_392 (O_392,N_19828,N_19795);
nand UO_393 (O_393,N_19757,N_19979);
nor UO_394 (O_394,N_19875,N_19821);
nand UO_395 (O_395,N_19850,N_19937);
nor UO_396 (O_396,N_19839,N_19831);
nand UO_397 (O_397,N_19941,N_19853);
nor UO_398 (O_398,N_19778,N_19758);
or UO_399 (O_399,N_19858,N_19792);
nor UO_400 (O_400,N_19897,N_19825);
nand UO_401 (O_401,N_19851,N_19800);
nand UO_402 (O_402,N_19880,N_19938);
nand UO_403 (O_403,N_19889,N_19901);
nand UO_404 (O_404,N_19897,N_19761);
or UO_405 (O_405,N_19804,N_19966);
nor UO_406 (O_406,N_19859,N_19819);
nand UO_407 (O_407,N_19938,N_19974);
nand UO_408 (O_408,N_19964,N_19846);
and UO_409 (O_409,N_19886,N_19862);
and UO_410 (O_410,N_19993,N_19808);
nor UO_411 (O_411,N_19926,N_19961);
xnor UO_412 (O_412,N_19778,N_19850);
nor UO_413 (O_413,N_19994,N_19815);
or UO_414 (O_414,N_19780,N_19994);
nand UO_415 (O_415,N_19772,N_19973);
xnor UO_416 (O_416,N_19877,N_19881);
or UO_417 (O_417,N_19981,N_19953);
or UO_418 (O_418,N_19780,N_19779);
or UO_419 (O_419,N_19998,N_19826);
xnor UO_420 (O_420,N_19994,N_19914);
and UO_421 (O_421,N_19937,N_19760);
or UO_422 (O_422,N_19903,N_19750);
nand UO_423 (O_423,N_19969,N_19881);
and UO_424 (O_424,N_19991,N_19752);
nand UO_425 (O_425,N_19856,N_19973);
and UO_426 (O_426,N_19883,N_19853);
and UO_427 (O_427,N_19943,N_19783);
nor UO_428 (O_428,N_19878,N_19955);
and UO_429 (O_429,N_19862,N_19795);
or UO_430 (O_430,N_19788,N_19885);
nand UO_431 (O_431,N_19851,N_19965);
nand UO_432 (O_432,N_19881,N_19839);
and UO_433 (O_433,N_19984,N_19965);
nor UO_434 (O_434,N_19804,N_19774);
or UO_435 (O_435,N_19924,N_19884);
nor UO_436 (O_436,N_19908,N_19969);
nand UO_437 (O_437,N_19808,N_19842);
and UO_438 (O_438,N_19855,N_19818);
nor UO_439 (O_439,N_19767,N_19781);
nand UO_440 (O_440,N_19866,N_19862);
or UO_441 (O_441,N_19839,N_19814);
and UO_442 (O_442,N_19780,N_19911);
or UO_443 (O_443,N_19897,N_19816);
nor UO_444 (O_444,N_19905,N_19991);
nor UO_445 (O_445,N_19763,N_19852);
nor UO_446 (O_446,N_19789,N_19841);
nand UO_447 (O_447,N_19936,N_19885);
xor UO_448 (O_448,N_19772,N_19848);
nand UO_449 (O_449,N_19971,N_19944);
or UO_450 (O_450,N_19873,N_19911);
and UO_451 (O_451,N_19870,N_19780);
nor UO_452 (O_452,N_19892,N_19967);
nor UO_453 (O_453,N_19907,N_19843);
nand UO_454 (O_454,N_19984,N_19764);
and UO_455 (O_455,N_19925,N_19829);
nand UO_456 (O_456,N_19839,N_19882);
or UO_457 (O_457,N_19917,N_19787);
and UO_458 (O_458,N_19925,N_19817);
and UO_459 (O_459,N_19875,N_19936);
xor UO_460 (O_460,N_19798,N_19895);
and UO_461 (O_461,N_19958,N_19845);
or UO_462 (O_462,N_19939,N_19894);
or UO_463 (O_463,N_19916,N_19768);
or UO_464 (O_464,N_19762,N_19843);
and UO_465 (O_465,N_19963,N_19995);
or UO_466 (O_466,N_19773,N_19837);
nor UO_467 (O_467,N_19951,N_19945);
nand UO_468 (O_468,N_19817,N_19959);
nor UO_469 (O_469,N_19908,N_19928);
nor UO_470 (O_470,N_19931,N_19798);
or UO_471 (O_471,N_19938,N_19919);
or UO_472 (O_472,N_19984,N_19782);
nor UO_473 (O_473,N_19800,N_19806);
and UO_474 (O_474,N_19958,N_19862);
and UO_475 (O_475,N_19788,N_19910);
and UO_476 (O_476,N_19811,N_19903);
nor UO_477 (O_477,N_19833,N_19778);
and UO_478 (O_478,N_19989,N_19824);
nand UO_479 (O_479,N_19876,N_19757);
nor UO_480 (O_480,N_19921,N_19751);
or UO_481 (O_481,N_19899,N_19773);
nor UO_482 (O_482,N_19857,N_19828);
or UO_483 (O_483,N_19979,N_19766);
nand UO_484 (O_484,N_19856,N_19826);
nor UO_485 (O_485,N_19773,N_19810);
nor UO_486 (O_486,N_19850,N_19916);
or UO_487 (O_487,N_19751,N_19889);
xnor UO_488 (O_488,N_19860,N_19758);
and UO_489 (O_489,N_19788,N_19803);
nor UO_490 (O_490,N_19890,N_19786);
nor UO_491 (O_491,N_19792,N_19887);
and UO_492 (O_492,N_19941,N_19780);
or UO_493 (O_493,N_19791,N_19873);
nor UO_494 (O_494,N_19768,N_19877);
and UO_495 (O_495,N_19789,N_19819);
xor UO_496 (O_496,N_19857,N_19992);
nand UO_497 (O_497,N_19754,N_19796);
and UO_498 (O_498,N_19874,N_19991);
xor UO_499 (O_499,N_19944,N_19765);
nand UO_500 (O_500,N_19761,N_19843);
xnor UO_501 (O_501,N_19941,N_19973);
xnor UO_502 (O_502,N_19833,N_19978);
and UO_503 (O_503,N_19861,N_19853);
nor UO_504 (O_504,N_19951,N_19808);
and UO_505 (O_505,N_19951,N_19845);
nor UO_506 (O_506,N_19793,N_19771);
nor UO_507 (O_507,N_19765,N_19889);
nand UO_508 (O_508,N_19894,N_19975);
nor UO_509 (O_509,N_19948,N_19884);
nor UO_510 (O_510,N_19773,N_19788);
and UO_511 (O_511,N_19768,N_19782);
or UO_512 (O_512,N_19889,N_19912);
nor UO_513 (O_513,N_19786,N_19867);
or UO_514 (O_514,N_19879,N_19937);
nor UO_515 (O_515,N_19840,N_19951);
xor UO_516 (O_516,N_19934,N_19941);
or UO_517 (O_517,N_19836,N_19857);
or UO_518 (O_518,N_19940,N_19999);
nand UO_519 (O_519,N_19949,N_19963);
or UO_520 (O_520,N_19913,N_19921);
and UO_521 (O_521,N_19908,N_19865);
and UO_522 (O_522,N_19765,N_19933);
and UO_523 (O_523,N_19872,N_19994);
nand UO_524 (O_524,N_19881,N_19956);
nand UO_525 (O_525,N_19890,N_19887);
and UO_526 (O_526,N_19957,N_19900);
nand UO_527 (O_527,N_19959,N_19938);
and UO_528 (O_528,N_19794,N_19947);
and UO_529 (O_529,N_19945,N_19980);
and UO_530 (O_530,N_19824,N_19867);
nand UO_531 (O_531,N_19868,N_19827);
or UO_532 (O_532,N_19916,N_19825);
nand UO_533 (O_533,N_19978,N_19917);
or UO_534 (O_534,N_19899,N_19799);
or UO_535 (O_535,N_19791,N_19816);
nand UO_536 (O_536,N_19768,N_19784);
xnor UO_537 (O_537,N_19774,N_19789);
nand UO_538 (O_538,N_19899,N_19833);
nand UO_539 (O_539,N_19916,N_19998);
or UO_540 (O_540,N_19880,N_19774);
or UO_541 (O_541,N_19921,N_19794);
nand UO_542 (O_542,N_19999,N_19854);
or UO_543 (O_543,N_19892,N_19918);
or UO_544 (O_544,N_19968,N_19879);
or UO_545 (O_545,N_19814,N_19927);
nand UO_546 (O_546,N_19979,N_19838);
nor UO_547 (O_547,N_19823,N_19956);
nand UO_548 (O_548,N_19813,N_19963);
nand UO_549 (O_549,N_19818,N_19922);
nand UO_550 (O_550,N_19938,N_19918);
xnor UO_551 (O_551,N_19970,N_19887);
or UO_552 (O_552,N_19798,N_19936);
or UO_553 (O_553,N_19759,N_19855);
or UO_554 (O_554,N_19943,N_19869);
nor UO_555 (O_555,N_19760,N_19936);
nor UO_556 (O_556,N_19895,N_19978);
nand UO_557 (O_557,N_19797,N_19924);
nor UO_558 (O_558,N_19879,N_19995);
nor UO_559 (O_559,N_19913,N_19949);
or UO_560 (O_560,N_19803,N_19762);
or UO_561 (O_561,N_19895,N_19953);
and UO_562 (O_562,N_19944,N_19925);
nand UO_563 (O_563,N_19984,N_19763);
nor UO_564 (O_564,N_19889,N_19927);
and UO_565 (O_565,N_19840,N_19872);
or UO_566 (O_566,N_19915,N_19827);
or UO_567 (O_567,N_19769,N_19812);
or UO_568 (O_568,N_19996,N_19753);
or UO_569 (O_569,N_19914,N_19956);
or UO_570 (O_570,N_19937,N_19752);
and UO_571 (O_571,N_19936,N_19964);
nor UO_572 (O_572,N_19873,N_19921);
nand UO_573 (O_573,N_19985,N_19831);
and UO_574 (O_574,N_19978,N_19788);
and UO_575 (O_575,N_19797,N_19794);
xor UO_576 (O_576,N_19783,N_19756);
nand UO_577 (O_577,N_19972,N_19823);
or UO_578 (O_578,N_19946,N_19964);
nand UO_579 (O_579,N_19995,N_19873);
nor UO_580 (O_580,N_19911,N_19946);
and UO_581 (O_581,N_19807,N_19826);
or UO_582 (O_582,N_19948,N_19767);
and UO_583 (O_583,N_19809,N_19834);
nor UO_584 (O_584,N_19823,N_19915);
xnor UO_585 (O_585,N_19862,N_19769);
xnor UO_586 (O_586,N_19783,N_19950);
nand UO_587 (O_587,N_19890,N_19889);
and UO_588 (O_588,N_19804,N_19809);
and UO_589 (O_589,N_19769,N_19801);
and UO_590 (O_590,N_19808,N_19865);
nand UO_591 (O_591,N_19888,N_19827);
nand UO_592 (O_592,N_19936,N_19768);
nand UO_593 (O_593,N_19750,N_19771);
nor UO_594 (O_594,N_19835,N_19805);
nand UO_595 (O_595,N_19902,N_19874);
or UO_596 (O_596,N_19761,N_19763);
nand UO_597 (O_597,N_19855,N_19840);
or UO_598 (O_598,N_19954,N_19757);
and UO_599 (O_599,N_19761,N_19960);
xor UO_600 (O_600,N_19843,N_19923);
or UO_601 (O_601,N_19990,N_19868);
nand UO_602 (O_602,N_19966,N_19771);
or UO_603 (O_603,N_19825,N_19769);
and UO_604 (O_604,N_19963,N_19838);
nor UO_605 (O_605,N_19782,N_19850);
and UO_606 (O_606,N_19984,N_19883);
nor UO_607 (O_607,N_19909,N_19830);
nor UO_608 (O_608,N_19987,N_19774);
nand UO_609 (O_609,N_19916,N_19843);
or UO_610 (O_610,N_19763,N_19791);
nand UO_611 (O_611,N_19943,N_19860);
and UO_612 (O_612,N_19784,N_19850);
or UO_613 (O_613,N_19811,N_19919);
nor UO_614 (O_614,N_19866,N_19843);
xor UO_615 (O_615,N_19776,N_19897);
nand UO_616 (O_616,N_19906,N_19820);
and UO_617 (O_617,N_19840,N_19895);
nand UO_618 (O_618,N_19766,N_19948);
nand UO_619 (O_619,N_19966,N_19926);
or UO_620 (O_620,N_19785,N_19958);
or UO_621 (O_621,N_19843,N_19883);
or UO_622 (O_622,N_19787,N_19833);
xnor UO_623 (O_623,N_19773,N_19961);
or UO_624 (O_624,N_19907,N_19775);
and UO_625 (O_625,N_19877,N_19928);
and UO_626 (O_626,N_19910,N_19977);
nand UO_627 (O_627,N_19986,N_19821);
nand UO_628 (O_628,N_19846,N_19882);
nor UO_629 (O_629,N_19919,N_19851);
xor UO_630 (O_630,N_19982,N_19782);
nor UO_631 (O_631,N_19940,N_19961);
nand UO_632 (O_632,N_19947,N_19772);
and UO_633 (O_633,N_19861,N_19985);
nor UO_634 (O_634,N_19930,N_19960);
nor UO_635 (O_635,N_19850,N_19993);
nand UO_636 (O_636,N_19788,N_19982);
and UO_637 (O_637,N_19816,N_19832);
nor UO_638 (O_638,N_19798,N_19878);
nor UO_639 (O_639,N_19867,N_19996);
xnor UO_640 (O_640,N_19874,N_19808);
or UO_641 (O_641,N_19948,N_19913);
and UO_642 (O_642,N_19983,N_19911);
or UO_643 (O_643,N_19860,N_19766);
and UO_644 (O_644,N_19949,N_19800);
nand UO_645 (O_645,N_19834,N_19920);
nand UO_646 (O_646,N_19873,N_19931);
xor UO_647 (O_647,N_19836,N_19938);
nand UO_648 (O_648,N_19833,N_19972);
nand UO_649 (O_649,N_19835,N_19763);
nor UO_650 (O_650,N_19932,N_19759);
and UO_651 (O_651,N_19754,N_19797);
nor UO_652 (O_652,N_19835,N_19762);
nor UO_653 (O_653,N_19753,N_19948);
nor UO_654 (O_654,N_19849,N_19796);
nor UO_655 (O_655,N_19828,N_19907);
or UO_656 (O_656,N_19800,N_19899);
nor UO_657 (O_657,N_19771,N_19829);
nor UO_658 (O_658,N_19978,N_19918);
nor UO_659 (O_659,N_19947,N_19854);
and UO_660 (O_660,N_19753,N_19903);
and UO_661 (O_661,N_19941,N_19797);
and UO_662 (O_662,N_19808,N_19981);
or UO_663 (O_663,N_19980,N_19924);
or UO_664 (O_664,N_19920,N_19891);
nand UO_665 (O_665,N_19777,N_19878);
nand UO_666 (O_666,N_19877,N_19930);
or UO_667 (O_667,N_19934,N_19973);
nand UO_668 (O_668,N_19920,N_19959);
nor UO_669 (O_669,N_19799,N_19862);
xnor UO_670 (O_670,N_19873,N_19773);
and UO_671 (O_671,N_19953,N_19794);
nor UO_672 (O_672,N_19932,N_19811);
and UO_673 (O_673,N_19857,N_19933);
xnor UO_674 (O_674,N_19908,N_19805);
and UO_675 (O_675,N_19785,N_19861);
and UO_676 (O_676,N_19780,N_19904);
nand UO_677 (O_677,N_19816,N_19945);
nor UO_678 (O_678,N_19767,N_19850);
or UO_679 (O_679,N_19820,N_19815);
xor UO_680 (O_680,N_19841,N_19768);
or UO_681 (O_681,N_19756,N_19842);
nor UO_682 (O_682,N_19978,N_19904);
xor UO_683 (O_683,N_19787,N_19870);
and UO_684 (O_684,N_19766,N_19943);
nand UO_685 (O_685,N_19907,N_19855);
xor UO_686 (O_686,N_19942,N_19809);
nor UO_687 (O_687,N_19808,N_19923);
or UO_688 (O_688,N_19952,N_19796);
and UO_689 (O_689,N_19981,N_19901);
xnor UO_690 (O_690,N_19852,N_19832);
nor UO_691 (O_691,N_19928,N_19925);
nor UO_692 (O_692,N_19872,N_19798);
or UO_693 (O_693,N_19793,N_19756);
or UO_694 (O_694,N_19983,N_19761);
nor UO_695 (O_695,N_19982,N_19957);
nand UO_696 (O_696,N_19806,N_19995);
and UO_697 (O_697,N_19900,N_19847);
nand UO_698 (O_698,N_19865,N_19772);
and UO_699 (O_699,N_19790,N_19953);
and UO_700 (O_700,N_19898,N_19855);
xor UO_701 (O_701,N_19878,N_19968);
or UO_702 (O_702,N_19916,N_19854);
nand UO_703 (O_703,N_19994,N_19783);
nor UO_704 (O_704,N_19848,N_19836);
and UO_705 (O_705,N_19905,N_19936);
or UO_706 (O_706,N_19780,N_19849);
and UO_707 (O_707,N_19750,N_19952);
or UO_708 (O_708,N_19811,N_19942);
nor UO_709 (O_709,N_19869,N_19751);
nand UO_710 (O_710,N_19995,N_19813);
or UO_711 (O_711,N_19948,N_19994);
nand UO_712 (O_712,N_19938,N_19903);
nor UO_713 (O_713,N_19886,N_19884);
nor UO_714 (O_714,N_19857,N_19833);
nand UO_715 (O_715,N_19976,N_19959);
nor UO_716 (O_716,N_19870,N_19863);
nor UO_717 (O_717,N_19924,N_19997);
and UO_718 (O_718,N_19769,N_19911);
and UO_719 (O_719,N_19806,N_19906);
and UO_720 (O_720,N_19860,N_19813);
nand UO_721 (O_721,N_19833,N_19895);
nand UO_722 (O_722,N_19830,N_19978);
and UO_723 (O_723,N_19800,N_19793);
nand UO_724 (O_724,N_19972,N_19889);
nand UO_725 (O_725,N_19847,N_19930);
and UO_726 (O_726,N_19829,N_19996);
nor UO_727 (O_727,N_19930,N_19798);
or UO_728 (O_728,N_19904,N_19960);
or UO_729 (O_729,N_19912,N_19943);
and UO_730 (O_730,N_19752,N_19931);
or UO_731 (O_731,N_19936,N_19896);
and UO_732 (O_732,N_19947,N_19758);
nor UO_733 (O_733,N_19869,N_19835);
nand UO_734 (O_734,N_19786,N_19800);
and UO_735 (O_735,N_19796,N_19838);
and UO_736 (O_736,N_19853,N_19780);
nor UO_737 (O_737,N_19917,N_19984);
and UO_738 (O_738,N_19767,N_19899);
nor UO_739 (O_739,N_19922,N_19939);
and UO_740 (O_740,N_19890,N_19855);
or UO_741 (O_741,N_19838,N_19942);
or UO_742 (O_742,N_19952,N_19901);
nand UO_743 (O_743,N_19922,N_19949);
and UO_744 (O_744,N_19915,N_19794);
nand UO_745 (O_745,N_19812,N_19986);
and UO_746 (O_746,N_19928,N_19849);
or UO_747 (O_747,N_19831,N_19865);
nor UO_748 (O_748,N_19832,N_19795);
and UO_749 (O_749,N_19804,N_19820);
or UO_750 (O_750,N_19909,N_19968);
and UO_751 (O_751,N_19899,N_19973);
nor UO_752 (O_752,N_19786,N_19985);
nand UO_753 (O_753,N_19869,N_19904);
nor UO_754 (O_754,N_19842,N_19789);
or UO_755 (O_755,N_19827,N_19991);
nor UO_756 (O_756,N_19991,N_19923);
or UO_757 (O_757,N_19908,N_19992);
nor UO_758 (O_758,N_19760,N_19915);
or UO_759 (O_759,N_19922,N_19998);
and UO_760 (O_760,N_19869,N_19782);
xnor UO_761 (O_761,N_19854,N_19907);
nand UO_762 (O_762,N_19768,N_19844);
nor UO_763 (O_763,N_19974,N_19941);
and UO_764 (O_764,N_19903,N_19796);
and UO_765 (O_765,N_19896,N_19923);
xnor UO_766 (O_766,N_19864,N_19782);
and UO_767 (O_767,N_19895,N_19763);
xor UO_768 (O_768,N_19816,N_19960);
or UO_769 (O_769,N_19774,N_19998);
and UO_770 (O_770,N_19797,N_19945);
or UO_771 (O_771,N_19857,N_19776);
nand UO_772 (O_772,N_19768,N_19783);
xnor UO_773 (O_773,N_19880,N_19779);
and UO_774 (O_774,N_19908,N_19975);
xor UO_775 (O_775,N_19823,N_19817);
nor UO_776 (O_776,N_19930,N_19982);
or UO_777 (O_777,N_19857,N_19846);
nand UO_778 (O_778,N_19834,N_19922);
nor UO_779 (O_779,N_19799,N_19990);
xor UO_780 (O_780,N_19884,N_19772);
nor UO_781 (O_781,N_19861,N_19937);
and UO_782 (O_782,N_19889,N_19903);
nor UO_783 (O_783,N_19780,N_19987);
nor UO_784 (O_784,N_19906,N_19826);
nand UO_785 (O_785,N_19786,N_19779);
or UO_786 (O_786,N_19755,N_19776);
nor UO_787 (O_787,N_19958,N_19765);
xnor UO_788 (O_788,N_19973,N_19759);
nor UO_789 (O_789,N_19871,N_19915);
nand UO_790 (O_790,N_19891,N_19791);
or UO_791 (O_791,N_19949,N_19872);
nor UO_792 (O_792,N_19825,N_19778);
and UO_793 (O_793,N_19969,N_19774);
or UO_794 (O_794,N_19795,N_19903);
nand UO_795 (O_795,N_19796,N_19779);
and UO_796 (O_796,N_19828,N_19941);
xor UO_797 (O_797,N_19791,N_19885);
xor UO_798 (O_798,N_19949,N_19876);
and UO_799 (O_799,N_19896,N_19960);
and UO_800 (O_800,N_19846,N_19945);
nand UO_801 (O_801,N_19927,N_19780);
nor UO_802 (O_802,N_19842,N_19978);
or UO_803 (O_803,N_19872,N_19894);
xnor UO_804 (O_804,N_19983,N_19903);
nand UO_805 (O_805,N_19966,N_19878);
nand UO_806 (O_806,N_19780,N_19814);
and UO_807 (O_807,N_19752,N_19775);
and UO_808 (O_808,N_19785,N_19928);
or UO_809 (O_809,N_19877,N_19824);
and UO_810 (O_810,N_19956,N_19994);
nand UO_811 (O_811,N_19852,N_19901);
and UO_812 (O_812,N_19787,N_19857);
xnor UO_813 (O_813,N_19947,N_19839);
or UO_814 (O_814,N_19934,N_19932);
or UO_815 (O_815,N_19757,N_19980);
nor UO_816 (O_816,N_19968,N_19828);
and UO_817 (O_817,N_19762,N_19879);
nand UO_818 (O_818,N_19808,N_19780);
nand UO_819 (O_819,N_19879,N_19775);
xnor UO_820 (O_820,N_19945,N_19843);
or UO_821 (O_821,N_19939,N_19758);
and UO_822 (O_822,N_19913,N_19834);
nand UO_823 (O_823,N_19918,N_19776);
or UO_824 (O_824,N_19944,N_19847);
nand UO_825 (O_825,N_19843,N_19960);
xor UO_826 (O_826,N_19951,N_19820);
nor UO_827 (O_827,N_19809,N_19794);
xnor UO_828 (O_828,N_19893,N_19755);
nor UO_829 (O_829,N_19777,N_19852);
and UO_830 (O_830,N_19853,N_19986);
or UO_831 (O_831,N_19852,N_19819);
and UO_832 (O_832,N_19852,N_19892);
xor UO_833 (O_833,N_19923,N_19929);
xor UO_834 (O_834,N_19987,N_19755);
xnor UO_835 (O_835,N_19899,N_19882);
or UO_836 (O_836,N_19926,N_19875);
nand UO_837 (O_837,N_19795,N_19822);
nand UO_838 (O_838,N_19791,N_19888);
nor UO_839 (O_839,N_19930,N_19814);
and UO_840 (O_840,N_19907,N_19957);
or UO_841 (O_841,N_19971,N_19958);
xor UO_842 (O_842,N_19815,N_19764);
nor UO_843 (O_843,N_19915,N_19933);
or UO_844 (O_844,N_19995,N_19944);
nor UO_845 (O_845,N_19909,N_19983);
or UO_846 (O_846,N_19909,N_19953);
or UO_847 (O_847,N_19777,N_19845);
nor UO_848 (O_848,N_19872,N_19818);
and UO_849 (O_849,N_19922,N_19975);
nand UO_850 (O_850,N_19947,N_19994);
nand UO_851 (O_851,N_19831,N_19935);
and UO_852 (O_852,N_19985,N_19841);
and UO_853 (O_853,N_19825,N_19776);
and UO_854 (O_854,N_19970,N_19976);
and UO_855 (O_855,N_19957,N_19788);
and UO_856 (O_856,N_19971,N_19777);
nor UO_857 (O_857,N_19827,N_19762);
nand UO_858 (O_858,N_19770,N_19771);
or UO_859 (O_859,N_19931,N_19849);
or UO_860 (O_860,N_19972,N_19947);
nor UO_861 (O_861,N_19867,N_19904);
xor UO_862 (O_862,N_19955,N_19798);
nand UO_863 (O_863,N_19823,N_19953);
nand UO_864 (O_864,N_19924,N_19983);
xor UO_865 (O_865,N_19766,N_19919);
or UO_866 (O_866,N_19861,N_19812);
nand UO_867 (O_867,N_19820,N_19977);
nand UO_868 (O_868,N_19849,N_19894);
and UO_869 (O_869,N_19985,N_19864);
or UO_870 (O_870,N_19892,N_19973);
nand UO_871 (O_871,N_19860,N_19993);
nand UO_872 (O_872,N_19916,N_19932);
and UO_873 (O_873,N_19814,N_19821);
nand UO_874 (O_874,N_19944,N_19933);
or UO_875 (O_875,N_19820,N_19832);
or UO_876 (O_876,N_19897,N_19779);
nand UO_877 (O_877,N_19923,N_19794);
nand UO_878 (O_878,N_19765,N_19894);
and UO_879 (O_879,N_19883,N_19891);
nor UO_880 (O_880,N_19836,N_19757);
nand UO_881 (O_881,N_19884,N_19848);
nor UO_882 (O_882,N_19841,N_19843);
and UO_883 (O_883,N_19759,N_19865);
or UO_884 (O_884,N_19795,N_19938);
and UO_885 (O_885,N_19906,N_19955);
nand UO_886 (O_886,N_19866,N_19977);
nand UO_887 (O_887,N_19997,N_19947);
and UO_888 (O_888,N_19941,N_19758);
xor UO_889 (O_889,N_19919,N_19822);
nand UO_890 (O_890,N_19772,N_19891);
and UO_891 (O_891,N_19933,N_19757);
nor UO_892 (O_892,N_19782,N_19993);
xnor UO_893 (O_893,N_19787,N_19792);
or UO_894 (O_894,N_19810,N_19844);
nand UO_895 (O_895,N_19952,N_19832);
and UO_896 (O_896,N_19833,N_19854);
and UO_897 (O_897,N_19867,N_19784);
and UO_898 (O_898,N_19859,N_19925);
nor UO_899 (O_899,N_19985,N_19796);
or UO_900 (O_900,N_19795,N_19773);
and UO_901 (O_901,N_19869,N_19965);
nor UO_902 (O_902,N_19847,N_19850);
nor UO_903 (O_903,N_19830,N_19848);
xnor UO_904 (O_904,N_19851,N_19989);
xor UO_905 (O_905,N_19802,N_19758);
nand UO_906 (O_906,N_19988,N_19796);
and UO_907 (O_907,N_19954,N_19837);
nand UO_908 (O_908,N_19998,N_19975);
nand UO_909 (O_909,N_19820,N_19859);
nand UO_910 (O_910,N_19946,N_19805);
and UO_911 (O_911,N_19783,N_19792);
nor UO_912 (O_912,N_19786,N_19805);
or UO_913 (O_913,N_19933,N_19927);
or UO_914 (O_914,N_19946,N_19827);
nand UO_915 (O_915,N_19994,N_19851);
nor UO_916 (O_916,N_19944,N_19894);
nor UO_917 (O_917,N_19759,N_19874);
nand UO_918 (O_918,N_19886,N_19936);
xor UO_919 (O_919,N_19852,N_19895);
nand UO_920 (O_920,N_19896,N_19790);
and UO_921 (O_921,N_19792,N_19972);
nor UO_922 (O_922,N_19793,N_19829);
nor UO_923 (O_923,N_19799,N_19959);
nand UO_924 (O_924,N_19793,N_19965);
nand UO_925 (O_925,N_19802,N_19922);
or UO_926 (O_926,N_19831,N_19863);
or UO_927 (O_927,N_19753,N_19951);
nand UO_928 (O_928,N_19965,N_19858);
nor UO_929 (O_929,N_19993,N_19832);
nor UO_930 (O_930,N_19804,N_19791);
nor UO_931 (O_931,N_19844,N_19992);
nor UO_932 (O_932,N_19944,N_19848);
nor UO_933 (O_933,N_19979,N_19812);
nor UO_934 (O_934,N_19812,N_19922);
and UO_935 (O_935,N_19772,N_19771);
nand UO_936 (O_936,N_19932,N_19989);
and UO_937 (O_937,N_19899,N_19896);
or UO_938 (O_938,N_19915,N_19839);
or UO_939 (O_939,N_19921,N_19962);
or UO_940 (O_940,N_19886,N_19828);
nand UO_941 (O_941,N_19819,N_19757);
xnor UO_942 (O_942,N_19782,N_19845);
xor UO_943 (O_943,N_19838,N_19758);
and UO_944 (O_944,N_19978,N_19803);
nand UO_945 (O_945,N_19831,N_19928);
nor UO_946 (O_946,N_19948,N_19764);
nor UO_947 (O_947,N_19796,N_19894);
nor UO_948 (O_948,N_19814,N_19867);
or UO_949 (O_949,N_19860,N_19961);
and UO_950 (O_950,N_19931,N_19760);
nand UO_951 (O_951,N_19807,N_19798);
nand UO_952 (O_952,N_19993,N_19990);
and UO_953 (O_953,N_19973,N_19914);
or UO_954 (O_954,N_19817,N_19809);
xor UO_955 (O_955,N_19909,N_19759);
nor UO_956 (O_956,N_19867,N_19783);
nand UO_957 (O_957,N_19866,N_19871);
and UO_958 (O_958,N_19887,N_19865);
nor UO_959 (O_959,N_19886,N_19760);
and UO_960 (O_960,N_19872,N_19942);
nand UO_961 (O_961,N_19995,N_19942);
and UO_962 (O_962,N_19866,N_19910);
nand UO_963 (O_963,N_19812,N_19903);
nand UO_964 (O_964,N_19759,N_19840);
and UO_965 (O_965,N_19765,N_19973);
or UO_966 (O_966,N_19774,N_19943);
or UO_967 (O_967,N_19806,N_19894);
or UO_968 (O_968,N_19769,N_19839);
nor UO_969 (O_969,N_19780,N_19977);
and UO_970 (O_970,N_19986,N_19762);
nor UO_971 (O_971,N_19806,N_19936);
and UO_972 (O_972,N_19999,N_19894);
nor UO_973 (O_973,N_19965,N_19790);
and UO_974 (O_974,N_19784,N_19915);
nor UO_975 (O_975,N_19827,N_19849);
and UO_976 (O_976,N_19863,N_19829);
nand UO_977 (O_977,N_19961,N_19833);
nand UO_978 (O_978,N_19914,N_19796);
or UO_979 (O_979,N_19886,N_19969);
xnor UO_980 (O_980,N_19900,N_19851);
nand UO_981 (O_981,N_19763,N_19995);
and UO_982 (O_982,N_19949,N_19937);
nand UO_983 (O_983,N_19881,N_19842);
nand UO_984 (O_984,N_19770,N_19919);
and UO_985 (O_985,N_19858,N_19892);
nor UO_986 (O_986,N_19869,N_19779);
nand UO_987 (O_987,N_19759,N_19933);
and UO_988 (O_988,N_19760,N_19960);
or UO_989 (O_989,N_19959,N_19826);
nand UO_990 (O_990,N_19975,N_19895);
or UO_991 (O_991,N_19903,N_19790);
and UO_992 (O_992,N_19987,N_19891);
nor UO_993 (O_993,N_19863,N_19855);
nand UO_994 (O_994,N_19787,N_19853);
or UO_995 (O_995,N_19918,N_19841);
nand UO_996 (O_996,N_19807,N_19820);
or UO_997 (O_997,N_19851,N_19779);
nor UO_998 (O_998,N_19818,N_19779);
nor UO_999 (O_999,N_19856,N_19978);
nand UO_1000 (O_1000,N_19967,N_19926);
or UO_1001 (O_1001,N_19949,N_19878);
or UO_1002 (O_1002,N_19799,N_19962);
or UO_1003 (O_1003,N_19802,N_19972);
nor UO_1004 (O_1004,N_19796,N_19964);
nor UO_1005 (O_1005,N_19873,N_19909);
and UO_1006 (O_1006,N_19984,N_19955);
nor UO_1007 (O_1007,N_19897,N_19870);
nand UO_1008 (O_1008,N_19823,N_19874);
nor UO_1009 (O_1009,N_19827,N_19764);
nand UO_1010 (O_1010,N_19911,N_19827);
or UO_1011 (O_1011,N_19992,N_19859);
or UO_1012 (O_1012,N_19797,N_19811);
xor UO_1013 (O_1013,N_19777,N_19944);
and UO_1014 (O_1014,N_19793,N_19971);
and UO_1015 (O_1015,N_19984,N_19865);
or UO_1016 (O_1016,N_19828,N_19956);
nand UO_1017 (O_1017,N_19932,N_19775);
xor UO_1018 (O_1018,N_19862,N_19914);
and UO_1019 (O_1019,N_19816,N_19878);
nand UO_1020 (O_1020,N_19925,N_19947);
or UO_1021 (O_1021,N_19843,N_19751);
and UO_1022 (O_1022,N_19972,N_19844);
nand UO_1023 (O_1023,N_19920,N_19778);
or UO_1024 (O_1024,N_19838,N_19818);
xnor UO_1025 (O_1025,N_19911,N_19850);
or UO_1026 (O_1026,N_19813,N_19949);
nor UO_1027 (O_1027,N_19807,N_19914);
or UO_1028 (O_1028,N_19824,N_19820);
or UO_1029 (O_1029,N_19833,N_19808);
nor UO_1030 (O_1030,N_19946,N_19810);
nor UO_1031 (O_1031,N_19835,N_19940);
nand UO_1032 (O_1032,N_19997,N_19961);
and UO_1033 (O_1033,N_19875,N_19846);
or UO_1034 (O_1034,N_19807,N_19957);
nand UO_1035 (O_1035,N_19908,N_19824);
and UO_1036 (O_1036,N_19842,N_19775);
or UO_1037 (O_1037,N_19908,N_19915);
and UO_1038 (O_1038,N_19859,N_19906);
nor UO_1039 (O_1039,N_19929,N_19932);
or UO_1040 (O_1040,N_19949,N_19790);
nand UO_1041 (O_1041,N_19852,N_19787);
nor UO_1042 (O_1042,N_19948,N_19988);
or UO_1043 (O_1043,N_19909,N_19901);
nor UO_1044 (O_1044,N_19999,N_19847);
or UO_1045 (O_1045,N_19994,N_19927);
and UO_1046 (O_1046,N_19809,N_19879);
xor UO_1047 (O_1047,N_19924,N_19927);
or UO_1048 (O_1048,N_19763,N_19987);
nand UO_1049 (O_1049,N_19925,N_19971);
or UO_1050 (O_1050,N_19756,N_19880);
nor UO_1051 (O_1051,N_19808,N_19863);
or UO_1052 (O_1052,N_19774,N_19946);
nand UO_1053 (O_1053,N_19982,N_19780);
nor UO_1054 (O_1054,N_19880,N_19841);
and UO_1055 (O_1055,N_19775,N_19997);
nor UO_1056 (O_1056,N_19804,N_19944);
nor UO_1057 (O_1057,N_19804,N_19766);
nand UO_1058 (O_1058,N_19999,N_19934);
or UO_1059 (O_1059,N_19994,N_19878);
and UO_1060 (O_1060,N_19858,N_19889);
and UO_1061 (O_1061,N_19869,N_19790);
nand UO_1062 (O_1062,N_19915,N_19907);
nand UO_1063 (O_1063,N_19936,N_19894);
and UO_1064 (O_1064,N_19857,N_19942);
nor UO_1065 (O_1065,N_19769,N_19779);
nor UO_1066 (O_1066,N_19937,N_19961);
and UO_1067 (O_1067,N_19888,N_19886);
or UO_1068 (O_1068,N_19924,N_19912);
and UO_1069 (O_1069,N_19895,N_19829);
or UO_1070 (O_1070,N_19991,N_19765);
and UO_1071 (O_1071,N_19806,N_19944);
or UO_1072 (O_1072,N_19982,N_19927);
nand UO_1073 (O_1073,N_19940,N_19966);
nand UO_1074 (O_1074,N_19927,N_19873);
and UO_1075 (O_1075,N_19786,N_19771);
nor UO_1076 (O_1076,N_19833,N_19844);
nor UO_1077 (O_1077,N_19917,N_19845);
or UO_1078 (O_1078,N_19879,N_19910);
or UO_1079 (O_1079,N_19847,N_19869);
and UO_1080 (O_1080,N_19888,N_19923);
and UO_1081 (O_1081,N_19885,N_19844);
nor UO_1082 (O_1082,N_19762,N_19896);
nor UO_1083 (O_1083,N_19766,N_19954);
nor UO_1084 (O_1084,N_19966,N_19817);
nand UO_1085 (O_1085,N_19953,N_19888);
nor UO_1086 (O_1086,N_19984,N_19809);
nor UO_1087 (O_1087,N_19957,N_19969);
or UO_1088 (O_1088,N_19960,N_19979);
nand UO_1089 (O_1089,N_19898,N_19854);
and UO_1090 (O_1090,N_19845,N_19979);
and UO_1091 (O_1091,N_19772,N_19837);
nand UO_1092 (O_1092,N_19766,N_19848);
and UO_1093 (O_1093,N_19948,N_19893);
and UO_1094 (O_1094,N_19931,N_19783);
and UO_1095 (O_1095,N_19778,N_19782);
nand UO_1096 (O_1096,N_19957,N_19816);
or UO_1097 (O_1097,N_19858,N_19855);
and UO_1098 (O_1098,N_19973,N_19868);
nand UO_1099 (O_1099,N_19836,N_19844);
and UO_1100 (O_1100,N_19833,N_19836);
or UO_1101 (O_1101,N_19903,N_19878);
or UO_1102 (O_1102,N_19947,N_19829);
or UO_1103 (O_1103,N_19945,N_19881);
or UO_1104 (O_1104,N_19830,N_19777);
xnor UO_1105 (O_1105,N_19966,N_19866);
and UO_1106 (O_1106,N_19871,N_19808);
nor UO_1107 (O_1107,N_19776,N_19933);
xor UO_1108 (O_1108,N_19769,N_19964);
nor UO_1109 (O_1109,N_19784,N_19871);
and UO_1110 (O_1110,N_19912,N_19918);
and UO_1111 (O_1111,N_19809,N_19867);
and UO_1112 (O_1112,N_19826,N_19974);
nor UO_1113 (O_1113,N_19833,N_19928);
or UO_1114 (O_1114,N_19976,N_19847);
nand UO_1115 (O_1115,N_19984,N_19972);
or UO_1116 (O_1116,N_19789,N_19990);
or UO_1117 (O_1117,N_19859,N_19950);
xnor UO_1118 (O_1118,N_19953,N_19901);
nor UO_1119 (O_1119,N_19814,N_19952);
nor UO_1120 (O_1120,N_19833,N_19758);
nand UO_1121 (O_1121,N_19988,N_19763);
and UO_1122 (O_1122,N_19953,N_19937);
nor UO_1123 (O_1123,N_19898,N_19843);
or UO_1124 (O_1124,N_19957,N_19844);
nor UO_1125 (O_1125,N_19797,N_19787);
nand UO_1126 (O_1126,N_19917,N_19761);
and UO_1127 (O_1127,N_19897,N_19784);
and UO_1128 (O_1128,N_19773,N_19803);
nand UO_1129 (O_1129,N_19820,N_19868);
nor UO_1130 (O_1130,N_19787,N_19915);
xnor UO_1131 (O_1131,N_19778,N_19949);
and UO_1132 (O_1132,N_19997,N_19880);
and UO_1133 (O_1133,N_19782,N_19780);
nand UO_1134 (O_1134,N_19846,N_19789);
or UO_1135 (O_1135,N_19820,N_19943);
nor UO_1136 (O_1136,N_19865,N_19955);
or UO_1137 (O_1137,N_19937,N_19857);
xnor UO_1138 (O_1138,N_19788,N_19828);
and UO_1139 (O_1139,N_19949,N_19903);
nand UO_1140 (O_1140,N_19943,N_19942);
and UO_1141 (O_1141,N_19953,N_19920);
nor UO_1142 (O_1142,N_19962,N_19770);
or UO_1143 (O_1143,N_19852,N_19781);
or UO_1144 (O_1144,N_19775,N_19755);
or UO_1145 (O_1145,N_19856,N_19986);
nand UO_1146 (O_1146,N_19862,N_19980);
nand UO_1147 (O_1147,N_19752,N_19970);
and UO_1148 (O_1148,N_19822,N_19858);
xnor UO_1149 (O_1149,N_19917,N_19758);
and UO_1150 (O_1150,N_19936,N_19780);
nor UO_1151 (O_1151,N_19919,N_19884);
nand UO_1152 (O_1152,N_19879,N_19854);
and UO_1153 (O_1153,N_19813,N_19830);
or UO_1154 (O_1154,N_19785,N_19881);
and UO_1155 (O_1155,N_19993,N_19937);
or UO_1156 (O_1156,N_19996,N_19921);
nor UO_1157 (O_1157,N_19787,N_19765);
xor UO_1158 (O_1158,N_19811,N_19965);
and UO_1159 (O_1159,N_19986,N_19916);
and UO_1160 (O_1160,N_19827,N_19912);
nor UO_1161 (O_1161,N_19778,N_19760);
nand UO_1162 (O_1162,N_19940,N_19974);
nand UO_1163 (O_1163,N_19843,N_19937);
nand UO_1164 (O_1164,N_19845,N_19947);
nand UO_1165 (O_1165,N_19986,N_19822);
nor UO_1166 (O_1166,N_19815,N_19892);
xor UO_1167 (O_1167,N_19929,N_19854);
nor UO_1168 (O_1168,N_19808,N_19986);
nor UO_1169 (O_1169,N_19823,N_19884);
nor UO_1170 (O_1170,N_19993,N_19822);
nand UO_1171 (O_1171,N_19835,N_19779);
nor UO_1172 (O_1172,N_19804,N_19943);
and UO_1173 (O_1173,N_19866,N_19961);
and UO_1174 (O_1174,N_19960,N_19765);
nand UO_1175 (O_1175,N_19885,N_19993);
or UO_1176 (O_1176,N_19757,N_19784);
nor UO_1177 (O_1177,N_19959,N_19766);
nand UO_1178 (O_1178,N_19901,N_19982);
or UO_1179 (O_1179,N_19823,N_19976);
and UO_1180 (O_1180,N_19795,N_19965);
nand UO_1181 (O_1181,N_19770,N_19815);
or UO_1182 (O_1182,N_19935,N_19830);
xnor UO_1183 (O_1183,N_19909,N_19826);
or UO_1184 (O_1184,N_19914,N_19779);
or UO_1185 (O_1185,N_19857,N_19974);
nor UO_1186 (O_1186,N_19966,N_19758);
or UO_1187 (O_1187,N_19957,N_19978);
and UO_1188 (O_1188,N_19779,N_19844);
nor UO_1189 (O_1189,N_19863,N_19848);
and UO_1190 (O_1190,N_19949,N_19822);
nor UO_1191 (O_1191,N_19872,N_19958);
nand UO_1192 (O_1192,N_19968,N_19782);
nand UO_1193 (O_1193,N_19971,N_19784);
or UO_1194 (O_1194,N_19810,N_19892);
nor UO_1195 (O_1195,N_19924,N_19767);
nor UO_1196 (O_1196,N_19937,N_19839);
xor UO_1197 (O_1197,N_19761,N_19945);
nand UO_1198 (O_1198,N_19766,N_19945);
or UO_1199 (O_1199,N_19886,N_19874);
nand UO_1200 (O_1200,N_19874,N_19765);
nand UO_1201 (O_1201,N_19849,N_19836);
and UO_1202 (O_1202,N_19948,N_19962);
nand UO_1203 (O_1203,N_19993,N_19851);
xnor UO_1204 (O_1204,N_19985,N_19895);
or UO_1205 (O_1205,N_19787,N_19776);
nand UO_1206 (O_1206,N_19817,N_19912);
and UO_1207 (O_1207,N_19944,N_19815);
and UO_1208 (O_1208,N_19990,N_19856);
and UO_1209 (O_1209,N_19983,N_19762);
or UO_1210 (O_1210,N_19757,N_19837);
nand UO_1211 (O_1211,N_19774,N_19918);
xnor UO_1212 (O_1212,N_19869,N_19946);
nand UO_1213 (O_1213,N_19767,N_19938);
nor UO_1214 (O_1214,N_19922,N_19794);
or UO_1215 (O_1215,N_19849,N_19882);
nor UO_1216 (O_1216,N_19887,N_19776);
nand UO_1217 (O_1217,N_19969,N_19854);
and UO_1218 (O_1218,N_19754,N_19901);
nand UO_1219 (O_1219,N_19868,N_19929);
nand UO_1220 (O_1220,N_19927,N_19839);
and UO_1221 (O_1221,N_19863,N_19873);
nor UO_1222 (O_1222,N_19873,N_19924);
and UO_1223 (O_1223,N_19989,N_19887);
nor UO_1224 (O_1224,N_19947,N_19929);
or UO_1225 (O_1225,N_19943,N_19995);
and UO_1226 (O_1226,N_19928,N_19774);
or UO_1227 (O_1227,N_19769,N_19844);
and UO_1228 (O_1228,N_19917,N_19770);
nor UO_1229 (O_1229,N_19941,N_19977);
and UO_1230 (O_1230,N_19936,N_19950);
xnor UO_1231 (O_1231,N_19924,N_19801);
xor UO_1232 (O_1232,N_19943,N_19992);
and UO_1233 (O_1233,N_19863,N_19797);
and UO_1234 (O_1234,N_19900,N_19980);
nand UO_1235 (O_1235,N_19953,N_19824);
nor UO_1236 (O_1236,N_19955,N_19924);
nor UO_1237 (O_1237,N_19960,N_19906);
and UO_1238 (O_1238,N_19968,N_19765);
nand UO_1239 (O_1239,N_19909,N_19936);
and UO_1240 (O_1240,N_19803,N_19755);
nand UO_1241 (O_1241,N_19848,N_19959);
nor UO_1242 (O_1242,N_19804,N_19923);
or UO_1243 (O_1243,N_19835,N_19798);
nand UO_1244 (O_1244,N_19827,N_19810);
and UO_1245 (O_1245,N_19811,N_19842);
or UO_1246 (O_1246,N_19800,N_19850);
nand UO_1247 (O_1247,N_19992,N_19951);
nand UO_1248 (O_1248,N_19831,N_19838);
xnor UO_1249 (O_1249,N_19854,N_19817);
nand UO_1250 (O_1250,N_19831,N_19976);
xor UO_1251 (O_1251,N_19936,N_19897);
nor UO_1252 (O_1252,N_19812,N_19778);
nor UO_1253 (O_1253,N_19986,N_19900);
nor UO_1254 (O_1254,N_19940,N_19900);
nand UO_1255 (O_1255,N_19874,N_19813);
nand UO_1256 (O_1256,N_19941,N_19946);
nor UO_1257 (O_1257,N_19878,N_19909);
or UO_1258 (O_1258,N_19826,N_19842);
xor UO_1259 (O_1259,N_19811,N_19841);
nor UO_1260 (O_1260,N_19812,N_19760);
or UO_1261 (O_1261,N_19845,N_19936);
nor UO_1262 (O_1262,N_19766,N_19985);
and UO_1263 (O_1263,N_19911,N_19797);
xnor UO_1264 (O_1264,N_19776,N_19773);
nand UO_1265 (O_1265,N_19833,N_19947);
nor UO_1266 (O_1266,N_19979,N_19854);
nor UO_1267 (O_1267,N_19795,N_19896);
or UO_1268 (O_1268,N_19760,N_19854);
or UO_1269 (O_1269,N_19778,N_19830);
and UO_1270 (O_1270,N_19888,N_19947);
or UO_1271 (O_1271,N_19953,N_19777);
nand UO_1272 (O_1272,N_19878,N_19826);
and UO_1273 (O_1273,N_19798,N_19842);
nor UO_1274 (O_1274,N_19911,N_19845);
or UO_1275 (O_1275,N_19752,N_19945);
nor UO_1276 (O_1276,N_19819,N_19988);
or UO_1277 (O_1277,N_19831,N_19846);
nand UO_1278 (O_1278,N_19841,N_19964);
nor UO_1279 (O_1279,N_19835,N_19846);
and UO_1280 (O_1280,N_19761,N_19793);
and UO_1281 (O_1281,N_19986,N_19828);
and UO_1282 (O_1282,N_19764,N_19803);
nand UO_1283 (O_1283,N_19946,N_19950);
and UO_1284 (O_1284,N_19814,N_19788);
or UO_1285 (O_1285,N_19869,N_19863);
nor UO_1286 (O_1286,N_19768,N_19779);
nor UO_1287 (O_1287,N_19949,N_19917);
or UO_1288 (O_1288,N_19886,N_19981);
and UO_1289 (O_1289,N_19966,N_19753);
xor UO_1290 (O_1290,N_19807,N_19855);
and UO_1291 (O_1291,N_19891,N_19989);
or UO_1292 (O_1292,N_19973,N_19911);
nor UO_1293 (O_1293,N_19798,N_19801);
nor UO_1294 (O_1294,N_19860,N_19862);
nor UO_1295 (O_1295,N_19907,N_19983);
or UO_1296 (O_1296,N_19886,N_19983);
nor UO_1297 (O_1297,N_19868,N_19810);
or UO_1298 (O_1298,N_19821,N_19944);
xnor UO_1299 (O_1299,N_19815,N_19798);
nand UO_1300 (O_1300,N_19845,N_19985);
and UO_1301 (O_1301,N_19951,N_19985);
or UO_1302 (O_1302,N_19853,N_19920);
or UO_1303 (O_1303,N_19889,N_19921);
or UO_1304 (O_1304,N_19853,N_19913);
or UO_1305 (O_1305,N_19972,N_19763);
and UO_1306 (O_1306,N_19903,N_19785);
xor UO_1307 (O_1307,N_19755,N_19761);
nand UO_1308 (O_1308,N_19851,N_19824);
and UO_1309 (O_1309,N_19891,N_19804);
nor UO_1310 (O_1310,N_19980,N_19803);
nor UO_1311 (O_1311,N_19809,N_19899);
xor UO_1312 (O_1312,N_19779,N_19802);
xor UO_1313 (O_1313,N_19854,N_19902);
nor UO_1314 (O_1314,N_19853,N_19781);
or UO_1315 (O_1315,N_19913,N_19860);
or UO_1316 (O_1316,N_19830,N_19755);
and UO_1317 (O_1317,N_19849,N_19941);
or UO_1318 (O_1318,N_19835,N_19782);
xnor UO_1319 (O_1319,N_19946,N_19791);
or UO_1320 (O_1320,N_19760,N_19861);
and UO_1321 (O_1321,N_19777,N_19998);
xor UO_1322 (O_1322,N_19803,N_19970);
or UO_1323 (O_1323,N_19918,N_19923);
and UO_1324 (O_1324,N_19856,N_19774);
or UO_1325 (O_1325,N_19885,N_19917);
and UO_1326 (O_1326,N_19821,N_19802);
nor UO_1327 (O_1327,N_19828,N_19926);
nand UO_1328 (O_1328,N_19986,N_19874);
nor UO_1329 (O_1329,N_19875,N_19870);
and UO_1330 (O_1330,N_19843,N_19871);
nor UO_1331 (O_1331,N_19899,N_19872);
nand UO_1332 (O_1332,N_19854,N_19845);
or UO_1333 (O_1333,N_19822,N_19980);
xor UO_1334 (O_1334,N_19842,N_19976);
and UO_1335 (O_1335,N_19944,N_19997);
or UO_1336 (O_1336,N_19870,N_19842);
nor UO_1337 (O_1337,N_19889,N_19891);
nor UO_1338 (O_1338,N_19864,N_19833);
nor UO_1339 (O_1339,N_19936,N_19914);
and UO_1340 (O_1340,N_19788,N_19968);
nor UO_1341 (O_1341,N_19932,N_19867);
nand UO_1342 (O_1342,N_19889,N_19764);
nand UO_1343 (O_1343,N_19772,N_19858);
or UO_1344 (O_1344,N_19835,N_19913);
nor UO_1345 (O_1345,N_19927,N_19959);
nand UO_1346 (O_1346,N_19927,N_19779);
or UO_1347 (O_1347,N_19922,N_19846);
nand UO_1348 (O_1348,N_19788,N_19768);
nand UO_1349 (O_1349,N_19780,N_19998);
or UO_1350 (O_1350,N_19917,N_19902);
and UO_1351 (O_1351,N_19784,N_19811);
and UO_1352 (O_1352,N_19808,N_19913);
nor UO_1353 (O_1353,N_19940,N_19932);
nor UO_1354 (O_1354,N_19981,N_19929);
nand UO_1355 (O_1355,N_19884,N_19920);
nand UO_1356 (O_1356,N_19922,N_19868);
nand UO_1357 (O_1357,N_19831,N_19833);
or UO_1358 (O_1358,N_19872,N_19925);
xor UO_1359 (O_1359,N_19876,N_19839);
and UO_1360 (O_1360,N_19781,N_19857);
or UO_1361 (O_1361,N_19947,N_19757);
nand UO_1362 (O_1362,N_19758,N_19831);
nor UO_1363 (O_1363,N_19909,N_19951);
xnor UO_1364 (O_1364,N_19880,N_19993);
and UO_1365 (O_1365,N_19760,N_19875);
nand UO_1366 (O_1366,N_19919,N_19918);
nand UO_1367 (O_1367,N_19883,N_19826);
or UO_1368 (O_1368,N_19887,N_19751);
nor UO_1369 (O_1369,N_19818,N_19870);
and UO_1370 (O_1370,N_19844,N_19805);
nor UO_1371 (O_1371,N_19768,N_19968);
xnor UO_1372 (O_1372,N_19931,N_19762);
nand UO_1373 (O_1373,N_19962,N_19866);
nand UO_1374 (O_1374,N_19804,N_19985);
nor UO_1375 (O_1375,N_19960,N_19944);
or UO_1376 (O_1376,N_19972,N_19890);
or UO_1377 (O_1377,N_19779,N_19881);
nand UO_1378 (O_1378,N_19948,N_19861);
and UO_1379 (O_1379,N_19787,N_19769);
nand UO_1380 (O_1380,N_19759,N_19818);
nor UO_1381 (O_1381,N_19792,N_19773);
or UO_1382 (O_1382,N_19909,N_19794);
and UO_1383 (O_1383,N_19879,N_19892);
and UO_1384 (O_1384,N_19942,N_19795);
nand UO_1385 (O_1385,N_19865,N_19761);
or UO_1386 (O_1386,N_19913,N_19992);
or UO_1387 (O_1387,N_19844,N_19882);
nand UO_1388 (O_1388,N_19980,N_19915);
and UO_1389 (O_1389,N_19926,N_19956);
and UO_1390 (O_1390,N_19909,N_19882);
or UO_1391 (O_1391,N_19992,N_19750);
nor UO_1392 (O_1392,N_19892,N_19937);
and UO_1393 (O_1393,N_19952,N_19990);
nor UO_1394 (O_1394,N_19959,N_19883);
nand UO_1395 (O_1395,N_19995,N_19760);
or UO_1396 (O_1396,N_19872,N_19898);
and UO_1397 (O_1397,N_19789,N_19835);
nand UO_1398 (O_1398,N_19751,N_19987);
xnor UO_1399 (O_1399,N_19879,N_19884);
nor UO_1400 (O_1400,N_19919,N_19759);
or UO_1401 (O_1401,N_19823,N_19813);
or UO_1402 (O_1402,N_19904,N_19936);
or UO_1403 (O_1403,N_19797,N_19818);
and UO_1404 (O_1404,N_19861,N_19772);
nand UO_1405 (O_1405,N_19891,N_19953);
nor UO_1406 (O_1406,N_19759,N_19809);
xnor UO_1407 (O_1407,N_19952,N_19997);
and UO_1408 (O_1408,N_19905,N_19767);
nor UO_1409 (O_1409,N_19777,N_19925);
and UO_1410 (O_1410,N_19951,N_19965);
nor UO_1411 (O_1411,N_19808,N_19791);
and UO_1412 (O_1412,N_19926,N_19984);
nand UO_1413 (O_1413,N_19858,N_19817);
nand UO_1414 (O_1414,N_19936,N_19853);
or UO_1415 (O_1415,N_19895,N_19914);
nand UO_1416 (O_1416,N_19909,N_19908);
xor UO_1417 (O_1417,N_19886,N_19777);
nor UO_1418 (O_1418,N_19893,N_19986);
xnor UO_1419 (O_1419,N_19919,N_19849);
nor UO_1420 (O_1420,N_19830,N_19827);
or UO_1421 (O_1421,N_19933,N_19905);
or UO_1422 (O_1422,N_19756,N_19887);
nor UO_1423 (O_1423,N_19832,N_19988);
and UO_1424 (O_1424,N_19843,N_19872);
or UO_1425 (O_1425,N_19964,N_19976);
xnor UO_1426 (O_1426,N_19844,N_19764);
nor UO_1427 (O_1427,N_19923,N_19908);
xnor UO_1428 (O_1428,N_19865,N_19847);
nand UO_1429 (O_1429,N_19868,N_19781);
and UO_1430 (O_1430,N_19808,N_19797);
nand UO_1431 (O_1431,N_19902,N_19916);
or UO_1432 (O_1432,N_19940,N_19907);
and UO_1433 (O_1433,N_19950,N_19835);
and UO_1434 (O_1434,N_19945,N_19770);
xnor UO_1435 (O_1435,N_19790,N_19757);
nor UO_1436 (O_1436,N_19845,N_19934);
and UO_1437 (O_1437,N_19941,N_19945);
nor UO_1438 (O_1438,N_19851,N_19868);
and UO_1439 (O_1439,N_19768,N_19878);
nand UO_1440 (O_1440,N_19817,N_19881);
or UO_1441 (O_1441,N_19770,N_19798);
nor UO_1442 (O_1442,N_19805,N_19991);
nand UO_1443 (O_1443,N_19987,N_19997);
xor UO_1444 (O_1444,N_19866,N_19781);
nor UO_1445 (O_1445,N_19817,N_19840);
or UO_1446 (O_1446,N_19877,N_19825);
and UO_1447 (O_1447,N_19950,N_19935);
and UO_1448 (O_1448,N_19801,N_19973);
nor UO_1449 (O_1449,N_19772,N_19867);
or UO_1450 (O_1450,N_19949,N_19989);
nand UO_1451 (O_1451,N_19761,N_19787);
xor UO_1452 (O_1452,N_19939,N_19895);
or UO_1453 (O_1453,N_19840,N_19810);
nand UO_1454 (O_1454,N_19805,N_19965);
and UO_1455 (O_1455,N_19971,N_19887);
and UO_1456 (O_1456,N_19867,N_19864);
nand UO_1457 (O_1457,N_19809,N_19947);
and UO_1458 (O_1458,N_19771,N_19845);
and UO_1459 (O_1459,N_19766,N_19764);
and UO_1460 (O_1460,N_19826,N_19804);
nand UO_1461 (O_1461,N_19812,N_19864);
and UO_1462 (O_1462,N_19928,N_19982);
nor UO_1463 (O_1463,N_19952,N_19866);
nand UO_1464 (O_1464,N_19958,N_19972);
or UO_1465 (O_1465,N_19925,N_19808);
xor UO_1466 (O_1466,N_19929,N_19861);
or UO_1467 (O_1467,N_19947,N_19977);
xnor UO_1468 (O_1468,N_19878,N_19750);
nand UO_1469 (O_1469,N_19803,N_19985);
nand UO_1470 (O_1470,N_19773,N_19777);
and UO_1471 (O_1471,N_19768,N_19899);
and UO_1472 (O_1472,N_19987,N_19869);
nor UO_1473 (O_1473,N_19789,N_19988);
nor UO_1474 (O_1474,N_19975,N_19976);
and UO_1475 (O_1475,N_19850,N_19776);
nor UO_1476 (O_1476,N_19876,N_19824);
xnor UO_1477 (O_1477,N_19908,N_19931);
nand UO_1478 (O_1478,N_19775,N_19783);
nand UO_1479 (O_1479,N_19983,N_19783);
nand UO_1480 (O_1480,N_19812,N_19878);
and UO_1481 (O_1481,N_19857,N_19926);
xnor UO_1482 (O_1482,N_19781,N_19842);
and UO_1483 (O_1483,N_19751,N_19871);
nor UO_1484 (O_1484,N_19940,N_19967);
and UO_1485 (O_1485,N_19859,N_19898);
nor UO_1486 (O_1486,N_19765,N_19848);
xor UO_1487 (O_1487,N_19827,N_19872);
nor UO_1488 (O_1488,N_19826,N_19900);
and UO_1489 (O_1489,N_19948,N_19789);
nand UO_1490 (O_1490,N_19821,N_19827);
and UO_1491 (O_1491,N_19953,N_19911);
and UO_1492 (O_1492,N_19922,N_19810);
and UO_1493 (O_1493,N_19760,N_19761);
nand UO_1494 (O_1494,N_19804,N_19816);
nand UO_1495 (O_1495,N_19856,N_19912);
nor UO_1496 (O_1496,N_19974,N_19949);
or UO_1497 (O_1497,N_19867,N_19820);
or UO_1498 (O_1498,N_19964,N_19981);
nand UO_1499 (O_1499,N_19841,N_19930);
nor UO_1500 (O_1500,N_19779,N_19893);
nor UO_1501 (O_1501,N_19883,N_19769);
or UO_1502 (O_1502,N_19997,N_19969);
nand UO_1503 (O_1503,N_19869,N_19895);
or UO_1504 (O_1504,N_19874,N_19837);
nor UO_1505 (O_1505,N_19819,N_19898);
nor UO_1506 (O_1506,N_19824,N_19991);
nand UO_1507 (O_1507,N_19859,N_19803);
nand UO_1508 (O_1508,N_19969,N_19866);
nand UO_1509 (O_1509,N_19915,N_19917);
or UO_1510 (O_1510,N_19902,N_19756);
or UO_1511 (O_1511,N_19810,N_19764);
or UO_1512 (O_1512,N_19910,N_19990);
nor UO_1513 (O_1513,N_19841,N_19929);
nor UO_1514 (O_1514,N_19875,N_19776);
or UO_1515 (O_1515,N_19998,N_19997);
nor UO_1516 (O_1516,N_19885,N_19833);
nand UO_1517 (O_1517,N_19897,N_19932);
nand UO_1518 (O_1518,N_19831,N_19951);
nor UO_1519 (O_1519,N_19796,N_19787);
and UO_1520 (O_1520,N_19841,N_19975);
nor UO_1521 (O_1521,N_19892,N_19995);
and UO_1522 (O_1522,N_19834,N_19985);
nand UO_1523 (O_1523,N_19944,N_19921);
or UO_1524 (O_1524,N_19779,N_19811);
nor UO_1525 (O_1525,N_19918,N_19963);
xor UO_1526 (O_1526,N_19887,N_19907);
nor UO_1527 (O_1527,N_19780,N_19879);
nand UO_1528 (O_1528,N_19957,N_19845);
nor UO_1529 (O_1529,N_19919,N_19857);
or UO_1530 (O_1530,N_19860,N_19922);
nor UO_1531 (O_1531,N_19854,N_19821);
nand UO_1532 (O_1532,N_19897,N_19812);
or UO_1533 (O_1533,N_19885,N_19974);
or UO_1534 (O_1534,N_19924,N_19981);
or UO_1535 (O_1535,N_19855,N_19769);
and UO_1536 (O_1536,N_19756,N_19869);
nor UO_1537 (O_1537,N_19884,N_19923);
xor UO_1538 (O_1538,N_19835,N_19877);
nand UO_1539 (O_1539,N_19797,N_19777);
nor UO_1540 (O_1540,N_19931,N_19935);
nor UO_1541 (O_1541,N_19945,N_19868);
or UO_1542 (O_1542,N_19875,N_19909);
or UO_1543 (O_1543,N_19969,N_19952);
nor UO_1544 (O_1544,N_19984,N_19986);
nor UO_1545 (O_1545,N_19831,N_19870);
or UO_1546 (O_1546,N_19768,N_19789);
nand UO_1547 (O_1547,N_19813,N_19810);
and UO_1548 (O_1548,N_19775,N_19908);
or UO_1549 (O_1549,N_19859,N_19971);
or UO_1550 (O_1550,N_19765,N_19981);
nor UO_1551 (O_1551,N_19767,N_19886);
nor UO_1552 (O_1552,N_19824,N_19795);
and UO_1553 (O_1553,N_19757,N_19856);
and UO_1554 (O_1554,N_19992,N_19945);
or UO_1555 (O_1555,N_19915,N_19941);
or UO_1556 (O_1556,N_19824,N_19800);
and UO_1557 (O_1557,N_19864,N_19789);
and UO_1558 (O_1558,N_19938,N_19891);
or UO_1559 (O_1559,N_19987,N_19958);
or UO_1560 (O_1560,N_19813,N_19790);
nor UO_1561 (O_1561,N_19989,N_19849);
nand UO_1562 (O_1562,N_19824,N_19895);
nand UO_1563 (O_1563,N_19850,N_19996);
nor UO_1564 (O_1564,N_19926,N_19897);
nor UO_1565 (O_1565,N_19765,N_19911);
or UO_1566 (O_1566,N_19985,N_19958);
nor UO_1567 (O_1567,N_19775,N_19817);
or UO_1568 (O_1568,N_19803,N_19996);
or UO_1569 (O_1569,N_19935,N_19866);
nand UO_1570 (O_1570,N_19793,N_19879);
nor UO_1571 (O_1571,N_19865,N_19854);
or UO_1572 (O_1572,N_19790,N_19781);
nand UO_1573 (O_1573,N_19860,N_19856);
and UO_1574 (O_1574,N_19970,N_19963);
nor UO_1575 (O_1575,N_19926,N_19915);
nor UO_1576 (O_1576,N_19751,N_19965);
and UO_1577 (O_1577,N_19916,N_19890);
and UO_1578 (O_1578,N_19772,N_19869);
nand UO_1579 (O_1579,N_19804,N_19872);
or UO_1580 (O_1580,N_19815,N_19882);
nand UO_1581 (O_1581,N_19856,N_19994);
nor UO_1582 (O_1582,N_19821,N_19893);
nand UO_1583 (O_1583,N_19776,N_19834);
nand UO_1584 (O_1584,N_19841,N_19981);
nor UO_1585 (O_1585,N_19973,N_19913);
nor UO_1586 (O_1586,N_19996,N_19814);
nand UO_1587 (O_1587,N_19884,N_19916);
and UO_1588 (O_1588,N_19823,N_19995);
nor UO_1589 (O_1589,N_19970,N_19847);
nor UO_1590 (O_1590,N_19882,N_19847);
nand UO_1591 (O_1591,N_19829,N_19875);
or UO_1592 (O_1592,N_19906,N_19915);
xnor UO_1593 (O_1593,N_19998,N_19917);
and UO_1594 (O_1594,N_19958,N_19753);
nand UO_1595 (O_1595,N_19802,N_19834);
nor UO_1596 (O_1596,N_19913,N_19896);
or UO_1597 (O_1597,N_19814,N_19787);
nand UO_1598 (O_1598,N_19858,N_19765);
nand UO_1599 (O_1599,N_19973,N_19849);
nand UO_1600 (O_1600,N_19973,N_19838);
and UO_1601 (O_1601,N_19837,N_19897);
or UO_1602 (O_1602,N_19899,N_19815);
xor UO_1603 (O_1603,N_19836,N_19926);
or UO_1604 (O_1604,N_19758,N_19760);
and UO_1605 (O_1605,N_19796,N_19888);
nand UO_1606 (O_1606,N_19888,N_19927);
nand UO_1607 (O_1607,N_19949,N_19891);
nor UO_1608 (O_1608,N_19849,N_19862);
and UO_1609 (O_1609,N_19778,N_19923);
nor UO_1610 (O_1610,N_19810,N_19879);
or UO_1611 (O_1611,N_19858,N_19976);
xor UO_1612 (O_1612,N_19884,N_19847);
and UO_1613 (O_1613,N_19939,N_19870);
nand UO_1614 (O_1614,N_19754,N_19886);
nand UO_1615 (O_1615,N_19944,N_19918);
nand UO_1616 (O_1616,N_19880,N_19945);
xnor UO_1617 (O_1617,N_19766,N_19773);
or UO_1618 (O_1618,N_19994,N_19926);
nor UO_1619 (O_1619,N_19999,N_19912);
nor UO_1620 (O_1620,N_19929,N_19984);
nand UO_1621 (O_1621,N_19805,N_19966);
nor UO_1622 (O_1622,N_19946,N_19997);
nand UO_1623 (O_1623,N_19909,N_19888);
xor UO_1624 (O_1624,N_19971,N_19998);
xor UO_1625 (O_1625,N_19928,N_19992);
or UO_1626 (O_1626,N_19944,N_19874);
nor UO_1627 (O_1627,N_19824,N_19934);
and UO_1628 (O_1628,N_19989,N_19975);
or UO_1629 (O_1629,N_19764,N_19782);
xor UO_1630 (O_1630,N_19917,N_19847);
nand UO_1631 (O_1631,N_19789,N_19934);
nor UO_1632 (O_1632,N_19863,N_19958);
xor UO_1633 (O_1633,N_19884,N_19938);
or UO_1634 (O_1634,N_19963,N_19974);
nor UO_1635 (O_1635,N_19816,N_19812);
nor UO_1636 (O_1636,N_19901,N_19934);
or UO_1637 (O_1637,N_19995,N_19912);
and UO_1638 (O_1638,N_19975,N_19768);
or UO_1639 (O_1639,N_19925,N_19848);
xnor UO_1640 (O_1640,N_19985,N_19860);
or UO_1641 (O_1641,N_19920,N_19878);
and UO_1642 (O_1642,N_19910,N_19923);
or UO_1643 (O_1643,N_19795,N_19755);
nand UO_1644 (O_1644,N_19756,N_19798);
and UO_1645 (O_1645,N_19775,N_19936);
and UO_1646 (O_1646,N_19883,N_19808);
nand UO_1647 (O_1647,N_19848,N_19939);
nor UO_1648 (O_1648,N_19972,N_19982);
xnor UO_1649 (O_1649,N_19982,N_19843);
xnor UO_1650 (O_1650,N_19860,N_19964);
nand UO_1651 (O_1651,N_19944,N_19829);
and UO_1652 (O_1652,N_19918,N_19826);
and UO_1653 (O_1653,N_19965,N_19918);
nor UO_1654 (O_1654,N_19791,N_19869);
nand UO_1655 (O_1655,N_19999,N_19841);
nor UO_1656 (O_1656,N_19964,N_19807);
xor UO_1657 (O_1657,N_19983,N_19945);
nor UO_1658 (O_1658,N_19931,N_19844);
and UO_1659 (O_1659,N_19935,N_19841);
nand UO_1660 (O_1660,N_19840,N_19985);
nand UO_1661 (O_1661,N_19976,N_19882);
or UO_1662 (O_1662,N_19880,N_19764);
and UO_1663 (O_1663,N_19994,N_19933);
or UO_1664 (O_1664,N_19884,N_19769);
and UO_1665 (O_1665,N_19770,N_19881);
or UO_1666 (O_1666,N_19935,N_19873);
nand UO_1667 (O_1667,N_19762,N_19838);
and UO_1668 (O_1668,N_19932,N_19777);
or UO_1669 (O_1669,N_19847,N_19859);
or UO_1670 (O_1670,N_19962,N_19885);
nor UO_1671 (O_1671,N_19875,N_19899);
xnor UO_1672 (O_1672,N_19944,N_19957);
or UO_1673 (O_1673,N_19864,N_19803);
nor UO_1674 (O_1674,N_19890,N_19799);
nand UO_1675 (O_1675,N_19878,N_19773);
nand UO_1676 (O_1676,N_19768,N_19758);
and UO_1677 (O_1677,N_19879,N_19911);
or UO_1678 (O_1678,N_19909,N_19843);
nand UO_1679 (O_1679,N_19804,N_19812);
xor UO_1680 (O_1680,N_19807,N_19933);
xnor UO_1681 (O_1681,N_19883,N_19938);
and UO_1682 (O_1682,N_19901,N_19984);
nand UO_1683 (O_1683,N_19796,N_19813);
nor UO_1684 (O_1684,N_19842,N_19956);
or UO_1685 (O_1685,N_19893,N_19837);
or UO_1686 (O_1686,N_19989,N_19761);
nor UO_1687 (O_1687,N_19858,N_19984);
and UO_1688 (O_1688,N_19763,N_19907);
or UO_1689 (O_1689,N_19898,N_19890);
nor UO_1690 (O_1690,N_19818,N_19995);
nor UO_1691 (O_1691,N_19828,N_19751);
and UO_1692 (O_1692,N_19920,N_19837);
or UO_1693 (O_1693,N_19875,N_19921);
nor UO_1694 (O_1694,N_19960,N_19916);
nand UO_1695 (O_1695,N_19809,N_19853);
and UO_1696 (O_1696,N_19754,N_19872);
and UO_1697 (O_1697,N_19958,N_19788);
nand UO_1698 (O_1698,N_19999,N_19759);
and UO_1699 (O_1699,N_19757,N_19814);
and UO_1700 (O_1700,N_19764,N_19982);
and UO_1701 (O_1701,N_19879,N_19754);
nand UO_1702 (O_1702,N_19814,N_19776);
nor UO_1703 (O_1703,N_19877,N_19952);
nand UO_1704 (O_1704,N_19801,N_19887);
nand UO_1705 (O_1705,N_19890,N_19965);
nand UO_1706 (O_1706,N_19954,N_19989);
or UO_1707 (O_1707,N_19781,N_19929);
or UO_1708 (O_1708,N_19815,N_19762);
and UO_1709 (O_1709,N_19771,N_19752);
or UO_1710 (O_1710,N_19980,N_19857);
or UO_1711 (O_1711,N_19816,N_19799);
and UO_1712 (O_1712,N_19930,N_19951);
or UO_1713 (O_1713,N_19906,N_19814);
nand UO_1714 (O_1714,N_19916,N_19756);
xnor UO_1715 (O_1715,N_19964,N_19814);
or UO_1716 (O_1716,N_19832,N_19836);
nand UO_1717 (O_1717,N_19771,N_19809);
and UO_1718 (O_1718,N_19793,N_19774);
nor UO_1719 (O_1719,N_19773,N_19836);
or UO_1720 (O_1720,N_19802,N_19877);
or UO_1721 (O_1721,N_19997,N_19862);
nor UO_1722 (O_1722,N_19841,N_19907);
nand UO_1723 (O_1723,N_19779,N_19760);
nor UO_1724 (O_1724,N_19823,N_19912);
nand UO_1725 (O_1725,N_19881,N_19986);
or UO_1726 (O_1726,N_19846,N_19761);
and UO_1727 (O_1727,N_19874,N_19786);
and UO_1728 (O_1728,N_19786,N_19860);
and UO_1729 (O_1729,N_19781,N_19861);
nor UO_1730 (O_1730,N_19960,N_19970);
and UO_1731 (O_1731,N_19895,N_19945);
nand UO_1732 (O_1732,N_19878,N_19988);
or UO_1733 (O_1733,N_19963,N_19941);
nand UO_1734 (O_1734,N_19766,N_19808);
nand UO_1735 (O_1735,N_19853,N_19841);
and UO_1736 (O_1736,N_19911,N_19836);
nand UO_1737 (O_1737,N_19828,N_19925);
nor UO_1738 (O_1738,N_19954,N_19836);
nand UO_1739 (O_1739,N_19952,N_19948);
or UO_1740 (O_1740,N_19910,N_19943);
or UO_1741 (O_1741,N_19782,N_19936);
xnor UO_1742 (O_1742,N_19898,N_19790);
or UO_1743 (O_1743,N_19998,N_19873);
nand UO_1744 (O_1744,N_19968,N_19875);
nand UO_1745 (O_1745,N_19923,N_19995);
and UO_1746 (O_1746,N_19967,N_19961);
nor UO_1747 (O_1747,N_19831,N_19809);
and UO_1748 (O_1748,N_19987,N_19829);
or UO_1749 (O_1749,N_19924,N_19945);
xor UO_1750 (O_1750,N_19825,N_19933);
or UO_1751 (O_1751,N_19958,N_19758);
nand UO_1752 (O_1752,N_19838,N_19813);
xnor UO_1753 (O_1753,N_19944,N_19844);
nor UO_1754 (O_1754,N_19895,N_19807);
and UO_1755 (O_1755,N_19943,N_19935);
or UO_1756 (O_1756,N_19985,N_19965);
or UO_1757 (O_1757,N_19798,N_19876);
and UO_1758 (O_1758,N_19753,N_19846);
xnor UO_1759 (O_1759,N_19853,N_19956);
and UO_1760 (O_1760,N_19857,N_19906);
nand UO_1761 (O_1761,N_19935,N_19898);
xnor UO_1762 (O_1762,N_19973,N_19834);
and UO_1763 (O_1763,N_19948,N_19931);
nor UO_1764 (O_1764,N_19992,N_19812);
xor UO_1765 (O_1765,N_19831,N_19909);
and UO_1766 (O_1766,N_19763,N_19977);
nor UO_1767 (O_1767,N_19793,N_19961);
nor UO_1768 (O_1768,N_19866,N_19783);
xor UO_1769 (O_1769,N_19971,N_19843);
and UO_1770 (O_1770,N_19968,N_19959);
nand UO_1771 (O_1771,N_19917,N_19860);
and UO_1772 (O_1772,N_19990,N_19977);
and UO_1773 (O_1773,N_19836,N_19772);
and UO_1774 (O_1774,N_19831,N_19966);
and UO_1775 (O_1775,N_19790,N_19929);
xnor UO_1776 (O_1776,N_19767,N_19907);
nand UO_1777 (O_1777,N_19867,N_19920);
and UO_1778 (O_1778,N_19753,N_19841);
and UO_1779 (O_1779,N_19787,N_19808);
nand UO_1780 (O_1780,N_19867,N_19777);
nand UO_1781 (O_1781,N_19885,N_19919);
or UO_1782 (O_1782,N_19751,N_19841);
or UO_1783 (O_1783,N_19929,N_19987);
nor UO_1784 (O_1784,N_19865,N_19750);
nand UO_1785 (O_1785,N_19899,N_19959);
nor UO_1786 (O_1786,N_19818,N_19821);
and UO_1787 (O_1787,N_19888,N_19808);
xor UO_1788 (O_1788,N_19778,N_19931);
nor UO_1789 (O_1789,N_19917,N_19813);
and UO_1790 (O_1790,N_19808,N_19772);
and UO_1791 (O_1791,N_19790,N_19764);
or UO_1792 (O_1792,N_19908,N_19994);
nand UO_1793 (O_1793,N_19835,N_19875);
nand UO_1794 (O_1794,N_19792,N_19966);
nand UO_1795 (O_1795,N_19998,N_19813);
xnor UO_1796 (O_1796,N_19950,N_19887);
nor UO_1797 (O_1797,N_19921,N_19880);
and UO_1798 (O_1798,N_19978,N_19899);
or UO_1799 (O_1799,N_19899,N_19753);
or UO_1800 (O_1800,N_19918,N_19845);
nand UO_1801 (O_1801,N_19831,N_19879);
or UO_1802 (O_1802,N_19965,N_19915);
xor UO_1803 (O_1803,N_19984,N_19837);
and UO_1804 (O_1804,N_19961,N_19751);
or UO_1805 (O_1805,N_19902,N_19798);
and UO_1806 (O_1806,N_19884,N_19781);
or UO_1807 (O_1807,N_19983,N_19841);
or UO_1808 (O_1808,N_19879,N_19962);
or UO_1809 (O_1809,N_19876,N_19956);
nand UO_1810 (O_1810,N_19961,N_19863);
and UO_1811 (O_1811,N_19916,N_19947);
or UO_1812 (O_1812,N_19953,N_19755);
or UO_1813 (O_1813,N_19910,N_19903);
or UO_1814 (O_1814,N_19822,N_19785);
or UO_1815 (O_1815,N_19871,N_19955);
and UO_1816 (O_1816,N_19838,N_19794);
or UO_1817 (O_1817,N_19869,N_19780);
and UO_1818 (O_1818,N_19771,N_19807);
or UO_1819 (O_1819,N_19838,N_19839);
nor UO_1820 (O_1820,N_19766,N_19870);
and UO_1821 (O_1821,N_19829,N_19880);
nor UO_1822 (O_1822,N_19935,N_19778);
and UO_1823 (O_1823,N_19911,N_19758);
and UO_1824 (O_1824,N_19929,N_19973);
nor UO_1825 (O_1825,N_19887,N_19833);
nand UO_1826 (O_1826,N_19954,N_19769);
and UO_1827 (O_1827,N_19965,N_19912);
or UO_1828 (O_1828,N_19867,N_19987);
and UO_1829 (O_1829,N_19965,N_19959);
nand UO_1830 (O_1830,N_19786,N_19973);
xnor UO_1831 (O_1831,N_19761,N_19868);
nor UO_1832 (O_1832,N_19893,N_19941);
nor UO_1833 (O_1833,N_19853,N_19843);
nor UO_1834 (O_1834,N_19968,N_19786);
or UO_1835 (O_1835,N_19754,N_19758);
nand UO_1836 (O_1836,N_19763,N_19759);
nor UO_1837 (O_1837,N_19972,N_19835);
nand UO_1838 (O_1838,N_19853,N_19882);
or UO_1839 (O_1839,N_19909,N_19768);
and UO_1840 (O_1840,N_19982,N_19803);
or UO_1841 (O_1841,N_19939,N_19919);
nand UO_1842 (O_1842,N_19826,N_19811);
nor UO_1843 (O_1843,N_19946,N_19877);
nand UO_1844 (O_1844,N_19753,N_19795);
nand UO_1845 (O_1845,N_19867,N_19937);
nor UO_1846 (O_1846,N_19983,N_19937);
nand UO_1847 (O_1847,N_19959,N_19888);
and UO_1848 (O_1848,N_19987,N_19788);
nor UO_1849 (O_1849,N_19866,N_19902);
and UO_1850 (O_1850,N_19807,N_19838);
nor UO_1851 (O_1851,N_19926,N_19964);
and UO_1852 (O_1852,N_19982,N_19920);
or UO_1853 (O_1853,N_19926,N_19882);
or UO_1854 (O_1854,N_19943,N_19929);
or UO_1855 (O_1855,N_19997,N_19758);
and UO_1856 (O_1856,N_19777,N_19820);
nand UO_1857 (O_1857,N_19813,N_19895);
nor UO_1858 (O_1858,N_19843,N_19959);
xor UO_1859 (O_1859,N_19905,N_19915);
nor UO_1860 (O_1860,N_19761,N_19750);
xnor UO_1861 (O_1861,N_19997,N_19921);
or UO_1862 (O_1862,N_19785,N_19792);
and UO_1863 (O_1863,N_19798,N_19837);
xnor UO_1864 (O_1864,N_19960,N_19863);
xnor UO_1865 (O_1865,N_19983,N_19795);
nor UO_1866 (O_1866,N_19791,N_19753);
and UO_1867 (O_1867,N_19940,N_19927);
nor UO_1868 (O_1868,N_19867,N_19902);
nand UO_1869 (O_1869,N_19968,N_19916);
nor UO_1870 (O_1870,N_19970,N_19806);
xor UO_1871 (O_1871,N_19864,N_19797);
and UO_1872 (O_1872,N_19761,N_19946);
and UO_1873 (O_1873,N_19827,N_19838);
and UO_1874 (O_1874,N_19842,N_19894);
and UO_1875 (O_1875,N_19965,N_19973);
and UO_1876 (O_1876,N_19955,N_19784);
or UO_1877 (O_1877,N_19953,N_19929);
or UO_1878 (O_1878,N_19894,N_19938);
nand UO_1879 (O_1879,N_19951,N_19906);
nor UO_1880 (O_1880,N_19863,N_19769);
xor UO_1881 (O_1881,N_19942,N_19922);
nand UO_1882 (O_1882,N_19973,N_19815);
or UO_1883 (O_1883,N_19857,N_19978);
xor UO_1884 (O_1884,N_19828,N_19966);
or UO_1885 (O_1885,N_19998,N_19874);
xnor UO_1886 (O_1886,N_19785,N_19975);
xnor UO_1887 (O_1887,N_19804,N_19873);
or UO_1888 (O_1888,N_19832,N_19898);
or UO_1889 (O_1889,N_19769,N_19842);
nor UO_1890 (O_1890,N_19817,N_19989);
nand UO_1891 (O_1891,N_19813,N_19883);
nor UO_1892 (O_1892,N_19800,N_19883);
nand UO_1893 (O_1893,N_19966,N_19785);
xnor UO_1894 (O_1894,N_19916,N_19817);
xnor UO_1895 (O_1895,N_19869,N_19911);
nand UO_1896 (O_1896,N_19872,N_19852);
or UO_1897 (O_1897,N_19781,N_19872);
and UO_1898 (O_1898,N_19940,N_19947);
nor UO_1899 (O_1899,N_19993,N_19869);
nand UO_1900 (O_1900,N_19757,N_19995);
nor UO_1901 (O_1901,N_19893,N_19866);
nand UO_1902 (O_1902,N_19861,N_19835);
nor UO_1903 (O_1903,N_19988,N_19926);
or UO_1904 (O_1904,N_19767,N_19831);
xnor UO_1905 (O_1905,N_19889,N_19893);
nor UO_1906 (O_1906,N_19952,N_19876);
nor UO_1907 (O_1907,N_19815,N_19911);
nand UO_1908 (O_1908,N_19831,N_19896);
or UO_1909 (O_1909,N_19780,N_19863);
nor UO_1910 (O_1910,N_19877,N_19915);
xnor UO_1911 (O_1911,N_19789,N_19796);
or UO_1912 (O_1912,N_19889,N_19792);
nor UO_1913 (O_1913,N_19985,N_19875);
and UO_1914 (O_1914,N_19927,N_19863);
nand UO_1915 (O_1915,N_19753,N_19860);
nand UO_1916 (O_1916,N_19952,N_19777);
and UO_1917 (O_1917,N_19895,N_19905);
nand UO_1918 (O_1918,N_19878,N_19970);
nand UO_1919 (O_1919,N_19962,N_19788);
or UO_1920 (O_1920,N_19916,N_19796);
xor UO_1921 (O_1921,N_19837,N_19884);
xnor UO_1922 (O_1922,N_19885,N_19877);
nand UO_1923 (O_1923,N_19919,N_19758);
nand UO_1924 (O_1924,N_19928,N_19753);
and UO_1925 (O_1925,N_19763,N_19954);
and UO_1926 (O_1926,N_19794,N_19887);
and UO_1927 (O_1927,N_19929,N_19821);
and UO_1928 (O_1928,N_19859,N_19879);
nor UO_1929 (O_1929,N_19756,N_19994);
nor UO_1930 (O_1930,N_19766,N_19847);
or UO_1931 (O_1931,N_19899,N_19954);
and UO_1932 (O_1932,N_19844,N_19845);
nor UO_1933 (O_1933,N_19907,N_19809);
or UO_1934 (O_1934,N_19904,N_19828);
xor UO_1935 (O_1935,N_19802,N_19797);
and UO_1936 (O_1936,N_19781,N_19786);
nand UO_1937 (O_1937,N_19868,N_19801);
nand UO_1938 (O_1938,N_19822,N_19781);
nand UO_1939 (O_1939,N_19839,N_19954);
and UO_1940 (O_1940,N_19944,N_19992);
nand UO_1941 (O_1941,N_19936,N_19807);
nor UO_1942 (O_1942,N_19970,N_19904);
or UO_1943 (O_1943,N_19970,N_19867);
xnor UO_1944 (O_1944,N_19921,N_19825);
and UO_1945 (O_1945,N_19976,N_19979);
or UO_1946 (O_1946,N_19867,N_19763);
xnor UO_1947 (O_1947,N_19826,N_19867);
and UO_1948 (O_1948,N_19829,N_19897);
or UO_1949 (O_1949,N_19852,N_19921);
and UO_1950 (O_1950,N_19823,N_19974);
nor UO_1951 (O_1951,N_19815,N_19781);
or UO_1952 (O_1952,N_19988,N_19853);
or UO_1953 (O_1953,N_19916,N_19878);
xnor UO_1954 (O_1954,N_19898,N_19846);
or UO_1955 (O_1955,N_19858,N_19871);
or UO_1956 (O_1956,N_19939,N_19867);
xor UO_1957 (O_1957,N_19919,N_19827);
nand UO_1958 (O_1958,N_19956,N_19963);
or UO_1959 (O_1959,N_19819,N_19802);
nand UO_1960 (O_1960,N_19957,N_19751);
and UO_1961 (O_1961,N_19819,N_19818);
and UO_1962 (O_1962,N_19830,N_19799);
nor UO_1963 (O_1963,N_19852,N_19804);
and UO_1964 (O_1964,N_19882,N_19935);
nor UO_1965 (O_1965,N_19965,N_19761);
nand UO_1966 (O_1966,N_19895,N_19901);
or UO_1967 (O_1967,N_19958,N_19825);
or UO_1968 (O_1968,N_19985,N_19887);
or UO_1969 (O_1969,N_19806,N_19835);
xor UO_1970 (O_1970,N_19832,N_19947);
nor UO_1971 (O_1971,N_19856,N_19761);
nor UO_1972 (O_1972,N_19916,N_19858);
and UO_1973 (O_1973,N_19912,N_19986);
nand UO_1974 (O_1974,N_19868,N_19981);
nor UO_1975 (O_1975,N_19785,N_19855);
nand UO_1976 (O_1976,N_19935,N_19770);
and UO_1977 (O_1977,N_19919,N_19787);
or UO_1978 (O_1978,N_19914,N_19872);
or UO_1979 (O_1979,N_19975,N_19752);
and UO_1980 (O_1980,N_19914,N_19833);
nand UO_1981 (O_1981,N_19850,N_19958);
nand UO_1982 (O_1982,N_19793,N_19977);
or UO_1983 (O_1983,N_19919,N_19778);
or UO_1984 (O_1984,N_19875,N_19993);
nor UO_1985 (O_1985,N_19813,N_19914);
or UO_1986 (O_1986,N_19787,N_19892);
or UO_1987 (O_1987,N_19869,N_19821);
and UO_1988 (O_1988,N_19752,N_19808);
and UO_1989 (O_1989,N_19838,N_19894);
and UO_1990 (O_1990,N_19750,N_19816);
and UO_1991 (O_1991,N_19972,N_19813);
and UO_1992 (O_1992,N_19751,N_19914);
or UO_1993 (O_1993,N_19754,N_19884);
and UO_1994 (O_1994,N_19767,N_19931);
nor UO_1995 (O_1995,N_19836,N_19891);
nand UO_1996 (O_1996,N_19877,N_19798);
nand UO_1997 (O_1997,N_19778,N_19994);
nor UO_1998 (O_1998,N_19786,N_19899);
or UO_1999 (O_1999,N_19756,N_19790);
nor UO_2000 (O_2000,N_19828,N_19900);
nand UO_2001 (O_2001,N_19758,N_19788);
or UO_2002 (O_2002,N_19914,N_19888);
xnor UO_2003 (O_2003,N_19792,N_19821);
nor UO_2004 (O_2004,N_19955,N_19872);
nand UO_2005 (O_2005,N_19965,N_19768);
nand UO_2006 (O_2006,N_19868,N_19757);
or UO_2007 (O_2007,N_19800,N_19777);
or UO_2008 (O_2008,N_19750,N_19906);
nand UO_2009 (O_2009,N_19960,N_19889);
nand UO_2010 (O_2010,N_19964,N_19985);
and UO_2011 (O_2011,N_19928,N_19950);
or UO_2012 (O_2012,N_19878,N_19919);
or UO_2013 (O_2013,N_19859,N_19942);
nand UO_2014 (O_2014,N_19930,N_19967);
nor UO_2015 (O_2015,N_19997,N_19970);
and UO_2016 (O_2016,N_19870,N_19803);
or UO_2017 (O_2017,N_19801,N_19804);
nor UO_2018 (O_2018,N_19913,N_19869);
nand UO_2019 (O_2019,N_19961,N_19762);
and UO_2020 (O_2020,N_19787,N_19887);
nor UO_2021 (O_2021,N_19753,N_19985);
nor UO_2022 (O_2022,N_19959,N_19809);
nand UO_2023 (O_2023,N_19819,N_19933);
and UO_2024 (O_2024,N_19998,N_19928);
nor UO_2025 (O_2025,N_19823,N_19842);
nand UO_2026 (O_2026,N_19935,N_19856);
nand UO_2027 (O_2027,N_19976,N_19974);
nand UO_2028 (O_2028,N_19864,N_19785);
nand UO_2029 (O_2029,N_19901,N_19803);
nor UO_2030 (O_2030,N_19797,N_19791);
nand UO_2031 (O_2031,N_19758,N_19988);
nor UO_2032 (O_2032,N_19838,N_19816);
and UO_2033 (O_2033,N_19978,N_19798);
xor UO_2034 (O_2034,N_19908,N_19813);
nand UO_2035 (O_2035,N_19761,N_19973);
and UO_2036 (O_2036,N_19982,N_19859);
nand UO_2037 (O_2037,N_19882,N_19796);
or UO_2038 (O_2038,N_19988,N_19856);
and UO_2039 (O_2039,N_19944,N_19864);
nand UO_2040 (O_2040,N_19859,N_19780);
or UO_2041 (O_2041,N_19836,N_19961);
or UO_2042 (O_2042,N_19761,N_19992);
nor UO_2043 (O_2043,N_19956,N_19836);
and UO_2044 (O_2044,N_19796,N_19860);
nor UO_2045 (O_2045,N_19860,N_19986);
nor UO_2046 (O_2046,N_19934,N_19823);
or UO_2047 (O_2047,N_19893,N_19885);
xnor UO_2048 (O_2048,N_19922,N_19876);
or UO_2049 (O_2049,N_19992,N_19924);
and UO_2050 (O_2050,N_19818,N_19928);
nor UO_2051 (O_2051,N_19830,N_19894);
or UO_2052 (O_2052,N_19798,N_19954);
and UO_2053 (O_2053,N_19955,N_19940);
and UO_2054 (O_2054,N_19787,N_19785);
nand UO_2055 (O_2055,N_19873,N_19964);
xnor UO_2056 (O_2056,N_19993,N_19802);
and UO_2057 (O_2057,N_19873,N_19906);
nor UO_2058 (O_2058,N_19753,N_19969);
nand UO_2059 (O_2059,N_19918,N_19981);
or UO_2060 (O_2060,N_19917,N_19890);
nor UO_2061 (O_2061,N_19887,N_19982);
and UO_2062 (O_2062,N_19972,N_19989);
nor UO_2063 (O_2063,N_19825,N_19866);
or UO_2064 (O_2064,N_19903,N_19832);
or UO_2065 (O_2065,N_19939,N_19810);
xnor UO_2066 (O_2066,N_19969,N_19844);
nand UO_2067 (O_2067,N_19803,N_19806);
nand UO_2068 (O_2068,N_19940,N_19858);
or UO_2069 (O_2069,N_19974,N_19932);
nor UO_2070 (O_2070,N_19911,N_19889);
nand UO_2071 (O_2071,N_19954,N_19981);
nand UO_2072 (O_2072,N_19814,N_19862);
and UO_2073 (O_2073,N_19905,N_19823);
nor UO_2074 (O_2074,N_19832,N_19904);
nor UO_2075 (O_2075,N_19881,N_19907);
nand UO_2076 (O_2076,N_19791,N_19894);
nor UO_2077 (O_2077,N_19758,N_19752);
or UO_2078 (O_2078,N_19955,N_19915);
nand UO_2079 (O_2079,N_19933,N_19870);
and UO_2080 (O_2080,N_19791,N_19921);
xor UO_2081 (O_2081,N_19908,N_19934);
nor UO_2082 (O_2082,N_19908,N_19788);
nand UO_2083 (O_2083,N_19826,N_19775);
or UO_2084 (O_2084,N_19923,N_19795);
or UO_2085 (O_2085,N_19915,N_19920);
and UO_2086 (O_2086,N_19876,N_19924);
nand UO_2087 (O_2087,N_19970,N_19896);
nand UO_2088 (O_2088,N_19942,N_19761);
nor UO_2089 (O_2089,N_19945,N_19987);
and UO_2090 (O_2090,N_19952,N_19808);
nor UO_2091 (O_2091,N_19954,N_19884);
and UO_2092 (O_2092,N_19812,N_19904);
or UO_2093 (O_2093,N_19865,N_19807);
and UO_2094 (O_2094,N_19889,N_19886);
or UO_2095 (O_2095,N_19979,N_19852);
nand UO_2096 (O_2096,N_19992,N_19786);
xor UO_2097 (O_2097,N_19845,N_19789);
and UO_2098 (O_2098,N_19930,N_19856);
nor UO_2099 (O_2099,N_19750,N_19869);
and UO_2100 (O_2100,N_19919,N_19786);
nor UO_2101 (O_2101,N_19965,N_19820);
nor UO_2102 (O_2102,N_19867,N_19885);
nand UO_2103 (O_2103,N_19872,N_19988);
and UO_2104 (O_2104,N_19943,N_19953);
xnor UO_2105 (O_2105,N_19939,N_19851);
nand UO_2106 (O_2106,N_19989,N_19948);
nand UO_2107 (O_2107,N_19793,N_19889);
nor UO_2108 (O_2108,N_19993,N_19760);
nor UO_2109 (O_2109,N_19941,N_19959);
and UO_2110 (O_2110,N_19867,N_19802);
xor UO_2111 (O_2111,N_19903,N_19992);
or UO_2112 (O_2112,N_19782,N_19856);
and UO_2113 (O_2113,N_19903,N_19905);
and UO_2114 (O_2114,N_19779,N_19813);
and UO_2115 (O_2115,N_19987,N_19838);
or UO_2116 (O_2116,N_19773,N_19898);
and UO_2117 (O_2117,N_19785,N_19932);
nand UO_2118 (O_2118,N_19900,N_19830);
nor UO_2119 (O_2119,N_19822,N_19927);
and UO_2120 (O_2120,N_19798,N_19974);
and UO_2121 (O_2121,N_19803,N_19958);
nand UO_2122 (O_2122,N_19869,N_19834);
nor UO_2123 (O_2123,N_19760,N_19782);
or UO_2124 (O_2124,N_19988,N_19947);
and UO_2125 (O_2125,N_19896,N_19774);
or UO_2126 (O_2126,N_19757,N_19756);
xor UO_2127 (O_2127,N_19885,N_19834);
and UO_2128 (O_2128,N_19937,N_19769);
nor UO_2129 (O_2129,N_19908,N_19871);
and UO_2130 (O_2130,N_19896,N_19784);
or UO_2131 (O_2131,N_19838,N_19773);
or UO_2132 (O_2132,N_19795,N_19985);
or UO_2133 (O_2133,N_19968,N_19837);
and UO_2134 (O_2134,N_19997,N_19753);
and UO_2135 (O_2135,N_19964,N_19918);
nand UO_2136 (O_2136,N_19847,N_19787);
nor UO_2137 (O_2137,N_19934,N_19933);
and UO_2138 (O_2138,N_19909,N_19889);
xor UO_2139 (O_2139,N_19812,N_19983);
nor UO_2140 (O_2140,N_19908,N_19956);
nor UO_2141 (O_2141,N_19845,N_19924);
nand UO_2142 (O_2142,N_19805,N_19827);
or UO_2143 (O_2143,N_19937,N_19804);
or UO_2144 (O_2144,N_19816,N_19911);
nand UO_2145 (O_2145,N_19778,N_19966);
and UO_2146 (O_2146,N_19905,N_19780);
nand UO_2147 (O_2147,N_19888,N_19975);
or UO_2148 (O_2148,N_19833,N_19892);
or UO_2149 (O_2149,N_19950,N_19805);
and UO_2150 (O_2150,N_19929,N_19906);
nor UO_2151 (O_2151,N_19986,N_19795);
nor UO_2152 (O_2152,N_19963,N_19754);
or UO_2153 (O_2153,N_19875,N_19922);
nand UO_2154 (O_2154,N_19878,N_19941);
nand UO_2155 (O_2155,N_19978,N_19954);
and UO_2156 (O_2156,N_19929,N_19968);
nor UO_2157 (O_2157,N_19812,N_19762);
or UO_2158 (O_2158,N_19828,N_19917);
nor UO_2159 (O_2159,N_19761,N_19832);
nand UO_2160 (O_2160,N_19906,N_19998);
or UO_2161 (O_2161,N_19929,N_19899);
nand UO_2162 (O_2162,N_19987,N_19845);
or UO_2163 (O_2163,N_19925,N_19774);
nor UO_2164 (O_2164,N_19864,N_19779);
or UO_2165 (O_2165,N_19782,N_19891);
xnor UO_2166 (O_2166,N_19886,N_19774);
and UO_2167 (O_2167,N_19767,N_19836);
nor UO_2168 (O_2168,N_19958,N_19993);
or UO_2169 (O_2169,N_19824,N_19963);
and UO_2170 (O_2170,N_19911,N_19922);
and UO_2171 (O_2171,N_19930,N_19804);
and UO_2172 (O_2172,N_19779,N_19892);
or UO_2173 (O_2173,N_19974,N_19782);
xor UO_2174 (O_2174,N_19966,N_19751);
nor UO_2175 (O_2175,N_19778,N_19752);
nor UO_2176 (O_2176,N_19850,N_19885);
and UO_2177 (O_2177,N_19912,N_19956);
and UO_2178 (O_2178,N_19971,N_19826);
nand UO_2179 (O_2179,N_19943,N_19845);
nor UO_2180 (O_2180,N_19829,N_19949);
nor UO_2181 (O_2181,N_19927,N_19991);
or UO_2182 (O_2182,N_19897,N_19791);
nor UO_2183 (O_2183,N_19830,N_19855);
and UO_2184 (O_2184,N_19793,N_19888);
or UO_2185 (O_2185,N_19856,N_19934);
nand UO_2186 (O_2186,N_19999,N_19762);
and UO_2187 (O_2187,N_19920,N_19750);
and UO_2188 (O_2188,N_19994,N_19986);
xnor UO_2189 (O_2189,N_19914,N_19944);
and UO_2190 (O_2190,N_19750,N_19795);
xor UO_2191 (O_2191,N_19828,N_19982);
or UO_2192 (O_2192,N_19759,N_19755);
or UO_2193 (O_2193,N_19807,N_19811);
xnor UO_2194 (O_2194,N_19853,N_19943);
and UO_2195 (O_2195,N_19982,N_19949);
nor UO_2196 (O_2196,N_19899,N_19964);
nor UO_2197 (O_2197,N_19924,N_19882);
or UO_2198 (O_2198,N_19884,N_19870);
nor UO_2199 (O_2199,N_19927,N_19847);
nor UO_2200 (O_2200,N_19843,N_19939);
nand UO_2201 (O_2201,N_19976,N_19861);
and UO_2202 (O_2202,N_19982,N_19857);
xnor UO_2203 (O_2203,N_19971,N_19795);
and UO_2204 (O_2204,N_19915,N_19901);
nor UO_2205 (O_2205,N_19883,N_19779);
nor UO_2206 (O_2206,N_19930,N_19845);
and UO_2207 (O_2207,N_19927,N_19787);
nor UO_2208 (O_2208,N_19920,N_19967);
nand UO_2209 (O_2209,N_19918,N_19807);
nand UO_2210 (O_2210,N_19852,N_19888);
or UO_2211 (O_2211,N_19928,N_19794);
or UO_2212 (O_2212,N_19801,N_19857);
and UO_2213 (O_2213,N_19990,N_19911);
xor UO_2214 (O_2214,N_19998,N_19919);
or UO_2215 (O_2215,N_19939,N_19981);
and UO_2216 (O_2216,N_19994,N_19839);
xnor UO_2217 (O_2217,N_19873,N_19818);
and UO_2218 (O_2218,N_19933,N_19947);
and UO_2219 (O_2219,N_19983,N_19765);
nor UO_2220 (O_2220,N_19999,N_19855);
or UO_2221 (O_2221,N_19841,N_19879);
or UO_2222 (O_2222,N_19953,N_19827);
nor UO_2223 (O_2223,N_19889,N_19828);
or UO_2224 (O_2224,N_19972,N_19992);
xor UO_2225 (O_2225,N_19944,N_19793);
nor UO_2226 (O_2226,N_19949,N_19915);
or UO_2227 (O_2227,N_19760,N_19919);
xnor UO_2228 (O_2228,N_19758,N_19834);
and UO_2229 (O_2229,N_19865,N_19960);
nand UO_2230 (O_2230,N_19977,N_19988);
and UO_2231 (O_2231,N_19916,N_19928);
xnor UO_2232 (O_2232,N_19944,N_19801);
nor UO_2233 (O_2233,N_19802,N_19926);
nor UO_2234 (O_2234,N_19975,N_19850);
and UO_2235 (O_2235,N_19980,N_19849);
nor UO_2236 (O_2236,N_19937,N_19787);
nor UO_2237 (O_2237,N_19953,N_19887);
xor UO_2238 (O_2238,N_19794,N_19882);
nand UO_2239 (O_2239,N_19903,N_19952);
or UO_2240 (O_2240,N_19811,N_19952);
and UO_2241 (O_2241,N_19773,N_19783);
or UO_2242 (O_2242,N_19911,N_19952);
nand UO_2243 (O_2243,N_19775,N_19782);
nand UO_2244 (O_2244,N_19840,N_19967);
or UO_2245 (O_2245,N_19854,N_19925);
nand UO_2246 (O_2246,N_19934,N_19804);
nand UO_2247 (O_2247,N_19808,N_19965);
and UO_2248 (O_2248,N_19815,N_19834);
or UO_2249 (O_2249,N_19858,N_19937);
and UO_2250 (O_2250,N_19970,N_19930);
and UO_2251 (O_2251,N_19878,N_19951);
or UO_2252 (O_2252,N_19872,N_19788);
or UO_2253 (O_2253,N_19808,N_19829);
and UO_2254 (O_2254,N_19799,N_19868);
nand UO_2255 (O_2255,N_19942,N_19806);
nand UO_2256 (O_2256,N_19968,N_19907);
or UO_2257 (O_2257,N_19844,N_19835);
xor UO_2258 (O_2258,N_19867,N_19785);
or UO_2259 (O_2259,N_19960,N_19811);
nor UO_2260 (O_2260,N_19942,N_19853);
nor UO_2261 (O_2261,N_19929,N_19856);
nand UO_2262 (O_2262,N_19859,N_19850);
xor UO_2263 (O_2263,N_19903,N_19870);
and UO_2264 (O_2264,N_19773,N_19893);
or UO_2265 (O_2265,N_19803,N_19751);
or UO_2266 (O_2266,N_19836,N_19898);
or UO_2267 (O_2267,N_19891,N_19862);
or UO_2268 (O_2268,N_19876,N_19906);
and UO_2269 (O_2269,N_19905,N_19864);
and UO_2270 (O_2270,N_19989,N_19873);
nand UO_2271 (O_2271,N_19907,N_19771);
or UO_2272 (O_2272,N_19840,N_19842);
or UO_2273 (O_2273,N_19974,N_19846);
nor UO_2274 (O_2274,N_19757,N_19863);
nor UO_2275 (O_2275,N_19772,N_19755);
xor UO_2276 (O_2276,N_19811,N_19970);
or UO_2277 (O_2277,N_19947,N_19807);
and UO_2278 (O_2278,N_19953,N_19815);
xor UO_2279 (O_2279,N_19764,N_19915);
nand UO_2280 (O_2280,N_19945,N_19832);
or UO_2281 (O_2281,N_19908,N_19933);
nand UO_2282 (O_2282,N_19902,N_19818);
or UO_2283 (O_2283,N_19872,N_19906);
or UO_2284 (O_2284,N_19757,N_19894);
and UO_2285 (O_2285,N_19920,N_19835);
nand UO_2286 (O_2286,N_19845,N_19864);
nand UO_2287 (O_2287,N_19928,N_19834);
nor UO_2288 (O_2288,N_19868,N_19838);
xnor UO_2289 (O_2289,N_19796,N_19959);
or UO_2290 (O_2290,N_19945,N_19753);
nand UO_2291 (O_2291,N_19937,N_19934);
nor UO_2292 (O_2292,N_19842,N_19791);
or UO_2293 (O_2293,N_19828,N_19955);
nand UO_2294 (O_2294,N_19956,N_19938);
nor UO_2295 (O_2295,N_19903,N_19830);
and UO_2296 (O_2296,N_19876,N_19859);
nor UO_2297 (O_2297,N_19830,N_19824);
or UO_2298 (O_2298,N_19780,N_19873);
nor UO_2299 (O_2299,N_19916,N_19887);
xor UO_2300 (O_2300,N_19824,N_19782);
nand UO_2301 (O_2301,N_19990,N_19767);
nand UO_2302 (O_2302,N_19811,N_19817);
or UO_2303 (O_2303,N_19943,N_19940);
xor UO_2304 (O_2304,N_19974,N_19813);
nand UO_2305 (O_2305,N_19987,N_19912);
nand UO_2306 (O_2306,N_19808,N_19816);
and UO_2307 (O_2307,N_19990,N_19894);
or UO_2308 (O_2308,N_19833,N_19868);
xor UO_2309 (O_2309,N_19757,N_19916);
and UO_2310 (O_2310,N_19757,N_19932);
nor UO_2311 (O_2311,N_19948,N_19990);
or UO_2312 (O_2312,N_19992,N_19986);
nor UO_2313 (O_2313,N_19892,N_19846);
or UO_2314 (O_2314,N_19780,N_19837);
nand UO_2315 (O_2315,N_19892,N_19925);
and UO_2316 (O_2316,N_19751,N_19880);
xor UO_2317 (O_2317,N_19821,N_19997);
or UO_2318 (O_2318,N_19997,N_19858);
and UO_2319 (O_2319,N_19806,N_19875);
nor UO_2320 (O_2320,N_19871,N_19950);
nor UO_2321 (O_2321,N_19885,N_19971);
or UO_2322 (O_2322,N_19903,N_19873);
nand UO_2323 (O_2323,N_19928,N_19964);
and UO_2324 (O_2324,N_19804,N_19904);
nand UO_2325 (O_2325,N_19940,N_19843);
and UO_2326 (O_2326,N_19881,N_19859);
nand UO_2327 (O_2327,N_19983,N_19832);
xor UO_2328 (O_2328,N_19753,N_19989);
or UO_2329 (O_2329,N_19982,N_19893);
nor UO_2330 (O_2330,N_19947,N_19804);
or UO_2331 (O_2331,N_19847,N_19901);
xnor UO_2332 (O_2332,N_19766,N_19975);
nand UO_2333 (O_2333,N_19850,N_19811);
nor UO_2334 (O_2334,N_19827,N_19995);
nor UO_2335 (O_2335,N_19913,N_19898);
or UO_2336 (O_2336,N_19840,N_19981);
or UO_2337 (O_2337,N_19820,N_19993);
and UO_2338 (O_2338,N_19901,N_19991);
or UO_2339 (O_2339,N_19850,N_19981);
nand UO_2340 (O_2340,N_19989,N_19776);
and UO_2341 (O_2341,N_19985,N_19919);
nor UO_2342 (O_2342,N_19822,N_19882);
nor UO_2343 (O_2343,N_19768,N_19923);
and UO_2344 (O_2344,N_19965,N_19976);
and UO_2345 (O_2345,N_19783,N_19759);
or UO_2346 (O_2346,N_19906,N_19937);
or UO_2347 (O_2347,N_19788,N_19834);
nand UO_2348 (O_2348,N_19981,N_19988);
nor UO_2349 (O_2349,N_19928,N_19978);
nor UO_2350 (O_2350,N_19870,N_19783);
nand UO_2351 (O_2351,N_19925,N_19868);
nor UO_2352 (O_2352,N_19892,N_19837);
nand UO_2353 (O_2353,N_19910,N_19858);
nor UO_2354 (O_2354,N_19942,N_19998);
nand UO_2355 (O_2355,N_19915,N_19855);
nand UO_2356 (O_2356,N_19905,N_19875);
and UO_2357 (O_2357,N_19942,N_19829);
xor UO_2358 (O_2358,N_19903,N_19757);
or UO_2359 (O_2359,N_19852,N_19978);
nand UO_2360 (O_2360,N_19971,N_19911);
and UO_2361 (O_2361,N_19857,N_19981);
nor UO_2362 (O_2362,N_19764,N_19847);
and UO_2363 (O_2363,N_19754,N_19804);
and UO_2364 (O_2364,N_19923,N_19807);
or UO_2365 (O_2365,N_19934,N_19834);
and UO_2366 (O_2366,N_19963,N_19992);
nor UO_2367 (O_2367,N_19754,N_19987);
or UO_2368 (O_2368,N_19975,N_19999);
or UO_2369 (O_2369,N_19847,N_19861);
or UO_2370 (O_2370,N_19973,N_19908);
and UO_2371 (O_2371,N_19954,N_19759);
or UO_2372 (O_2372,N_19956,N_19843);
nor UO_2373 (O_2373,N_19975,N_19890);
and UO_2374 (O_2374,N_19904,N_19855);
nand UO_2375 (O_2375,N_19810,N_19883);
nand UO_2376 (O_2376,N_19883,N_19836);
and UO_2377 (O_2377,N_19909,N_19906);
nor UO_2378 (O_2378,N_19930,N_19918);
nand UO_2379 (O_2379,N_19865,N_19996);
or UO_2380 (O_2380,N_19832,N_19973);
and UO_2381 (O_2381,N_19924,N_19994);
nand UO_2382 (O_2382,N_19829,N_19751);
nand UO_2383 (O_2383,N_19856,N_19895);
nor UO_2384 (O_2384,N_19770,N_19836);
and UO_2385 (O_2385,N_19847,N_19813);
nor UO_2386 (O_2386,N_19832,N_19878);
and UO_2387 (O_2387,N_19914,N_19923);
nand UO_2388 (O_2388,N_19928,N_19995);
nor UO_2389 (O_2389,N_19945,N_19985);
nand UO_2390 (O_2390,N_19777,N_19884);
or UO_2391 (O_2391,N_19782,N_19881);
and UO_2392 (O_2392,N_19969,N_19872);
nor UO_2393 (O_2393,N_19908,N_19899);
and UO_2394 (O_2394,N_19769,N_19941);
and UO_2395 (O_2395,N_19776,N_19799);
or UO_2396 (O_2396,N_19947,N_19971);
nand UO_2397 (O_2397,N_19978,N_19962);
nor UO_2398 (O_2398,N_19816,N_19939);
nand UO_2399 (O_2399,N_19896,N_19877);
nand UO_2400 (O_2400,N_19833,N_19963);
and UO_2401 (O_2401,N_19825,N_19948);
nor UO_2402 (O_2402,N_19995,N_19869);
nand UO_2403 (O_2403,N_19783,N_19861);
xnor UO_2404 (O_2404,N_19948,N_19782);
nor UO_2405 (O_2405,N_19984,N_19942);
or UO_2406 (O_2406,N_19903,N_19937);
or UO_2407 (O_2407,N_19948,N_19982);
nand UO_2408 (O_2408,N_19908,N_19951);
nand UO_2409 (O_2409,N_19966,N_19988);
or UO_2410 (O_2410,N_19861,N_19883);
and UO_2411 (O_2411,N_19915,N_19765);
and UO_2412 (O_2412,N_19903,N_19948);
nor UO_2413 (O_2413,N_19883,N_19897);
or UO_2414 (O_2414,N_19948,N_19752);
nor UO_2415 (O_2415,N_19938,N_19838);
xnor UO_2416 (O_2416,N_19989,N_19884);
and UO_2417 (O_2417,N_19974,N_19860);
and UO_2418 (O_2418,N_19813,N_19798);
and UO_2419 (O_2419,N_19755,N_19957);
and UO_2420 (O_2420,N_19853,N_19800);
nand UO_2421 (O_2421,N_19963,N_19907);
nor UO_2422 (O_2422,N_19893,N_19877);
and UO_2423 (O_2423,N_19884,N_19958);
or UO_2424 (O_2424,N_19898,N_19902);
nor UO_2425 (O_2425,N_19970,N_19860);
nand UO_2426 (O_2426,N_19785,N_19807);
nand UO_2427 (O_2427,N_19989,N_19866);
nand UO_2428 (O_2428,N_19974,N_19975);
nand UO_2429 (O_2429,N_19795,N_19955);
nor UO_2430 (O_2430,N_19865,N_19948);
nor UO_2431 (O_2431,N_19938,N_19858);
nor UO_2432 (O_2432,N_19991,N_19812);
or UO_2433 (O_2433,N_19988,N_19938);
nand UO_2434 (O_2434,N_19790,N_19880);
or UO_2435 (O_2435,N_19760,N_19900);
and UO_2436 (O_2436,N_19947,N_19750);
and UO_2437 (O_2437,N_19977,N_19856);
xor UO_2438 (O_2438,N_19937,N_19750);
xnor UO_2439 (O_2439,N_19914,N_19873);
nand UO_2440 (O_2440,N_19786,N_19906);
nor UO_2441 (O_2441,N_19923,N_19776);
nand UO_2442 (O_2442,N_19895,N_19887);
or UO_2443 (O_2443,N_19994,N_19991);
nand UO_2444 (O_2444,N_19911,N_19851);
and UO_2445 (O_2445,N_19989,N_19856);
xnor UO_2446 (O_2446,N_19889,N_19939);
and UO_2447 (O_2447,N_19888,N_19883);
and UO_2448 (O_2448,N_19935,N_19766);
and UO_2449 (O_2449,N_19953,N_19874);
xor UO_2450 (O_2450,N_19778,N_19879);
and UO_2451 (O_2451,N_19982,N_19880);
xnor UO_2452 (O_2452,N_19783,N_19825);
nand UO_2453 (O_2453,N_19967,N_19769);
nand UO_2454 (O_2454,N_19818,N_19811);
nor UO_2455 (O_2455,N_19770,N_19982);
and UO_2456 (O_2456,N_19823,N_19814);
and UO_2457 (O_2457,N_19776,N_19960);
nand UO_2458 (O_2458,N_19890,N_19853);
nand UO_2459 (O_2459,N_19928,N_19881);
nor UO_2460 (O_2460,N_19842,N_19865);
and UO_2461 (O_2461,N_19950,N_19803);
or UO_2462 (O_2462,N_19925,N_19905);
nor UO_2463 (O_2463,N_19839,N_19846);
nor UO_2464 (O_2464,N_19946,N_19813);
or UO_2465 (O_2465,N_19958,N_19963);
or UO_2466 (O_2466,N_19981,N_19905);
and UO_2467 (O_2467,N_19960,N_19968);
nor UO_2468 (O_2468,N_19875,N_19808);
and UO_2469 (O_2469,N_19871,N_19801);
and UO_2470 (O_2470,N_19792,N_19806);
and UO_2471 (O_2471,N_19803,N_19955);
nand UO_2472 (O_2472,N_19957,N_19863);
nor UO_2473 (O_2473,N_19900,N_19833);
or UO_2474 (O_2474,N_19963,N_19898);
and UO_2475 (O_2475,N_19875,N_19957);
nand UO_2476 (O_2476,N_19960,N_19763);
nor UO_2477 (O_2477,N_19836,N_19933);
and UO_2478 (O_2478,N_19998,N_19773);
nand UO_2479 (O_2479,N_19797,N_19925);
and UO_2480 (O_2480,N_19984,N_19894);
nand UO_2481 (O_2481,N_19764,N_19967);
nand UO_2482 (O_2482,N_19801,N_19830);
nor UO_2483 (O_2483,N_19952,N_19910);
or UO_2484 (O_2484,N_19811,N_19867);
or UO_2485 (O_2485,N_19841,N_19844);
nor UO_2486 (O_2486,N_19899,N_19784);
or UO_2487 (O_2487,N_19927,N_19849);
xnor UO_2488 (O_2488,N_19851,N_19915);
and UO_2489 (O_2489,N_19905,N_19779);
nand UO_2490 (O_2490,N_19917,N_19851);
nand UO_2491 (O_2491,N_19931,N_19843);
or UO_2492 (O_2492,N_19995,N_19796);
and UO_2493 (O_2493,N_19976,N_19940);
or UO_2494 (O_2494,N_19863,N_19825);
nand UO_2495 (O_2495,N_19871,N_19756);
nand UO_2496 (O_2496,N_19827,N_19898);
nand UO_2497 (O_2497,N_19754,N_19948);
and UO_2498 (O_2498,N_19755,N_19948);
or UO_2499 (O_2499,N_19976,N_19840);
endmodule