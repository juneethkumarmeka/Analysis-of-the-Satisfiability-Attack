module basic_2500_25000_3000_50_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1203,In_2335);
nor U1 (N_1,In_503,In_2105);
nand U2 (N_2,In_1715,In_2266);
nand U3 (N_3,In_819,In_471);
or U4 (N_4,In_583,In_1359);
and U5 (N_5,In_2233,In_345);
xor U6 (N_6,In_2040,In_522);
and U7 (N_7,In_263,In_2141);
or U8 (N_8,In_1869,In_2048);
and U9 (N_9,In_2384,In_123);
nor U10 (N_10,In_2244,In_2329);
nand U11 (N_11,In_298,In_2164);
nor U12 (N_12,In_2173,In_1010);
and U13 (N_13,In_184,In_1561);
or U14 (N_14,In_1563,In_2341);
xnor U15 (N_15,In_910,In_1683);
or U16 (N_16,In_1427,In_1199);
nand U17 (N_17,In_1914,In_2369);
xnor U18 (N_18,In_549,In_647);
or U19 (N_19,In_1933,In_2063);
nand U20 (N_20,In_576,In_1170);
nand U21 (N_21,In_1982,In_1850);
or U22 (N_22,In_2235,In_1278);
nand U23 (N_23,In_1056,In_1755);
or U24 (N_24,In_39,In_1688);
and U25 (N_25,In_1326,In_1773);
nor U26 (N_26,In_2316,In_1034);
and U27 (N_27,In_967,In_698);
nand U28 (N_28,In_565,In_954);
nand U29 (N_29,In_2184,In_988);
nor U30 (N_30,In_2143,In_831);
nand U31 (N_31,In_1100,In_1525);
or U32 (N_32,In_2339,In_461);
nor U33 (N_33,In_1699,In_1239);
or U34 (N_34,In_2411,In_305);
and U35 (N_35,In_224,In_450);
and U36 (N_36,In_1319,In_2267);
nor U37 (N_37,In_310,In_198);
nor U38 (N_38,In_1618,In_1904);
nand U39 (N_39,In_1084,In_837);
and U40 (N_40,In_719,In_2431);
nor U41 (N_41,In_741,In_1925);
or U42 (N_42,In_750,In_1210);
and U43 (N_43,In_2125,In_1114);
nor U44 (N_44,In_1268,In_1208);
nand U45 (N_45,In_1674,In_2206);
nand U46 (N_46,In_361,In_2292);
xnor U47 (N_47,In_1031,In_1002);
nand U48 (N_48,In_1197,In_1856);
and U49 (N_49,In_2491,In_408);
nand U50 (N_50,In_1201,In_248);
nand U51 (N_51,In_435,In_1454);
or U52 (N_52,In_1596,In_1644);
and U53 (N_53,In_1472,In_1445);
and U54 (N_54,In_1779,In_149);
and U55 (N_55,In_508,In_753);
and U56 (N_56,In_1901,In_2163);
nand U57 (N_57,In_1703,In_330);
nor U58 (N_58,In_2452,In_178);
nor U59 (N_59,In_1250,In_564);
nand U60 (N_60,In_365,In_2211);
nor U61 (N_61,In_1587,In_1556);
or U62 (N_62,In_1189,In_1775);
or U63 (N_63,In_1527,In_771);
or U64 (N_64,In_2152,In_1336);
xor U65 (N_65,In_824,In_2458);
or U66 (N_66,In_1424,In_2247);
or U67 (N_67,In_518,In_1416);
nor U68 (N_68,In_1630,In_2301);
and U69 (N_69,In_1829,In_1501);
nor U70 (N_70,In_1870,In_2187);
and U71 (N_71,In_2189,In_434);
or U72 (N_72,In_462,In_2137);
nor U73 (N_73,In_2407,In_2272);
nor U74 (N_74,In_1656,In_47);
nand U75 (N_75,In_431,In_845);
and U76 (N_76,In_88,In_92);
and U77 (N_77,In_321,In_869);
xor U78 (N_78,In_513,In_2304);
xor U79 (N_79,In_390,In_1626);
nand U80 (N_80,In_2002,In_1781);
and U81 (N_81,In_418,In_2228);
and U82 (N_82,In_1449,In_113);
or U83 (N_83,In_2471,In_1269);
or U84 (N_84,In_707,In_1037);
nor U85 (N_85,In_151,In_1685);
nand U86 (N_86,In_812,In_12);
xor U87 (N_87,In_1185,In_1207);
xnor U88 (N_88,In_889,In_1743);
or U89 (N_89,In_798,In_162);
nor U90 (N_90,In_282,In_2053);
and U91 (N_91,In_1428,In_356);
nor U92 (N_92,In_0,In_43);
xor U93 (N_93,In_1811,In_2019);
or U94 (N_94,In_1568,In_923);
xor U95 (N_95,In_2317,In_1158);
and U96 (N_96,In_2380,In_2386);
nand U97 (N_97,In_2483,In_748);
nand U98 (N_98,In_813,In_1079);
or U99 (N_99,In_2481,In_1886);
and U100 (N_100,In_903,In_732);
nand U101 (N_101,In_504,In_966);
and U102 (N_102,In_402,In_957);
or U103 (N_103,In_28,In_1083);
nor U104 (N_104,In_2179,In_1431);
or U105 (N_105,In_677,In_554);
or U106 (N_106,In_1019,In_419);
or U107 (N_107,In_601,In_497);
nor U108 (N_108,In_2410,In_1680);
nand U109 (N_109,In_1602,In_255);
nand U110 (N_110,In_2284,In_2416);
and U111 (N_111,In_2007,In_2006);
or U112 (N_112,In_1337,In_219);
or U113 (N_113,In_706,In_2364);
and U114 (N_114,In_687,In_117);
xor U115 (N_115,In_2277,In_484);
nand U116 (N_116,In_1749,In_2234);
nor U117 (N_117,In_476,In_104);
nand U118 (N_118,In_441,In_1394);
and U119 (N_119,In_1752,In_2077);
nand U120 (N_120,In_317,In_512);
nand U121 (N_121,In_458,In_2475);
and U122 (N_122,In_448,In_1857);
and U123 (N_123,In_2276,In_1795);
and U124 (N_124,In_169,In_2379);
nor U125 (N_125,In_1074,In_2221);
and U126 (N_126,In_1629,In_912);
nand U127 (N_127,In_621,In_2375);
nand U128 (N_128,In_1796,In_1619);
nor U129 (N_129,In_929,In_1774);
nor U130 (N_130,In_1710,In_1138);
or U131 (N_131,In_1273,In_909);
nand U132 (N_132,In_668,In_2037);
nor U133 (N_133,In_1279,In_2367);
or U134 (N_134,In_1382,In_166);
xnor U135 (N_135,In_2132,In_1997);
and U136 (N_136,In_977,In_2102);
or U137 (N_137,In_1046,In_1579);
nor U138 (N_138,In_992,In_1924);
or U139 (N_139,In_7,In_1800);
xnor U140 (N_140,In_896,In_1999);
nor U141 (N_141,In_1689,In_314);
or U142 (N_142,In_126,In_1132);
nor U143 (N_143,In_1754,In_56);
nor U144 (N_144,In_1168,In_1162);
nand U145 (N_145,In_492,In_1885);
xor U146 (N_146,In_120,In_1011);
nor U147 (N_147,In_1669,In_849);
nand U148 (N_148,In_1860,In_15);
nor U149 (N_149,In_1875,In_713);
or U150 (N_150,In_1953,In_2114);
or U151 (N_151,In_1569,In_412);
and U152 (N_152,In_1729,In_1330);
or U153 (N_153,In_1632,In_1276);
nand U154 (N_154,In_980,In_1589);
or U155 (N_155,In_284,In_2360);
xor U156 (N_156,In_2171,In_981);
nor U157 (N_157,In_651,In_1045);
nor U158 (N_158,In_2089,In_1890);
nand U159 (N_159,In_1888,In_1701);
nor U160 (N_160,In_1607,In_2172);
nand U161 (N_161,In_1971,In_1955);
nor U162 (N_162,In_1038,In_1893);
or U163 (N_163,In_1522,In_873);
nor U164 (N_164,In_2197,In_1897);
or U165 (N_165,In_1183,In_1735);
nor U166 (N_166,In_78,In_2287);
nand U167 (N_167,In_2154,In_972);
nand U168 (N_168,In_860,In_1673);
nand U169 (N_169,In_469,In_1747);
nand U170 (N_170,In_618,In_1530);
or U171 (N_171,In_355,In_1111);
or U172 (N_172,In_944,In_573);
and U173 (N_173,In_1960,In_1731);
nand U174 (N_174,In_1603,In_35);
or U175 (N_175,In_1164,In_1967);
and U176 (N_176,In_1966,In_993);
and U177 (N_177,In_1545,In_1756);
nor U178 (N_178,In_363,In_2196);
and U179 (N_179,In_1842,In_342);
and U180 (N_180,In_1894,In_2413);
nand U181 (N_181,In_1861,In_1557);
or U182 (N_182,In_787,In_1266);
nand U183 (N_183,In_1837,In_574);
nor U184 (N_184,In_2273,In_751);
nor U185 (N_185,In_1863,In_2011);
and U186 (N_186,In_905,In_1469);
and U187 (N_187,In_1661,In_1512);
and U188 (N_188,In_1020,In_67);
or U189 (N_189,In_792,In_1347);
nor U190 (N_190,In_1913,In_353);
nand U191 (N_191,In_1766,In_1161);
nand U192 (N_192,In_1108,In_2406);
or U193 (N_193,In_1050,In_2209);
nor U194 (N_194,In_274,In_1306);
nor U195 (N_195,In_1093,In_636);
and U196 (N_196,In_1400,In_24);
nand U197 (N_197,In_2162,In_313);
or U198 (N_198,In_2299,In_1565);
or U199 (N_199,In_2049,In_464);
or U200 (N_200,In_505,In_1116);
or U201 (N_201,In_2240,In_577);
nand U202 (N_202,In_1312,In_2027);
and U203 (N_203,In_163,In_782);
nand U204 (N_204,In_2357,In_1814);
or U205 (N_205,In_1601,In_2440);
or U206 (N_206,In_1687,In_146);
nand U207 (N_207,In_828,In_267);
and U208 (N_208,In_2430,In_2437);
and U209 (N_209,In_351,In_2351);
nor U210 (N_210,In_742,In_1434);
nor U211 (N_211,In_1004,In_1932);
nand U212 (N_212,In_1912,In_319);
or U213 (N_213,In_159,In_602);
and U214 (N_214,In_2004,In_273);
nor U215 (N_215,In_1395,In_1128);
and U216 (N_216,In_1243,In_1282);
nand U217 (N_217,In_83,In_95);
or U218 (N_218,In_2024,In_2098);
xnor U219 (N_219,In_140,In_1152);
nand U220 (N_220,In_1694,In_2438);
nand U221 (N_221,In_662,In_2282);
nor U222 (N_222,In_1973,In_223);
and U223 (N_223,In_2237,In_332);
and U224 (N_224,In_375,In_2322);
nand U225 (N_225,In_2227,In_1588);
nor U226 (N_226,In_347,In_1213);
or U227 (N_227,In_2409,In_2252);
nor U228 (N_228,In_1738,In_2298);
and U229 (N_229,In_1836,In_2484);
nor U230 (N_230,In_1057,In_1113);
and U231 (N_231,In_615,In_478);
or U232 (N_232,In_403,In_1780);
nor U233 (N_233,In_1003,In_1221);
or U234 (N_234,In_116,In_724);
xor U235 (N_235,In_2307,In_1098);
nand U236 (N_236,In_745,In_623);
nand U237 (N_237,In_139,In_585);
nor U238 (N_238,In_1249,In_2337);
and U239 (N_239,In_1172,In_1817);
and U240 (N_240,In_611,In_1753);
or U241 (N_241,In_2257,In_2338);
nor U242 (N_242,In_951,In_2314);
nor U243 (N_243,In_1041,In_1044);
nor U244 (N_244,In_1553,In_1290);
or U245 (N_245,In_109,In_407);
or U246 (N_246,In_609,In_1786);
nor U247 (N_247,In_718,In_1981);
or U248 (N_248,In_1574,In_2133);
or U249 (N_249,In_1797,In_1702);
nor U250 (N_250,In_1493,In_1389);
or U251 (N_251,In_1181,In_733);
nand U252 (N_252,In_1898,In_171);
nor U253 (N_253,In_2156,In_1272);
nand U254 (N_254,In_2183,In_1102);
or U255 (N_255,In_68,In_941);
xnor U256 (N_256,In_272,In_1280);
nand U257 (N_257,In_244,In_709);
or U258 (N_258,In_2450,In_1346);
xnor U259 (N_259,In_2248,In_422);
xor U260 (N_260,In_1304,In_661);
and U261 (N_261,In_1135,In_1819);
or U262 (N_262,In_1302,In_1824);
and U263 (N_263,In_1583,In_1483);
and U264 (N_264,In_1918,In_1670);
and U265 (N_265,In_2123,In_1495);
xnor U266 (N_266,In_2265,In_1645);
nor U267 (N_267,In_892,In_50);
and U268 (N_268,In_2117,In_1867);
nand U269 (N_269,In_791,In_1463);
nor U270 (N_270,In_1926,In_848);
nor U271 (N_271,In_1295,In_1976);
nor U272 (N_272,In_697,In_2015);
nand U273 (N_273,In_1,In_1834);
nor U274 (N_274,In_1492,In_1147);
and U275 (N_275,In_1484,In_776);
nand U276 (N_276,In_772,In_640);
and U277 (N_277,In_1062,In_1146);
nand U278 (N_278,In_1235,In_920);
and U279 (N_279,In_1672,In_1115);
and U280 (N_280,In_2111,In_1818);
and U281 (N_281,In_1532,In_1684);
nand U282 (N_282,In_550,In_1307);
or U283 (N_283,In_1040,In_1145);
and U284 (N_284,In_1435,In_757);
nand U285 (N_285,In_1071,In_535);
nand U286 (N_286,In_1992,In_2195);
nor U287 (N_287,In_998,In_1223);
nand U288 (N_288,In_1091,In_1001);
xor U289 (N_289,In_105,In_301);
nand U290 (N_290,In_372,In_1090);
xor U291 (N_291,In_2054,In_1939);
nor U292 (N_292,In_31,In_1027);
and U293 (N_293,In_1746,In_2081);
and U294 (N_294,In_2095,In_194);
nor U295 (N_295,In_1957,In_4);
or U296 (N_296,In_52,In_1081);
and U297 (N_297,In_1174,In_593);
and U298 (N_298,In_256,In_213);
nor U299 (N_299,In_532,In_770);
and U300 (N_300,In_1948,In_727);
nor U301 (N_301,In_2368,In_265);
and U302 (N_302,In_1977,In_173);
and U303 (N_303,In_886,In_234);
nand U304 (N_304,In_1772,In_2175);
xor U305 (N_305,In_879,In_1092);
and U306 (N_306,In_610,In_843);
nor U307 (N_307,In_451,In_1163);
and U308 (N_308,In_2488,In_1622);
nor U309 (N_309,In_1810,In_1544);
and U310 (N_310,In_102,In_414);
and U311 (N_311,In_2336,In_1720);
and U312 (N_312,In_1776,In_2436);
and U313 (N_313,In_2250,In_2318);
nand U314 (N_314,In_1486,In_71);
nor U315 (N_315,In_1119,In_1157);
and U316 (N_316,In_1457,In_2071);
or U317 (N_317,In_1101,In_1335);
nor U318 (N_318,In_1399,In_562);
and U319 (N_319,In_996,In_594);
nand U320 (N_320,In_898,In_934);
or U321 (N_321,In_2327,In_135);
or U322 (N_322,In_190,In_2457);
nor U323 (N_323,In_1740,In_2108);
nand U324 (N_324,In_2347,In_2426);
nand U325 (N_325,In_1641,In_1832);
nand U326 (N_326,In_1442,In_2487);
xor U327 (N_327,In_820,In_1505);
nor U328 (N_328,In_2356,In_1984);
and U329 (N_329,In_93,In_536);
and U330 (N_330,In_287,In_1790);
and U331 (N_331,In_271,In_936);
nor U332 (N_332,In_2468,In_2434);
nor U333 (N_333,In_165,In_1049);
and U334 (N_334,In_1432,In_290);
nand U335 (N_335,In_1464,In_2366);
nand U336 (N_336,In_876,In_439);
and U337 (N_337,In_334,In_888);
xnor U338 (N_338,In_32,In_1838);
and U339 (N_339,In_2151,In_1120);
nor U340 (N_340,In_2005,In_208);
or U341 (N_341,In_1891,In_2365);
nor U342 (N_342,In_654,In_211);
nand U343 (N_343,In_2062,In_333);
nor U344 (N_344,In_100,In_145);
nand U345 (N_345,In_1851,In_1535);
or U346 (N_346,In_2190,In_138);
xnor U347 (N_347,In_1730,In_1691);
nand U348 (N_348,In_150,In_1853);
nor U349 (N_349,In_2289,In_421);
or U350 (N_350,In_1309,In_129);
and U351 (N_351,In_1708,In_2078);
and U352 (N_352,In_875,In_2290);
xor U353 (N_353,In_856,In_2178);
and U354 (N_354,In_1066,In_1864);
nand U355 (N_355,In_2448,In_1274);
and U356 (N_356,In_1865,In_229);
or U357 (N_357,In_1620,In_1663);
and U358 (N_358,In_1778,In_130);
xnor U359 (N_359,In_2136,In_261);
nor U360 (N_360,In_632,In_584);
xor U361 (N_361,In_708,In_952);
and U362 (N_362,In_182,In_1363);
or U363 (N_363,In_2447,In_1537);
or U364 (N_364,In_595,In_1193);
xor U365 (N_365,In_231,In_1154);
nand U366 (N_366,In_19,In_1647);
nor U367 (N_367,In_767,In_1156);
nor U368 (N_368,In_468,In_1112);
or U369 (N_369,In_588,In_2119);
nand U370 (N_370,In_1671,In_1627);
nand U371 (N_371,In_2417,In_1825);
xor U372 (N_372,In_1440,In_2215);
or U373 (N_373,In_1323,In_1012);
nor U374 (N_374,In_38,In_1721);
and U375 (N_375,In_1131,In_49);
or U376 (N_376,In_1375,In_1256);
nor U377 (N_377,In_380,In_1546);
nor U378 (N_378,In_57,In_2100);
and U379 (N_379,In_1209,In_1808);
or U380 (N_380,In_1757,In_1234);
nor U381 (N_381,In_481,In_1809);
and U382 (N_382,In_477,In_1067);
or U383 (N_383,In_2180,In_2218);
nand U384 (N_384,In_2067,In_37);
nand U385 (N_385,In_1725,In_1889);
and U386 (N_386,In_884,In_1030);
and U387 (N_387,In_1451,In_23);
nand U388 (N_388,In_420,In_1471);
nor U389 (N_389,In_153,In_1718);
or U390 (N_390,In_22,In_877);
nand U391 (N_391,In_761,In_2432);
nand U392 (N_392,In_855,In_2383);
and U393 (N_393,In_656,In_1650);
and U394 (N_394,In_1169,In_1065);
or U395 (N_395,In_2388,In_2074);
and U396 (N_396,In_1419,In_1257);
and U397 (N_397,In_950,In_1621);
and U398 (N_398,In_1129,In_2405);
and U399 (N_399,In_2499,In_486);
nand U400 (N_400,In_1059,In_1515);
and U401 (N_401,In_1233,In_215);
nand U402 (N_402,In_2349,In_2275);
nor U403 (N_403,In_930,In_1241);
and U404 (N_404,In_2047,In_620);
nand U405 (N_405,In_1297,In_1386);
and U406 (N_406,In_36,In_1402);
or U407 (N_407,In_976,In_2070);
or U408 (N_408,In_2490,In_669);
nor U409 (N_409,In_409,In_887);
or U410 (N_410,In_1777,In_1783);
xnor U411 (N_411,In_586,In_587);
nor U412 (N_412,In_1998,In_1491);
and U413 (N_413,In_125,In_1764);
and U414 (N_414,In_704,In_1008);
and U415 (N_415,In_2008,In_962);
nand U416 (N_416,In_299,In_259);
nand U417 (N_417,In_459,In_1247);
nor U418 (N_418,In_2096,In_596);
nand U419 (N_419,In_2076,In_2231);
or U420 (N_420,In_1315,In_1087);
or U421 (N_421,In_986,In_1379);
xnor U422 (N_422,In_1868,In_1225);
nand U423 (N_423,In_2449,In_1543);
or U424 (N_424,In_2200,In_685);
or U425 (N_425,In_1230,In_2168);
nor U426 (N_426,In_449,In_191);
nand U427 (N_427,In_247,In_2442);
or U428 (N_428,In_2285,In_17);
nor U429 (N_429,In_1334,In_1762);
xnor U430 (N_430,In_281,In_1060);
or U431 (N_431,In_2497,In_2274);
nand U432 (N_432,In_559,In_2253);
and U433 (N_433,In_510,In_2198);
nor U434 (N_434,In_1640,In_1013);
nand U435 (N_435,In_2455,In_245);
nand U436 (N_436,In_1662,In_2372);
nor U437 (N_437,In_1763,In_1639);
and U438 (N_438,In_1513,In_991);
nand U439 (N_439,In_1608,In_21);
nand U440 (N_440,In_913,In_2262);
and U441 (N_441,In_2112,In_1069);
and U442 (N_442,In_346,In_2391);
nand U443 (N_443,In_1651,In_1965);
nor U444 (N_444,In_1370,In_1910);
nor U445 (N_445,In_107,In_1734);
and U446 (N_446,In_254,In_1453);
xnor U447 (N_447,In_371,In_2121);
nor U448 (N_448,In_1942,In_160);
nand U449 (N_449,In_1785,In_735);
nand U450 (N_450,In_1813,In_279);
xnor U451 (N_451,In_1109,In_2315);
nand U452 (N_452,In_1009,In_1541);
nor U453 (N_453,In_1341,In_2118);
xor U454 (N_454,In_1499,In_756);
and U455 (N_455,In_1840,In_1270);
and U456 (N_456,In_1294,In_2045);
or U457 (N_457,In_514,In_2026);
or U458 (N_458,In_1974,In_8);
nand U459 (N_459,In_715,In_714);
or U460 (N_460,In_10,In_2381);
and U461 (N_461,In_628,In_2138);
and U462 (N_462,In_1919,In_711);
nor U463 (N_463,In_2238,In_61);
or U464 (N_464,In_774,In_1693);
nand U465 (N_465,In_379,In_567);
and U466 (N_466,In_2361,In_1231);
or U467 (N_467,In_627,In_1633);
nand U468 (N_468,In_2226,In_94);
nor U469 (N_469,In_2496,In_1745);
nor U470 (N_470,In_2344,In_2099);
nand U471 (N_471,In_1528,In_1139);
or U472 (N_472,In_1481,In_2495);
nand U473 (N_473,In_309,In_1920);
nand U474 (N_474,In_1951,In_1305);
nor U475 (N_475,In_847,In_664);
nand U476 (N_476,In_2330,In_2398);
or U477 (N_477,In_404,In_30);
nand U478 (N_478,In_1166,In_1187);
and U479 (N_479,In_1993,In_79);
nand U480 (N_480,In_1823,In_63);
xnor U481 (N_481,In_341,In_168);
nor U482 (N_482,In_343,In_366);
xor U483 (N_483,In_963,In_1907);
nor U484 (N_484,In_1787,In_2092);
xor U485 (N_485,In_200,In_1063);
nand U486 (N_486,In_2176,In_960);
nand U487 (N_487,In_827,In_251);
nand U488 (N_488,In_1724,In_1042);
xor U489 (N_489,In_2232,In_2306);
nor U490 (N_490,In_1996,In_793);
and U491 (N_491,In_556,In_2308);
and U492 (N_492,In_1255,In_721);
nand U493 (N_493,In_561,In_1356);
and U494 (N_494,In_466,In_385);
xnor U495 (N_495,In_457,In_1381);
nand U496 (N_496,In_260,In_2427);
nor U497 (N_497,In_376,In_1252);
xnor U498 (N_498,In_2177,In_2286);
or U499 (N_499,In_633,In_1956);
and U500 (N_500,In_425,In_1401);
nand U501 (N_501,In_599,In_1529);
and U502 (N_502,N_144,In_1127);
nor U503 (N_503,In_1521,N_459);
and U504 (N_504,In_1459,N_7);
or U505 (N_505,In_1643,In_175);
nand U506 (N_506,N_325,In_2331);
or U507 (N_507,In_1106,In_838);
nand U508 (N_508,In_1732,In_597);
nor U509 (N_509,N_184,In_320);
nor U510 (N_510,In_1118,In_1947);
nor U511 (N_511,N_105,In_1903);
or U512 (N_512,N_36,In_253);
nor U513 (N_513,In_2142,N_341);
nor U514 (N_514,In_97,N_78);
nand U515 (N_515,In_746,In_1103);
or U516 (N_516,In_187,N_131);
xnor U517 (N_517,In_1324,In_1333);
nor U518 (N_518,In_1498,In_2161);
nor U519 (N_519,In_316,In_349);
nor U520 (N_520,In_1659,In_27);
nand U521 (N_521,In_1068,In_1872);
nand U522 (N_522,N_77,In_54);
xnor U523 (N_523,N_197,In_740);
nor U524 (N_524,In_60,In_2480);
and U525 (N_525,N_98,In_540);
nand U526 (N_526,In_2088,In_91);
or U527 (N_527,In_1600,In_1934);
or U528 (N_528,N_442,In_1686);
xor U529 (N_529,In_127,In_1478);
nor U530 (N_530,N_236,N_237);
or U531 (N_531,In_2193,N_170);
nand U532 (N_532,In_1329,In_904);
or U533 (N_533,In_1711,In_897);
or U534 (N_534,N_25,In_2342);
and U535 (N_535,In_465,In_2073);
nand U536 (N_536,In_1859,In_895);
xnor U537 (N_537,In_2101,N_432);
or U538 (N_538,N_60,In_1364);
nand U539 (N_539,N_122,In_1141);
nand U540 (N_540,In_2464,In_1595);
and U541 (N_541,In_581,N_259);
nor U542 (N_542,In_1547,In_275);
or U543 (N_543,N_20,In_940);
and U544 (N_544,In_297,In_98);
nand U545 (N_545,N_199,N_319);
and U546 (N_546,In_46,In_2323);
nand U547 (N_547,In_648,In_1523);
nand U548 (N_548,In_2363,In_695);
nand U549 (N_549,In_455,In_2346);
xor U550 (N_550,In_164,In_850);
and U551 (N_551,In_1342,N_95);
or U552 (N_552,In_89,In_671);
nor U553 (N_553,In_526,In_1460);
nor U554 (N_554,In_193,N_106);
or U555 (N_555,In_1476,In_866);
nand U556 (N_556,In_1831,In_1877);
or U557 (N_557,In_1503,In_1204);
nor U558 (N_558,In_802,N_446);
or U559 (N_559,In_2397,In_511);
nor U560 (N_560,In_1806,In_1423);
or U561 (N_561,In_1945,In_397);
nand U562 (N_562,In_328,In_1820);
and U563 (N_563,In_202,In_572);
and U564 (N_564,N_393,In_1550);
nor U565 (N_565,In_426,In_2036);
xor U566 (N_566,In_1862,In_1648);
nor U567 (N_567,In_189,In_1979);
and U568 (N_568,In_1107,In_1655);
and U569 (N_569,In_1612,In_300);
nor U570 (N_570,N_457,In_1150);
or U571 (N_571,In_20,In_1418);
xnor U572 (N_572,N_149,In_207);
nor U573 (N_573,In_395,In_306);
and U574 (N_574,In_738,In_818);
and U575 (N_575,In_916,In_1938);
xor U576 (N_576,In_357,In_2044);
nand U577 (N_577,In_1909,In_786);
nor U578 (N_578,N_128,N_348);
nor U579 (N_579,In_1318,In_2041);
and U580 (N_580,In_730,N_491);
and U581 (N_581,In_2472,In_147);
xnor U582 (N_582,N_90,In_1344);
nor U583 (N_583,In_558,N_167);
nor U584 (N_584,In_2167,N_83);
or U585 (N_585,In_1206,In_1950);
or U586 (N_586,In_1802,In_515);
or U587 (N_587,In_1229,N_431);
xnor U588 (N_588,In_1990,N_246);
xnor U589 (N_589,In_218,In_1317);
or U590 (N_590,In_766,In_1064);
or U591 (N_591,In_399,In_1219);
or U592 (N_592,In_1261,In_2009);
nor U593 (N_593,In_293,N_69);
nand U594 (N_594,N_439,In_509);
nor U595 (N_595,N_357,In_578);
nor U596 (N_596,N_322,N_157);
and U597 (N_597,In_1217,In_788);
nor U598 (N_598,In_686,N_18);
nand U599 (N_599,In_2454,In_1258);
and U600 (N_600,N_80,In_1299);
or U601 (N_601,In_6,In_1182);
and U602 (N_602,N_435,In_373);
or U603 (N_603,N_412,In_552);
and U604 (N_604,In_1858,In_1482);
or U605 (N_605,N_407,In_1717);
xor U606 (N_606,In_1931,In_2283);
or U607 (N_607,N_494,In_984);
nor U608 (N_608,In_1200,In_672);
nand U609 (N_609,In_1228,In_666);
xnor U610 (N_610,In_1338,N_355);
nor U611 (N_611,In_1360,In_1039);
or U612 (N_612,N_151,In_2354);
and U613 (N_613,N_293,N_472);
nand U614 (N_614,In_295,In_358);
and U615 (N_615,In_655,N_159);
nor U616 (N_616,N_231,In_479);
nand U617 (N_617,In_1123,In_496);
and U618 (N_618,In_1794,In_1741);
nand U619 (N_619,N_99,In_527);
or U620 (N_620,In_1409,In_438);
and U621 (N_621,In_1771,In_283);
nand U622 (N_622,N_294,In_429);
or U623 (N_623,In_2203,In_1705);
xor U624 (N_624,In_1542,In_382);
or U625 (N_625,N_460,In_1211);
or U626 (N_626,In_307,In_2429);
nand U627 (N_627,N_338,In_652);
and U628 (N_628,N_245,In_1357);
nand U629 (N_629,In_2207,In_1043);
xor U630 (N_630,In_26,In_874);
xnor U631 (N_631,N_162,In_947);
and U632 (N_632,In_192,In_720);
nor U633 (N_633,In_2473,N_356);
nor U634 (N_634,In_1534,N_3);
and U635 (N_635,In_1425,In_2446);
nand U636 (N_636,In_606,In_1277);
xor U637 (N_637,In_1377,In_688);
nor U638 (N_638,N_468,In_285);
and U639 (N_639,N_448,In_1308);
or U640 (N_640,In_1303,In_1559);
and U641 (N_641,In_1636,N_209);
nor U642 (N_642,In_681,N_256);
and U643 (N_643,In_520,N_428);
xnor U644 (N_644,In_1846,In_2281);
or U645 (N_645,N_306,In_2489);
or U646 (N_646,In_70,N_311);
or U647 (N_647,In_2103,In_548);
nand U648 (N_648,N_299,In_268);
or U649 (N_649,N_146,In_338);
nand U650 (N_650,In_62,N_372);
nor U651 (N_651,In_1876,In_2353);
nand U652 (N_652,N_206,In_45);
or U653 (N_653,In_2120,In_2166);
nor U654 (N_654,In_2186,In_2439);
and U655 (N_655,In_1052,In_968);
nor U656 (N_656,In_1026,In_560);
xor U657 (N_657,In_865,In_2461);
and U658 (N_658,In_643,In_1830);
and U659 (N_659,In_1061,In_359);
nor U660 (N_660,In_423,N_11);
nand U661 (N_661,In_1089,In_2288);
nand U662 (N_662,In_780,In_204);
nor U663 (N_663,In_589,In_1184);
nand U664 (N_664,In_2017,In_1887);
and U665 (N_665,In_659,In_1366);
nand U666 (N_666,N_214,In_1668);
and U667 (N_667,In_1972,In_840);
or U668 (N_668,In_971,In_675);
xor U669 (N_669,N_21,In_1758);
and U670 (N_670,N_488,In_999);
nor U671 (N_671,N_447,In_1855);
nor U672 (N_672,In_1900,N_340);
or U673 (N_673,In_1314,In_1291);
or U674 (N_674,In_1511,In_2109);
nor U675 (N_675,In_1218,In_131);
nand U676 (N_676,In_167,In_185);
nor U677 (N_677,In_2115,In_1343);
or U678 (N_678,In_2038,In_871);
and U679 (N_679,N_309,In_658);
and U680 (N_680,In_1022,In_480);
nor U681 (N_681,N_292,In_716);
and U682 (N_682,In_808,In_181);
and U683 (N_683,N_375,In_1954);
nor U684 (N_684,In_1117,In_1551);
and U685 (N_685,N_211,In_155);
nand U686 (N_686,In_489,In_288);
and U687 (N_687,In_111,N_483);
nor U688 (N_688,In_543,In_398);
and U689 (N_689,In_1430,In_1994);
and U690 (N_690,In_1029,In_1552);
xnor U691 (N_691,In_73,In_1358);
xor U692 (N_692,N_160,N_89);
nand U693 (N_693,In_755,N_458);
nand U694 (N_694,In_1845,N_76);
nor U695 (N_695,In_841,In_1035);
or U696 (N_696,N_202,N_300);
nand U697 (N_697,In_326,In_180);
nand U698 (N_698,In_1637,In_1352);
nor U699 (N_699,In_534,In_541);
or U700 (N_700,N_163,In_2385);
nor U701 (N_701,N_239,In_1980);
and U702 (N_702,In_604,N_70);
nand U703 (N_703,In_2104,In_1941);
nand U704 (N_704,In_2319,In_2082);
and U705 (N_705,N_187,In_237);
nand U706 (N_706,N_327,In_809);
xor U707 (N_707,N_317,In_1576);
nand U708 (N_708,In_80,N_28);
nand U709 (N_709,In_2093,In_436);
and U710 (N_710,In_236,In_1695);
or U711 (N_711,In_1287,In_1179);
nor U712 (N_712,In_1236,In_765);
nor U713 (N_713,In_1456,In_1654);
nor U714 (N_714,In_1369,In_490);
nor U715 (N_715,In_227,N_22);
nand U716 (N_716,N_499,In_852);
nor U717 (N_717,N_32,N_188);
nor U718 (N_718,N_476,In_1404);
and U719 (N_719,N_478,In_2302);
or U720 (N_720,In_571,In_725);
or U721 (N_721,In_801,N_427);
xor U722 (N_722,N_480,In_142);
and U723 (N_723,In_1053,In_312);
xnor U724 (N_724,In_924,In_600);
xor U725 (N_725,In_1070,In_2003);
nor U726 (N_726,In_673,In_1332);
and U727 (N_727,In_1310,In_2422);
nor U728 (N_728,In_1488,In_2016);
nor U729 (N_729,In_835,In_1096);
xnor U730 (N_730,In_2023,N_382);
nor U731 (N_731,In_1477,In_1097);
and U732 (N_732,In_2057,In_694);
xor U733 (N_733,In_1140,In_2377);
or U734 (N_734,In_752,In_318);
or U735 (N_735,In_294,In_132);
and U736 (N_736,In_829,In_1944);
nand U737 (N_737,N_365,N_273);
nand U738 (N_738,N_475,In_156);
nand U739 (N_739,In_705,In_1959);
nor U740 (N_740,In_1110,In_1094);
nand U741 (N_741,N_454,In_1384);
nand U742 (N_742,In_2328,N_425);
or U743 (N_743,In_2241,In_1222);
nor U744 (N_744,In_350,In_1970);
nor U745 (N_745,N_180,In_99);
nand U746 (N_746,N_337,N_141);
and U747 (N_747,In_2034,In_1176);
or U748 (N_748,N_29,In_642);
xor U749 (N_749,In_388,In_216);
or U750 (N_750,N_362,N_320);
and U751 (N_751,In_2080,N_226);
nor U752 (N_752,In_302,In_1591);
nor U753 (N_753,In_2256,In_86);
or U754 (N_754,N_384,N_436);
xnor U755 (N_755,In_935,In_1054);
and U756 (N_756,In_1387,In_2412);
or U757 (N_757,N_248,N_367);
nand U758 (N_758,In_555,In_1871);
and U759 (N_759,In_203,In_292);
nand U760 (N_760,In_401,N_242);
nor U761 (N_761,In_228,In_1167);
nand U762 (N_762,In_1392,N_174);
nand U763 (N_763,N_398,In_1968);
xor U764 (N_764,In_797,In_1226);
and U765 (N_765,In_832,In_2494);
nor U766 (N_766,In_475,In_805);
and U767 (N_767,In_822,In_501);
and U768 (N_768,In_494,In_34);
and U769 (N_769,In_763,In_580);
nand U770 (N_770,In_2039,In_880);
nand U771 (N_771,In_1788,In_1675);
nand U772 (N_772,In_775,In_1374);
xnor U773 (N_773,In_1516,In_1298);
nor U774 (N_774,In_1350,In_867);
and U775 (N_775,N_185,In_758);
nand U776 (N_776,N_59,In_949);
and U777 (N_777,N_381,In_2216);
xnor U778 (N_778,N_181,In_885);
or U779 (N_779,In_853,N_464);
nand U780 (N_780,N_240,In_1812);
or U781 (N_781,N_15,N_177);
or U782 (N_782,In_616,In_499);
or U783 (N_783,N_114,In_2191);
nor U784 (N_784,In_1978,In_2147);
nand U785 (N_785,In_2486,In_1712);
nor U786 (N_786,In_396,N_258);
or U787 (N_787,N_373,In_3);
nor U788 (N_788,In_1458,In_1422);
and U789 (N_789,In_2159,In_381);
or U790 (N_790,In_989,In_2097);
or U791 (N_791,In_901,In_973);
nand U792 (N_792,In_1895,In_815);
and U793 (N_793,In_2245,In_2106);
and U794 (N_794,In_183,N_196);
or U795 (N_795,N_54,In_1554);
nand U796 (N_796,In_943,In_2165);
and U797 (N_797,N_383,In_2144);
or U798 (N_798,N_473,N_39);
xnor U799 (N_799,In_460,N_429);
nand U800 (N_800,N_262,In_323);
nor U801 (N_801,N_388,In_152);
or U802 (N_802,N_397,N_218);
or U803 (N_803,In_1700,In_389);
nand U804 (N_804,In_737,In_286);
or U805 (N_805,N_38,In_84);
nor U806 (N_806,In_5,In_128);
nand U807 (N_807,In_1024,In_1224);
and U808 (N_808,In_2033,In_1613);
nand U809 (N_809,In_1125,In_2131);
or U810 (N_810,In_2469,In_2170);
xnor U811 (N_811,N_307,In_1227);
nor U812 (N_812,In_1192,In_1292);
nand U813 (N_813,In_1597,N_119);
and U814 (N_814,In_2157,In_1406);
nand U815 (N_815,N_125,In_1540);
nand U816 (N_816,N_64,N_461);
xnor U817 (N_817,In_199,In_1835);
or U818 (N_818,In_1262,In_1617);
or U819 (N_819,In_1412,In_2043);
nor U820 (N_820,In_1873,In_1572);
nor U821 (N_821,In_2493,In_1144);
xnor U822 (N_822,N_8,N_385);
nand U823 (N_823,In_537,N_112);
and U824 (N_824,N_434,In_1077);
or U825 (N_825,In_861,In_2320);
and U826 (N_826,In_1339,In_394);
or U827 (N_827,In_614,N_17);
nor U828 (N_828,In_1393,N_441);
or U829 (N_829,In_2268,N_403);
and U830 (N_830,In_990,In_2456);
nor U831 (N_831,In_1929,In_1190);
nand U832 (N_832,In_1055,N_423);
nand U833 (N_833,In_18,In_2374);
nor U834 (N_834,In_2294,In_626);
nor U835 (N_835,In_2478,In_783);
or U836 (N_836,In_1610,In_2083);
nand U837 (N_837,In_335,In_257);
nand U838 (N_838,In_933,In_1564);
nor U839 (N_839,In_1188,In_81);
nand U840 (N_840,N_455,In_2113);
xor U841 (N_841,In_1383,In_304);
or U842 (N_842,In_1288,N_166);
nand U843 (N_843,In_59,In_582);
xor U844 (N_844,N_335,In_1690);
nand U845 (N_845,In_2058,N_154);
xor U846 (N_846,N_126,N_276);
nor U847 (N_847,In_789,In_1765);
nor U848 (N_848,In_590,N_73);
nor U849 (N_849,In_277,In_473);
and U850 (N_850,N_191,In_488);
nand U851 (N_851,In_2358,N_201);
nor U852 (N_852,In_918,In_2225);
and U853 (N_853,In_158,In_1593);
or U854 (N_854,N_308,In_2188);
and U855 (N_855,N_195,In_369);
or U856 (N_856,In_2158,In_1609);
xor U857 (N_857,N_111,In_2271);
or U858 (N_858,In_1649,N_158);
nand U859 (N_859,In_1709,In_2192);
nor U860 (N_860,N_324,In_579);
and U861 (N_861,In_1391,N_310);
nor U862 (N_862,N_369,In_547);
nor U863 (N_863,In_1413,N_422);
nor U864 (N_864,In_1949,N_272);
and U865 (N_865,N_97,In_747);
xnor U866 (N_866,In_1058,In_868);
and U867 (N_867,In_1088,In_1259);
nand U868 (N_868,N_94,In_2482);
or U869 (N_869,In_1371,N_2);
xor U870 (N_870,In_2052,N_61);
and U871 (N_871,N_74,In_66);
or U872 (N_872,In_55,In_1679);
and U873 (N_873,In_1995,In_1822);
xor U874 (N_874,In_1594,In_2465);
and U875 (N_875,In_325,In_821);
or U876 (N_876,In_1558,In_2423);
or U877 (N_877,In_362,In_1080);
nor U878 (N_878,In_1841,In_739);
and U879 (N_879,In_225,N_216);
and U880 (N_880,In_1410,N_93);
or U881 (N_881,N_352,In_2086);
nand U882 (N_882,In_374,In_1566);
and U883 (N_883,In_1878,In_1232);
nand U884 (N_884,In_2462,N_68);
or U885 (N_885,In_176,In_1604);
nand U886 (N_886,In_768,N_378);
and U887 (N_887,In_942,In_1076);
and U888 (N_888,In_696,In_2370);
nor U889 (N_889,In_1354,In_948);
nand U890 (N_890,N_127,In_779);
and U891 (N_891,In_2014,N_463);
and U892 (N_892,In_911,In_811);
or U893 (N_893,In_1803,In_266);
nand U894 (N_894,N_104,N_453);
nor U895 (N_895,In_2148,In_232);
nor U896 (N_896,In_483,N_401);
nor U897 (N_897,N_67,In_890);
or U898 (N_898,In_1411,In_2293);
or U899 (N_899,In_1420,In_1638);
xor U900 (N_900,N_264,In_1828);
nand U901 (N_901,In_1137,In_1681);
and U902 (N_902,N_27,N_416);
nand U903 (N_903,In_42,In_1130);
or U904 (N_904,In_689,In_863);
and U905 (N_905,In_762,N_363);
and U906 (N_906,In_2390,In_1014);
and U907 (N_907,N_215,In_2466);
nor U908 (N_908,N_406,N_331);
and U909 (N_909,In_778,N_135);
nand U910 (N_910,In_1036,N_279);
nand U911 (N_911,In_1175,In_833);
nor U912 (N_912,N_394,In_1507);
nor U913 (N_913,In_58,N_12);
nor U914 (N_914,In_1826,In_524);
nand U915 (N_915,N_88,In_1023);
and U916 (N_916,In_2091,In_1625);
and U917 (N_917,N_138,In_336);
or U918 (N_918,N_489,In_1051);
or U919 (N_919,In_344,N_498);
or U920 (N_920,In_2259,In_2066);
and U921 (N_921,In_1883,N_26);
or U922 (N_922,In_914,In_2130);
nor U923 (N_923,In_1590,N_116);
nand U924 (N_924,N_277,In_212);
nor U925 (N_925,In_1584,N_16);
xor U926 (N_926,In_978,In_1704);
and U927 (N_927,In_900,N_238);
nand U928 (N_928,N_145,In_530);
nor U929 (N_929,In_608,In_1124);
nor U930 (N_930,N_470,N_351);
or U931 (N_931,In_1549,In_1538);
nor U932 (N_932,In_1186,In_1726);
nor U933 (N_933,In_1570,In_1881);
nor U934 (N_934,N_302,In_2020);
nor U935 (N_935,In_769,In_842);
nand U936 (N_936,In_1378,In_101);
or U937 (N_937,In_985,N_313);
and U938 (N_938,In_331,N_465);
nand U939 (N_939,In_995,N_203);
or U940 (N_940,In_1414,N_165);
nand U941 (N_941,In_1719,In_1265);
and U942 (N_942,In_1153,In_1349);
or U943 (N_943,In_472,In_2404);
and U944 (N_944,In_722,In_1028);
nand U945 (N_945,In_882,In_157);
or U946 (N_946,N_379,In_591);
and U947 (N_947,In_270,In_2498);
and U948 (N_948,N_410,In_1770);
or U949 (N_949,In_1191,In_592);
or U950 (N_950,In_210,In_1248);
nor U951 (N_951,In_692,N_437);
and U952 (N_952,In_2352,In_1623);
and U953 (N_953,In_364,N_42);
nand U954 (N_954,In_638,In_230);
nand U955 (N_955,In_531,In_872);
and U956 (N_956,N_91,In_1592);
nand U957 (N_957,In_945,In_387);
nor U958 (N_958,N_482,N_14);
nand U959 (N_959,In_1896,N_295);
nor U960 (N_960,N_182,In_348);
nor U961 (N_961,In_2264,N_449);
or U962 (N_962,In_134,In_1722);
nor U963 (N_963,N_479,In_1555);
or U964 (N_964,In_470,N_387);
xnor U965 (N_965,N_47,In_220);
and U966 (N_966,N_303,In_2291);
or U967 (N_967,In_1021,In_1367);
or U968 (N_968,In_1682,In_851);
xor U969 (N_969,In_2160,In_1438);
and U970 (N_970,In_1450,In_1852);
and U971 (N_971,In_1517,N_452);
and U972 (N_972,In_205,N_134);
nand U973 (N_973,N_45,In_1727);
nor U974 (N_974,N_13,In_1791);
nor U975 (N_975,N_376,In_1991);
nand U976 (N_976,In_2477,N_217);
xor U977 (N_977,In_1936,In_322);
and U978 (N_978,In_2068,In_1465);
nor U979 (N_979,N_31,N_344);
nand U980 (N_980,In_2217,In_1122);
nor U981 (N_981,In_1930,In_2064);
nor U982 (N_982,In_542,In_96);
nand U983 (N_983,In_1696,N_377);
xor U984 (N_984,In_1085,In_2251);
nand U985 (N_985,In_922,In_2332);
and U986 (N_986,In_1536,N_329);
nand U987 (N_987,In_2451,N_120);
xor U988 (N_988,N_124,N_466);
or U989 (N_989,In_1178,In_2428);
nor U990 (N_990,N_252,In_2297);
and U991 (N_991,N_278,In_69);
nor U992 (N_992,In_1429,In_759);
nor U993 (N_993,N_96,N_49);
xnor U994 (N_994,N_34,In_124);
or U995 (N_995,In_921,In_1398);
and U996 (N_996,In_2394,In_1815);
nor U997 (N_997,In_2185,In_712);
or U998 (N_998,N_430,In_1015);
nand U999 (N_999,In_2345,In_1455);
nor U1000 (N_1000,In_1736,In_700);
nand U1001 (N_1001,In_1173,N_596);
or U1002 (N_1002,In_1793,N_580);
xnor U1003 (N_1003,In_214,In_1099);
or U1004 (N_1004,In_955,In_442);
xnor U1005 (N_1005,N_130,In_2050);
or U1006 (N_1006,In_2061,N_832);
and U1007 (N_1007,N_493,In_106);
nand U1008 (N_1008,N_670,In_1985);
nand U1009 (N_1009,N_921,N_615);
and U1010 (N_1010,N_731,N_749);
and U1011 (N_1011,In_2387,N_702);
nor U1012 (N_1012,N_200,In_1165);
xor U1013 (N_1013,N_958,In_1275);
and U1014 (N_1014,N_595,In_64);
xnor U1015 (N_1015,N_443,N_993);
nor U1016 (N_1016,N_831,In_956);
or U1017 (N_1017,N_847,N_502);
nor U1018 (N_1018,N_708,N_769);
or U1019 (N_1019,In_619,In_607);
nor U1020 (N_1020,N_176,In_174);
and U1021 (N_1021,N_880,In_1496);
nand U1022 (N_1022,In_1821,N_729);
and U1023 (N_1023,N_0,In_646);
nor U1024 (N_1024,N_129,In_1284);
nand U1025 (N_1025,N_72,N_996);
and U1026 (N_1026,In_2174,N_805);
and U1027 (N_1027,In_1577,N_767);
nor U1028 (N_1028,In_1007,In_1415);
nor U1029 (N_1029,N_678,N_190);
nand U1030 (N_1030,In_2219,N_321);
and U1031 (N_1031,N_288,N_213);
nor U1032 (N_1032,N_546,In_1616);
or U1033 (N_1033,In_1518,In_1293);
or U1034 (N_1034,N_598,N_208);
and U1035 (N_1035,In_803,In_1373);
nor U1036 (N_1036,In_2392,In_1882);
and U1037 (N_1037,In_634,In_1526);
nand U1038 (N_1038,In_635,In_1915);
nor U1039 (N_1039,N_763,N_680);
xor U1040 (N_1040,N_495,In_1254);
nand U1041 (N_1041,In_1142,N_524);
or U1042 (N_1042,N_314,In_528);
and U1043 (N_1043,In_1606,In_1605);
nand U1044 (N_1044,N_518,N_528);
nor U1045 (N_1045,N_552,N_793);
and U1046 (N_1046,In_258,N_757);
or U1047 (N_1047,In_994,In_1961);
and U1048 (N_1048,N_396,In_118);
nand U1049 (N_1049,In_2371,In_1500);
nor U1050 (N_1050,In_2069,In_201);
and U1051 (N_1051,In_143,N_40);
nand U1052 (N_1052,In_1421,In_327);
nor U1053 (N_1053,N_616,In_2046);
xnor U1054 (N_1054,In_1989,N_56);
nand U1055 (N_1055,N_646,In_974);
nor U1056 (N_1056,N_705,N_940);
nand U1057 (N_1057,N_792,N_339);
and U1058 (N_1058,In_2075,In_1479);
nand U1059 (N_1059,N_123,In_539);
nor U1060 (N_1060,In_1908,In_1761);
or U1061 (N_1061,N_913,In_108);
or U1062 (N_1062,In_2028,N_799);
nor U1063 (N_1063,In_467,In_1666);
nand U1064 (N_1064,In_2444,In_233);
nand U1065 (N_1065,In_1737,N_746);
nor U1066 (N_1066,In_1676,In_2230);
and U1067 (N_1067,In_1921,In_428);
and U1068 (N_1068,N_600,In_1462);
nand U1069 (N_1069,N_632,In_1642);
xor U1070 (N_1070,N_759,In_262);
nand U1071 (N_1071,In_1467,In_1376);
or U1072 (N_1072,In_800,In_1271);
nor U1073 (N_1073,N_156,In_1759);
xor U1074 (N_1074,In_177,In_799);
and U1075 (N_1075,N_990,N_578);
nor U1076 (N_1076,N_970,N_718);
nor U1077 (N_1077,N_950,N_304);
nand U1078 (N_1078,N_33,In_1849);
nor U1079 (N_1079,In_315,In_1260);
and U1080 (N_1080,In_2325,In_777);
or U1081 (N_1081,N_699,In_2421);
nand U1082 (N_1082,N_175,In_538);
or U1083 (N_1083,N_789,N_153);
or U1084 (N_1084,N_467,In_1854);
and U1085 (N_1085,In_1678,N_147);
nor U1086 (N_1086,N_654,In_246);
nor U1087 (N_1087,In_1631,N_694);
nand U1088 (N_1088,N_618,N_490);
xor U1089 (N_1089,N_280,N_931);
or U1090 (N_1090,N_400,In_75);
or U1091 (N_1091,N_863,N_517);
and U1092 (N_1092,N_684,N_612);
and U1093 (N_1093,In_360,In_1506);
and U1094 (N_1094,N_421,N_148);
xnor U1095 (N_1095,In_393,In_1899);
and U1096 (N_1096,In_2199,In_2239);
nand U1097 (N_1097,N_802,In_2312);
and U1098 (N_1098,In_1032,N_63);
nand U1099 (N_1099,In_2146,In_1874);
xnor U1100 (N_1100,N_856,N_703);
nand U1101 (N_1101,In_90,In_1286);
nor U1102 (N_1102,N_819,In_2270);
nor U1103 (N_1103,In_1692,N_583);
and U1104 (N_1104,In_1136,N_593);
nand U1105 (N_1105,In_2059,N_700);
xnor U1106 (N_1106,N_263,N_41);
nand U1107 (N_1107,In_1397,In_702);
nand U1108 (N_1108,N_587,In_432);
nand U1109 (N_1109,In_927,N_982);
nand U1110 (N_1110,In_2333,N_509);
nor U1111 (N_1111,In_810,N_933);
xnor U1112 (N_1112,In_794,N_834);
or U1113 (N_1113,N_814,N_927);
and U1114 (N_1114,In_1585,In_1075);
nor U1115 (N_1115,In_340,N_143);
nor U1116 (N_1116,In_2310,In_553);
nor U1117 (N_1117,N_959,N_102);
xor U1118 (N_1118,N_888,N_567);
and U1119 (N_1119,In_2402,In_329);
nand U1120 (N_1120,In_533,In_613);
and U1121 (N_1121,In_378,In_1143);
or U1122 (N_1122,N_768,In_844);
and U1123 (N_1123,N_878,In_1799);
and U1124 (N_1124,In_1220,N_445);
nor U1125 (N_1125,In_500,N_777);
nand U1126 (N_1126,N_906,In_1975);
nand U1127 (N_1127,In_2414,In_1713);
and U1128 (N_1128,N_361,In_186);
nand U1129 (N_1129,In_1466,N_658);
or U1130 (N_1130,N_444,N_576);
nor U1131 (N_1131,N_512,In_2124);
nand U1132 (N_1132,N_286,N_350);
nand U1133 (N_1133,In_2150,In_487);
nand U1134 (N_1134,N_765,N_810);
and U1135 (N_1135,N_301,N_243);
and U1136 (N_1136,In_440,N_922);
and U1137 (N_1137,In_691,In_1244);
or U1138 (N_1138,In_1697,In_1739);
nor U1139 (N_1139,In_2400,In_650);
or U1140 (N_1140,In_683,N_456);
xnor U1141 (N_1141,In_463,N_743);
or U1142 (N_1142,In_2260,N_771);
and U1143 (N_1143,N_219,In_1816);
xnor U1144 (N_1144,In_983,In_2441);
nor U1145 (N_1145,In_1017,N_811);
and U1146 (N_1146,In_1533,N_661);
nand U1147 (N_1147,N_347,N_839);
xnor U1148 (N_1148,In_1148,N_469);
nor U1149 (N_1149,In_804,In_1242);
nor U1150 (N_1150,N_669,N_693);
and U1151 (N_1151,In_1289,In_2350);
and U1152 (N_1152,N_837,In_1439);
nand U1153 (N_1153,N_774,In_1567);
and U1154 (N_1154,N_969,N_5);
nand U1155 (N_1155,In_1760,In_1000);
and U1156 (N_1156,N_671,In_1750);
or U1157 (N_1157,In_1461,N_275);
or U1158 (N_1158,N_107,In_2139);
and U1159 (N_1159,N_515,N_391);
nor U1160 (N_1160,N_233,In_979);
nand U1161 (N_1161,N_626,N_904);
or U1162 (N_1162,In_2022,In_1205);
and U1163 (N_1163,N_513,N_169);
nor U1164 (N_1164,In_1792,In_1916);
nand U1165 (N_1165,N_591,N_782);
or U1166 (N_1166,N_1,In_665);
nor U1167 (N_1167,N_254,In_726);
nand U1168 (N_1168,In_1361,N_672);
xnor U1169 (N_1169,In_29,N_508);
xor U1170 (N_1170,N_142,In_1652);
nand U1171 (N_1171,In_2084,In_1149);
and U1172 (N_1172,N_627,N_850);
nor U1173 (N_1173,N_800,In_575);
or U1174 (N_1174,N_884,N_836);
nor U1175 (N_1175,In_217,N_988);
nor U1176 (N_1176,N_250,N_696);
nand U1177 (N_1177,N_649,In_452);
nor U1178 (N_1178,In_2229,N_642);
xor U1179 (N_1179,N_634,N_9);
xor U1180 (N_1180,In_144,In_670);
nor U1181 (N_1181,N_869,N_812);
and U1182 (N_1182,In_1902,In_1263);
or U1183 (N_1183,N_650,N_797);
xnor U1184 (N_1184,N_909,N_395);
nor U1185 (N_1185,In_937,In_1839);
and U1186 (N_1186,In_1879,In_1504);
nor U1187 (N_1187,In_830,N_544);
or U1188 (N_1188,In_2223,In_76);
nor U1189 (N_1189,N_784,N_336);
or U1190 (N_1190,In_926,In_1212);
and U1191 (N_1191,N_930,In_773);
nor U1192 (N_1192,N_52,N_249);
or U1193 (N_1193,In_946,N_282);
and U1194 (N_1194,In_1215,N_999);
nand U1195 (N_1195,In_2128,N_870);
or U1196 (N_1196,In_1782,In_2376);
nand U1197 (N_1197,N_605,N_323);
nand U1198 (N_1198,N_366,In_2261);
xnor U1199 (N_1199,N_750,N_891);
xnor U1200 (N_1200,In_2242,In_243);
or U1201 (N_1201,N_758,N_636);
or U1202 (N_1202,N_977,In_2202);
or U1203 (N_1203,In_1322,In_122);
nor U1204 (N_1204,In_1742,In_870);
nor U1205 (N_1205,N_677,N_798);
or U1206 (N_1206,In_1441,N_326);
nand U1207 (N_1207,N_944,In_1408);
nor U1208 (N_1208,N_505,In_1155);
and U1209 (N_1209,N_978,In_878);
or U1210 (N_1210,In_482,N_79);
or U1211 (N_1211,In_2056,In_1313);
nand U1212 (N_1212,N_620,In_1880);
or U1213 (N_1213,N_232,N_617);
xnor U1214 (N_1214,N_115,N_916);
nor U1215 (N_1215,N_548,N_701);
and U1216 (N_1216,In_2208,N_579);
xnor U1217 (N_1217,In_1433,In_519);
and U1218 (N_1218,N_803,In_1497);
and U1219 (N_1219,In_9,N_46);
or U1220 (N_1220,N_564,N_543);
or U1221 (N_1221,N_589,N_861);
or U1222 (N_1222,In_2025,N_523);
or U1223 (N_1223,In_197,In_41);
nor U1224 (N_1224,In_703,In_1940);
or U1225 (N_1225,In_2065,N_796);
nand U1226 (N_1226,N_328,In_1325);
xor U1227 (N_1227,In_764,In_16);
nor U1228 (N_1228,In_1962,In_1345);
and U1229 (N_1229,N_625,In_1987);
and U1230 (N_1230,N_534,N_961);
nand U1231 (N_1231,N_735,N_657);
and U1232 (N_1232,In_1562,N_934);
or U1233 (N_1233,N_161,N_297);
or U1234 (N_1234,In_754,In_1983);
nand U1235 (N_1235,In_1784,In_883);
or U1236 (N_1236,In_2140,In_1452);
nand U1237 (N_1237,N_712,N_776);
nor U1238 (N_1238,N_81,In_2408);
and U1239 (N_1239,N_965,In_2090);
or U1240 (N_1240,N_786,N_24);
nand U1241 (N_1241,In_690,In_1372);
nor U1242 (N_1242,In_1664,N_225);
nand U1243 (N_1243,N_137,N_845);
and U1244 (N_1244,In_65,In_2);
and U1245 (N_1245,N_736,In_970);
xor U1246 (N_1246,N_915,N_984);
xnor U1247 (N_1247,N_266,N_840);
xnor U1248 (N_1248,N_898,N_644);
and U1249 (N_1249,N_569,N_848);
nor U1250 (N_1250,N_737,N_537);
nand U1251 (N_1251,In_1407,N_808);
nand U1252 (N_1252,N_53,In_919);
xor U1253 (N_1253,In_2094,In_2030);
nand U1254 (N_1254,In_1598,In_2401);
and U1255 (N_1255,N_474,In_1238);
and U1256 (N_1256,In_453,N_873);
xor U1257 (N_1257,N_868,In_823);
nand U1258 (N_1258,N_575,N_597);
nor U1259 (N_1259,N_539,N_963);
and U1260 (N_1260,N_562,In_141);
nor U1261 (N_1261,N_622,N_588);
nor U1262 (N_1262,N_954,In_1847);
or U1263 (N_1263,N_289,In_1958);
nor U1264 (N_1264,N_10,In_2155);
and U1265 (N_1265,In_846,In_2204);
nor U1266 (N_1266,N_791,In_2029);
nor U1267 (N_1267,N_715,N_409);
nand U1268 (N_1268,N_140,N_484);
and U1269 (N_1269,In_430,N_841);
nand U1270 (N_1270,N_720,N_770);
or U1271 (N_1271,In_1707,In_1509);
and U1272 (N_1272,In_2072,In_631);
or U1273 (N_1273,N_752,N_168);
nand U1274 (N_1274,In_1390,N_917);
xor U1275 (N_1275,In_1426,N_210);
and U1276 (N_1276,In_2079,N_481);
and U1277 (N_1277,In_932,In_569);
or U1278 (N_1278,N_222,In_857);
xor U1279 (N_1279,In_2214,N_519);
xor U1280 (N_1280,N_714,In_367);
and U1281 (N_1281,In_1751,N_241);
nand U1282 (N_1282,In_2309,N_566);
or U1283 (N_1283,In_115,In_1805);
nor U1284 (N_1284,N_496,N_973);
nand U1285 (N_1285,In_308,In_1362);
xor U1286 (N_1286,In_2300,N_860);
xor U1287 (N_1287,N_725,N_635);
or U1288 (N_1288,In_1804,N_251);
nand U1289 (N_1289,N_885,In_2459);
or U1290 (N_1290,In_249,N_882);
xnor U1291 (N_1291,In_1253,In_699);
or U1292 (N_1292,In_1906,In_1789);
or U1293 (N_1293,N_829,In_2435);
or U1294 (N_1294,In_680,In_206);
nor U1295 (N_1295,In_965,In_1575);
nand U1296 (N_1296,N_521,In_415);
xor U1297 (N_1297,In_114,In_2031);
nor U1298 (N_1298,In_1281,N_986);
xnor U1299 (N_1299,In_1923,N_937);
or U1300 (N_1300,N_507,N_925);
or U1301 (N_1301,N_173,N_641);
nor U1302 (N_1302,N_924,N_865);
nor U1303 (N_1303,In_1025,N_345);
nor U1304 (N_1304,N_604,N_957);
nand U1305 (N_1305,N_881,In_1171);
or U1306 (N_1306,In_133,In_1928);
nor U1307 (N_1307,In_1714,In_1006);
nand U1308 (N_1308,In_1514,N_433);
nand U1309 (N_1309,In_40,N_926);
or U1310 (N_1310,In_446,In_2485);
nand U1311 (N_1311,In_649,In_2145);
or U1312 (N_1312,N_551,In_1833);
and U1313 (N_1313,N_451,N_371);
nor U1314 (N_1314,N_899,N_44);
nor U1315 (N_1315,N_573,In_1246);
or U1316 (N_1316,In_72,In_2010);
nand U1317 (N_1317,N_438,In_1385);
nor U1318 (N_1318,In_276,N_257);
nor U1319 (N_1319,In_196,N_610);
nor U1320 (N_1320,In_2269,In_11);
xnor U1321 (N_1321,N_806,In_807);
nor U1322 (N_1322,N_908,N_716);
nor U1323 (N_1323,N_665,In_2134);
xnor U1324 (N_1324,N_664,In_1614);
and U1325 (N_1325,N_655,In_2415);
and U1326 (N_1326,N_619,N_540);
xor U1327 (N_1327,N_267,N_951);
nor U1328 (N_1328,N_150,In_641);
nor U1329 (N_1329,N_374,In_2213);
nand U1330 (N_1330,N_709,N_581);
nor U1331 (N_1331,N_666,N_471);
nand U1332 (N_1332,N_189,N_651);
or U1333 (N_1333,In_2000,In_1331);
and U1334 (N_1334,In_1078,In_1946);
or U1335 (N_1335,In_252,In_1474);
and U1336 (N_1336,N_285,In_2396);
nor U1337 (N_1337,N_823,N_592);
or U1338 (N_1338,N_717,N_603);
nand U1339 (N_1339,N_283,N_945);
and U1340 (N_1340,In_1969,In_2326);
and U1341 (N_1341,In_85,In_1494);
and U1342 (N_1342,N_526,In_1480);
xor U1343 (N_1343,N_101,In_1073);
and U1344 (N_1344,In_242,N_887);
and U1345 (N_1345,In_1396,N_815);
or U1346 (N_1346,N_849,N_639);
nand U1347 (N_1347,N_942,In_551);
xor U1348 (N_1348,N_943,In_77);
or U1349 (N_1349,N_689,In_383);
and U1350 (N_1350,N_955,In_339);
or U1351 (N_1351,In_2279,In_997);
nand U1352 (N_1352,In_2013,In_188);
xor U1353 (N_1353,N_205,N_876);
or U1354 (N_1354,In_1963,N_713);
xnor U1355 (N_1355,N_186,N_773);
nand U1356 (N_1356,N_192,N_609);
or U1357 (N_1357,N_477,N_872);
nor U1358 (N_1358,N_133,In_410);
or U1359 (N_1359,In_1104,N_974);
xnor U1360 (N_1360,N_998,In_864);
and U1361 (N_1361,In_506,N_529);
nand U1362 (N_1362,In_728,In_734);
xor U1363 (N_1363,In_289,N_305);
or U1364 (N_1364,N_392,N_911);
nand U1365 (N_1365,In_1151,N_938);
or U1366 (N_1366,N_660,In_1646);
and U1367 (N_1367,N_952,N_762);
and U1368 (N_1368,N_807,N_785);
nor U1369 (N_1369,N_662,In_859);
nor U1370 (N_1370,In_1316,N_570);
or U1371 (N_1371,N_724,N_602);
nand U1372 (N_1372,N_66,N_695);
xor U1373 (N_1373,N_48,N_674);
nand U1374 (N_1374,N_795,N_525);
or U1375 (N_1375,In_1798,N_65);
or U1376 (N_1376,N_907,In_1072);
nand U1377 (N_1377,N_359,N_844);
nor U1378 (N_1378,N_334,N_462);
and U1379 (N_1379,N_966,N_902);
nand U1380 (N_1380,N_647,N_404);
or U1381 (N_1381,N_230,N_867);
or U1382 (N_1382,In_834,In_521);
and U1383 (N_1383,N_753,In_546);
xor U1384 (N_1384,In_1581,N_228);
xor U1385 (N_1385,In_982,In_1964);
nand U1386 (N_1386,In_1468,In_1611);
and U1387 (N_1387,In_1733,In_1365);
nand U1388 (N_1388,In_1768,In_2249);
nand U1389 (N_1389,N_405,N_554);
or U1390 (N_1390,In_226,In_1767);
xnor U1391 (N_1391,In_529,In_2246);
or U1392 (N_1392,N_287,In_1884);
xnor U1393 (N_1393,In_2453,N_402);
nand U1394 (N_1394,N_659,In_796);
or U1395 (N_1395,In_2042,In_637);
nand U1396 (N_1396,N_486,N_676);
xnor U1397 (N_1397,In_2343,In_907);
nand U1398 (N_1398,N_682,In_1214);
nor U1399 (N_1399,In_570,N_360);
nand U1400 (N_1400,In_2321,In_474);
or U1401 (N_1401,N_653,N_164);
nor U1402 (N_1402,N_740,N_772);
or U1403 (N_1403,In_1769,In_2110);
or U1404 (N_1404,In_2254,N_500);
or U1405 (N_1405,N_804,N_920);
xor U1406 (N_1406,In_1133,N_172);
and U1407 (N_1407,N_706,In_1519);
nor U1408 (N_1408,In_858,N_183);
nor U1409 (N_1409,In_303,In_1524);
nor U1410 (N_1410,N_992,In_925);
or U1411 (N_1411,N_281,In_264);
and U1412 (N_1412,In_456,In_915);
nor U1413 (N_1413,N_261,In_51);
nand U1414 (N_1414,In_678,N_346);
nor U1415 (N_1415,In_790,N_440);
and U1416 (N_1416,In_2403,N_809);
nand U1417 (N_1417,In_48,In_1353);
nor U1418 (N_1418,In_629,N_599);
and U1419 (N_1419,N_892,N_981);
or U1420 (N_1420,N_613,N_745);
and U1421 (N_1421,In_2305,In_2395);
nand U1422 (N_1422,In_1905,N_516);
and U1423 (N_1423,In_1748,N_656);
and U1424 (N_1424,In_368,N_889);
nor U1425 (N_1425,N_155,N_37);
and U1426 (N_1426,In_743,In_241);
xor U1427 (N_1427,N_235,N_726);
nand U1428 (N_1428,N_825,N_851);
nor U1429 (N_1429,In_1580,In_2012);
nand U1430 (N_1430,In_179,N_614);
xnor U1431 (N_1431,In_917,N_586);
nor U1432 (N_1432,In_239,In_405);
nor U1433 (N_1433,In_2373,In_1624);
nor U1434 (N_1434,N_914,N_550);
or U1435 (N_1435,In_445,N_419);
nor U1436 (N_1436,In_836,In_1548);
nand U1437 (N_1437,In_391,In_2085);
xnor U1438 (N_1438,In_1340,N_390);
nor U1439 (N_1439,In_784,N_895);
nand U1440 (N_1440,N_935,N_685);
and U1441 (N_1441,In_1196,In_1417);
nand U1442 (N_1442,In_2399,N_584);
nor U1443 (N_1443,N_817,N_590);
nand U1444 (N_1444,In_1195,In_386);
or U1445 (N_1445,In_622,In_969);
nor U1446 (N_1446,In_2443,N_207);
and U1447 (N_1447,N_901,N_864);
nor U1448 (N_1448,N_948,N_103);
and U1449 (N_1449,In_400,In_278);
nand U1450 (N_1450,In_893,N_989);
and U1451 (N_1451,In_1911,In_324);
or U1452 (N_1452,In_1300,N_318);
xnor U1453 (N_1453,In_1531,N_585);
or U1454 (N_1454,In_1943,In_1134);
xor U1455 (N_1455,In_291,In_624);
nor U1456 (N_1456,In_352,N_987);
xnor U1457 (N_1457,N_354,N_820);
xnor U1458 (N_1458,In_2425,In_1105);
and U1459 (N_1459,In_1848,In_1283);
nor U1460 (N_1460,In_2313,In_1660);
nand U1461 (N_1461,N_290,In_1264);
nor U1462 (N_1462,N_722,In_1095);
or U1463 (N_1463,In_1628,N_707);
xor U1464 (N_1464,N_691,N_533);
nor U1465 (N_1465,In_544,In_485);
nor U1466 (N_1466,In_370,In_2418);
nand U1467 (N_1467,In_2324,In_413);
or U1468 (N_1468,In_2222,N_890);
nor U1469 (N_1469,In_1677,N_751);
nand U1470 (N_1470,In_437,N_50);
and U1471 (N_1471,N_742,N_721);
or U1472 (N_1472,N_683,N_417);
and U1473 (N_1473,In_2032,N_883);
xnor U1474 (N_1474,N_608,N_628);
and U1475 (N_1475,N_962,N_547);
or U1476 (N_1476,In_653,In_1658);
nor U1477 (N_1477,N_556,In_517);
or U1478 (N_1478,In_2470,N_673);
nor U1479 (N_1479,N_910,N_754);
nand U1480 (N_1480,In_2210,N_535);
and U1481 (N_1481,In_1728,N_755);
or U1482 (N_1482,N_298,N_284);
or U1483 (N_1483,N_900,N_734);
nor U1484 (N_1484,N_688,N_511);
and U1485 (N_1485,In_1571,N_739);
xnor U1486 (N_1486,In_1005,In_1194);
or U1487 (N_1487,N_723,N_358);
nor U1488 (N_1488,In_1744,In_1634);
xor U1489 (N_1489,N_221,In_2194);
nand U1490 (N_1490,In_2355,N_624);
and U1491 (N_1491,N_100,In_902);
or U1492 (N_1492,N_788,In_839);
or U1493 (N_1493,N_342,N_370);
xor U1494 (N_1494,In_1665,In_1843);
and U1495 (N_1495,In_2359,N_853);
and U1496 (N_1496,N_23,N_818);
nor U1497 (N_1497,N_947,In_491);
nand U1498 (N_1498,In_112,N_794);
or U1499 (N_1499,In_630,In_862);
nand U1500 (N_1500,N_936,N_1058);
or U1501 (N_1501,N_645,In_311);
xnor U1502 (N_1502,N_1093,N_1232);
and U1503 (N_1503,N_1204,N_1210);
or U1504 (N_1504,N_1092,N_1485);
xnor U1505 (N_1505,N_1476,N_58);
nor U1506 (N_1506,N_687,In_1047);
and U1507 (N_1507,N_918,N_1088);
nand U1508 (N_1508,N_1444,In_411);
nand U1509 (N_1509,N_1394,N_1446);
and U1510 (N_1510,N_1033,N_1487);
xnor U1511 (N_1511,In_605,N_1284);
nand U1512 (N_1512,N_1097,N_949);
and U1513 (N_1513,N_1360,N_532);
and U1514 (N_1514,N_260,N_577);
xor U1515 (N_1515,N_1380,N_1491);
xor U1516 (N_1516,In_2051,In_195);
nand U1517 (N_1517,N_1280,In_2258);
and U1518 (N_1518,In_2129,N_879);
nor U1519 (N_1519,N_1013,N_1313);
and U1520 (N_1520,N_1340,N_652);
nand U1521 (N_1521,N_1197,In_1121);
or U1522 (N_1522,N_1129,In_1473);
xor U1523 (N_1523,N_1163,N_1483);
nand U1524 (N_1524,N_1264,N_1249);
and U1525 (N_1525,N_1403,N_821);
nand U1526 (N_1526,N_565,N_82);
nor U1527 (N_1527,N_1416,N_1443);
or U1528 (N_1528,N_1477,N_813);
nor U1529 (N_1529,N_1332,N_1229);
xnor U1530 (N_1530,N_1192,N_1381);
nand U1531 (N_1531,N_522,N_253);
nand U1532 (N_1532,In_2126,N_1470);
nor U1533 (N_1533,N_1304,In_1403);
and U1534 (N_1534,N_1318,N_1302);
and U1535 (N_1535,N_855,N_1005);
or U1536 (N_1536,N_690,N_415);
and U1537 (N_1537,In_598,N_194);
nand U1538 (N_1538,N_1344,N_1306);
xor U1539 (N_1539,N_1189,In_1706);
nor U1540 (N_1540,N_1140,N_1326);
or U1541 (N_1541,In_2135,N_866);
nor U1542 (N_1542,N_19,N_995);
and U1543 (N_1543,N_1037,N_538);
xnor U1544 (N_1544,In_495,N_86);
and U1545 (N_1545,N_1267,N_204);
nand U1546 (N_1546,N_389,N_1365);
nor U1547 (N_1547,In_679,N_1274);
or U1548 (N_1548,N_728,N_1172);
nor U1549 (N_1549,N_1373,In_1801);
nor U1550 (N_1550,N_1110,N_1357);
and U1551 (N_1551,In_238,N_1199);
nand U1552 (N_1552,N_1074,In_1086);
and U1553 (N_1553,N_824,N_1301);
or U1554 (N_1554,In_2311,N_1227);
nor U1555 (N_1555,N_1029,N_1134);
and U1556 (N_1556,N_1475,In_1586);
or U1557 (N_1557,N_1495,N_1441);
and U1558 (N_1558,N_748,In_2224);
and U1559 (N_1559,N_1269,N_1182);
nand U1560 (N_1560,N_1109,N_1174);
and U1561 (N_1561,In_221,N_1328);
nand U1562 (N_1562,N_1261,N_1399);
and U1563 (N_1563,In_1582,In_617);
and U1564 (N_1564,In_172,N_1464);
nand U1565 (N_1565,N_265,N_1171);
nor U1566 (N_1566,N_629,In_444);
and U1567 (N_1567,In_2334,N_1356);
nand U1568 (N_1568,N_1202,N_675);
xor U1569 (N_1569,N_1014,N_553);
nor U1570 (N_1570,N_756,N_1218);
and U1571 (N_1571,In_392,N_1370);
or U1572 (N_1572,N_846,N_816);
nor U1573 (N_1573,N_582,N_55);
nor U1574 (N_1574,In_908,In_25);
nand U1575 (N_1575,N_1244,In_603);
nor U1576 (N_1576,N_1004,N_1224);
and U1577 (N_1577,In_1240,N_783);
or U1578 (N_1578,In_74,N_1025);
or U1579 (N_1579,N_692,N_1392);
nor U1580 (N_1580,N_1179,In_1485);
nand U1581 (N_1581,N_1283,N_1063);
or U1582 (N_1582,N_1308,N_1463);
nand U1583 (N_1583,In_2018,N_1488);
nor U1584 (N_1584,N_1119,N_1415);
and U1585 (N_1585,N_1075,In_1489);
nor U1586 (N_1586,In_33,N_1402);
nor U1587 (N_1587,In_2255,N_1042);
or U1588 (N_1588,N_760,N_1299);
nor U1589 (N_1589,N_1233,N_1474);
and U1590 (N_1590,In_1599,N_1011);
and U1591 (N_1591,N_1070,In_814);
or U1592 (N_1592,N_857,N_1354);
and U1593 (N_1593,N_1193,N_1294);
and U1594 (N_1594,In_1615,N_1177);
and U1595 (N_1595,In_148,N_623);
nor U1596 (N_1596,N_775,N_108);
nand U1597 (N_1597,N_1143,In_2116);
nor U1598 (N_1598,In_2280,N_1240);
xor U1599 (N_1599,N_1116,N_1012);
nand U1600 (N_1600,N_1103,N_1288);
nand U1601 (N_1601,N_43,N_1237);
and U1602 (N_1602,N_1314,N_621);
nor U1603 (N_1603,In_2212,N_871);
or U1604 (N_1604,N_1167,In_2205);
and U1605 (N_1605,N_1164,In_2389);
and U1606 (N_1606,In_121,N_730);
nand U1607 (N_1607,N_1041,In_235);
nand U1608 (N_1608,In_744,N_964);
nand U1609 (N_1609,N_822,N_1317);
nand U1610 (N_1610,In_660,N_1405);
nand U1611 (N_1611,N_57,N_1462);
nor U1612 (N_1612,In_1216,N_1432);
nand U1613 (N_1613,N_1239,N_1124);
xor U1614 (N_1614,N_1351,N_905);
and U1615 (N_1615,N_1466,In_2303);
xnor U1616 (N_1616,In_1935,N_179);
or U1617 (N_1617,N_1161,N_679);
nand U1618 (N_1618,N_1449,N_1260);
or U1619 (N_1619,In_1573,N_897);
nand U1620 (N_1620,In_507,N_503);
nor U1621 (N_1621,N_1083,N_1343);
or U1622 (N_1622,In_14,N_779);
nor U1623 (N_1623,N_1067,N_198);
nor U1624 (N_1624,N_1438,In_566);
nor U1625 (N_1625,N_1121,N_572);
nor U1626 (N_1626,N_558,N_1324);
and U1627 (N_1627,N_1125,N_1022);
nor U1628 (N_1628,In_1892,N_1203);
nor U1629 (N_1629,N_1236,N_801);
xor U1630 (N_1630,N_1321,N_1278);
nand U1631 (N_1631,N_1217,In_1937);
nand U1632 (N_1632,In_958,N_631);
or U1633 (N_1633,N_1408,In_209);
and U1634 (N_1634,N_399,N_1157);
or U1635 (N_1635,N_527,N_1461);
nor U1636 (N_1636,In_1355,N_1243);
and U1637 (N_1637,In_2001,N_1238);
and U1638 (N_1638,N_1419,N_1247);
and U1639 (N_1639,N_1078,N_1122);
nor U1640 (N_1640,In_1448,N_1128);
xnor U1641 (N_1641,N_833,N_1468);
and U1642 (N_1642,In_1560,N_1158);
nand U1643 (N_1643,N_193,N_1417);
nor U1644 (N_1644,N_719,N_1170);
and U1645 (N_1645,N_1099,N_1338);
or U1646 (N_1646,In_906,N_1337);
nor U1647 (N_1647,In_1657,N_1152);
nand U1648 (N_1648,N_514,N_1266);
nor U1649 (N_1649,In_1922,N_939);
nor U1650 (N_1650,N_1256,N_979);
nor U1651 (N_1651,N_1453,N_1034);
or U1652 (N_1652,N_315,N_842);
or U1653 (N_1653,N_1286,N_1433);
nor U1654 (N_1654,N_611,In_110);
nand U1655 (N_1655,In_2362,N_1205);
nor U1656 (N_1656,N_541,In_2220);
and U1657 (N_1657,N_1389,N_1149);
nand U1658 (N_1658,N_1160,N_1084);
xor U1659 (N_1659,N_247,N_1333);
nand U1660 (N_1660,N_1465,N_1358);
nand U1661 (N_1661,N_780,N_1220);
and U1662 (N_1662,In_2243,N_1138);
nor U1663 (N_1663,N_985,In_1251);
nor U1664 (N_1664,N_1010,In_2278);
and U1665 (N_1665,N_1054,N_1498);
nand U1666 (N_1666,N_1126,N_1076);
nor U1667 (N_1667,N_859,N_408);
and U1668 (N_1668,In_1296,N_411);
nor U1669 (N_1669,N_1281,N_1020);
and U1670 (N_1670,N_975,N_1413);
nand U1671 (N_1671,N_1346,N_1082);
and U1672 (N_1672,In_785,N_1311);
nor U1673 (N_1673,N_648,N_1342);
and U1674 (N_1674,N_994,N_152);
or U1675 (N_1675,N_1307,In_1328);
xor U1676 (N_1676,In_2393,N_530);
nor U1677 (N_1677,N_35,N_741);
nor U1678 (N_1678,N_967,In_1470);
xnor U1679 (N_1679,In_1443,N_420);
nand U1680 (N_1680,N_1018,N_1410);
or U1681 (N_1681,N_1079,In_1160);
nor U1682 (N_1682,N_747,N_971);
and U1683 (N_1683,In_2169,N_62);
nor U1684 (N_1684,N_1457,N_1407);
and U1685 (N_1685,N_1426,N_1211);
nor U1686 (N_1686,In_891,N_1372);
or U1687 (N_1687,N_1245,N_941);
xor U1688 (N_1688,N_1345,N_274);
nand U1689 (N_1689,N_1398,N_1101);
nor U1690 (N_1690,N_1072,N_501);
nor U1691 (N_1691,In_2479,N_1480);
or U1692 (N_1692,N_497,N_1290);
xor U1693 (N_1693,In_894,N_766);
or U1694 (N_1694,N_1420,N_1216);
or U1695 (N_1695,N_1439,N_1492);
nand U1696 (N_1696,N_426,N_912);
xnor U1697 (N_1697,In_2340,N_1479);
nand U1698 (N_1698,N_1303,N_1366);
or U1699 (N_1699,N_269,N_1336);
nor U1700 (N_1700,N_413,N_667);
or U1701 (N_1701,N_1265,N_1362);
nor U1702 (N_1702,In_975,N_1077);
nand U1703 (N_1703,N_1327,In_2296);
or U1704 (N_1704,N_1309,N_1061);
or U1705 (N_1705,N_1431,N_117);
and U1706 (N_1706,N_1363,N_332);
and U1707 (N_1707,N_1044,N_698);
nor U1708 (N_1708,N_1183,N_560);
nor U1709 (N_1709,In_710,N_1031);
nand U1710 (N_1710,N_1150,In_612);
nor U1711 (N_1711,In_854,N_1268);
and U1712 (N_1712,N_875,N_1409);
and U1713 (N_1713,N_1201,N_761);
nor U1714 (N_1714,In_1245,In_1502);
nor U1715 (N_1715,N_1348,In_170);
and U1716 (N_1716,N_956,N_1108);
and U1717 (N_1717,In_2087,N_790);
nor U1718 (N_1718,N_704,N_643);
or U1719 (N_1719,N_1454,N_764);
and U1720 (N_1720,In_525,N_1154);
nor U1721 (N_1721,In_682,In_2419);
nand U1722 (N_1722,N_1206,N_1335);
nand U1723 (N_1723,N_1310,N_1055);
or U1724 (N_1724,In_667,N_1400);
and U1725 (N_1725,N_1359,N_1325);
and U1726 (N_1726,N_1291,N_1339);
nor U1727 (N_1727,N_1147,In_1510);
xor U1728 (N_1728,N_1428,N_1250);
xor U1729 (N_1729,N_710,N_136);
nand U1730 (N_1730,N_121,N_1445);
nand U1731 (N_1731,N_1496,N_1030);
and U1732 (N_1732,In_1475,N_1251);
nand U1733 (N_1733,In_1988,N_1257);
and U1734 (N_1734,N_1455,N_1208);
nor U1735 (N_1735,N_1168,In_729);
or U1736 (N_1736,N_1440,In_2153);
and U1737 (N_1737,N_1185,N_1478);
xor U1738 (N_1738,In_1723,N_1484);
nor U1739 (N_1739,N_960,N_75);
xnor U1740 (N_1740,In_781,In_2055);
nor U1741 (N_1741,N_212,N_1422);
and U1742 (N_1742,In_1126,N_1200);
and U1743 (N_1743,N_1258,N_6);
nor U1744 (N_1744,In_2476,N_380);
nor U1745 (N_1745,N_1329,N_1102);
nand U1746 (N_1746,In_1301,In_2460);
and U1747 (N_1747,N_312,In_222);
nand U1748 (N_1748,N_858,N_1016);
xor U1749 (N_1749,N_1285,N_1017);
xnor U1750 (N_1750,N_1047,In_2420);
nand U1751 (N_1751,N_877,In_806);
nand U1752 (N_1752,N_1190,In_2433);
or U1753 (N_1753,N_1040,N_1412);
nand U1754 (N_1754,N_364,N_1493);
nand U1755 (N_1755,N_972,N_1277);
xor U1756 (N_1756,N_113,In_1380);
nor U1757 (N_1757,N_781,N_830);
and U1758 (N_1758,In_749,N_1068);
or U1759 (N_1759,N_1424,N_1316);
and U1760 (N_1760,N_1027,In_493);
and U1761 (N_1761,N_1127,N_976);
and U1762 (N_1762,N_1297,In_1327);
or U1763 (N_1763,N_1141,In_795);
nand U1764 (N_1764,N_787,In_1198);
xnor U1765 (N_1765,N_1252,N_946);
nor U1766 (N_1766,In_2201,In_447);
or U1767 (N_1767,N_894,N_1352);
nor U1768 (N_1768,In_568,N_637);
and U1769 (N_1769,N_1430,N_1353);
or U1770 (N_1770,N_1436,N_330);
or U1771 (N_1771,N_1048,N_697);
nand U1772 (N_1772,N_893,In_674);
xnor U1773 (N_1773,In_1267,N_1112);
nor U1774 (N_1774,N_487,N_1322);
and U1775 (N_1775,N_51,In_417);
and U1776 (N_1776,N_1139,N_1458);
and U1777 (N_1777,In_1348,N_1385);
nor U1778 (N_1778,N_1374,N_1153);
or U1779 (N_1779,In_931,N_1123);
nor U1780 (N_1780,N_668,N_1038);
and U1781 (N_1781,N_343,N_1305);
and U1782 (N_1782,N_1471,N_316);
or U1783 (N_1783,N_928,N_1181);
or U1784 (N_1784,N_980,N_1225);
nand U1785 (N_1785,N_418,In_53);
nand U1786 (N_1786,N_559,In_1578);
or U1787 (N_1787,In_817,N_1007);
and U1788 (N_1788,N_1397,N_1071);
nor U1789 (N_1789,N_1223,In_881);
and U1790 (N_1790,N_1401,In_545);
nand U1791 (N_1791,N_633,In_1487);
or U1792 (N_1792,N_1191,N_1395);
or U1793 (N_1793,N_1226,N_549);
and U1794 (N_1794,In_701,N_1489);
and U1795 (N_1795,In_103,N_1246);
nand U1796 (N_1796,N_574,N_1046);
nand U1797 (N_1797,In_1508,N_118);
nand U1798 (N_1798,N_1132,In_443);
or U1799 (N_1799,In_625,N_1375);
nand U1800 (N_1800,N_1024,N_1032);
nor U1801 (N_1801,N_1212,N_1118);
or U1802 (N_1802,In_1180,In_1444);
nand U1803 (N_1803,In_516,N_1215);
xnor U1804 (N_1804,N_386,N_1035);
nor U1805 (N_1805,In_161,N_271);
xnor U1806 (N_1806,N_1272,N_1151);
xor U1807 (N_1807,N_1276,In_557);
and U1808 (N_1808,N_1263,N_1490);
or U1809 (N_1809,N_1221,In_1177);
nand U1810 (N_1810,In_1321,N_1106);
or U1811 (N_1811,N_132,N_1098);
or U1812 (N_1812,N_1086,N_1051);
and U1813 (N_1813,In_1917,In_693);
and U1814 (N_1814,N_1131,N_178);
or U1815 (N_1815,N_1028,N_1056);
or U1816 (N_1816,N_1039,N_1388);
and U1817 (N_1817,N_896,In_959);
and U1818 (N_1818,In_657,In_2474);
nand U1819 (N_1819,N_854,In_1490);
nor U1820 (N_1820,N_1050,N_30);
or U1821 (N_1821,N_1002,N_663);
or U1822 (N_1822,In_1018,In_1927);
nor U1823 (N_1823,In_736,N_1271);
and U1824 (N_1824,In_1016,In_523);
and U1825 (N_1825,N_92,N_1391);
nand U1826 (N_1826,N_1222,N_1282);
nor U1827 (N_1827,In_684,N_1451);
and U1828 (N_1828,In_928,In_2182);
nand U1829 (N_1829,N_1350,N_1198);
and U1830 (N_1830,N_1341,N_353);
or U1831 (N_1831,N_1006,N_835);
or U1832 (N_1832,In_427,N_1015);
nor U1833 (N_1833,N_1472,In_1698);
or U1834 (N_1834,N_110,N_1090);
nand U1835 (N_1835,In_250,N_1213);
nand U1836 (N_1836,N_1052,N_1406);
or U1837 (N_1837,In_899,In_498);
or U1838 (N_1838,N_1133,N_1043);
nor U1839 (N_1839,N_1379,N_1254);
nand U1840 (N_1840,In_416,N_1384);
xor U1841 (N_1841,N_1499,N_1361);
and U1842 (N_1842,N_1393,In_964);
nor U1843 (N_1843,N_1060,In_825);
and U1844 (N_1844,N_1023,In_1986);
xnor U1845 (N_1845,In_1311,N_1442);
or U1846 (N_1846,N_1289,N_1195);
and U1847 (N_1847,N_1196,N_1315);
and U1848 (N_1848,In_354,In_2127);
xnor U1849 (N_1849,N_1057,N_1323);
nor U1850 (N_1850,N_1104,N_1241);
or U1851 (N_1851,In_1520,N_1270);
and U1852 (N_1852,In_2107,N_1298);
nor U1853 (N_1853,In_424,N_1008);
nor U1854 (N_1854,In_136,N_1473);
nor U1855 (N_1855,N_1095,N_733);
or U1856 (N_1856,In_2021,N_601);
or U1857 (N_1857,N_1094,N_1188);
or U1858 (N_1858,N_1437,N_1378);
or U1859 (N_1859,N_1287,N_953);
nand U1860 (N_1860,N_1355,N_1111);
nor U1861 (N_1861,N_1467,N_1231);
and U1862 (N_1862,N_520,In_82);
nor U1863 (N_1863,In_1446,In_1952);
or U1864 (N_1864,In_137,In_1827);
and U1865 (N_1865,In_296,N_1165);
or U1866 (N_1866,In_1866,In_1159);
nor U1867 (N_1867,N_109,N_1144);
or U1868 (N_1868,N_1275,N_1066);
and U1869 (N_1869,N_531,N_1460);
nand U1870 (N_1870,In_1844,N_778);
nand U1871 (N_1871,N_1135,In_2236);
or U1872 (N_1872,N_711,N_1418);
nand U1873 (N_1873,N_997,N_234);
or U1874 (N_1874,N_1146,N_485);
nor U1875 (N_1875,In_502,N_71);
nand U1876 (N_1876,In_938,N_607);
or U1877 (N_1877,In_2060,N_270);
nor U1878 (N_1878,N_968,In_2035);
and U1879 (N_1879,In_280,N_1049);
or U1880 (N_1880,N_1334,In_2463);
or U1881 (N_1881,N_492,N_296);
nand U1882 (N_1882,N_1162,N_1136);
or U1883 (N_1883,N_506,N_368);
nand U1884 (N_1884,N_1175,N_450);
nor U1885 (N_1885,N_1497,N_1368);
xor U1886 (N_1886,In_1351,N_1228);
nand U1887 (N_1887,N_1320,N_827);
or U1888 (N_1888,N_1259,N_268);
and U1889 (N_1889,N_1069,N_838);
and U1890 (N_1890,In_731,N_1481);
xor U1891 (N_1891,N_727,N_220);
xor U1892 (N_1892,N_84,In_1436);
nand U1893 (N_1893,N_1367,N_1159);
and U1894 (N_1894,In_2181,In_44);
nor U1895 (N_1895,N_983,In_240);
nand U1896 (N_1896,N_1295,N_1296);
nand U1897 (N_1897,N_738,In_953);
nand U1898 (N_1898,N_1089,In_2378);
and U1899 (N_1899,N_87,In_663);
or U1900 (N_1900,N_1156,N_1194);
or U1901 (N_1901,N_1447,N_1456);
nor U1902 (N_1902,In_1437,N_561);
nor U1903 (N_1903,In_2445,N_1214);
nor U1904 (N_1904,N_1021,N_563);
and U1905 (N_1905,N_414,N_1117);
xor U1906 (N_1906,N_1142,N_1113);
nor U1907 (N_1907,N_1255,N_1169);
or U1908 (N_1908,N_862,N_843);
or U1909 (N_1909,N_224,N_630);
nor U1910 (N_1910,N_1230,In_1202);
nand U1911 (N_1911,N_1486,N_1234);
nand U1912 (N_1912,In_2149,N_1115);
nand U1913 (N_1913,In_433,N_638);
nor U1914 (N_1914,N_1100,N_1045);
nor U1915 (N_1915,In_2492,N_1423);
nand U1916 (N_1916,N_886,N_1376);
or U1917 (N_1917,N_1421,N_640);
and U1918 (N_1918,N_1469,N_1331);
or U1919 (N_1919,N_1137,N_555);
xnor U1920 (N_1920,In_1405,N_1180);
or U1921 (N_1921,N_1404,N_1105);
or U1922 (N_1922,N_1148,N_1000);
and U1923 (N_1923,N_568,N_1187);
and U1924 (N_1924,N_903,N_1386);
or U1925 (N_1925,N_1434,N_1003);
or U1926 (N_1926,N_1450,N_571);
and U1927 (N_1927,N_1248,In_1716);
or U1928 (N_1928,N_1347,In_939);
nor U1929 (N_1929,N_244,In_1285);
or U1930 (N_1930,N_1429,N_1173);
or U1931 (N_1931,N_1009,N_1064);
xnor U1932 (N_1932,In_2424,N_1494);
nand U1933 (N_1933,N_349,In_1082);
and U1934 (N_1934,N_681,N_1300);
nand U1935 (N_1935,N_594,In_645);
or U1936 (N_1936,In_1033,N_1448);
nor U1937 (N_1937,In_454,N_1130);
or U1938 (N_1938,N_1166,N_424);
nand U1939 (N_1939,N_1459,In_1237);
and U1940 (N_1940,N_255,N_1085);
nor U1941 (N_1941,In_1653,N_1091);
nor U1942 (N_1942,N_1414,N_1387);
nor U1943 (N_1943,N_1026,N_1235);
nand U1944 (N_1944,In_639,N_1081);
nor U1945 (N_1945,N_1242,In_1388);
nor U1946 (N_1946,In_563,In_269);
or U1947 (N_1947,N_291,N_1312);
or U1948 (N_1948,N_223,In_961);
xor U1949 (N_1949,In_760,N_1292);
or U1950 (N_1950,In_717,N_1452);
nor U1951 (N_1951,In_377,N_1107);
nand U1952 (N_1952,N_1435,N_1273);
xnor U1953 (N_1953,N_4,In_2295);
or U1954 (N_1954,N_1330,N_1364);
or U1955 (N_1955,N_606,N_1001);
or U1956 (N_1956,N_1155,N_1411);
or U1957 (N_1957,N_536,N_1396);
nand U1958 (N_1958,N_1390,In_119);
nor U1959 (N_1959,N_686,In_644);
nand U1960 (N_1960,N_1279,N_1114);
nand U1961 (N_1961,In_1635,N_1145);
nor U1962 (N_1962,N_1036,In_676);
and U1963 (N_1963,N_1262,N_85);
or U1964 (N_1964,In_1320,N_171);
and U1965 (N_1965,N_826,In_13);
nor U1966 (N_1966,N_1186,N_1065);
and U1967 (N_1967,N_1319,In_2122);
and U1968 (N_1968,N_1059,N_545);
xor U1969 (N_1969,N_1425,N_1382);
xor U1970 (N_1970,N_1207,In_723);
nand U1971 (N_1971,In_384,N_1383);
nand U1972 (N_1972,N_1062,N_919);
or U1973 (N_1973,In_1807,N_1209);
and U1974 (N_1974,N_1087,N_1080);
and U1975 (N_1975,N_1073,In_2467);
nor U1976 (N_1976,In_987,N_1219);
or U1977 (N_1977,N_1053,In_87);
xor U1978 (N_1978,N_744,N_557);
nor U1979 (N_1979,In_816,N_1253);
or U1980 (N_1980,N_1178,In_826);
or U1981 (N_1981,In_154,N_929);
nor U1982 (N_1982,In_337,N_932);
nand U1983 (N_1983,N_1371,N_333);
and U1984 (N_1984,N_1482,In_1048);
nor U1985 (N_1985,N_542,N_828);
xor U1986 (N_1986,In_406,N_923);
nor U1987 (N_1987,In_2263,In_1447);
and U1988 (N_1988,N_1377,N_1019);
xor U1989 (N_1989,N_229,In_2382);
and U1990 (N_1990,N_1184,N_139);
nand U1991 (N_1991,N_1120,N_1293);
or U1992 (N_1992,N_504,N_510);
xnor U1993 (N_1993,N_852,N_1096);
nand U1994 (N_1994,N_991,N_1349);
nand U1995 (N_1995,In_1539,N_874);
or U1996 (N_1996,N_1427,N_1176);
nor U1997 (N_1997,In_2348,N_227);
and U1998 (N_1998,N_732,N_1369);
nor U1999 (N_1999,In_1368,In_1667);
nand U2000 (N_2000,N_1650,N_1586);
or U2001 (N_2001,N_1868,N_1700);
and U2002 (N_2002,N_1720,N_1929);
nor U2003 (N_2003,N_1948,N_1511);
and U2004 (N_2004,N_1734,N_1595);
nor U2005 (N_2005,N_1900,N_1596);
or U2006 (N_2006,N_1616,N_1551);
nor U2007 (N_2007,N_1764,N_1600);
xnor U2008 (N_2008,N_1591,N_1837);
and U2009 (N_2009,N_1906,N_1961);
and U2010 (N_2010,N_1791,N_1537);
nor U2011 (N_2011,N_1944,N_1880);
nor U2012 (N_2012,N_1725,N_1621);
nor U2013 (N_2013,N_1699,N_1573);
nor U2014 (N_2014,N_1937,N_1631);
nand U2015 (N_2015,N_1803,N_1854);
or U2016 (N_2016,N_1793,N_1506);
nor U2017 (N_2017,N_1902,N_1851);
nand U2018 (N_2018,N_1715,N_1896);
and U2019 (N_2019,N_1912,N_1986);
nand U2020 (N_2020,N_1608,N_1624);
and U2021 (N_2021,N_1761,N_1992);
or U2022 (N_2022,N_1776,N_1863);
and U2023 (N_2023,N_1972,N_1669);
and U2024 (N_2024,N_1812,N_1686);
and U2025 (N_2025,N_1566,N_1982);
nor U2026 (N_2026,N_1947,N_1641);
nor U2027 (N_2027,N_1640,N_1694);
nand U2028 (N_2028,N_1876,N_1701);
nor U2029 (N_2029,N_1781,N_1664);
and U2030 (N_2030,N_1999,N_1894);
nor U2031 (N_2031,N_1996,N_1557);
nor U2032 (N_2032,N_1878,N_1530);
nor U2033 (N_2033,N_1866,N_1717);
xor U2034 (N_2034,N_1558,N_1702);
and U2035 (N_2035,N_1800,N_1731);
nand U2036 (N_2036,N_1960,N_1535);
nor U2037 (N_2037,N_1517,N_1716);
nand U2038 (N_2038,N_1954,N_1626);
nor U2039 (N_2039,N_1553,N_1941);
nor U2040 (N_2040,N_1648,N_1974);
nand U2041 (N_2041,N_1763,N_1835);
or U2042 (N_2042,N_1963,N_1849);
nor U2043 (N_2043,N_1684,N_1625);
and U2044 (N_2044,N_1945,N_1698);
nor U2045 (N_2045,N_1501,N_1507);
and U2046 (N_2046,N_1922,N_1886);
nor U2047 (N_2047,N_1949,N_1636);
or U2048 (N_2048,N_1555,N_1713);
and U2049 (N_2049,N_1615,N_1879);
xnor U2050 (N_2050,N_1955,N_1799);
nand U2051 (N_2051,N_1512,N_1674);
nand U2052 (N_2052,N_1749,N_1989);
and U2053 (N_2053,N_1897,N_1677);
and U2054 (N_2054,N_1516,N_1829);
and U2055 (N_2055,N_1521,N_1842);
nand U2056 (N_2056,N_1697,N_1620);
nor U2057 (N_2057,N_1518,N_1790);
nand U2058 (N_2058,N_1861,N_1565);
or U2059 (N_2059,N_1690,N_1743);
xnor U2060 (N_2060,N_1827,N_1617);
and U2061 (N_2061,N_1561,N_1578);
or U2062 (N_2062,N_1576,N_1718);
or U2063 (N_2063,N_1593,N_1884);
nand U2064 (N_2064,N_1704,N_1735);
and U2065 (N_2065,N_1695,N_1783);
or U2066 (N_2066,N_1574,N_1809);
or U2067 (N_2067,N_1659,N_1895);
and U2068 (N_2068,N_1634,N_1738);
or U2069 (N_2069,N_1838,N_1856);
nand U2070 (N_2070,N_1752,N_1582);
nor U2071 (N_2071,N_1782,N_1755);
and U2072 (N_2072,N_1872,N_1795);
xnor U2073 (N_2073,N_1644,N_1592);
xor U2074 (N_2074,N_1924,N_1811);
nor U2075 (N_2075,N_1657,N_1509);
or U2076 (N_2076,N_1881,N_1639);
nand U2077 (N_2077,N_1911,N_1770);
nor U2078 (N_2078,N_1691,N_1768);
or U2079 (N_2079,N_1550,N_1970);
and U2080 (N_2080,N_1587,N_1719);
nor U2081 (N_2081,N_1899,N_1769);
and U2082 (N_2082,N_1660,N_1870);
xnor U2083 (N_2083,N_1540,N_1789);
nor U2084 (N_2084,N_1532,N_1662);
nand U2085 (N_2085,N_1693,N_1977);
nand U2086 (N_2086,N_1794,N_1831);
nand U2087 (N_2087,N_1729,N_1796);
nand U2088 (N_2088,N_1844,N_1687);
nand U2089 (N_2089,N_1773,N_1936);
nor U2090 (N_2090,N_1806,N_1602);
nor U2091 (N_2091,N_1556,N_1885);
nor U2092 (N_2092,N_1584,N_1500);
nand U2093 (N_2093,N_1520,N_1546);
nand U2094 (N_2094,N_1871,N_1552);
nor U2095 (N_2095,N_1746,N_1820);
xor U2096 (N_2096,N_1708,N_1741);
and U2097 (N_2097,N_1765,N_1685);
or U2098 (N_2098,N_1706,N_1762);
nor U2099 (N_2099,N_1601,N_1824);
xor U2100 (N_2100,N_1751,N_1819);
or U2101 (N_2101,N_1581,N_1607);
nand U2102 (N_2102,N_1721,N_1926);
nand U2103 (N_2103,N_1562,N_1938);
or U2104 (N_2104,N_1850,N_1801);
nand U2105 (N_2105,N_1575,N_1672);
nand U2106 (N_2106,N_1547,N_1767);
and U2107 (N_2107,N_1877,N_1671);
and U2108 (N_2108,N_1745,N_1610);
xnor U2109 (N_2109,N_1932,N_1737);
nor U2110 (N_2110,N_1888,N_1971);
nand U2111 (N_2111,N_1920,N_1663);
and U2112 (N_2112,N_1930,N_1661);
and U2113 (N_2113,N_1942,N_1676);
and U2114 (N_2114,N_1559,N_1654);
nor U2115 (N_2115,N_1946,N_1524);
nor U2116 (N_2116,N_1632,N_1703);
xor U2117 (N_2117,N_1712,N_1748);
or U2118 (N_2118,N_1709,N_1689);
and U2119 (N_2119,N_1679,N_1688);
xor U2120 (N_2120,N_1774,N_1825);
and U2121 (N_2121,N_1612,N_1798);
nand U2122 (N_2122,N_1822,N_1728);
and U2123 (N_2123,N_1655,N_1536);
and U2124 (N_2124,N_1554,N_1785);
nor U2125 (N_2125,N_1980,N_1523);
nor U2126 (N_2126,N_1533,N_1991);
and U2127 (N_2127,N_1505,N_1780);
and U2128 (N_2128,N_1777,N_1613);
or U2129 (N_2129,N_1904,N_1784);
nand U2130 (N_2130,N_1993,N_1665);
nor U2131 (N_2131,N_1513,N_1867);
or U2132 (N_2132,N_1858,N_1990);
xnor U2133 (N_2133,N_1652,N_1771);
nor U2134 (N_2134,N_1840,N_1653);
nor U2135 (N_2135,N_1692,N_1987);
or U2136 (N_2136,N_1673,N_1649);
nand U2137 (N_2137,N_1571,N_1696);
or U2138 (N_2138,N_1915,N_1935);
and U2139 (N_2139,N_1647,N_1808);
and U2140 (N_2140,N_1680,N_1514);
or U2141 (N_2141,N_1726,N_1622);
or U2142 (N_2142,N_1797,N_1710);
xnor U2143 (N_2143,N_1913,N_1964);
and U2144 (N_2144,N_1599,N_1775);
nor U2145 (N_2145,N_1848,N_1637);
nor U2146 (N_2146,N_1860,N_1853);
nor U2147 (N_2147,N_1564,N_1979);
nor U2148 (N_2148,N_1953,N_1570);
and U2149 (N_2149,N_1678,N_1508);
or U2150 (N_2150,N_1818,N_1943);
xnor U2151 (N_2151,N_1510,N_1502);
or U2152 (N_2152,N_1609,N_1759);
xor U2153 (N_2153,N_1847,N_1747);
nand U2154 (N_2154,N_1614,N_1569);
nor U2155 (N_2155,N_1543,N_1969);
and U2156 (N_2156,N_1957,N_1522);
nand U2157 (N_2157,N_1817,N_1869);
nand U2158 (N_2158,N_1905,N_1766);
and U2159 (N_2159,N_1670,N_1816);
nor U2160 (N_2160,N_1864,N_1628);
nand U2161 (N_2161,N_1638,N_1778);
or U2162 (N_2162,N_1925,N_1841);
and U2163 (N_2163,N_1952,N_1740);
nor U2164 (N_2164,N_1901,N_1968);
nand U2165 (N_2165,N_1604,N_1833);
nor U2166 (N_2166,N_1642,N_1927);
or U2167 (N_2167,N_1750,N_1830);
nor U2168 (N_2168,N_1722,N_1802);
nor U2169 (N_2169,N_1643,N_1732);
nor U2170 (N_2170,N_1959,N_1988);
and U2171 (N_2171,N_1939,N_1810);
nor U2172 (N_2172,N_1733,N_1619);
nor U2173 (N_2173,N_1984,N_1973);
and U2174 (N_2174,N_1723,N_1779);
nor U2175 (N_2175,N_1859,N_1668);
or U2176 (N_2176,N_1623,N_1966);
or U2177 (N_2177,N_1846,N_1635);
or U2178 (N_2178,N_1978,N_1792);
and U2179 (N_2179,N_1956,N_1529);
nand U2180 (N_2180,N_1525,N_1539);
and U2181 (N_2181,N_1589,N_1597);
nand U2182 (N_2182,N_1898,N_1645);
nor U2183 (N_2183,N_1940,N_1908);
and U2184 (N_2184,N_1588,N_1606);
nand U2185 (N_2185,N_1577,N_1629);
nand U2186 (N_2186,N_1627,N_1658);
nand U2187 (N_2187,N_1962,N_1909);
and U2188 (N_2188,N_1845,N_1923);
xnor U2189 (N_2189,N_1560,N_1843);
or U2190 (N_2190,N_1772,N_1931);
nor U2191 (N_2191,N_1756,N_1994);
and U2192 (N_2192,N_1528,N_1786);
and U2193 (N_2193,N_1882,N_1804);
nand U2194 (N_2194,N_1983,N_1891);
or U2195 (N_2195,N_1548,N_1744);
nor U2196 (N_2196,N_1997,N_1515);
and U2197 (N_2197,N_1857,N_1958);
and U2198 (N_2198,N_1646,N_1760);
and U2199 (N_2199,N_1545,N_1727);
or U2200 (N_2200,N_1807,N_1893);
and U2201 (N_2201,N_1757,N_1950);
nor U2202 (N_2202,N_1873,N_1742);
or U2203 (N_2203,N_1519,N_1585);
and U2204 (N_2204,N_1874,N_1736);
and U2205 (N_2205,N_1985,N_1633);
or U2206 (N_2206,N_1583,N_1503);
nor U2207 (N_2207,N_1865,N_1875);
or U2208 (N_2208,N_1730,N_1707);
or U2209 (N_2209,N_1714,N_1724);
or U2210 (N_2210,N_1531,N_1666);
xnor U2211 (N_2211,N_1967,N_1618);
xor U2212 (N_2212,N_1568,N_1526);
or U2213 (N_2213,N_1951,N_1563);
nand U2214 (N_2214,N_1917,N_1981);
and U2215 (N_2215,N_1855,N_1527);
nand U2216 (N_2216,N_1889,N_1852);
or U2217 (N_2217,N_1921,N_1542);
and U2218 (N_2218,N_1828,N_1538);
or U2219 (N_2219,N_1976,N_1823);
or U2220 (N_2220,N_1928,N_1683);
nor U2221 (N_2221,N_1892,N_1836);
nand U2222 (N_2222,N_1998,N_1541);
nor U2223 (N_2223,N_1907,N_1656);
nand U2224 (N_2224,N_1682,N_1630);
and U2225 (N_2225,N_1903,N_1603);
or U2226 (N_2226,N_1534,N_1975);
or U2227 (N_2227,N_1890,N_1813);
and U2228 (N_2228,N_1590,N_1862);
and U2229 (N_2229,N_1651,N_1995);
and U2230 (N_2230,N_1544,N_1826);
and U2231 (N_2231,N_1675,N_1572);
or U2232 (N_2232,N_1933,N_1815);
nand U2233 (N_2233,N_1681,N_1934);
nor U2234 (N_2234,N_1910,N_1611);
nor U2235 (N_2235,N_1834,N_1594);
nand U2236 (N_2236,N_1504,N_1883);
and U2237 (N_2237,N_1821,N_1605);
and U2238 (N_2238,N_1598,N_1567);
nand U2239 (N_2239,N_1839,N_1753);
or U2240 (N_2240,N_1739,N_1667);
nor U2241 (N_2241,N_1758,N_1805);
nand U2242 (N_2242,N_1787,N_1918);
xnor U2243 (N_2243,N_1887,N_1549);
and U2244 (N_2244,N_1916,N_1580);
or U2245 (N_2245,N_1754,N_1711);
nor U2246 (N_2246,N_1919,N_1579);
xnor U2247 (N_2247,N_1705,N_1914);
nand U2248 (N_2248,N_1788,N_1814);
xor U2249 (N_2249,N_1965,N_1832);
and U2250 (N_2250,N_1904,N_1901);
xnor U2251 (N_2251,N_1696,N_1714);
or U2252 (N_2252,N_1943,N_1598);
and U2253 (N_2253,N_1679,N_1802);
nor U2254 (N_2254,N_1537,N_1999);
nand U2255 (N_2255,N_1734,N_1834);
nand U2256 (N_2256,N_1826,N_1641);
nand U2257 (N_2257,N_1598,N_1580);
or U2258 (N_2258,N_1651,N_1771);
or U2259 (N_2259,N_1964,N_1785);
nor U2260 (N_2260,N_1720,N_1790);
or U2261 (N_2261,N_1992,N_1608);
and U2262 (N_2262,N_1544,N_1709);
and U2263 (N_2263,N_1777,N_1935);
nor U2264 (N_2264,N_1824,N_1957);
or U2265 (N_2265,N_1852,N_1626);
and U2266 (N_2266,N_1554,N_1786);
or U2267 (N_2267,N_1924,N_1790);
or U2268 (N_2268,N_1502,N_1816);
nand U2269 (N_2269,N_1971,N_1517);
and U2270 (N_2270,N_1742,N_1850);
nand U2271 (N_2271,N_1545,N_1698);
xor U2272 (N_2272,N_1892,N_1569);
or U2273 (N_2273,N_1559,N_1652);
nor U2274 (N_2274,N_1730,N_1968);
or U2275 (N_2275,N_1875,N_1588);
nor U2276 (N_2276,N_1976,N_1975);
and U2277 (N_2277,N_1630,N_1912);
nor U2278 (N_2278,N_1734,N_1592);
or U2279 (N_2279,N_1819,N_1574);
and U2280 (N_2280,N_1774,N_1563);
or U2281 (N_2281,N_1627,N_1803);
nor U2282 (N_2282,N_1841,N_1725);
nor U2283 (N_2283,N_1776,N_1960);
nor U2284 (N_2284,N_1929,N_1969);
or U2285 (N_2285,N_1993,N_1868);
nand U2286 (N_2286,N_1654,N_1530);
nor U2287 (N_2287,N_1591,N_1804);
and U2288 (N_2288,N_1983,N_1794);
nor U2289 (N_2289,N_1856,N_1671);
and U2290 (N_2290,N_1571,N_1702);
nor U2291 (N_2291,N_1899,N_1912);
nor U2292 (N_2292,N_1618,N_1859);
nor U2293 (N_2293,N_1958,N_1783);
and U2294 (N_2294,N_1615,N_1725);
or U2295 (N_2295,N_1612,N_1614);
and U2296 (N_2296,N_1590,N_1725);
nor U2297 (N_2297,N_1903,N_1563);
nor U2298 (N_2298,N_1973,N_1820);
nand U2299 (N_2299,N_1921,N_1721);
or U2300 (N_2300,N_1782,N_1995);
xnor U2301 (N_2301,N_1580,N_1573);
or U2302 (N_2302,N_1810,N_1882);
nand U2303 (N_2303,N_1997,N_1788);
nor U2304 (N_2304,N_1840,N_1610);
and U2305 (N_2305,N_1574,N_1784);
nand U2306 (N_2306,N_1953,N_1916);
nand U2307 (N_2307,N_1682,N_1529);
nand U2308 (N_2308,N_1900,N_1811);
or U2309 (N_2309,N_1650,N_1577);
nand U2310 (N_2310,N_1773,N_1891);
nand U2311 (N_2311,N_1599,N_1696);
nand U2312 (N_2312,N_1835,N_1597);
nor U2313 (N_2313,N_1946,N_1843);
nand U2314 (N_2314,N_1969,N_1724);
nand U2315 (N_2315,N_1704,N_1685);
or U2316 (N_2316,N_1577,N_1511);
xnor U2317 (N_2317,N_1694,N_1850);
xor U2318 (N_2318,N_1524,N_1890);
and U2319 (N_2319,N_1538,N_1577);
nor U2320 (N_2320,N_1706,N_1896);
nand U2321 (N_2321,N_1743,N_1941);
nor U2322 (N_2322,N_1534,N_1997);
nand U2323 (N_2323,N_1975,N_1939);
nand U2324 (N_2324,N_1664,N_1685);
nor U2325 (N_2325,N_1865,N_1814);
nand U2326 (N_2326,N_1848,N_1688);
or U2327 (N_2327,N_1993,N_1823);
nand U2328 (N_2328,N_1593,N_1932);
or U2329 (N_2329,N_1665,N_1961);
or U2330 (N_2330,N_1655,N_1794);
nand U2331 (N_2331,N_1505,N_1809);
or U2332 (N_2332,N_1752,N_1834);
nor U2333 (N_2333,N_1974,N_1955);
and U2334 (N_2334,N_1804,N_1568);
or U2335 (N_2335,N_1807,N_1623);
nand U2336 (N_2336,N_1799,N_1506);
nor U2337 (N_2337,N_1981,N_1588);
nand U2338 (N_2338,N_1581,N_1745);
and U2339 (N_2339,N_1869,N_1907);
nand U2340 (N_2340,N_1689,N_1536);
and U2341 (N_2341,N_1519,N_1641);
nor U2342 (N_2342,N_1586,N_1786);
and U2343 (N_2343,N_1811,N_1779);
nor U2344 (N_2344,N_1897,N_1807);
nand U2345 (N_2345,N_1697,N_1769);
nor U2346 (N_2346,N_1784,N_1979);
nor U2347 (N_2347,N_1780,N_1763);
or U2348 (N_2348,N_1630,N_1803);
nand U2349 (N_2349,N_1985,N_1714);
nor U2350 (N_2350,N_1698,N_1958);
and U2351 (N_2351,N_1505,N_1775);
nand U2352 (N_2352,N_1570,N_1554);
or U2353 (N_2353,N_1769,N_1859);
nor U2354 (N_2354,N_1574,N_1559);
nand U2355 (N_2355,N_1989,N_1502);
nand U2356 (N_2356,N_1989,N_1637);
nand U2357 (N_2357,N_1684,N_1806);
nand U2358 (N_2358,N_1552,N_1799);
or U2359 (N_2359,N_1659,N_1666);
or U2360 (N_2360,N_1686,N_1648);
and U2361 (N_2361,N_1958,N_1664);
or U2362 (N_2362,N_1742,N_1731);
xor U2363 (N_2363,N_1594,N_1685);
nor U2364 (N_2364,N_1814,N_1690);
or U2365 (N_2365,N_1791,N_1566);
nand U2366 (N_2366,N_1957,N_1563);
nand U2367 (N_2367,N_1722,N_1944);
and U2368 (N_2368,N_1660,N_1924);
nor U2369 (N_2369,N_1998,N_1604);
or U2370 (N_2370,N_1877,N_1555);
and U2371 (N_2371,N_1835,N_1667);
and U2372 (N_2372,N_1892,N_1609);
and U2373 (N_2373,N_1803,N_1788);
or U2374 (N_2374,N_1649,N_1645);
nand U2375 (N_2375,N_1796,N_1978);
or U2376 (N_2376,N_1726,N_1793);
nand U2377 (N_2377,N_1965,N_1559);
nor U2378 (N_2378,N_1843,N_1671);
or U2379 (N_2379,N_1530,N_1600);
nor U2380 (N_2380,N_1690,N_1945);
nor U2381 (N_2381,N_1685,N_1538);
nand U2382 (N_2382,N_1646,N_1635);
or U2383 (N_2383,N_1764,N_1578);
or U2384 (N_2384,N_1670,N_1989);
or U2385 (N_2385,N_1965,N_1783);
and U2386 (N_2386,N_1779,N_1804);
nand U2387 (N_2387,N_1618,N_1950);
nor U2388 (N_2388,N_1538,N_1594);
or U2389 (N_2389,N_1588,N_1696);
xor U2390 (N_2390,N_1552,N_1618);
nand U2391 (N_2391,N_1951,N_1605);
xnor U2392 (N_2392,N_1694,N_1530);
or U2393 (N_2393,N_1963,N_1513);
nor U2394 (N_2394,N_1843,N_1913);
or U2395 (N_2395,N_1777,N_1582);
nand U2396 (N_2396,N_1532,N_1822);
or U2397 (N_2397,N_1697,N_1589);
or U2398 (N_2398,N_1818,N_1596);
and U2399 (N_2399,N_1951,N_1717);
nor U2400 (N_2400,N_1917,N_1647);
nor U2401 (N_2401,N_1811,N_1694);
and U2402 (N_2402,N_1685,N_1847);
nand U2403 (N_2403,N_1654,N_1799);
and U2404 (N_2404,N_1997,N_1507);
nor U2405 (N_2405,N_1894,N_1550);
nand U2406 (N_2406,N_1972,N_1890);
and U2407 (N_2407,N_1876,N_1979);
or U2408 (N_2408,N_1684,N_1722);
xor U2409 (N_2409,N_1662,N_1933);
or U2410 (N_2410,N_1885,N_1638);
and U2411 (N_2411,N_1640,N_1828);
nor U2412 (N_2412,N_1961,N_1681);
and U2413 (N_2413,N_1654,N_1811);
or U2414 (N_2414,N_1560,N_1845);
or U2415 (N_2415,N_1672,N_1971);
xnor U2416 (N_2416,N_1545,N_1661);
nand U2417 (N_2417,N_1526,N_1626);
nor U2418 (N_2418,N_1799,N_1850);
nor U2419 (N_2419,N_1581,N_1767);
nand U2420 (N_2420,N_1516,N_1734);
nor U2421 (N_2421,N_1990,N_1847);
xor U2422 (N_2422,N_1740,N_1566);
or U2423 (N_2423,N_1505,N_1509);
nand U2424 (N_2424,N_1993,N_1597);
and U2425 (N_2425,N_1509,N_1532);
or U2426 (N_2426,N_1815,N_1878);
nor U2427 (N_2427,N_1889,N_1705);
nor U2428 (N_2428,N_1762,N_1942);
xnor U2429 (N_2429,N_1669,N_1808);
nor U2430 (N_2430,N_1601,N_1795);
nand U2431 (N_2431,N_1875,N_1502);
and U2432 (N_2432,N_1862,N_1536);
xor U2433 (N_2433,N_1900,N_1687);
nand U2434 (N_2434,N_1597,N_1621);
nand U2435 (N_2435,N_1580,N_1821);
or U2436 (N_2436,N_1973,N_1647);
xor U2437 (N_2437,N_1882,N_1815);
nand U2438 (N_2438,N_1684,N_1819);
and U2439 (N_2439,N_1540,N_1994);
and U2440 (N_2440,N_1837,N_1895);
or U2441 (N_2441,N_1982,N_1955);
nand U2442 (N_2442,N_1715,N_1839);
nor U2443 (N_2443,N_1984,N_1619);
or U2444 (N_2444,N_1701,N_1639);
xnor U2445 (N_2445,N_1899,N_1666);
and U2446 (N_2446,N_1744,N_1538);
nand U2447 (N_2447,N_1644,N_1634);
and U2448 (N_2448,N_1707,N_1901);
or U2449 (N_2449,N_1942,N_1644);
nor U2450 (N_2450,N_1982,N_1788);
nand U2451 (N_2451,N_1566,N_1521);
and U2452 (N_2452,N_1643,N_1960);
or U2453 (N_2453,N_1843,N_1630);
and U2454 (N_2454,N_1931,N_1935);
nand U2455 (N_2455,N_1844,N_1905);
or U2456 (N_2456,N_1813,N_1931);
and U2457 (N_2457,N_1564,N_1759);
nor U2458 (N_2458,N_1674,N_1883);
nand U2459 (N_2459,N_1579,N_1620);
nand U2460 (N_2460,N_1713,N_1894);
and U2461 (N_2461,N_1610,N_1751);
nand U2462 (N_2462,N_1729,N_1990);
or U2463 (N_2463,N_1892,N_1751);
xnor U2464 (N_2464,N_1958,N_1992);
and U2465 (N_2465,N_1767,N_1805);
nand U2466 (N_2466,N_1627,N_1818);
or U2467 (N_2467,N_1709,N_1672);
or U2468 (N_2468,N_1986,N_1784);
or U2469 (N_2469,N_1555,N_1742);
xnor U2470 (N_2470,N_1756,N_1730);
nand U2471 (N_2471,N_1536,N_1532);
nor U2472 (N_2472,N_1943,N_1908);
nor U2473 (N_2473,N_1742,N_1908);
or U2474 (N_2474,N_1715,N_1750);
xnor U2475 (N_2475,N_1520,N_1954);
and U2476 (N_2476,N_1682,N_1961);
nand U2477 (N_2477,N_1695,N_1820);
or U2478 (N_2478,N_1830,N_1856);
nor U2479 (N_2479,N_1982,N_1707);
nand U2480 (N_2480,N_1703,N_1966);
nand U2481 (N_2481,N_1896,N_1653);
or U2482 (N_2482,N_1923,N_1686);
nor U2483 (N_2483,N_1676,N_1683);
or U2484 (N_2484,N_1929,N_1892);
or U2485 (N_2485,N_1507,N_1796);
nand U2486 (N_2486,N_1568,N_1896);
and U2487 (N_2487,N_1560,N_1750);
and U2488 (N_2488,N_1979,N_1993);
nor U2489 (N_2489,N_1836,N_1873);
and U2490 (N_2490,N_1960,N_1880);
nor U2491 (N_2491,N_1874,N_1615);
nor U2492 (N_2492,N_1841,N_1583);
and U2493 (N_2493,N_1673,N_1707);
xnor U2494 (N_2494,N_1597,N_1940);
xnor U2495 (N_2495,N_1735,N_1594);
and U2496 (N_2496,N_1777,N_1611);
nor U2497 (N_2497,N_1951,N_1665);
or U2498 (N_2498,N_1867,N_1929);
nand U2499 (N_2499,N_1845,N_1891);
xor U2500 (N_2500,N_2111,N_2089);
or U2501 (N_2501,N_2131,N_2039);
and U2502 (N_2502,N_2276,N_2442);
and U2503 (N_2503,N_2412,N_2355);
nand U2504 (N_2504,N_2090,N_2108);
xnor U2505 (N_2505,N_2298,N_2058);
nor U2506 (N_2506,N_2386,N_2024);
nand U2507 (N_2507,N_2356,N_2289);
or U2508 (N_2508,N_2278,N_2093);
nand U2509 (N_2509,N_2489,N_2147);
xnor U2510 (N_2510,N_2311,N_2119);
and U2511 (N_2511,N_2008,N_2116);
nand U2512 (N_2512,N_2395,N_2344);
or U2513 (N_2513,N_2085,N_2308);
or U2514 (N_2514,N_2491,N_2018);
nor U2515 (N_2515,N_2127,N_2270);
and U2516 (N_2516,N_2142,N_2248);
nor U2517 (N_2517,N_2385,N_2316);
nand U2518 (N_2518,N_2079,N_2424);
xor U2519 (N_2519,N_2411,N_2397);
or U2520 (N_2520,N_2103,N_2241);
and U2521 (N_2521,N_2493,N_2138);
and U2522 (N_2522,N_2230,N_2307);
nor U2523 (N_2523,N_2281,N_2359);
or U2524 (N_2524,N_2244,N_2306);
nor U2525 (N_2525,N_2498,N_2291);
or U2526 (N_2526,N_2486,N_2026);
or U2527 (N_2527,N_2256,N_2333);
or U2528 (N_2528,N_2065,N_2321);
and U2529 (N_2529,N_2364,N_2312);
xor U2530 (N_2530,N_2201,N_2328);
or U2531 (N_2531,N_2099,N_2123);
nor U2532 (N_2532,N_2372,N_2151);
nand U2533 (N_2533,N_2141,N_2242);
or U2534 (N_2534,N_2438,N_2461);
nand U2535 (N_2535,N_2129,N_2071);
and U2536 (N_2536,N_2143,N_2433);
or U2537 (N_2537,N_2114,N_2014);
or U2538 (N_2538,N_2404,N_2408);
or U2539 (N_2539,N_2224,N_2113);
nand U2540 (N_2540,N_2189,N_2440);
nor U2541 (N_2541,N_2254,N_2346);
and U2542 (N_2542,N_2416,N_2013);
and U2543 (N_2543,N_2236,N_2221);
nor U2544 (N_2544,N_2112,N_2052);
nor U2545 (N_2545,N_2252,N_2032);
or U2546 (N_2546,N_2290,N_2341);
nand U2547 (N_2547,N_2219,N_2296);
and U2548 (N_2548,N_2294,N_2302);
and U2549 (N_2549,N_2020,N_2309);
and U2550 (N_2550,N_2492,N_2028);
nand U2551 (N_2551,N_2188,N_2177);
and U2552 (N_2552,N_2470,N_2063);
nand U2553 (N_2553,N_2334,N_2390);
xor U2554 (N_2554,N_2444,N_2484);
nor U2555 (N_2555,N_2250,N_2200);
nor U2556 (N_2556,N_2448,N_2184);
nand U2557 (N_2557,N_2207,N_2443);
nor U2558 (N_2558,N_2027,N_2050);
and U2559 (N_2559,N_2384,N_2365);
or U2560 (N_2560,N_2011,N_2391);
nor U2561 (N_2561,N_2418,N_2148);
and U2562 (N_2562,N_2451,N_2392);
xnor U2563 (N_2563,N_2406,N_2343);
nand U2564 (N_2564,N_2313,N_2042);
nand U2565 (N_2565,N_2399,N_2047);
or U2566 (N_2566,N_2432,N_2156);
nor U2567 (N_2567,N_2109,N_2358);
nor U2568 (N_2568,N_2351,N_2382);
or U2569 (N_2569,N_2387,N_2087);
nor U2570 (N_2570,N_2314,N_2354);
nand U2571 (N_2571,N_2429,N_2367);
or U2572 (N_2572,N_2213,N_2135);
and U2573 (N_2573,N_2191,N_2455);
nor U2574 (N_2574,N_2258,N_2231);
or U2575 (N_2575,N_2419,N_2240);
and U2576 (N_2576,N_2192,N_2454);
nor U2577 (N_2577,N_2490,N_2046);
and U2578 (N_2578,N_2379,N_2479);
nand U2579 (N_2579,N_2318,N_2245);
and U2580 (N_2580,N_2036,N_2423);
or U2581 (N_2581,N_2226,N_2457);
nand U2582 (N_2582,N_2260,N_2217);
nand U2583 (N_2583,N_2170,N_2209);
and U2584 (N_2584,N_2081,N_2082);
nand U2585 (N_2585,N_2465,N_2004);
nor U2586 (N_2586,N_2259,N_2257);
and U2587 (N_2587,N_2439,N_2169);
and U2588 (N_2588,N_2165,N_2060);
nand U2589 (N_2589,N_2202,N_2167);
nor U2590 (N_2590,N_2352,N_2292);
nand U2591 (N_2591,N_2273,N_2373);
nor U2592 (N_2592,N_2474,N_2105);
nor U2593 (N_2593,N_2064,N_2096);
nor U2594 (N_2594,N_2195,N_2293);
or U2595 (N_2595,N_2153,N_2057);
nand U2596 (N_2596,N_2371,N_2137);
nand U2597 (N_2597,N_2173,N_2488);
nand U2598 (N_2598,N_2381,N_2069);
and U2599 (N_2599,N_2473,N_2253);
xor U2600 (N_2600,N_2239,N_2172);
nor U2601 (N_2601,N_2130,N_2080);
nor U2602 (N_2602,N_2277,N_2227);
nor U2603 (N_2603,N_2140,N_2427);
nor U2604 (N_2604,N_2310,N_2218);
or U2605 (N_2605,N_2297,N_2075);
or U2606 (N_2606,N_2009,N_2447);
and U2607 (N_2607,N_2185,N_2271);
nor U2608 (N_2608,N_2025,N_2073);
and U2609 (N_2609,N_2054,N_2325);
xnor U2610 (N_2610,N_2033,N_2401);
and U2611 (N_2611,N_2441,N_2181);
or U2612 (N_2612,N_2329,N_2146);
nor U2613 (N_2613,N_2186,N_2215);
or U2614 (N_2614,N_2496,N_2094);
or U2615 (N_2615,N_2414,N_2171);
and U2616 (N_2616,N_2300,N_2037);
nand U2617 (N_2617,N_2118,N_2198);
and U2618 (N_2618,N_2317,N_2499);
nor U2619 (N_2619,N_2066,N_2166);
or U2620 (N_2620,N_2394,N_2268);
and U2621 (N_2621,N_2158,N_2287);
nand U2622 (N_2622,N_2249,N_2174);
nand U2623 (N_2623,N_2012,N_2005);
nor U2624 (N_2624,N_2377,N_2428);
nand U2625 (N_2625,N_2475,N_2366);
nand U2626 (N_2626,N_2086,N_2262);
and U2627 (N_2627,N_2349,N_2251);
and U2628 (N_2628,N_2061,N_2104);
and U2629 (N_2629,N_2178,N_2403);
nor U2630 (N_2630,N_2204,N_2107);
nor U2631 (N_2631,N_2445,N_2168);
nand U2632 (N_2632,N_2115,N_2223);
nor U2633 (N_2633,N_2348,N_2120);
xor U2634 (N_2634,N_2001,N_2162);
or U2635 (N_2635,N_2487,N_2208);
nand U2636 (N_2636,N_2450,N_2339);
nand U2637 (N_2637,N_2003,N_2234);
nand U2638 (N_2638,N_2106,N_2092);
and U2639 (N_2639,N_2396,N_2182);
and U2640 (N_2640,N_2097,N_2431);
nor U2641 (N_2641,N_2464,N_2160);
and U2642 (N_2642,N_2459,N_2456);
and U2643 (N_2643,N_2286,N_2121);
nor U2644 (N_2644,N_2015,N_2323);
and U2645 (N_2645,N_2045,N_2229);
nand U2646 (N_2646,N_2436,N_2393);
xor U2647 (N_2647,N_2163,N_2139);
nand U2648 (N_2648,N_2155,N_2303);
nor U2649 (N_2649,N_2477,N_2067);
nand U2650 (N_2650,N_2144,N_2161);
xor U2651 (N_2651,N_2006,N_2038);
or U2652 (N_2652,N_2136,N_2337);
and U2653 (N_2653,N_2255,N_2481);
or U2654 (N_2654,N_2340,N_2280);
or U2655 (N_2655,N_2246,N_2369);
or U2656 (N_2656,N_2288,N_2361);
nor U2657 (N_2657,N_2157,N_2388);
or U2658 (N_2658,N_2019,N_2084);
or U2659 (N_2659,N_2035,N_2210);
nand U2660 (N_2660,N_2194,N_2212);
and U2661 (N_2661,N_2410,N_2098);
and U2662 (N_2662,N_2247,N_2110);
or U2663 (N_2663,N_2345,N_2233);
nor U2664 (N_2664,N_2261,N_2152);
or U2665 (N_2665,N_2421,N_2336);
or U2666 (N_2666,N_2134,N_2062);
and U2667 (N_2667,N_2324,N_2353);
nand U2668 (N_2668,N_2468,N_2305);
and U2669 (N_2669,N_2088,N_2274);
and U2670 (N_2670,N_2374,N_2220);
nor U2671 (N_2671,N_2347,N_2338);
or U2672 (N_2672,N_2409,N_2124);
and U2673 (N_2673,N_2007,N_2010);
nand U2674 (N_2674,N_2048,N_2193);
nand U2675 (N_2675,N_2154,N_2083);
or U2676 (N_2676,N_2023,N_2452);
nand U2677 (N_2677,N_2145,N_2331);
and U2678 (N_2678,N_2176,N_2000);
nand U2679 (N_2679,N_2376,N_2332);
and U2680 (N_2680,N_2472,N_2016);
and U2681 (N_2681,N_2034,N_2301);
or U2682 (N_2682,N_2180,N_2049);
nand U2683 (N_2683,N_2471,N_2434);
xor U2684 (N_2684,N_2285,N_2150);
nor U2685 (N_2685,N_2022,N_2405);
nor U2686 (N_2686,N_2463,N_2342);
or U2687 (N_2687,N_2402,N_2237);
and U2688 (N_2688,N_2190,N_2077);
nand U2689 (N_2689,N_2021,N_2304);
and U2690 (N_2690,N_2357,N_2380);
xnor U2691 (N_2691,N_2206,N_2199);
and U2692 (N_2692,N_2322,N_2149);
nor U2693 (N_2693,N_2159,N_2315);
or U2694 (N_2694,N_2417,N_2056);
xor U2695 (N_2695,N_2398,N_2279);
nor U2696 (N_2696,N_2460,N_2378);
or U2697 (N_2697,N_2478,N_2327);
nand U2698 (N_2698,N_2480,N_2426);
nand U2699 (N_2699,N_2383,N_2183);
nand U2700 (N_2700,N_2102,N_2299);
nand U2701 (N_2701,N_2494,N_2122);
nand U2702 (N_2702,N_2101,N_2187);
nand U2703 (N_2703,N_2126,N_2389);
nor U2704 (N_2704,N_2453,N_2040);
or U2705 (N_2705,N_2044,N_2133);
and U2706 (N_2706,N_2078,N_2041);
and U2707 (N_2707,N_2030,N_2495);
nand U2708 (N_2708,N_2326,N_2068);
and U2709 (N_2709,N_2400,N_2100);
or U2710 (N_2710,N_2164,N_2017);
and U2711 (N_2711,N_2320,N_2466);
nand U2712 (N_2712,N_2476,N_2420);
xnor U2713 (N_2713,N_2282,N_2132);
xor U2714 (N_2714,N_2225,N_2179);
nor U2715 (N_2715,N_2263,N_2362);
nand U2716 (N_2716,N_2363,N_2482);
xnor U2717 (N_2717,N_2235,N_2449);
or U2718 (N_2718,N_2413,N_2059);
nor U2719 (N_2719,N_2275,N_2497);
xnor U2720 (N_2720,N_2055,N_2232);
and U2721 (N_2721,N_2330,N_2272);
nand U2722 (N_2722,N_2214,N_2243);
or U2723 (N_2723,N_2072,N_2125);
nor U2724 (N_2724,N_2070,N_2360);
or U2725 (N_2725,N_2074,N_2467);
or U2726 (N_2726,N_2375,N_2284);
xnor U2727 (N_2727,N_2002,N_2076);
xor U2728 (N_2728,N_2051,N_2091);
nand U2729 (N_2729,N_2422,N_2462);
nor U2730 (N_2730,N_2435,N_2370);
nand U2731 (N_2731,N_2117,N_2483);
or U2732 (N_2732,N_2425,N_2266);
xor U2733 (N_2733,N_2415,N_2095);
and U2734 (N_2734,N_2196,N_2485);
or U2735 (N_2735,N_2228,N_2295);
nand U2736 (N_2736,N_2283,N_2350);
nor U2737 (N_2737,N_2238,N_2335);
or U2738 (N_2738,N_2269,N_2264);
nor U2739 (N_2739,N_2319,N_2031);
and U2740 (N_2740,N_2368,N_2043);
nand U2741 (N_2741,N_2437,N_2205);
xor U2742 (N_2742,N_2265,N_2469);
nand U2743 (N_2743,N_2458,N_2216);
nand U2744 (N_2744,N_2430,N_2029);
nor U2745 (N_2745,N_2446,N_2197);
nand U2746 (N_2746,N_2407,N_2175);
and U2747 (N_2747,N_2222,N_2053);
or U2748 (N_2748,N_2128,N_2203);
or U2749 (N_2749,N_2267,N_2211);
or U2750 (N_2750,N_2420,N_2081);
or U2751 (N_2751,N_2299,N_2239);
nor U2752 (N_2752,N_2441,N_2137);
and U2753 (N_2753,N_2164,N_2038);
nor U2754 (N_2754,N_2171,N_2347);
nor U2755 (N_2755,N_2205,N_2279);
nor U2756 (N_2756,N_2150,N_2066);
and U2757 (N_2757,N_2340,N_2081);
nand U2758 (N_2758,N_2263,N_2250);
nand U2759 (N_2759,N_2367,N_2198);
nor U2760 (N_2760,N_2005,N_2493);
or U2761 (N_2761,N_2420,N_2097);
or U2762 (N_2762,N_2287,N_2021);
or U2763 (N_2763,N_2251,N_2259);
and U2764 (N_2764,N_2339,N_2260);
nand U2765 (N_2765,N_2049,N_2478);
or U2766 (N_2766,N_2325,N_2048);
nand U2767 (N_2767,N_2326,N_2466);
and U2768 (N_2768,N_2097,N_2173);
nand U2769 (N_2769,N_2280,N_2362);
nand U2770 (N_2770,N_2094,N_2349);
nor U2771 (N_2771,N_2352,N_2091);
and U2772 (N_2772,N_2325,N_2207);
nor U2773 (N_2773,N_2326,N_2058);
and U2774 (N_2774,N_2452,N_2399);
xor U2775 (N_2775,N_2399,N_2114);
nand U2776 (N_2776,N_2381,N_2297);
or U2777 (N_2777,N_2352,N_2215);
and U2778 (N_2778,N_2474,N_2217);
or U2779 (N_2779,N_2259,N_2084);
nor U2780 (N_2780,N_2136,N_2431);
xnor U2781 (N_2781,N_2428,N_2034);
nor U2782 (N_2782,N_2367,N_2024);
nand U2783 (N_2783,N_2440,N_2407);
or U2784 (N_2784,N_2302,N_2088);
nand U2785 (N_2785,N_2496,N_2087);
nand U2786 (N_2786,N_2422,N_2032);
nand U2787 (N_2787,N_2435,N_2440);
and U2788 (N_2788,N_2455,N_2348);
xor U2789 (N_2789,N_2327,N_2442);
or U2790 (N_2790,N_2465,N_2468);
nor U2791 (N_2791,N_2389,N_2337);
nor U2792 (N_2792,N_2010,N_2106);
and U2793 (N_2793,N_2131,N_2259);
or U2794 (N_2794,N_2053,N_2321);
and U2795 (N_2795,N_2183,N_2213);
xnor U2796 (N_2796,N_2421,N_2396);
nand U2797 (N_2797,N_2443,N_2238);
and U2798 (N_2798,N_2123,N_2033);
nor U2799 (N_2799,N_2132,N_2066);
xor U2800 (N_2800,N_2135,N_2459);
and U2801 (N_2801,N_2031,N_2007);
nor U2802 (N_2802,N_2408,N_2054);
and U2803 (N_2803,N_2233,N_2135);
xnor U2804 (N_2804,N_2203,N_2013);
or U2805 (N_2805,N_2094,N_2248);
xor U2806 (N_2806,N_2267,N_2011);
and U2807 (N_2807,N_2390,N_2247);
nand U2808 (N_2808,N_2429,N_2155);
nand U2809 (N_2809,N_2240,N_2162);
or U2810 (N_2810,N_2134,N_2019);
xnor U2811 (N_2811,N_2350,N_2274);
xnor U2812 (N_2812,N_2081,N_2005);
or U2813 (N_2813,N_2069,N_2340);
nor U2814 (N_2814,N_2202,N_2431);
and U2815 (N_2815,N_2326,N_2152);
nor U2816 (N_2816,N_2434,N_2335);
nand U2817 (N_2817,N_2293,N_2013);
nand U2818 (N_2818,N_2177,N_2302);
xor U2819 (N_2819,N_2487,N_2124);
and U2820 (N_2820,N_2321,N_2424);
xor U2821 (N_2821,N_2137,N_2339);
xnor U2822 (N_2822,N_2093,N_2495);
nor U2823 (N_2823,N_2093,N_2310);
xnor U2824 (N_2824,N_2212,N_2452);
or U2825 (N_2825,N_2176,N_2109);
or U2826 (N_2826,N_2209,N_2152);
xnor U2827 (N_2827,N_2099,N_2151);
or U2828 (N_2828,N_2271,N_2081);
or U2829 (N_2829,N_2089,N_2336);
nand U2830 (N_2830,N_2117,N_2265);
nor U2831 (N_2831,N_2152,N_2240);
or U2832 (N_2832,N_2360,N_2230);
and U2833 (N_2833,N_2441,N_2442);
nand U2834 (N_2834,N_2418,N_2266);
nand U2835 (N_2835,N_2213,N_2219);
and U2836 (N_2836,N_2037,N_2442);
and U2837 (N_2837,N_2214,N_2010);
and U2838 (N_2838,N_2157,N_2439);
nand U2839 (N_2839,N_2345,N_2232);
nor U2840 (N_2840,N_2299,N_2420);
nor U2841 (N_2841,N_2367,N_2230);
and U2842 (N_2842,N_2043,N_2075);
or U2843 (N_2843,N_2026,N_2024);
or U2844 (N_2844,N_2191,N_2183);
nand U2845 (N_2845,N_2249,N_2359);
or U2846 (N_2846,N_2179,N_2122);
nor U2847 (N_2847,N_2404,N_2204);
xnor U2848 (N_2848,N_2160,N_2321);
or U2849 (N_2849,N_2111,N_2349);
nor U2850 (N_2850,N_2438,N_2131);
or U2851 (N_2851,N_2027,N_2440);
and U2852 (N_2852,N_2284,N_2007);
nor U2853 (N_2853,N_2393,N_2351);
nand U2854 (N_2854,N_2120,N_2119);
nor U2855 (N_2855,N_2328,N_2465);
xor U2856 (N_2856,N_2473,N_2220);
xor U2857 (N_2857,N_2310,N_2352);
and U2858 (N_2858,N_2216,N_2031);
or U2859 (N_2859,N_2199,N_2212);
nand U2860 (N_2860,N_2300,N_2494);
xnor U2861 (N_2861,N_2433,N_2154);
nor U2862 (N_2862,N_2292,N_2259);
and U2863 (N_2863,N_2381,N_2415);
or U2864 (N_2864,N_2156,N_2014);
nor U2865 (N_2865,N_2489,N_2450);
nand U2866 (N_2866,N_2215,N_2187);
nand U2867 (N_2867,N_2357,N_2150);
nand U2868 (N_2868,N_2367,N_2491);
or U2869 (N_2869,N_2306,N_2012);
or U2870 (N_2870,N_2370,N_2236);
nor U2871 (N_2871,N_2002,N_2024);
and U2872 (N_2872,N_2066,N_2389);
nor U2873 (N_2873,N_2452,N_2373);
nand U2874 (N_2874,N_2035,N_2447);
nor U2875 (N_2875,N_2381,N_2043);
and U2876 (N_2876,N_2015,N_2494);
or U2877 (N_2877,N_2041,N_2415);
and U2878 (N_2878,N_2335,N_2277);
nand U2879 (N_2879,N_2191,N_2305);
nor U2880 (N_2880,N_2399,N_2294);
and U2881 (N_2881,N_2213,N_2137);
nor U2882 (N_2882,N_2072,N_2130);
nand U2883 (N_2883,N_2194,N_2410);
nor U2884 (N_2884,N_2306,N_2438);
and U2885 (N_2885,N_2357,N_2458);
nand U2886 (N_2886,N_2201,N_2444);
nand U2887 (N_2887,N_2373,N_2143);
nand U2888 (N_2888,N_2086,N_2328);
nand U2889 (N_2889,N_2205,N_2229);
or U2890 (N_2890,N_2495,N_2440);
xnor U2891 (N_2891,N_2496,N_2407);
and U2892 (N_2892,N_2146,N_2195);
nand U2893 (N_2893,N_2352,N_2433);
and U2894 (N_2894,N_2267,N_2472);
and U2895 (N_2895,N_2455,N_2174);
xnor U2896 (N_2896,N_2440,N_2171);
nor U2897 (N_2897,N_2072,N_2078);
nor U2898 (N_2898,N_2384,N_2407);
nand U2899 (N_2899,N_2271,N_2045);
and U2900 (N_2900,N_2414,N_2100);
nor U2901 (N_2901,N_2397,N_2111);
or U2902 (N_2902,N_2147,N_2404);
nand U2903 (N_2903,N_2450,N_2140);
nand U2904 (N_2904,N_2286,N_2148);
nand U2905 (N_2905,N_2000,N_2216);
and U2906 (N_2906,N_2283,N_2041);
nor U2907 (N_2907,N_2274,N_2430);
nor U2908 (N_2908,N_2018,N_2444);
nand U2909 (N_2909,N_2353,N_2395);
xor U2910 (N_2910,N_2056,N_2407);
or U2911 (N_2911,N_2302,N_2370);
and U2912 (N_2912,N_2218,N_2433);
xor U2913 (N_2913,N_2402,N_2014);
nor U2914 (N_2914,N_2467,N_2111);
nand U2915 (N_2915,N_2307,N_2383);
and U2916 (N_2916,N_2209,N_2182);
and U2917 (N_2917,N_2095,N_2234);
nand U2918 (N_2918,N_2065,N_2409);
or U2919 (N_2919,N_2382,N_2474);
nor U2920 (N_2920,N_2389,N_2302);
xnor U2921 (N_2921,N_2006,N_2179);
nand U2922 (N_2922,N_2278,N_2201);
and U2923 (N_2923,N_2003,N_2336);
nand U2924 (N_2924,N_2306,N_2245);
nor U2925 (N_2925,N_2212,N_2378);
and U2926 (N_2926,N_2249,N_2294);
nor U2927 (N_2927,N_2397,N_2077);
or U2928 (N_2928,N_2291,N_2358);
and U2929 (N_2929,N_2359,N_2291);
nand U2930 (N_2930,N_2351,N_2103);
nand U2931 (N_2931,N_2348,N_2109);
nor U2932 (N_2932,N_2195,N_2469);
and U2933 (N_2933,N_2040,N_2480);
nand U2934 (N_2934,N_2434,N_2155);
and U2935 (N_2935,N_2141,N_2360);
nor U2936 (N_2936,N_2151,N_2219);
nor U2937 (N_2937,N_2015,N_2315);
nand U2938 (N_2938,N_2067,N_2355);
xor U2939 (N_2939,N_2297,N_2353);
xnor U2940 (N_2940,N_2008,N_2433);
nand U2941 (N_2941,N_2012,N_2322);
and U2942 (N_2942,N_2473,N_2467);
or U2943 (N_2943,N_2458,N_2143);
or U2944 (N_2944,N_2247,N_2255);
nand U2945 (N_2945,N_2402,N_2082);
nand U2946 (N_2946,N_2405,N_2261);
nor U2947 (N_2947,N_2130,N_2126);
xor U2948 (N_2948,N_2143,N_2272);
nor U2949 (N_2949,N_2210,N_2368);
or U2950 (N_2950,N_2142,N_2452);
or U2951 (N_2951,N_2289,N_2213);
and U2952 (N_2952,N_2368,N_2201);
and U2953 (N_2953,N_2345,N_2330);
nor U2954 (N_2954,N_2124,N_2114);
or U2955 (N_2955,N_2097,N_2142);
nand U2956 (N_2956,N_2167,N_2338);
or U2957 (N_2957,N_2196,N_2355);
xor U2958 (N_2958,N_2052,N_2279);
nand U2959 (N_2959,N_2376,N_2402);
and U2960 (N_2960,N_2165,N_2006);
nor U2961 (N_2961,N_2015,N_2264);
nand U2962 (N_2962,N_2041,N_2065);
or U2963 (N_2963,N_2225,N_2080);
and U2964 (N_2964,N_2413,N_2398);
xor U2965 (N_2965,N_2407,N_2062);
xnor U2966 (N_2966,N_2009,N_2156);
xor U2967 (N_2967,N_2437,N_2042);
and U2968 (N_2968,N_2131,N_2381);
nand U2969 (N_2969,N_2041,N_2149);
or U2970 (N_2970,N_2352,N_2466);
nand U2971 (N_2971,N_2108,N_2067);
nor U2972 (N_2972,N_2105,N_2411);
nor U2973 (N_2973,N_2084,N_2467);
and U2974 (N_2974,N_2457,N_2438);
xnor U2975 (N_2975,N_2027,N_2421);
nand U2976 (N_2976,N_2382,N_2353);
xor U2977 (N_2977,N_2330,N_2211);
nand U2978 (N_2978,N_2349,N_2404);
nand U2979 (N_2979,N_2144,N_2300);
or U2980 (N_2980,N_2331,N_2174);
nand U2981 (N_2981,N_2272,N_2140);
nand U2982 (N_2982,N_2154,N_2072);
or U2983 (N_2983,N_2366,N_2152);
nand U2984 (N_2984,N_2493,N_2104);
and U2985 (N_2985,N_2201,N_2259);
nand U2986 (N_2986,N_2239,N_2021);
or U2987 (N_2987,N_2008,N_2026);
nor U2988 (N_2988,N_2456,N_2438);
xor U2989 (N_2989,N_2190,N_2300);
xnor U2990 (N_2990,N_2021,N_2078);
nor U2991 (N_2991,N_2338,N_2383);
nand U2992 (N_2992,N_2161,N_2353);
and U2993 (N_2993,N_2347,N_2233);
and U2994 (N_2994,N_2029,N_2245);
or U2995 (N_2995,N_2411,N_2360);
and U2996 (N_2996,N_2248,N_2165);
nor U2997 (N_2997,N_2451,N_2351);
and U2998 (N_2998,N_2387,N_2177);
or U2999 (N_2999,N_2498,N_2245);
xnor U3000 (N_3000,N_2756,N_2919);
and U3001 (N_3001,N_2621,N_2616);
and U3002 (N_3002,N_2559,N_2906);
nand U3003 (N_3003,N_2887,N_2830);
and U3004 (N_3004,N_2568,N_2913);
nand U3005 (N_3005,N_2805,N_2813);
nand U3006 (N_3006,N_2845,N_2920);
and U3007 (N_3007,N_2723,N_2950);
xnor U3008 (N_3008,N_2793,N_2938);
xnor U3009 (N_3009,N_2580,N_2758);
nor U3010 (N_3010,N_2860,N_2940);
and U3011 (N_3011,N_2992,N_2914);
xor U3012 (N_3012,N_2754,N_2874);
or U3013 (N_3013,N_2833,N_2869);
nand U3014 (N_3014,N_2625,N_2923);
nor U3015 (N_3015,N_2769,N_2942);
nor U3016 (N_3016,N_2853,N_2900);
and U3017 (N_3017,N_2708,N_2542);
nor U3018 (N_3018,N_2522,N_2789);
and U3019 (N_3019,N_2885,N_2979);
nor U3020 (N_3020,N_2948,N_2589);
or U3021 (N_3021,N_2868,N_2560);
nor U3022 (N_3022,N_2893,N_2693);
or U3023 (N_3023,N_2867,N_2840);
or U3024 (N_3024,N_2533,N_2976);
nor U3025 (N_3025,N_2683,N_2815);
nand U3026 (N_3026,N_2788,N_2565);
nor U3027 (N_3027,N_2806,N_2669);
xnor U3028 (N_3028,N_2782,N_2932);
nor U3029 (N_3029,N_2956,N_2516);
and U3030 (N_3030,N_2988,N_2578);
nor U3031 (N_3031,N_2768,N_2643);
and U3032 (N_3032,N_2785,N_2753);
nand U3033 (N_3033,N_2779,N_2912);
nor U3034 (N_3034,N_2889,N_2891);
nand U3035 (N_3035,N_2841,N_2777);
and U3036 (N_3036,N_2811,N_2528);
nand U3037 (N_3037,N_2743,N_2575);
and U3038 (N_3038,N_2663,N_2604);
and U3039 (N_3039,N_2832,N_2744);
or U3040 (N_3040,N_2807,N_2918);
and U3041 (N_3041,N_2761,N_2986);
nor U3042 (N_3042,N_2958,N_2687);
or U3043 (N_3043,N_2558,N_2509);
xor U3044 (N_3044,N_2981,N_2762);
nor U3045 (N_3045,N_2880,N_2549);
or U3046 (N_3046,N_2664,N_2633);
xor U3047 (N_3047,N_2883,N_2968);
nor U3048 (N_3048,N_2747,N_2757);
and U3049 (N_3049,N_2775,N_2943);
nand U3050 (N_3050,N_2688,N_2978);
nand U3051 (N_3051,N_2639,N_2704);
or U3052 (N_3052,N_2573,N_2917);
and U3053 (N_3053,N_2530,N_2647);
and U3054 (N_3054,N_2847,N_2929);
xnor U3055 (N_3055,N_2725,N_2588);
or U3056 (N_3056,N_2982,N_2784);
nor U3057 (N_3057,N_2962,N_2545);
or U3058 (N_3058,N_2836,N_2718);
or U3059 (N_3059,N_2995,N_2808);
nand U3060 (N_3060,N_2652,N_2823);
nor U3061 (N_3061,N_2872,N_2554);
nor U3062 (N_3062,N_2724,N_2595);
and U3063 (N_3063,N_2925,N_2812);
xor U3064 (N_3064,N_2682,N_2680);
and U3065 (N_3065,N_2671,N_2760);
and U3066 (N_3066,N_2577,N_2928);
and U3067 (N_3067,N_2649,N_2609);
nand U3068 (N_3068,N_2751,N_2571);
nand U3069 (N_3069,N_2967,N_2903);
and U3070 (N_3070,N_2878,N_2644);
and U3071 (N_3071,N_2865,N_2689);
nand U3072 (N_3072,N_2921,N_2701);
nor U3073 (N_3073,N_2875,N_2745);
nor U3074 (N_3074,N_2692,N_2684);
and U3075 (N_3075,N_2896,N_2628);
nor U3076 (N_3076,N_2685,N_2630);
and U3077 (N_3077,N_2966,N_2672);
nor U3078 (N_3078,N_2722,N_2646);
xnor U3079 (N_3079,N_2977,N_2697);
and U3080 (N_3080,N_2567,N_2668);
nor U3081 (N_3081,N_2935,N_2716);
or U3082 (N_3082,N_2505,N_2947);
or U3083 (N_3083,N_2766,N_2907);
or U3084 (N_3084,N_2615,N_2605);
or U3085 (N_3085,N_2667,N_2892);
and U3086 (N_3086,N_2746,N_2719);
nor U3087 (N_3087,N_2911,N_2705);
and U3088 (N_3088,N_2820,N_2791);
or U3089 (N_3089,N_2537,N_2711);
nor U3090 (N_3090,N_2500,N_2710);
xor U3091 (N_3091,N_2698,N_2562);
nor U3092 (N_3092,N_2946,N_2957);
nor U3093 (N_3093,N_2737,N_2510);
xor U3094 (N_3094,N_2729,N_2518);
or U3095 (N_3095,N_2980,N_2648);
or U3096 (N_3096,N_2521,N_2608);
nor U3097 (N_3097,N_2749,N_2690);
or U3098 (N_3098,N_2894,N_2563);
and U3099 (N_3099,N_2694,N_2764);
and U3100 (N_3100,N_2547,N_2534);
nand U3101 (N_3101,N_2674,N_2888);
xor U3102 (N_3102,N_2984,N_2770);
nor U3103 (N_3103,N_2787,N_2863);
nor U3104 (N_3104,N_2582,N_2622);
xor U3105 (N_3105,N_2733,N_2679);
or U3106 (N_3106,N_2523,N_2797);
nor U3107 (N_3107,N_2798,N_2862);
nand U3108 (N_3108,N_2792,N_2529);
nor U3109 (N_3109,N_2842,N_2598);
and U3110 (N_3110,N_2513,N_2816);
nor U3111 (N_3111,N_2910,N_2707);
nor U3112 (N_3112,N_2996,N_2546);
and U3113 (N_3113,N_2606,N_2959);
nor U3114 (N_3114,N_2810,N_2566);
and U3115 (N_3115,N_2825,N_2656);
or U3116 (N_3116,N_2517,N_2717);
or U3117 (N_3117,N_2802,N_2826);
or U3118 (N_3118,N_2944,N_2933);
and U3119 (N_3119,N_2972,N_2819);
xnor U3120 (N_3120,N_2613,N_2673);
and U3121 (N_3121,N_2866,N_2829);
and U3122 (N_3122,N_2964,N_2817);
and U3123 (N_3123,N_2736,N_2922);
nor U3124 (N_3124,N_2607,N_2963);
nand U3125 (N_3125,N_2501,N_2596);
nand U3126 (N_3126,N_2991,N_2678);
nand U3127 (N_3127,N_2583,N_2709);
or U3128 (N_3128,N_2654,N_2650);
and U3129 (N_3129,N_2726,N_2532);
or U3130 (N_3130,N_2740,N_2732);
xor U3131 (N_3131,N_2601,N_2702);
xor U3132 (N_3132,N_2844,N_2540);
nor U3133 (N_3133,N_2640,N_2965);
or U3134 (N_3134,N_2850,N_2994);
and U3135 (N_3135,N_2626,N_2548);
nand U3136 (N_3136,N_2783,N_2750);
or U3137 (N_3137,N_2727,N_2586);
or U3138 (N_3138,N_2954,N_2666);
and U3139 (N_3139,N_2553,N_2610);
or U3140 (N_3140,N_2511,N_2675);
nor U3141 (N_3141,N_2951,N_2855);
or U3142 (N_3142,N_2795,N_2773);
nand U3143 (N_3143,N_2949,N_2915);
nand U3144 (N_3144,N_2641,N_2712);
or U3145 (N_3145,N_2902,N_2508);
nor U3146 (N_3146,N_2636,N_2945);
or U3147 (N_3147,N_2786,N_2714);
xor U3148 (N_3148,N_2552,N_2818);
and U3149 (N_3149,N_2801,N_2585);
or U3150 (N_3150,N_2512,N_2550);
nand U3151 (N_3151,N_2635,N_2752);
and U3152 (N_3152,N_2890,N_2504);
or U3153 (N_3153,N_2642,N_2857);
or U3154 (N_3154,N_2882,N_2557);
or U3155 (N_3155,N_2539,N_2824);
nor U3156 (N_3156,N_2846,N_2686);
and U3157 (N_3157,N_2941,N_2765);
nand U3158 (N_3158,N_2561,N_2515);
nand U3159 (N_3159,N_2720,N_2657);
and U3160 (N_3160,N_2527,N_2843);
or U3161 (N_3161,N_2973,N_2771);
nand U3162 (N_3162,N_2936,N_2871);
and U3163 (N_3163,N_2937,N_2898);
nand U3164 (N_3164,N_2838,N_2570);
and U3165 (N_3165,N_2612,N_2828);
and U3166 (N_3166,N_2519,N_2993);
or U3167 (N_3167,N_2763,N_2873);
nor U3168 (N_3168,N_2955,N_2681);
and U3169 (N_3169,N_2886,N_2879);
nand U3170 (N_3170,N_2658,N_2877);
and U3171 (N_3171,N_2634,N_2631);
nor U3172 (N_3172,N_2599,N_2526);
or U3173 (N_3173,N_2574,N_2696);
xor U3174 (N_3174,N_2627,N_2555);
or U3175 (N_3175,N_2971,N_2794);
nand U3176 (N_3176,N_2904,N_2572);
or U3177 (N_3177,N_2854,N_2861);
nand U3178 (N_3178,N_2593,N_2576);
and U3179 (N_3179,N_2677,N_2665);
nor U3180 (N_3180,N_2809,N_2541);
or U3181 (N_3181,N_2556,N_2632);
and U3182 (N_3182,N_2901,N_2551);
nand U3183 (N_3183,N_2790,N_2738);
or U3184 (N_3184,N_2543,N_2905);
nand U3185 (N_3185,N_2776,N_2623);
nand U3186 (N_3186,N_2975,N_2876);
nand U3187 (N_3187,N_2742,N_2638);
or U3188 (N_3188,N_2662,N_2590);
xnor U3189 (N_3189,N_2602,N_2814);
or U3190 (N_3190,N_2730,N_2870);
nor U3191 (N_3191,N_2864,N_2660);
or U3192 (N_3192,N_2939,N_2772);
nor U3193 (N_3193,N_2858,N_2659);
xor U3194 (N_3194,N_2617,N_2579);
and U3195 (N_3195,N_2587,N_2803);
and U3196 (N_3196,N_2895,N_2952);
nor U3197 (N_3197,N_2859,N_2851);
nand U3198 (N_3198,N_2848,N_2759);
nand U3199 (N_3199,N_2594,N_2969);
and U3200 (N_3200,N_2849,N_2503);
nor U3201 (N_3201,N_2620,N_2734);
or U3202 (N_3202,N_2974,N_2603);
or U3203 (N_3203,N_2931,N_2739);
and U3204 (N_3204,N_2999,N_2600);
xnor U3205 (N_3205,N_2514,N_2611);
and U3206 (N_3206,N_2591,N_2998);
nand U3207 (N_3207,N_2597,N_2804);
nor U3208 (N_3208,N_2691,N_2767);
and U3209 (N_3209,N_2834,N_2645);
or U3210 (N_3210,N_2524,N_2970);
xnor U3211 (N_3211,N_2655,N_2520);
or U3212 (N_3212,N_2525,N_2897);
nor U3213 (N_3213,N_2584,N_2507);
nor U3214 (N_3214,N_2569,N_2721);
and U3215 (N_3215,N_2989,N_2637);
or U3216 (N_3216,N_2629,N_2731);
and U3217 (N_3217,N_2695,N_2884);
xnor U3218 (N_3218,N_2661,N_2748);
or U3219 (N_3219,N_2618,N_2837);
xor U3220 (N_3220,N_2899,N_2778);
xnor U3221 (N_3221,N_2839,N_2916);
nand U3222 (N_3222,N_2699,N_2735);
nor U3223 (N_3223,N_2960,N_2755);
nand U3224 (N_3224,N_2502,N_2651);
nor U3225 (N_3225,N_2535,N_2983);
nor U3226 (N_3226,N_2592,N_2536);
nor U3227 (N_3227,N_2531,N_2835);
or U3228 (N_3228,N_2822,N_2506);
nor U3229 (N_3229,N_2653,N_2619);
or U3230 (N_3230,N_2852,N_2713);
nand U3231 (N_3231,N_2796,N_2728);
or U3232 (N_3232,N_2924,N_2715);
nand U3233 (N_3233,N_2538,N_2703);
and U3234 (N_3234,N_2544,N_2961);
nand U3235 (N_3235,N_2953,N_2706);
or U3236 (N_3236,N_2614,N_2827);
nor U3237 (N_3237,N_2676,N_2997);
and U3238 (N_3238,N_2799,N_2881);
nor U3239 (N_3239,N_2856,N_2927);
or U3240 (N_3240,N_2564,N_2930);
nor U3241 (N_3241,N_2985,N_2774);
nand U3242 (N_3242,N_2800,N_2581);
and U3243 (N_3243,N_2909,N_2781);
and U3244 (N_3244,N_2780,N_2908);
nand U3245 (N_3245,N_2987,N_2934);
xnor U3246 (N_3246,N_2990,N_2831);
and U3247 (N_3247,N_2624,N_2741);
or U3248 (N_3248,N_2821,N_2926);
nand U3249 (N_3249,N_2670,N_2700);
and U3250 (N_3250,N_2733,N_2967);
or U3251 (N_3251,N_2746,N_2560);
and U3252 (N_3252,N_2617,N_2606);
and U3253 (N_3253,N_2647,N_2707);
nor U3254 (N_3254,N_2652,N_2765);
nand U3255 (N_3255,N_2585,N_2548);
nor U3256 (N_3256,N_2820,N_2899);
xor U3257 (N_3257,N_2938,N_2520);
xor U3258 (N_3258,N_2954,N_2765);
and U3259 (N_3259,N_2500,N_2828);
nand U3260 (N_3260,N_2881,N_2935);
nor U3261 (N_3261,N_2897,N_2846);
and U3262 (N_3262,N_2688,N_2588);
or U3263 (N_3263,N_2880,N_2503);
nand U3264 (N_3264,N_2955,N_2691);
and U3265 (N_3265,N_2913,N_2692);
or U3266 (N_3266,N_2852,N_2720);
and U3267 (N_3267,N_2740,N_2769);
nand U3268 (N_3268,N_2781,N_2972);
nand U3269 (N_3269,N_2732,N_2835);
nand U3270 (N_3270,N_2820,N_2787);
nor U3271 (N_3271,N_2612,N_2574);
or U3272 (N_3272,N_2898,N_2801);
nor U3273 (N_3273,N_2772,N_2510);
or U3274 (N_3274,N_2976,N_2570);
and U3275 (N_3275,N_2555,N_2798);
nor U3276 (N_3276,N_2910,N_2663);
or U3277 (N_3277,N_2852,N_2693);
and U3278 (N_3278,N_2665,N_2512);
nand U3279 (N_3279,N_2929,N_2696);
nor U3280 (N_3280,N_2589,N_2651);
nor U3281 (N_3281,N_2698,N_2735);
nand U3282 (N_3282,N_2647,N_2764);
nand U3283 (N_3283,N_2819,N_2923);
or U3284 (N_3284,N_2956,N_2716);
nor U3285 (N_3285,N_2726,N_2800);
nor U3286 (N_3286,N_2752,N_2803);
nand U3287 (N_3287,N_2996,N_2824);
and U3288 (N_3288,N_2662,N_2579);
nand U3289 (N_3289,N_2773,N_2522);
and U3290 (N_3290,N_2946,N_2945);
nand U3291 (N_3291,N_2857,N_2532);
nor U3292 (N_3292,N_2959,N_2739);
or U3293 (N_3293,N_2805,N_2701);
nand U3294 (N_3294,N_2818,N_2970);
and U3295 (N_3295,N_2514,N_2516);
nor U3296 (N_3296,N_2648,N_2948);
or U3297 (N_3297,N_2935,N_2693);
or U3298 (N_3298,N_2635,N_2955);
nand U3299 (N_3299,N_2847,N_2667);
nor U3300 (N_3300,N_2730,N_2865);
xor U3301 (N_3301,N_2900,N_2808);
or U3302 (N_3302,N_2986,N_2520);
nand U3303 (N_3303,N_2501,N_2614);
nor U3304 (N_3304,N_2541,N_2629);
nor U3305 (N_3305,N_2757,N_2732);
and U3306 (N_3306,N_2890,N_2585);
nor U3307 (N_3307,N_2968,N_2913);
nor U3308 (N_3308,N_2910,N_2966);
or U3309 (N_3309,N_2743,N_2963);
nor U3310 (N_3310,N_2539,N_2615);
nand U3311 (N_3311,N_2905,N_2913);
or U3312 (N_3312,N_2609,N_2519);
xor U3313 (N_3313,N_2730,N_2609);
nand U3314 (N_3314,N_2897,N_2516);
nor U3315 (N_3315,N_2963,N_2537);
nor U3316 (N_3316,N_2770,N_2980);
nand U3317 (N_3317,N_2507,N_2921);
or U3318 (N_3318,N_2648,N_2750);
and U3319 (N_3319,N_2907,N_2557);
nand U3320 (N_3320,N_2999,N_2647);
and U3321 (N_3321,N_2592,N_2763);
nor U3322 (N_3322,N_2710,N_2818);
nand U3323 (N_3323,N_2681,N_2808);
nand U3324 (N_3324,N_2501,N_2955);
and U3325 (N_3325,N_2722,N_2757);
and U3326 (N_3326,N_2577,N_2610);
or U3327 (N_3327,N_2883,N_2738);
nand U3328 (N_3328,N_2803,N_2741);
or U3329 (N_3329,N_2686,N_2560);
nand U3330 (N_3330,N_2864,N_2887);
nor U3331 (N_3331,N_2606,N_2871);
or U3332 (N_3332,N_2534,N_2948);
nand U3333 (N_3333,N_2831,N_2735);
nor U3334 (N_3334,N_2978,N_2987);
xnor U3335 (N_3335,N_2665,N_2648);
nor U3336 (N_3336,N_2576,N_2573);
and U3337 (N_3337,N_2936,N_2510);
or U3338 (N_3338,N_2857,N_2965);
or U3339 (N_3339,N_2934,N_2911);
nor U3340 (N_3340,N_2638,N_2558);
nor U3341 (N_3341,N_2904,N_2626);
or U3342 (N_3342,N_2549,N_2873);
nor U3343 (N_3343,N_2994,N_2913);
and U3344 (N_3344,N_2766,N_2930);
and U3345 (N_3345,N_2823,N_2506);
and U3346 (N_3346,N_2956,N_2964);
or U3347 (N_3347,N_2533,N_2741);
and U3348 (N_3348,N_2563,N_2693);
or U3349 (N_3349,N_2718,N_2813);
nor U3350 (N_3350,N_2926,N_2728);
or U3351 (N_3351,N_2759,N_2559);
and U3352 (N_3352,N_2792,N_2507);
and U3353 (N_3353,N_2856,N_2544);
and U3354 (N_3354,N_2521,N_2576);
or U3355 (N_3355,N_2998,N_2936);
nand U3356 (N_3356,N_2552,N_2627);
or U3357 (N_3357,N_2570,N_2843);
nor U3358 (N_3358,N_2617,N_2652);
or U3359 (N_3359,N_2593,N_2843);
nor U3360 (N_3360,N_2982,N_2570);
nand U3361 (N_3361,N_2982,N_2552);
or U3362 (N_3362,N_2946,N_2867);
or U3363 (N_3363,N_2866,N_2645);
xnor U3364 (N_3364,N_2629,N_2984);
nor U3365 (N_3365,N_2692,N_2945);
and U3366 (N_3366,N_2633,N_2926);
or U3367 (N_3367,N_2907,N_2662);
and U3368 (N_3368,N_2630,N_2798);
xor U3369 (N_3369,N_2814,N_2771);
xnor U3370 (N_3370,N_2906,N_2790);
or U3371 (N_3371,N_2525,N_2544);
xor U3372 (N_3372,N_2595,N_2698);
xnor U3373 (N_3373,N_2560,N_2678);
or U3374 (N_3374,N_2511,N_2910);
nor U3375 (N_3375,N_2868,N_2672);
xnor U3376 (N_3376,N_2748,N_2610);
nand U3377 (N_3377,N_2842,N_2509);
or U3378 (N_3378,N_2568,N_2814);
nand U3379 (N_3379,N_2705,N_2726);
xnor U3380 (N_3380,N_2824,N_2965);
nand U3381 (N_3381,N_2713,N_2778);
or U3382 (N_3382,N_2707,N_2713);
nor U3383 (N_3383,N_2710,N_2810);
nor U3384 (N_3384,N_2817,N_2821);
or U3385 (N_3385,N_2756,N_2597);
and U3386 (N_3386,N_2588,N_2627);
nor U3387 (N_3387,N_2535,N_2814);
or U3388 (N_3388,N_2632,N_2842);
or U3389 (N_3389,N_2788,N_2665);
and U3390 (N_3390,N_2753,N_2951);
and U3391 (N_3391,N_2726,N_2740);
and U3392 (N_3392,N_2531,N_2637);
or U3393 (N_3393,N_2595,N_2631);
or U3394 (N_3394,N_2556,N_2553);
nor U3395 (N_3395,N_2601,N_2752);
or U3396 (N_3396,N_2816,N_2518);
and U3397 (N_3397,N_2726,N_2612);
nand U3398 (N_3398,N_2730,N_2680);
and U3399 (N_3399,N_2934,N_2702);
nand U3400 (N_3400,N_2792,N_2858);
nand U3401 (N_3401,N_2548,N_2721);
and U3402 (N_3402,N_2624,N_2869);
nor U3403 (N_3403,N_2627,N_2636);
or U3404 (N_3404,N_2554,N_2774);
and U3405 (N_3405,N_2631,N_2817);
nor U3406 (N_3406,N_2568,N_2808);
nand U3407 (N_3407,N_2588,N_2983);
and U3408 (N_3408,N_2719,N_2829);
nor U3409 (N_3409,N_2857,N_2752);
or U3410 (N_3410,N_2624,N_2526);
nand U3411 (N_3411,N_2666,N_2804);
xor U3412 (N_3412,N_2842,N_2514);
nor U3413 (N_3413,N_2684,N_2887);
nor U3414 (N_3414,N_2829,N_2585);
nand U3415 (N_3415,N_2743,N_2767);
nor U3416 (N_3416,N_2579,N_2651);
nand U3417 (N_3417,N_2545,N_2771);
and U3418 (N_3418,N_2579,N_2895);
and U3419 (N_3419,N_2634,N_2643);
nand U3420 (N_3420,N_2837,N_2512);
nor U3421 (N_3421,N_2660,N_2904);
nor U3422 (N_3422,N_2651,N_2653);
nor U3423 (N_3423,N_2892,N_2756);
nand U3424 (N_3424,N_2720,N_2583);
and U3425 (N_3425,N_2890,N_2992);
or U3426 (N_3426,N_2988,N_2545);
and U3427 (N_3427,N_2888,N_2996);
nor U3428 (N_3428,N_2623,N_2793);
or U3429 (N_3429,N_2792,N_2588);
and U3430 (N_3430,N_2500,N_2628);
and U3431 (N_3431,N_2954,N_2699);
nor U3432 (N_3432,N_2656,N_2895);
or U3433 (N_3433,N_2710,N_2980);
nor U3434 (N_3434,N_2827,N_2551);
xor U3435 (N_3435,N_2727,N_2645);
and U3436 (N_3436,N_2640,N_2651);
nand U3437 (N_3437,N_2996,N_2902);
nand U3438 (N_3438,N_2631,N_2909);
xnor U3439 (N_3439,N_2635,N_2692);
and U3440 (N_3440,N_2809,N_2869);
nor U3441 (N_3441,N_2950,N_2771);
and U3442 (N_3442,N_2871,N_2777);
nor U3443 (N_3443,N_2576,N_2711);
xor U3444 (N_3444,N_2706,N_2611);
nand U3445 (N_3445,N_2600,N_2795);
or U3446 (N_3446,N_2813,N_2590);
nor U3447 (N_3447,N_2923,N_2561);
or U3448 (N_3448,N_2504,N_2971);
and U3449 (N_3449,N_2736,N_2902);
xnor U3450 (N_3450,N_2614,N_2746);
or U3451 (N_3451,N_2621,N_2917);
or U3452 (N_3452,N_2690,N_2607);
xnor U3453 (N_3453,N_2864,N_2950);
or U3454 (N_3454,N_2873,N_2972);
xnor U3455 (N_3455,N_2675,N_2684);
or U3456 (N_3456,N_2570,N_2736);
xor U3457 (N_3457,N_2930,N_2665);
xnor U3458 (N_3458,N_2915,N_2503);
nand U3459 (N_3459,N_2951,N_2554);
and U3460 (N_3460,N_2897,N_2644);
nor U3461 (N_3461,N_2991,N_2985);
nor U3462 (N_3462,N_2705,N_2928);
and U3463 (N_3463,N_2689,N_2533);
or U3464 (N_3464,N_2832,N_2772);
nand U3465 (N_3465,N_2593,N_2707);
or U3466 (N_3466,N_2503,N_2976);
and U3467 (N_3467,N_2771,N_2925);
nand U3468 (N_3468,N_2873,N_2806);
nand U3469 (N_3469,N_2695,N_2691);
or U3470 (N_3470,N_2515,N_2884);
and U3471 (N_3471,N_2883,N_2696);
nor U3472 (N_3472,N_2680,N_2573);
nor U3473 (N_3473,N_2645,N_2702);
or U3474 (N_3474,N_2988,N_2899);
nand U3475 (N_3475,N_2692,N_2753);
nand U3476 (N_3476,N_2732,N_2958);
nand U3477 (N_3477,N_2888,N_2659);
xnor U3478 (N_3478,N_2635,N_2564);
or U3479 (N_3479,N_2598,N_2823);
or U3480 (N_3480,N_2937,N_2790);
and U3481 (N_3481,N_2576,N_2833);
nor U3482 (N_3482,N_2881,N_2904);
or U3483 (N_3483,N_2599,N_2598);
nand U3484 (N_3484,N_2963,N_2806);
and U3485 (N_3485,N_2862,N_2653);
nor U3486 (N_3486,N_2874,N_2780);
and U3487 (N_3487,N_2833,N_2960);
and U3488 (N_3488,N_2825,N_2932);
and U3489 (N_3489,N_2581,N_2514);
nor U3490 (N_3490,N_2905,N_2814);
and U3491 (N_3491,N_2685,N_2976);
or U3492 (N_3492,N_2591,N_2749);
xor U3493 (N_3493,N_2901,N_2624);
xor U3494 (N_3494,N_2939,N_2567);
nor U3495 (N_3495,N_2792,N_2581);
and U3496 (N_3496,N_2880,N_2872);
nand U3497 (N_3497,N_2605,N_2844);
nand U3498 (N_3498,N_2510,N_2943);
nor U3499 (N_3499,N_2721,N_2768);
and U3500 (N_3500,N_3483,N_3008);
nand U3501 (N_3501,N_3127,N_3305);
xor U3502 (N_3502,N_3321,N_3031);
xnor U3503 (N_3503,N_3353,N_3476);
and U3504 (N_3504,N_3465,N_3237);
or U3505 (N_3505,N_3281,N_3067);
and U3506 (N_3506,N_3295,N_3063);
nor U3507 (N_3507,N_3470,N_3482);
and U3508 (N_3508,N_3184,N_3011);
or U3509 (N_3509,N_3021,N_3265);
nor U3510 (N_3510,N_3005,N_3309);
or U3511 (N_3511,N_3491,N_3259);
nand U3512 (N_3512,N_3124,N_3484);
nor U3513 (N_3513,N_3410,N_3350);
or U3514 (N_3514,N_3172,N_3173);
and U3515 (N_3515,N_3022,N_3444);
and U3516 (N_3516,N_3210,N_3039);
xnor U3517 (N_3517,N_3085,N_3159);
nor U3518 (N_3518,N_3406,N_3232);
nor U3519 (N_3519,N_3280,N_3479);
nor U3520 (N_3520,N_3270,N_3264);
nand U3521 (N_3521,N_3017,N_3466);
or U3522 (N_3522,N_3393,N_3004);
nand U3523 (N_3523,N_3453,N_3267);
nand U3524 (N_3524,N_3083,N_3103);
or U3525 (N_3525,N_3474,N_3449);
or U3526 (N_3526,N_3035,N_3409);
and U3527 (N_3527,N_3056,N_3024);
xnor U3528 (N_3528,N_3025,N_3358);
and U3529 (N_3529,N_3020,N_3101);
or U3530 (N_3530,N_3268,N_3219);
and U3531 (N_3531,N_3236,N_3002);
or U3532 (N_3532,N_3390,N_3057);
nor U3533 (N_3533,N_3338,N_3034);
or U3534 (N_3534,N_3272,N_3007);
nor U3535 (N_3535,N_3445,N_3100);
or U3536 (N_3536,N_3239,N_3447);
nor U3537 (N_3537,N_3140,N_3015);
or U3538 (N_3538,N_3443,N_3455);
and U3539 (N_3539,N_3128,N_3274);
nand U3540 (N_3540,N_3045,N_3402);
or U3541 (N_3541,N_3432,N_3260);
nor U3542 (N_3542,N_3388,N_3417);
xor U3543 (N_3543,N_3030,N_3302);
and U3544 (N_3544,N_3171,N_3487);
nand U3545 (N_3545,N_3009,N_3311);
xnor U3546 (N_3546,N_3473,N_3446);
nor U3547 (N_3547,N_3387,N_3069);
or U3548 (N_3548,N_3076,N_3053);
nor U3549 (N_3549,N_3434,N_3122);
or U3550 (N_3550,N_3148,N_3166);
and U3551 (N_3551,N_3425,N_3411);
nand U3552 (N_3552,N_3190,N_3458);
xor U3553 (N_3553,N_3277,N_3316);
or U3554 (N_3554,N_3431,N_3426);
xnor U3555 (N_3555,N_3111,N_3467);
and U3556 (N_3556,N_3208,N_3248);
nand U3557 (N_3557,N_3462,N_3396);
nor U3558 (N_3558,N_3163,N_3217);
and U3559 (N_3559,N_3240,N_3271);
and U3560 (N_3560,N_3322,N_3154);
xnor U3561 (N_3561,N_3399,N_3486);
nor U3562 (N_3562,N_3419,N_3028);
nand U3563 (N_3563,N_3266,N_3206);
and U3564 (N_3564,N_3098,N_3223);
and U3565 (N_3565,N_3414,N_3436);
nand U3566 (N_3566,N_3060,N_3430);
nand U3567 (N_3567,N_3093,N_3359);
nand U3568 (N_3568,N_3125,N_3139);
and U3569 (N_3569,N_3293,N_3253);
nor U3570 (N_3570,N_3241,N_3243);
nand U3571 (N_3571,N_3463,N_3178);
nor U3572 (N_3572,N_3003,N_3318);
or U3573 (N_3573,N_3200,N_3347);
nor U3574 (N_3574,N_3183,N_3228);
and U3575 (N_3575,N_3108,N_3481);
nor U3576 (N_3576,N_3498,N_3335);
xnor U3577 (N_3577,N_3255,N_3055);
and U3578 (N_3578,N_3169,N_3469);
nor U3579 (N_3579,N_3314,N_3349);
nand U3580 (N_3580,N_3168,N_3102);
nor U3581 (N_3581,N_3304,N_3494);
xor U3582 (N_3582,N_3164,N_3459);
and U3583 (N_3583,N_3294,N_3418);
nor U3584 (N_3584,N_3084,N_3475);
nor U3585 (N_3585,N_3114,N_3152);
xor U3586 (N_3586,N_3218,N_3392);
nand U3587 (N_3587,N_3221,N_3345);
xnor U3588 (N_3588,N_3010,N_3119);
and U3589 (N_3589,N_3420,N_3279);
nand U3590 (N_3590,N_3497,N_3339);
nand U3591 (N_3591,N_3061,N_3456);
or U3592 (N_3592,N_3105,N_3049);
nor U3593 (N_3593,N_3068,N_3450);
and U3594 (N_3594,N_3263,N_3495);
or U3595 (N_3595,N_3027,N_3110);
xnor U3596 (N_3596,N_3251,N_3033);
and U3597 (N_3597,N_3472,N_3023);
xnor U3598 (N_3598,N_3401,N_3234);
nor U3599 (N_3599,N_3386,N_3300);
and U3600 (N_3600,N_3029,N_3046);
nor U3601 (N_3601,N_3136,N_3220);
xnor U3602 (N_3602,N_3365,N_3490);
and U3603 (N_3603,N_3192,N_3207);
nand U3604 (N_3604,N_3079,N_3161);
or U3605 (N_3605,N_3089,N_3073);
or U3606 (N_3606,N_3433,N_3000);
xor U3607 (N_3607,N_3372,N_3205);
nand U3608 (N_3608,N_3346,N_3117);
and U3609 (N_3609,N_3341,N_3363);
nor U3610 (N_3610,N_3202,N_3109);
xor U3611 (N_3611,N_3471,N_3429);
nand U3612 (N_3612,N_3229,N_3249);
nand U3613 (N_3613,N_3325,N_3222);
nand U3614 (N_3614,N_3397,N_3216);
nand U3615 (N_3615,N_3380,N_3242);
nor U3616 (N_3616,N_3016,N_3323);
or U3617 (N_3617,N_3224,N_3158);
nand U3618 (N_3618,N_3464,N_3231);
nand U3619 (N_3619,N_3047,N_3080);
and U3620 (N_3620,N_3400,N_3442);
xnor U3621 (N_3621,N_3106,N_3367);
xor U3622 (N_3622,N_3489,N_3308);
nand U3623 (N_3623,N_3330,N_3340);
nor U3624 (N_3624,N_3496,N_3037);
or U3625 (N_3625,N_3376,N_3099);
and U3626 (N_3626,N_3226,N_3375);
nand U3627 (N_3627,N_3227,N_3317);
nand U3628 (N_3628,N_3097,N_3132);
xnor U3629 (N_3629,N_3160,N_3273);
or U3630 (N_3630,N_3478,N_3278);
nand U3631 (N_3631,N_3187,N_3048);
and U3632 (N_3632,N_3062,N_3120);
and U3633 (N_3633,N_3324,N_3452);
and U3634 (N_3634,N_3146,N_3343);
and U3635 (N_3635,N_3040,N_3244);
nand U3636 (N_3636,N_3195,N_3041);
nor U3637 (N_3637,N_3312,N_3213);
and U3638 (N_3638,N_3329,N_3189);
or U3639 (N_3639,N_3403,N_3215);
and U3640 (N_3640,N_3014,N_3133);
or U3641 (N_3641,N_3082,N_3254);
and U3642 (N_3642,N_3269,N_3121);
or U3643 (N_3643,N_3356,N_3332);
or U3644 (N_3644,N_3175,N_3174);
and U3645 (N_3645,N_3460,N_3369);
and U3646 (N_3646,N_3019,N_3135);
nand U3647 (N_3647,N_3087,N_3246);
or U3648 (N_3648,N_3182,N_3112);
and U3649 (N_3649,N_3282,N_3129);
and U3650 (N_3650,N_3437,N_3477);
nor U3651 (N_3651,N_3233,N_3147);
and U3652 (N_3652,N_3247,N_3032);
nand U3653 (N_3653,N_3156,N_3485);
nand U3654 (N_3654,N_3198,N_3499);
nand U3655 (N_3655,N_3086,N_3492);
nand U3656 (N_3656,N_3179,N_3299);
xnor U3657 (N_3657,N_3404,N_3395);
nand U3658 (N_3658,N_3131,N_3012);
and U3659 (N_3659,N_3326,N_3454);
nand U3660 (N_3660,N_3275,N_3252);
or U3661 (N_3661,N_3351,N_3026);
nand U3662 (N_3662,N_3389,N_3370);
nand U3663 (N_3663,N_3310,N_3036);
or U3664 (N_3664,N_3371,N_3075);
or U3665 (N_3665,N_3107,N_3385);
nand U3666 (N_3666,N_3441,N_3438);
nor U3667 (N_3667,N_3336,N_3188);
nand U3668 (N_3668,N_3448,N_3289);
and U3669 (N_3669,N_3211,N_3151);
nand U3670 (N_3670,N_3368,N_3081);
or U3671 (N_3671,N_3285,N_3162);
or U3672 (N_3672,N_3394,N_3126);
or U3673 (N_3673,N_3145,N_3209);
and U3674 (N_3674,N_3422,N_3071);
or U3675 (N_3675,N_3078,N_3018);
nor U3676 (N_3676,N_3288,N_3257);
or U3677 (N_3677,N_3451,N_3043);
nor U3678 (N_3678,N_3165,N_3428);
xor U3679 (N_3679,N_3423,N_3167);
nand U3680 (N_3680,N_3070,N_3230);
nor U3681 (N_3681,N_3439,N_3261);
nand U3682 (N_3682,N_3123,N_3357);
nand U3683 (N_3683,N_3201,N_3134);
xor U3684 (N_3684,N_3421,N_3424);
or U3685 (N_3685,N_3348,N_3342);
nor U3686 (N_3686,N_3203,N_3096);
and U3687 (N_3687,N_3225,N_3362);
nand U3688 (N_3688,N_3006,N_3276);
nand U3689 (N_3689,N_3170,N_3292);
nand U3690 (N_3690,N_3262,N_3435);
or U3691 (N_3691,N_3191,N_3290);
and U3692 (N_3692,N_3398,N_3457);
nor U3693 (N_3693,N_3177,N_3383);
or U3694 (N_3694,N_3149,N_3141);
or U3695 (N_3695,N_3050,N_3307);
nor U3696 (N_3696,N_3407,N_3258);
nor U3697 (N_3697,N_3042,N_3256);
nand U3698 (N_3698,N_3153,N_3104);
or U3699 (N_3699,N_3077,N_3118);
xnor U3700 (N_3700,N_3144,N_3058);
nor U3701 (N_3701,N_3038,N_3091);
or U3702 (N_3702,N_3327,N_3354);
nand U3703 (N_3703,N_3095,N_3405);
or U3704 (N_3704,N_3142,N_3361);
nand U3705 (N_3705,N_3378,N_3374);
nand U3706 (N_3706,N_3296,N_3137);
nor U3707 (N_3707,N_3054,N_3301);
nand U3708 (N_3708,N_3352,N_3157);
and U3709 (N_3709,N_3130,N_3072);
and U3710 (N_3710,N_3059,N_3488);
and U3711 (N_3711,N_3051,N_3013);
or U3712 (N_3712,N_3331,N_3180);
or U3713 (N_3713,N_3364,N_3194);
nor U3714 (N_3714,N_3116,N_3186);
and U3715 (N_3715,N_3313,N_3287);
or U3716 (N_3716,N_3052,N_3360);
nand U3717 (N_3717,N_3328,N_3344);
nand U3718 (N_3718,N_3150,N_3212);
xor U3719 (N_3719,N_3238,N_3427);
xnor U3720 (N_3720,N_3416,N_3379);
nand U3721 (N_3721,N_3138,N_3065);
nor U3722 (N_3722,N_3355,N_3245);
and U3723 (N_3723,N_3381,N_3286);
and U3724 (N_3724,N_3382,N_3250);
and U3725 (N_3725,N_3064,N_3283);
and U3726 (N_3726,N_3001,N_3413);
nand U3727 (N_3727,N_3066,N_3440);
xor U3728 (N_3728,N_3319,N_3408);
nor U3729 (N_3729,N_3199,N_3196);
nor U3730 (N_3730,N_3143,N_3204);
nand U3731 (N_3731,N_3155,N_3333);
xnor U3732 (N_3732,N_3094,N_3115);
and U3733 (N_3733,N_3181,N_3092);
nor U3734 (N_3734,N_3384,N_3088);
xor U3735 (N_3735,N_3214,N_3176);
and U3736 (N_3736,N_3185,N_3377);
xor U3737 (N_3737,N_3297,N_3303);
and U3738 (N_3738,N_3235,N_3315);
and U3739 (N_3739,N_3461,N_3480);
nor U3740 (N_3740,N_3415,N_3298);
xor U3741 (N_3741,N_3373,N_3412);
nor U3742 (N_3742,N_3334,N_3468);
nand U3743 (N_3743,N_3090,N_3391);
and U3744 (N_3744,N_3306,N_3193);
or U3745 (N_3745,N_3366,N_3337);
or U3746 (N_3746,N_3493,N_3044);
xor U3747 (N_3747,N_3291,N_3284);
and U3748 (N_3748,N_3197,N_3074);
and U3749 (N_3749,N_3113,N_3320);
or U3750 (N_3750,N_3034,N_3496);
xor U3751 (N_3751,N_3143,N_3317);
or U3752 (N_3752,N_3352,N_3342);
nand U3753 (N_3753,N_3090,N_3191);
nor U3754 (N_3754,N_3456,N_3437);
xnor U3755 (N_3755,N_3395,N_3440);
nor U3756 (N_3756,N_3012,N_3010);
xnor U3757 (N_3757,N_3429,N_3491);
or U3758 (N_3758,N_3033,N_3026);
or U3759 (N_3759,N_3480,N_3469);
or U3760 (N_3760,N_3401,N_3338);
or U3761 (N_3761,N_3084,N_3069);
nor U3762 (N_3762,N_3021,N_3161);
xor U3763 (N_3763,N_3273,N_3083);
and U3764 (N_3764,N_3285,N_3488);
nor U3765 (N_3765,N_3423,N_3425);
or U3766 (N_3766,N_3478,N_3252);
nor U3767 (N_3767,N_3037,N_3073);
nand U3768 (N_3768,N_3091,N_3310);
or U3769 (N_3769,N_3273,N_3397);
xnor U3770 (N_3770,N_3402,N_3218);
xor U3771 (N_3771,N_3298,N_3202);
or U3772 (N_3772,N_3055,N_3128);
nand U3773 (N_3773,N_3212,N_3013);
nor U3774 (N_3774,N_3257,N_3117);
nand U3775 (N_3775,N_3245,N_3192);
nand U3776 (N_3776,N_3240,N_3028);
nor U3777 (N_3777,N_3401,N_3133);
and U3778 (N_3778,N_3299,N_3435);
nor U3779 (N_3779,N_3215,N_3246);
and U3780 (N_3780,N_3351,N_3496);
and U3781 (N_3781,N_3480,N_3326);
nor U3782 (N_3782,N_3075,N_3167);
nand U3783 (N_3783,N_3291,N_3259);
or U3784 (N_3784,N_3211,N_3227);
or U3785 (N_3785,N_3455,N_3237);
nor U3786 (N_3786,N_3232,N_3214);
nand U3787 (N_3787,N_3486,N_3016);
nand U3788 (N_3788,N_3121,N_3443);
nand U3789 (N_3789,N_3087,N_3471);
or U3790 (N_3790,N_3066,N_3160);
xor U3791 (N_3791,N_3388,N_3194);
nor U3792 (N_3792,N_3179,N_3150);
and U3793 (N_3793,N_3270,N_3372);
and U3794 (N_3794,N_3014,N_3464);
nand U3795 (N_3795,N_3427,N_3383);
and U3796 (N_3796,N_3334,N_3160);
nor U3797 (N_3797,N_3057,N_3185);
nand U3798 (N_3798,N_3254,N_3138);
nand U3799 (N_3799,N_3119,N_3482);
nor U3800 (N_3800,N_3394,N_3488);
or U3801 (N_3801,N_3232,N_3057);
and U3802 (N_3802,N_3013,N_3325);
nand U3803 (N_3803,N_3436,N_3291);
or U3804 (N_3804,N_3422,N_3155);
nand U3805 (N_3805,N_3289,N_3198);
xnor U3806 (N_3806,N_3149,N_3271);
and U3807 (N_3807,N_3397,N_3204);
nand U3808 (N_3808,N_3006,N_3138);
nand U3809 (N_3809,N_3285,N_3212);
xnor U3810 (N_3810,N_3363,N_3061);
or U3811 (N_3811,N_3320,N_3044);
xnor U3812 (N_3812,N_3172,N_3082);
nor U3813 (N_3813,N_3070,N_3475);
xor U3814 (N_3814,N_3200,N_3028);
xnor U3815 (N_3815,N_3213,N_3338);
nand U3816 (N_3816,N_3317,N_3449);
or U3817 (N_3817,N_3282,N_3275);
or U3818 (N_3818,N_3311,N_3457);
nand U3819 (N_3819,N_3367,N_3297);
or U3820 (N_3820,N_3131,N_3068);
nor U3821 (N_3821,N_3254,N_3188);
and U3822 (N_3822,N_3436,N_3141);
nand U3823 (N_3823,N_3113,N_3145);
nor U3824 (N_3824,N_3203,N_3178);
nand U3825 (N_3825,N_3238,N_3160);
and U3826 (N_3826,N_3476,N_3440);
nand U3827 (N_3827,N_3079,N_3338);
or U3828 (N_3828,N_3047,N_3351);
xor U3829 (N_3829,N_3245,N_3042);
nor U3830 (N_3830,N_3295,N_3335);
nor U3831 (N_3831,N_3318,N_3468);
nand U3832 (N_3832,N_3204,N_3025);
nor U3833 (N_3833,N_3275,N_3496);
and U3834 (N_3834,N_3144,N_3383);
or U3835 (N_3835,N_3180,N_3496);
nand U3836 (N_3836,N_3385,N_3495);
nor U3837 (N_3837,N_3424,N_3438);
or U3838 (N_3838,N_3215,N_3247);
nand U3839 (N_3839,N_3266,N_3346);
and U3840 (N_3840,N_3338,N_3086);
nand U3841 (N_3841,N_3309,N_3327);
or U3842 (N_3842,N_3093,N_3450);
xor U3843 (N_3843,N_3035,N_3241);
and U3844 (N_3844,N_3395,N_3085);
and U3845 (N_3845,N_3285,N_3293);
nor U3846 (N_3846,N_3244,N_3310);
nand U3847 (N_3847,N_3147,N_3439);
nor U3848 (N_3848,N_3287,N_3182);
nand U3849 (N_3849,N_3422,N_3429);
xor U3850 (N_3850,N_3081,N_3456);
nand U3851 (N_3851,N_3025,N_3398);
nand U3852 (N_3852,N_3460,N_3179);
nand U3853 (N_3853,N_3269,N_3275);
nand U3854 (N_3854,N_3021,N_3038);
nor U3855 (N_3855,N_3221,N_3208);
nor U3856 (N_3856,N_3234,N_3345);
xor U3857 (N_3857,N_3029,N_3325);
nand U3858 (N_3858,N_3483,N_3332);
nand U3859 (N_3859,N_3165,N_3290);
nor U3860 (N_3860,N_3183,N_3440);
nor U3861 (N_3861,N_3249,N_3395);
and U3862 (N_3862,N_3004,N_3339);
nand U3863 (N_3863,N_3338,N_3166);
nand U3864 (N_3864,N_3302,N_3441);
nor U3865 (N_3865,N_3383,N_3412);
or U3866 (N_3866,N_3261,N_3155);
and U3867 (N_3867,N_3305,N_3386);
nor U3868 (N_3868,N_3441,N_3142);
nand U3869 (N_3869,N_3172,N_3248);
or U3870 (N_3870,N_3431,N_3415);
nand U3871 (N_3871,N_3365,N_3320);
or U3872 (N_3872,N_3323,N_3297);
and U3873 (N_3873,N_3030,N_3004);
xor U3874 (N_3874,N_3489,N_3179);
nor U3875 (N_3875,N_3477,N_3220);
and U3876 (N_3876,N_3197,N_3160);
and U3877 (N_3877,N_3162,N_3441);
nor U3878 (N_3878,N_3387,N_3423);
or U3879 (N_3879,N_3139,N_3219);
xor U3880 (N_3880,N_3369,N_3294);
and U3881 (N_3881,N_3408,N_3068);
and U3882 (N_3882,N_3429,N_3144);
nor U3883 (N_3883,N_3169,N_3481);
and U3884 (N_3884,N_3410,N_3031);
and U3885 (N_3885,N_3435,N_3487);
or U3886 (N_3886,N_3364,N_3220);
or U3887 (N_3887,N_3359,N_3275);
nor U3888 (N_3888,N_3132,N_3109);
or U3889 (N_3889,N_3400,N_3312);
and U3890 (N_3890,N_3008,N_3232);
xor U3891 (N_3891,N_3271,N_3386);
or U3892 (N_3892,N_3067,N_3066);
xor U3893 (N_3893,N_3140,N_3217);
nor U3894 (N_3894,N_3296,N_3057);
and U3895 (N_3895,N_3458,N_3015);
nand U3896 (N_3896,N_3117,N_3367);
xor U3897 (N_3897,N_3174,N_3158);
xor U3898 (N_3898,N_3453,N_3050);
or U3899 (N_3899,N_3127,N_3466);
nand U3900 (N_3900,N_3461,N_3081);
nand U3901 (N_3901,N_3444,N_3216);
and U3902 (N_3902,N_3081,N_3036);
nand U3903 (N_3903,N_3344,N_3036);
or U3904 (N_3904,N_3037,N_3375);
and U3905 (N_3905,N_3355,N_3208);
or U3906 (N_3906,N_3446,N_3265);
nor U3907 (N_3907,N_3493,N_3465);
or U3908 (N_3908,N_3407,N_3003);
and U3909 (N_3909,N_3262,N_3131);
xnor U3910 (N_3910,N_3159,N_3187);
or U3911 (N_3911,N_3383,N_3408);
or U3912 (N_3912,N_3413,N_3037);
nor U3913 (N_3913,N_3243,N_3417);
and U3914 (N_3914,N_3499,N_3275);
and U3915 (N_3915,N_3391,N_3471);
nor U3916 (N_3916,N_3126,N_3147);
nor U3917 (N_3917,N_3329,N_3058);
nor U3918 (N_3918,N_3450,N_3369);
and U3919 (N_3919,N_3306,N_3124);
or U3920 (N_3920,N_3488,N_3071);
and U3921 (N_3921,N_3273,N_3441);
and U3922 (N_3922,N_3190,N_3454);
or U3923 (N_3923,N_3375,N_3442);
and U3924 (N_3924,N_3144,N_3101);
xor U3925 (N_3925,N_3297,N_3173);
or U3926 (N_3926,N_3258,N_3425);
nand U3927 (N_3927,N_3226,N_3391);
nor U3928 (N_3928,N_3364,N_3373);
nand U3929 (N_3929,N_3298,N_3492);
and U3930 (N_3930,N_3123,N_3040);
nor U3931 (N_3931,N_3078,N_3054);
nor U3932 (N_3932,N_3035,N_3398);
or U3933 (N_3933,N_3061,N_3117);
and U3934 (N_3934,N_3466,N_3137);
nor U3935 (N_3935,N_3092,N_3199);
nor U3936 (N_3936,N_3451,N_3290);
xor U3937 (N_3937,N_3082,N_3499);
or U3938 (N_3938,N_3060,N_3434);
nand U3939 (N_3939,N_3026,N_3129);
and U3940 (N_3940,N_3341,N_3009);
and U3941 (N_3941,N_3489,N_3464);
or U3942 (N_3942,N_3062,N_3431);
and U3943 (N_3943,N_3497,N_3414);
nor U3944 (N_3944,N_3477,N_3156);
xor U3945 (N_3945,N_3272,N_3419);
or U3946 (N_3946,N_3135,N_3025);
nand U3947 (N_3947,N_3097,N_3413);
nand U3948 (N_3948,N_3034,N_3326);
or U3949 (N_3949,N_3301,N_3039);
nor U3950 (N_3950,N_3046,N_3270);
nand U3951 (N_3951,N_3180,N_3060);
nor U3952 (N_3952,N_3037,N_3151);
nand U3953 (N_3953,N_3409,N_3007);
xnor U3954 (N_3954,N_3277,N_3410);
and U3955 (N_3955,N_3351,N_3176);
xor U3956 (N_3956,N_3102,N_3157);
or U3957 (N_3957,N_3367,N_3052);
nor U3958 (N_3958,N_3129,N_3198);
or U3959 (N_3959,N_3285,N_3306);
xor U3960 (N_3960,N_3187,N_3389);
or U3961 (N_3961,N_3381,N_3094);
nand U3962 (N_3962,N_3264,N_3432);
xnor U3963 (N_3963,N_3081,N_3088);
nor U3964 (N_3964,N_3149,N_3015);
nor U3965 (N_3965,N_3483,N_3076);
and U3966 (N_3966,N_3403,N_3190);
nor U3967 (N_3967,N_3386,N_3234);
and U3968 (N_3968,N_3462,N_3269);
and U3969 (N_3969,N_3203,N_3479);
and U3970 (N_3970,N_3122,N_3225);
nand U3971 (N_3971,N_3375,N_3192);
nor U3972 (N_3972,N_3089,N_3164);
nor U3973 (N_3973,N_3217,N_3043);
nor U3974 (N_3974,N_3180,N_3178);
and U3975 (N_3975,N_3116,N_3494);
and U3976 (N_3976,N_3263,N_3229);
nand U3977 (N_3977,N_3241,N_3409);
nor U3978 (N_3978,N_3267,N_3123);
and U3979 (N_3979,N_3175,N_3340);
nand U3980 (N_3980,N_3037,N_3137);
xor U3981 (N_3981,N_3201,N_3249);
xor U3982 (N_3982,N_3151,N_3414);
and U3983 (N_3983,N_3343,N_3284);
and U3984 (N_3984,N_3076,N_3452);
nand U3985 (N_3985,N_3271,N_3477);
and U3986 (N_3986,N_3176,N_3194);
nor U3987 (N_3987,N_3395,N_3012);
nor U3988 (N_3988,N_3302,N_3281);
nor U3989 (N_3989,N_3322,N_3275);
nor U3990 (N_3990,N_3298,N_3300);
nand U3991 (N_3991,N_3495,N_3198);
and U3992 (N_3992,N_3214,N_3373);
and U3993 (N_3993,N_3425,N_3463);
nor U3994 (N_3994,N_3392,N_3220);
nor U3995 (N_3995,N_3494,N_3140);
nor U3996 (N_3996,N_3215,N_3417);
nand U3997 (N_3997,N_3291,N_3184);
nand U3998 (N_3998,N_3416,N_3027);
nor U3999 (N_3999,N_3213,N_3076);
or U4000 (N_4000,N_3746,N_3987);
nor U4001 (N_4001,N_3718,N_3971);
and U4002 (N_4002,N_3548,N_3918);
or U4003 (N_4003,N_3824,N_3635);
and U4004 (N_4004,N_3964,N_3711);
nor U4005 (N_4005,N_3776,N_3917);
or U4006 (N_4006,N_3881,N_3817);
xor U4007 (N_4007,N_3965,N_3617);
nor U4008 (N_4008,N_3590,N_3579);
and U4009 (N_4009,N_3603,N_3594);
nor U4010 (N_4010,N_3688,N_3840);
or U4011 (N_4011,N_3736,N_3831);
nor U4012 (N_4012,N_3519,N_3937);
and U4013 (N_4013,N_3698,N_3611);
xor U4014 (N_4014,N_3798,N_3605);
or U4015 (N_4015,N_3753,N_3620);
nand U4016 (N_4016,N_3695,N_3512);
xor U4017 (N_4017,N_3810,N_3511);
nor U4018 (N_4018,N_3939,N_3676);
and U4019 (N_4019,N_3781,N_3959);
nor U4020 (N_4020,N_3822,N_3670);
nand U4021 (N_4021,N_3503,N_3516);
or U4022 (N_4022,N_3553,N_3575);
nand U4023 (N_4023,N_3991,N_3581);
nor U4024 (N_4024,N_3597,N_3802);
nand U4025 (N_4025,N_3535,N_3838);
or U4026 (N_4026,N_3723,N_3812);
and U4027 (N_4027,N_3685,N_3513);
or U4028 (N_4028,N_3976,N_3880);
nor U4029 (N_4029,N_3515,N_3910);
or U4030 (N_4030,N_3842,N_3848);
nand U4031 (N_4031,N_3924,N_3993);
xnor U4032 (N_4032,N_3803,N_3945);
or U4033 (N_4033,N_3889,N_3554);
xnor U4034 (N_4034,N_3958,N_3974);
nor U4035 (N_4035,N_3702,N_3639);
nor U4036 (N_4036,N_3556,N_3830);
or U4037 (N_4037,N_3806,N_3844);
and U4038 (N_4038,N_3829,N_3808);
or U4039 (N_4039,N_3867,N_3893);
nor U4040 (N_4040,N_3645,N_3518);
nand U4041 (N_4041,N_3583,N_3841);
and U4042 (N_4042,N_3853,N_3782);
xnor U4043 (N_4043,N_3527,N_3750);
nor U4044 (N_4044,N_3682,N_3681);
and U4045 (N_4045,N_3843,N_3788);
nor U4046 (N_4046,N_3668,N_3962);
nand U4047 (N_4047,N_3877,N_3538);
xor U4048 (N_4048,N_3957,N_3664);
nor U4049 (N_4049,N_3858,N_3839);
xor U4050 (N_4050,N_3805,N_3759);
nand U4051 (N_4051,N_3978,N_3735);
or U4052 (N_4052,N_3992,N_3891);
nor U4053 (N_4053,N_3628,N_3607);
nand U4054 (N_4054,N_3989,N_3618);
and U4055 (N_4055,N_3821,N_3592);
or U4056 (N_4056,N_3990,N_3689);
or U4057 (N_4057,N_3526,N_3561);
and U4058 (N_4058,N_3567,N_3994);
nor U4059 (N_4059,N_3565,N_3784);
and U4060 (N_4060,N_3970,N_3814);
or U4061 (N_4061,N_3520,N_3796);
nand U4062 (N_4062,N_3525,N_3551);
and U4063 (N_4063,N_3981,N_3609);
or U4064 (N_4064,N_3675,N_3799);
and U4065 (N_4065,N_3537,N_3601);
or U4066 (N_4066,N_3623,N_3598);
and U4067 (N_4067,N_3568,N_3986);
nor U4068 (N_4068,N_3789,N_3602);
or U4069 (N_4069,N_3774,N_3655);
or U4070 (N_4070,N_3928,N_3919);
or U4071 (N_4071,N_3783,N_3902);
nor U4072 (N_4072,N_3706,N_3778);
or U4073 (N_4073,N_3524,N_3818);
or U4074 (N_4074,N_3528,N_3543);
nor U4075 (N_4075,N_3973,N_3522);
nand U4076 (N_4076,N_3564,N_3773);
and U4077 (N_4077,N_3815,N_3691);
xnor U4078 (N_4078,N_3577,N_3916);
or U4079 (N_4079,N_3825,N_3813);
nand U4080 (N_4080,N_3909,N_3758);
xor U4081 (N_4081,N_3947,N_3741);
nor U4082 (N_4082,N_3604,N_3876);
nand U4083 (N_4083,N_3755,N_3517);
and U4084 (N_4084,N_3612,N_3828);
nand U4085 (N_4085,N_3610,N_3762);
or U4086 (N_4086,N_3508,N_3864);
nor U4087 (N_4087,N_3509,N_3627);
and U4088 (N_4088,N_3638,N_3887);
or U4089 (N_4089,N_3930,N_3679);
nand U4090 (N_4090,N_3692,N_3683);
and U4091 (N_4091,N_3742,N_3576);
and U4092 (N_4092,N_3878,N_3866);
and U4093 (N_4093,N_3927,N_3745);
and U4094 (N_4094,N_3795,N_3785);
nand U4095 (N_4095,N_3644,N_3980);
and U4096 (N_4096,N_3975,N_3640);
or U4097 (N_4097,N_3729,N_3772);
or U4098 (N_4098,N_3665,N_3642);
or U4099 (N_4099,N_3500,N_3501);
xor U4100 (N_4100,N_3673,N_3851);
nand U4101 (N_4101,N_3832,N_3700);
nand U4102 (N_4102,N_3854,N_3787);
xnor U4103 (N_4103,N_3558,N_3716);
nand U4104 (N_4104,N_3633,N_3580);
or U4105 (N_4105,N_3775,N_3827);
nor U4106 (N_4106,N_3862,N_3714);
or U4107 (N_4107,N_3699,N_3907);
nor U4108 (N_4108,N_3949,N_3906);
nand U4109 (N_4109,N_3649,N_3593);
nand U4110 (N_4110,N_3896,N_3748);
nand U4111 (N_4111,N_3826,N_3613);
nor U4112 (N_4112,N_3721,N_3886);
nand U4113 (N_4113,N_3935,N_3710);
nand U4114 (N_4114,N_3544,N_3911);
nor U4115 (N_4115,N_3730,N_3940);
xor U4116 (N_4116,N_3868,N_3760);
nand U4117 (N_4117,N_3571,N_3632);
nor U4118 (N_4118,N_3800,N_3652);
or U4119 (N_4119,N_3658,N_3953);
nor U4120 (N_4120,N_3703,N_3629);
and U4121 (N_4121,N_3534,N_3694);
and U4122 (N_4122,N_3983,N_3636);
nor U4123 (N_4123,N_3715,N_3977);
or U4124 (N_4124,N_3897,N_3726);
and U4125 (N_4125,N_3969,N_3619);
and U4126 (N_4126,N_3728,N_3797);
nor U4127 (N_4127,N_3546,N_3532);
nand U4128 (N_4128,N_3834,N_3733);
nand U4129 (N_4129,N_3861,N_3540);
and U4130 (N_4130,N_3662,N_3545);
xnor U4131 (N_4131,N_3998,N_3560);
nand U4132 (N_4132,N_3739,N_3536);
nand U4133 (N_4133,N_3942,N_3510);
nand U4134 (N_4134,N_3616,N_3740);
nand U4135 (N_4135,N_3771,N_3634);
or U4136 (N_4136,N_3988,N_3563);
nor U4137 (N_4137,N_3712,N_3530);
nand U4138 (N_4138,N_3624,N_3719);
nor U4139 (N_4139,N_3856,N_3833);
or U4140 (N_4140,N_3790,N_3550);
or U4141 (N_4141,N_3879,N_3898);
nor U4142 (N_4142,N_3967,N_3650);
nand U4143 (N_4143,N_3587,N_3859);
or U4144 (N_4144,N_3722,N_3562);
or U4145 (N_4145,N_3816,N_3849);
or U4146 (N_4146,N_3539,N_3667);
nand U4147 (N_4147,N_3621,N_3903);
and U4148 (N_4148,N_3677,N_3908);
or U4149 (N_4149,N_3531,N_3507);
or U4150 (N_4150,N_3865,N_3523);
nor U4151 (N_4151,N_3654,N_3643);
nor U4152 (N_4152,N_3696,N_3572);
nand U4153 (N_4153,N_3820,N_3870);
or U4154 (N_4154,N_3678,N_3653);
and U4155 (N_4155,N_3705,N_3837);
nand U4156 (N_4156,N_3555,N_3549);
or U4157 (N_4157,N_3690,N_3920);
or U4158 (N_4158,N_3573,N_3595);
or U4159 (N_4159,N_3954,N_3857);
or U4160 (N_4160,N_3926,N_3660);
or U4161 (N_4161,N_3923,N_3894);
nand U4162 (N_4162,N_3960,N_3985);
nand U4163 (N_4163,N_3709,N_3780);
and U4164 (N_4164,N_3769,N_3727);
or U4165 (N_4165,N_3899,N_3765);
nor U4166 (N_4166,N_3591,N_3938);
nor U4167 (N_4167,N_3669,N_3914);
and U4168 (N_4168,N_3836,N_3997);
nand U4169 (N_4169,N_3596,N_3845);
or U4170 (N_4170,N_3751,N_3557);
or U4171 (N_4171,N_3925,N_3871);
nand U4172 (N_4172,N_3514,N_3589);
xor U4173 (N_4173,N_3885,N_3793);
xnor U4174 (N_4174,N_3811,N_3541);
nand U4175 (N_4175,N_3763,N_3946);
or U4176 (N_4176,N_3963,N_3863);
nand U4177 (N_4177,N_3804,N_3666);
nor U4178 (N_4178,N_3888,N_3529);
or U4179 (N_4179,N_3873,N_3651);
nor U4180 (N_4180,N_3948,N_3941);
nor U4181 (N_4181,N_3955,N_3671);
xor U4182 (N_4182,N_3892,N_3521);
nand U4183 (N_4183,N_3757,N_3752);
nor U4184 (N_4184,N_3704,N_3850);
nor U4185 (N_4185,N_3770,N_3578);
or U4186 (N_4186,N_3625,N_3582);
nor U4187 (N_4187,N_3913,N_3630);
or U4188 (N_4188,N_3982,N_3717);
nor U4189 (N_4189,N_3961,N_3855);
xnor U4190 (N_4190,N_3950,N_3995);
and U4191 (N_4191,N_3852,N_3932);
or U4192 (N_4192,N_3943,N_3792);
and U4193 (N_4193,N_3807,N_3713);
and U4194 (N_4194,N_3749,N_3966);
xnor U4195 (N_4195,N_3884,N_3883);
nor U4196 (N_4196,N_3502,N_3680);
and U4197 (N_4197,N_3707,N_3761);
or U4198 (N_4198,N_3606,N_3933);
and U4199 (N_4199,N_3767,N_3929);
and U4200 (N_4200,N_3697,N_3738);
nand U4201 (N_4201,N_3979,N_3701);
nand U4202 (N_4202,N_3584,N_3744);
or U4203 (N_4203,N_3659,N_3922);
nand U4204 (N_4204,N_3984,N_3779);
or U4205 (N_4205,N_3794,N_3835);
xor U4206 (N_4206,N_3777,N_3956);
nor U4207 (N_4207,N_3951,N_3934);
nand U4208 (N_4208,N_3552,N_3972);
nor U4209 (N_4209,N_3674,N_3641);
nor U4210 (N_4210,N_3687,N_3900);
or U4211 (N_4211,N_3895,N_3686);
and U4212 (N_4212,N_3872,N_3720);
or U4213 (N_4213,N_3614,N_3754);
nor U4214 (N_4214,N_3952,N_3725);
nand U4215 (N_4215,N_3505,N_3766);
nor U4216 (N_4216,N_3743,N_3823);
nand U4217 (N_4217,N_3631,N_3574);
and U4218 (N_4218,N_3882,N_3747);
nor U4219 (N_4219,N_3559,N_3569);
and U4220 (N_4220,N_3566,N_3999);
nand U4221 (N_4221,N_3542,N_3615);
and U4222 (N_4222,N_3732,N_3648);
nand U4223 (N_4223,N_3904,N_3901);
nand U4224 (N_4224,N_3570,N_3708);
nand U4225 (N_4225,N_3921,N_3847);
nand U4226 (N_4226,N_3905,N_3600);
xor U4227 (N_4227,N_3869,N_3936);
nor U4228 (N_4228,N_3809,N_3506);
and U4229 (N_4229,N_3846,N_3599);
nand U4230 (N_4230,N_3915,N_3533);
nand U4231 (N_4231,N_3874,N_3622);
or U4232 (N_4232,N_3646,N_3944);
or U4233 (N_4233,N_3586,N_3731);
xnor U4234 (N_4234,N_3663,N_3860);
nor U4235 (N_4235,N_3768,N_3724);
nand U4236 (N_4236,N_3672,N_3588);
nand U4237 (N_4237,N_3637,N_3756);
nor U4238 (N_4238,N_3657,N_3764);
and U4239 (N_4239,N_3734,N_3875);
or U4240 (N_4240,N_3547,N_3656);
or U4241 (N_4241,N_3693,N_3737);
nand U4242 (N_4242,N_3912,N_3931);
xnor U4243 (N_4243,N_3801,N_3504);
nand U4244 (N_4244,N_3968,N_3996);
and U4245 (N_4245,N_3585,N_3890);
nand U4246 (N_4246,N_3626,N_3819);
or U4247 (N_4247,N_3661,N_3791);
nor U4248 (N_4248,N_3684,N_3647);
or U4249 (N_4249,N_3608,N_3786);
nor U4250 (N_4250,N_3601,N_3795);
or U4251 (N_4251,N_3837,N_3574);
or U4252 (N_4252,N_3560,N_3527);
nand U4253 (N_4253,N_3530,N_3917);
nor U4254 (N_4254,N_3602,N_3946);
or U4255 (N_4255,N_3926,N_3836);
and U4256 (N_4256,N_3945,N_3987);
nor U4257 (N_4257,N_3516,N_3906);
nor U4258 (N_4258,N_3581,N_3658);
or U4259 (N_4259,N_3774,N_3913);
and U4260 (N_4260,N_3643,N_3793);
nand U4261 (N_4261,N_3932,N_3661);
xor U4262 (N_4262,N_3519,N_3943);
or U4263 (N_4263,N_3738,N_3907);
nor U4264 (N_4264,N_3807,N_3701);
nand U4265 (N_4265,N_3565,N_3900);
nor U4266 (N_4266,N_3733,N_3840);
and U4267 (N_4267,N_3715,N_3899);
nor U4268 (N_4268,N_3874,N_3644);
nand U4269 (N_4269,N_3597,N_3831);
or U4270 (N_4270,N_3663,N_3883);
xor U4271 (N_4271,N_3709,N_3731);
nand U4272 (N_4272,N_3775,N_3837);
nand U4273 (N_4273,N_3635,N_3804);
nor U4274 (N_4274,N_3888,N_3862);
nand U4275 (N_4275,N_3735,N_3966);
and U4276 (N_4276,N_3837,N_3673);
nand U4277 (N_4277,N_3867,N_3788);
nand U4278 (N_4278,N_3765,N_3912);
or U4279 (N_4279,N_3724,N_3728);
nor U4280 (N_4280,N_3635,N_3746);
and U4281 (N_4281,N_3847,N_3924);
or U4282 (N_4282,N_3918,N_3867);
or U4283 (N_4283,N_3909,N_3968);
xnor U4284 (N_4284,N_3630,N_3561);
and U4285 (N_4285,N_3755,N_3883);
and U4286 (N_4286,N_3549,N_3581);
and U4287 (N_4287,N_3826,N_3996);
and U4288 (N_4288,N_3560,N_3625);
or U4289 (N_4289,N_3652,N_3866);
nor U4290 (N_4290,N_3820,N_3531);
nand U4291 (N_4291,N_3684,N_3598);
nand U4292 (N_4292,N_3830,N_3503);
nand U4293 (N_4293,N_3545,N_3624);
nand U4294 (N_4294,N_3695,N_3962);
nor U4295 (N_4295,N_3720,N_3535);
nand U4296 (N_4296,N_3620,N_3903);
and U4297 (N_4297,N_3609,N_3933);
and U4298 (N_4298,N_3719,N_3704);
and U4299 (N_4299,N_3855,N_3865);
nand U4300 (N_4300,N_3683,N_3559);
or U4301 (N_4301,N_3554,N_3604);
nor U4302 (N_4302,N_3523,N_3789);
xor U4303 (N_4303,N_3591,N_3892);
nand U4304 (N_4304,N_3691,N_3878);
or U4305 (N_4305,N_3916,N_3608);
nand U4306 (N_4306,N_3521,N_3834);
or U4307 (N_4307,N_3604,N_3569);
nor U4308 (N_4308,N_3527,N_3556);
xnor U4309 (N_4309,N_3850,N_3612);
nor U4310 (N_4310,N_3752,N_3808);
and U4311 (N_4311,N_3516,N_3765);
xnor U4312 (N_4312,N_3647,N_3934);
nand U4313 (N_4313,N_3862,N_3870);
nand U4314 (N_4314,N_3551,N_3766);
nor U4315 (N_4315,N_3853,N_3592);
and U4316 (N_4316,N_3605,N_3926);
xor U4317 (N_4317,N_3728,N_3607);
nor U4318 (N_4318,N_3649,N_3775);
or U4319 (N_4319,N_3779,N_3918);
nand U4320 (N_4320,N_3827,N_3554);
nand U4321 (N_4321,N_3568,N_3619);
or U4322 (N_4322,N_3584,N_3921);
or U4323 (N_4323,N_3638,N_3723);
nand U4324 (N_4324,N_3655,N_3786);
and U4325 (N_4325,N_3837,N_3701);
and U4326 (N_4326,N_3522,N_3909);
or U4327 (N_4327,N_3819,N_3717);
xor U4328 (N_4328,N_3551,N_3601);
and U4329 (N_4329,N_3923,N_3716);
and U4330 (N_4330,N_3512,N_3819);
nand U4331 (N_4331,N_3545,N_3581);
and U4332 (N_4332,N_3848,N_3768);
and U4333 (N_4333,N_3567,N_3663);
and U4334 (N_4334,N_3578,N_3635);
or U4335 (N_4335,N_3984,N_3808);
nand U4336 (N_4336,N_3677,N_3544);
and U4337 (N_4337,N_3957,N_3796);
nor U4338 (N_4338,N_3922,N_3961);
or U4339 (N_4339,N_3674,N_3713);
or U4340 (N_4340,N_3601,N_3715);
nand U4341 (N_4341,N_3639,N_3652);
or U4342 (N_4342,N_3891,N_3637);
nor U4343 (N_4343,N_3828,N_3844);
nand U4344 (N_4344,N_3699,N_3582);
nor U4345 (N_4345,N_3795,N_3890);
nand U4346 (N_4346,N_3522,N_3906);
nor U4347 (N_4347,N_3550,N_3892);
xor U4348 (N_4348,N_3890,N_3555);
and U4349 (N_4349,N_3913,N_3945);
and U4350 (N_4350,N_3768,N_3556);
and U4351 (N_4351,N_3579,N_3714);
or U4352 (N_4352,N_3845,N_3996);
nor U4353 (N_4353,N_3741,N_3506);
nand U4354 (N_4354,N_3910,N_3574);
nor U4355 (N_4355,N_3992,N_3571);
nor U4356 (N_4356,N_3817,N_3847);
nand U4357 (N_4357,N_3681,N_3975);
and U4358 (N_4358,N_3761,N_3887);
nand U4359 (N_4359,N_3962,N_3806);
or U4360 (N_4360,N_3666,N_3985);
nor U4361 (N_4361,N_3812,N_3864);
or U4362 (N_4362,N_3848,N_3567);
and U4363 (N_4363,N_3610,N_3758);
nand U4364 (N_4364,N_3582,N_3789);
and U4365 (N_4365,N_3625,N_3613);
and U4366 (N_4366,N_3678,N_3633);
and U4367 (N_4367,N_3766,N_3555);
xnor U4368 (N_4368,N_3691,N_3887);
or U4369 (N_4369,N_3541,N_3760);
and U4370 (N_4370,N_3845,N_3774);
and U4371 (N_4371,N_3672,N_3717);
or U4372 (N_4372,N_3534,N_3844);
nand U4373 (N_4373,N_3523,N_3961);
and U4374 (N_4374,N_3852,N_3859);
or U4375 (N_4375,N_3813,N_3549);
or U4376 (N_4376,N_3933,N_3652);
and U4377 (N_4377,N_3920,N_3656);
nor U4378 (N_4378,N_3784,N_3721);
or U4379 (N_4379,N_3851,N_3531);
nand U4380 (N_4380,N_3752,N_3666);
and U4381 (N_4381,N_3931,N_3810);
nor U4382 (N_4382,N_3733,N_3569);
nand U4383 (N_4383,N_3764,N_3673);
or U4384 (N_4384,N_3749,N_3888);
or U4385 (N_4385,N_3659,N_3958);
nand U4386 (N_4386,N_3809,N_3869);
or U4387 (N_4387,N_3743,N_3545);
and U4388 (N_4388,N_3772,N_3885);
nor U4389 (N_4389,N_3842,N_3692);
nor U4390 (N_4390,N_3738,N_3843);
or U4391 (N_4391,N_3699,N_3782);
nor U4392 (N_4392,N_3763,N_3764);
nand U4393 (N_4393,N_3590,N_3747);
and U4394 (N_4394,N_3912,N_3657);
or U4395 (N_4395,N_3690,N_3985);
nand U4396 (N_4396,N_3572,N_3829);
nand U4397 (N_4397,N_3831,N_3808);
nand U4398 (N_4398,N_3707,N_3560);
nor U4399 (N_4399,N_3953,N_3950);
nor U4400 (N_4400,N_3796,N_3874);
nor U4401 (N_4401,N_3786,N_3512);
and U4402 (N_4402,N_3888,N_3524);
and U4403 (N_4403,N_3862,N_3597);
nand U4404 (N_4404,N_3960,N_3608);
xor U4405 (N_4405,N_3848,N_3620);
nand U4406 (N_4406,N_3851,N_3955);
or U4407 (N_4407,N_3568,N_3523);
xnor U4408 (N_4408,N_3524,N_3700);
and U4409 (N_4409,N_3985,N_3531);
or U4410 (N_4410,N_3680,N_3869);
xor U4411 (N_4411,N_3862,N_3659);
or U4412 (N_4412,N_3640,N_3693);
nor U4413 (N_4413,N_3822,N_3961);
or U4414 (N_4414,N_3904,N_3543);
xor U4415 (N_4415,N_3863,N_3599);
or U4416 (N_4416,N_3922,N_3674);
nand U4417 (N_4417,N_3524,N_3900);
or U4418 (N_4418,N_3714,N_3947);
nor U4419 (N_4419,N_3767,N_3772);
xor U4420 (N_4420,N_3927,N_3828);
and U4421 (N_4421,N_3962,N_3968);
nor U4422 (N_4422,N_3764,N_3501);
or U4423 (N_4423,N_3645,N_3963);
or U4424 (N_4424,N_3846,N_3513);
nand U4425 (N_4425,N_3501,N_3664);
or U4426 (N_4426,N_3660,N_3578);
or U4427 (N_4427,N_3612,N_3968);
xor U4428 (N_4428,N_3620,N_3666);
and U4429 (N_4429,N_3989,N_3628);
nand U4430 (N_4430,N_3705,N_3961);
xor U4431 (N_4431,N_3720,N_3604);
nor U4432 (N_4432,N_3816,N_3822);
and U4433 (N_4433,N_3517,N_3873);
nor U4434 (N_4434,N_3735,N_3912);
or U4435 (N_4435,N_3665,N_3999);
and U4436 (N_4436,N_3918,N_3502);
and U4437 (N_4437,N_3820,N_3858);
nor U4438 (N_4438,N_3781,N_3981);
nand U4439 (N_4439,N_3624,N_3552);
nor U4440 (N_4440,N_3641,N_3946);
and U4441 (N_4441,N_3687,N_3700);
or U4442 (N_4442,N_3930,N_3520);
and U4443 (N_4443,N_3775,N_3934);
xor U4444 (N_4444,N_3865,N_3682);
nor U4445 (N_4445,N_3687,N_3803);
and U4446 (N_4446,N_3920,N_3594);
or U4447 (N_4447,N_3996,N_3664);
and U4448 (N_4448,N_3508,N_3690);
nor U4449 (N_4449,N_3842,N_3768);
nor U4450 (N_4450,N_3984,N_3617);
nor U4451 (N_4451,N_3812,N_3511);
xor U4452 (N_4452,N_3729,N_3794);
nor U4453 (N_4453,N_3879,N_3754);
or U4454 (N_4454,N_3932,N_3578);
and U4455 (N_4455,N_3961,N_3864);
nand U4456 (N_4456,N_3873,N_3576);
nor U4457 (N_4457,N_3801,N_3757);
or U4458 (N_4458,N_3700,N_3938);
nor U4459 (N_4459,N_3685,N_3951);
or U4460 (N_4460,N_3888,N_3732);
or U4461 (N_4461,N_3536,N_3671);
nand U4462 (N_4462,N_3662,N_3612);
and U4463 (N_4463,N_3537,N_3747);
nor U4464 (N_4464,N_3774,N_3758);
nand U4465 (N_4465,N_3716,N_3882);
nor U4466 (N_4466,N_3864,N_3856);
and U4467 (N_4467,N_3670,N_3737);
nand U4468 (N_4468,N_3797,N_3883);
nor U4469 (N_4469,N_3523,N_3730);
nand U4470 (N_4470,N_3996,N_3854);
xnor U4471 (N_4471,N_3657,N_3783);
nand U4472 (N_4472,N_3550,N_3890);
nand U4473 (N_4473,N_3660,N_3885);
and U4474 (N_4474,N_3734,N_3858);
nor U4475 (N_4475,N_3658,N_3757);
nand U4476 (N_4476,N_3620,N_3711);
nand U4477 (N_4477,N_3933,N_3596);
and U4478 (N_4478,N_3691,N_3512);
nor U4479 (N_4479,N_3948,N_3720);
nand U4480 (N_4480,N_3929,N_3734);
nand U4481 (N_4481,N_3851,N_3965);
nor U4482 (N_4482,N_3842,N_3755);
or U4483 (N_4483,N_3883,N_3537);
and U4484 (N_4484,N_3516,N_3939);
and U4485 (N_4485,N_3954,N_3983);
or U4486 (N_4486,N_3899,N_3555);
nand U4487 (N_4487,N_3984,N_3847);
xnor U4488 (N_4488,N_3975,N_3956);
nand U4489 (N_4489,N_3656,N_3977);
xnor U4490 (N_4490,N_3893,N_3935);
or U4491 (N_4491,N_3555,N_3699);
and U4492 (N_4492,N_3896,N_3773);
or U4493 (N_4493,N_3632,N_3586);
xnor U4494 (N_4494,N_3822,N_3921);
and U4495 (N_4495,N_3829,N_3895);
xor U4496 (N_4496,N_3627,N_3933);
nand U4497 (N_4497,N_3551,N_3786);
or U4498 (N_4498,N_3501,N_3680);
nor U4499 (N_4499,N_3692,N_3717);
or U4500 (N_4500,N_4354,N_4400);
xnor U4501 (N_4501,N_4372,N_4100);
or U4502 (N_4502,N_4072,N_4238);
and U4503 (N_4503,N_4351,N_4419);
nor U4504 (N_4504,N_4135,N_4492);
nor U4505 (N_4505,N_4139,N_4281);
and U4506 (N_4506,N_4491,N_4335);
and U4507 (N_4507,N_4343,N_4480);
or U4508 (N_4508,N_4498,N_4114);
nor U4509 (N_4509,N_4048,N_4120);
nand U4510 (N_4510,N_4373,N_4174);
nand U4511 (N_4511,N_4079,N_4111);
and U4512 (N_4512,N_4476,N_4325);
nor U4513 (N_4513,N_4395,N_4307);
or U4514 (N_4514,N_4332,N_4209);
nand U4515 (N_4515,N_4399,N_4387);
nand U4516 (N_4516,N_4087,N_4166);
xor U4517 (N_4517,N_4165,N_4308);
nand U4518 (N_4518,N_4499,N_4167);
and U4519 (N_4519,N_4271,N_4040);
nor U4520 (N_4520,N_4294,N_4277);
and U4521 (N_4521,N_4276,N_4097);
nand U4522 (N_4522,N_4088,N_4229);
nor U4523 (N_4523,N_4105,N_4326);
nor U4524 (N_4524,N_4226,N_4030);
xnor U4525 (N_4525,N_4024,N_4228);
and U4526 (N_4526,N_4394,N_4316);
nand U4527 (N_4527,N_4129,N_4002);
or U4528 (N_4528,N_4485,N_4392);
or U4529 (N_4529,N_4446,N_4213);
nand U4530 (N_4530,N_4283,N_4412);
nor U4531 (N_4531,N_4184,N_4258);
or U4532 (N_4532,N_4356,N_4149);
xnor U4533 (N_4533,N_4108,N_4192);
or U4534 (N_4534,N_4443,N_4011);
nor U4535 (N_4535,N_4101,N_4303);
nor U4536 (N_4536,N_4198,N_4451);
or U4537 (N_4537,N_4455,N_4243);
nor U4538 (N_4538,N_4159,N_4094);
nand U4539 (N_4539,N_4224,N_4241);
and U4540 (N_4540,N_4104,N_4145);
and U4541 (N_4541,N_4337,N_4244);
or U4542 (N_4542,N_4235,N_4185);
nand U4543 (N_4543,N_4413,N_4342);
nand U4544 (N_4544,N_4080,N_4403);
nor U4545 (N_4545,N_4046,N_4219);
or U4546 (N_4546,N_4274,N_4363);
nand U4547 (N_4547,N_4423,N_4099);
nor U4548 (N_4548,N_4312,N_4171);
and U4549 (N_4549,N_4338,N_4310);
nor U4550 (N_4550,N_4218,N_4160);
or U4551 (N_4551,N_4324,N_4035);
nand U4552 (N_4552,N_4267,N_4256);
nand U4553 (N_4553,N_4411,N_4306);
or U4554 (N_4554,N_4428,N_4345);
and U4555 (N_4555,N_4078,N_4297);
nand U4556 (N_4556,N_4031,N_4453);
or U4557 (N_4557,N_4199,N_4128);
nand U4558 (N_4558,N_4062,N_4421);
or U4559 (N_4559,N_4234,N_4300);
and U4560 (N_4560,N_4298,N_4318);
nand U4561 (N_4561,N_4003,N_4414);
nor U4562 (N_4562,N_4045,N_4489);
and U4563 (N_4563,N_4207,N_4056);
nor U4564 (N_4564,N_4064,N_4071);
and U4565 (N_4565,N_4393,N_4315);
or U4566 (N_4566,N_4349,N_4469);
nor U4567 (N_4567,N_4254,N_4361);
nand U4568 (N_4568,N_4242,N_4010);
nand U4569 (N_4569,N_4019,N_4376);
nor U4570 (N_4570,N_4470,N_4378);
nand U4571 (N_4571,N_4210,N_4435);
nor U4572 (N_4572,N_4295,N_4117);
nand U4573 (N_4573,N_4278,N_4331);
and U4574 (N_4574,N_4494,N_4482);
xor U4575 (N_4575,N_4313,N_4465);
or U4576 (N_4576,N_4050,N_4475);
and U4577 (N_4577,N_4444,N_4196);
and U4578 (N_4578,N_4102,N_4144);
and U4579 (N_4579,N_4442,N_4405);
nand U4580 (N_4580,N_4156,N_4216);
xnor U4581 (N_4581,N_4366,N_4365);
nand U4582 (N_4582,N_4259,N_4425);
or U4583 (N_4583,N_4106,N_4454);
nand U4584 (N_4584,N_4176,N_4113);
xor U4585 (N_4585,N_4076,N_4248);
nand U4586 (N_4586,N_4270,N_4095);
and U4587 (N_4587,N_4023,N_4146);
or U4588 (N_4588,N_4181,N_4367);
or U4589 (N_4589,N_4397,N_4127);
nor U4590 (N_4590,N_4118,N_4293);
nand U4591 (N_4591,N_4320,N_4066);
xor U4592 (N_4592,N_4410,N_4246);
or U4593 (N_4593,N_4255,N_4473);
xor U4594 (N_4594,N_4460,N_4092);
xnor U4595 (N_4595,N_4093,N_4404);
and U4596 (N_4596,N_4347,N_4236);
or U4597 (N_4597,N_4340,N_4057);
and U4598 (N_4598,N_4344,N_4091);
nor U4599 (N_4599,N_4452,N_4264);
or U4600 (N_4600,N_4205,N_4377);
xor U4601 (N_4601,N_4039,N_4291);
and U4602 (N_4602,N_4440,N_4427);
xnor U4603 (N_4603,N_4287,N_4309);
nand U4604 (N_4604,N_4483,N_4286);
or U4605 (N_4605,N_4133,N_4112);
or U4606 (N_4606,N_4371,N_4382);
nand U4607 (N_4607,N_4245,N_4402);
xor U4608 (N_4608,N_4038,N_4257);
nand U4609 (N_4609,N_4014,N_4004);
nand U4610 (N_4610,N_4022,N_4124);
or U4611 (N_4611,N_4082,N_4052);
xnor U4612 (N_4612,N_4265,N_4268);
nand U4613 (N_4613,N_4339,N_4116);
nor U4614 (N_4614,N_4169,N_4081);
and U4615 (N_4615,N_4383,N_4231);
and U4616 (N_4616,N_4186,N_4292);
nor U4617 (N_4617,N_4302,N_4075);
nor U4618 (N_4618,N_4047,N_4358);
and U4619 (N_4619,N_4379,N_4152);
and U4620 (N_4620,N_4136,N_4333);
nand U4621 (N_4621,N_4261,N_4032);
nand U4622 (N_4622,N_4468,N_4005);
nor U4623 (N_4623,N_4190,N_4179);
nor U4624 (N_4624,N_4466,N_4479);
nor U4625 (N_4625,N_4329,N_4138);
and U4626 (N_4626,N_4493,N_4009);
or U4627 (N_4627,N_4249,N_4086);
and U4628 (N_4628,N_4001,N_4305);
or U4629 (N_4629,N_4422,N_4222);
and U4630 (N_4630,N_4107,N_4158);
and U4631 (N_4631,N_4006,N_4330);
or U4632 (N_4632,N_4362,N_4073);
nand U4633 (N_4633,N_4183,N_4061);
or U4634 (N_4634,N_4177,N_4098);
nor U4635 (N_4635,N_4155,N_4284);
nand U4636 (N_4636,N_4497,N_4122);
and U4637 (N_4637,N_4280,N_4360);
nand U4638 (N_4638,N_4279,N_4457);
nor U4639 (N_4639,N_4153,N_4203);
nand U4640 (N_4640,N_4407,N_4083);
nand U4641 (N_4641,N_4389,N_4323);
and U4642 (N_4642,N_4364,N_4175);
nand U4643 (N_4643,N_4041,N_4008);
nand U4644 (N_4644,N_4195,N_4408);
nand U4645 (N_4645,N_4467,N_4143);
xor U4646 (N_4646,N_4201,N_4237);
or U4647 (N_4647,N_4348,N_4449);
and U4648 (N_4648,N_4161,N_4266);
nand U4649 (N_4649,N_4015,N_4434);
and U4650 (N_4650,N_4487,N_4194);
nor U4651 (N_4651,N_4123,N_4227);
nand U4652 (N_4652,N_4125,N_4285);
and U4653 (N_4653,N_4426,N_4142);
xnor U4654 (N_4654,N_4458,N_4021);
and U4655 (N_4655,N_4486,N_4130);
and U4656 (N_4656,N_4432,N_4020);
nand U4657 (N_4657,N_4275,N_4350);
nor U4658 (N_4658,N_4437,N_4439);
nor U4659 (N_4659,N_4007,N_4406);
and U4660 (N_4660,N_4162,N_4121);
and U4661 (N_4661,N_4202,N_4028);
nand U4662 (N_4662,N_4063,N_4193);
nor U4663 (N_4663,N_4396,N_4172);
nand U4664 (N_4664,N_4441,N_4250);
xor U4665 (N_4665,N_4059,N_4027);
or U4666 (N_4666,N_4018,N_4012);
nand U4667 (N_4667,N_4481,N_4311);
or U4668 (N_4668,N_4200,N_4384);
nor U4669 (N_4669,N_4390,N_4074);
and U4670 (N_4670,N_4137,N_4187);
nor U4671 (N_4671,N_4418,N_4416);
and U4672 (N_4672,N_4409,N_4141);
nor U4673 (N_4673,N_4206,N_4474);
nand U4674 (N_4674,N_4368,N_4462);
nor U4675 (N_4675,N_4401,N_4110);
or U4676 (N_4676,N_4191,N_4429);
nor U4677 (N_4677,N_4208,N_4215);
or U4678 (N_4678,N_4164,N_4036);
nand U4679 (N_4679,N_4464,N_4353);
nand U4680 (N_4680,N_4084,N_4272);
nand U4681 (N_4681,N_4025,N_4431);
nor U4682 (N_4682,N_4447,N_4496);
nand U4683 (N_4683,N_4060,N_4239);
nor U4684 (N_4684,N_4296,N_4051);
or U4685 (N_4685,N_4433,N_4370);
xnor U4686 (N_4686,N_4260,N_4214);
or U4687 (N_4687,N_4178,N_4314);
nand U4688 (N_4688,N_4067,N_4484);
nand U4689 (N_4689,N_4119,N_4230);
nand U4690 (N_4690,N_4150,N_4381);
and U4691 (N_4691,N_4478,N_4044);
xnor U4692 (N_4692,N_4319,N_4134);
nand U4693 (N_4693,N_4301,N_4355);
and U4694 (N_4694,N_4000,N_4420);
nor U4695 (N_4695,N_4336,N_4131);
nand U4696 (N_4696,N_4415,N_4450);
and U4697 (N_4697,N_4334,N_4077);
or U4698 (N_4698,N_4252,N_4217);
nor U4699 (N_4699,N_4033,N_4026);
nor U4700 (N_4700,N_4157,N_4398);
nand U4701 (N_4701,N_4225,N_4380);
xnor U4702 (N_4702,N_4170,N_4448);
nor U4703 (N_4703,N_4090,N_4154);
and U4704 (N_4704,N_4043,N_4352);
nand U4705 (N_4705,N_4438,N_4289);
and U4706 (N_4706,N_4357,N_4037);
nand U4707 (N_4707,N_4232,N_4321);
and U4708 (N_4708,N_4269,N_4240);
nor U4709 (N_4709,N_4029,N_4463);
and U4710 (N_4710,N_4263,N_4328);
and U4711 (N_4711,N_4459,N_4042);
nor U4712 (N_4712,N_4282,N_4299);
and U4713 (N_4713,N_4430,N_4290);
xor U4714 (N_4714,N_4251,N_4070);
or U4715 (N_4715,N_4374,N_4188);
xor U4716 (N_4716,N_4189,N_4197);
or U4717 (N_4717,N_4288,N_4273);
and U4718 (N_4718,N_4212,N_4103);
xnor U4719 (N_4719,N_4495,N_4147);
and U4720 (N_4720,N_4304,N_4211);
nand U4721 (N_4721,N_4055,N_4317);
nand U4722 (N_4722,N_4085,N_4359);
or U4723 (N_4723,N_4253,N_4115);
nand U4724 (N_4724,N_4058,N_4132);
nor U4725 (N_4725,N_4221,N_4375);
and U4726 (N_4726,N_4385,N_4151);
nor U4727 (N_4727,N_4126,N_4388);
and U4728 (N_4728,N_4233,N_4069);
nor U4729 (N_4729,N_4391,N_4204);
and U4730 (N_4730,N_4054,N_4017);
or U4731 (N_4731,N_4247,N_4327);
nor U4732 (N_4732,N_4341,N_4262);
and U4733 (N_4733,N_4053,N_4173);
nand U4734 (N_4734,N_4089,N_4477);
xnor U4735 (N_4735,N_4220,N_4346);
xor U4736 (N_4736,N_4471,N_4445);
and U4737 (N_4737,N_4182,N_4168);
nor U4738 (N_4738,N_4034,N_4424);
and U4739 (N_4739,N_4488,N_4140);
and U4740 (N_4740,N_4386,N_4436);
and U4741 (N_4741,N_4016,N_4417);
nand U4742 (N_4742,N_4109,N_4096);
nand U4743 (N_4743,N_4068,N_4049);
nand U4744 (N_4744,N_4461,N_4472);
nand U4745 (N_4745,N_4490,N_4322);
nand U4746 (N_4746,N_4223,N_4065);
nand U4747 (N_4747,N_4456,N_4148);
nand U4748 (N_4748,N_4013,N_4369);
nand U4749 (N_4749,N_4180,N_4163);
or U4750 (N_4750,N_4181,N_4051);
or U4751 (N_4751,N_4116,N_4444);
nand U4752 (N_4752,N_4107,N_4078);
nand U4753 (N_4753,N_4029,N_4234);
or U4754 (N_4754,N_4435,N_4193);
and U4755 (N_4755,N_4143,N_4234);
and U4756 (N_4756,N_4497,N_4363);
nor U4757 (N_4757,N_4246,N_4152);
or U4758 (N_4758,N_4236,N_4427);
nand U4759 (N_4759,N_4170,N_4035);
nor U4760 (N_4760,N_4309,N_4199);
xor U4761 (N_4761,N_4392,N_4491);
or U4762 (N_4762,N_4102,N_4255);
and U4763 (N_4763,N_4094,N_4414);
and U4764 (N_4764,N_4265,N_4196);
and U4765 (N_4765,N_4257,N_4105);
xor U4766 (N_4766,N_4325,N_4327);
nand U4767 (N_4767,N_4215,N_4119);
and U4768 (N_4768,N_4261,N_4018);
nand U4769 (N_4769,N_4252,N_4303);
and U4770 (N_4770,N_4471,N_4442);
or U4771 (N_4771,N_4325,N_4381);
and U4772 (N_4772,N_4116,N_4458);
xor U4773 (N_4773,N_4385,N_4000);
nor U4774 (N_4774,N_4458,N_4233);
nand U4775 (N_4775,N_4233,N_4471);
nand U4776 (N_4776,N_4218,N_4436);
or U4777 (N_4777,N_4353,N_4147);
nand U4778 (N_4778,N_4408,N_4355);
and U4779 (N_4779,N_4495,N_4356);
and U4780 (N_4780,N_4400,N_4016);
and U4781 (N_4781,N_4134,N_4180);
and U4782 (N_4782,N_4480,N_4309);
nor U4783 (N_4783,N_4393,N_4038);
and U4784 (N_4784,N_4166,N_4405);
and U4785 (N_4785,N_4459,N_4106);
xnor U4786 (N_4786,N_4019,N_4356);
or U4787 (N_4787,N_4149,N_4413);
or U4788 (N_4788,N_4098,N_4044);
or U4789 (N_4789,N_4244,N_4330);
nand U4790 (N_4790,N_4309,N_4035);
or U4791 (N_4791,N_4216,N_4162);
and U4792 (N_4792,N_4387,N_4324);
nand U4793 (N_4793,N_4027,N_4109);
or U4794 (N_4794,N_4100,N_4420);
and U4795 (N_4795,N_4456,N_4336);
nor U4796 (N_4796,N_4005,N_4031);
and U4797 (N_4797,N_4433,N_4238);
xnor U4798 (N_4798,N_4022,N_4444);
and U4799 (N_4799,N_4309,N_4448);
or U4800 (N_4800,N_4058,N_4476);
and U4801 (N_4801,N_4207,N_4040);
or U4802 (N_4802,N_4237,N_4040);
or U4803 (N_4803,N_4351,N_4136);
xor U4804 (N_4804,N_4123,N_4217);
nor U4805 (N_4805,N_4387,N_4219);
nand U4806 (N_4806,N_4270,N_4145);
and U4807 (N_4807,N_4017,N_4394);
nand U4808 (N_4808,N_4291,N_4423);
nand U4809 (N_4809,N_4364,N_4285);
or U4810 (N_4810,N_4015,N_4353);
and U4811 (N_4811,N_4281,N_4224);
or U4812 (N_4812,N_4406,N_4299);
and U4813 (N_4813,N_4238,N_4375);
nor U4814 (N_4814,N_4294,N_4409);
nor U4815 (N_4815,N_4395,N_4323);
or U4816 (N_4816,N_4184,N_4152);
or U4817 (N_4817,N_4235,N_4124);
or U4818 (N_4818,N_4127,N_4275);
or U4819 (N_4819,N_4097,N_4437);
or U4820 (N_4820,N_4267,N_4299);
nor U4821 (N_4821,N_4252,N_4313);
nand U4822 (N_4822,N_4335,N_4354);
nand U4823 (N_4823,N_4414,N_4208);
or U4824 (N_4824,N_4323,N_4033);
or U4825 (N_4825,N_4345,N_4097);
xor U4826 (N_4826,N_4421,N_4173);
and U4827 (N_4827,N_4245,N_4013);
or U4828 (N_4828,N_4450,N_4333);
xor U4829 (N_4829,N_4477,N_4436);
nor U4830 (N_4830,N_4438,N_4196);
nand U4831 (N_4831,N_4425,N_4462);
nand U4832 (N_4832,N_4131,N_4146);
or U4833 (N_4833,N_4443,N_4036);
nor U4834 (N_4834,N_4003,N_4153);
nor U4835 (N_4835,N_4498,N_4352);
or U4836 (N_4836,N_4313,N_4161);
nand U4837 (N_4837,N_4298,N_4264);
nor U4838 (N_4838,N_4001,N_4419);
xnor U4839 (N_4839,N_4057,N_4385);
or U4840 (N_4840,N_4378,N_4309);
and U4841 (N_4841,N_4304,N_4350);
nor U4842 (N_4842,N_4451,N_4128);
and U4843 (N_4843,N_4315,N_4282);
nor U4844 (N_4844,N_4224,N_4096);
and U4845 (N_4845,N_4247,N_4050);
or U4846 (N_4846,N_4285,N_4074);
or U4847 (N_4847,N_4214,N_4478);
nor U4848 (N_4848,N_4331,N_4136);
or U4849 (N_4849,N_4187,N_4420);
xor U4850 (N_4850,N_4317,N_4397);
nor U4851 (N_4851,N_4195,N_4376);
nand U4852 (N_4852,N_4189,N_4253);
and U4853 (N_4853,N_4268,N_4271);
nor U4854 (N_4854,N_4053,N_4169);
nand U4855 (N_4855,N_4053,N_4154);
nand U4856 (N_4856,N_4154,N_4198);
and U4857 (N_4857,N_4163,N_4397);
nand U4858 (N_4858,N_4224,N_4298);
nor U4859 (N_4859,N_4134,N_4416);
or U4860 (N_4860,N_4041,N_4162);
and U4861 (N_4861,N_4085,N_4302);
or U4862 (N_4862,N_4223,N_4327);
or U4863 (N_4863,N_4385,N_4302);
and U4864 (N_4864,N_4330,N_4010);
nand U4865 (N_4865,N_4037,N_4110);
or U4866 (N_4866,N_4315,N_4188);
xor U4867 (N_4867,N_4462,N_4343);
or U4868 (N_4868,N_4422,N_4352);
or U4869 (N_4869,N_4468,N_4106);
and U4870 (N_4870,N_4312,N_4068);
nand U4871 (N_4871,N_4120,N_4013);
or U4872 (N_4872,N_4412,N_4214);
nor U4873 (N_4873,N_4209,N_4090);
or U4874 (N_4874,N_4286,N_4405);
nand U4875 (N_4875,N_4054,N_4329);
nor U4876 (N_4876,N_4135,N_4344);
xor U4877 (N_4877,N_4377,N_4448);
or U4878 (N_4878,N_4109,N_4451);
and U4879 (N_4879,N_4292,N_4157);
nor U4880 (N_4880,N_4243,N_4278);
nor U4881 (N_4881,N_4184,N_4192);
xnor U4882 (N_4882,N_4111,N_4330);
and U4883 (N_4883,N_4404,N_4372);
nand U4884 (N_4884,N_4186,N_4266);
nand U4885 (N_4885,N_4111,N_4141);
nor U4886 (N_4886,N_4457,N_4239);
nor U4887 (N_4887,N_4236,N_4084);
and U4888 (N_4888,N_4150,N_4133);
nor U4889 (N_4889,N_4021,N_4285);
and U4890 (N_4890,N_4444,N_4140);
and U4891 (N_4891,N_4459,N_4235);
and U4892 (N_4892,N_4499,N_4178);
or U4893 (N_4893,N_4156,N_4236);
or U4894 (N_4894,N_4018,N_4398);
nand U4895 (N_4895,N_4286,N_4214);
or U4896 (N_4896,N_4327,N_4226);
nor U4897 (N_4897,N_4254,N_4251);
and U4898 (N_4898,N_4246,N_4112);
or U4899 (N_4899,N_4174,N_4154);
or U4900 (N_4900,N_4470,N_4355);
nand U4901 (N_4901,N_4308,N_4017);
or U4902 (N_4902,N_4096,N_4185);
and U4903 (N_4903,N_4001,N_4366);
or U4904 (N_4904,N_4004,N_4122);
xor U4905 (N_4905,N_4188,N_4438);
nand U4906 (N_4906,N_4454,N_4037);
and U4907 (N_4907,N_4138,N_4248);
nor U4908 (N_4908,N_4409,N_4441);
nand U4909 (N_4909,N_4051,N_4369);
nand U4910 (N_4910,N_4069,N_4374);
and U4911 (N_4911,N_4386,N_4128);
nor U4912 (N_4912,N_4113,N_4417);
and U4913 (N_4913,N_4238,N_4210);
nor U4914 (N_4914,N_4241,N_4194);
nor U4915 (N_4915,N_4466,N_4339);
and U4916 (N_4916,N_4121,N_4209);
nor U4917 (N_4917,N_4224,N_4419);
nand U4918 (N_4918,N_4213,N_4308);
nor U4919 (N_4919,N_4088,N_4306);
nand U4920 (N_4920,N_4095,N_4001);
and U4921 (N_4921,N_4294,N_4283);
xor U4922 (N_4922,N_4276,N_4378);
or U4923 (N_4923,N_4209,N_4351);
nand U4924 (N_4924,N_4452,N_4290);
and U4925 (N_4925,N_4385,N_4252);
nand U4926 (N_4926,N_4235,N_4191);
or U4927 (N_4927,N_4193,N_4336);
nand U4928 (N_4928,N_4080,N_4412);
or U4929 (N_4929,N_4450,N_4178);
and U4930 (N_4930,N_4446,N_4276);
and U4931 (N_4931,N_4410,N_4296);
nand U4932 (N_4932,N_4319,N_4052);
xnor U4933 (N_4933,N_4122,N_4169);
xnor U4934 (N_4934,N_4387,N_4016);
or U4935 (N_4935,N_4489,N_4309);
and U4936 (N_4936,N_4150,N_4418);
nand U4937 (N_4937,N_4314,N_4301);
nand U4938 (N_4938,N_4067,N_4274);
and U4939 (N_4939,N_4435,N_4314);
and U4940 (N_4940,N_4045,N_4343);
xnor U4941 (N_4941,N_4123,N_4448);
nor U4942 (N_4942,N_4025,N_4297);
nor U4943 (N_4943,N_4405,N_4025);
nor U4944 (N_4944,N_4101,N_4309);
nor U4945 (N_4945,N_4218,N_4405);
and U4946 (N_4946,N_4023,N_4311);
nand U4947 (N_4947,N_4307,N_4263);
xnor U4948 (N_4948,N_4477,N_4200);
xor U4949 (N_4949,N_4477,N_4281);
or U4950 (N_4950,N_4034,N_4151);
or U4951 (N_4951,N_4172,N_4079);
nor U4952 (N_4952,N_4195,N_4213);
or U4953 (N_4953,N_4045,N_4017);
and U4954 (N_4954,N_4034,N_4096);
and U4955 (N_4955,N_4185,N_4272);
or U4956 (N_4956,N_4420,N_4320);
nand U4957 (N_4957,N_4208,N_4223);
xnor U4958 (N_4958,N_4141,N_4213);
nand U4959 (N_4959,N_4498,N_4453);
or U4960 (N_4960,N_4332,N_4308);
and U4961 (N_4961,N_4273,N_4440);
nand U4962 (N_4962,N_4427,N_4100);
nor U4963 (N_4963,N_4161,N_4241);
nor U4964 (N_4964,N_4217,N_4346);
or U4965 (N_4965,N_4024,N_4180);
xnor U4966 (N_4966,N_4087,N_4352);
and U4967 (N_4967,N_4274,N_4327);
nor U4968 (N_4968,N_4300,N_4202);
and U4969 (N_4969,N_4388,N_4434);
and U4970 (N_4970,N_4092,N_4045);
and U4971 (N_4971,N_4366,N_4048);
and U4972 (N_4972,N_4350,N_4399);
nand U4973 (N_4973,N_4379,N_4444);
nor U4974 (N_4974,N_4165,N_4072);
nand U4975 (N_4975,N_4189,N_4105);
nor U4976 (N_4976,N_4429,N_4251);
and U4977 (N_4977,N_4438,N_4266);
or U4978 (N_4978,N_4345,N_4207);
nor U4979 (N_4979,N_4451,N_4189);
and U4980 (N_4980,N_4374,N_4335);
nor U4981 (N_4981,N_4164,N_4009);
or U4982 (N_4982,N_4021,N_4071);
xnor U4983 (N_4983,N_4367,N_4366);
or U4984 (N_4984,N_4198,N_4460);
and U4985 (N_4985,N_4180,N_4081);
nand U4986 (N_4986,N_4205,N_4397);
or U4987 (N_4987,N_4176,N_4431);
nor U4988 (N_4988,N_4428,N_4412);
or U4989 (N_4989,N_4063,N_4065);
nand U4990 (N_4990,N_4370,N_4468);
and U4991 (N_4991,N_4271,N_4204);
and U4992 (N_4992,N_4212,N_4255);
or U4993 (N_4993,N_4028,N_4082);
xor U4994 (N_4994,N_4374,N_4350);
xor U4995 (N_4995,N_4148,N_4469);
nand U4996 (N_4996,N_4036,N_4236);
nand U4997 (N_4997,N_4343,N_4414);
nor U4998 (N_4998,N_4356,N_4367);
and U4999 (N_4999,N_4227,N_4336);
xnor U5000 (N_5000,N_4994,N_4894);
nand U5001 (N_5001,N_4860,N_4587);
or U5002 (N_5002,N_4917,N_4825);
and U5003 (N_5003,N_4715,N_4929);
xnor U5004 (N_5004,N_4651,N_4501);
nor U5005 (N_5005,N_4827,N_4553);
or U5006 (N_5006,N_4741,N_4882);
nand U5007 (N_5007,N_4661,N_4500);
and U5008 (N_5008,N_4566,N_4508);
nor U5009 (N_5009,N_4601,N_4757);
nor U5010 (N_5010,N_4855,N_4898);
nand U5011 (N_5011,N_4779,N_4516);
and U5012 (N_5012,N_4828,N_4678);
or U5013 (N_5013,N_4576,N_4796);
or U5014 (N_5014,N_4534,N_4765);
nand U5015 (N_5015,N_4841,N_4972);
and U5016 (N_5016,N_4591,N_4902);
or U5017 (N_5017,N_4676,N_4778);
nor U5018 (N_5018,N_4912,N_4689);
and U5019 (N_5019,N_4936,N_4667);
and U5020 (N_5020,N_4908,N_4890);
xor U5021 (N_5021,N_4829,N_4671);
and U5022 (N_5022,N_4598,N_4750);
nand U5023 (N_5023,N_4982,N_4948);
and U5024 (N_5024,N_4627,N_4990);
and U5025 (N_5025,N_4571,N_4680);
or U5026 (N_5026,N_4710,N_4513);
nand U5027 (N_5027,N_4998,N_4851);
and U5028 (N_5028,N_4502,N_4714);
xor U5029 (N_5029,N_4790,N_4704);
and U5030 (N_5030,N_4589,N_4970);
and U5031 (N_5031,N_4533,N_4547);
xor U5032 (N_5032,N_4599,N_4536);
or U5033 (N_5033,N_4938,N_4723);
nor U5034 (N_5034,N_4803,N_4614);
xor U5035 (N_5035,N_4694,N_4885);
and U5036 (N_5036,N_4818,N_4717);
or U5037 (N_5037,N_4563,N_4849);
and U5038 (N_5038,N_4783,N_4942);
or U5039 (N_5039,N_4659,N_4840);
nand U5040 (N_5040,N_4760,N_4868);
or U5041 (N_5041,N_4976,N_4672);
nand U5042 (N_5042,N_4570,N_4688);
and U5043 (N_5043,N_4557,N_4657);
or U5044 (N_5044,N_4558,N_4629);
nor U5045 (N_5045,N_4978,N_4742);
nand U5046 (N_5046,N_4679,N_4916);
nand U5047 (N_5047,N_4620,N_4837);
and U5048 (N_5048,N_4621,N_4945);
nor U5049 (N_5049,N_4539,N_4865);
xor U5050 (N_5050,N_4612,N_4517);
and U5051 (N_5051,N_4969,N_4608);
xor U5052 (N_5052,N_4867,N_4977);
and U5053 (N_5053,N_4718,N_4652);
xnor U5054 (N_5054,N_4858,N_4791);
or U5055 (N_5055,N_4550,N_4705);
and U5056 (N_5056,N_4737,N_4719);
or U5057 (N_5057,N_4919,N_4583);
and U5058 (N_5058,N_4896,N_4766);
xor U5059 (N_5059,N_4656,N_4979);
xnor U5060 (N_5060,N_4879,N_4707);
nor U5061 (N_5061,N_4792,N_4654);
or U5062 (N_5062,N_4987,N_4843);
and U5063 (N_5063,N_4826,N_4506);
and U5064 (N_5064,N_4693,N_4626);
xor U5065 (N_5065,N_4915,N_4909);
xnor U5066 (N_5066,N_4992,N_4997);
nor U5067 (N_5067,N_4615,N_4922);
and U5068 (N_5068,N_4594,N_4649);
or U5069 (N_5069,N_4716,N_4971);
and U5070 (N_5070,N_4875,N_4686);
and U5071 (N_5071,N_4895,N_4965);
and U5072 (N_5072,N_4511,N_4899);
xnor U5073 (N_5073,N_4930,N_4691);
and U5074 (N_5074,N_4735,N_4995);
nand U5075 (N_5075,N_4763,N_4876);
and U5076 (N_5076,N_4666,N_4546);
or U5077 (N_5077,N_4893,N_4815);
or U5078 (N_5078,N_4639,N_4759);
and U5079 (N_5079,N_4973,N_4607);
nor U5080 (N_5080,N_4838,N_4781);
and U5081 (N_5081,N_4728,N_4947);
nand U5082 (N_5082,N_4555,N_4519);
nand U5083 (N_5083,N_4952,N_4644);
nor U5084 (N_5084,N_4712,N_4526);
or U5085 (N_5085,N_4883,N_4623);
xnor U5086 (N_5086,N_4923,N_4761);
and U5087 (N_5087,N_4523,N_4640);
and U5088 (N_5088,N_4758,N_4762);
and U5089 (N_5089,N_4584,N_4634);
or U5090 (N_5090,N_4698,N_4812);
or U5091 (N_5091,N_4795,N_4920);
and U5092 (N_5092,N_4549,N_4525);
nand U5093 (N_5093,N_4518,N_4632);
nand U5094 (N_5094,N_4844,N_4537);
and U5095 (N_5095,N_4560,N_4753);
and U5096 (N_5096,N_4515,N_4754);
nor U5097 (N_5097,N_4673,N_4820);
nor U5098 (N_5098,N_4806,N_4535);
and U5099 (N_5099,N_4572,N_4805);
nand U5100 (N_5100,N_4903,N_4959);
or U5101 (N_5101,N_4586,N_4701);
nor U5102 (N_5102,N_4565,N_4552);
nor U5103 (N_5103,N_4824,N_4708);
and U5104 (N_5104,N_4776,N_4747);
nor U5105 (N_5105,N_4579,N_4692);
and U5106 (N_5106,N_4787,N_4514);
or U5107 (N_5107,N_4870,N_4703);
xor U5108 (N_5108,N_4683,N_4745);
xnor U5109 (N_5109,N_4813,N_4677);
nand U5110 (N_5110,N_4736,N_4551);
or U5111 (N_5111,N_4772,N_4530);
nand U5112 (N_5112,N_4748,N_4648);
nor U5113 (N_5113,N_4642,N_4799);
nand U5114 (N_5114,N_4630,N_4600);
nand U5115 (N_5115,N_4582,N_4684);
xnor U5116 (N_5116,N_4574,N_4524);
nand U5117 (N_5117,N_4907,N_4988);
nand U5118 (N_5118,N_4906,N_4764);
nand U5119 (N_5119,N_4853,N_4854);
and U5120 (N_5120,N_4605,N_4768);
nor U5121 (N_5121,N_4665,N_4996);
xnor U5122 (N_5122,N_4633,N_4789);
xor U5123 (N_5123,N_4538,N_4588);
nor U5124 (N_5124,N_4821,N_4880);
nand U5125 (N_5125,N_4732,N_4749);
or U5126 (N_5126,N_4562,N_4556);
and U5127 (N_5127,N_4842,N_4985);
nor U5128 (N_5128,N_4911,N_4784);
nand U5129 (N_5129,N_4581,N_4709);
xor U5130 (N_5130,N_4541,N_4956);
and U5131 (N_5131,N_4848,N_4733);
or U5132 (N_5132,N_4863,N_4738);
nand U5133 (N_5133,N_4554,N_4967);
or U5134 (N_5134,N_4986,N_4613);
nor U5135 (N_5135,N_4662,N_4674);
or U5136 (N_5136,N_4963,N_4816);
nand U5137 (N_5137,N_4878,N_4962);
nand U5138 (N_5138,N_4725,N_4528);
or U5139 (N_5139,N_4960,N_4527);
or U5140 (N_5140,N_4850,N_4597);
xnor U5141 (N_5141,N_4808,N_4881);
and U5142 (N_5142,N_4846,N_4833);
and U5143 (N_5143,N_4618,N_4951);
and U5144 (N_5144,N_4729,N_4924);
nand U5145 (N_5145,N_4713,N_4873);
nor U5146 (N_5146,N_4585,N_4617);
nand U5147 (N_5147,N_4811,N_4658);
nand U5148 (N_5148,N_4505,N_4869);
xnor U5149 (N_5149,N_4943,N_4577);
nor U5150 (N_5150,N_4578,N_4775);
xnor U5151 (N_5151,N_4940,N_4522);
nand U5152 (N_5152,N_4609,N_4625);
or U5153 (N_5153,N_4934,N_4981);
or U5154 (N_5154,N_4700,N_4567);
nand U5155 (N_5155,N_4905,N_4636);
xnor U5156 (N_5156,N_4975,N_4722);
xnor U5157 (N_5157,N_4509,N_4835);
nor U5158 (N_5158,N_4830,N_4966);
nand U5159 (N_5159,N_4797,N_4711);
or U5160 (N_5160,N_4660,N_4702);
and U5161 (N_5161,N_4993,N_4794);
nor U5162 (N_5162,N_4770,N_4690);
and U5163 (N_5163,N_4682,N_4961);
nor U5164 (N_5164,N_4592,N_4933);
and U5165 (N_5165,N_4918,N_4755);
or U5166 (N_5166,N_4569,N_4543);
nor U5167 (N_5167,N_4647,N_4891);
and U5168 (N_5168,N_4681,N_4974);
nor U5169 (N_5169,N_4596,N_4983);
or U5170 (N_5170,N_4769,N_4610);
nor U5171 (N_5171,N_4897,N_4889);
or U5172 (N_5172,N_4544,N_4675);
and U5173 (N_5173,N_4696,N_4635);
nand U5174 (N_5174,N_4801,N_4695);
nand U5175 (N_5175,N_4958,N_4980);
or U5176 (N_5176,N_4752,N_4595);
nand U5177 (N_5177,N_4872,N_4548);
xnor U5178 (N_5178,N_4886,N_4809);
nor U5179 (N_5179,N_4575,N_4545);
nand U5180 (N_5180,N_4941,N_4611);
nand U5181 (N_5181,N_4503,N_4670);
nor U5182 (N_5182,N_4939,N_4564);
xnor U5183 (N_5183,N_4646,N_4520);
nor U5184 (N_5184,N_4823,N_4726);
nor U5185 (N_5185,N_4871,N_4561);
and U5186 (N_5186,N_4914,N_4669);
and U5187 (N_5187,N_4932,N_4877);
xor U5188 (N_5188,N_4989,N_4730);
nand U5189 (N_5189,N_4913,N_4663);
and U5190 (N_5190,N_4955,N_4834);
nor U5191 (N_5191,N_4831,N_4857);
nand U5192 (N_5192,N_4756,N_4935);
nand U5193 (N_5193,N_4999,N_4743);
xnor U5194 (N_5194,N_4861,N_4814);
nand U5195 (N_5195,N_4847,N_4532);
nor U5196 (N_5196,N_4706,N_4624);
nand U5197 (N_5197,N_4862,N_4650);
and U5198 (N_5198,N_4653,N_4859);
or U5199 (N_5199,N_4817,N_4628);
and U5200 (N_5200,N_4602,N_4968);
and U5201 (N_5201,N_4949,N_4721);
or U5202 (N_5202,N_4800,N_4944);
nand U5203 (N_5203,N_4946,N_4641);
and U5204 (N_5204,N_4786,N_4740);
or U5205 (N_5205,N_4836,N_4773);
nand U5206 (N_5206,N_4874,N_4782);
nor U5207 (N_5207,N_4622,N_4852);
and U5208 (N_5208,N_4685,N_4788);
nand U5209 (N_5209,N_4751,N_4839);
nor U5210 (N_5210,N_4645,N_4631);
nor U5211 (N_5211,N_4904,N_4832);
or U5212 (N_5212,N_4668,N_4785);
or U5213 (N_5213,N_4606,N_4931);
nor U5214 (N_5214,N_4793,N_4746);
nand U5215 (N_5215,N_4655,N_4643);
or U5216 (N_5216,N_4542,N_4928);
nand U5217 (N_5217,N_4984,N_4529);
xor U5218 (N_5218,N_4910,N_4638);
or U5219 (N_5219,N_4925,N_4991);
or U5220 (N_5220,N_4568,N_4744);
xnor U5221 (N_5221,N_4510,N_4619);
or U5222 (N_5222,N_4864,N_4767);
nor U5223 (N_5223,N_4888,N_4798);
nor U5224 (N_5224,N_4504,N_4856);
or U5225 (N_5225,N_4964,N_4720);
nand U5226 (N_5226,N_4954,N_4774);
nor U5227 (N_5227,N_4687,N_4512);
or U5228 (N_5228,N_4921,N_4616);
or U5229 (N_5229,N_4540,N_4804);
nor U5230 (N_5230,N_4822,N_4573);
and U5231 (N_5231,N_4845,N_4771);
nor U5232 (N_5232,N_4777,N_4699);
nor U5233 (N_5233,N_4810,N_4900);
nor U5234 (N_5234,N_4892,N_4950);
nand U5235 (N_5235,N_4604,N_4637);
and U5236 (N_5236,N_4780,N_4531);
or U5237 (N_5237,N_4724,N_4866);
nand U5238 (N_5238,N_4507,N_4937);
nor U5239 (N_5239,N_4926,N_4884);
nor U5240 (N_5240,N_4887,N_4727);
nand U5241 (N_5241,N_4593,N_4734);
xor U5242 (N_5242,N_4603,N_4664);
or U5243 (N_5243,N_4953,N_4731);
nor U5244 (N_5244,N_4802,N_4819);
nor U5245 (N_5245,N_4957,N_4559);
nor U5246 (N_5246,N_4807,N_4590);
and U5247 (N_5247,N_4580,N_4927);
or U5248 (N_5248,N_4739,N_4901);
nand U5249 (N_5249,N_4697,N_4521);
or U5250 (N_5250,N_4541,N_4768);
nor U5251 (N_5251,N_4981,N_4511);
xnor U5252 (N_5252,N_4802,N_4974);
or U5253 (N_5253,N_4783,N_4714);
and U5254 (N_5254,N_4875,N_4690);
nor U5255 (N_5255,N_4643,N_4761);
nor U5256 (N_5256,N_4947,N_4667);
nor U5257 (N_5257,N_4916,N_4959);
and U5258 (N_5258,N_4660,N_4515);
nor U5259 (N_5259,N_4696,N_4873);
or U5260 (N_5260,N_4772,N_4841);
or U5261 (N_5261,N_4585,N_4860);
nor U5262 (N_5262,N_4618,N_4886);
nand U5263 (N_5263,N_4983,N_4730);
or U5264 (N_5264,N_4666,N_4978);
xor U5265 (N_5265,N_4725,N_4924);
or U5266 (N_5266,N_4637,N_4853);
nor U5267 (N_5267,N_4737,N_4662);
or U5268 (N_5268,N_4625,N_4970);
and U5269 (N_5269,N_4972,N_4878);
nor U5270 (N_5270,N_4636,N_4847);
nor U5271 (N_5271,N_4602,N_4945);
and U5272 (N_5272,N_4807,N_4784);
nor U5273 (N_5273,N_4873,N_4995);
nor U5274 (N_5274,N_4982,N_4983);
nand U5275 (N_5275,N_4660,N_4807);
and U5276 (N_5276,N_4652,N_4623);
and U5277 (N_5277,N_4961,N_4723);
nand U5278 (N_5278,N_4931,N_4737);
nand U5279 (N_5279,N_4990,N_4618);
nand U5280 (N_5280,N_4739,N_4693);
and U5281 (N_5281,N_4740,N_4964);
and U5282 (N_5282,N_4650,N_4784);
and U5283 (N_5283,N_4906,N_4710);
nand U5284 (N_5284,N_4898,N_4924);
nor U5285 (N_5285,N_4686,N_4867);
and U5286 (N_5286,N_4826,N_4979);
xnor U5287 (N_5287,N_4603,N_4992);
nor U5288 (N_5288,N_4871,N_4544);
or U5289 (N_5289,N_4538,N_4583);
or U5290 (N_5290,N_4689,N_4671);
xor U5291 (N_5291,N_4588,N_4615);
nor U5292 (N_5292,N_4577,N_4905);
and U5293 (N_5293,N_4505,N_4852);
nand U5294 (N_5294,N_4808,N_4937);
nand U5295 (N_5295,N_4888,N_4603);
and U5296 (N_5296,N_4840,N_4794);
xnor U5297 (N_5297,N_4836,N_4749);
or U5298 (N_5298,N_4700,N_4525);
or U5299 (N_5299,N_4870,N_4893);
nand U5300 (N_5300,N_4753,N_4874);
nor U5301 (N_5301,N_4996,N_4949);
xor U5302 (N_5302,N_4961,N_4750);
and U5303 (N_5303,N_4810,N_4523);
nand U5304 (N_5304,N_4772,N_4659);
nand U5305 (N_5305,N_4876,N_4574);
and U5306 (N_5306,N_4635,N_4854);
nor U5307 (N_5307,N_4864,N_4969);
nor U5308 (N_5308,N_4708,N_4590);
or U5309 (N_5309,N_4535,N_4584);
and U5310 (N_5310,N_4957,N_4539);
nor U5311 (N_5311,N_4672,N_4977);
nor U5312 (N_5312,N_4618,N_4532);
and U5313 (N_5313,N_4730,N_4685);
and U5314 (N_5314,N_4993,N_4996);
or U5315 (N_5315,N_4982,N_4848);
and U5316 (N_5316,N_4955,N_4994);
and U5317 (N_5317,N_4959,N_4810);
and U5318 (N_5318,N_4502,N_4770);
nor U5319 (N_5319,N_4928,N_4607);
nor U5320 (N_5320,N_4892,N_4902);
and U5321 (N_5321,N_4580,N_4878);
and U5322 (N_5322,N_4782,N_4603);
nand U5323 (N_5323,N_4722,N_4955);
and U5324 (N_5324,N_4754,N_4867);
nand U5325 (N_5325,N_4931,N_4739);
and U5326 (N_5326,N_4588,N_4529);
nor U5327 (N_5327,N_4692,N_4553);
and U5328 (N_5328,N_4526,N_4970);
xor U5329 (N_5329,N_4798,N_4577);
and U5330 (N_5330,N_4981,N_4650);
xor U5331 (N_5331,N_4697,N_4925);
or U5332 (N_5332,N_4687,N_4550);
and U5333 (N_5333,N_4912,N_4613);
or U5334 (N_5334,N_4569,N_4711);
nor U5335 (N_5335,N_4950,N_4828);
nand U5336 (N_5336,N_4617,N_4859);
nand U5337 (N_5337,N_4756,N_4667);
or U5338 (N_5338,N_4766,N_4704);
and U5339 (N_5339,N_4501,N_4642);
nor U5340 (N_5340,N_4981,N_4550);
xor U5341 (N_5341,N_4856,N_4611);
nor U5342 (N_5342,N_4926,N_4640);
and U5343 (N_5343,N_4827,N_4549);
nand U5344 (N_5344,N_4687,N_4843);
nor U5345 (N_5345,N_4569,N_4740);
and U5346 (N_5346,N_4548,N_4703);
and U5347 (N_5347,N_4803,N_4751);
nor U5348 (N_5348,N_4847,N_4654);
or U5349 (N_5349,N_4878,N_4825);
or U5350 (N_5350,N_4684,N_4777);
nand U5351 (N_5351,N_4523,N_4776);
or U5352 (N_5352,N_4584,N_4917);
and U5353 (N_5353,N_4791,N_4859);
nor U5354 (N_5354,N_4519,N_4920);
or U5355 (N_5355,N_4963,N_4922);
nor U5356 (N_5356,N_4732,N_4929);
nor U5357 (N_5357,N_4761,N_4558);
and U5358 (N_5358,N_4891,N_4854);
or U5359 (N_5359,N_4798,N_4911);
or U5360 (N_5360,N_4794,N_4557);
nand U5361 (N_5361,N_4703,N_4624);
nand U5362 (N_5362,N_4960,N_4952);
xnor U5363 (N_5363,N_4631,N_4960);
or U5364 (N_5364,N_4966,N_4598);
xnor U5365 (N_5365,N_4768,N_4564);
and U5366 (N_5366,N_4668,N_4804);
nor U5367 (N_5367,N_4885,N_4775);
or U5368 (N_5368,N_4962,N_4615);
and U5369 (N_5369,N_4885,N_4558);
and U5370 (N_5370,N_4565,N_4528);
nor U5371 (N_5371,N_4637,N_4979);
or U5372 (N_5372,N_4853,N_4641);
and U5373 (N_5373,N_4556,N_4875);
nor U5374 (N_5374,N_4708,N_4947);
nand U5375 (N_5375,N_4899,N_4892);
or U5376 (N_5376,N_4897,N_4903);
nand U5377 (N_5377,N_4573,N_4582);
nor U5378 (N_5378,N_4646,N_4964);
nor U5379 (N_5379,N_4587,N_4531);
nor U5380 (N_5380,N_4932,N_4695);
nor U5381 (N_5381,N_4803,N_4514);
nor U5382 (N_5382,N_4623,N_4711);
nand U5383 (N_5383,N_4734,N_4857);
xor U5384 (N_5384,N_4548,N_4841);
nor U5385 (N_5385,N_4557,N_4790);
nor U5386 (N_5386,N_4914,N_4811);
or U5387 (N_5387,N_4762,N_4948);
and U5388 (N_5388,N_4518,N_4885);
xor U5389 (N_5389,N_4881,N_4871);
or U5390 (N_5390,N_4558,N_4679);
nand U5391 (N_5391,N_4661,N_4681);
nand U5392 (N_5392,N_4544,N_4823);
nor U5393 (N_5393,N_4641,N_4943);
nand U5394 (N_5394,N_4539,N_4849);
xor U5395 (N_5395,N_4783,N_4979);
nor U5396 (N_5396,N_4570,N_4605);
nor U5397 (N_5397,N_4902,N_4936);
nor U5398 (N_5398,N_4848,N_4930);
nor U5399 (N_5399,N_4553,N_4733);
nor U5400 (N_5400,N_4970,N_4963);
xor U5401 (N_5401,N_4598,N_4811);
xor U5402 (N_5402,N_4956,N_4763);
nand U5403 (N_5403,N_4903,N_4768);
nor U5404 (N_5404,N_4684,N_4845);
nor U5405 (N_5405,N_4861,N_4691);
nand U5406 (N_5406,N_4678,N_4689);
or U5407 (N_5407,N_4508,N_4970);
or U5408 (N_5408,N_4635,N_4862);
nand U5409 (N_5409,N_4604,N_4543);
nand U5410 (N_5410,N_4956,N_4612);
nand U5411 (N_5411,N_4889,N_4774);
nand U5412 (N_5412,N_4598,N_4715);
or U5413 (N_5413,N_4821,N_4871);
and U5414 (N_5414,N_4751,N_4994);
nor U5415 (N_5415,N_4966,N_4683);
and U5416 (N_5416,N_4928,N_4855);
nand U5417 (N_5417,N_4788,N_4503);
nand U5418 (N_5418,N_4854,N_4982);
or U5419 (N_5419,N_4874,N_4536);
and U5420 (N_5420,N_4731,N_4627);
or U5421 (N_5421,N_4738,N_4665);
or U5422 (N_5422,N_4570,N_4653);
nand U5423 (N_5423,N_4929,N_4966);
nand U5424 (N_5424,N_4698,N_4720);
or U5425 (N_5425,N_4948,N_4803);
or U5426 (N_5426,N_4657,N_4836);
and U5427 (N_5427,N_4915,N_4508);
or U5428 (N_5428,N_4908,N_4837);
or U5429 (N_5429,N_4706,N_4572);
nor U5430 (N_5430,N_4869,N_4510);
or U5431 (N_5431,N_4868,N_4901);
nor U5432 (N_5432,N_4822,N_4821);
nand U5433 (N_5433,N_4834,N_4642);
nand U5434 (N_5434,N_4673,N_4535);
nor U5435 (N_5435,N_4698,N_4794);
or U5436 (N_5436,N_4774,N_4815);
and U5437 (N_5437,N_4750,N_4755);
or U5438 (N_5438,N_4543,N_4678);
nand U5439 (N_5439,N_4949,N_4592);
and U5440 (N_5440,N_4818,N_4819);
xnor U5441 (N_5441,N_4585,N_4711);
nor U5442 (N_5442,N_4857,N_4850);
or U5443 (N_5443,N_4536,N_4650);
and U5444 (N_5444,N_4876,N_4672);
and U5445 (N_5445,N_4774,N_4670);
nand U5446 (N_5446,N_4516,N_4822);
nand U5447 (N_5447,N_4538,N_4571);
or U5448 (N_5448,N_4660,N_4597);
or U5449 (N_5449,N_4639,N_4714);
nand U5450 (N_5450,N_4995,N_4945);
and U5451 (N_5451,N_4744,N_4842);
nand U5452 (N_5452,N_4730,N_4801);
or U5453 (N_5453,N_4592,N_4904);
and U5454 (N_5454,N_4751,N_4528);
and U5455 (N_5455,N_4569,N_4881);
and U5456 (N_5456,N_4773,N_4810);
nor U5457 (N_5457,N_4500,N_4863);
nor U5458 (N_5458,N_4995,N_4731);
or U5459 (N_5459,N_4775,N_4842);
nor U5460 (N_5460,N_4502,N_4580);
and U5461 (N_5461,N_4620,N_4614);
nor U5462 (N_5462,N_4971,N_4681);
or U5463 (N_5463,N_4854,N_4809);
and U5464 (N_5464,N_4864,N_4530);
or U5465 (N_5465,N_4719,N_4616);
xor U5466 (N_5466,N_4861,N_4982);
and U5467 (N_5467,N_4764,N_4732);
nor U5468 (N_5468,N_4998,N_4812);
or U5469 (N_5469,N_4713,N_4885);
and U5470 (N_5470,N_4932,N_4682);
xnor U5471 (N_5471,N_4977,N_4780);
or U5472 (N_5472,N_4968,N_4634);
and U5473 (N_5473,N_4855,N_4530);
and U5474 (N_5474,N_4687,N_4674);
or U5475 (N_5475,N_4866,N_4930);
or U5476 (N_5476,N_4730,N_4824);
xnor U5477 (N_5477,N_4603,N_4930);
nor U5478 (N_5478,N_4892,N_4817);
nand U5479 (N_5479,N_4933,N_4686);
and U5480 (N_5480,N_4627,N_4685);
xnor U5481 (N_5481,N_4776,N_4808);
and U5482 (N_5482,N_4732,N_4814);
xnor U5483 (N_5483,N_4597,N_4528);
nand U5484 (N_5484,N_4979,N_4903);
nor U5485 (N_5485,N_4542,N_4665);
nand U5486 (N_5486,N_4508,N_4885);
and U5487 (N_5487,N_4753,N_4574);
and U5488 (N_5488,N_4886,N_4628);
nand U5489 (N_5489,N_4935,N_4995);
nand U5490 (N_5490,N_4601,N_4821);
or U5491 (N_5491,N_4807,N_4869);
and U5492 (N_5492,N_4962,N_4544);
and U5493 (N_5493,N_4669,N_4973);
xor U5494 (N_5494,N_4641,N_4746);
xnor U5495 (N_5495,N_4942,N_4562);
nand U5496 (N_5496,N_4521,N_4787);
nor U5497 (N_5497,N_4508,N_4959);
nand U5498 (N_5498,N_4677,N_4521);
xor U5499 (N_5499,N_4915,N_4977);
or U5500 (N_5500,N_5263,N_5446);
or U5501 (N_5501,N_5053,N_5361);
nand U5502 (N_5502,N_5416,N_5138);
nand U5503 (N_5503,N_5316,N_5388);
or U5504 (N_5504,N_5418,N_5354);
nand U5505 (N_5505,N_5050,N_5267);
or U5506 (N_5506,N_5006,N_5124);
or U5507 (N_5507,N_5114,N_5450);
nand U5508 (N_5508,N_5429,N_5087);
and U5509 (N_5509,N_5023,N_5355);
or U5510 (N_5510,N_5403,N_5194);
and U5511 (N_5511,N_5382,N_5379);
nand U5512 (N_5512,N_5497,N_5183);
or U5513 (N_5513,N_5166,N_5414);
or U5514 (N_5514,N_5494,N_5459);
nand U5515 (N_5515,N_5454,N_5412);
nor U5516 (N_5516,N_5490,N_5219);
and U5517 (N_5517,N_5499,N_5251);
and U5518 (N_5518,N_5203,N_5034);
xor U5519 (N_5519,N_5482,N_5280);
xor U5520 (N_5520,N_5109,N_5027);
nor U5521 (N_5521,N_5223,N_5299);
nor U5522 (N_5522,N_5464,N_5275);
and U5523 (N_5523,N_5004,N_5322);
nand U5524 (N_5524,N_5070,N_5365);
xor U5525 (N_5525,N_5484,N_5082);
nor U5526 (N_5526,N_5302,N_5474);
or U5527 (N_5527,N_5029,N_5139);
nand U5528 (N_5528,N_5468,N_5417);
nor U5529 (N_5529,N_5340,N_5231);
and U5530 (N_5530,N_5310,N_5432);
nor U5531 (N_5531,N_5458,N_5297);
and U5532 (N_5532,N_5154,N_5237);
and U5533 (N_5533,N_5160,N_5091);
or U5534 (N_5534,N_5366,N_5157);
nor U5535 (N_5535,N_5456,N_5448);
or U5536 (N_5536,N_5402,N_5329);
and U5537 (N_5537,N_5054,N_5017);
and U5538 (N_5538,N_5117,N_5009);
and U5539 (N_5539,N_5304,N_5397);
nand U5540 (N_5540,N_5031,N_5281);
or U5541 (N_5541,N_5073,N_5296);
xnor U5542 (N_5542,N_5074,N_5106);
nor U5543 (N_5543,N_5457,N_5318);
nand U5544 (N_5544,N_5003,N_5099);
and U5545 (N_5545,N_5171,N_5016);
nand U5546 (N_5546,N_5202,N_5442);
nand U5547 (N_5547,N_5420,N_5462);
or U5548 (N_5548,N_5078,N_5118);
nand U5549 (N_5549,N_5368,N_5426);
or U5550 (N_5550,N_5007,N_5151);
nand U5551 (N_5551,N_5390,N_5461);
xnor U5552 (N_5552,N_5039,N_5463);
or U5553 (N_5553,N_5327,N_5077);
or U5554 (N_5554,N_5019,N_5069);
or U5555 (N_5555,N_5348,N_5192);
nand U5556 (N_5556,N_5015,N_5083);
and U5557 (N_5557,N_5057,N_5294);
or U5558 (N_5558,N_5000,N_5059);
nand U5559 (N_5559,N_5066,N_5245);
and U5560 (N_5560,N_5048,N_5303);
and U5561 (N_5561,N_5313,N_5277);
and U5562 (N_5562,N_5234,N_5274);
xor U5563 (N_5563,N_5123,N_5162);
or U5564 (N_5564,N_5349,N_5481);
or U5565 (N_5565,N_5206,N_5384);
or U5566 (N_5566,N_5147,N_5400);
xnor U5567 (N_5567,N_5172,N_5197);
or U5568 (N_5568,N_5269,N_5063);
nor U5569 (N_5569,N_5467,N_5079);
nor U5570 (N_5570,N_5145,N_5150);
xnor U5571 (N_5571,N_5037,N_5451);
and U5572 (N_5572,N_5127,N_5434);
and U5573 (N_5573,N_5419,N_5359);
nand U5574 (N_5574,N_5170,N_5184);
or U5575 (N_5575,N_5014,N_5328);
and U5576 (N_5576,N_5265,N_5360);
or U5577 (N_5577,N_5026,N_5307);
and U5578 (N_5578,N_5258,N_5421);
nand U5579 (N_5579,N_5239,N_5092);
nand U5580 (N_5580,N_5438,N_5301);
nand U5581 (N_5581,N_5075,N_5097);
nand U5582 (N_5582,N_5187,N_5241);
nor U5583 (N_5583,N_5080,N_5407);
and U5584 (N_5584,N_5144,N_5324);
and U5585 (N_5585,N_5248,N_5319);
nand U5586 (N_5586,N_5475,N_5222);
nor U5587 (N_5587,N_5393,N_5049);
or U5588 (N_5588,N_5242,N_5404);
or U5589 (N_5589,N_5305,N_5378);
nand U5590 (N_5590,N_5093,N_5455);
xnor U5591 (N_5591,N_5047,N_5444);
or U5592 (N_5592,N_5344,N_5411);
nor U5593 (N_5593,N_5196,N_5369);
or U5594 (N_5594,N_5220,N_5210);
nand U5595 (N_5595,N_5282,N_5189);
nand U5596 (N_5596,N_5396,N_5221);
nand U5597 (N_5597,N_5096,N_5142);
nand U5598 (N_5598,N_5363,N_5244);
nor U5599 (N_5599,N_5065,N_5428);
xnor U5600 (N_5600,N_5051,N_5169);
nor U5601 (N_5601,N_5067,N_5094);
and U5602 (N_5602,N_5317,N_5071);
and U5603 (N_5603,N_5140,N_5387);
xor U5604 (N_5604,N_5246,N_5178);
nor U5605 (N_5605,N_5135,N_5216);
nor U5606 (N_5606,N_5290,N_5121);
and U5607 (N_5607,N_5158,N_5370);
nor U5608 (N_5608,N_5035,N_5249);
xnor U5609 (N_5609,N_5110,N_5413);
and U5610 (N_5610,N_5001,N_5300);
and U5611 (N_5611,N_5466,N_5181);
nand U5612 (N_5612,N_5072,N_5055);
or U5613 (N_5613,N_5089,N_5153);
nor U5614 (N_5614,N_5453,N_5264);
or U5615 (N_5615,N_5351,N_5141);
nor U5616 (N_5616,N_5104,N_5250);
or U5617 (N_5617,N_5152,N_5218);
and U5618 (N_5618,N_5295,N_5149);
nand U5619 (N_5619,N_5228,N_5256);
nand U5620 (N_5620,N_5217,N_5491);
and U5621 (N_5621,N_5209,N_5227);
nor U5622 (N_5622,N_5460,N_5289);
or U5623 (N_5623,N_5389,N_5308);
nor U5624 (N_5624,N_5101,N_5284);
or U5625 (N_5625,N_5131,N_5052);
or U5626 (N_5626,N_5156,N_5408);
nand U5627 (N_5627,N_5298,N_5122);
and U5628 (N_5628,N_5350,N_5473);
and U5629 (N_5629,N_5410,N_5425);
and U5630 (N_5630,N_5060,N_5112);
or U5631 (N_5631,N_5155,N_5163);
or U5632 (N_5632,N_5485,N_5291);
and U5633 (N_5633,N_5364,N_5424);
nor U5634 (N_5634,N_5010,N_5115);
and U5635 (N_5635,N_5032,N_5386);
nand U5636 (N_5636,N_5020,N_5041);
xnor U5637 (N_5637,N_5180,N_5175);
nand U5638 (N_5638,N_5266,N_5174);
nor U5639 (N_5639,N_5190,N_5038);
nand U5640 (N_5640,N_5230,N_5452);
or U5641 (N_5641,N_5102,N_5312);
nand U5642 (N_5642,N_5492,N_5286);
nor U5643 (N_5643,N_5111,N_5213);
nor U5644 (N_5644,N_5084,N_5343);
nor U5645 (N_5645,N_5188,N_5042);
nand U5646 (N_5646,N_5323,N_5415);
and U5647 (N_5647,N_5431,N_5341);
or U5648 (N_5648,N_5377,N_5443);
and U5649 (N_5649,N_5168,N_5357);
and U5650 (N_5650,N_5285,N_5044);
nand U5651 (N_5651,N_5129,N_5165);
nand U5652 (N_5652,N_5385,N_5191);
nor U5653 (N_5653,N_5198,N_5214);
nor U5654 (N_5654,N_5201,N_5086);
and U5655 (N_5655,N_5476,N_5440);
or U5656 (N_5656,N_5119,N_5254);
nand U5657 (N_5657,N_5148,N_5236);
or U5658 (N_5658,N_5113,N_5100);
nand U5659 (N_5659,N_5381,N_5480);
and U5660 (N_5660,N_5478,N_5205);
nor U5661 (N_5661,N_5233,N_5422);
nor U5662 (N_5662,N_5179,N_5283);
nand U5663 (N_5663,N_5471,N_5371);
and U5664 (N_5664,N_5392,N_5098);
nand U5665 (N_5665,N_5208,N_5333);
nand U5666 (N_5666,N_5200,N_5182);
nand U5667 (N_5667,N_5173,N_5224);
nor U5668 (N_5668,N_5345,N_5081);
or U5669 (N_5669,N_5430,N_5043);
or U5670 (N_5670,N_5394,N_5225);
nor U5671 (N_5671,N_5268,N_5235);
nand U5672 (N_5672,N_5331,N_5433);
and U5673 (N_5673,N_5068,N_5347);
nor U5674 (N_5674,N_5030,N_5133);
and U5675 (N_5675,N_5399,N_5212);
nand U5676 (N_5676,N_5391,N_5332);
or U5677 (N_5677,N_5445,N_5279);
or U5678 (N_5678,N_5215,N_5186);
nand U5679 (N_5679,N_5489,N_5398);
and U5680 (N_5680,N_5271,N_5493);
or U5681 (N_5681,N_5103,N_5314);
or U5682 (N_5682,N_5335,N_5406);
and U5683 (N_5683,N_5409,N_5204);
nor U5684 (N_5684,N_5229,N_5177);
and U5685 (N_5685,N_5012,N_5105);
and U5686 (N_5686,N_5159,N_5401);
or U5687 (N_5687,N_5436,N_5374);
or U5688 (N_5688,N_5257,N_5176);
or U5689 (N_5689,N_5085,N_5108);
or U5690 (N_5690,N_5270,N_5018);
and U5691 (N_5691,N_5321,N_5477);
or U5692 (N_5692,N_5346,N_5496);
nor U5693 (N_5693,N_5375,N_5226);
nor U5694 (N_5694,N_5498,N_5326);
or U5695 (N_5695,N_5356,N_5252);
nand U5696 (N_5696,N_5146,N_5362);
nor U5697 (N_5697,N_5002,N_5336);
or U5698 (N_5698,N_5243,N_5259);
nor U5699 (N_5699,N_5207,N_5056);
and U5700 (N_5700,N_5260,N_5353);
nor U5701 (N_5701,N_5107,N_5447);
and U5702 (N_5702,N_5372,N_5488);
nand U5703 (N_5703,N_5276,N_5383);
and U5704 (N_5704,N_5376,N_5021);
and U5705 (N_5705,N_5465,N_5185);
nand U5706 (N_5706,N_5320,N_5358);
or U5707 (N_5707,N_5046,N_5132);
xnor U5708 (N_5708,N_5334,N_5022);
nor U5709 (N_5709,N_5199,N_5143);
nand U5710 (N_5710,N_5287,N_5293);
or U5711 (N_5711,N_5441,N_5193);
nor U5712 (N_5712,N_5278,N_5045);
nor U5713 (N_5713,N_5273,N_5126);
nand U5714 (N_5714,N_5373,N_5423);
nand U5715 (N_5715,N_5380,N_5011);
and U5716 (N_5716,N_5120,N_5449);
or U5717 (N_5717,N_5338,N_5125);
or U5718 (N_5718,N_5090,N_5330);
and U5719 (N_5719,N_5076,N_5405);
nand U5720 (N_5720,N_5483,N_5136);
and U5721 (N_5721,N_5342,N_5028);
nand U5722 (N_5722,N_5337,N_5325);
and U5723 (N_5723,N_5253,N_5062);
nor U5724 (N_5724,N_5247,N_5311);
or U5725 (N_5725,N_5013,N_5352);
nand U5726 (N_5726,N_5240,N_5261);
nor U5727 (N_5727,N_5195,N_5495);
xnor U5728 (N_5728,N_5061,N_5427);
or U5729 (N_5729,N_5306,N_5487);
and U5730 (N_5730,N_5088,N_5435);
nand U5731 (N_5731,N_5134,N_5469);
and U5732 (N_5732,N_5161,N_5232);
nand U5733 (N_5733,N_5128,N_5292);
nand U5734 (N_5734,N_5005,N_5064);
nor U5735 (N_5735,N_5040,N_5211);
and U5736 (N_5736,N_5479,N_5167);
nor U5737 (N_5737,N_5437,N_5008);
or U5738 (N_5738,N_5130,N_5262);
nor U5739 (N_5739,N_5164,N_5367);
or U5740 (N_5740,N_5288,N_5309);
xnor U5741 (N_5741,N_5238,N_5339);
nand U5742 (N_5742,N_5470,N_5439);
nor U5743 (N_5743,N_5095,N_5116);
or U5744 (N_5744,N_5395,N_5472);
and U5745 (N_5745,N_5036,N_5255);
nor U5746 (N_5746,N_5058,N_5025);
or U5747 (N_5747,N_5033,N_5024);
and U5748 (N_5748,N_5315,N_5486);
nand U5749 (N_5749,N_5137,N_5272);
and U5750 (N_5750,N_5086,N_5427);
and U5751 (N_5751,N_5445,N_5325);
nand U5752 (N_5752,N_5318,N_5444);
and U5753 (N_5753,N_5321,N_5330);
xnor U5754 (N_5754,N_5254,N_5133);
and U5755 (N_5755,N_5419,N_5174);
nor U5756 (N_5756,N_5183,N_5129);
or U5757 (N_5757,N_5215,N_5462);
and U5758 (N_5758,N_5043,N_5274);
nand U5759 (N_5759,N_5381,N_5348);
xnor U5760 (N_5760,N_5320,N_5414);
nor U5761 (N_5761,N_5116,N_5264);
or U5762 (N_5762,N_5216,N_5206);
nor U5763 (N_5763,N_5201,N_5382);
and U5764 (N_5764,N_5153,N_5481);
nor U5765 (N_5765,N_5059,N_5330);
nand U5766 (N_5766,N_5307,N_5148);
xnor U5767 (N_5767,N_5214,N_5449);
or U5768 (N_5768,N_5279,N_5111);
or U5769 (N_5769,N_5378,N_5480);
and U5770 (N_5770,N_5065,N_5364);
nand U5771 (N_5771,N_5489,N_5122);
nand U5772 (N_5772,N_5147,N_5021);
nor U5773 (N_5773,N_5282,N_5485);
nand U5774 (N_5774,N_5441,N_5432);
nand U5775 (N_5775,N_5104,N_5297);
and U5776 (N_5776,N_5426,N_5315);
or U5777 (N_5777,N_5064,N_5151);
nor U5778 (N_5778,N_5120,N_5179);
xnor U5779 (N_5779,N_5205,N_5392);
nor U5780 (N_5780,N_5287,N_5049);
xor U5781 (N_5781,N_5261,N_5209);
nor U5782 (N_5782,N_5314,N_5162);
or U5783 (N_5783,N_5323,N_5213);
nand U5784 (N_5784,N_5439,N_5014);
nand U5785 (N_5785,N_5393,N_5230);
nor U5786 (N_5786,N_5476,N_5312);
nand U5787 (N_5787,N_5043,N_5300);
nor U5788 (N_5788,N_5235,N_5008);
nand U5789 (N_5789,N_5061,N_5399);
or U5790 (N_5790,N_5026,N_5022);
nand U5791 (N_5791,N_5444,N_5363);
or U5792 (N_5792,N_5064,N_5349);
or U5793 (N_5793,N_5081,N_5270);
or U5794 (N_5794,N_5147,N_5065);
and U5795 (N_5795,N_5298,N_5418);
nand U5796 (N_5796,N_5478,N_5120);
and U5797 (N_5797,N_5329,N_5117);
nor U5798 (N_5798,N_5028,N_5452);
xor U5799 (N_5799,N_5053,N_5259);
or U5800 (N_5800,N_5050,N_5214);
and U5801 (N_5801,N_5161,N_5220);
or U5802 (N_5802,N_5287,N_5290);
or U5803 (N_5803,N_5176,N_5456);
and U5804 (N_5804,N_5433,N_5175);
and U5805 (N_5805,N_5347,N_5301);
xor U5806 (N_5806,N_5123,N_5266);
nand U5807 (N_5807,N_5104,N_5112);
and U5808 (N_5808,N_5281,N_5375);
or U5809 (N_5809,N_5085,N_5022);
or U5810 (N_5810,N_5381,N_5263);
and U5811 (N_5811,N_5029,N_5193);
and U5812 (N_5812,N_5074,N_5458);
nand U5813 (N_5813,N_5057,N_5033);
and U5814 (N_5814,N_5314,N_5253);
nand U5815 (N_5815,N_5328,N_5291);
nand U5816 (N_5816,N_5154,N_5177);
and U5817 (N_5817,N_5455,N_5344);
nor U5818 (N_5818,N_5188,N_5454);
nor U5819 (N_5819,N_5427,N_5022);
nand U5820 (N_5820,N_5388,N_5448);
or U5821 (N_5821,N_5369,N_5213);
xor U5822 (N_5822,N_5142,N_5323);
nor U5823 (N_5823,N_5340,N_5341);
xnor U5824 (N_5824,N_5183,N_5493);
nand U5825 (N_5825,N_5023,N_5361);
and U5826 (N_5826,N_5232,N_5151);
nand U5827 (N_5827,N_5068,N_5356);
nor U5828 (N_5828,N_5313,N_5049);
nor U5829 (N_5829,N_5128,N_5210);
or U5830 (N_5830,N_5329,N_5110);
nand U5831 (N_5831,N_5147,N_5411);
nor U5832 (N_5832,N_5466,N_5348);
xnor U5833 (N_5833,N_5440,N_5083);
nor U5834 (N_5834,N_5130,N_5445);
nor U5835 (N_5835,N_5132,N_5106);
nand U5836 (N_5836,N_5367,N_5341);
and U5837 (N_5837,N_5318,N_5170);
nand U5838 (N_5838,N_5463,N_5161);
or U5839 (N_5839,N_5085,N_5120);
or U5840 (N_5840,N_5379,N_5213);
xor U5841 (N_5841,N_5217,N_5450);
nor U5842 (N_5842,N_5110,N_5084);
and U5843 (N_5843,N_5195,N_5423);
nor U5844 (N_5844,N_5389,N_5270);
nor U5845 (N_5845,N_5468,N_5327);
and U5846 (N_5846,N_5487,N_5429);
nand U5847 (N_5847,N_5326,N_5110);
nand U5848 (N_5848,N_5490,N_5080);
nor U5849 (N_5849,N_5016,N_5252);
nor U5850 (N_5850,N_5120,N_5482);
nand U5851 (N_5851,N_5333,N_5273);
or U5852 (N_5852,N_5019,N_5306);
nand U5853 (N_5853,N_5067,N_5071);
and U5854 (N_5854,N_5338,N_5444);
or U5855 (N_5855,N_5144,N_5490);
nand U5856 (N_5856,N_5112,N_5349);
nand U5857 (N_5857,N_5093,N_5249);
or U5858 (N_5858,N_5373,N_5194);
nand U5859 (N_5859,N_5051,N_5439);
or U5860 (N_5860,N_5250,N_5084);
xor U5861 (N_5861,N_5064,N_5443);
nand U5862 (N_5862,N_5033,N_5227);
xor U5863 (N_5863,N_5197,N_5084);
nand U5864 (N_5864,N_5480,N_5079);
nand U5865 (N_5865,N_5447,N_5339);
and U5866 (N_5866,N_5469,N_5498);
xnor U5867 (N_5867,N_5132,N_5235);
nor U5868 (N_5868,N_5454,N_5396);
nor U5869 (N_5869,N_5398,N_5012);
or U5870 (N_5870,N_5377,N_5493);
or U5871 (N_5871,N_5101,N_5477);
xor U5872 (N_5872,N_5452,N_5056);
nor U5873 (N_5873,N_5013,N_5375);
xor U5874 (N_5874,N_5375,N_5143);
nand U5875 (N_5875,N_5084,N_5451);
nand U5876 (N_5876,N_5027,N_5389);
and U5877 (N_5877,N_5266,N_5103);
or U5878 (N_5878,N_5173,N_5349);
nor U5879 (N_5879,N_5355,N_5361);
or U5880 (N_5880,N_5445,N_5435);
or U5881 (N_5881,N_5131,N_5001);
nand U5882 (N_5882,N_5306,N_5252);
nand U5883 (N_5883,N_5055,N_5378);
or U5884 (N_5884,N_5004,N_5359);
nor U5885 (N_5885,N_5150,N_5177);
xnor U5886 (N_5886,N_5182,N_5140);
nand U5887 (N_5887,N_5412,N_5427);
or U5888 (N_5888,N_5223,N_5365);
nand U5889 (N_5889,N_5262,N_5122);
or U5890 (N_5890,N_5086,N_5499);
nor U5891 (N_5891,N_5396,N_5051);
nand U5892 (N_5892,N_5200,N_5378);
nor U5893 (N_5893,N_5325,N_5472);
and U5894 (N_5894,N_5173,N_5395);
and U5895 (N_5895,N_5487,N_5229);
nand U5896 (N_5896,N_5219,N_5299);
xor U5897 (N_5897,N_5447,N_5222);
and U5898 (N_5898,N_5341,N_5208);
nor U5899 (N_5899,N_5335,N_5321);
xnor U5900 (N_5900,N_5239,N_5201);
nand U5901 (N_5901,N_5168,N_5225);
or U5902 (N_5902,N_5304,N_5461);
xor U5903 (N_5903,N_5366,N_5408);
xnor U5904 (N_5904,N_5049,N_5489);
or U5905 (N_5905,N_5443,N_5251);
nor U5906 (N_5906,N_5096,N_5313);
nor U5907 (N_5907,N_5028,N_5077);
and U5908 (N_5908,N_5376,N_5117);
or U5909 (N_5909,N_5242,N_5270);
xor U5910 (N_5910,N_5189,N_5083);
and U5911 (N_5911,N_5247,N_5422);
nand U5912 (N_5912,N_5176,N_5239);
or U5913 (N_5913,N_5272,N_5061);
nor U5914 (N_5914,N_5033,N_5239);
or U5915 (N_5915,N_5113,N_5220);
nor U5916 (N_5916,N_5134,N_5363);
nand U5917 (N_5917,N_5040,N_5034);
nor U5918 (N_5918,N_5318,N_5241);
nor U5919 (N_5919,N_5333,N_5117);
xor U5920 (N_5920,N_5230,N_5237);
and U5921 (N_5921,N_5031,N_5093);
and U5922 (N_5922,N_5086,N_5292);
and U5923 (N_5923,N_5232,N_5001);
or U5924 (N_5924,N_5026,N_5283);
nand U5925 (N_5925,N_5232,N_5201);
and U5926 (N_5926,N_5017,N_5094);
nand U5927 (N_5927,N_5334,N_5317);
and U5928 (N_5928,N_5414,N_5054);
nor U5929 (N_5929,N_5337,N_5063);
nand U5930 (N_5930,N_5400,N_5052);
or U5931 (N_5931,N_5421,N_5104);
nand U5932 (N_5932,N_5277,N_5468);
xor U5933 (N_5933,N_5154,N_5309);
nor U5934 (N_5934,N_5181,N_5095);
nand U5935 (N_5935,N_5426,N_5424);
and U5936 (N_5936,N_5052,N_5128);
nor U5937 (N_5937,N_5273,N_5495);
or U5938 (N_5938,N_5312,N_5064);
or U5939 (N_5939,N_5296,N_5297);
and U5940 (N_5940,N_5156,N_5022);
nand U5941 (N_5941,N_5008,N_5251);
or U5942 (N_5942,N_5065,N_5409);
and U5943 (N_5943,N_5155,N_5038);
xnor U5944 (N_5944,N_5178,N_5389);
nand U5945 (N_5945,N_5356,N_5096);
and U5946 (N_5946,N_5379,N_5431);
or U5947 (N_5947,N_5262,N_5066);
and U5948 (N_5948,N_5337,N_5058);
and U5949 (N_5949,N_5261,N_5092);
and U5950 (N_5950,N_5260,N_5307);
or U5951 (N_5951,N_5165,N_5022);
nor U5952 (N_5952,N_5409,N_5043);
nor U5953 (N_5953,N_5375,N_5046);
or U5954 (N_5954,N_5474,N_5097);
and U5955 (N_5955,N_5331,N_5489);
nor U5956 (N_5956,N_5369,N_5215);
nand U5957 (N_5957,N_5253,N_5005);
xnor U5958 (N_5958,N_5460,N_5414);
and U5959 (N_5959,N_5237,N_5266);
and U5960 (N_5960,N_5333,N_5020);
nor U5961 (N_5961,N_5091,N_5001);
or U5962 (N_5962,N_5406,N_5249);
nand U5963 (N_5963,N_5223,N_5005);
nand U5964 (N_5964,N_5477,N_5445);
or U5965 (N_5965,N_5376,N_5298);
nor U5966 (N_5966,N_5429,N_5302);
or U5967 (N_5967,N_5439,N_5324);
nand U5968 (N_5968,N_5328,N_5226);
or U5969 (N_5969,N_5249,N_5073);
nand U5970 (N_5970,N_5110,N_5043);
nor U5971 (N_5971,N_5104,N_5033);
nor U5972 (N_5972,N_5248,N_5424);
nor U5973 (N_5973,N_5193,N_5414);
nand U5974 (N_5974,N_5219,N_5172);
and U5975 (N_5975,N_5289,N_5352);
nor U5976 (N_5976,N_5193,N_5426);
nand U5977 (N_5977,N_5285,N_5233);
xor U5978 (N_5978,N_5221,N_5362);
or U5979 (N_5979,N_5144,N_5365);
nor U5980 (N_5980,N_5353,N_5460);
and U5981 (N_5981,N_5379,N_5217);
or U5982 (N_5982,N_5137,N_5455);
or U5983 (N_5983,N_5141,N_5199);
and U5984 (N_5984,N_5078,N_5163);
nor U5985 (N_5985,N_5049,N_5486);
nor U5986 (N_5986,N_5370,N_5200);
xnor U5987 (N_5987,N_5338,N_5289);
xor U5988 (N_5988,N_5435,N_5136);
nand U5989 (N_5989,N_5142,N_5453);
and U5990 (N_5990,N_5187,N_5454);
or U5991 (N_5991,N_5440,N_5220);
or U5992 (N_5992,N_5481,N_5270);
or U5993 (N_5993,N_5222,N_5372);
nand U5994 (N_5994,N_5133,N_5337);
xor U5995 (N_5995,N_5476,N_5091);
or U5996 (N_5996,N_5185,N_5315);
or U5997 (N_5997,N_5015,N_5053);
nand U5998 (N_5998,N_5372,N_5139);
nor U5999 (N_5999,N_5010,N_5325);
nor U6000 (N_6000,N_5779,N_5608);
and U6001 (N_6001,N_5899,N_5833);
nor U6002 (N_6002,N_5829,N_5832);
or U6003 (N_6003,N_5906,N_5970);
nor U6004 (N_6004,N_5712,N_5768);
nand U6005 (N_6005,N_5851,N_5793);
or U6006 (N_6006,N_5972,N_5905);
nor U6007 (N_6007,N_5859,N_5950);
nand U6008 (N_6008,N_5576,N_5914);
and U6009 (N_6009,N_5936,N_5740);
xor U6010 (N_6010,N_5589,N_5605);
nand U6011 (N_6011,N_5979,N_5864);
nor U6012 (N_6012,N_5573,N_5858);
and U6013 (N_6013,N_5765,N_5989);
and U6014 (N_6014,N_5562,N_5944);
nand U6015 (N_6015,N_5582,N_5898);
and U6016 (N_6016,N_5949,N_5901);
and U6017 (N_6017,N_5560,N_5511);
or U6018 (N_6018,N_5971,N_5506);
nor U6019 (N_6019,N_5913,N_5633);
nand U6020 (N_6020,N_5788,N_5964);
or U6021 (N_6021,N_5609,N_5615);
and U6022 (N_6022,N_5504,N_5996);
nor U6023 (N_6023,N_5919,N_5885);
nor U6024 (N_6024,N_5692,N_5939);
nand U6025 (N_6025,N_5715,N_5694);
or U6026 (N_6026,N_5755,N_5565);
xor U6027 (N_6027,N_5522,N_5850);
and U6028 (N_6028,N_5528,N_5719);
xor U6029 (N_6029,N_5714,N_5963);
and U6030 (N_6030,N_5763,N_5678);
nand U6031 (N_6031,N_5874,N_5670);
xnor U6032 (N_6032,N_5772,N_5521);
nand U6033 (N_6033,N_5805,N_5546);
nand U6034 (N_6034,N_5697,N_5978);
nor U6035 (N_6035,N_5975,N_5876);
nand U6036 (N_6036,N_5544,N_5778);
or U6037 (N_6037,N_5908,N_5904);
xor U6038 (N_6038,N_5951,N_5825);
and U6039 (N_6039,N_5983,N_5619);
nor U6040 (N_6040,N_5928,N_5533);
nand U6041 (N_6041,N_5541,N_5593);
nor U6042 (N_6042,N_5551,N_5747);
and U6043 (N_6043,N_5759,N_5785);
or U6044 (N_6044,N_5806,N_5746);
or U6045 (N_6045,N_5836,N_5616);
xnor U6046 (N_6046,N_5705,N_5563);
xnor U6047 (N_6047,N_5770,N_5696);
nor U6048 (N_6048,N_5642,N_5802);
nor U6049 (N_6049,N_5910,N_5568);
nand U6050 (N_6050,N_5947,N_5826);
or U6051 (N_6051,N_5809,N_5869);
and U6052 (N_6052,N_5967,N_5875);
xor U6053 (N_6053,N_5830,N_5984);
nor U6054 (N_6054,N_5915,N_5995);
xnor U6055 (N_6055,N_5517,N_5912);
and U6056 (N_6056,N_5753,N_5916);
or U6057 (N_6057,N_5634,N_5854);
or U6058 (N_6058,N_5959,N_5668);
or U6059 (N_6059,N_5860,N_5695);
or U6060 (N_6060,N_5501,N_5515);
and U6061 (N_6061,N_5636,N_5985);
nor U6062 (N_6062,N_5643,N_5617);
nand U6063 (N_6063,N_5855,N_5811);
or U6064 (N_6064,N_5709,N_5725);
or U6065 (N_6065,N_5844,N_5784);
and U6066 (N_6066,N_5552,N_5766);
nand U6067 (N_6067,N_5952,N_5958);
or U6068 (N_6068,N_5786,N_5956);
or U6069 (N_6069,N_5790,N_5691);
nor U6070 (N_6070,N_5835,N_5856);
or U6071 (N_6071,N_5679,N_5942);
and U6072 (N_6072,N_5953,N_5867);
nand U6073 (N_6073,N_5520,N_5626);
nand U6074 (N_6074,N_5940,N_5597);
nor U6075 (N_6075,N_5706,N_5661);
and U6076 (N_6076,N_5516,N_5902);
or U6077 (N_6077,N_5641,N_5798);
nor U6078 (N_6078,N_5801,N_5583);
or U6079 (N_6079,N_5976,N_5594);
and U6080 (N_6080,N_5644,N_5657);
and U6081 (N_6081,N_5673,N_5726);
nand U6082 (N_6082,N_5539,N_5815);
nor U6083 (N_6083,N_5883,N_5586);
nand U6084 (N_6084,N_5820,N_5807);
and U6085 (N_6085,N_5839,N_5873);
xnor U6086 (N_6086,N_5926,N_5827);
or U6087 (N_6087,N_5866,N_5781);
xnor U6088 (N_6088,N_5771,N_5665);
nor U6089 (N_6089,N_5669,N_5675);
or U6090 (N_6090,N_5502,N_5693);
or U6091 (N_6091,N_5553,N_5812);
nand U6092 (N_6092,N_5738,N_5871);
nand U6093 (N_6093,N_5804,N_5505);
or U6094 (N_6094,N_5587,N_5532);
or U6095 (N_6095,N_5818,N_5998);
and U6096 (N_6096,N_5930,N_5795);
nand U6097 (N_6097,N_5723,N_5702);
or U6098 (N_6098,N_5613,N_5549);
xor U6099 (N_6099,N_5846,N_5757);
nand U6100 (N_6100,N_5838,N_5577);
nand U6101 (N_6101,N_5567,N_5966);
and U6102 (N_6102,N_5981,N_5720);
or U6103 (N_6103,N_5922,N_5965);
and U6104 (N_6104,N_5584,N_5853);
and U6105 (N_6105,N_5588,N_5897);
nor U6106 (N_6106,N_5843,N_5819);
or U6107 (N_6107,N_5711,N_5537);
xor U6108 (N_6108,N_5748,N_5625);
or U6109 (N_6109,N_5623,N_5736);
or U6110 (N_6110,N_5848,N_5704);
nor U6111 (N_6111,N_5686,N_5894);
or U6112 (N_6112,N_5782,N_5646);
or U6113 (N_6113,N_5775,N_5672);
and U6114 (N_6114,N_5895,N_5917);
and U6115 (N_6115,N_5776,N_5580);
xnor U6116 (N_6116,N_5624,N_5557);
and U6117 (N_6117,N_5934,N_5896);
nor U6118 (N_6118,N_5822,N_5513);
or U6119 (N_6119,N_5638,N_5534);
nor U6120 (N_6120,N_5857,N_5741);
or U6121 (N_6121,N_5758,N_5687);
xor U6122 (N_6122,N_5685,N_5890);
nand U6123 (N_6123,N_5703,N_5993);
nand U6124 (N_6124,N_5681,N_5509);
nor U6125 (N_6125,N_5612,N_5680);
nor U6126 (N_6126,N_5828,N_5994);
xor U6127 (N_6127,N_5841,N_5783);
or U6128 (N_6128,N_5724,N_5566);
nor U6129 (N_6129,N_5721,N_5962);
or U6130 (N_6130,N_5749,N_5664);
nand U6131 (N_6131,N_5764,N_5526);
and U6132 (N_6132,N_5637,N_5888);
xor U6133 (N_6133,N_5500,N_5650);
or U6134 (N_6134,N_5713,N_5558);
nor U6135 (N_6135,N_5925,N_5561);
nor U6136 (N_6136,N_5538,N_5777);
nand U6137 (N_6137,N_5799,N_5663);
and U6138 (N_6138,N_5655,N_5700);
and U6139 (N_6139,N_5525,N_5870);
or U6140 (N_6140,N_5957,N_5861);
xor U6141 (N_6141,N_5507,N_5519);
and U6142 (N_6142,N_5731,N_5973);
nor U6143 (N_6143,N_5977,N_5774);
and U6144 (N_6144,N_5632,N_5531);
or U6145 (N_6145,N_5773,N_5813);
xnor U6146 (N_6146,N_5542,N_5969);
and U6147 (N_6147,N_5933,N_5974);
nand U6148 (N_6148,N_5540,N_5654);
nor U6149 (N_6149,N_5992,N_5941);
xnor U6150 (N_6150,N_5999,N_5817);
nor U6151 (N_6151,N_5635,N_5954);
nor U6152 (N_6152,N_5732,N_5760);
xor U6153 (N_6153,N_5893,N_5647);
and U6154 (N_6154,N_5824,N_5518);
nor U6155 (N_6155,N_5920,N_5660);
or U6156 (N_6156,N_5629,N_5545);
and U6157 (N_6157,N_5780,N_5823);
and U6158 (N_6158,N_5658,N_5892);
or U6159 (N_6159,N_5960,N_5701);
nand U6160 (N_6160,N_5931,N_5847);
or U6161 (N_6161,N_5752,N_5676);
nor U6162 (N_6162,N_5907,N_5667);
nand U6163 (N_6163,N_5868,N_5767);
nor U6164 (N_6164,N_5729,N_5649);
nor U6165 (N_6165,N_5743,N_5816);
nor U6166 (N_6166,N_5645,N_5945);
nor U6167 (N_6167,N_5756,N_5622);
or U6168 (N_6168,N_5599,N_5514);
and U6169 (N_6169,N_5674,N_5581);
or U6170 (N_6170,N_5900,N_5834);
and U6171 (N_6171,N_5716,N_5707);
nand U6172 (N_6172,N_5968,N_5570);
nand U6173 (N_6173,N_5924,N_5879);
or U6174 (N_6174,N_5877,N_5728);
nand U6175 (N_6175,N_5938,N_5718);
xnor U6176 (N_6176,N_5590,N_5742);
or U6177 (N_6177,N_5671,N_5842);
and U6178 (N_6178,N_5683,N_5591);
nor U6179 (N_6179,N_5508,N_5659);
and U6180 (N_6180,N_5948,N_5717);
nand U6181 (N_6181,N_5881,N_5761);
or U6182 (N_6182,N_5909,N_5997);
and U6183 (N_6183,N_5730,N_5648);
or U6184 (N_6184,N_5651,N_5739);
and U6185 (N_6185,N_5598,N_5787);
xnor U6186 (N_6186,N_5733,N_5796);
xor U6187 (N_6187,N_5662,N_5555);
and U6188 (N_6188,N_5880,N_5872);
or U6189 (N_6189,N_5929,N_5602);
nor U6190 (N_6190,N_5792,N_5810);
or U6191 (N_6191,N_5510,N_5762);
or U6192 (N_6192,N_5512,N_5621);
nand U6193 (N_6193,N_5574,N_5556);
nor U6194 (N_6194,N_5955,N_5831);
nand U6195 (N_6195,N_5630,N_5600);
nor U6196 (N_6196,N_5988,N_5640);
xnor U6197 (N_6197,N_5980,N_5803);
nor U6198 (N_6198,N_5606,N_5987);
xor U6199 (N_6199,N_5564,N_5882);
nand U6200 (N_6200,N_5789,N_5927);
nor U6201 (N_6201,N_5610,N_5575);
nor U6202 (N_6202,N_5821,N_5791);
nor U6203 (N_6203,N_5536,N_5524);
or U6204 (N_6204,N_5611,N_5865);
nor U6205 (N_6205,N_5535,N_5639);
and U6206 (N_6206,N_5891,N_5699);
nand U6207 (N_6207,N_5620,N_5684);
and U6208 (N_6208,N_5585,N_5708);
xnor U6209 (N_6209,N_5921,N_5889);
nand U6210 (N_6210,N_5601,N_5886);
or U6211 (N_6211,N_5814,N_5604);
or U6212 (N_6212,N_5656,N_5614);
and U6213 (N_6213,N_5618,N_5961);
nor U6214 (N_6214,N_5529,N_5547);
nor U6215 (N_6215,N_5523,N_5698);
and U6216 (N_6216,N_5991,N_5652);
or U6217 (N_6217,N_5794,N_5840);
or U6218 (N_6218,N_5690,N_5849);
and U6219 (N_6219,N_5569,N_5937);
xor U6220 (N_6220,N_5548,N_5990);
and U6221 (N_6221,N_5982,N_5631);
nor U6222 (N_6222,N_5878,N_5751);
nor U6223 (N_6223,N_5530,N_5754);
nand U6224 (N_6224,N_5578,N_5628);
nor U6225 (N_6225,N_5923,N_5710);
nor U6226 (N_6226,N_5845,N_5903);
xor U6227 (N_6227,N_5554,N_5527);
and U6228 (N_6228,N_5918,N_5572);
nor U6229 (N_6229,N_5550,N_5559);
and U6230 (N_6230,N_5800,N_5744);
nor U6231 (N_6231,N_5627,N_5607);
or U6232 (N_6232,N_5797,N_5735);
nor U6233 (N_6233,N_5769,N_5689);
and U6234 (N_6234,N_5666,N_5596);
xor U6235 (N_6235,N_5935,N_5595);
nand U6236 (N_6236,N_5884,N_5571);
nand U6237 (N_6237,N_5579,N_5750);
and U6238 (N_6238,N_5603,N_5862);
and U6239 (N_6239,N_5837,N_5543);
or U6240 (N_6240,N_5932,N_5688);
nor U6241 (N_6241,N_5727,N_5734);
and U6242 (N_6242,N_5946,N_5745);
nand U6243 (N_6243,N_5592,N_5677);
and U6244 (N_6244,N_5887,N_5682);
nor U6245 (N_6245,N_5722,N_5503);
or U6246 (N_6246,N_5653,N_5986);
nor U6247 (N_6247,N_5911,N_5943);
nor U6248 (N_6248,N_5852,N_5863);
nor U6249 (N_6249,N_5737,N_5808);
nand U6250 (N_6250,N_5734,N_5952);
and U6251 (N_6251,N_5639,N_5709);
nor U6252 (N_6252,N_5683,N_5662);
nor U6253 (N_6253,N_5608,N_5774);
nand U6254 (N_6254,N_5669,N_5890);
and U6255 (N_6255,N_5579,N_5552);
or U6256 (N_6256,N_5588,N_5688);
nand U6257 (N_6257,N_5724,N_5760);
xnor U6258 (N_6258,N_5662,N_5596);
and U6259 (N_6259,N_5915,N_5582);
or U6260 (N_6260,N_5895,N_5800);
xor U6261 (N_6261,N_5692,N_5978);
or U6262 (N_6262,N_5859,N_5577);
xnor U6263 (N_6263,N_5801,N_5507);
and U6264 (N_6264,N_5557,N_5820);
xnor U6265 (N_6265,N_5729,N_5659);
nor U6266 (N_6266,N_5944,N_5816);
nor U6267 (N_6267,N_5756,N_5668);
nor U6268 (N_6268,N_5601,N_5741);
nor U6269 (N_6269,N_5576,N_5615);
nand U6270 (N_6270,N_5628,N_5837);
and U6271 (N_6271,N_5579,N_5749);
or U6272 (N_6272,N_5617,N_5719);
and U6273 (N_6273,N_5773,N_5519);
or U6274 (N_6274,N_5861,N_5714);
and U6275 (N_6275,N_5981,N_5529);
nor U6276 (N_6276,N_5541,N_5560);
nor U6277 (N_6277,N_5670,N_5553);
nor U6278 (N_6278,N_5536,N_5825);
and U6279 (N_6279,N_5793,N_5768);
xnor U6280 (N_6280,N_5689,N_5565);
or U6281 (N_6281,N_5622,N_5772);
nor U6282 (N_6282,N_5737,N_5966);
or U6283 (N_6283,N_5835,N_5834);
nor U6284 (N_6284,N_5550,N_5990);
nand U6285 (N_6285,N_5807,N_5847);
nand U6286 (N_6286,N_5705,N_5846);
and U6287 (N_6287,N_5782,N_5710);
xnor U6288 (N_6288,N_5789,N_5571);
or U6289 (N_6289,N_5747,N_5787);
nor U6290 (N_6290,N_5900,N_5757);
nor U6291 (N_6291,N_5654,N_5938);
or U6292 (N_6292,N_5862,N_5734);
nand U6293 (N_6293,N_5707,N_5914);
nor U6294 (N_6294,N_5741,N_5884);
nor U6295 (N_6295,N_5595,N_5740);
nor U6296 (N_6296,N_5980,N_5759);
nand U6297 (N_6297,N_5884,N_5586);
nand U6298 (N_6298,N_5954,N_5537);
nand U6299 (N_6299,N_5971,N_5678);
and U6300 (N_6300,N_5596,N_5956);
nand U6301 (N_6301,N_5988,N_5531);
nand U6302 (N_6302,N_5746,N_5695);
nand U6303 (N_6303,N_5971,N_5951);
and U6304 (N_6304,N_5568,N_5687);
nor U6305 (N_6305,N_5834,N_5881);
xnor U6306 (N_6306,N_5638,N_5647);
and U6307 (N_6307,N_5746,N_5910);
nand U6308 (N_6308,N_5914,N_5588);
nor U6309 (N_6309,N_5800,N_5671);
or U6310 (N_6310,N_5927,N_5630);
nand U6311 (N_6311,N_5822,N_5628);
xor U6312 (N_6312,N_5528,N_5750);
nand U6313 (N_6313,N_5999,N_5878);
or U6314 (N_6314,N_5611,N_5841);
or U6315 (N_6315,N_5863,N_5873);
and U6316 (N_6316,N_5789,N_5836);
nand U6317 (N_6317,N_5660,N_5719);
and U6318 (N_6318,N_5538,N_5596);
and U6319 (N_6319,N_5677,N_5521);
nand U6320 (N_6320,N_5846,N_5927);
and U6321 (N_6321,N_5671,N_5876);
xor U6322 (N_6322,N_5736,N_5533);
nor U6323 (N_6323,N_5762,N_5857);
nor U6324 (N_6324,N_5780,N_5621);
nor U6325 (N_6325,N_5806,N_5639);
or U6326 (N_6326,N_5781,N_5909);
or U6327 (N_6327,N_5947,N_5746);
or U6328 (N_6328,N_5593,N_5968);
nor U6329 (N_6329,N_5735,N_5541);
nand U6330 (N_6330,N_5823,N_5591);
or U6331 (N_6331,N_5579,N_5936);
and U6332 (N_6332,N_5803,N_5743);
or U6333 (N_6333,N_5647,N_5864);
or U6334 (N_6334,N_5749,N_5769);
or U6335 (N_6335,N_5783,N_5784);
nor U6336 (N_6336,N_5562,N_5806);
and U6337 (N_6337,N_5598,N_5625);
nand U6338 (N_6338,N_5769,N_5638);
nand U6339 (N_6339,N_5619,N_5821);
nand U6340 (N_6340,N_5507,N_5729);
and U6341 (N_6341,N_5715,N_5599);
and U6342 (N_6342,N_5662,N_5687);
nor U6343 (N_6343,N_5776,N_5536);
xnor U6344 (N_6344,N_5695,N_5924);
nor U6345 (N_6345,N_5517,N_5651);
nand U6346 (N_6346,N_5666,N_5626);
and U6347 (N_6347,N_5907,N_5573);
xnor U6348 (N_6348,N_5988,N_5997);
and U6349 (N_6349,N_5728,N_5853);
nor U6350 (N_6350,N_5875,N_5756);
nand U6351 (N_6351,N_5611,N_5543);
nor U6352 (N_6352,N_5847,N_5942);
and U6353 (N_6353,N_5887,N_5532);
and U6354 (N_6354,N_5962,N_5544);
and U6355 (N_6355,N_5916,N_5885);
and U6356 (N_6356,N_5575,N_5536);
and U6357 (N_6357,N_5651,N_5553);
nand U6358 (N_6358,N_5547,N_5914);
nor U6359 (N_6359,N_5822,N_5696);
nand U6360 (N_6360,N_5621,N_5618);
and U6361 (N_6361,N_5807,N_5896);
or U6362 (N_6362,N_5999,N_5956);
xnor U6363 (N_6363,N_5924,N_5921);
nand U6364 (N_6364,N_5920,N_5850);
nor U6365 (N_6365,N_5957,N_5988);
or U6366 (N_6366,N_5656,N_5898);
and U6367 (N_6367,N_5616,N_5675);
or U6368 (N_6368,N_5536,N_5587);
nand U6369 (N_6369,N_5609,N_5887);
nand U6370 (N_6370,N_5967,N_5953);
nor U6371 (N_6371,N_5836,N_5627);
nand U6372 (N_6372,N_5681,N_5548);
and U6373 (N_6373,N_5633,N_5919);
and U6374 (N_6374,N_5831,N_5569);
and U6375 (N_6375,N_5754,N_5846);
nor U6376 (N_6376,N_5569,N_5984);
nor U6377 (N_6377,N_5743,N_5819);
or U6378 (N_6378,N_5688,N_5953);
nand U6379 (N_6379,N_5662,N_5536);
or U6380 (N_6380,N_5810,N_5796);
nor U6381 (N_6381,N_5784,N_5735);
and U6382 (N_6382,N_5784,N_5752);
or U6383 (N_6383,N_5818,N_5601);
or U6384 (N_6384,N_5974,N_5551);
nand U6385 (N_6385,N_5655,N_5888);
nor U6386 (N_6386,N_5972,N_5773);
nand U6387 (N_6387,N_5970,N_5709);
nand U6388 (N_6388,N_5881,N_5720);
and U6389 (N_6389,N_5565,N_5717);
nor U6390 (N_6390,N_5538,N_5610);
or U6391 (N_6391,N_5799,N_5952);
or U6392 (N_6392,N_5988,N_5675);
and U6393 (N_6393,N_5548,N_5999);
and U6394 (N_6394,N_5597,N_5508);
nor U6395 (N_6395,N_5757,N_5991);
nor U6396 (N_6396,N_5508,N_5655);
xnor U6397 (N_6397,N_5684,N_5691);
nor U6398 (N_6398,N_5964,N_5733);
nand U6399 (N_6399,N_5826,N_5544);
or U6400 (N_6400,N_5682,N_5589);
xnor U6401 (N_6401,N_5574,N_5710);
nor U6402 (N_6402,N_5814,N_5699);
xor U6403 (N_6403,N_5961,N_5572);
and U6404 (N_6404,N_5829,N_5837);
and U6405 (N_6405,N_5706,N_5722);
nand U6406 (N_6406,N_5879,N_5788);
xor U6407 (N_6407,N_5686,N_5673);
and U6408 (N_6408,N_5854,N_5715);
nor U6409 (N_6409,N_5903,N_5755);
xor U6410 (N_6410,N_5588,N_5894);
nor U6411 (N_6411,N_5645,N_5649);
nand U6412 (N_6412,N_5728,N_5901);
and U6413 (N_6413,N_5926,N_5547);
and U6414 (N_6414,N_5679,N_5521);
or U6415 (N_6415,N_5737,N_5735);
nand U6416 (N_6416,N_5538,N_5672);
nand U6417 (N_6417,N_5967,N_5987);
or U6418 (N_6418,N_5830,N_5533);
or U6419 (N_6419,N_5729,N_5870);
nor U6420 (N_6420,N_5887,N_5672);
and U6421 (N_6421,N_5665,N_5787);
nor U6422 (N_6422,N_5918,N_5718);
nor U6423 (N_6423,N_5502,N_5565);
xor U6424 (N_6424,N_5890,N_5772);
xnor U6425 (N_6425,N_5658,N_5623);
nor U6426 (N_6426,N_5566,N_5852);
nand U6427 (N_6427,N_5743,N_5678);
xnor U6428 (N_6428,N_5998,N_5634);
nor U6429 (N_6429,N_5825,N_5631);
nand U6430 (N_6430,N_5772,N_5967);
xnor U6431 (N_6431,N_5967,N_5548);
nand U6432 (N_6432,N_5597,N_5988);
nand U6433 (N_6433,N_5652,N_5777);
nor U6434 (N_6434,N_5637,N_5503);
or U6435 (N_6435,N_5666,N_5872);
or U6436 (N_6436,N_5720,N_5644);
and U6437 (N_6437,N_5572,N_5864);
nand U6438 (N_6438,N_5543,N_5711);
nand U6439 (N_6439,N_5696,N_5631);
nand U6440 (N_6440,N_5937,N_5626);
or U6441 (N_6441,N_5854,N_5547);
and U6442 (N_6442,N_5959,N_5974);
or U6443 (N_6443,N_5507,N_5970);
nand U6444 (N_6444,N_5619,N_5918);
nand U6445 (N_6445,N_5655,N_5763);
xor U6446 (N_6446,N_5918,N_5803);
or U6447 (N_6447,N_5929,N_5831);
or U6448 (N_6448,N_5537,N_5808);
or U6449 (N_6449,N_5589,N_5677);
nor U6450 (N_6450,N_5893,N_5623);
and U6451 (N_6451,N_5590,N_5596);
nand U6452 (N_6452,N_5759,N_5818);
nor U6453 (N_6453,N_5823,N_5520);
xnor U6454 (N_6454,N_5988,N_5890);
nand U6455 (N_6455,N_5523,N_5735);
or U6456 (N_6456,N_5924,N_5923);
nor U6457 (N_6457,N_5781,N_5724);
nand U6458 (N_6458,N_5943,N_5809);
and U6459 (N_6459,N_5993,N_5798);
xor U6460 (N_6460,N_5539,N_5742);
nand U6461 (N_6461,N_5858,N_5969);
and U6462 (N_6462,N_5587,N_5812);
nor U6463 (N_6463,N_5564,N_5893);
or U6464 (N_6464,N_5795,N_5792);
or U6465 (N_6465,N_5997,N_5816);
or U6466 (N_6466,N_5763,N_5879);
nand U6467 (N_6467,N_5617,N_5757);
nand U6468 (N_6468,N_5684,N_5674);
or U6469 (N_6469,N_5852,N_5580);
and U6470 (N_6470,N_5743,N_5890);
nand U6471 (N_6471,N_5559,N_5834);
and U6472 (N_6472,N_5910,N_5743);
and U6473 (N_6473,N_5854,N_5982);
nor U6474 (N_6474,N_5671,N_5627);
nand U6475 (N_6475,N_5748,N_5825);
nor U6476 (N_6476,N_5627,N_5945);
and U6477 (N_6477,N_5790,N_5576);
or U6478 (N_6478,N_5656,N_5978);
nand U6479 (N_6479,N_5608,N_5976);
nand U6480 (N_6480,N_5700,N_5801);
nand U6481 (N_6481,N_5925,N_5755);
nor U6482 (N_6482,N_5815,N_5933);
nand U6483 (N_6483,N_5808,N_5548);
nand U6484 (N_6484,N_5678,N_5772);
nor U6485 (N_6485,N_5937,N_5508);
nand U6486 (N_6486,N_5541,N_5602);
or U6487 (N_6487,N_5597,N_5864);
and U6488 (N_6488,N_5572,N_5836);
or U6489 (N_6489,N_5735,N_5843);
nand U6490 (N_6490,N_5899,N_5958);
or U6491 (N_6491,N_5602,N_5952);
and U6492 (N_6492,N_5507,N_5505);
nor U6493 (N_6493,N_5920,N_5787);
or U6494 (N_6494,N_5528,N_5779);
and U6495 (N_6495,N_5557,N_5621);
or U6496 (N_6496,N_5795,N_5802);
nor U6497 (N_6497,N_5864,N_5730);
or U6498 (N_6498,N_5802,N_5711);
or U6499 (N_6499,N_5962,N_5625);
or U6500 (N_6500,N_6073,N_6149);
or U6501 (N_6501,N_6159,N_6053);
nand U6502 (N_6502,N_6030,N_6369);
xnor U6503 (N_6503,N_6274,N_6289);
nor U6504 (N_6504,N_6313,N_6119);
nand U6505 (N_6505,N_6206,N_6464);
and U6506 (N_6506,N_6096,N_6263);
nor U6507 (N_6507,N_6420,N_6423);
or U6508 (N_6508,N_6154,N_6403);
nand U6509 (N_6509,N_6430,N_6102);
and U6510 (N_6510,N_6110,N_6432);
nand U6511 (N_6511,N_6328,N_6434);
or U6512 (N_6512,N_6201,N_6390);
or U6513 (N_6513,N_6281,N_6287);
nor U6514 (N_6514,N_6439,N_6486);
nand U6515 (N_6515,N_6317,N_6142);
nor U6516 (N_6516,N_6008,N_6214);
nor U6517 (N_6517,N_6043,N_6334);
and U6518 (N_6518,N_6463,N_6202);
or U6519 (N_6519,N_6060,N_6185);
nand U6520 (N_6520,N_6271,N_6006);
nand U6521 (N_6521,N_6446,N_6231);
nor U6522 (N_6522,N_6057,N_6198);
or U6523 (N_6523,N_6347,N_6192);
xnor U6524 (N_6524,N_6194,N_6460);
nand U6525 (N_6525,N_6381,N_6478);
nor U6526 (N_6526,N_6078,N_6151);
nand U6527 (N_6527,N_6184,N_6356);
or U6528 (N_6528,N_6480,N_6071);
or U6529 (N_6529,N_6098,N_6324);
xnor U6530 (N_6530,N_6285,N_6384);
and U6531 (N_6531,N_6443,N_6130);
nor U6532 (N_6532,N_6092,N_6469);
or U6533 (N_6533,N_6150,N_6243);
nor U6534 (N_6534,N_6373,N_6445);
or U6535 (N_6535,N_6027,N_6134);
or U6536 (N_6536,N_6181,N_6321);
nand U6537 (N_6537,N_6459,N_6306);
and U6538 (N_6538,N_6264,N_6323);
nand U6539 (N_6539,N_6332,N_6056);
or U6540 (N_6540,N_6426,N_6409);
or U6541 (N_6541,N_6302,N_6031);
and U6542 (N_6542,N_6499,N_6496);
nand U6543 (N_6543,N_6303,N_6353);
or U6544 (N_6544,N_6273,N_6018);
and U6545 (N_6545,N_6166,N_6256);
xor U6546 (N_6546,N_6244,N_6153);
nor U6547 (N_6547,N_6229,N_6470);
and U6548 (N_6548,N_6000,N_6288);
or U6549 (N_6549,N_6492,N_6300);
nand U6550 (N_6550,N_6377,N_6010);
nand U6551 (N_6551,N_6455,N_6322);
nand U6552 (N_6552,N_6035,N_6396);
nor U6553 (N_6553,N_6065,N_6363);
nand U6554 (N_6554,N_6352,N_6419);
or U6555 (N_6555,N_6236,N_6029);
nand U6556 (N_6556,N_6069,N_6320);
nand U6557 (N_6557,N_6144,N_6022);
nor U6558 (N_6558,N_6415,N_6171);
nor U6559 (N_6559,N_6215,N_6160);
nand U6560 (N_6560,N_6136,N_6367);
nor U6561 (N_6561,N_6112,N_6371);
xnor U6562 (N_6562,N_6075,N_6090);
or U6563 (N_6563,N_6032,N_6345);
or U6564 (N_6564,N_6167,N_6168);
nor U6565 (N_6565,N_6079,N_6487);
nand U6566 (N_6566,N_6309,N_6392);
nand U6567 (N_6567,N_6483,N_6427);
xor U6568 (N_6568,N_6123,N_6195);
or U6569 (N_6569,N_6489,N_6210);
or U6570 (N_6570,N_6341,N_6205);
or U6571 (N_6571,N_6114,N_6041);
or U6572 (N_6572,N_6212,N_6174);
or U6573 (N_6573,N_6054,N_6380);
or U6574 (N_6574,N_6397,N_6133);
and U6575 (N_6575,N_6011,N_6466);
nand U6576 (N_6576,N_6132,N_6095);
nor U6577 (N_6577,N_6044,N_6180);
xnor U6578 (N_6578,N_6222,N_6346);
or U6579 (N_6579,N_6177,N_6226);
nor U6580 (N_6580,N_6479,N_6405);
nor U6581 (N_6581,N_6232,N_6428);
nand U6582 (N_6582,N_6218,N_6003);
nand U6583 (N_6583,N_6070,N_6002);
and U6584 (N_6584,N_6311,N_6333);
nand U6585 (N_6585,N_6351,N_6097);
or U6586 (N_6586,N_6389,N_6337);
nor U6587 (N_6587,N_6406,N_6276);
or U6588 (N_6588,N_6284,N_6196);
nor U6589 (N_6589,N_6137,N_6305);
nor U6590 (N_6590,N_6354,N_6152);
xor U6591 (N_6591,N_6083,N_6474);
xor U6592 (N_6592,N_6360,N_6355);
nor U6593 (N_6593,N_6211,N_6190);
or U6594 (N_6594,N_6146,N_6413);
or U6595 (N_6595,N_6485,N_6085);
nor U6596 (N_6596,N_6475,N_6424);
or U6597 (N_6597,N_6312,N_6339);
and U6598 (N_6598,N_6066,N_6183);
nand U6599 (N_6599,N_6316,N_6014);
nand U6600 (N_6600,N_6037,N_6265);
and U6601 (N_6601,N_6161,N_6051);
or U6602 (N_6602,N_6076,N_6310);
nor U6603 (N_6603,N_6441,N_6062);
and U6604 (N_6604,N_6047,N_6462);
nand U6605 (N_6605,N_6108,N_6219);
xnor U6606 (N_6606,N_6457,N_6366);
and U6607 (N_6607,N_6064,N_6275);
nor U6608 (N_6608,N_6178,N_6107);
nor U6609 (N_6609,N_6402,N_6128);
or U6610 (N_6610,N_6148,N_6453);
nand U6611 (N_6611,N_6417,N_6111);
nand U6612 (N_6612,N_6315,N_6291);
nor U6613 (N_6613,N_6401,N_6394);
or U6614 (N_6614,N_6141,N_6225);
and U6615 (N_6615,N_6127,N_6348);
nand U6616 (N_6616,N_6013,N_6370);
nor U6617 (N_6617,N_6407,N_6121);
and U6618 (N_6618,N_6458,N_6372);
nand U6619 (N_6619,N_6208,N_6145);
nand U6620 (N_6620,N_6314,N_6235);
nor U6621 (N_6621,N_6368,N_6042);
xor U6622 (N_6622,N_6498,N_6336);
and U6623 (N_6623,N_6262,N_6105);
xnor U6624 (N_6624,N_6376,N_6131);
and U6625 (N_6625,N_6259,N_6077);
nor U6626 (N_6626,N_6021,N_6290);
and U6627 (N_6627,N_6040,N_6036);
or U6628 (N_6628,N_6068,N_6143);
or U6629 (N_6629,N_6456,N_6468);
nor U6630 (N_6630,N_6307,N_6362);
nand U6631 (N_6631,N_6217,N_6220);
nand U6632 (N_6632,N_6412,N_6357);
and U6633 (N_6633,N_6237,N_6117);
and U6634 (N_6634,N_6452,N_6012);
and U6635 (N_6635,N_6228,N_6400);
nor U6636 (N_6636,N_6325,N_6282);
nor U6637 (N_6637,N_6147,N_6286);
xnor U6638 (N_6638,N_6129,N_6398);
or U6639 (N_6639,N_6388,N_6207);
nor U6640 (N_6640,N_6199,N_6484);
xor U6641 (N_6641,N_6074,N_6411);
or U6642 (N_6642,N_6138,N_6497);
and U6643 (N_6643,N_6422,N_6087);
nor U6644 (N_6644,N_6326,N_6279);
nand U6645 (N_6645,N_6327,N_6451);
nand U6646 (N_6646,N_6024,N_6182);
xor U6647 (N_6647,N_6017,N_6431);
nor U6648 (N_6648,N_6104,N_6239);
and U6649 (N_6649,N_6258,N_6113);
nor U6650 (N_6650,N_6476,N_6124);
nand U6651 (N_6651,N_6386,N_6209);
or U6652 (N_6652,N_6242,N_6319);
and U6653 (N_6653,N_6421,N_6408);
nor U6654 (N_6654,N_6465,N_6188);
nor U6655 (N_6655,N_6101,N_6296);
or U6656 (N_6656,N_6299,N_6193);
nand U6657 (N_6657,N_6100,N_6088);
and U6658 (N_6658,N_6488,N_6447);
xor U6659 (N_6659,N_6061,N_6046);
or U6660 (N_6660,N_6248,N_6416);
xor U6661 (N_6661,N_6072,N_6086);
or U6662 (N_6662,N_6039,N_6163);
xor U6663 (N_6663,N_6081,N_6358);
or U6664 (N_6664,N_6382,N_6364);
nand U6665 (N_6665,N_6454,N_6234);
or U6666 (N_6666,N_6301,N_6294);
and U6667 (N_6667,N_6126,N_6135);
nand U6668 (N_6668,N_6005,N_6467);
nand U6669 (N_6669,N_6254,N_6378);
xnor U6670 (N_6670,N_6444,N_6246);
or U6671 (N_6671,N_6089,N_6435);
and U6672 (N_6672,N_6058,N_6249);
or U6673 (N_6673,N_6442,N_6473);
nor U6674 (N_6674,N_6374,N_6034);
xnor U6675 (N_6675,N_6383,N_6280);
and U6676 (N_6676,N_6094,N_6349);
or U6677 (N_6677,N_6450,N_6247);
nand U6678 (N_6678,N_6395,N_6404);
nand U6679 (N_6679,N_6216,N_6429);
nor U6680 (N_6680,N_6385,N_6433);
and U6681 (N_6681,N_6245,N_6471);
nand U6682 (N_6682,N_6170,N_6391);
nor U6683 (N_6683,N_6266,N_6308);
xor U6684 (N_6684,N_6359,N_6350);
nand U6685 (N_6685,N_6493,N_6241);
nand U6686 (N_6686,N_6007,N_6257);
nor U6687 (N_6687,N_6204,N_6399);
nor U6688 (N_6688,N_6251,N_6261);
nand U6689 (N_6689,N_6140,N_6091);
nor U6690 (N_6690,N_6162,N_6270);
nor U6691 (N_6691,N_6344,N_6227);
or U6692 (N_6692,N_6001,N_6203);
nor U6693 (N_6693,N_6082,N_6187);
nor U6694 (N_6694,N_6223,N_6015);
and U6695 (N_6695,N_6033,N_6125);
and U6696 (N_6696,N_6268,N_6252);
and U6697 (N_6697,N_6048,N_6025);
or U6698 (N_6698,N_6109,N_6063);
nor U6699 (N_6699,N_6139,N_6331);
nor U6700 (N_6700,N_6318,N_6179);
and U6701 (N_6701,N_6267,N_6026);
nand U6702 (N_6702,N_6093,N_6490);
nand U6703 (N_6703,N_6293,N_6055);
and U6704 (N_6704,N_6297,N_6253);
nand U6705 (N_6705,N_6272,N_6186);
nor U6706 (N_6706,N_6375,N_6004);
or U6707 (N_6707,N_6414,N_6045);
xnor U6708 (N_6708,N_6436,N_6169);
nor U6709 (N_6709,N_6115,N_6292);
or U6710 (N_6710,N_6038,N_6295);
or U6711 (N_6711,N_6165,N_6304);
and U6712 (N_6712,N_6023,N_6365);
nand U6713 (N_6713,N_6418,N_6019);
xor U6714 (N_6714,N_6335,N_6052);
nor U6715 (N_6715,N_6298,N_6009);
or U6716 (N_6716,N_6449,N_6106);
and U6717 (N_6717,N_6156,N_6080);
nor U6718 (N_6718,N_6175,N_6116);
or U6719 (N_6719,N_6084,N_6269);
xor U6720 (N_6720,N_6338,N_6233);
or U6721 (N_6721,N_6437,N_6050);
nor U6722 (N_6722,N_6379,N_6250);
xnor U6723 (N_6723,N_6173,N_6238);
nand U6724 (N_6724,N_6067,N_6393);
or U6725 (N_6725,N_6277,N_6340);
nand U6726 (N_6726,N_6164,N_6197);
or U6727 (N_6727,N_6255,N_6118);
and U6728 (N_6728,N_6343,N_6122);
and U6729 (N_6729,N_6191,N_6278);
xnor U6730 (N_6730,N_6410,N_6482);
nand U6731 (N_6731,N_6472,N_6494);
or U6732 (N_6732,N_6329,N_6224);
nand U6733 (N_6733,N_6189,N_6260);
xnor U6734 (N_6734,N_6425,N_6016);
xor U6735 (N_6735,N_6221,N_6330);
nand U6736 (N_6736,N_6230,N_6020);
nor U6737 (N_6737,N_6481,N_6103);
nand U6738 (N_6738,N_6059,N_6387);
nor U6739 (N_6739,N_6440,N_6120);
nand U6740 (N_6740,N_6240,N_6448);
and U6741 (N_6741,N_6438,N_6176);
and U6742 (N_6742,N_6213,N_6361);
xor U6743 (N_6743,N_6200,N_6028);
nand U6744 (N_6744,N_6461,N_6049);
or U6745 (N_6745,N_6172,N_6491);
and U6746 (N_6746,N_6283,N_6495);
and U6747 (N_6747,N_6157,N_6158);
nor U6748 (N_6748,N_6099,N_6155);
or U6749 (N_6749,N_6477,N_6342);
or U6750 (N_6750,N_6299,N_6252);
and U6751 (N_6751,N_6488,N_6263);
nor U6752 (N_6752,N_6037,N_6473);
and U6753 (N_6753,N_6146,N_6026);
nand U6754 (N_6754,N_6116,N_6064);
and U6755 (N_6755,N_6039,N_6488);
and U6756 (N_6756,N_6125,N_6231);
nor U6757 (N_6757,N_6297,N_6172);
nand U6758 (N_6758,N_6232,N_6016);
or U6759 (N_6759,N_6257,N_6027);
nor U6760 (N_6760,N_6173,N_6183);
or U6761 (N_6761,N_6123,N_6287);
and U6762 (N_6762,N_6148,N_6379);
nor U6763 (N_6763,N_6229,N_6291);
nor U6764 (N_6764,N_6141,N_6142);
nand U6765 (N_6765,N_6319,N_6061);
nand U6766 (N_6766,N_6076,N_6382);
nand U6767 (N_6767,N_6053,N_6249);
nand U6768 (N_6768,N_6187,N_6283);
nor U6769 (N_6769,N_6337,N_6265);
or U6770 (N_6770,N_6255,N_6071);
nand U6771 (N_6771,N_6260,N_6322);
or U6772 (N_6772,N_6329,N_6185);
or U6773 (N_6773,N_6492,N_6380);
nand U6774 (N_6774,N_6019,N_6246);
and U6775 (N_6775,N_6172,N_6220);
or U6776 (N_6776,N_6307,N_6083);
nor U6777 (N_6777,N_6162,N_6338);
nand U6778 (N_6778,N_6229,N_6307);
and U6779 (N_6779,N_6457,N_6140);
nor U6780 (N_6780,N_6495,N_6458);
nor U6781 (N_6781,N_6430,N_6336);
or U6782 (N_6782,N_6010,N_6314);
or U6783 (N_6783,N_6192,N_6038);
nand U6784 (N_6784,N_6066,N_6104);
or U6785 (N_6785,N_6490,N_6481);
nor U6786 (N_6786,N_6142,N_6010);
nor U6787 (N_6787,N_6257,N_6107);
nor U6788 (N_6788,N_6476,N_6459);
nor U6789 (N_6789,N_6476,N_6027);
and U6790 (N_6790,N_6110,N_6012);
nand U6791 (N_6791,N_6447,N_6396);
and U6792 (N_6792,N_6446,N_6404);
nand U6793 (N_6793,N_6098,N_6176);
nand U6794 (N_6794,N_6388,N_6349);
nor U6795 (N_6795,N_6205,N_6398);
nand U6796 (N_6796,N_6458,N_6087);
or U6797 (N_6797,N_6237,N_6472);
nand U6798 (N_6798,N_6450,N_6477);
or U6799 (N_6799,N_6156,N_6055);
nor U6800 (N_6800,N_6260,N_6161);
nor U6801 (N_6801,N_6295,N_6020);
nand U6802 (N_6802,N_6096,N_6315);
nor U6803 (N_6803,N_6479,N_6174);
or U6804 (N_6804,N_6239,N_6313);
and U6805 (N_6805,N_6112,N_6117);
nor U6806 (N_6806,N_6049,N_6154);
nand U6807 (N_6807,N_6300,N_6275);
nor U6808 (N_6808,N_6088,N_6291);
nand U6809 (N_6809,N_6289,N_6055);
and U6810 (N_6810,N_6447,N_6067);
nor U6811 (N_6811,N_6383,N_6327);
or U6812 (N_6812,N_6049,N_6044);
or U6813 (N_6813,N_6028,N_6086);
and U6814 (N_6814,N_6442,N_6234);
and U6815 (N_6815,N_6312,N_6411);
nor U6816 (N_6816,N_6060,N_6433);
and U6817 (N_6817,N_6421,N_6119);
nand U6818 (N_6818,N_6133,N_6377);
or U6819 (N_6819,N_6383,N_6299);
or U6820 (N_6820,N_6252,N_6468);
or U6821 (N_6821,N_6367,N_6257);
nor U6822 (N_6822,N_6401,N_6460);
nand U6823 (N_6823,N_6183,N_6231);
xor U6824 (N_6824,N_6371,N_6456);
and U6825 (N_6825,N_6392,N_6121);
xor U6826 (N_6826,N_6077,N_6042);
or U6827 (N_6827,N_6103,N_6334);
and U6828 (N_6828,N_6188,N_6112);
or U6829 (N_6829,N_6008,N_6417);
and U6830 (N_6830,N_6422,N_6188);
nor U6831 (N_6831,N_6300,N_6385);
nand U6832 (N_6832,N_6119,N_6125);
nor U6833 (N_6833,N_6163,N_6217);
nor U6834 (N_6834,N_6099,N_6142);
nor U6835 (N_6835,N_6184,N_6015);
nand U6836 (N_6836,N_6239,N_6424);
and U6837 (N_6837,N_6316,N_6348);
or U6838 (N_6838,N_6197,N_6282);
and U6839 (N_6839,N_6149,N_6092);
nand U6840 (N_6840,N_6150,N_6460);
nor U6841 (N_6841,N_6115,N_6321);
or U6842 (N_6842,N_6218,N_6235);
nor U6843 (N_6843,N_6471,N_6380);
nand U6844 (N_6844,N_6477,N_6419);
and U6845 (N_6845,N_6230,N_6103);
nand U6846 (N_6846,N_6194,N_6128);
nor U6847 (N_6847,N_6023,N_6384);
nor U6848 (N_6848,N_6401,N_6101);
nor U6849 (N_6849,N_6450,N_6321);
and U6850 (N_6850,N_6395,N_6424);
nand U6851 (N_6851,N_6077,N_6371);
xor U6852 (N_6852,N_6367,N_6024);
or U6853 (N_6853,N_6113,N_6481);
or U6854 (N_6854,N_6373,N_6352);
nand U6855 (N_6855,N_6442,N_6323);
nor U6856 (N_6856,N_6103,N_6361);
and U6857 (N_6857,N_6018,N_6212);
and U6858 (N_6858,N_6363,N_6274);
nand U6859 (N_6859,N_6058,N_6032);
nor U6860 (N_6860,N_6447,N_6479);
and U6861 (N_6861,N_6069,N_6266);
or U6862 (N_6862,N_6086,N_6005);
xor U6863 (N_6863,N_6224,N_6283);
nor U6864 (N_6864,N_6420,N_6324);
or U6865 (N_6865,N_6243,N_6265);
nand U6866 (N_6866,N_6215,N_6406);
nand U6867 (N_6867,N_6044,N_6225);
and U6868 (N_6868,N_6419,N_6275);
xor U6869 (N_6869,N_6372,N_6337);
and U6870 (N_6870,N_6449,N_6437);
and U6871 (N_6871,N_6273,N_6258);
and U6872 (N_6872,N_6035,N_6031);
nor U6873 (N_6873,N_6115,N_6405);
nand U6874 (N_6874,N_6261,N_6104);
nand U6875 (N_6875,N_6425,N_6007);
nand U6876 (N_6876,N_6172,N_6439);
or U6877 (N_6877,N_6019,N_6357);
xor U6878 (N_6878,N_6408,N_6236);
xnor U6879 (N_6879,N_6370,N_6104);
nor U6880 (N_6880,N_6298,N_6030);
and U6881 (N_6881,N_6128,N_6258);
nand U6882 (N_6882,N_6295,N_6471);
and U6883 (N_6883,N_6276,N_6257);
and U6884 (N_6884,N_6418,N_6179);
nor U6885 (N_6885,N_6213,N_6373);
or U6886 (N_6886,N_6423,N_6044);
nand U6887 (N_6887,N_6250,N_6024);
nor U6888 (N_6888,N_6178,N_6267);
nand U6889 (N_6889,N_6019,N_6030);
nor U6890 (N_6890,N_6243,N_6402);
nand U6891 (N_6891,N_6312,N_6450);
nor U6892 (N_6892,N_6355,N_6499);
nor U6893 (N_6893,N_6394,N_6022);
or U6894 (N_6894,N_6486,N_6071);
nand U6895 (N_6895,N_6241,N_6002);
and U6896 (N_6896,N_6289,N_6327);
nor U6897 (N_6897,N_6376,N_6035);
nand U6898 (N_6898,N_6244,N_6260);
or U6899 (N_6899,N_6426,N_6183);
nor U6900 (N_6900,N_6433,N_6468);
and U6901 (N_6901,N_6280,N_6225);
nor U6902 (N_6902,N_6493,N_6379);
nor U6903 (N_6903,N_6273,N_6090);
and U6904 (N_6904,N_6216,N_6307);
xor U6905 (N_6905,N_6391,N_6212);
nand U6906 (N_6906,N_6038,N_6069);
xor U6907 (N_6907,N_6230,N_6037);
and U6908 (N_6908,N_6406,N_6404);
nor U6909 (N_6909,N_6279,N_6375);
nor U6910 (N_6910,N_6296,N_6431);
nor U6911 (N_6911,N_6428,N_6082);
xor U6912 (N_6912,N_6048,N_6244);
nand U6913 (N_6913,N_6134,N_6438);
nor U6914 (N_6914,N_6232,N_6111);
and U6915 (N_6915,N_6302,N_6174);
and U6916 (N_6916,N_6025,N_6429);
and U6917 (N_6917,N_6336,N_6494);
or U6918 (N_6918,N_6107,N_6210);
or U6919 (N_6919,N_6142,N_6046);
or U6920 (N_6920,N_6007,N_6126);
or U6921 (N_6921,N_6022,N_6042);
nor U6922 (N_6922,N_6202,N_6092);
or U6923 (N_6923,N_6073,N_6443);
and U6924 (N_6924,N_6343,N_6158);
nor U6925 (N_6925,N_6372,N_6205);
nand U6926 (N_6926,N_6114,N_6392);
and U6927 (N_6927,N_6427,N_6005);
or U6928 (N_6928,N_6298,N_6377);
and U6929 (N_6929,N_6430,N_6278);
or U6930 (N_6930,N_6350,N_6498);
nor U6931 (N_6931,N_6488,N_6016);
nor U6932 (N_6932,N_6382,N_6193);
xor U6933 (N_6933,N_6086,N_6266);
or U6934 (N_6934,N_6049,N_6011);
and U6935 (N_6935,N_6270,N_6359);
or U6936 (N_6936,N_6094,N_6492);
or U6937 (N_6937,N_6309,N_6035);
nor U6938 (N_6938,N_6432,N_6214);
and U6939 (N_6939,N_6402,N_6204);
or U6940 (N_6940,N_6351,N_6386);
xnor U6941 (N_6941,N_6384,N_6112);
and U6942 (N_6942,N_6220,N_6023);
xor U6943 (N_6943,N_6459,N_6427);
nor U6944 (N_6944,N_6094,N_6129);
xor U6945 (N_6945,N_6098,N_6002);
nand U6946 (N_6946,N_6244,N_6433);
and U6947 (N_6947,N_6499,N_6134);
nor U6948 (N_6948,N_6405,N_6247);
xnor U6949 (N_6949,N_6051,N_6427);
xnor U6950 (N_6950,N_6337,N_6420);
xor U6951 (N_6951,N_6180,N_6198);
and U6952 (N_6952,N_6318,N_6187);
nand U6953 (N_6953,N_6035,N_6040);
nand U6954 (N_6954,N_6071,N_6453);
nand U6955 (N_6955,N_6308,N_6497);
nand U6956 (N_6956,N_6412,N_6191);
nor U6957 (N_6957,N_6322,N_6456);
and U6958 (N_6958,N_6142,N_6261);
or U6959 (N_6959,N_6204,N_6274);
nor U6960 (N_6960,N_6206,N_6196);
nor U6961 (N_6961,N_6326,N_6110);
nand U6962 (N_6962,N_6018,N_6259);
nor U6963 (N_6963,N_6120,N_6239);
or U6964 (N_6964,N_6097,N_6481);
and U6965 (N_6965,N_6384,N_6195);
nor U6966 (N_6966,N_6379,N_6369);
nor U6967 (N_6967,N_6140,N_6386);
nand U6968 (N_6968,N_6215,N_6201);
or U6969 (N_6969,N_6427,N_6070);
or U6970 (N_6970,N_6367,N_6068);
nand U6971 (N_6971,N_6186,N_6075);
and U6972 (N_6972,N_6033,N_6283);
and U6973 (N_6973,N_6206,N_6184);
xor U6974 (N_6974,N_6337,N_6106);
and U6975 (N_6975,N_6232,N_6391);
nor U6976 (N_6976,N_6257,N_6135);
and U6977 (N_6977,N_6263,N_6356);
nand U6978 (N_6978,N_6036,N_6346);
xor U6979 (N_6979,N_6489,N_6337);
or U6980 (N_6980,N_6361,N_6349);
nand U6981 (N_6981,N_6054,N_6433);
nor U6982 (N_6982,N_6374,N_6458);
and U6983 (N_6983,N_6351,N_6016);
or U6984 (N_6984,N_6156,N_6372);
nand U6985 (N_6985,N_6005,N_6207);
or U6986 (N_6986,N_6379,N_6422);
nand U6987 (N_6987,N_6452,N_6125);
or U6988 (N_6988,N_6182,N_6432);
or U6989 (N_6989,N_6407,N_6311);
xor U6990 (N_6990,N_6124,N_6120);
nor U6991 (N_6991,N_6128,N_6137);
or U6992 (N_6992,N_6358,N_6085);
nand U6993 (N_6993,N_6362,N_6256);
and U6994 (N_6994,N_6102,N_6391);
nand U6995 (N_6995,N_6471,N_6272);
nor U6996 (N_6996,N_6283,N_6491);
and U6997 (N_6997,N_6132,N_6018);
and U6998 (N_6998,N_6356,N_6125);
nor U6999 (N_6999,N_6230,N_6039);
nor U7000 (N_7000,N_6806,N_6606);
and U7001 (N_7001,N_6711,N_6635);
or U7002 (N_7002,N_6738,N_6573);
nor U7003 (N_7003,N_6912,N_6589);
or U7004 (N_7004,N_6919,N_6845);
and U7005 (N_7005,N_6528,N_6637);
nand U7006 (N_7006,N_6581,N_6902);
and U7007 (N_7007,N_6855,N_6555);
or U7008 (N_7008,N_6934,N_6751);
or U7009 (N_7009,N_6976,N_6930);
or U7010 (N_7010,N_6772,N_6612);
nand U7011 (N_7011,N_6885,N_6697);
or U7012 (N_7012,N_6599,N_6915);
nor U7013 (N_7013,N_6675,N_6650);
nor U7014 (N_7014,N_6792,N_6770);
and U7015 (N_7015,N_6800,N_6516);
or U7016 (N_7016,N_6990,N_6506);
nor U7017 (N_7017,N_6859,N_6578);
nand U7018 (N_7018,N_6881,N_6672);
or U7019 (N_7019,N_6632,N_6636);
nor U7020 (N_7020,N_6793,N_6878);
and U7021 (N_7021,N_6674,N_6576);
or U7022 (N_7022,N_6744,N_6529);
nor U7023 (N_7023,N_6525,N_6535);
nand U7024 (N_7024,N_6691,N_6549);
nand U7025 (N_7025,N_6513,N_6510);
or U7026 (N_7026,N_6988,N_6960);
or U7027 (N_7027,N_6729,N_6822);
nand U7028 (N_7028,N_6821,N_6973);
and U7029 (N_7029,N_6896,N_6677);
or U7030 (N_7030,N_6785,N_6723);
or U7031 (N_7031,N_6541,N_6895);
or U7032 (N_7032,N_6783,N_6667);
and U7033 (N_7033,N_6634,N_6843);
or U7034 (N_7034,N_6561,N_6811);
nor U7035 (N_7035,N_6850,N_6907);
nor U7036 (N_7036,N_6605,N_6985);
or U7037 (N_7037,N_6730,N_6649);
xnor U7038 (N_7038,N_6903,N_6666);
xor U7039 (N_7039,N_6601,N_6777);
and U7040 (N_7040,N_6810,N_6813);
or U7041 (N_7041,N_6540,N_6998);
nor U7042 (N_7042,N_6608,N_6712);
or U7043 (N_7043,N_6921,N_6553);
nor U7044 (N_7044,N_6779,N_6773);
xnor U7045 (N_7045,N_6527,N_6786);
nor U7046 (N_7046,N_6820,N_6987);
nand U7047 (N_7047,N_6737,N_6966);
nand U7048 (N_7048,N_6898,N_6593);
nor U7049 (N_7049,N_6542,N_6518);
xor U7050 (N_7050,N_6630,N_6989);
nor U7051 (N_7051,N_6710,N_6787);
xnor U7052 (N_7052,N_6570,N_6782);
or U7053 (N_7053,N_6974,N_6798);
xor U7054 (N_7054,N_6877,N_6734);
or U7055 (N_7055,N_6586,N_6889);
nand U7056 (N_7056,N_6621,N_6847);
and U7057 (N_7057,N_6975,N_6696);
xor U7058 (N_7058,N_6836,N_6590);
xor U7059 (N_7059,N_6900,N_6757);
or U7060 (N_7060,N_6954,N_6834);
or U7061 (N_7061,N_6817,N_6548);
and U7062 (N_7062,N_6670,N_6550);
and U7063 (N_7063,N_6842,N_6687);
xor U7064 (N_7064,N_6685,N_6959);
and U7065 (N_7065,N_6695,N_6991);
nor U7066 (N_7066,N_6707,N_6673);
or U7067 (N_7067,N_6603,N_6888);
or U7068 (N_7068,N_6933,N_6764);
and U7069 (N_7069,N_6718,N_6940);
or U7070 (N_7070,N_6564,N_6926);
xor U7071 (N_7071,N_6882,N_6958);
and U7072 (N_7072,N_6755,N_6780);
nor U7073 (N_7073,N_6760,N_6676);
or U7074 (N_7074,N_6914,N_6699);
and U7075 (N_7075,N_6661,N_6501);
nand U7076 (N_7076,N_6962,N_6597);
and U7077 (N_7077,N_6981,N_6771);
nand U7078 (N_7078,N_6874,N_6828);
nand U7079 (N_7079,N_6722,N_6706);
nor U7080 (N_7080,N_6752,N_6514);
nor U7081 (N_7081,N_6747,N_6598);
nor U7082 (N_7082,N_6844,N_6731);
nand U7083 (N_7083,N_6862,N_6851);
nor U7084 (N_7084,N_6536,N_6922);
nand U7085 (N_7085,N_6524,N_6971);
or U7086 (N_7086,N_6665,N_6623);
nand U7087 (N_7087,N_6521,N_6716);
and U7088 (N_7088,N_6533,N_6887);
and U7089 (N_7089,N_6702,N_6538);
or U7090 (N_7090,N_6788,N_6663);
and U7091 (N_7091,N_6852,N_6965);
and U7092 (N_7092,N_6867,N_6897);
nand U7093 (N_7093,N_6617,N_6972);
or U7094 (N_7094,N_6761,N_6928);
nand U7095 (N_7095,N_6920,N_6567);
nor U7096 (N_7096,N_6993,N_6931);
or U7097 (N_7097,N_6583,N_6824);
nand U7098 (N_7098,N_6803,N_6908);
xnor U7099 (N_7099,N_6875,N_6544);
or U7100 (N_7100,N_6704,N_6886);
or U7101 (N_7101,N_6812,N_6656);
and U7102 (N_7102,N_6628,N_6776);
or U7103 (N_7103,N_6997,N_6618);
or U7104 (N_7104,N_6627,N_6577);
or U7105 (N_7105,N_6643,N_6502);
nand U7106 (N_7106,N_6853,N_6648);
nor U7107 (N_7107,N_6986,N_6584);
or U7108 (N_7108,N_6582,N_6652);
and U7109 (N_7109,N_6858,N_6999);
nand U7110 (N_7110,N_6551,N_6517);
or U7111 (N_7111,N_6728,N_6941);
xnor U7112 (N_7112,N_6591,N_6952);
xor U7113 (N_7113,N_6532,N_6996);
and U7114 (N_7114,N_6936,N_6951);
xnor U7115 (N_7115,N_6693,N_6899);
and U7116 (N_7116,N_6758,N_6864);
and U7117 (N_7117,N_6505,N_6511);
or U7118 (N_7118,N_6831,N_6778);
xor U7119 (N_7119,N_6805,N_6688);
nor U7120 (N_7120,N_6714,N_6560);
nand U7121 (N_7121,N_6840,N_6607);
and U7122 (N_7122,N_6733,N_6891);
nor U7123 (N_7123,N_6775,N_6917);
or U7124 (N_7124,N_6641,N_6507);
and U7125 (N_7125,N_6892,N_6841);
nand U7126 (N_7126,N_6816,N_6969);
nor U7127 (N_7127,N_6807,N_6742);
nand U7128 (N_7128,N_6943,N_6705);
nand U7129 (N_7129,N_6768,N_6592);
nand U7130 (N_7130,N_6503,N_6938);
nand U7131 (N_7131,N_6992,N_6614);
and U7132 (N_7132,N_6546,N_6537);
or U7133 (N_7133,N_6565,N_6715);
or U7134 (N_7134,N_6609,N_6748);
or U7135 (N_7135,N_6604,N_6616);
or U7136 (N_7136,N_6849,N_6935);
or U7137 (N_7137,N_6682,N_6745);
xnor U7138 (N_7138,N_6890,N_6789);
and U7139 (N_7139,N_6547,N_6825);
and U7140 (N_7140,N_6683,N_6808);
xnor U7141 (N_7141,N_6937,N_6569);
xnor U7142 (N_7142,N_6575,N_6644);
nand U7143 (N_7143,N_6719,N_6631);
nand U7144 (N_7144,N_6619,N_6512);
nor U7145 (N_7145,N_6504,N_6804);
and U7146 (N_7146,N_6963,N_6791);
nor U7147 (N_7147,N_6796,N_6689);
nand U7148 (N_7148,N_6995,N_6743);
or U7149 (N_7149,N_6911,N_6871);
nand U7150 (N_7150,N_6955,N_6563);
and U7151 (N_7151,N_6873,N_6880);
and U7152 (N_7152,N_6692,N_6658);
nor U7153 (N_7153,N_6982,N_6709);
or U7154 (N_7154,N_6700,N_6750);
and U7155 (N_7155,N_6918,N_6984);
or U7156 (N_7156,N_6949,N_6839);
xor U7157 (N_7157,N_6629,N_6508);
or U7158 (N_7158,N_6797,N_6732);
and U7159 (N_7159,N_6727,N_6756);
nor U7160 (N_7160,N_6657,N_6967);
or U7161 (N_7161,N_6901,N_6827);
nand U7162 (N_7162,N_6913,N_6762);
nand U7163 (N_7163,N_6556,N_6924);
nor U7164 (N_7164,N_6651,N_6659);
and U7165 (N_7165,N_6978,N_6884);
nor U7166 (N_7166,N_6894,N_6620);
or U7167 (N_7167,N_6708,N_6767);
nand U7168 (N_7168,N_6947,N_6678);
nor U7169 (N_7169,N_6579,N_6815);
nand U7170 (N_7170,N_6929,N_6879);
nand U7171 (N_7171,N_6814,N_6939);
nand U7172 (N_7172,N_6857,N_6863);
and U7173 (N_7173,N_6725,N_6686);
or U7174 (N_7174,N_6968,N_6713);
nor U7175 (N_7175,N_6876,N_6622);
and U7176 (N_7176,N_6945,N_6600);
and U7177 (N_7177,N_6753,N_6522);
or U7178 (N_7178,N_6534,N_6763);
and U7179 (N_7179,N_6653,N_6610);
nand U7180 (N_7180,N_6515,N_6979);
and U7181 (N_7181,N_6801,N_6646);
or U7182 (N_7182,N_6923,N_6594);
or U7183 (N_7183,N_6953,N_6662);
xnor U7184 (N_7184,N_6741,N_6749);
nand U7185 (N_7185,N_6950,N_6694);
nor U7186 (N_7186,N_6671,N_6531);
or U7187 (N_7187,N_6588,N_6856);
nor U7188 (N_7188,N_6909,N_6944);
nor U7189 (N_7189,N_6946,N_6829);
xor U7190 (N_7190,N_6654,N_6625);
nand U7191 (N_7191,N_6660,N_6872);
nand U7192 (N_7192,N_6554,N_6769);
nand U7193 (N_7193,N_6509,N_6765);
or U7194 (N_7194,N_6970,N_6848);
or U7195 (N_7195,N_6739,N_6595);
nand U7196 (N_7196,N_6860,N_6865);
nand U7197 (N_7197,N_6562,N_6558);
xor U7198 (N_7198,N_6956,N_6870);
nand U7199 (N_7199,N_6585,N_6559);
or U7200 (N_7200,N_6854,N_6526);
nor U7201 (N_7201,N_6680,N_6611);
or U7202 (N_7202,N_6639,N_6774);
nor U7203 (N_7203,N_6746,N_6754);
or U7204 (N_7204,N_6905,N_6964);
nor U7205 (N_7205,N_6566,N_6647);
nor U7206 (N_7206,N_6830,N_6596);
nor U7207 (N_7207,N_6906,N_6932);
nor U7208 (N_7208,N_6523,N_6642);
or U7209 (N_7209,N_6645,N_6519);
or U7210 (N_7210,N_6866,N_6655);
or U7211 (N_7211,N_6809,N_6698);
or U7212 (N_7212,N_6668,N_6818);
nor U7213 (N_7213,N_6961,N_6832);
or U7214 (N_7214,N_6690,N_6587);
xnor U7215 (N_7215,N_6568,N_6994);
or U7216 (N_7216,N_6861,N_6640);
or U7217 (N_7217,N_6846,N_6736);
nor U7218 (N_7218,N_6574,N_6983);
and U7219 (N_7219,N_6957,N_6927);
nand U7220 (N_7220,N_6826,N_6948);
nor U7221 (N_7221,N_6838,N_6543);
and U7222 (N_7222,N_6835,N_6703);
or U7223 (N_7223,N_6833,N_6545);
or U7224 (N_7224,N_6802,N_6819);
or U7225 (N_7225,N_6795,N_6624);
nor U7226 (N_7226,N_6500,N_6615);
and U7227 (N_7227,N_6664,N_6638);
and U7228 (N_7228,N_6980,N_6794);
and U7229 (N_7229,N_6681,N_6717);
nand U7230 (N_7230,N_6942,N_6613);
or U7231 (N_7231,N_6869,N_6684);
or U7232 (N_7232,N_6669,N_6580);
nand U7233 (N_7233,N_6823,N_6552);
or U7234 (N_7234,N_6977,N_6557);
or U7235 (N_7235,N_6735,N_6883);
nand U7236 (N_7236,N_6701,N_6781);
xor U7237 (N_7237,N_6799,N_6893);
or U7238 (N_7238,N_6626,N_6759);
xnor U7239 (N_7239,N_6726,N_6837);
xnor U7240 (N_7240,N_6740,N_6720);
nor U7241 (N_7241,N_6724,N_6679);
or U7242 (N_7242,N_6530,N_6916);
nor U7243 (N_7243,N_6520,N_6572);
or U7244 (N_7244,N_6925,N_6904);
or U7245 (N_7245,N_6790,N_6868);
xnor U7246 (N_7246,N_6721,N_6633);
or U7247 (N_7247,N_6766,N_6571);
nor U7248 (N_7248,N_6784,N_6539);
nor U7249 (N_7249,N_6602,N_6910);
and U7250 (N_7250,N_6953,N_6776);
and U7251 (N_7251,N_6535,N_6956);
nand U7252 (N_7252,N_6623,N_6891);
or U7253 (N_7253,N_6853,N_6825);
nor U7254 (N_7254,N_6878,N_6531);
or U7255 (N_7255,N_6877,N_6594);
nand U7256 (N_7256,N_6812,N_6657);
nor U7257 (N_7257,N_6655,N_6917);
and U7258 (N_7258,N_6502,N_6850);
and U7259 (N_7259,N_6844,N_6507);
nor U7260 (N_7260,N_6785,N_6886);
xnor U7261 (N_7261,N_6815,N_6757);
and U7262 (N_7262,N_6853,N_6856);
and U7263 (N_7263,N_6732,N_6632);
xor U7264 (N_7264,N_6805,N_6566);
nand U7265 (N_7265,N_6986,N_6792);
nor U7266 (N_7266,N_6893,N_6616);
xnor U7267 (N_7267,N_6500,N_6719);
xnor U7268 (N_7268,N_6792,N_6923);
and U7269 (N_7269,N_6661,N_6595);
nor U7270 (N_7270,N_6607,N_6883);
or U7271 (N_7271,N_6584,N_6773);
xnor U7272 (N_7272,N_6772,N_6645);
or U7273 (N_7273,N_6768,N_6719);
and U7274 (N_7274,N_6564,N_6969);
and U7275 (N_7275,N_6945,N_6527);
nand U7276 (N_7276,N_6810,N_6594);
nor U7277 (N_7277,N_6793,N_6685);
and U7278 (N_7278,N_6920,N_6728);
nand U7279 (N_7279,N_6613,N_6778);
xor U7280 (N_7280,N_6947,N_6716);
nand U7281 (N_7281,N_6731,N_6725);
nor U7282 (N_7282,N_6680,N_6959);
and U7283 (N_7283,N_6761,N_6712);
and U7284 (N_7284,N_6553,N_6801);
nor U7285 (N_7285,N_6845,N_6507);
nand U7286 (N_7286,N_6944,N_6596);
and U7287 (N_7287,N_6974,N_6864);
xor U7288 (N_7288,N_6866,N_6962);
nor U7289 (N_7289,N_6716,N_6900);
and U7290 (N_7290,N_6746,N_6970);
nor U7291 (N_7291,N_6561,N_6988);
nor U7292 (N_7292,N_6673,N_6541);
xor U7293 (N_7293,N_6881,N_6827);
nand U7294 (N_7294,N_6549,N_6958);
nor U7295 (N_7295,N_6606,N_6553);
and U7296 (N_7296,N_6618,N_6577);
nor U7297 (N_7297,N_6872,N_6978);
or U7298 (N_7298,N_6568,N_6830);
or U7299 (N_7299,N_6516,N_6746);
nand U7300 (N_7300,N_6817,N_6813);
nor U7301 (N_7301,N_6905,N_6686);
xnor U7302 (N_7302,N_6785,N_6808);
nand U7303 (N_7303,N_6725,N_6716);
or U7304 (N_7304,N_6726,N_6936);
or U7305 (N_7305,N_6931,N_6971);
nand U7306 (N_7306,N_6602,N_6872);
and U7307 (N_7307,N_6768,N_6827);
and U7308 (N_7308,N_6662,N_6758);
and U7309 (N_7309,N_6861,N_6769);
nor U7310 (N_7310,N_6502,N_6774);
or U7311 (N_7311,N_6858,N_6674);
xnor U7312 (N_7312,N_6737,N_6887);
and U7313 (N_7313,N_6825,N_6936);
and U7314 (N_7314,N_6871,N_6664);
and U7315 (N_7315,N_6526,N_6699);
and U7316 (N_7316,N_6892,N_6732);
and U7317 (N_7317,N_6717,N_6525);
nor U7318 (N_7318,N_6541,N_6871);
nand U7319 (N_7319,N_6846,N_6641);
nor U7320 (N_7320,N_6862,N_6511);
or U7321 (N_7321,N_6595,N_6871);
nor U7322 (N_7322,N_6552,N_6781);
or U7323 (N_7323,N_6834,N_6674);
and U7324 (N_7324,N_6956,N_6575);
nor U7325 (N_7325,N_6840,N_6610);
or U7326 (N_7326,N_6897,N_6728);
nand U7327 (N_7327,N_6594,N_6845);
nor U7328 (N_7328,N_6614,N_6928);
and U7329 (N_7329,N_6813,N_6863);
nor U7330 (N_7330,N_6905,N_6722);
nand U7331 (N_7331,N_6671,N_6604);
nand U7332 (N_7332,N_6875,N_6754);
xnor U7333 (N_7333,N_6596,N_6952);
nand U7334 (N_7334,N_6724,N_6823);
or U7335 (N_7335,N_6904,N_6962);
or U7336 (N_7336,N_6952,N_6921);
nor U7337 (N_7337,N_6587,N_6642);
or U7338 (N_7338,N_6699,N_6538);
nor U7339 (N_7339,N_6942,N_6593);
or U7340 (N_7340,N_6697,N_6822);
nand U7341 (N_7341,N_6646,N_6954);
and U7342 (N_7342,N_6671,N_6916);
nand U7343 (N_7343,N_6895,N_6865);
or U7344 (N_7344,N_6845,N_6591);
nand U7345 (N_7345,N_6638,N_6772);
and U7346 (N_7346,N_6972,N_6675);
nor U7347 (N_7347,N_6859,N_6787);
nor U7348 (N_7348,N_6574,N_6601);
and U7349 (N_7349,N_6876,N_6844);
nand U7350 (N_7350,N_6923,N_6696);
and U7351 (N_7351,N_6872,N_6886);
or U7352 (N_7352,N_6817,N_6975);
or U7353 (N_7353,N_6522,N_6842);
xor U7354 (N_7354,N_6847,N_6741);
and U7355 (N_7355,N_6584,N_6598);
nor U7356 (N_7356,N_6968,N_6896);
nor U7357 (N_7357,N_6964,N_6526);
nand U7358 (N_7358,N_6715,N_6751);
nor U7359 (N_7359,N_6975,N_6866);
xor U7360 (N_7360,N_6765,N_6929);
and U7361 (N_7361,N_6801,N_6942);
xnor U7362 (N_7362,N_6864,N_6876);
nor U7363 (N_7363,N_6748,N_6711);
and U7364 (N_7364,N_6737,N_6541);
and U7365 (N_7365,N_6529,N_6586);
nand U7366 (N_7366,N_6672,N_6898);
or U7367 (N_7367,N_6646,N_6598);
nor U7368 (N_7368,N_6927,N_6972);
nor U7369 (N_7369,N_6962,N_6648);
nor U7370 (N_7370,N_6943,N_6844);
or U7371 (N_7371,N_6943,N_6873);
nor U7372 (N_7372,N_6971,N_6930);
and U7373 (N_7373,N_6888,N_6914);
nand U7374 (N_7374,N_6805,N_6655);
nand U7375 (N_7375,N_6726,N_6833);
nor U7376 (N_7376,N_6545,N_6552);
or U7377 (N_7377,N_6804,N_6773);
nand U7378 (N_7378,N_6960,N_6838);
and U7379 (N_7379,N_6647,N_6817);
nor U7380 (N_7380,N_6924,N_6959);
or U7381 (N_7381,N_6592,N_6776);
nand U7382 (N_7382,N_6846,N_6649);
nand U7383 (N_7383,N_6657,N_6906);
nand U7384 (N_7384,N_6725,N_6746);
and U7385 (N_7385,N_6926,N_6746);
nand U7386 (N_7386,N_6943,N_6834);
or U7387 (N_7387,N_6918,N_6841);
nor U7388 (N_7388,N_6703,N_6864);
and U7389 (N_7389,N_6560,N_6981);
nand U7390 (N_7390,N_6641,N_6990);
nand U7391 (N_7391,N_6792,N_6991);
and U7392 (N_7392,N_6876,N_6939);
or U7393 (N_7393,N_6583,N_6826);
or U7394 (N_7394,N_6988,N_6835);
or U7395 (N_7395,N_6560,N_6742);
nor U7396 (N_7396,N_6619,N_6826);
or U7397 (N_7397,N_6743,N_6966);
or U7398 (N_7398,N_6539,N_6525);
or U7399 (N_7399,N_6528,N_6769);
nor U7400 (N_7400,N_6877,N_6785);
or U7401 (N_7401,N_6627,N_6696);
or U7402 (N_7402,N_6783,N_6505);
nand U7403 (N_7403,N_6638,N_6760);
or U7404 (N_7404,N_6838,N_6971);
nor U7405 (N_7405,N_6597,N_6712);
xnor U7406 (N_7406,N_6737,N_6956);
nor U7407 (N_7407,N_6950,N_6710);
xor U7408 (N_7408,N_6572,N_6810);
nand U7409 (N_7409,N_6505,N_6563);
or U7410 (N_7410,N_6621,N_6547);
or U7411 (N_7411,N_6869,N_6934);
or U7412 (N_7412,N_6731,N_6511);
and U7413 (N_7413,N_6816,N_6571);
or U7414 (N_7414,N_6539,N_6501);
nand U7415 (N_7415,N_6984,N_6865);
nor U7416 (N_7416,N_6998,N_6904);
nand U7417 (N_7417,N_6881,N_6519);
xor U7418 (N_7418,N_6786,N_6607);
or U7419 (N_7419,N_6568,N_6885);
and U7420 (N_7420,N_6893,N_6626);
xnor U7421 (N_7421,N_6879,N_6688);
or U7422 (N_7422,N_6863,N_6553);
nor U7423 (N_7423,N_6990,N_6563);
and U7424 (N_7424,N_6888,N_6840);
or U7425 (N_7425,N_6650,N_6809);
nor U7426 (N_7426,N_6990,N_6780);
nor U7427 (N_7427,N_6665,N_6533);
nor U7428 (N_7428,N_6684,N_6529);
or U7429 (N_7429,N_6871,N_6692);
or U7430 (N_7430,N_6811,N_6665);
nor U7431 (N_7431,N_6726,N_6999);
xor U7432 (N_7432,N_6727,N_6587);
and U7433 (N_7433,N_6967,N_6696);
or U7434 (N_7434,N_6513,N_6666);
or U7435 (N_7435,N_6776,N_6518);
nand U7436 (N_7436,N_6541,N_6547);
or U7437 (N_7437,N_6951,N_6847);
or U7438 (N_7438,N_6811,N_6615);
xor U7439 (N_7439,N_6768,N_6708);
or U7440 (N_7440,N_6830,N_6855);
nand U7441 (N_7441,N_6787,N_6688);
and U7442 (N_7442,N_6988,N_6756);
or U7443 (N_7443,N_6665,N_6580);
and U7444 (N_7444,N_6598,N_6620);
and U7445 (N_7445,N_6824,N_6826);
and U7446 (N_7446,N_6869,N_6593);
or U7447 (N_7447,N_6739,N_6627);
nand U7448 (N_7448,N_6773,N_6862);
nand U7449 (N_7449,N_6981,N_6722);
nand U7450 (N_7450,N_6991,N_6993);
nor U7451 (N_7451,N_6854,N_6637);
nor U7452 (N_7452,N_6820,N_6729);
nand U7453 (N_7453,N_6952,N_6603);
and U7454 (N_7454,N_6914,N_6688);
nand U7455 (N_7455,N_6953,N_6546);
nand U7456 (N_7456,N_6880,N_6613);
and U7457 (N_7457,N_6908,N_6661);
or U7458 (N_7458,N_6546,N_6780);
and U7459 (N_7459,N_6733,N_6746);
nor U7460 (N_7460,N_6730,N_6810);
and U7461 (N_7461,N_6547,N_6941);
nor U7462 (N_7462,N_6934,N_6746);
xnor U7463 (N_7463,N_6605,N_6546);
and U7464 (N_7464,N_6812,N_6510);
or U7465 (N_7465,N_6621,N_6734);
xor U7466 (N_7466,N_6738,N_6759);
nand U7467 (N_7467,N_6728,N_6501);
and U7468 (N_7468,N_6895,N_6946);
and U7469 (N_7469,N_6838,N_6900);
nand U7470 (N_7470,N_6938,N_6631);
or U7471 (N_7471,N_6661,N_6772);
nand U7472 (N_7472,N_6685,N_6619);
or U7473 (N_7473,N_6805,N_6952);
xor U7474 (N_7474,N_6872,N_6958);
xor U7475 (N_7475,N_6805,N_6505);
xnor U7476 (N_7476,N_6658,N_6994);
xnor U7477 (N_7477,N_6630,N_6594);
and U7478 (N_7478,N_6561,N_6850);
or U7479 (N_7479,N_6662,N_6549);
xnor U7480 (N_7480,N_6671,N_6841);
nor U7481 (N_7481,N_6893,N_6516);
or U7482 (N_7482,N_6701,N_6690);
xnor U7483 (N_7483,N_6763,N_6966);
or U7484 (N_7484,N_6902,N_6680);
nand U7485 (N_7485,N_6641,N_6971);
and U7486 (N_7486,N_6703,N_6829);
nor U7487 (N_7487,N_6897,N_6933);
and U7488 (N_7488,N_6661,N_6993);
or U7489 (N_7489,N_6815,N_6645);
or U7490 (N_7490,N_6566,N_6747);
and U7491 (N_7491,N_6699,N_6844);
or U7492 (N_7492,N_6529,N_6863);
and U7493 (N_7493,N_6626,N_6958);
and U7494 (N_7494,N_6669,N_6943);
nor U7495 (N_7495,N_6753,N_6536);
and U7496 (N_7496,N_6699,N_6745);
nor U7497 (N_7497,N_6782,N_6960);
nor U7498 (N_7498,N_6919,N_6938);
xnor U7499 (N_7499,N_6772,N_6756);
xor U7500 (N_7500,N_7084,N_7022);
and U7501 (N_7501,N_7449,N_7309);
nand U7502 (N_7502,N_7356,N_7214);
nand U7503 (N_7503,N_7135,N_7336);
nor U7504 (N_7504,N_7152,N_7430);
or U7505 (N_7505,N_7429,N_7381);
nand U7506 (N_7506,N_7434,N_7198);
and U7507 (N_7507,N_7141,N_7451);
nor U7508 (N_7508,N_7438,N_7377);
or U7509 (N_7509,N_7458,N_7019);
nor U7510 (N_7510,N_7357,N_7126);
nor U7511 (N_7511,N_7128,N_7024);
or U7512 (N_7512,N_7132,N_7111);
and U7513 (N_7513,N_7178,N_7319);
and U7514 (N_7514,N_7172,N_7042);
nand U7515 (N_7515,N_7065,N_7256);
nand U7516 (N_7516,N_7162,N_7064);
nand U7517 (N_7517,N_7026,N_7428);
and U7518 (N_7518,N_7410,N_7183);
nand U7519 (N_7519,N_7139,N_7484);
nand U7520 (N_7520,N_7032,N_7234);
nor U7521 (N_7521,N_7277,N_7237);
and U7522 (N_7522,N_7313,N_7071);
nand U7523 (N_7523,N_7292,N_7118);
and U7524 (N_7524,N_7415,N_7337);
nor U7525 (N_7525,N_7191,N_7279);
nor U7526 (N_7526,N_7268,N_7035);
nor U7527 (N_7527,N_7364,N_7348);
or U7528 (N_7528,N_7325,N_7460);
nand U7529 (N_7529,N_7366,N_7146);
and U7530 (N_7530,N_7184,N_7195);
nor U7531 (N_7531,N_7487,N_7383);
or U7532 (N_7532,N_7252,N_7243);
and U7533 (N_7533,N_7299,N_7359);
or U7534 (N_7534,N_7416,N_7029);
nor U7535 (N_7535,N_7335,N_7455);
nor U7536 (N_7536,N_7367,N_7002);
or U7537 (N_7537,N_7389,N_7239);
and U7538 (N_7538,N_7296,N_7280);
or U7539 (N_7539,N_7185,N_7499);
nor U7540 (N_7540,N_7267,N_7238);
nor U7541 (N_7541,N_7074,N_7161);
and U7542 (N_7542,N_7230,N_7261);
nor U7543 (N_7543,N_7350,N_7046);
nor U7544 (N_7544,N_7332,N_7173);
nand U7545 (N_7545,N_7082,N_7482);
xor U7546 (N_7546,N_7117,N_7331);
nand U7547 (N_7547,N_7355,N_7067);
and U7548 (N_7548,N_7113,N_7303);
xor U7549 (N_7549,N_7255,N_7311);
nand U7550 (N_7550,N_7121,N_7360);
and U7551 (N_7551,N_7246,N_7137);
nand U7552 (N_7552,N_7436,N_7119);
and U7553 (N_7553,N_7199,N_7180);
or U7554 (N_7554,N_7401,N_7260);
or U7555 (N_7555,N_7386,N_7147);
or U7556 (N_7556,N_7403,N_7140);
and U7557 (N_7557,N_7201,N_7495);
nand U7558 (N_7558,N_7101,N_7088);
nor U7559 (N_7559,N_7069,N_7008);
and U7560 (N_7560,N_7106,N_7073);
and U7561 (N_7561,N_7320,N_7054);
and U7562 (N_7562,N_7170,N_7225);
nor U7563 (N_7563,N_7131,N_7282);
nor U7564 (N_7564,N_7116,N_7354);
or U7565 (N_7565,N_7400,N_7248);
nor U7566 (N_7566,N_7154,N_7294);
and U7567 (N_7567,N_7276,N_7143);
and U7568 (N_7568,N_7473,N_7028);
nor U7569 (N_7569,N_7006,N_7109);
or U7570 (N_7570,N_7329,N_7258);
xor U7571 (N_7571,N_7417,N_7095);
xnor U7572 (N_7572,N_7156,N_7264);
and U7573 (N_7573,N_7130,N_7293);
or U7574 (N_7574,N_7150,N_7437);
or U7575 (N_7575,N_7070,N_7039);
or U7576 (N_7576,N_7058,N_7287);
or U7577 (N_7577,N_7457,N_7250);
or U7578 (N_7578,N_7012,N_7259);
nand U7579 (N_7579,N_7402,N_7194);
nor U7580 (N_7580,N_7440,N_7203);
nand U7581 (N_7581,N_7308,N_7052);
nand U7582 (N_7582,N_7371,N_7444);
nand U7583 (N_7583,N_7392,N_7425);
or U7584 (N_7584,N_7010,N_7466);
nor U7585 (N_7585,N_7391,N_7363);
xor U7586 (N_7586,N_7136,N_7323);
nand U7587 (N_7587,N_7398,N_7431);
nor U7588 (N_7588,N_7213,N_7091);
nor U7589 (N_7589,N_7212,N_7489);
or U7590 (N_7590,N_7447,N_7125);
nor U7591 (N_7591,N_7468,N_7343);
or U7592 (N_7592,N_7186,N_7376);
or U7593 (N_7593,N_7285,N_7060);
and U7594 (N_7594,N_7157,N_7483);
nor U7595 (N_7595,N_7291,N_7102);
and U7596 (N_7596,N_7247,N_7083);
and U7597 (N_7597,N_7159,N_7003);
nor U7598 (N_7598,N_7275,N_7000);
or U7599 (N_7599,N_7271,N_7253);
and U7600 (N_7600,N_7025,N_7314);
and U7601 (N_7601,N_7103,N_7200);
and U7602 (N_7602,N_7096,N_7066);
or U7603 (N_7603,N_7050,N_7413);
nand U7604 (N_7604,N_7051,N_7055);
and U7605 (N_7605,N_7472,N_7378);
nor U7606 (N_7606,N_7063,N_7433);
or U7607 (N_7607,N_7036,N_7441);
and U7608 (N_7608,N_7412,N_7189);
xor U7609 (N_7609,N_7228,N_7465);
or U7610 (N_7610,N_7420,N_7171);
nor U7611 (N_7611,N_7160,N_7009);
and U7612 (N_7612,N_7432,N_7474);
nand U7613 (N_7613,N_7094,N_7148);
or U7614 (N_7614,N_7344,N_7076);
nor U7615 (N_7615,N_7347,N_7016);
or U7616 (N_7616,N_7450,N_7404);
nand U7617 (N_7617,N_7182,N_7223);
nand U7618 (N_7618,N_7375,N_7321);
nand U7619 (N_7619,N_7215,N_7205);
and U7620 (N_7620,N_7075,N_7358);
or U7621 (N_7621,N_7176,N_7423);
nand U7622 (N_7622,N_7272,N_7089);
and U7623 (N_7623,N_7044,N_7001);
and U7624 (N_7624,N_7334,N_7476);
nor U7625 (N_7625,N_7369,N_7361);
or U7626 (N_7626,N_7164,N_7405);
nor U7627 (N_7627,N_7222,N_7013);
or U7628 (N_7628,N_7414,N_7167);
nor U7629 (N_7629,N_7351,N_7353);
nand U7630 (N_7630,N_7384,N_7079);
or U7631 (N_7631,N_7040,N_7333);
and U7632 (N_7632,N_7373,N_7494);
or U7633 (N_7633,N_7030,N_7077);
xnor U7634 (N_7634,N_7045,N_7057);
or U7635 (N_7635,N_7216,N_7396);
xnor U7636 (N_7636,N_7227,N_7453);
or U7637 (N_7637,N_7422,N_7219);
nand U7638 (N_7638,N_7339,N_7426);
xor U7639 (N_7639,N_7318,N_7244);
or U7640 (N_7640,N_7409,N_7210);
nor U7641 (N_7641,N_7442,N_7362);
nand U7642 (N_7642,N_7326,N_7007);
or U7643 (N_7643,N_7283,N_7493);
nand U7644 (N_7644,N_7341,N_7316);
nand U7645 (N_7645,N_7262,N_7078);
nand U7646 (N_7646,N_7048,N_7107);
nor U7647 (N_7647,N_7221,N_7491);
and U7648 (N_7648,N_7467,N_7123);
nand U7649 (N_7649,N_7390,N_7187);
nor U7650 (N_7650,N_7127,N_7481);
or U7651 (N_7651,N_7352,N_7249);
xor U7652 (N_7652,N_7427,N_7310);
nand U7653 (N_7653,N_7446,N_7245);
nand U7654 (N_7654,N_7174,N_7419);
nor U7655 (N_7655,N_7469,N_7011);
and U7656 (N_7656,N_7380,N_7115);
nand U7657 (N_7657,N_7317,N_7492);
and U7658 (N_7658,N_7454,N_7217);
or U7659 (N_7659,N_7462,N_7023);
nor U7660 (N_7660,N_7098,N_7105);
nor U7661 (N_7661,N_7211,N_7459);
or U7662 (N_7662,N_7181,N_7068);
and U7663 (N_7663,N_7100,N_7177);
and U7664 (N_7664,N_7004,N_7349);
nand U7665 (N_7665,N_7193,N_7328);
or U7666 (N_7666,N_7269,N_7163);
and U7667 (N_7667,N_7315,N_7153);
nor U7668 (N_7668,N_7497,N_7443);
nand U7669 (N_7669,N_7298,N_7397);
and U7670 (N_7670,N_7424,N_7448);
nor U7671 (N_7671,N_7059,N_7478);
or U7672 (N_7672,N_7486,N_7374);
nor U7673 (N_7673,N_7047,N_7122);
and U7674 (N_7674,N_7251,N_7220);
nand U7675 (N_7675,N_7477,N_7086);
nand U7676 (N_7676,N_7056,N_7169);
nor U7677 (N_7677,N_7190,N_7043);
and U7678 (N_7678,N_7072,N_7188);
and U7679 (N_7679,N_7295,N_7488);
nand U7680 (N_7680,N_7196,N_7471);
and U7681 (N_7681,N_7340,N_7470);
nand U7682 (N_7682,N_7439,N_7286);
nand U7683 (N_7683,N_7204,N_7061);
nor U7684 (N_7684,N_7209,N_7254);
nand U7685 (N_7685,N_7406,N_7192);
nor U7686 (N_7686,N_7155,N_7338);
nand U7687 (N_7687,N_7242,N_7490);
or U7688 (N_7688,N_7168,N_7005);
nand U7689 (N_7689,N_7290,N_7475);
nand U7690 (N_7690,N_7037,N_7281);
nor U7691 (N_7691,N_7456,N_7038);
or U7692 (N_7692,N_7085,N_7263);
and U7693 (N_7693,N_7099,N_7129);
or U7694 (N_7694,N_7020,N_7092);
nor U7695 (N_7695,N_7120,N_7330);
nor U7696 (N_7696,N_7158,N_7240);
or U7697 (N_7697,N_7452,N_7062);
nor U7698 (N_7698,N_7112,N_7151);
or U7699 (N_7699,N_7408,N_7202);
nor U7700 (N_7700,N_7265,N_7015);
nor U7701 (N_7701,N_7399,N_7093);
and U7702 (N_7702,N_7387,N_7346);
or U7703 (N_7703,N_7306,N_7418);
nand U7704 (N_7704,N_7485,N_7370);
nand U7705 (N_7705,N_7327,N_7395);
nand U7706 (N_7706,N_7270,N_7145);
nand U7707 (N_7707,N_7379,N_7226);
and U7708 (N_7708,N_7018,N_7388);
nor U7709 (N_7709,N_7104,N_7014);
nor U7710 (N_7710,N_7393,N_7017);
nor U7711 (N_7711,N_7053,N_7229);
and U7712 (N_7712,N_7034,N_7166);
and U7713 (N_7713,N_7394,N_7232);
and U7714 (N_7714,N_7461,N_7231);
and U7715 (N_7715,N_7097,N_7197);
or U7716 (N_7716,N_7411,N_7175);
or U7717 (N_7717,N_7049,N_7300);
or U7718 (N_7718,N_7307,N_7322);
nand U7719 (N_7719,N_7342,N_7297);
or U7720 (N_7720,N_7124,N_7273);
nand U7721 (N_7721,N_7288,N_7206);
xnor U7722 (N_7722,N_7033,N_7031);
and U7723 (N_7723,N_7266,N_7365);
nor U7724 (N_7724,N_7304,N_7110);
nor U7725 (N_7725,N_7027,N_7235);
nor U7726 (N_7726,N_7324,N_7345);
xor U7727 (N_7727,N_7368,N_7041);
nor U7728 (N_7728,N_7496,N_7144);
or U7729 (N_7729,N_7302,N_7312);
nand U7730 (N_7730,N_7257,N_7464);
xor U7731 (N_7731,N_7289,N_7278);
or U7732 (N_7732,N_7421,N_7372);
nand U7733 (N_7733,N_7133,N_7087);
nor U7734 (N_7734,N_7274,N_7165);
and U7735 (N_7735,N_7134,N_7149);
nand U7736 (N_7736,N_7305,N_7138);
nor U7737 (N_7737,N_7233,N_7179);
nand U7738 (N_7738,N_7301,N_7241);
or U7739 (N_7739,N_7498,N_7435);
nand U7740 (N_7740,N_7224,N_7479);
nor U7741 (N_7741,N_7081,N_7445);
and U7742 (N_7742,N_7142,N_7385);
nand U7743 (N_7743,N_7090,N_7407);
nor U7744 (N_7744,N_7080,N_7480);
and U7745 (N_7745,N_7114,N_7463);
or U7746 (N_7746,N_7207,N_7284);
nor U7747 (N_7747,N_7236,N_7208);
nand U7748 (N_7748,N_7108,N_7218);
nand U7749 (N_7749,N_7021,N_7382);
and U7750 (N_7750,N_7322,N_7330);
xor U7751 (N_7751,N_7186,N_7467);
xnor U7752 (N_7752,N_7007,N_7333);
xnor U7753 (N_7753,N_7318,N_7118);
and U7754 (N_7754,N_7303,N_7287);
and U7755 (N_7755,N_7149,N_7206);
or U7756 (N_7756,N_7322,N_7115);
and U7757 (N_7757,N_7245,N_7318);
nand U7758 (N_7758,N_7423,N_7005);
and U7759 (N_7759,N_7086,N_7388);
nand U7760 (N_7760,N_7071,N_7209);
nor U7761 (N_7761,N_7469,N_7186);
and U7762 (N_7762,N_7318,N_7022);
nor U7763 (N_7763,N_7318,N_7378);
nor U7764 (N_7764,N_7030,N_7159);
nand U7765 (N_7765,N_7287,N_7251);
and U7766 (N_7766,N_7006,N_7396);
nor U7767 (N_7767,N_7485,N_7473);
or U7768 (N_7768,N_7279,N_7398);
nand U7769 (N_7769,N_7459,N_7186);
nand U7770 (N_7770,N_7378,N_7391);
and U7771 (N_7771,N_7135,N_7053);
xor U7772 (N_7772,N_7203,N_7076);
and U7773 (N_7773,N_7391,N_7434);
and U7774 (N_7774,N_7479,N_7084);
and U7775 (N_7775,N_7454,N_7030);
nor U7776 (N_7776,N_7480,N_7386);
nor U7777 (N_7777,N_7147,N_7240);
nor U7778 (N_7778,N_7326,N_7195);
or U7779 (N_7779,N_7096,N_7251);
nor U7780 (N_7780,N_7155,N_7172);
or U7781 (N_7781,N_7150,N_7158);
nand U7782 (N_7782,N_7333,N_7495);
nor U7783 (N_7783,N_7360,N_7399);
nand U7784 (N_7784,N_7375,N_7058);
nand U7785 (N_7785,N_7246,N_7308);
and U7786 (N_7786,N_7281,N_7391);
and U7787 (N_7787,N_7123,N_7061);
nor U7788 (N_7788,N_7391,N_7493);
nor U7789 (N_7789,N_7334,N_7486);
or U7790 (N_7790,N_7165,N_7300);
nor U7791 (N_7791,N_7096,N_7471);
nor U7792 (N_7792,N_7275,N_7255);
and U7793 (N_7793,N_7277,N_7264);
or U7794 (N_7794,N_7157,N_7286);
or U7795 (N_7795,N_7192,N_7337);
xor U7796 (N_7796,N_7059,N_7189);
nand U7797 (N_7797,N_7195,N_7213);
and U7798 (N_7798,N_7166,N_7253);
or U7799 (N_7799,N_7098,N_7008);
nor U7800 (N_7800,N_7312,N_7118);
nand U7801 (N_7801,N_7346,N_7330);
and U7802 (N_7802,N_7085,N_7298);
or U7803 (N_7803,N_7090,N_7258);
nor U7804 (N_7804,N_7467,N_7142);
or U7805 (N_7805,N_7388,N_7199);
and U7806 (N_7806,N_7493,N_7458);
nand U7807 (N_7807,N_7016,N_7219);
nand U7808 (N_7808,N_7111,N_7415);
and U7809 (N_7809,N_7000,N_7014);
nor U7810 (N_7810,N_7133,N_7388);
xnor U7811 (N_7811,N_7486,N_7298);
and U7812 (N_7812,N_7485,N_7224);
nand U7813 (N_7813,N_7100,N_7232);
nand U7814 (N_7814,N_7355,N_7414);
nand U7815 (N_7815,N_7084,N_7105);
nand U7816 (N_7816,N_7340,N_7204);
nand U7817 (N_7817,N_7283,N_7130);
nand U7818 (N_7818,N_7466,N_7338);
nand U7819 (N_7819,N_7074,N_7398);
nor U7820 (N_7820,N_7319,N_7455);
or U7821 (N_7821,N_7042,N_7488);
nor U7822 (N_7822,N_7269,N_7064);
and U7823 (N_7823,N_7100,N_7031);
nor U7824 (N_7824,N_7159,N_7334);
and U7825 (N_7825,N_7174,N_7442);
nand U7826 (N_7826,N_7041,N_7253);
nor U7827 (N_7827,N_7430,N_7437);
and U7828 (N_7828,N_7467,N_7289);
xnor U7829 (N_7829,N_7393,N_7330);
and U7830 (N_7830,N_7094,N_7240);
or U7831 (N_7831,N_7365,N_7181);
nand U7832 (N_7832,N_7317,N_7345);
nand U7833 (N_7833,N_7358,N_7117);
nor U7834 (N_7834,N_7420,N_7408);
nand U7835 (N_7835,N_7440,N_7068);
and U7836 (N_7836,N_7435,N_7224);
and U7837 (N_7837,N_7156,N_7401);
nand U7838 (N_7838,N_7311,N_7173);
or U7839 (N_7839,N_7327,N_7287);
or U7840 (N_7840,N_7322,N_7266);
and U7841 (N_7841,N_7153,N_7244);
nor U7842 (N_7842,N_7351,N_7243);
nor U7843 (N_7843,N_7203,N_7048);
or U7844 (N_7844,N_7434,N_7272);
and U7845 (N_7845,N_7247,N_7384);
nor U7846 (N_7846,N_7019,N_7120);
nand U7847 (N_7847,N_7320,N_7495);
xnor U7848 (N_7848,N_7372,N_7208);
nor U7849 (N_7849,N_7283,N_7242);
nand U7850 (N_7850,N_7233,N_7007);
nand U7851 (N_7851,N_7455,N_7440);
and U7852 (N_7852,N_7338,N_7014);
or U7853 (N_7853,N_7172,N_7275);
nand U7854 (N_7854,N_7261,N_7405);
nor U7855 (N_7855,N_7446,N_7022);
and U7856 (N_7856,N_7470,N_7498);
nand U7857 (N_7857,N_7015,N_7370);
and U7858 (N_7858,N_7229,N_7119);
nor U7859 (N_7859,N_7314,N_7242);
and U7860 (N_7860,N_7286,N_7416);
nor U7861 (N_7861,N_7376,N_7009);
and U7862 (N_7862,N_7493,N_7266);
nand U7863 (N_7863,N_7424,N_7073);
nand U7864 (N_7864,N_7069,N_7028);
nand U7865 (N_7865,N_7366,N_7232);
xnor U7866 (N_7866,N_7155,N_7050);
or U7867 (N_7867,N_7367,N_7169);
nand U7868 (N_7868,N_7267,N_7100);
nor U7869 (N_7869,N_7144,N_7145);
and U7870 (N_7870,N_7234,N_7496);
nand U7871 (N_7871,N_7354,N_7053);
and U7872 (N_7872,N_7053,N_7104);
nand U7873 (N_7873,N_7498,N_7437);
xor U7874 (N_7874,N_7015,N_7452);
or U7875 (N_7875,N_7363,N_7481);
or U7876 (N_7876,N_7454,N_7226);
and U7877 (N_7877,N_7388,N_7439);
xnor U7878 (N_7878,N_7175,N_7302);
or U7879 (N_7879,N_7475,N_7494);
and U7880 (N_7880,N_7137,N_7223);
and U7881 (N_7881,N_7029,N_7373);
nand U7882 (N_7882,N_7017,N_7209);
nand U7883 (N_7883,N_7136,N_7294);
nor U7884 (N_7884,N_7184,N_7388);
nand U7885 (N_7885,N_7258,N_7361);
xnor U7886 (N_7886,N_7043,N_7362);
xor U7887 (N_7887,N_7022,N_7440);
and U7888 (N_7888,N_7101,N_7022);
nor U7889 (N_7889,N_7372,N_7494);
nand U7890 (N_7890,N_7435,N_7329);
xnor U7891 (N_7891,N_7425,N_7296);
nor U7892 (N_7892,N_7005,N_7057);
or U7893 (N_7893,N_7405,N_7182);
and U7894 (N_7894,N_7156,N_7464);
nor U7895 (N_7895,N_7090,N_7231);
nor U7896 (N_7896,N_7394,N_7130);
nor U7897 (N_7897,N_7431,N_7134);
xnor U7898 (N_7898,N_7322,N_7431);
nand U7899 (N_7899,N_7254,N_7136);
nand U7900 (N_7900,N_7273,N_7480);
and U7901 (N_7901,N_7420,N_7396);
nor U7902 (N_7902,N_7166,N_7387);
nor U7903 (N_7903,N_7300,N_7275);
or U7904 (N_7904,N_7172,N_7394);
nand U7905 (N_7905,N_7170,N_7018);
nand U7906 (N_7906,N_7157,N_7438);
or U7907 (N_7907,N_7028,N_7166);
nor U7908 (N_7908,N_7164,N_7173);
nor U7909 (N_7909,N_7426,N_7055);
or U7910 (N_7910,N_7419,N_7286);
nor U7911 (N_7911,N_7081,N_7297);
nand U7912 (N_7912,N_7358,N_7466);
and U7913 (N_7913,N_7025,N_7119);
and U7914 (N_7914,N_7441,N_7280);
or U7915 (N_7915,N_7457,N_7499);
nor U7916 (N_7916,N_7085,N_7035);
nor U7917 (N_7917,N_7204,N_7004);
and U7918 (N_7918,N_7389,N_7217);
and U7919 (N_7919,N_7200,N_7091);
and U7920 (N_7920,N_7172,N_7460);
and U7921 (N_7921,N_7431,N_7463);
nor U7922 (N_7922,N_7374,N_7316);
and U7923 (N_7923,N_7227,N_7037);
and U7924 (N_7924,N_7239,N_7312);
and U7925 (N_7925,N_7231,N_7330);
nand U7926 (N_7926,N_7442,N_7495);
nor U7927 (N_7927,N_7393,N_7464);
or U7928 (N_7928,N_7183,N_7076);
nor U7929 (N_7929,N_7283,N_7140);
and U7930 (N_7930,N_7081,N_7467);
and U7931 (N_7931,N_7310,N_7051);
xor U7932 (N_7932,N_7311,N_7137);
nand U7933 (N_7933,N_7033,N_7378);
and U7934 (N_7934,N_7487,N_7224);
nor U7935 (N_7935,N_7167,N_7243);
nor U7936 (N_7936,N_7308,N_7278);
nor U7937 (N_7937,N_7210,N_7054);
and U7938 (N_7938,N_7040,N_7194);
or U7939 (N_7939,N_7193,N_7444);
nand U7940 (N_7940,N_7208,N_7452);
or U7941 (N_7941,N_7287,N_7367);
and U7942 (N_7942,N_7158,N_7363);
and U7943 (N_7943,N_7278,N_7444);
or U7944 (N_7944,N_7041,N_7351);
or U7945 (N_7945,N_7099,N_7493);
xnor U7946 (N_7946,N_7427,N_7284);
and U7947 (N_7947,N_7310,N_7170);
or U7948 (N_7948,N_7218,N_7157);
nand U7949 (N_7949,N_7211,N_7484);
or U7950 (N_7950,N_7050,N_7019);
nor U7951 (N_7951,N_7142,N_7370);
and U7952 (N_7952,N_7441,N_7171);
and U7953 (N_7953,N_7315,N_7425);
nand U7954 (N_7954,N_7120,N_7423);
and U7955 (N_7955,N_7215,N_7411);
and U7956 (N_7956,N_7048,N_7444);
and U7957 (N_7957,N_7359,N_7317);
nor U7958 (N_7958,N_7052,N_7359);
nand U7959 (N_7959,N_7391,N_7185);
nand U7960 (N_7960,N_7158,N_7217);
or U7961 (N_7961,N_7295,N_7053);
and U7962 (N_7962,N_7022,N_7115);
xor U7963 (N_7963,N_7020,N_7110);
and U7964 (N_7964,N_7292,N_7013);
nor U7965 (N_7965,N_7096,N_7260);
nor U7966 (N_7966,N_7077,N_7406);
xnor U7967 (N_7967,N_7074,N_7068);
nor U7968 (N_7968,N_7054,N_7399);
nor U7969 (N_7969,N_7249,N_7396);
or U7970 (N_7970,N_7317,N_7423);
xor U7971 (N_7971,N_7476,N_7153);
nand U7972 (N_7972,N_7111,N_7065);
and U7973 (N_7973,N_7144,N_7107);
nand U7974 (N_7974,N_7412,N_7376);
or U7975 (N_7975,N_7086,N_7033);
or U7976 (N_7976,N_7427,N_7074);
or U7977 (N_7977,N_7405,N_7252);
and U7978 (N_7978,N_7093,N_7490);
nand U7979 (N_7979,N_7342,N_7352);
nand U7980 (N_7980,N_7435,N_7118);
nor U7981 (N_7981,N_7209,N_7048);
or U7982 (N_7982,N_7289,N_7196);
and U7983 (N_7983,N_7446,N_7070);
or U7984 (N_7984,N_7477,N_7084);
nand U7985 (N_7985,N_7032,N_7491);
nand U7986 (N_7986,N_7467,N_7324);
and U7987 (N_7987,N_7050,N_7304);
and U7988 (N_7988,N_7244,N_7272);
or U7989 (N_7989,N_7216,N_7245);
nand U7990 (N_7990,N_7337,N_7023);
nand U7991 (N_7991,N_7409,N_7079);
and U7992 (N_7992,N_7291,N_7223);
or U7993 (N_7993,N_7204,N_7444);
or U7994 (N_7994,N_7124,N_7247);
nand U7995 (N_7995,N_7201,N_7000);
and U7996 (N_7996,N_7316,N_7369);
or U7997 (N_7997,N_7306,N_7124);
nor U7998 (N_7998,N_7202,N_7479);
or U7999 (N_7999,N_7268,N_7093);
nor U8000 (N_8000,N_7907,N_7790);
nor U8001 (N_8001,N_7787,N_7829);
nor U8002 (N_8002,N_7624,N_7839);
or U8003 (N_8003,N_7658,N_7841);
nor U8004 (N_8004,N_7830,N_7634);
or U8005 (N_8005,N_7759,N_7855);
or U8006 (N_8006,N_7638,N_7568);
xnor U8007 (N_8007,N_7690,N_7663);
or U8008 (N_8008,N_7869,N_7898);
nor U8009 (N_8009,N_7604,N_7513);
or U8010 (N_8010,N_7552,N_7571);
xnor U8011 (N_8011,N_7609,N_7934);
or U8012 (N_8012,N_7861,N_7810);
and U8013 (N_8013,N_7626,N_7928);
xnor U8014 (N_8014,N_7915,N_7738);
nor U8015 (N_8015,N_7577,N_7742);
nand U8016 (N_8016,N_7923,N_7516);
and U8017 (N_8017,N_7851,N_7548);
or U8018 (N_8018,N_7677,N_7884);
or U8019 (N_8019,N_7675,N_7925);
nand U8020 (N_8020,N_7756,N_7909);
or U8021 (N_8021,N_7900,N_7801);
nand U8022 (N_8022,N_7969,N_7629);
nand U8023 (N_8023,N_7959,N_7671);
xor U8024 (N_8024,N_7992,N_7666);
nand U8025 (N_8025,N_7741,N_7961);
nor U8026 (N_8026,N_7795,N_7730);
and U8027 (N_8027,N_7501,N_7768);
or U8028 (N_8028,N_7797,N_7971);
and U8029 (N_8029,N_7650,N_7786);
or U8030 (N_8030,N_7581,N_7845);
xnor U8031 (N_8031,N_7957,N_7892);
nor U8032 (N_8032,N_7789,N_7942);
nor U8033 (N_8033,N_7659,N_7931);
or U8034 (N_8034,N_7937,N_7974);
and U8035 (N_8035,N_7550,N_7602);
nand U8036 (N_8036,N_7990,N_7968);
xor U8037 (N_8037,N_7733,N_7521);
or U8038 (N_8038,N_7509,N_7710);
xor U8039 (N_8039,N_7665,N_7958);
and U8040 (N_8040,N_7676,N_7922);
nor U8041 (N_8041,N_7570,N_7559);
nor U8042 (N_8042,N_7821,N_7582);
and U8043 (N_8043,N_7611,N_7938);
nor U8044 (N_8044,N_7960,N_7712);
and U8045 (N_8045,N_7988,N_7536);
nor U8046 (N_8046,N_7895,N_7586);
nor U8047 (N_8047,N_7952,N_7773);
nand U8048 (N_8048,N_7983,N_7596);
nand U8049 (N_8049,N_7963,N_7522);
nor U8050 (N_8050,N_7950,N_7860);
nand U8051 (N_8051,N_7554,N_7747);
or U8052 (N_8052,N_7679,N_7544);
nor U8053 (N_8053,N_7534,N_7887);
nand U8054 (N_8054,N_7635,N_7962);
and U8055 (N_8055,N_7966,N_7770);
nand U8056 (N_8056,N_7836,N_7893);
nor U8057 (N_8057,N_7930,N_7500);
nor U8058 (N_8058,N_7798,N_7914);
or U8059 (N_8059,N_7776,N_7538);
nand U8060 (N_8060,N_7902,N_7637);
nor U8061 (N_8061,N_7542,N_7881);
nand U8062 (N_8062,N_7653,N_7649);
nand U8063 (N_8063,N_7739,N_7504);
or U8064 (N_8064,N_7998,N_7728);
and U8065 (N_8065,N_7615,N_7751);
nor U8066 (N_8066,N_7796,N_7846);
nand U8067 (N_8067,N_7605,N_7965);
nor U8068 (N_8068,N_7578,N_7686);
and U8069 (N_8069,N_7600,N_7540);
and U8070 (N_8070,N_7744,N_7643);
xor U8071 (N_8071,N_7621,N_7802);
and U8072 (N_8072,N_7694,N_7867);
and U8073 (N_8073,N_7511,N_7834);
and U8074 (N_8074,N_7883,N_7720);
nand U8075 (N_8075,N_7817,N_7655);
nand U8076 (N_8076,N_7681,N_7535);
nand U8077 (N_8077,N_7627,N_7980);
nand U8078 (N_8078,N_7917,N_7619);
nor U8079 (N_8079,N_7606,N_7657);
xnor U8080 (N_8080,N_7953,N_7593);
nand U8081 (N_8081,N_7826,N_7858);
and U8082 (N_8082,N_7729,N_7654);
and U8083 (N_8083,N_7847,N_7644);
and U8084 (N_8084,N_7603,N_7889);
or U8085 (N_8085,N_7505,N_7954);
and U8086 (N_8086,N_7614,N_7631);
nor U8087 (N_8087,N_7967,N_7610);
nand U8088 (N_8088,N_7918,N_7986);
or U8089 (N_8089,N_7997,N_7981);
and U8090 (N_8090,N_7760,N_7857);
or U8091 (N_8091,N_7572,N_7612);
or U8092 (N_8092,N_7734,N_7926);
and U8093 (N_8093,N_7868,N_7678);
and U8094 (N_8094,N_7662,N_7775);
nor U8095 (N_8095,N_7890,N_7794);
nand U8096 (N_8096,N_7748,N_7780);
nand U8097 (N_8097,N_7667,N_7545);
nand U8098 (N_8098,N_7502,N_7749);
and U8099 (N_8099,N_7819,N_7716);
or U8100 (N_8100,N_7595,N_7987);
nand U8101 (N_8101,N_7639,N_7523);
and U8102 (N_8102,N_7707,N_7862);
nand U8103 (N_8103,N_7824,N_7680);
or U8104 (N_8104,N_7964,N_7708);
nand U8105 (N_8105,N_7685,N_7588);
and U8106 (N_8106,N_7706,N_7517);
nor U8107 (N_8107,N_7575,N_7592);
or U8108 (N_8108,N_7896,N_7921);
nor U8109 (N_8109,N_7555,N_7640);
and U8110 (N_8110,N_7779,N_7563);
nand U8111 (N_8111,N_7725,N_7850);
nand U8112 (N_8112,N_7806,N_7977);
and U8113 (N_8113,N_7723,N_7698);
nor U8114 (N_8114,N_7673,N_7804);
or U8115 (N_8115,N_7622,N_7558);
or U8116 (N_8116,N_7761,N_7837);
or U8117 (N_8117,N_7674,N_7731);
or U8118 (N_8118,N_7777,N_7539);
nor U8119 (N_8119,N_7908,N_7647);
or U8120 (N_8120,N_7785,N_7506);
nor U8121 (N_8121,N_7994,N_7863);
and U8122 (N_8122,N_7701,N_7591);
and U8123 (N_8123,N_7935,N_7507);
xor U8124 (N_8124,N_7510,N_7746);
or U8125 (N_8125,N_7519,N_7736);
and U8126 (N_8126,N_7689,N_7692);
xor U8127 (N_8127,N_7866,N_7633);
xnor U8128 (N_8128,N_7625,N_7813);
nand U8129 (N_8129,N_7993,N_7891);
and U8130 (N_8130,N_7842,N_7512);
or U8131 (N_8131,N_7745,N_7533);
or U8132 (N_8132,N_7995,N_7947);
or U8133 (N_8133,N_7515,N_7672);
nand U8134 (N_8134,N_7752,N_7929);
nand U8135 (N_8135,N_7835,N_7668);
or U8136 (N_8136,N_7771,N_7553);
nor U8137 (N_8137,N_7943,N_7878);
nand U8138 (N_8138,N_7503,N_7765);
and U8139 (N_8139,N_7549,N_7975);
nand U8140 (N_8140,N_7976,N_7583);
and U8141 (N_8141,N_7949,N_7946);
nand U8142 (N_8142,N_7541,N_7772);
nor U8143 (N_8143,N_7556,N_7576);
xor U8144 (N_8144,N_7764,N_7693);
nand U8145 (N_8145,N_7573,N_7715);
nand U8146 (N_8146,N_7562,N_7831);
xnor U8147 (N_8147,N_7551,N_7514);
and U8148 (N_8148,N_7816,N_7608);
xor U8149 (N_8149,N_7940,N_7955);
xnor U8150 (N_8150,N_7695,N_7880);
and U8151 (N_8151,N_7546,N_7901);
nand U8152 (N_8152,N_7856,N_7691);
or U8153 (N_8153,N_7941,N_7569);
or U8154 (N_8154,N_7956,N_7520);
and U8155 (N_8155,N_7597,N_7833);
or U8156 (N_8156,N_7853,N_7822);
or U8157 (N_8157,N_7973,N_7652);
nor U8158 (N_8158,N_7815,N_7778);
and U8159 (N_8159,N_7844,N_7670);
nor U8160 (N_8160,N_7788,N_7530);
nor U8161 (N_8161,N_7820,N_7948);
nand U8162 (N_8162,N_7913,N_7721);
and U8163 (N_8163,N_7740,N_7599);
xor U8164 (N_8164,N_7518,N_7899);
or U8165 (N_8165,N_7879,N_7601);
xor U8166 (N_8166,N_7714,N_7557);
nor U8167 (N_8167,N_7808,N_7528);
or U8168 (N_8168,N_7894,N_7832);
or U8169 (N_8169,N_7849,N_7618);
or U8170 (N_8170,N_7711,N_7924);
nand U8171 (N_8171,N_7565,N_7996);
nand U8172 (N_8172,N_7903,N_7970);
and U8173 (N_8173,N_7537,N_7783);
nand U8174 (N_8174,N_7607,N_7598);
nor U8175 (N_8175,N_7874,N_7805);
and U8176 (N_8176,N_7683,N_7628);
and U8177 (N_8177,N_7724,N_7766);
or U8178 (N_8178,N_7755,N_7508);
nor U8179 (N_8179,N_7916,N_7648);
nand U8180 (N_8180,N_7717,N_7905);
nor U8181 (N_8181,N_7718,N_7684);
or U8182 (N_8182,N_7774,N_7527);
nor U8183 (N_8183,N_7840,N_7933);
nor U8184 (N_8184,N_7561,N_7871);
nand U8185 (N_8185,N_7906,N_7623);
nand U8186 (N_8186,N_7656,N_7978);
and U8187 (N_8187,N_7696,N_7660);
and U8188 (N_8188,N_7753,N_7703);
nor U8189 (N_8189,N_7859,N_7985);
nor U8190 (N_8190,N_7543,N_7792);
or U8191 (N_8191,N_7632,N_7704);
or U8192 (N_8192,N_7864,N_7682);
or U8193 (N_8193,N_7594,N_7564);
or U8194 (N_8194,N_7574,N_7809);
nor U8195 (N_8195,N_7531,N_7828);
or U8196 (N_8196,N_7700,N_7727);
nor U8197 (N_8197,N_7877,N_7793);
or U8198 (N_8198,N_7807,N_7823);
or U8199 (N_8199,N_7566,N_7932);
or U8200 (N_8200,N_7873,N_7927);
or U8201 (N_8201,N_7646,N_7560);
nor U8202 (N_8202,N_7580,N_7547);
nor U8203 (N_8203,N_7636,N_7750);
xor U8204 (N_8204,N_7897,N_7945);
or U8205 (N_8205,N_7664,N_7782);
nand U8206 (N_8206,N_7910,N_7758);
nand U8207 (N_8207,N_7661,N_7584);
nor U8208 (N_8208,N_7617,N_7989);
nand U8209 (N_8209,N_7818,N_7722);
and U8210 (N_8210,N_7999,N_7825);
nand U8211 (N_8211,N_7767,N_7699);
and U8212 (N_8212,N_7920,N_7726);
or U8213 (N_8213,N_7791,N_7526);
or U8214 (N_8214,N_7882,N_7811);
and U8215 (N_8215,N_7743,N_7769);
or U8216 (N_8216,N_7800,N_7709);
nor U8217 (N_8217,N_7585,N_7843);
nor U8218 (N_8218,N_7529,N_7984);
and U8219 (N_8219,N_7944,N_7972);
and U8220 (N_8220,N_7757,N_7991);
nand U8221 (N_8221,N_7532,N_7904);
xnor U8222 (N_8222,N_7567,N_7936);
and U8223 (N_8223,N_7781,N_7705);
and U8224 (N_8224,N_7848,N_7763);
or U8225 (N_8225,N_7827,N_7911);
nor U8226 (N_8226,N_7838,N_7875);
or U8227 (N_8227,N_7630,N_7939);
and U8228 (N_8228,N_7951,N_7613);
nor U8229 (N_8229,N_7919,N_7888);
and U8230 (N_8230,N_7620,N_7737);
nand U8231 (N_8231,N_7697,N_7524);
nor U8232 (N_8232,N_7784,N_7669);
xor U8233 (N_8233,N_7713,N_7589);
nand U8234 (N_8234,N_7762,N_7886);
or U8235 (N_8235,N_7719,N_7735);
or U8236 (N_8236,N_7885,N_7642);
nand U8237 (N_8237,N_7645,N_7870);
or U8238 (N_8238,N_7799,N_7702);
nor U8239 (N_8239,N_7579,N_7912);
or U8240 (N_8240,N_7803,N_7876);
xor U8241 (N_8241,N_7754,N_7587);
or U8242 (N_8242,N_7854,N_7651);
and U8243 (N_8243,N_7641,N_7590);
xnor U8244 (N_8244,N_7732,N_7812);
nor U8245 (N_8245,N_7814,N_7616);
and U8246 (N_8246,N_7852,N_7982);
nand U8247 (N_8247,N_7865,N_7525);
nor U8248 (N_8248,N_7688,N_7687);
nand U8249 (N_8249,N_7979,N_7872);
nor U8250 (N_8250,N_7517,N_7549);
xor U8251 (N_8251,N_7892,N_7847);
or U8252 (N_8252,N_7605,N_7973);
or U8253 (N_8253,N_7793,N_7518);
xnor U8254 (N_8254,N_7841,N_7946);
or U8255 (N_8255,N_7592,N_7923);
or U8256 (N_8256,N_7658,N_7938);
nand U8257 (N_8257,N_7568,N_7946);
or U8258 (N_8258,N_7644,N_7662);
or U8259 (N_8259,N_7830,N_7823);
and U8260 (N_8260,N_7681,N_7649);
nor U8261 (N_8261,N_7574,N_7636);
nand U8262 (N_8262,N_7670,N_7706);
and U8263 (N_8263,N_7565,N_7918);
nor U8264 (N_8264,N_7678,N_7502);
and U8265 (N_8265,N_7847,N_7782);
nand U8266 (N_8266,N_7598,N_7621);
or U8267 (N_8267,N_7780,N_7538);
and U8268 (N_8268,N_7835,N_7815);
nor U8269 (N_8269,N_7545,N_7663);
and U8270 (N_8270,N_7500,N_7619);
and U8271 (N_8271,N_7725,N_7825);
and U8272 (N_8272,N_7594,N_7688);
and U8273 (N_8273,N_7595,N_7553);
or U8274 (N_8274,N_7910,N_7634);
nor U8275 (N_8275,N_7767,N_7686);
nand U8276 (N_8276,N_7986,N_7629);
or U8277 (N_8277,N_7955,N_7971);
or U8278 (N_8278,N_7590,N_7528);
nand U8279 (N_8279,N_7682,N_7563);
or U8280 (N_8280,N_7805,N_7985);
nor U8281 (N_8281,N_7904,N_7999);
or U8282 (N_8282,N_7583,N_7807);
nor U8283 (N_8283,N_7755,N_7531);
nor U8284 (N_8284,N_7916,N_7529);
and U8285 (N_8285,N_7613,N_7920);
or U8286 (N_8286,N_7911,N_7846);
nor U8287 (N_8287,N_7967,N_7966);
nor U8288 (N_8288,N_7959,N_7628);
nor U8289 (N_8289,N_7602,N_7566);
nand U8290 (N_8290,N_7706,N_7947);
or U8291 (N_8291,N_7650,N_7512);
and U8292 (N_8292,N_7692,N_7531);
nor U8293 (N_8293,N_7931,N_7854);
nor U8294 (N_8294,N_7925,N_7794);
or U8295 (N_8295,N_7621,N_7640);
nand U8296 (N_8296,N_7825,N_7927);
nand U8297 (N_8297,N_7813,N_7875);
xnor U8298 (N_8298,N_7956,N_7664);
nor U8299 (N_8299,N_7574,N_7645);
nor U8300 (N_8300,N_7633,N_7579);
or U8301 (N_8301,N_7898,N_7631);
and U8302 (N_8302,N_7635,N_7968);
or U8303 (N_8303,N_7901,N_7727);
nor U8304 (N_8304,N_7957,N_7731);
nor U8305 (N_8305,N_7879,N_7803);
or U8306 (N_8306,N_7501,N_7675);
nor U8307 (N_8307,N_7652,N_7596);
and U8308 (N_8308,N_7529,N_7689);
and U8309 (N_8309,N_7632,N_7716);
nand U8310 (N_8310,N_7938,N_7579);
nand U8311 (N_8311,N_7998,N_7801);
nand U8312 (N_8312,N_7908,N_7617);
or U8313 (N_8313,N_7896,N_7557);
and U8314 (N_8314,N_7522,N_7754);
and U8315 (N_8315,N_7584,N_7559);
or U8316 (N_8316,N_7505,N_7898);
and U8317 (N_8317,N_7632,N_7828);
or U8318 (N_8318,N_7611,N_7814);
and U8319 (N_8319,N_7878,N_7602);
and U8320 (N_8320,N_7813,N_7716);
nand U8321 (N_8321,N_7929,N_7614);
nand U8322 (N_8322,N_7696,N_7580);
nor U8323 (N_8323,N_7746,N_7686);
nor U8324 (N_8324,N_7876,N_7809);
nor U8325 (N_8325,N_7901,N_7517);
nand U8326 (N_8326,N_7688,N_7862);
and U8327 (N_8327,N_7559,N_7569);
and U8328 (N_8328,N_7792,N_7798);
nand U8329 (N_8329,N_7994,N_7641);
nor U8330 (N_8330,N_7878,N_7897);
and U8331 (N_8331,N_7514,N_7515);
or U8332 (N_8332,N_7724,N_7523);
and U8333 (N_8333,N_7535,N_7969);
and U8334 (N_8334,N_7512,N_7834);
and U8335 (N_8335,N_7721,N_7744);
xnor U8336 (N_8336,N_7865,N_7770);
nand U8337 (N_8337,N_7575,N_7548);
and U8338 (N_8338,N_7944,N_7865);
xnor U8339 (N_8339,N_7899,N_7748);
or U8340 (N_8340,N_7569,N_7807);
and U8341 (N_8341,N_7807,N_7906);
and U8342 (N_8342,N_7746,N_7568);
and U8343 (N_8343,N_7830,N_7901);
nand U8344 (N_8344,N_7610,N_7601);
nor U8345 (N_8345,N_7596,N_7733);
nor U8346 (N_8346,N_7522,N_7591);
xnor U8347 (N_8347,N_7811,N_7616);
and U8348 (N_8348,N_7594,N_7848);
xor U8349 (N_8349,N_7892,N_7776);
and U8350 (N_8350,N_7938,N_7846);
nand U8351 (N_8351,N_7974,N_7559);
and U8352 (N_8352,N_7761,N_7879);
nor U8353 (N_8353,N_7875,N_7582);
or U8354 (N_8354,N_7727,N_7773);
and U8355 (N_8355,N_7995,N_7538);
or U8356 (N_8356,N_7736,N_7981);
and U8357 (N_8357,N_7679,N_7978);
xnor U8358 (N_8358,N_7972,N_7923);
or U8359 (N_8359,N_7524,N_7633);
or U8360 (N_8360,N_7952,N_7893);
or U8361 (N_8361,N_7606,N_7904);
or U8362 (N_8362,N_7776,N_7743);
or U8363 (N_8363,N_7747,N_7896);
and U8364 (N_8364,N_7766,N_7956);
nand U8365 (N_8365,N_7909,N_7717);
nand U8366 (N_8366,N_7839,N_7735);
or U8367 (N_8367,N_7767,N_7746);
nand U8368 (N_8368,N_7942,N_7684);
xnor U8369 (N_8369,N_7856,N_7593);
nand U8370 (N_8370,N_7608,N_7713);
or U8371 (N_8371,N_7541,N_7524);
nand U8372 (N_8372,N_7979,N_7682);
nor U8373 (N_8373,N_7842,N_7920);
xnor U8374 (N_8374,N_7853,N_7703);
and U8375 (N_8375,N_7691,N_7916);
nand U8376 (N_8376,N_7667,N_7564);
nand U8377 (N_8377,N_7783,N_7825);
nor U8378 (N_8378,N_7508,N_7521);
nand U8379 (N_8379,N_7692,N_7856);
and U8380 (N_8380,N_7774,N_7868);
and U8381 (N_8381,N_7567,N_7623);
or U8382 (N_8382,N_7735,N_7754);
and U8383 (N_8383,N_7886,N_7786);
and U8384 (N_8384,N_7587,N_7858);
nor U8385 (N_8385,N_7719,N_7881);
or U8386 (N_8386,N_7832,N_7677);
nand U8387 (N_8387,N_7910,N_7883);
nand U8388 (N_8388,N_7541,N_7938);
nand U8389 (N_8389,N_7693,N_7679);
nand U8390 (N_8390,N_7826,N_7873);
nand U8391 (N_8391,N_7883,N_7708);
or U8392 (N_8392,N_7682,N_7765);
nor U8393 (N_8393,N_7760,N_7672);
and U8394 (N_8394,N_7833,N_7732);
or U8395 (N_8395,N_7865,N_7514);
xnor U8396 (N_8396,N_7967,N_7702);
nor U8397 (N_8397,N_7613,N_7532);
or U8398 (N_8398,N_7625,N_7629);
and U8399 (N_8399,N_7666,N_7879);
nor U8400 (N_8400,N_7704,N_7705);
and U8401 (N_8401,N_7776,N_7707);
xnor U8402 (N_8402,N_7868,N_7870);
nor U8403 (N_8403,N_7903,N_7796);
nand U8404 (N_8404,N_7854,N_7774);
and U8405 (N_8405,N_7809,N_7709);
and U8406 (N_8406,N_7946,N_7879);
and U8407 (N_8407,N_7672,N_7973);
nor U8408 (N_8408,N_7988,N_7957);
or U8409 (N_8409,N_7890,N_7796);
and U8410 (N_8410,N_7851,N_7691);
or U8411 (N_8411,N_7599,N_7626);
xor U8412 (N_8412,N_7677,N_7529);
or U8413 (N_8413,N_7602,N_7660);
nor U8414 (N_8414,N_7985,N_7973);
nor U8415 (N_8415,N_7543,N_7740);
nor U8416 (N_8416,N_7847,N_7751);
nor U8417 (N_8417,N_7708,N_7837);
nand U8418 (N_8418,N_7533,N_7739);
nor U8419 (N_8419,N_7563,N_7544);
xnor U8420 (N_8420,N_7825,N_7599);
nor U8421 (N_8421,N_7754,N_7686);
nor U8422 (N_8422,N_7730,N_7558);
xnor U8423 (N_8423,N_7664,N_7969);
nand U8424 (N_8424,N_7821,N_7752);
nand U8425 (N_8425,N_7677,N_7654);
xnor U8426 (N_8426,N_7508,N_7786);
and U8427 (N_8427,N_7595,N_7947);
nand U8428 (N_8428,N_7897,N_7990);
or U8429 (N_8429,N_7615,N_7678);
and U8430 (N_8430,N_7743,N_7668);
or U8431 (N_8431,N_7515,N_7933);
nor U8432 (N_8432,N_7536,N_7791);
or U8433 (N_8433,N_7929,N_7761);
and U8434 (N_8434,N_7790,N_7986);
nor U8435 (N_8435,N_7950,N_7895);
nor U8436 (N_8436,N_7679,N_7746);
and U8437 (N_8437,N_7989,N_7786);
nand U8438 (N_8438,N_7706,N_7660);
nor U8439 (N_8439,N_7580,N_7757);
or U8440 (N_8440,N_7606,N_7720);
nor U8441 (N_8441,N_7569,N_7738);
nand U8442 (N_8442,N_7736,N_7561);
and U8443 (N_8443,N_7767,N_7892);
xor U8444 (N_8444,N_7940,N_7791);
and U8445 (N_8445,N_7610,N_7778);
nand U8446 (N_8446,N_7965,N_7822);
nor U8447 (N_8447,N_7733,N_7915);
or U8448 (N_8448,N_7679,N_7552);
or U8449 (N_8449,N_7728,N_7868);
nand U8450 (N_8450,N_7803,N_7608);
nand U8451 (N_8451,N_7886,N_7811);
and U8452 (N_8452,N_7971,N_7999);
nand U8453 (N_8453,N_7799,N_7720);
or U8454 (N_8454,N_7995,N_7877);
and U8455 (N_8455,N_7724,N_7677);
nand U8456 (N_8456,N_7649,N_7834);
and U8457 (N_8457,N_7641,N_7887);
and U8458 (N_8458,N_7519,N_7692);
xnor U8459 (N_8459,N_7549,N_7773);
or U8460 (N_8460,N_7859,N_7940);
nand U8461 (N_8461,N_7519,N_7843);
nor U8462 (N_8462,N_7902,N_7910);
nand U8463 (N_8463,N_7917,N_7873);
nand U8464 (N_8464,N_7629,N_7976);
or U8465 (N_8465,N_7997,N_7622);
xnor U8466 (N_8466,N_7798,N_7592);
nand U8467 (N_8467,N_7901,N_7916);
and U8468 (N_8468,N_7526,N_7778);
and U8469 (N_8469,N_7751,N_7562);
and U8470 (N_8470,N_7931,N_7963);
nor U8471 (N_8471,N_7736,N_7532);
xor U8472 (N_8472,N_7647,N_7690);
nor U8473 (N_8473,N_7739,N_7972);
nor U8474 (N_8474,N_7641,N_7869);
nand U8475 (N_8475,N_7671,N_7952);
nor U8476 (N_8476,N_7974,N_7580);
and U8477 (N_8477,N_7975,N_7744);
nor U8478 (N_8478,N_7976,N_7567);
nor U8479 (N_8479,N_7771,N_7938);
or U8480 (N_8480,N_7971,N_7661);
and U8481 (N_8481,N_7683,N_7506);
or U8482 (N_8482,N_7548,N_7917);
xor U8483 (N_8483,N_7505,N_7890);
and U8484 (N_8484,N_7760,N_7791);
nand U8485 (N_8485,N_7686,N_7866);
nand U8486 (N_8486,N_7543,N_7680);
or U8487 (N_8487,N_7827,N_7536);
or U8488 (N_8488,N_7567,N_7854);
nor U8489 (N_8489,N_7964,N_7563);
nor U8490 (N_8490,N_7864,N_7553);
nand U8491 (N_8491,N_7617,N_7966);
nand U8492 (N_8492,N_7912,N_7885);
xnor U8493 (N_8493,N_7758,N_7978);
nand U8494 (N_8494,N_7755,N_7670);
xnor U8495 (N_8495,N_7855,N_7914);
and U8496 (N_8496,N_7809,N_7989);
xnor U8497 (N_8497,N_7939,N_7672);
or U8498 (N_8498,N_7829,N_7776);
nor U8499 (N_8499,N_7813,N_7517);
nand U8500 (N_8500,N_8368,N_8314);
nor U8501 (N_8501,N_8244,N_8457);
or U8502 (N_8502,N_8237,N_8485);
nand U8503 (N_8503,N_8075,N_8439);
nor U8504 (N_8504,N_8419,N_8252);
nand U8505 (N_8505,N_8498,N_8270);
nor U8506 (N_8506,N_8305,N_8293);
or U8507 (N_8507,N_8183,N_8353);
nand U8508 (N_8508,N_8335,N_8477);
or U8509 (N_8509,N_8054,N_8389);
nor U8510 (N_8510,N_8351,N_8259);
or U8511 (N_8511,N_8376,N_8068);
nand U8512 (N_8512,N_8303,N_8493);
nor U8513 (N_8513,N_8484,N_8324);
or U8514 (N_8514,N_8122,N_8312);
nand U8515 (N_8515,N_8042,N_8339);
nand U8516 (N_8516,N_8322,N_8474);
nor U8517 (N_8517,N_8003,N_8289);
or U8518 (N_8518,N_8230,N_8082);
nand U8519 (N_8519,N_8148,N_8408);
and U8520 (N_8520,N_8479,N_8436);
nor U8521 (N_8521,N_8106,N_8294);
nand U8522 (N_8522,N_8184,N_8275);
and U8523 (N_8523,N_8059,N_8381);
nand U8524 (N_8524,N_8402,N_8409);
nor U8525 (N_8525,N_8097,N_8220);
xnor U8526 (N_8526,N_8386,N_8251);
nor U8527 (N_8527,N_8115,N_8064);
and U8528 (N_8528,N_8354,N_8169);
nand U8529 (N_8529,N_8411,N_8022);
or U8530 (N_8530,N_8103,N_8154);
nand U8531 (N_8531,N_8048,N_8273);
nor U8532 (N_8532,N_8483,N_8205);
nand U8533 (N_8533,N_8213,N_8356);
or U8534 (N_8534,N_8456,N_8168);
or U8535 (N_8535,N_8362,N_8441);
and U8536 (N_8536,N_8188,N_8127);
xor U8537 (N_8537,N_8421,N_8131);
nand U8538 (N_8538,N_8399,N_8442);
nor U8539 (N_8539,N_8111,N_8041);
or U8540 (N_8540,N_8004,N_8038);
or U8541 (N_8541,N_8327,N_8152);
xor U8542 (N_8542,N_8228,N_8404);
or U8543 (N_8543,N_8373,N_8066);
and U8544 (N_8544,N_8211,N_8242);
nor U8545 (N_8545,N_8288,N_8145);
nor U8546 (N_8546,N_8491,N_8248);
nor U8547 (N_8547,N_8443,N_8124);
or U8548 (N_8548,N_8119,N_8412);
and U8549 (N_8549,N_8380,N_8088);
xnor U8550 (N_8550,N_8410,N_8050);
or U8551 (N_8551,N_8086,N_8212);
nor U8552 (N_8552,N_8463,N_8138);
nor U8553 (N_8553,N_8157,N_8151);
nand U8554 (N_8554,N_8297,N_8392);
or U8555 (N_8555,N_8300,N_8102);
xnor U8556 (N_8556,N_8290,N_8121);
or U8557 (N_8557,N_8174,N_8182);
xnor U8558 (N_8558,N_8378,N_8034);
and U8559 (N_8559,N_8197,N_8049);
and U8560 (N_8560,N_8241,N_8274);
and U8561 (N_8561,N_8489,N_8417);
nand U8562 (N_8562,N_8236,N_8391);
nor U8563 (N_8563,N_8018,N_8135);
or U8564 (N_8564,N_8454,N_8191);
nand U8565 (N_8565,N_8167,N_8393);
nand U8566 (N_8566,N_8001,N_8447);
and U8567 (N_8567,N_8079,N_8071);
or U8568 (N_8568,N_8318,N_8080);
nor U8569 (N_8569,N_8030,N_8438);
and U8570 (N_8570,N_8087,N_8229);
and U8571 (N_8571,N_8035,N_8146);
and U8572 (N_8572,N_8344,N_8023);
xnor U8573 (N_8573,N_8308,N_8199);
nand U8574 (N_8574,N_8451,N_8488);
or U8575 (N_8575,N_8461,N_8235);
or U8576 (N_8576,N_8254,N_8406);
nor U8577 (N_8577,N_8377,N_8178);
nand U8578 (N_8578,N_8480,N_8141);
nor U8579 (N_8579,N_8129,N_8219);
nor U8580 (N_8580,N_8139,N_8158);
nor U8581 (N_8581,N_8427,N_8470);
and U8582 (N_8582,N_8194,N_8435);
and U8583 (N_8583,N_8047,N_8346);
and U8584 (N_8584,N_8045,N_8341);
xor U8585 (N_8585,N_8223,N_8455);
nand U8586 (N_8586,N_8093,N_8434);
nor U8587 (N_8587,N_8026,N_8495);
nand U8588 (N_8588,N_8008,N_8025);
nor U8589 (N_8589,N_8187,N_8382);
or U8590 (N_8590,N_8063,N_8478);
nor U8591 (N_8591,N_8096,N_8195);
nand U8592 (N_8592,N_8134,N_8385);
nor U8593 (N_8593,N_8136,N_8216);
xnor U8594 (N_8594,N_8051,N_8343);
or U8595 (N_8595,N_8067,N_8285);
or U8596 (N_8596,N_8232,N_8143);
or U8597 (N_8597,N_8245,N_8217);
nor U8598 (N_8598,N_8331,N_8144);
nor U8599 (N_8599,N_8202,N_8125);
nor U8600 (N_8600,N_8165,N_8114);
nand U8601 (N_8601,N_8448,N_8269);
nand U8602 (N_8602,N_8361,N_8424);
or U8603 (N_8603,N_8070,N_8283);
or U8604 (N_8604,N_8072,N_8163);
nand U8605 (N_8605,N_8364,N_8415);
and U8606 (N_8606,N_8092,N_8462);
or U8607 (N_8607,N_8403,N_8091);
nand U8608 (N_8608,N_8348,N_8473);
nand U8609 (N_8609,N_8272,N_8420);
or U8610 (N_8610,N_8323,N_8112);
nand U8611 (N_8611,N_8400,N_8065);
nor U8612 (N_8612,N_8055,N_8175);
xnor U8613 (N_8613,N_8014,N_8425);
nand U8614 (N_8614,N_8328,N_8078);
nand U8615 (N_8615,N_8264,N_8372);
or U8616 (N_8616,N_8298,N_8043);
and U8617 (N_8617,N_8471,N_8350);
or U8618 (N_8618,N_8180,N_8428);
nor U8619 (N_8619,N_8494,N_8309);
nor U8620 (N_8620,N_8084,N_8161);
xnor U8621 (N_8621,N_8039,N_8299);
and U8622 (N_8622,N_8390,N_8028);
nand U8623 (N_8623,N_8370,N_8153);
or U8624 (N_8624,N_8329,N_8422);
or U8625 (N_8625,N_8384,N_8416);
or U8626 (N_8626,N_8053,N_8061);
xnor U8627 (N_8627,N_8388,N_8433);
nor U8628 (N_8628,N_8077,N_8398);
and U8629 (N_8629,N_8109,N_8010);
or U8630 (N_8630,N_8118,N_8164);
or U8631 (N_8631,N_8449,N_8257);
nor U8632 (N_8632,N_8396,N_8226);
and U8633 (N_8633,N_8209,N_8268);
and U8634 (N_8634,N_8155,N_8340);
nor U8635 (N_8635,N_8379,N_8414);
nand U8636 (N_8636,N_8450,N_8295);
or U8637 (N_8637,N_8181,N_8044);
nand U8638 (N_8638,N_8458,N_8040);
or U8639 (N_8639,N_8334,N_8429);
nand U8640 (N_8640,N_8058,N_8374);
xnor U8641 (N_8641,N_8365,N_8358);
nand U8642 (N_8642,N_8367,N_8267);
xor U8643 (N_8643,N_8200,N_8006);
nand U8644 (N_8644,N_8156,N_8342);
nor U8645 (N_8645,N_8375,N_8310);
nor U8646 (N_8646,N_8263,N_8233);
nand U8647 (N_8647,N_8407,N_8060);
or U8648 (N_8648,N_8446,N_8029);
or U8649 (N_8649,N_8487,N_8475);
and U8650 (N_8650,N_8037,N_8395);
nor U8651 (N_8651,N_8467,N_8304);
nand U8652 (N_8652,N_8240,N_8173);
nand U8653 (N_8653,N_8469,N_8418);
nand U8654 (N_8654,N_8401,N_8387);
or U8655 (N_8655,N_8214,N_8177);
nor U8656 (N_8656,N_8284,N_8117);
or U8657 (N_8657,N_8179,N_8198);
and U8658 (N_8658,N_8201,N_8052);
nand U8659 (N_8659,N_8325,N_8355);
nor U8660 (N_8660,N_8430,N_8371);
xor U8661 (N_8661,N_8464,N_8497);
and U8662 (N_8662,N_8405,N_8315);
or U8663 (N_8663,N_8215,N_8330);
and U8664 (N_8664,N_8332,N_8445);
xnor U8665 (N_8665,N_8476,N_8147);
nor U8666 (N_8666,N_8033,N_8130);
or U8667 (N_8667,N_8281,N_8221);
or U8668 (N_8668,N_8260,N_8224);
nand U8669 (N_8669,N_8286,N_8017);
nor U8670 (N_8670,N_8258,N_8255);
or U8671 (N_8671,N_8250,N_8444);
and U8672 (N_8672,N_8466,N_8397);
or U8673 (N_8673,N_8311,N_8481);
and U8674 (N_8674,N_8296,N_8486);
nand U8675 (N_8675,N_8262,N_8196);
nand U8676 (N_8676,N_8094,N_8247);
nor U8677 (N_8677,N_8291,N_8171);
and U8678 (N_8678,N_8265,N_8320);
nor U8679 (N_8679,N_8349,N_8062);
nand U8680 (N_8680,N_8120,N_8276);
xor U8681 (N_8681,N_8140,N_8015);
nand U8682 (N_8682,N_8316,N_8176);
or U8683 (N_8683,N_8278,N_8012);
and U8684 (N_8684,N_8021,N_8095);
or U8685 (N_8685,N_8036,N_8189);
and U8686 (N_8686,N_8437,N_8090);
nand U8687 (N_8687,N_8338,N_8207);
nand U8688 (N_8688,N_8204,N_8016);
xnor U8689 (N_8689,N_8027,N_8468);
and U8690 (N_8690,N_8032,N_8193);
or U8691 (N_8691,N_8359,N_8307);
nor U8692 (N_8692,N_8108,N_8317);
or U8693 (N_8693,N_8360,N_8142);
nor U8694 (N_8694,N_8019,N_8326);
nor U8695 (N_8695,N_8482,N_8472);
xnor U8696 (N_8696,N_8313,N_8496);
nor U8697 (N_8697,N_8302,N_8336);
nand U8698 (N_8698,N_8306,N_8266);
nand U8699 (N_8699,N_8105,N_8100);
nor U8700 (N_8700,N_8011,N_8192);
and U8701 (N_8701,N_8413,N_8347);
nand U8702 (N_8702,N_8225,N_8203);
or U8703 (N_8703,N_8031,N_8431);
nor U8704 (N_8704,N_8465,N_8170);
nor U8705 (N_8705,N_8459,N_8432);
and U8706 (N_8706,N_8005,N_8133);
and U8707 (N_8707,N_8277,N_8081);
and U8708 (N_8708,N_8218,N_8366);
nor U8709 (N_8709,N_8098,N_8186);
and U8710 (N_8710,N_8279,N_8249);
nor U8711 (N_8711,N_8089,N_8208);
or U8712 (N_8712,N_8185,N_8253);
and U8713 (N_8713,N_8292,N_8460);
xor U8714 (N_8714,N_8000,N_8099);
or U8715 (N_8715,N_8057,N_8007);
nand U8716 (N_8716,N_8256,N_8287);
or U8717 (N_8717,N_8107,N_8159);
nor U8718 (N_8718,N_8069,N_8352);
nand U8719 (N_8719,N_8162,N_8261);
and U8720 (N_8720,N_8490,N_8301);
nand U8721 (N_8721,N_8073,N_8020);
or U8722 (N_8722,N_8101,N_8210);
nor U8723 (N_8723,N_8222,N_8234);
or U8724 (N_8724,N_8126,N_8238);
nor U8725 (N_8725,N_8085,N_8357);
and U8726 (N_8726,N_8166,N_8319);
and U8727 (N_8727,N_8337,N_8076);
nor U8728 (N_8728,N_8110,N_8150);
nor U8729 (N_8729,N_8492,N_8453);
nand U8730 (N_8730,N_8132,N_8056);
xnor U8731 (N_8731,N_8452,N_8206);
nor U8732 (N_8732,N_8369,N_8002);
nand U8733 (N_8733,N_8160,N_8024);
nand U8734 (N_8734,N_8009,N_8280);
nor U8735 (N_8735,N_8046,N_8123);
nand U8736 (N_8736,N_8149,N_8282);
and U8737 (N_8737,N_8172,N_8227);
or U8738 (N_8738,N_8239,N_8013);
xor U8739 (N_8739,N_8231,N_8137);
xor U8740 (N_8740,N_8271,N_8104);
nand U8741 (N_8741,N_8440,N_8333);
nand U8742 (N_8742,N_8394,N_8243);
nand U8743 (N_8743,N_8113,N_8246);
and U8744 (N_8744,N_8083,N_8321);
nor U8745 (N_8745,N_8423,N_8190);
nor U8746 (N_8746,N_8383,N_8363);
nor U8747 (N_8747,N_8116,N_8345);
nand U8748 (N_8748,N_8074,N_8499);
and U8749 (N_8749,N_8426,N_8128);
nand U8750 (N_8750,N_8324,N_8194);
nor U8751 (N_8751,N_8129,N_8317);
and U8752 (N_8752,N_8000,N_8177);
nand U8753 (N_8753,N_8330,N_8155);
and U8754 (N_8754,N_8332,N_8094);
nand U8755 (N_8755,N_8271,N_8116);
or U8756 (N_8756,N_8255,N_8449);
and U8757 (N_8757,N_8086,N_8213);
nand U8758 (N_8758,N_8008,N_8354);
and U8759 (N_8759,N_8115,N_8446);
nor U8760 (N_8760,N_8275,N_8032);
nand U8761 (N_8761,N_8250,N_8091);
nor U8762 (N_8762,N_8334,N_8364);
nand U8763 (N_8763,N_8352,N_8486);
and U8764 (N_8764,N_8317,N_8300);
and U8765 (N_8765,N_8206,N_8205);
or U8766 (N_8766,N_8423,N_8049);
or U8767 (N_8767,N_8387,N_8353);
or U8768 (N_8768,N_8077,N_8075);
or U8769 (N_8769,N_8465,N_8264);
or U8770 (N_8770,N_8094,N_8355);
nor U8771 (N_8771,N_8042,N_8418);
or U8772 (N_8772,N_8317,N_8166);
and U8773 (N_8773,N_8265,N_8316);
and U8774 (N_8774,N_8110,N_8066);
or U8775 (N_8775,N_8362,N_8328);
or U8776 (N_8776,N_8169,N_8219);
nand U8777 (N_8777,N_8434,N_8198);
nand U8778 (N_8778,N_8325,N_8338);
or U8779 (N_8779,N_8341,N_8281);
and U8780 (N_8780,N_8084,N_8415);
or U8781 (N_8781,N_8388,N_8246);
nand U8782 (N_8782,N_8111,N_8122);
xnor U8783 (N_8783,N_8345,N_8211);
or U8784 (N_8784,N_8010,N_8387);
nand U8785 (N_8785,N_8021,N_8494);
nand U8786 (N_8786,N_8128,N_8191);
nand U8787 (N_8787,N_8007,N_8004);
and U8788 (N_8788,N_8218,N_8009);
or U8789 (N_8789,N_8442,N_8116);
nand U8790 (N_8790,N_8109,N_8007);
nor U8791 (N_8791,N_8070,N_8287);
and U8792 (N_8792,N_8035,N_8151);
or U8793 (N_8793,N_8111,N_8327);
or U8794 (N_8794,N_8109,N_8162);
and U8795 (N_8795,N_8433,N_8056);
nand U8796 (N_8796,N_8164,N_8137);
nor U8797 (N_8797,N_8232,N_8085);
or U8798 (N_8798,N_8409,N_8422);
xnor U8799 (N_8799,N_8379,N_8245);
xnor U8800 (N_8800,N_8184,N_8236);
or U8801 (N_8801,N_8196,N_8254);
nand U8802 (N_8802,N_8411,N_8185);
and U8803 (N_8803,N_8442,N_8077);
and U8804 (N_8804,N_8456,N_8290);
nor U8805 (N_8805,N_8032,N_8006);
nand U8806 (N_8806,N_8272,N_8350);
nor U8807 (N_8807,N_8177,N_8043);
nor U8808 (N_8808,N_8397,N_8151);
or U8809 (N_8809,N_8080,N_8461);
nor U8810 (N_8810,N_8404,N_8403);
nor U8811 (N_8811,N_8007,N_8480);
and U8812 (N_8812,N_8368,N_8119);
nor U8813 (N_8813,N_8162,N_8302);
or U8814 (N_8814,N_8227,N_8049);
or U8815 (N_8815,N_8352,N_8274);
or U8816 (N_8816,N_8233,N_8088);
or U8817 (N_8817,N_8021,N_8374);
and U8818 (N_8818,N_8173,N_8014);
or U8819 (N_8819,N_8133,N_8388);
nand U8820 (N_8820,N_8338,N_8213);
and U8821 (N_8821,N_8192,N_8415);
nand U8822 (N_8822,N_8353,N_8339);
nand U8823 (N_8823,N_8175,N_8035);
and U8824 (N_8824,N_8171,N_8485);
nor U8825 (N_8825,N_8073,N_8087);
or U8826 (N_8826,N_8083,N_8137);
nor U8827 (N_8827,N_8074,N_8180);
or U8828 (N_8828,N_8413,N_8490);
and U8829 (N_8829,N_8409,N_8017);
or U8830 (N_8830,N_8453,N_8099);
nor U8831 (N_8831,N_8398,N_8428);
or U8832 (N_8832,N_8105,N_8489);
and U8833 (N_8833,N_8197,N_8194);
and U8834 (N_8834,N_8335,N_8304);
nand U8835 (N_8835,N_8496,N_8119);
and U8836 (N_8836,N_8138,N_8136);
nand U8837 (N_8837,N_8352,N_8398);
xnor U8838 (N_8838,N_8359,N_8491);
xnor U8839 (N_8839,N_8453,N_8057);
and U8840 (N_8840,N_8244,N_8464);
or U8841 (N_8841,N_8195,N_8285);
nor U8842 (N_8842,N_8485,N_8233);
nand U8843 (N_8843,N_8307,N_8440);
nor U8844 (N_8844,N_8112,N_8440);
nor U8845 (N_8845,N_8417,N_8341);
nor U8846 (N_8846,N_8387,N_8384);
nand U8847 (N_8847,N_8127,N_8251);
xor U8848 (N_8848,N_8378,N_8172);
or U8849 (N_8849,N_8464,N_8249);
nor U8850 (N_8850,N_8190,N_8048);
and U8851 (N_8851,N_8108,N_8070);
and U8852 (N_8852,N_8458,N_8365);
nand U8853 (N_8853,N_8040,N_8340);
nor U8854 (N_8854,N_8109,N_8464);
and U8855 (N_8855,N_8396,N_8345);
nor U8856 (N_8856,N_8343,N_8075);
nand U8857 (N_8857,N_8213,N_8224);
nand U8858 (N_8858,N_8259,N_8412);
and U8859 (N_8859,N_8053,N_8035);
and U8860 (N_8860,N_8465,N_8081);
xor U8861 (N_8861,N_8224,N_8369);
or U8862 (N_8862,N_8078,N_8379);
xor U8863 (N_8863,N_8223,N_8031);
nor U8864 (N_8864,N_8370,N_8078);
or U8865 (N_8865,N_8459,N_8158);
and U8866 (N_8866,N_8014,N_8436);
and U8867 (N_8867,N_8131,N_8438);
nor U8868 (N_8868,N_8496,N_8393);
or U8869 (N_8869,N_8279,N_8107);
nor U8870 (N_8870,N_8071,N_8389);
nand U8871 (N_8871,N_8377,N_8095);
or U8872 (N_8872,N_8142,N_8464);
or U8873 (N_8873,N_8240,N_8243);
nor U8874 (N_8874,N_8052,N_8057);
and U8875 (N_8875,N_8103,N_8462);
nor U8876 (N_8876,N_8403,N_8414);
nand U8877 (N_8877,N_8302,N_8392);
xor U8878 (N_8878,N_8374,N_8056);
or U8879 (N_8879,N_8052,N_8303);
or U8880 (N_8880,N_8470,N_8376);
or U8881 (N_8881,N_8417,N_8345);
nor U8882 (N_8882,N_8054,N_8199);
nor U8883 (N_8883,N_8206,N_8415);
xnor U8884 (N_8884,N_8335,N_8340);
or U8885 (N_8885,N_8358,N_8442);
and U8886 (N_8886,N_8023,N_8303);
nor U8887 (N_8887,N_8278,N_8277);
xnor U8888 (N_8888,N_8185,N_8275);
nand U8889 (N_8889,N_8270,N_8002);
nand U8890 (N_8890,N_8100,N_8170);
and U8891 (N_8891,N_8029,N_8376);
nor U8892 (N_8892,N_8142,N_8395);
xor U8893 (N_8893,N_8464,N_8341);
xor U8894 (N_8894,N_8106,N_8009);
nor U8895 (N_8895,N_8473,N_8265);
or U8896 (N_8896,N_8345,N_8222);
nor U8897 (N_8897,N_8402,N_8383);
nand U8898 (N_8898,N_8030,N_8312);
or U8899 (N_8899,N_8325,N_8394);
and U8900 (N_8900,N_8311,N_8363);
xor U8901 (N_8901,N_8003,N_8207);
and U8902 (N_8902,N_8303,N_8441);
xnor U8903 (N_8903,N_8072,N_8022);
or U8904 (N_8904,N_8064,N_8181);
nand U8905 (N_8905,N_8493,N_8137);
and U8906 (N_8906,N_8030,N_8325);
nor U8907 (N_8907,N_8126,N_8419);
nor U8908 (N_8908,N_8413,N_8156);
nor U8909 (N_8909,N_8097,N_8280);
and U8910 (N_8910,N_8353,N_8415);
nor U8911 (N_8911,N_8362,N_8381);
nand U8912 (N_8912,N_8305,N_8489);
nand U8913 (N_8913,N_8131,N_8444);
or U8914 (N_8914,N_8217,N_8421);
nand U8915 (N_8915,N_8001,N_8206);
nor U8916 (N_8916,N_8008,N_8124);
or U8917 (N_8917,N_8275,N_8414);
nor U8918 (N_8918,N_8451,N_8339);
and U8919 (N_8919,N_8025,N_8287);
nand U8920 (N_8920,N_8463,N_8101);
xor U8921 (N_8921,N_8346,N_8113);
or U8922 (N_8922,N_8007,N_8219);
nand U8923 (N_8923,N_8151,N_8455);
nor U8924 (N_8924,N_8432,N_8373);
xnor U8925 (N_8925,N_8003,N_8084);
nor U8926 (N_8926,N_8343,N_8323);
xor U8927 (N_8927,N_8239,N_8012);
and U8928 (N_8928,N_8398,N_8191);
nor U8929 (N_8929,N_8385,N_8060);
xnor U8930 (N_8930,N_8224,N_8220);
and U8931 (N_8931,N_8150,N_8233);
nand U8932 (N_8932,N_8037,N_8209);
or U8933 (N_8933,N_8272,N_8143);
and U8934 (N_8934,N_8102,N_8205);
and U8935 (N_8935,N_8030,N_8059);
and U8936 (N_8936,N_8480,N_8032);
nor U8937 (N_8937,N_8206,N_8072);
nor U8938 (N_8938,N_8342,N_8010);
nor U8939 (N_8939,N_8324,N_8293);
nor U8940 (N_8940,N_8353,N_8154);
or U8941 (N_8941,N_8425,N_8295);
or U8942 (N_8942,N_8132,N_8077);
nand U8943 (N_8943,N_8149,N_8498);
nand U8944 (N_8944,N_8125,N_8004);
xor U8945 (N_8945,N_8033,N_8333);
nor U8946 (N_8946,N_8341,N_8362);
nand U8947 (N_8947,N_8164,N_8124);
nand U8948 (N_8948,N_8221,N_8131);
and U8949 (N_8949,N_8102,N_8037);
xor U8950 (N_8950,N_8286,N_8419);
and U8951 (N_8951,N_8079,N_8325);
nand U8952 (N_8952,N_8498,N_8045);
nor U8953 (N_8953,N_8196,N_8465);
xor U8954 (N_8954,N_8050,N_8133);
nand U8955 (N_8955,N_8283,N_8208);
and U8956 (N_8956,N_8273,N_8496);
xor U8957 (N_8957,N_8402,N_8312);
and U8958 (N_8958,N_8086,N_8350);
nand U8959 (N_8959,N_8034,N_8212);
nor U8960 (N_8960,N_8091,N_8043);
or U8961 (N_8961,N_8029,N_8035);
nand U8962 (N_8962,N_8050,N_8477);
xnor U8963 (N_8963,N_8243,N_8390);
xnor U8964 (N_8964,N_8083,N_8324);
and U8965 (N_8965,N_8131,N_8393);
or U8966 (N_8966,N_8297,N_8334);
and U8967 (N_8967,N_8049,N_8194);
and U8968 (N_8968,N_8359,N_8235);
nor U8969 (N_8969,N_8494,N_8340);
nand U8970 (N_8970,N_8417,N_8018);
nor U8971 (N_8971,N_8256,N_8379);
or U8972 (N_8972,N_8139,N_8321);
or U8973 (N_8973,N_8386,N_8423);
nand U8974 (N_8974,N_8487,N_8132);
nor U8975 (N_8975,N_8057,N_8324);
xnor U8976 (N_8976,N_8372,N_8473);
and U8977 (N_8977,N_8248,N_8125);
and U8978 (N_8978,N_8076,N_8456);
or U8979 (N_8979,N_8296,N_8077);
or U8980 (N_8980,N_8200,N_8206);
and U8981 (N_8981,N_8462,N_8164);
and U8982 (N_8982,N_8046,N_8207);
or U8983 (N_8983,N_8385,N_8390);
or U8984 (N_8984,N_8174,N_8373);
nor U8985 (N_8985,N_8351,N_8200);
nand U8986 (N_8986,N_8303,N_8372);
and U8987 (N_8987,N_8111,N_8087);
and U8988 (N_8988,N_8459,N_8149);
or U8989 (N_8989,N_8423,N_8440);
nor U8990 (N_8990,N_8474,N_8200);
and U8991 (N_8991,N_8389,N_8112);
nand U8992 (N_8992,N_8164,N_8297);
nand U8993 (N_8993,N_8262,N_8420);
nand U8994 (N_8994,N_8099,N_8176);
or U8995 (N_8995,N_8305,N_8195);
nand U8996 (N_8996,N_8151,N_8329);
and U8997 (N_8997,N_8141,N_8178);
nand U8998 (N_8998,N_8002,N_8013);
nand U8999 (N_8999,N_8317,N_8377);
or U9000 (N_9000,N_8604,N_8550);
xnor U9001 (N_9001,N_8869,N_8817);
nand U9002 (N_9002,N_8612,N_8665);
or U9003 (N_9003,N_8794,N_8706);
nor U9004 (N_9004,N_8579,N_8692);
nor U9005 (N_9005,N_8603,N_8867);
and U9006 (N_9006,N_8752,N_8978);
or U9007 (N_9007,N_8721,N_8703);
or U9008 (N_9008,N_8740,N_8924);
nor U9009 (N_9009,N_8517,N_8634);
or U9010 (N_9010,N_8667,N_8628);
and U9011 (N_9011,N_8576,N_8950);
nand U9012 (N_9012,N_8729,N_8904);
and U9013 (N_9013,N_8882,N_8972);
nor U9014 (N_9014,N_8563,N_8872);
nor U9015 (N_9015,N_8656,N_8544);
nand U9016 (N_9016,N_8553,N_8774);
xor U9017 (N_9017,N_8986,N_8501);
xnor U9018 (N_9018,N_8806,N_8961);
or U9019 (N_9019,N_8698,N_8596);
and U9020 (N_9020,N_8876,N_8556);
or U9021 (N_9021,N_8525,N_8808);
nor U9022 (N_9022,N_8963,N_8565);
nor U9023 (N_9023,N_8929,N_8696);
or U9024 (N_9024,N_8900,N_8688);
xnor U9025 (N_9025,N_8605,N_8773);
nand U9026 (N_9026,N_8502,N_8932);
and U9027 (N_9027,N_8850,N_8951);
and U9028 (N_9028,N_8888,N_8922);
xnor U9029 (N_9029,N_8673,N_8906);
xnor U9030 (N_9030,N_8877,N_8662);
nand U9031 (N_9031,N_8704,N_8680);
nor U9032 (N_9032,N_8562,N_8857);
nor U9033 (N_9033,N_8652,N_8657);
or U9034 (N_9034,N_8841,N_8871);
nor U9035 (N_9035,N_8883,N_8503);
or U9036 (N_9036,N_8761,N_8925);
xnor U9037 (N_9037,N_8754,N_8685);
nor U9038 (N_9038,N_8514,N_8573);
nor U9039 (N_9039,N_8779,N_8759);
or U9040 (N_9040,N_8608,N_8694);
and U9041 (N_9041,N_8725,N_8957);
xor U9042 (N_9042,N_8783,N_8560);
nor U9043 (N_9043,N_8899,N_8955);
xor U9044 (N_9044,N_8934,N_8549);
nand U9045 (N_9045,N_8901,N_8691);
and U9046 (N_9046,N_8510,N_8973);
nor U9047 (N_9047,N_8533,N_8585);
nand U9048 (N_9048,N_8791,N_8992);
or U9049 (N_9049,N_8661,N_8814);
nand U9050 (N_9050,N_8891,N_8545);
nor U9051 (N_9051,N_8918,N_8647);
and U9052 (N_9052,N_8923,N_8930);
and U9053 (N_9053,N_8728,N_8666);
nand U9054 (N_9054,N_8548,N_8640);
nand U9055 (N_9055,N_8860,N_8726);
nor U9056 (N_9056,N_8509,N_8919);
nor U9057 (N_9057,N_8587,N_8641);
nand U9058 (N_9058,N_8873,N_8559);
and U9059 (N_9059,N_8821,N_8663);
or U9060 (N_9060,N_8845,N_8700);
and U9061 (N_9061,N_8583,N_8572);
and U9062 (N_9062,N_8785,N_8539);
or U9063 (N_9063,N_8672,N_8720);
and U9064 (N_9064,N_8938,N_8574);
nor U9065 (N_9065,N_8552,N_8546);
and U9066 (N_9066,N_8832,N_8743);
and U9067 (N_9067,N_8724,N_8770);
nor U9068 (N_9068,N_8970,N_8898);
nor U9069 (N_9069,N_8926,N_8980);
nand U9070 (N_9070,N_8621,N_8982);
nand U9071 (N_9071,N_8920,N_8981);
or U9072 (N_9072,N_8683,N_8676);
or U9073 (N_9073,N_8829,N_8902);
or U9074 (N_9074,N_8797,N_8964);
nand U9075 (N_9075,N_8916,N_8717);
xnor U9076 (N_9076,N_8578,N_8983);
xor U9077 (N_9077,N_8772,N_8591);
nand U9078 (N_9078,N_8997,N_8831);
nand U9079 (N_9079,N_8936,N_8984);
or U9080 (N_9080,N_8781,N_8849);
xor U9081 (N_9081,N_8631,N_8646);
xor U9082 (N_9082,N_8554,N_8649);
nand U9083 (N_9083,N_8737,N_8610);
nor U9084 (N_9084,N_8912,N_8856);
nor U9085 (N_9085,N_8697,N_8713);
xnor U9086 (N_9086,N_8708,N_8942);
or U9087 (N_9087,N_8868,N_8810);
nor U9088 (N_9088,N_8727,N_8535);
nor U9089 (N_9089,N_8690,N_8854);
nor U9090 (N_9090,N_8753,N_8944);
nand U9091 (N_9091,N_8954,N_8760);
and U9092 (N_9092,N_8707,N_8522);
xnor U9093 (N_9093,N_8624,N_8588);
or U9094 (N_9094,N_8648,N_8568);
nor U9095 (N_9095,N_8506,N_8818);
and U9096 (N_9096,N_8626,N_8541);
nand U9097 (N_9097,N_8633,N_8990);
or U9098 (N_9098,N_8682,N_8968);
nor U9099 (N_9099,N_8619,N_8825);
and U9100 (N_9100,N_8755,N_8564);
or U9101 (N_9101,N_8865,N_8505);
xnor U9102 (N_9102,N_8630,N_8977);
nand U9103 (N_9103,N_8875,N_8594);
nor U9104 (N_9104,N_8846,N_8569);
or U9105 (N_9105,N_8967,N_8756);
nor U9106 (N_9106,N_8807,N_8824);
xor U9107 (N_9107,N_8835,N_8763);
or U9108 (N_9108,N_8879,N_8826);
and U9109 (N_9109,N_8532,N_8540);
and U9110 (N_9110,N_8567,N_8751);
and U9111 (N_9111,N_8892,N_8645);
or U9112 (N_9112,N_8622,N_8748);
or U9113 (N_9113,N_8827,N_8636);
xnor U9114 (N_9114,N_8796,N_8858);
nand U9115 (N_9115,N_8880,N_8538);
or U9116 (N_9116,N_8935,N_8803);
nor U9117 (N_9117,N_8693,N_8744);
xnor U9118 (N_9118,N_8999,N_8679);
nand U9119 (N_9119,N_8595,N_8758);
nor U9120 (N_9120,N_8609,N_8991);
and U9121 (N_9121,N_8575,N_8848);
xor U9122 (N_9122,N_8811,N_8577);
and U9123 (N_9123,N_8741,N_8953);
nand U9124 (N_9124,N_8805,N_8613);
nor U9125 (N_9125,N_8861,N_8611);
and U9126 (N_9126,N_8884,N_8927);
nand U9127 (N_9127,N_8701,N_8620);
and U9128 (N_9128,N_8976,N_8523);
or U9129 (N_9129,N_8838,N_8940);
or U9130 (N_9130,N_8776,N_8671);
xor U9131 (N_9131,N_8948,N_8946);
nor U9132 (N_9132,N_8536,N_8747);
and U9133 (N_9133,N_8528,N_8543);
nand U9134 (N_9134,N_8987,N_8716);
xor U9135 (N_9135,N_8784,N_8702);
and U9136 (N_9136,N_8718,N_8837);
and U9137 (N_9137,N_8952,N_8910);
and U9138 (N_9138,N_8750,N_8816);
or U9139 (N_9139,N_8639,N_8844);
nor U9140 (N_9140,N_8802,N_8788);
nor U9141 (N_9141,N_8943,N_8616);
nor U9142 (N_9142,N_8928,N_8589);
nand U9143 (N_9143,N_8600,N_8689);
or U9144 (N_9144,N_8766,N_8586);
and U9145 (N_9145,N_8714,N_8659);
or U9146 (N_9146,N_8602,N_8842);
nand U9147 (N_9147,N_8778,N_8520);
nand U9148 (N_9148,N_8813,N_8907);
and U9149 (N_9149,N_8732,N_8995);
or U9150 (N_9150,N_8722,N_8500);
xnor U9151 (N_9151,N_8915,N_8681);
nand U9152 (N_9152,N_8792,N_8668);
nand U9153 (N_9153,N_8705,N_8931);
or U9154 (N_9154,N_8921,N_8710);
nand U9155 (N_9155,N_8765,N_8699);
nand U9156 (N_9156,N_8911,N_8993);
nand U9157 (N_9157,N_8733,N_8775);
nor U9158 (N_9158,N_8513,N_8833);
nor U9159 (N_9159,N_8996,N_8745);
or U9160 (N_9160,N_8917,N_8551);
nand U9161 (N_9161,N_8994,N_8599);
or U9162 (N_9162,N_8593,N_8787);
and U9163 (N_9163,N_8767,N_8966);
nor U9164 (N_9164,N_8903,N_8804);
nand U9165 (N_9165,N_8905,N_8885);
or U9166 (N_9166,N_8859,N_8895);
or U9167 (N_9167,N_8653,N_8843);
nor U9168 (N_9168,N_8937,N_8998);
or U9169 (N_9169,N_8945,N_8746);
or U9170 (N_9170,N_8512,N_8530);
nand U9171 (N_9171,N_8819,N_8913);
nor U9172 (N_9172,N_8786,N_8584);
or U9173 (N_9173,N_8637,N_8870);
nor U9174 (N_9174,N_8780,N_8985);
and U9175 (N_9175,N_8988,N_8894);
xor U9176 (N_9176,N_8508,N_8719);
or U9177 (N_9177,N_8547,N_8504);
nor U9178 (N_9178,N_8909,N_8557);
or U9179 (N_9179,N_8592,N_8615);
or U9180 (N_9180,N_8762,N_8852);
nor U9181 (N_9181,N_8828,N_8798);
or U9182 (N_9182,N_8558,N_8643);
nand U9183 (N_9183,N_8855,N_8555);
or U9184 (N_9184,N_8534,N_8887);
and U9185 (N_9185,N_8851,N_8969);
xor U9186 (N_9186,N_8670,N_8625);
and U9187 (N_9187,N_8958,N_8542);
or U9188 (N_9188,N_8830,N_8820);
and U9189 (N_9189,N_8782,N_8581);
or U9190 (N_9190,N_8658,N_8878);
and U9191 (N_9191,N_8777,N_8635);
nand U9192 (N_9192,N_8715,N_8711);
and U9193 (N_9193,N_8979,N_8939);
and U9194 (N_9194,N_8874,N_8655);
and U9195 (N_9195,N_8566,N_8960);
nand U9196 (N_9196,N_8956,N_8511);
or U9197 (N_9197,N_8650,N_8801);
nand U9198 (N_9198,N_8896,N_8933);
and U9199 (N_9199,N_8823,N_8949);
and U9200 (N_9200,N_8739,N_8597);
nor U9201 (N_9201,N_8771,N_8709);
nor U9202 (N_9202,N_8742,N_8764);
xor U9203 (N_9203,N_8526,N_8974);
or U9204 (N_9204,N_8614,N_8590);
and U9205 (N_9205,N_8730,N_8521);
or U9206 (N_9206,N_8840,N_8893);
and U9207 (N_9207,N_8686,N_8723);
xor U9208 (N_9208,N_8736,N_8678);
nand U9209 (N_9209,N_8795,N_8757);
nand U9210 (N_9210,N_8527,N_8617);
nor U9211 (N_9211,N_8606,N_8570);
or U9212 (N_9212,N_8790,N_8863);
nor U9213 (N_9213,N_8975,N_8897);
or U9214 (N_9214,N_8677,N_8862);
or U9215 (N_9215,N_8839,N_8822);
nand U9216 (N_9216,N_8989,N_8642);
nor U9217 (N_9217,N_8571,N_8674);
and U9218 (N_9218,N_8580,N_8731);
nand U9219 (N_9219,N_8749,N_8815);
or U9220 (N_9220,N_8531,N_8768);
and U9221 (N_9221,N_8524,N_8864);
and U9222 (N_9222,N_8629,N_8507);
nand U9223 (N_9223,N_8654,N_8638);
and U9224 (N_9224,N_8651,N_8660);
nor U9225 (N_9225,N_8687,N_8914);
nand U9226 (N_9226,N_8627,N_8971);
and U9227 (N_9227,N_8607,N_8812);
nor U9228 (N_9228,N_8582,N_8809);
nor U9229 (N_9229,N_8866,N_8516);
xor U9230 (N_9230,N_8738,N_8618);
nor U9231 (N_9231,N_8684,N_8793);
nor U9232 (N_9232,N_8941,N_8965);
and U9233 (N_9233,N_8789,N_8886);
xor U9234 (N_9234,N_8623,N_8735);
and U9235 (N_9235,N_8669,N_8644);
nand U9236 (N_9236,N_8890,N_8799);
nand U9237 (N_9237,N_8908,N_8881);
or U9238 (N_9238,N_8518,N_8695);
and U9239 (N_9239,N_8598,N_8632);
nor U9240 (N_9240,N_8834,N_8800);
and U9241 (N_9241,N_8561,N_8519);
nor U9242 (N_9242,N_8959,N_8675);
nand U9243 (N_9243,N_8664,N_8947);
nor U9244 (N_9244,N_8769,N_8836);
and U9245 (N_9245,N_8734,N_8515);
nor U9246 (N_9246,N_8537,N_8853);
nand U9247 (N_9247,N_8889,N_8601);
and U9248 (N_9248,N_8847,N_8529);
or U9249 (N_9249,N_8962,N_8712);
nand U9250 (N_9250,N_8670,N_8657);
nor U9251 (N_9251,N_8542,N_8750);
nor U9252 (N_9252,N_8827,N_8608);
and U9253 (N_9253,N_8870,N_8962);
and U9254 (N_9254,N_8953,N_8766);
nand U9255 (N_9255,N_8627,N_8747);
or U9256 (N_9256,N_8801,N_8771);
or U9257 (N_9257,N_8607,N_8946);
and U9258 (N_9258,N_8988,N_8628);
xnor U9259 (N_9259,N_8623,N_8630);
nor U9260 (N_9260,N_8687,N_8822);
or U9261 (N_9261,N_8528,N_8803);
and U9262 (N_9262,N_8882,N_8677);
or U9263 (N_9263,N_8578,N_8555);
xnor U9264 (N_9264,N_8995,N_8575);
xor U9265 (N_9265,N_8865,N_8530);
nand U9266 (N_9266,N_8626,N_8922);
or U9267 (N_9267,N_8862,N_8944);
xnor U9268 (N_9268,N_8989,N_8966);
or U9269 (N_9269,N_8561,N_8820);
and U9270 (N_9270,N_8979,N_8947);
nand U9271 (N_9271,N_8573,N_8562);
nor U9272 (N_9272,N_8619,N_8546);
and U9273 (N_9273,N_8797,N_8710);
nand U9274 (N_9274,N_8684,N_8614);
xnor U9275 (N_9275,N_8892,N_8698);
nor U9276 (N_9276,N_8653,N_8581);
or U9277 (N_9277,N_8548,N_8731);
nor U9278 (N_9278,N_8931,N_8686);
or U9279 (N_9279,N_8945,N_8723);
and U9280 (N_9280,N_8562,N_8739);
or U9281 (N_9281,N_8544,N_8673);
or U9282 (N_9282,N_8965,N_8601);
xnor U9283 (N_9283,N_8564,N_8638);
nor U9284 (N_9284,N_8827,N_8575);
and U9285 (N_9285,N_8682,N_8704);
nand U9286 (N_9286,N_8877,N_8912);
nand U9287 (N_9287,N_8993,N_8722);
nor U9288 (N_9288,N_8813,N_8660);
nand U9289 (N_9289,N_8891,N_8655);
nor U9290 (N_9290,N_8561,N_8598);
nor U9291 (N_9291,N_8846,N_8855);
nand U9292 (N_9292,N_8565,N_8715);
or U9293 (N_9293,N_8776,N_8636);
and U9294 (N_9294,N_8741,N_8623);
nand U9295 (N_9295,N_8641,N_8607);
or U9296 (N_9296,N_8769,N_8945);
nand U9297 (N_9297,N_8730,N_8779);
nand U9298 (N_9298,N_8922,N_8678);
and U9299 (N_9299,N_8642,N_8772);
or U9300 (N_9300,N_8619,N_8577);
and U9301 (N_9301,N_8671,N_8632);
xor U9302 (N_9302,N_8639,N_8851);
nand U9303 (N_9303,N_8875,N_8585);
nor U9304 (N_9304,N_8956,N_8826);
or U9305 (N_9305,N_8558,N_8791);
nor U9306 (N_9306,N_8670,N_8669);
nand U9307 (N_9307,N_8525,N_8823);
or U9308 (N_9308,N_8601,N_8580);
nand U9309 (N_9309,N_8843,N_8647);
nand U9310 (N_9310,N_8688,N_8924);
nand U9311 (N_9311,N_8926,N_8533);
and U9312 (N_9312,N_8918,N_8966);
nor U9313 (N_9313,N_8695,N_8818);
and U9314 (N_9314,N_8995,N_8522);
nand U9315 (N_9315,N_8621,N_8710);
nor U9316 (N_9316,N_8797,N_8627);
xor U9317 (N_9317,N_8962,N_8703);
nand U9318 (N_9318,N_8721,N_8580);
nand U9319 (N_9319,N_8655,N_8546);
and U9320 (N_9320,N_8882,N_8702);
and U9321 (N_9321,N_8580,N_8997);
xor U9322 (N_9322,N_8851,N_8716);
and U9323 (N_9323,N_8573,N_8728);
and U9324 (N_9324,N_8964,N_8794);
nand U9325 (N_9325,N_8580,N_8578);
or U9326 (N_9326,N_8849,N_8896);
nand U9327 (N_9327,N_8737,N_8761);
and U9328 (N_9328,N_8912,N_8720);
xnor U9329 (N_9329,N_8541,N_8689);
nand U9330 (N_9330,N_8668,N_8764);
or U9331 (N_9331,N_8901,N_8580);
xor U9332 (N_9332,N_8506,N_8694);
nor U9333 (N_9333,N_8775,N_8807);
and U9334 (N_9334,N_8500,N_8771);
nand U9335 (N_9335,N_8749,N_8658);
nor U9336 (N_9336,N_8620,N_8737);
and U9337 (N_9337,N_8952,N_8579);
nand U9338 (N_9338,N_8579,N_8510);
nor U9339 (N_9339,N_8588,N_8766);
xor U9340 (N_9340,N_8707,N_8534);
nor U9341 (N_9341,N_8664,N_8598);
or U9342 (N_9342,N_8926,N_8668);
nand U9343 (N_9343,N_8783,N_8873);
nand U9344 (N_9344,N_8959,N_8706);
nor U9345 (N_9345,N_8848,N_8688);
and U9346 (N_9346,N_8828,N_8814);
xnor U9347 (N_9347,N_8616,N_8656);
nor U9348 (N_9348,N_8889,N_8906);
or U9349 (N_9349,N_8826,N_8592);
and U9350 (N_9350,N_8640,N_8556);
nor U9351 (N_9351,N_8781,N_8850);
or U9352 (N_9352,N_8843,N_8681);
and U9353 (N_9353,N_8839,N_8666);
xor U9354 (N_9354,N_8898,N_8776);
and U9355 (N_9355,N_8512,N_8938);
or U9356 (N_9356,N_8871,N_8537);
xnor U9357 (N_9357,N_8552,N_8652);
or U9358 (N_9358,N_8658,N_8876);
and U9359 (N_9359,N_8964,N_8770);
xnor U9360 (N_9360,N_8880,N_8776);
nor U9361 (N_9361,N_8680,N_8912);
nand U9362 (N_9362,N_8711,N_8944);
nor U9363 (N_9363,N_8849,N_8505);
or U9364 (N_9364,N_8844,N_8860);
nor U9365 (N_9365,N_8786,N_8724);
or U9366 (N_9366,N_8904,N_8773);
and U9367 (N_9367,N_8746,N_8593);
and U9368 (N_9368,N_8863,N_8819);
and U9369 (N_9369,N_8742,N_8533);
nor U9370 (N_9370,N_8837,N_8978);
or U9371 (N_9371,N_8752,N_8846);
xor U9372 (N_9372,N_8790,N_8826);
nor U9373 (N_9373,N_8913,N_8556);
nor U9374 (N_9374,N_8899,N_8828);
or U9375 (N_9375,N_8532,N_8581);
xor U9376 (N_9376,N_8854,N_8826);
nor U9377 (N_9377,N_8893,N_8548);
nor U9378 (N_9378,N_8590,N_8727);
or U9379 (N_9379,N_8938,N_8957);
nand U9380 (N_9380,N_8657,N_8573);
nor U9381 (N_9381,N_8638,N_8925);
and U9382 (N_9382,N_8963,N_8971);
and U9383 (N_9383,N_8755,N_8634);
or U9384 (N_9384,N_8517,N_8522);
xor U9385 (N_9385,N_8510,N_8722);
nand U9386 (N_9386,N_8744,N_8602);
nand U9387 (N_9387,N_8684,N_8901);
nand U9388 (N_9388,N_8743,N_8997);
or U9389 (N_9389,N_8793,N_8783);
nor U9390 (N_9390,N_8713,N_8799);
nand U9391 (N_9391,N_8574,N_8533);
and U9392 (N_9392,N_8599,N_8784);
nand U9393 (N_9393,N_8815,N_8637);
nand U9394 (N_9394,N_8932,N_8815);
or U9395 (N_9395,N_8514,N_8919);
nand U9396 (N_9396,N_8837,N_8839);
or U9397 (N_9397,N_8500,N_8572);
and U9398 (N_9398,N_8516,N_8771);
and U9399 (N_9399,N_8924,N_8737);
nand U9400 (N_9400,N_8771,N_8533);
nor U9401 (N_9401,N_8687,N_8768);
xnor U9402 (N_9402,N_8772,N_8995);
nor U9403 (N_9403,N_8522,N_8742);
nor U9404 (N_9404,N_8937,N_8566);
nand U9405 (N_9405,N_8545,N_8770);
or U9406 (N_9406,N_8559,N_8900);
and U9407 (N_9407,N_8974,N_8550);
or U9408 (N_9408,N_8657,N_8568);
or U9409 (N_9409,N_8969,N_8689);
and U9410 (N_9410,N_8666,N_8926);
nor U9411 (N_9411,N_8585,N_8720);
nand U9412 (N_9412,N_8618,N_8558);
or U9413 (N_9413,N_8946,N_8717);
nor U9414 (N_9414,N_8885,N_8528);
and U9415 (N_9415,N_8887,N_8700);
nor U9416 (N_9416,N_8824,N_8838);
nand U9417 (N_9417,N_8842,N_8931);
nor U9418 (N_9418,N_8779,N_8743);
nand U9419 (N_9419,N_8711,N_8920);
or U9420 (N_9420,N_8687,N_8817);
or U9421 (N_9421,N_8727,N_8692);
xor U9422 (N_9422,N_8510,N_8765);
or U9423 (N_9423,N_8559,N_8983);
nand U9424 (N_9424,N_8663,N_8753);
or U9425 (N_9425,N_8584,N_8875);
and U9426 (N_9426,N_8929,N_8888);
or U9427 (N_9427,N_8920,N_8826);
or U9428 (N_9428,N_8879,N_8829);
or U9429 (N_9429,N_8759,N_8920);
or U9430 (N_9430,N_8572,N_8970);
nor U9431 (N_9431,N_8814,N_8804);
nand U9432 (N_9432,N_8503,N_8714);
xnor U9433 (N_9433,N_8584,N_8576);
nand U9434 (N_9434,N_8515,N_8699);
nor U9435 (N_9435,N_8845,N_8821);
and U9436 (N_9436,N_8789,N_8509);
or U9437 (N_9437,N_8857,N_8715);
or U9438 (N_9438,N_8701,N_8745);
nor U9439 (N_9439,N_8800,N_8615);
and U9440 (N_9440,N_8856,N_8764);
and U9441 (N_9441,N_8598,N_8631);
and U9442 (N_9442,N_8820,N_8892);
and U9443 (N_9443,N_8865,N_8873);
and U9444 (N_9444,N_8651,N_8585);
and U9445 (N_9445,N_8908,N_8853);
and U9446 (N_9446,N_8900,N_8830);
nor U9447 (N_9447,N_8700,N_8869);
nand U9448 (N_9448,N_8634,N_8908);
or U9449 (N_9449,N_8577,N_8943);
and U9450 (N_9450,N_8866,N_8993);
nor U9451 (N_9451,N_8792,N_8553);
nor U9452 (N_9452,N_8654,N_8725);
or U9453 (N_9453,N_8552,N_8594);
nand U9454 (N_9454,N_8770,N_8604);
nand U9455 (N_9455,N_8956,N_8824);
nand U9456 (N_9456,N_8512,N_8818);
and U9457 (N_9457,N_8637,N_8579);
or U9458 (N_9458,N_8678,N_8542);
or U9459 (N_9459,N_8989,N_8521);
nor U9460 (N_9460,N_8762,N_8885);
nor U9461 (N_9461,N_8673,N_8777);
nand U9462 (N_9462,N_8655,N_8511);
and U9463 (N_9463,N_8605,N_8928);
nand U9464 (N_9464,N_8921,N_8775);
and U9465 (N_9465,N_8722,N_8547);
or U9466 (N_9466,N_8819,N_8583);
xor U9467 (N_9467,N_8788,N_8686);
or U9468 (N_9468,N_8994,N_8898);
nand U9469 (N_9469,N_8602,N_8830);
and U9470 (N_9470,N_8848,N_8973);
and U9471 (N_9471,N_8604,N_8584);
or U9472 (N_9472,N_8658,N_8754);
nand U9473 (N_9473,N_8736,N_8509);
and U9474 (N_9474,N_8730,N_8781);
nand U9475 (N_9475,N_8682,N_8620);
xor U9476 (N_9476,N_8989,N_8777);
nor U9477 (N_9477,N_8940,N_8698);
nand U9478 (N_9478,N_8738,N_8570);
nor U9479 (N_9479,N_8568,N_8996);
nand U9480 (N_9480,N_8560,N_8631);
and U9481 (N_9481,N_8783,N_8523);
and U9482 (N_9482,N_8767,N_8928);
nand U9483 (N_9483,N_8523,N_8909);
nor U9484 (N_9484,N_8819,N_8750);
and U9485 (N_9485,N_8611,N_8711);
nor U9486 (N_9486,N_8728,N_8871);
or U9487 (N_9487,N_8739,N_8668);
nand U9488 (N_9488,N_8945,N_8659);
nand U9489 (N_9489,N_8552,N_8784);
nand U9490 (N_9490,N_8698,N_8922);
or U9491 (N_9491,N_8722,N_8961);
or U9492 (N_9492,N_8967,N_8646);
xor U9493 (N_9493,N_8500,N_8792);
nor U9494 (N_9494,N_8535,N_8984);
nor U9495 (N_9495,N_8777,N_8812);
and U9496 (N_9496,N_8703,N_8852);
nand U9497 (N_9497,N_8599,N_8929);
xor U9498 (N_9498,N_8767,N_8695);
nand U9499 (N_9499,N_8896,N_8599);
and U9500 (N_9500,N_9373,N_9212);
nor U9501 (N_9501,N_9497,N_9017);
or U9502 (N_9502,N_9467,N_9463);
nand U9503 (N_9503,N_9058,N_9132);
nor U9504 (N_9504,N_9073,N_9036);
and U9505 (N_9505,N_9136,N_9133);
nand U9506 (N_9506,N_9245,N_9433);
nand U9507 (N_9507,N_9458,N_9040);
or U9508 (N_9508,N_9317,N_9189);
nor U9509 (N_9509,N_9233,N_9422);
nand U9510 (N_9510,N_9261,N_9236);
or U9511 (N_9511,N_9401,N_9063);
and U9512 (N_9512,N_9171,N_9099);
nor U9513 (N_9513,N_9353,N_9417);
or U9514 (N_9514,N_9342,N_9115);
or U9515 (N_9515,N_9399,N_9195);
and U9516 (N_9516,N_9213,N_9468);
nand U9517 (N_9517,N_9310,N_9411);
nor U9518 (N_9518,N_9314,N_9348);
or U9519 (N_9519,N_9101,N_9203);
or U9520 (N_9520,N_9174,N_9252);
or U9521 (N_9521,N_9210,N_9100);
or U9522 (N_9522,N_9004,N_9486);
or U9523 (N_9523,N_9404,N_9387);
nand U9524 (N_9524,N_9379,N_9326);
or U9525 (N_9525,N_9278,N_9328);
and U9526 (N_9526,N_9388,N_9194);
nor U9527 (N_9527,N_9435,N_9138);
nor U9528 (N_9528,N_9472,N_9331);
nor U9529 (N_9529,N_9364,N_9475);
or U9530 (N_9530,N_9227,N_9391);
nand U9531 (N_9531,N_9144,N_9121);
nand U9532 (N_9532,N_9418,N_9449);
nor U9533 (N_9533,N_9325,N_9114);
or U9534 (N_9534,N_9222,N_9102);
nand U9535 (N_9535,N_9498,N_9157);
nor U9536 (N_9536,N_9406,N_9207);
nand U9537 (N_9537,N_9359,N_9262);
xnor U9538 (N_9538,N_9151,N_9442);
and U9539 (N_9539,N_9384,N_9251);
nand U9540 (N_9540,N_9035,N_9260);
or U9541 (N_9541,N_9088,N_9180);
nor U9542 (N_9542,N_9492,N_9028);
and U9543 (N_9543,N_9312,N_9053);
or U9544 (N_9544,N_9027,N_9340);
nand U9545 (N_9545,N_9407,N_9060);
or U9546 (N_9546,N_9270,N_9175);
nor U9547 (N_9547,N_9170,N_9003);
and U9548 (N_9548,N_9276,N_9007);
or U9549 (N_9549,N_9488,N_9134);
or U9550 (N_9550,N_9295,N_9358);
nor U9551 (N_9551,N_9034,N_9182);
nor U9552 (N_9552,N_9098,N_9108);
and U9553 (N_9553,N_9414,N_9072);
and U9554 (N_9554,N_9343,N_9464);
xor U9555 (N_9555,N_9452,N_9224);
or U9556 (N_9556,N_9499,N_9025);
and U9557 (N_9557,N_9131,N_9321);
nand U9558 (N_9558,N_9455,N_9327);
and U9559 (N_9559,N_9392,N_9226);
xnor U9560 (N_9560,N_9347,N_9275);
and U9561 (N_9561,N_9011,N_9309);
xor U9562 (N_9562,N_9029,N_9288);
xnor U9563 (N_9563,N_9427,N_9232);
or U9564 (N_9564,N_9292,N_9263);
or U9565 (N_9565,N_9443,N_9070);
and U9566 (N_9566,N_9061,N_9380);
xor U9567 (N_9567,N_9393,N_9265);
nand U9568 (N_9568,N_9448,N_9366);
and U9569 (N_9569,N_9487,N_9298);
nand U9570 (N_9570,N_9282,N_9211);
nand U9571 (N_9571,N_9377,N_9436);
and U9572 (N_9572,N_9480,N_9336);
and U9573 (N_9573,N_9112,N_9163);
xor U9574 (N_9574,N_9409,N_9390);
or U9575 (N_9575,N_9402,N_9009);
nor U9576 (N_9576,N_9272,N_9239);
and U9577 (N_9577,N_9301,N_9269);
xor U9578 (N_9578,N_9065,N_9357);
nand U9579 (N_9579,N_9005,N_9281);
nor U9580 (N_9580,N_9396,N_9051);
or U9581 (N_9581,N_9344,N_9014);
nor U9582 (N_9582,N_9473,N_9001);
or U9583 (N_9583,N_9451,N_9042);
and U9584 (N_9584,N_9367,N_9441);
nand U9585 (N_9585,N_9454,N_9188);
nand U9586 (N_9586,N_9316,N_9139);
nor U9587 (N_9587,N_9221,N_9395);
nand U9588 (N_9588,N_9071,N_9218);
nor U9589 (N_9589,N_9156,N_9438);
nor U9590 (N_9590,N_9320,N_9045);
nor U9591 (N_9591,N_9285,N_9111);
or U9592 (N_9592,N_9496,N_9032);
xor U9593 (N_9593,N_9471,N_9067);
xnor U9594 (N_9594,N_9081,N_9122);
nand U9595 (N_9595,N_9319,N_9062);
or U9596 (N_9596,N_9076,N_9290);
nand U9597 (N_9597,N_9318,N_9026);
xor U9598 (N_9598,N_9082,N_9123);
nand U9599 (N_9599,N_9225,N_9006);
nand U9600 (N_9600,N_9000,N_9378);
or U9601 (N_9601,N_9337,N_9477);
xor U9602 (N_9602,N_9079,N_9056);
or U9603 (N_9603,N_9087,N_9172);
or U9604 (N_9604,N_9179,N_9434);
and U9605 (N_9605,N_9117,N_9440);
and U9606 (N_9606,N_9015,N_9482);
or U9607 (N_9607,N_9185,N_9255);
or U9608 (N_9608,N_9246,N_9362);
or U9609 (N_9609,N_9462,N_9299);
nor U9610 (N_9610,N_9089,N_9303);
or U9611 (N_9611,N_9426,N_9141);
xor U9612 (N_9612,N_9247,N_9178);
nor U9613 (N_9613,N_9242,N_9368);
nand U9614 (N_9614,N_9116,N_9238);
nor U9615 (N_9615,N_9177,N_9375);
nand U9616 (N_9616,N_9168,N_9086);
xor U9617 (N_9617,N_9453,N_9104);
and U9618 (N_9618,N_9140,N_9080);
or U9619 (N_9619,N_9078,N_9191);
nor U9620 (N_9620,N_9147,N_9351);
and U9621 (N_9621,N_9478,N_9074);
and U9622 (N_9622,N_9383,N_9250);
nand U9623 (N_9623,N_9201,N_9332);
xnor U9624 (N_9624,N_9110,N_9193);
and U9625 (N_9625,N_9052,N_9165);
or U9626 (N_9626,N_9095,N_9125);
or U9627 (N_9627,N_9456,N_9302);
or U9628 (N_9628,N_9444,N_9322);
and U9629 (N_9629,N_9154,N_9491);
or U9630 (N_9630,N_9159,N_9012);
and U9631 (N_9631,N_9381,N_9127);
nand U9632 (N_9632,N_9217,N_9135);
or U9633 (N_9633,N_9046,N_9445);
and U9634 (N_9634,N_9044,N_9047);
and U9635 (N_9635,N_9184,N_9304);
and U9636 (N_9636,N_9169,N_9020);
nor U9637 (N_9637,N_9408,N_9405);
nor U9638 (N_9638,N_9173,N_9306);
nor U9639 (N_9639,N_9024,N_9216);
nor U9640 (N_9640,N_9258,N_9231);
nor U9641 (N_9641,N_9372,N_9280);
or U9642 (N_9642,N_9335,N_9385);
xor U9643 (N_9643,N_9106,N_9197);
or U9644 (N_9644,N_9018,N_9037);
or U9645 (N_9645,N_9267,N_9370);
and U9646 (N_9646,N_9397,N_9196);
nor U9647 (N_9647,N_9164,N_9248);
nand U9648 (N_9648,N_9214,N_9235);
and U9649 (N_9649,N_9243,N_9068);
or U9650 (N_9650,N_9489,N_9493);
xnor U9651 (N_9651,N_9143,N_9043);
nand U9652 (N_9652,N_9093,N_9479);
and U9653 (N_9653,N_9481,N_9162);
nor U9654 (N_9654,N_9066,N_9023);
nand U9655 (N_9655,N_9202,N_9289);
nor U9656 (N_9656,N_9160,N_9031);
nor U9657 (N_9657,N_9389,N_9187);
and U9658 (N_9658,N_9206,N_9176);
xnor U9659 (N_9659,N_9307,N_9096);
or U9660 (N_9660,N_9277,N_9155);
and U9661 (N_9661,N_9181,N_9167);
nand U9662 (N_9662,N_9274,N_9150);
nand U9663 (N_9663,N_9077,N_9356);
nand U9664 (N_9664,N_9446,N_9240);
nor U9665 (N_9665,N_9016,N_9410);
nand U9666 (N_9666,N_9257,N_9146);
nand U9667 (N_9667,N_9183,N_9416);
or U9668 (N_9668,N_9474,N_9279);
or U9669 (N_9669,N_9429,N_9228);
nor U9670 (N_9670,N_9350,N_9190);
and U9671 (N_9671,N_9339,N_9334);
xor U9672 (N_9672,N_9439,N_9120);
and U9673 (N_9673,N_9254,N_9363);
xor U9674 (N_9674,N_9145,N_9186);
and U9675 (N_9675,N_9158,N_9329);
or U9676 (N_9676,N_9039,N_9296);
or U9677 (N_9677,N_9403,N_9346);
and U9678 (N_9678,N_9431,N_9371);
nand U9679 (N_9679,N_9119,N_9054);
nor U9680 (N_9680,N_9354,N_9333);
or U9681 (N_9681,N_9420,N_9369);
or U9682 (N_9682,N_9097,N_9421);
nand U9683 (N_9683,N_9118,N_9415);
nand U9684 (N_9684,N_9294,N_9215);
nand U9685 (N_9685,N_9022,N_9094);
and U9686 (N_9686,N_9485,N_9008);
nor U9687 (N_9687,N_9283,N_9223);
nand U9688 (N_9688,N_9365,N_9041);
or U9689 (N_9689,N_9229,N_9209);
nor U9690 (N_9690,N_9019,N_9220);
and U9691 (N_9691,N_9048,N_9413);
nand U9692 (N_9692,N_9130,N_9128);
nand U9693 (N_9693,N_9386,N_9241);
xnor U9694 (N_9694,N_9447,N_9484);
and U9695 (N_9695,N_9148,N_9311);
xor U9696 (N_9696,N_9152,N_9419);
or U9697 (N_9697,N_9266,N_9244);
xor U9698 (N_9698,N_9166,N_9021);
or U9699 (N_9699,N_9374,N_9126);
nand U9700 (N_9700,N_9466,N_9460);
or U9701 (N_9701,N_9412,N_9149);
or U9702 (N_9702,N_9400,N_9208);
and U9703 (N_9703,N_9330,N_9033);
and U9704 (N_9704,N_9355,N_9253);
nand U9705 (N_9705,N_9382,N_9059);
or U9706 (N_9706,N_9469,N_9083);
nor U9707 (N_9707,N_9341,N_9450);
and U9708 (N_9708,N_9425,N_9234);
and U9709 (N_9709,N_9271,N_9476);
nand U9710 (N_9710,N_9230,N_9204);
and U9711 (N_9711,N_9075,N_9105);
nor U9712 (N_9712,N_9069,N_9494);
nand U9713 (N_9713,N_9084,N_9124);
and U9714 (N_9714,N_9259,N_9085);
nand U9715 (N_9715,N_9313,N_9428);
nand U9716 (N_9716,N_9268,N_9324);
or U9717 (N_9717,N_9291,N_9465);
and U9718 (N_9718,N_9113,N_9237);
nor U9719 (N_9719,N_9490,N_9064);
nand U9720 (N_9720,N_9256,N_9055);
nand U9721 (N_9721,N_9129,N_9091);
and U9722 (N_9722,N_9049,N_9424);
xor U9723 (N_9723,N_9345,N_9109);
nor U9724 (N_9724,N_9360,N_9361);
nand U9725 (N_9725,N_9092,N_9090);
nor U9726 (N_9726,N_9457,N_9293);
and U9727 (N_9727,N_9432,N_9137);
or U9728 (N_9728,N_9198,N_9142);
nand U9729 (N_9729,N_9192,N_9349);
nor U9730 (N_9730,N_9323,N_9013);
nor U9731 (N_9731,N_9297,N_9423);
nand U9732 (N_9732,N_9002,N_9483);
nand U9733 (N_9733,N_9103,N_9249);
nand U9734 (N_9734,N_9376,N_9430);
or U9735 (N_9735,N_9050,N_9219);
and U9736 (N_9736,N_9264,N_9352);
or U9737 (N_9737,N_9305,N_9161);
or U9738 (N_9738,N_9205,N_9287);
nand U9739 (N_9739,N_9338,N_9461);
nor U9740 (N_9740,N_9286,N_9107);
or U9741 (N_9741,N_9010,N_9284);
xnor U9742 (N_9742,N_9200,N_9057);
and U9743 (N_9743,N_9199,N_9038);
and U9744 (N_9744,N_9437,N_9273);
nor U9745 (N_9745,N_9153,N_9398);
nor U9746 (N_9746,N_9459,N_9030);
and U9747 (N_9747,N_9394,N_9300);
and U9748 (N_9748,N_9315,N_9495);
nor U9749 (N_9749,N_9308,N_9470);
nand U9750 (N_9750,N_9403,N_9492);
or U9751 (N_9751,N_9084,N_9432);
or U9752 (N_9752,N_9072,N_9051);
or U9753 (N_9753,N_9362,N_9132);
nand U9754 (N_9754,N_9203,N_9302);
xnor U9755 (N_9755,N_9145,N_9048);
and U9756 (N_9756,N_9289,N_9274);
or U9757 (N_9757,N_9088,N_9135);
or U9758 (N_9758,N_9215,N_9155);
or U9759 (N_9759,N_9128,N_9272);
xor U9760 (N_9760,N_9442,N_9160);
nand U9761 (N_9761,N_9252,N_9214);
xnor U9762 (N_9762,N_9436,N_9096);
nand U9763 (N_9763,N_9171,N_9357);
and U9764 (N_9764,N_9228,N_9065);
and U9765 (N_9765,N_9073,N_9442);
and U9766 (N_9766,N_9371,N_9275);
nor U9767 (N_9767,N_9119,N_9152);
nor U9768 (N_9768,N_9297,N_9162);
or U9769 (N_9769,N_9121,N_9390);
nor U9770 (N_9770,N_9363,N_9168);
and U9771 (N_9771,N_9430,N_9011);
nor U9772 (N_9772,N_9246,N_9176);
nand U9773 (N_9773,N_9097,N_9343);
nand U9774 (N_9774,N_9464,N_9365);
nor U9775 (N_9775,N_9102,N_9231);
and U9776 (N_9776,N_9045,N_9454);
nand U9777 (N_9777,N_9087,N_9050);
and U9778 (N_9778,N_9158,N_9167);
and U9779 (N_9779,N_9314,N_9447);
nor U9780 (N_9780,N_9222,N_9305);
nand U9781 (N_9781,N_9106,N_9026);
nand U9782 (N_9782,N_9204,N_9207);
and U9783 (N_9783,N_9110,N_9085);
nand U9784 (N_9784,N_9364,N_9384);
xor U9785 (N_9785,N_9318,N_9419);
nand U9786 (N_9786,N_9029,N_9061);
nand U9787 (N_9787,N_9284,N_9491);
and U9788 (N_9788,N_9012,N_9188);
xnor U9789 (N_9789,N_9172,N_9492);
nand U9790 (N_9790,N_9463,N_9480);
and U9791 (N_9791,N_9247,N_9499);
and U9792 (N_9792,N_9411,N_9171);
or U9793 (N_9793,N_9359,N_9349);
or U9794 (N_9794,N_9123,N_9129);
nor U9795 (N_9795,N_9159,N_9037);
and U9796 (N_9796,N_9071,N_9346);
nand U9797 (N_9797,N_9036,N_9309);
nor U9798 (N_9798,N_9291,N_9308);
or U9799 (N_9799,N_9364,N_9315);
nor U9800 (N_9800,N_9125,N_9177);
or U9801 (N_9801,N_9010,N_9329);
nand U9802 (N_9802,N_9390,N_9204);
and U9803 (N_9803,N_9003,N_9312);
or U9804 (N_9804,N_9482,N_9293);
or U9805 (N_9805,N_9487,N_9046);
xnor U9806 (N_9806,N_9222,N_9185);
nor U9807 (N_9807,N_9415,N_9064);
or U9808 (N_9808,N_9018,N_9446);
nor U9809 (N_9809,N_9295,N_9406);
or U9810 (N_9810,N_9227,N_9306);
nand U9811 (N_9811,N_9442,N_9121);
nand U9812 (N_9812,N_9036,N_9497);
and U9813 (N_9813,N_9482,N_9019);
or U9814 (N_9814,N_9171,N_9282);
nor U9815 (N_9815,N_9397,N_9357);
nor U9816 (N_9816,N_9091,N_9386);
or U9817 (N_9817,N_9284,N_9366);
or U9818 (N_9818,N_9351,N_9170);
nor U9819 (N_9819,N_9242,N_9162);
or U9820 (N_9820,N_9150,N_9334);
and U9821 (N_9821,N_9059,N_9295);
and U9822 (N_9822,N_9034,N_9033);
or U9823 (N_9823,N_9272,N_9490);
nand U9824 (N_9824,N_9418,N_9325);
nand U9825 (N_9825,N_9129,N_9484);
and U9826 (N_9826,N_9472,N_9264);
nand U9827 (N_9827,N_9153,N_9373);
nor U9828 (N_9828,N_9134,N_9374);
and U9829 (N_9829,N_9100,N_9420);
and U9830 (N_9830,N_9235,N_9229);
or U9831 (N_9831,N_9091,N_9351);
nand U9832 (N_9832,N_9465,N_9284);
or U9833 (N_9833,N_9116,N_9287);
nand U9834 (N_9834,N_9427,N_9302);
and U9835 (N_9835,N_9094,N_9126);
xor U9836 (N_9836,N_9206,N_9326);
and U9837 (N_9837,N_9204,N_9238);
and U9838 (N_9838,N_9300,N_9128);
or U9839 (N_9839,N_9262,N_9291);
nor U9840 (N_9840,N_9330,N_9421);
or U9841 (N_9841,N_9074,N_9239);
and U9842 (N_9842,N_9155,N_9351);
and U9843 (N_9843,N_9162,N_9416);
nor U9844 (N_9844,N_9075,N_9291);
nand U9845 (N_9845,N_9339,N_9220);
nor U9846 (N_9846,N_9449,N_9402);
or U9847 (N_9847,N_9327,N_9106);
nand U9848 (N_9848,N_9191,N_9439);
nor U9849 (N_9849,N_9251,N_9225);
nand U9850 (N_9850,N_9477,N_9083);
nand U9851 (N_9851,N_9368,N_9479);
nor U9852 (N_9852,N_9196,N_9127);
and U9853 (N_9853,N_9238,N_9434);
nand U9854 (N_9854,N_9192,N_9128);
or U9855 (N_9855,N_9390,N_9084);
and U9856 (N_9856,N_9149,N_9098);
or U9857 (N_9857,N_9127,N_9185);
or U9858 (N_9858,N_9359,N_9470);
or U9859 (N_9859,N_9236,N_9181);
and U9860 (N_9860,N_9453,N_9280);
xnor U9861 (N_9861,N_9110,N_9209);
xnor U9862 (N_9862,N_9135,N_9318);
nand U9863 (N_9863,N_9266,N_9182);
nor U9864 (N_9864,N_9364,N_9293);
nand U9865 (N_9865,N_9194,N_9079);
or U9866 (N_9866,N_9007,N_9494);
nand U9867 (N_9867,N_9189,N_9258);
nand U9868 (N_9868,N_9484,N_9205);
nor U9869 (N_9869,N_9030,N_9425);
or U9870 (N_9870,N_9177,N_9462);
nor U9871 (N_9871,N_9279,N_9213);
nor U9872 (N_9872,N_9364,N_9180);
or U9873 (N_9873,N_9364,N_9032);
or U9874 (N_9874,N_9233,N_9062);
nand U9875 (N_9875,N_9418,N_9116);
and U9876 (N_9876,N_9435,N_9373);
and U9877 (N_9877,N_9479,N_9467);
or U9878 (N_9878,N_9280,N_9351);
or U9879 (N_9879,N_9327,N_9025);
nand U9880 (N_9880,N_9008,N_9208);
and U9881 (N_9881,N_9168,N_9414);
or U9882 (N_9882,N_9313,N_9381);
and U9883 (N_9883,N_9113,N_9247);
or U9884 (N_9884,N_9440,N_9482);
and U9885 (N_9885,N_9170,N_9392);
nand U9886 (N_9886,N_9472,N_9037);
or U9887 (N_9887,N_9180,N_9397);
nand U9888 (N_9888,N_9157,N_9237);
and U9889 (N_9889,N_9270,N_9029);
and U9890 (N_9890,N_9385,N_9059);
nor U9891 (N_9891,N_9084,N_9322);
or U9892 (N_9892,N_9067,N_9141);
nor U9893 (N_9893,N_9276,N_9189);
and U9894 (N_9894,N_9002,N_9448);
nor U9895 (N_9895,N_9390,N_9040);
and U9896 (N_9896,N_9019,N_9433);
and U9897 (N_9897,N_9197,N_9292);
nor U9898 (N_9898,N_9127,N_9288);
and U9899 (N_9899,N_9258,N_9271);
and U9900 (N_9900,N_9042,N_9012);
nor U9901 (N_9901,N_9199,N_9074);
xnor U9902 (N_9902,N_9377,N_9395);
nor U9903 (N_9903,N_9124,N_9199);
nand U9904 (N_9904,N_9069,N_9005);
and U9905 (N_9905,N_9259,N_9454);
and U9906 (N_9906,N_9105,N_9387);
or U9907 (N_9907,N_9097,N_9275);
nand U9908 (N_9908,N_9045,N_9408);
nor U9909 (N_9909,N_9105,N_9067);
or U9910 (N_9910,N_9313,N_9470);
and U9911 (N_9911,N_9387,N_9274);
nand U9912 (N_9912,N_9334,N_9390);
or U9913 (N_9913,N_9060,N_9202);
xor U9914 (N_9914,N_9008,N_9454);
nand U9915 (N_9915,N_9400,N_9301);
nand U9916 (N_9916,N_9320,N_9293);
and U9917 (N_9917,N_9436,N_9094);
nand U9918 (N_9918,N_9359,N_9274);
and U9919 (N_9919,N_9046,N_9012);
and U9920 (N_9920,N_9359,N_9085);
nand U9921 (N_9921,N_9378,N_9234);
nand U9922 (N_9922,N_9233,N_9147);
nor U9923 (N_9923,N_9453,N_9388);
nand U9924 (N_9924,N_9416,N_9121);
and U9925 (N_9925,N_9339,N_9479);
or U9926 (N_9926,N_9383,N_9440);
or U9927 (N_9927,N_9430,N_9238);
and U9928 (N_9928,N_9192,N_9237);
or U9929 (N_9929,N_9452,N_9133);
nand U9930 (N_9930,N_9273,N_9487);
or U9931 (N_9931,N_9083,N_9012);
and U9932 (N_9932,N_9107,N_9089);
nand U9933 (N_9933,N_9178,N_9006);
and U9934 (N_9934,N_9299,N_9219);
or U9935 (N_9935,N_9003,N_9167);
and U9936 (N_9936,N_9150,N_9099);
or U9937 (N_9937,N_9226,N_9228);
nand U9938 (N_9938,N_9180,N_9120);
nand U9939 (N_9939,N_9415,N_9445);
or U9940 (N_9940,N_9008,N_9020);
or U9941 (N_9941,N_9150,N_9384);
nor U9942 (N_9942,N_9318,N_9027);
or U9943 (N_9943,N_9012,N_9240);
nand U9944 (N_9944,N_9008,N_9024);
and U9945 (N_9945,N_9054,N_9270);
or U9946 (N_9946,N_9315,N_9415);
nor U9947 (N_9947,N_9380,N_9174);
xnor U9948 (N_9948,N_9081,N_9484);
xor U9949 (N_9949,N_9369,N_9478);
or U9950 (N_9950,N_9081,N_9171);
nand U9951 (N_9951,N_9399,N_9194);
or U9952 (N_9952,N_9204,N_9313);
nor U9953 (N_9953,N_9186,N_9343);
or U9954 (N_9954,N_9087,N_9481);
nand U9955 (N_9955,N_9199,N_9072);
and U9956 (N_9956,N_9166,N_9485);
and U9957 (N_9957,N_9163,N_9290);
or U9958 (N_9958,N_9111,N_9146);
or U9959 (N_9959,N_9307,N_9301);
and U9960 (N_9960,N_9004,N_9305);
nand U9961 (N_9961,N_9213,N_9048);
nand U9962 (N_9962,N_9408,N_9320);
nand U9963 (N_9963,N_9464,N_9229);
nor U9964 (N_9964,N_9061,N_9295);
or U9965 (N_9965,N_9413,N_9455);
nor U9966 (N_9966,N_9204,N_9335);
or U9967 (N_9967,N_9386,N_9005);
and U9968 (N_9968,N_9340,N_9478);
nand U9969 (N_9969,N_9191,N_9177);
and U9970 (N_9970,N_9314,N_9229);
or U9971 (N_9971,N_9350,N_9482);
or U9972 (N_9972,N_9220,N_9323);
xor U9973 (N_9973,N_9095,N_9022);
or U9974 (N_9974,N_9080,N_9404);
nand U9975 (N_9975,N_9442,N_9499);
nor U9976 (N_9976,N_9293,N_9099);
nand U9977 (N_9977,N_9325,N_9244);
nor U9978 (N_9978,N_9242,N_9311);
nand U9979 (N_9979,N_9414,N_9015);
nor U9980 (N_9980,N_9376,N_9455);
or U9981 (N_9981,N_9076,N_9352);
xor U9982 (N_9982,N_9257,N_9315);
nand U9983 (N_9983,N_9266,N_9144);
nor U9984 (N_9984,N_9006,N_9101);
nand U9985 (N_9985,N_9096,N_9248);
nand U9986 (N_9986,N_9110,N_9010);
nand U9987 (N_9987,N_9471,N_9202);
and U9988 (N_9988,N_9321,N_9389);
nand U9989 (N_9989,N_9368,N_9334);
xnor U9990 (N_9990,N_9046,N_9058);
nor U9991 (N_9991,N_9379,N_9072);
and U9992 (N_9992,N_9084,N_9118);
and U9993 (N_9993,N_9335,N_9491);
xor U9994 (N_9994,N_9065,N_9020);
nor U9995 (N_9995,N_9176,N_9490);
or U9996 (N_9996,N_9006,N_9338);
and U9997 (N_9997,N_9072,N_9389);
nor U9998 (N_9998,N_9201,N_9124);
nand U9999 (N_9999,N_9457,N_9424);
nand U10000 (N_10000,N_9700,N_9697);
xnor U10001 (N_10001,N_9531,N_9525);
nand U10002 (N_10002,N_9970,N_9862);
or U10003 (N_10003,N_9930,N_9562);
nor U10004 (N_10004,N_9567,N_9580);
nor U10005 (N_10005,N_9711,N_9628);
nand U10006 (N_10006,N_9641,N_9516);
and U10007 (N_10007,N_9633,N_9514);
nand U10008 (N_10008,N_9672,N_9627);
or U10009 (N_10009,N_9594,N_9617);
nor U10010 (N_10010,N_9956,N_9554);
nand U10011 (N_10011,N_9847,N_9784);
nand U10012 (N_10012,N_9529,N_9863);
and U10013 (N_10013,N_9704,N_9714);
xor U10014 (N_10014,N_9873,N_9926);
or U10015 (N_10015,N_9935,N_9741);
or U10016 (N_10016,N_9619,N_9947);
nor U10017 (N_10017,N_9588,N_9522);
or U10018 (N_10018,N_9515,N_9945);
nand U10019 (N_10019,N_9671,N_9615);
xor U10020 (N_10020,N_9864,N_9960);
xnor U10021 (N_10021,N_9557,N_9844);
xnor U10022 (N_10022,N_9751,N_9528);
nand U10023 (N_10023,N_9600,N_9511);
and U10024 (N_10024,N_9551,N_9954);
nor U10025 (N_10025,N_9545,N_9882);
or U10026 (N_10026,N_9646,N_9716);
nor U10027 (N_10027,N_9823,N_9771);
and U10028 (N_10028,N_9684,N_9686);
xor U10029 (N_10029,N_9717,N_9931);
and U10030 (N_10030,N_9653,N_9650);
and U10031 (N_10031,N_9609,N_9502);
and U10032 (N_10032,N_9505,N_9821);
or U10033 (N_10033,N_9851,N_9572);
nor U10034 (N_10034,N_9907,N_9829);
nand U10035 (N_10035,N_9875,N_9585);
or U10036 (N_10036,N_9856,N_9839);
or U10037 (N_10037,N_9889,N_9659);
and U10038 (N_10038,N_9701,N_9749);
or U10039 (N_10039,N_9901,N_9988);
or U10040 (N_10040,N_9649,N_9836);
xor U10041 (N_10041,N_9637,N_9781);
or U10042 (N_10042,N_9950,N_9920);
and U10043 (N_10043,N_9718,N_9855);
or U10044 (N_10044,N_9974,N_9869);
and U10045 (N_10045,N_9799,N_9852);
or U10046 (N_10046,N_9730,N_9946);
nand U10047 (N_10047,N_9849,N_9807);
or U10048 (N_10048,N_9803,N_9993);
or U10049 (N_10049,N_9508,N_9890);
nor U10050 (N_10050,N_9512,N_9876);
and U10051 (N_10051,N_9984,N_9573);
or U10052 (N_10052,N_9929,N_9962);
or U10053 (N_10053,N_9584,N_9549);
nor U10054 (N_10054,N_9846,N_9842);
nor U10055 (N_10055,N_9828,N_9967);
or U10056 (N_10056,N_9552,N_9743);
nand U10057 (N_10057,N_9568,N_9958);
or U10058 (N_10058,N_9555,N_9520);
or U10059 (N_10059,N_9533,N_9558);
and U10060 (N_10060,N_9689,N_9918);
nor U10061 (N_10061,N_9699,N_9761);
or U10062 (N_10062,N_9998,N_9733);
nand U10063 (N_10063,N_9768,N_9859);
xnor U10064 (N_10064,N_9796,N_9786);
nand U10065 (N_10065,N_9804,N_9780);
nand U10066 (N_10066,N_9524,N_9660);
nor U10067 (N_10067,N_9640,N_9824);
nand U10068 (N_10068,N_9886,N_9861);
nor U10069 (N_10069,N_9675,N_9815);
nand U10070 (N_10070,N_9805,N_9978);
nor U10071 (N_10071,N_9759,N_9798);
nand U10072 (N_10072,N_9830,N_9995);
and U10073 (N_10073,N_9932,N_9850);
nor U10074 (N_10074,N_9544,N_9959);
and U10075 (N_10075,N_9613,N_9732);
nor U10076 (N_10076,N_9521,N_9854);
xnor U10077 (N_10077,N_9611,N_9953);
nor U10078 (N_10078,N_9695,N_9662);
or U10079 (N_10079,N_9589,N_9801);
or U10080 (N_10080,N_9972,N_9831);
nor U10081 (N_10081,N_9734,N_9802);
and U10082 (N_10082,N_9599,N_9602);
or U10083 (N_10083,N_9608,N_9534);
nor U10084 (N_10084,N_9651,N_9575);
and U10085 (N_10085,N_9832,N_9723);
or U10086 (N_10086,N_9778,N_9938);
nand U10087 (N_10087,N_9680,N_9944);
and U10088 (N_10088,N_9827,N_9527);
nand U10089 (N_10089,N_9586,N_9532);
nand U10090 (N_10090,N_9705,N_9957);
nand U10091 (N_10091,N_9756,N_9791);
or U10092 (N_10092,N_9503,N_9709);
nor U10093 (N_10093,N_9857,N_9987);
or U10094 (N_10094,N_9750,N_9858);
and U10095 (N_10095,N_9691,N_9840);
nor U10096 (N_10096,N_9725,N_9879);
or U10097 (N_10097,N_9763,N_9724);
or U10098 (N_10098,N_9665,N_9538);
nand U10099 (N_10099,N_9736,N_9677);
xnor U10100 (N_10100,N_9924,N_9674);
xor U10101 (N_10101,N_9645,N_9912);
or U10102 (N_10102,N_9727,N_9726);
xor U10103 (N_10103,N_9583,N_9712);
and U10104 (N_10104,N_9865,N_9603);
or U10105 (N_10105,N_9845,N_9587);
or U10106 (N_10106,N_9835,N_9765);
or U10107 (N_10107,N_9693,N_9698);
nor U10108 (N_10108,N_9510,N_9774);
nor U10109 (N_10109,N_9616,N_9744);
nor U10110 (N_10110,N_9578,N_9951);
or U10111 (N_10111,N_9574,N_9710);
nand U10112 (N_10112,N_9785,N_9537);
and U10113 (N_10113,N_9762,N_9994);
or U10114 (N_10114,N_9560,N_9919);
and U10115 (N_10115,N_9992,N_9990);
nand U10116 (N_10116,N_9794,N_9982);
nand U10117 (N_10117,N_9596,N_9639);
and U10118 (N_10118,N_9707,N_9908);
nor U10119 (N_10119,N_9841,N_9973);
and U10120 (N_10120,N_9971,N_9884);
nor U10121 (N_10121,N_9969,N_9687);
or U10122 (N_10122,N_9729,N_9655);
nand U10123 (N_10123,N_9610,N_9542);
nand U10124 (N_10124,N_9997,N_9891);
nand U10125 (N_10125,N_9739,N_9868);
and U10126 (N_10126,N_9652,N_9748);
or U10127 (N_10127,N_9731,N_9806);
and U10128 (N_10128,N_9916,N_9928);
xor U10129 (N_10129,N_9772,N_9764);
nand U10130 (N_10130,N_9728,N_9682);
nor U10131 (N_10131,N_9819,N_9788);
and U10132 (N_10132,N_9658,N_9941);
and U10133 (N_10133,N_9899,N_9892);
or U10134 (N_10134,N_9881,N_9666);
and U10135 (N_10135,N_9706,N_9563);
nand U10136 (N_10136,N_9925,N_9540);
or U10137 (N_10137,N_9777,N_9570);
and U10138 (N_10138,N_9745,N_9834);
nor U10139 (N_10139,N_9506,N_9738);
and U10140 (N_10140,N_9679,N_9933);
or U10141 (N_10141,N_9811,N_9746);
nand U10142 (N_10142,N_9817,N_9688);
nand U10143 (N_10143,N_9656,N_9797);
xnor U10144 (N_10144,N_9883,N_9880);
nand U10145 (N_10145,N_9979,N_9625);
nand U10146 (N_10146,N_9624,N_9775);
nand U10147 (N_10147,N_9690,N_9647);
nor U10148 (N_10148,N_9989,N_9571);
nand U10149 (N_10149,N_9713,N_9740);
or U10150 (N_10150,N_9668,N_9634);
xnor U10151 (N_10151,N_9898,N_9735);
or U10152 (N_10152,N_9719,N_9895);
xor U10153 (N_10153,N_9991,N_9871);
nor U10154 (N_10154,N_9536,N_9906);
and U10155 (N_10155,N_9535,N_9885);
and U10156 (N_10156,N_9681,N_9747);
or U10157 (N_10157,N_9636,N_9783);
nand U10158 (N_10158,N_9948,N_9800);
and U10159 (N_10159,N_9564,N_9635);
or U10160 (N_10160,N_9893,N_9769);
nor U10161 (N_10161,N_9943,N_9737);
nand U10162 (N_10162,N_9530,N_9838);
nor U10163 (N_10163,N_9721,N_9867);
or U10164 (N_10164,N_9519,N_9814);
nor U10165 (N_10165,N_9685,N_9605);
xor U10166 (N_10166,N_9631,N_9826);
nor U10167 (N_10167,N_9539,N_9526);
or U10168 (N_10168,N_9902,N_9678);
nand U10169 (N_10169,N_9614,N_9582);
nor U10170 (N_10170,N_9518,N_9683);
nand U10171 (N_10171,N_9722,N_9664);
nor U10172 (N_10172,N_9897,N_9661);
and U10173 (N_10173,N_9547,N_9913);
nor U10174 (N_10174,N_9911,N_9790);
nand U10175 (N_10175,N_9915,N_9964);
nand U10176 (N_10176,N_9900,N_9556);
and U10177 (N_10177,N_9757,N_9553);
xnor U10178 (N_10178,N_9601,N_9703);
or U10179 (N_10179,N_9896,N_9593);
or U10180 (N_10180,N_9509,N_9742);
xnor U10181 (N_10181,N_9853,N_9937);
or U10182 (N_10182,N_9961,N_9981);
nand U10183 (N_10183,N_9782,N_9630);
or U10184 (N_10184,N_9592,N_9669);
nor U10185 (N_10185,N_9986,N_9996);
nor U10186 (N_10186,N_9629,N_9934);
nor U10187 (N_10187,N_9626,N_9667);
nor U10188 (N_10188,N_9936,N_9597);
or U10189 (N_10189,N_9595,N_9810);
and U10190 (N_10190,N_9914,N_9657);
nand U10191 (N_10191,N_9887,N_9576);
nor U10192 (N_10192,N_9500,N_9980);
nand U10193 (N_10193,N_9939,N_9905);
and U10194 (N_10194,N_9999,N_9837);
xnor U10195 (N_10195,N_9921,N_9816);
nor U10196 (N_10196,N_9755,N_9692);
or U10197 (N_10197,N_9753,N_9708);
and U10198 (N_10198,N_9702,N_9654);
xnor U10199 (N_10199,N_9809,N_9696);
or U10200 (N_10200,N_9550,N_9808);
nor U10201 (N_10201,N_9910,N_9569);
or U10202 (N_10202,N_9874,N_9642);
nand U10203 (N_10203,N_9670,N_9591);
and U10204 (N_10204,N_9663,N_9517);
or U10205 (N_10205,N_9559,N_9541);
or U10206 (N_10206,N_9546,N_9860);
xnor U10207 (N_10207,N_9795,N_9507);
nand U10208 (N_10208,N_9923,N_9965);
or U10209 (N_10209,N_9966,N_9644);
and U10210 (N_10210,N_9622,N_9872);
and U10211 (N_10211,N_9820,N_9504);
nand U10212 (N_10212,N_9909,N_9985);
or U10213 (N_10213,N_9754,N_9940);
and U10214 (N_10214,N_9792,N_9776);
nand U10215 (N_10215,N_9949,N_9822);
nand U10216 (N_10216,N_9715,N_9648);
and U10217 (N_10217,N_9673,N_9623);
and U10218 (N_10218,N_9848,N_9579);
xnor U10219 (N_10219,N_9770,N_9904);
nor U10220 (N_10220,N_9825,N_9976);
nand U10221 (N_10221,N_9813,N_9638);
nand U10222 (N_10222,N_9590,N_9604);
nand U10223 (N_10223,N_9758,N_9773);
xnor U10224 (N_10224,N_9621,N_9870);
xnor U10225 (N_10225,N_9543,N_9606);
nand U10226 (N_10226,N_9843,N_9513);
nand U10227 (N_10227,N_9694,N_9878);
nor U10228 (N_10228,N_9833,N_9523);
nor U10229 (N_10229,N_9767,N_9977);
or U10230 (N_10230,N_9963,N_9620);
nand U10231 (N_10231,N_9903,N_9983);
and U10232 (N_10232,N_9793,N_9612);
or U10233 (N_10233,N_9975,N_9598);
or U10234 (N_10234,N_9618,N_9760);
nand U10235 (N_10235,N_9577,N_9607);
nor U10236 (N_10236,N_9565,N_9501);
or U10237 (N_10237,N_9787,N_9561);
nor U10238 (N_10238,N_9952,N_9779);
xor U10239 (N_10239,N_9752,N_9942);
nor U10240 (N_10240,N_9581,N_9676);
nand U10241 (N_10241,N_9877,N_9812);
or U10242 (N_10242,N_9818,N_9789);
nor U10243 (N_10243,N_9548,N_9720);
or U10244 (N_10244,N_9927,N_9643);
or U10245 (N_10245,N_9955,N_9922);
or U10246 (N_10246,N_9894,N_9632);
and U10247 (N_10247,N_9917,N_9766);
and U10248 (N_10248,N_9866,N_9968);
xor U10249 (N_10249,N_9888,N_9566);
nor U10250 (N_10250,N_9817,N_9734);
or U10251 (N_10251,N_9776,N_9946);
or U10252 (N_10252,N_9873,N_9736);
or U10253 (N_10253,N_9569,N_9994);
nor U10254 (N_10254,N_9994,N_9576);
nor U10255 (N_10255,N_9846,N_9956);
nand U10256 (N_10256,N_9746,N_9661);
nor U10257 (N_10257,N_9976,N_9650);
nor U10258 (N_10258,N_9596,N_9688);
or U10259 (N_10259,N_9529,N_9611);
nor U10260 (N_10260,N_9866,N_9865);
nor U10261 (N_10261,N_9972,N_9863);
or U10262 (N_10262,N_9809,N_9796);
and U10263 (N_10263,N_9918,N_9914);
nand U10264 (N_10264,N_9648,N_9796);
or U10265 (N_10265,N_9884,N_9925);
nand U10266 (N_10266,N_9708,N_9604);
nor U10267 (N_10267,N_9542,N_9672);
or U10268 (N_10268,N_9862,N_9831);
and U10269 (N_10269,N_9790,N_9979);
or U10270 (N_10270,N_9560,N_9853);
nand U10271 (N_10271,N_9661,N_9534);
or U10272 (N_10272,N_9786,N_9739);
nand U10273 (N_10273,N_9667,N_9753);
or U10274 (N_10274,N_9553,N_9646);
nor U10275 (N_10275,N_9534,N_9578);
and U10276 (N_10276,N_9770,N_9616);
nor U10277 (N_10277,N_9928,N_9598);
xnor U10278 (N_10278,N_9769,N_9656);
nand U10279 (N_10279,N_9561,N_9822);
or U10280 (N_10280,N_9796,N_9660);
or U10281 (N_10281,N_9671,N_9938);
xor U10282 (N_10282,N_9610,N_9979);
and U10283 (N_10283,N_9800,N_9730);
nor U10284 (N_10284,N_9548,N_9604);
nand U10285 (N_10285,N_9885,N_9857);
xor U10286 (N_10286,N_9773,N_9517);
nor U10287 (N_10287,N_9584,N_9757);
or U10288 (N_10288,N_9658,N_9572);
or U10289 (N_10289,N_9788,N_9909);
nand U10290 (N_10290,N_9802,N_9633);
xnor U10291 (N_10291,N_9556,N_9993);
and U10292 (N_10292,N_9548,N_9704);
nor U10293 (N_10293,N_9724,N_9977);
nand U10294 (N_10294,N_9726,N_9918);
and U10295 (N_10295,N_9969,N_9978);
or U10296 (N_10296,N_9873,N_9636);
and U10297 (N_10297,N_9682,N_9689);
xnor U10298 (N_10298,N_9777,N_9981);
or U10299 (N_10299,N_9768,N_9777);
or U10300 (N_10300,N_9914,N_9925);
and U10301 (N_10301,N_9876,N_9739);
and U10302 (N_10302,N_9620,N_9724);
xnor U10303 (N_10303,N_9749,N_9919);
and U10304 (N_10304,N_9886,N_9577);
xnor U10305 (N_10305,N_9742,N_9938);
nand U10306 (N_10306,N_9887,N_9597);
xnor U10307 (N_10307,N_9921,N_9769);
nand U10308 (N_10308,N_9590,N_9794);
nand U10309 (N_10309,N_9719,N_9697);
or U10310 (N_10310,N_9834,N_9890);
and U10311 (N_10311,N_9587,N_9559);
nand U10312 (N_10312,N_9724,N_9797);
or U10313 (N_10313,N_9593,N_9862);
or U10314 (N_10314,N_9903,N_9894);
xor U10315 (N_10315,N_9744,N_9735);
or U10316 (N_10316,N_9843,N_9948);
and U10317 (N_10317,N_9748,N_9712);
nor U10318 (N_10318,N_9839,N_9531);
and U10319 (N_10319,N_9839,N_9704);
nor U10320 (N_10320,N_9728,N_9851);
nand U10321 (N_10321,N_9825,N_9969);
nor U10322 (N_10322,N_9890,N_9930);
or U10323 (N_10323,N_9557,N_9927);
nor U10324 (N_10324,N_9631,N_9951);
nor U10325 (N_10325,N_9571,N_9645);
nand U10326 (N_10326,N_9682,N_9835);
xnor U10327 (N_10327,N_9851,N_9789);
and U10328 (N_10328,N_9895,N_9623);
and U10329 (N_10329,N_9741,N_9578);
xor U10330 (N_10330,N_9941,N_9875);
nand U10331 (N_10331,N_9533,N_9627);
xnor U10332 (N_10332,N_9836,N_9635);
and U10333 (N_10333,N_9537,N_9659);
or U10334 (N_10334,N_9970,N_9885);
and U10335 (N_10335,N_9936,N_9985);
or U10336 (N_10336,N_9689,N_9870);
or U10337 (N_10337,N_9691,N_9921);
nor U10338 (N_10338,N_9961,N_9788);
nor U10339 (N_10339,N_9812,N_9973);
nand U10340 (N_10340,N_9842,N_9515);
nor U10341 (N_10341,N_9871,N_9710);
nor U10342 (N_10342,N_9646,N_9939);
and U10343 (N_10343,N_9817,N_9619);
xor U10344 (N_10344,N_9606,N_9784);
and U10345 (N_10345,N_9543,N_9962);
nand U10346 (N_10346,N_9557,N_9649);
xor U10347 (N_10347,N_9976,N_9637);
or U10348 (N_10348,N_9624,N_9938);
and U10349 (N_10349,N_9842,N_9502);
nand U10350 (N_10350,N_9873,N_9893);
nor U10351 (N_10351,N_9964,N_9709);
and U10352 (N_10352,N_9928,N_9529);
nand U10353 (N_10353,N_9533,N_9978);
or U10354 (N_10354,N_9798,N_9702);
xnor U10355 (N_10355,N_9830,N_9879);
nor U10356 (N_10356,N_9991,N_9597);
or U10357 (N_10357,N_9742,N_9930);
or U10358 (N_10358,N_9858,N_9834);
or U10359 (N_10359,N_9511,N_9501);
xnor U10360 (N_10360,N_9526,N_9645);
or U10361 (N_10361,N_9651,N_9545);
nor U10362 (N_10362,N_9559,N_9923);
nor U10363 (N_10363,N_9557,N_9897);
or U10364 (N_10364,N_9739,N_9993);
nand U10365 (N_10365,N_9638,N_9779);
nor U10366 (N_10366,N_9997,N_9585);
and U10367 (N_10367,N_9646,N_9691);
nand U10368 (N_10368,N_9659,N_9914);
and U10369 (N_10369,N_9719,N_9968);
and U10370 (N_10370,N_9599,N_9871);
and U10371 (N_10371,N_9880,N_9622);
nand U10372 (N_10372,N_9773,N_9548);
and U10373 (N_10373,N_9766,N_9824);
xnor U10374 (N_10374,N_9765,N_9756);
nor U10375 (N_10375,N_9877,N_9576);
xor U10376 (N_10376,N_9542,N_9843);
nor U10377 (N_10377,N_9515,N_9507);
or U10378 (N_10378,N_9834,N_9598);
and U10379 (N_10379,N_9844,N_9866);
xor U10380 (N_10380,N_9547,N_9896);
or U10381 (N_10381,N_9740,N_9608);
nand U10382 (N_10382,N_9906,N_9690);
or U10383 (N_10383,N_9824,N_9508);
nand U10384 (N_10384,N_9736,N_9963);
or U10385 (N_10385,N_9538,N_9862);
and U10386 (N_10386,N_9857,N_9762);
nand U10387 (N_10387,N_9895,N_9981);
nor U10388 (N_10388,N_9631,N_9690);
xor U10389 (N_10389,N_9531,N_9746);
or U10390 (N_10390,N_9941,N_9501);
xor U10391 (N_10391,N_9762,N_9667);
nor U10392 (N_10392,N_9668,N_9962);
xor U10393 (N_10393,N_9686,N_9976);
nand U10394 (N_10394,N_9588,N_9645);
nand U10395 (N_10395,N_9533,N_9811);
and U10396 (N_10396,N_9612,N_9764);
nor U10397 (N_10397,N_9843,N_9611);
nor U10398 (N_10398,N_9748,N_9536);
and U10399 (N_10399,N_9779,N_9749);
nor U10400 (N_10400,N_9804,N_9550);
and U10401 (N_10401,N_9931,N_9811);
and U10402 (N_10402,N_9926,N_9810);
and U10403 (N_10403,N_9991,N_9652);
xor U10404 (N_10404,N_9853,N_9705);
nand U10405 (N_10405,N_9825,N_9709);
nor U10406 (N_10406,N_9972,N_9817);
and U10407 (N_10407,N_9561,N_9747);
nor U10408 (N_10408,N_9960,N_9949);
or U10409 (N_10409,N_9908,N_9913);
nor U10410 (N_10410,N_9803,N_9586);
or U10411 (N_10411,N_9664,N_9899);
nand U10412 (N_10412,N_9994,N_9878);
and U10413 (N_10413,N_9800,N_9575);
or U10414 (N_10414,N_9732,N_9837);
nor U10415 (N_10415,N_9683,N_9675);
or U10416 (N_10416,N_9965,N_9987);
and U10417 (N_10417,N_9571,N_9558);
nor U10418 (N_10418,N_9924,N_9825);
nor U10419 (N_10419,N_9645,N_9623);
nor U10420 (N_10420,N_9655,N_9803);
and U10421 (N_10421,N_9795,N_9717);
and U10422 (N_10422,N_9888,N_9637);
nand U10423 (N_10423,N_9639,N_9643);
nor U10424 (N_10424,N_9577,N_9939);
and U10425 (N_10425,N_9845,N_9772);
or U10426 (N_10426,N_9917,N_9602);
nand U10427 (N_10427,N_9554,N_9862);
and U10428 (N_10428,N_9941,N_9710);
nand U10429 (N_10429,N_9892,N_9614);
or U10430 (N_10430,N_9951,N_9921);
nand U10431 (N_10431,N_9612,N_9979);
nor U10432 (N_10432,N_9966,N_9521);
and U10433 (N_10433,N_9881,N_9919);
nor U10434 (N_10434,N_9998,N_9776);
nand U10435 (N_10435,N_9785,N_9766);
xor U10436 (N_10436,N_9897,N_9547);
and U10437 (N_10437,N_9841,N_9523);
nand U10438 (N_10438,N_9628,N_9572);
xor U10439 (N_10439,N_9715,N_9979);
nor U10440 (N_10440,N_9955,N_9628);
or U10441 (N_10441,N_9991,N_9913);
and U10442 (N_10442,N_9578,N_9977);
xnor U10443 (N_10443,N_9919,N_9832);
nand U10444 (N_10444,N_9551,N_9720);
or U10445 (N_10445,N_9854,N_9751);
or U10446 (N_10446,N_9968,N_9903);
or U10447 (N_10447,N_9950,N_9711);
nor U10448 (N_10448,N_9594,N_9899);
nor U10449 (N_10449,N_9791,N_9825);
nand U10450 (N_10450,N_9660,N_9634);
nand U10451 (N_10451,N_9780,N_9843);
or U10452 (N_10452,N_9628,N_9581);
nand U10453 (N_10453,N_9591,N_9700);
or U10454 (N_10454,N_9504,N_9682);
nand U10455 (N_10455,N_9733,N_9996);
or U10456 (N_10456,N_9650,N_9776);
nand U10457 (N_10457,N_9801,N_9605);
nand U10458 (N_10458,N_9795,N_9518);
or U10459 (N_10459,N_9673,N_9632);
or U10460 (N_10460,N_9942,N_9970);
nand U10461 (N_10461,N_9914,N_9883);
nor U10462 (N_10462,N_9978,N_9621);
or U10463 (N_10463,N_9774,N_9742);
nor U10464 (N_10464,N_9591,N_9943);
nand U10465 (N_10465,N_9516,N_9666);
or U10466 (N_10466,N_9875,N_9675);
nor U10467 (N_10467,N_9782,N_9728);
nand U10468 (N_10468,N_9528,N_9821);
nand U10469 (N_10469,N_9787,N_9630);
nor U10470 (N_10470,N_9775,N_9992);
and U10471 (N_10471,N_9932,N_9692);
and U10472 (N_10472,N_9683,N_9815);
or U10473 (N_10473,N_9632,N_9984);
and U10474 (N_10474,N_9651,N_9905);
nand U10475 (N_10475,N_9897,N_9680);
or U10476 (N_10476,N_9950,N_9687);
and U10477 (N_10477,N_9843,N_9553);
and U10478 (N_10478,N_9891,N_9527);
and U10479 (N_10479,N_9508,N_9672);
and U10480 (N_10480,N_9723,N_9949);
or U10481 (N_10481,N_9636,N_9525);
nor U10482 (N_10482,N_9791,N_9890);
and U10483 (N_10483,N_9968,N_9617);
and U10484 (N_10484,N_9887,N_9935);
and U10485 (N_10485,N_9623,N_9738);
nand U10486 (N_10486,N_9566,N_9775);
nand U10487 (N_10487,N_9510,N_9694);
nor U10488 (N_10488,N_9938,N_9910);
nand U10489 (N_10489,N_9818,N_9527);
and U10490 (N_10490,N_9577,N_9824);
nand U10491 (N_10491,N_9995,N_9903);
nand U10492 (N_10492,N_9765,N_9867);
or U10493 (N_10493,N_9848,N_9748);
and U10494 (N_10494,N_9680,N_9642);
and U10495 (N_10495,N_9743,N_9600);
and U10496 (N_10496,N_9858,N_9727);
or U10497 (N_10497,N_9785,N_9510);
and U10498 (N_10498,N_9928,N_9812);
or U10499 (N_10499,N_9617,N_9970);
nand U10500 (N_10500,N_10465,N_10394);
nand U10501 (N_10501,N_10086,N_10224);
nand U10502 (N_10502,N_10077,N_10450);
nand U10503 (N_10503,N_10326,N_10056);
xor U10504 (N_10504,N_10181,N_10017);
nand U10505 (N_10505,N_10333,N_10339);
nor U10506 (N_10506,N_10197,N_10310);
nor U10507 (N_10507,N_10360,N_10462);
or U10508 (N_10508,N_10327,N_10315);
nor U10509 (N_10509,N_10336,N_10428);
and U10510 (N_10510,N_10121,N_10150);
xnor U10511 (N_10511,N_10448,N_10129);
and U10512 (N_10512,N_10358,N_10031);
and U10513 (N_10513,N_10398,N_10328);
nor U10514 (N_10514,N_10455,N_10162);
nor U10515 (N_10515,N_10187,N_10020);
nor U10516 (N_10516,N_10477,N_10348);
or U10517 (N_10517,N_10209,N_10193);
or U10518 (N_10518,N_10332,N_10330);
nor U10519 (N_10519,N_10101,N_10494);
xor U10520 (N_10520,N_10228,N_10236);
or U10521 (N_10521,N_10104,N_10016);
nand U10522 (N_10522,N_10198,N_10436);
and U10523 (N_10523,N_10276,N_10222);
nand U10524 (N_10524,N_10279,N_10054);
nor U10525 (N_10525,N_10317,N_10269);
nand U10526 (N_10526,N_10190,N_10435);
or U10527 (N_10527,N_10124,N_10257);
nor U10528 (N_10528,N_10291,N_10030);
nand U10529 (N_10529,N_10148,N_10060);
nand U10530 (N_10530,N_10404,N_10309);
nor U10531 (N_10531,N_10136,N_10453);
nand U10532 (N_10532,N_10231,N_10180);
nor U10533 (N_10533,N_10367,N_10290);
nand U10534 (N_10534,N_10306,N_10137);
and U10535 (N_10535,N_10344,N_10161);
and U10536 (N_10536,N_10442,N_10140);
xnor U10537 (N_10537,N_10345,N_10475);
nor U10538 (N_10538,N_10454,N_10083);
nor U10539 (N_10539,N_10098,N_10079);
or U10540 (N_10540,N_10090,N_10250);
nor U10541 (N_10541,N_10211,N_10322);
nor U10542 (N_10542,N_10285,N_10007);
or U10543 (N_10543,N_10068,N_10210);
nor U10544 (N_10544,N_10130,N_10214);
or U10545 (N_10545,N_10029,N_10377);
nor U10546 (N_10546,N_10449,N_10258);
and U10547 (N_10547,N_10393,N_10271);
xor U10548 (N_10548,N_10318,N_10491);
or U10549 (N_10549,N_10260,N_10497);
nand U10550 (N_10550,N_10041,N_10433);
nand U10551 (N_10551,N_10218,N_10202);
nor U10552 (N_10552,N_10125,N_10416);
xor U10553 (N_10553,N_10082,N_10033);
nand U10554 (N_10554,N_10275,N_10414);
or U10555 (N_10555,N_10035,N_10078);
nand U10556 (N_10556,N_10153,N_10149);
nand U10557 (N_10557,N_10157,N_10251);
or U10558 (N_10558,N_10230,N_10468);
nor U10559 (N_10559,N_10429,N_10146);
and U10560 (N_10560,N_10390,N_10164);
nand U10561 (N_10561,N_10132,N_10143);
or U10562 (N_10562,N_10215,N_10112);
or U10563 (N_10563,N_10158,N_10201);
or U10564 (N_10564,N_10354,N_10032);
xnor U10565 (N_10565,N_10311,N_10381);
and U10566 (N_10566,N_10243,N_10365);
or U10567 (N_10567,N_10493,N_10488);
or U10568 (N_10568,N_10061,N_10070);
and U10569 (N_10569,N_10461,N_10034);
and U10570 (N_10570,N_10473,N_10113);
nand U10571 (N_10571,N_10195,N_10357);
nor U10572 (N_10572,N_10200,N_10024);
nor U10573 (N_10573,N_10423,N_10186);
nand U10574 (N_10574,N_10434,N_10019);
and U10575 (N_10575,N_10419,N_10107);
nand U10576 (N_10576,N_10000,N_10499);
or U10577 (N_10577,N_10323,N_10272);
or U10578 (N_10578,N_10350,N_10066);
or U10579 (N_10579,N_10457,N_10298);
and U10580 (N_10580,N_10259,N_10342);
or U10581 (N_10581,N_10430,N_10002);
and U10582 (N_10582,N_10174,N_10165);
nor U10583 (N_10583,N_10478,N_10444);
nor U10584 (N_10584,N_10026,N_10139);
or U10585 (N_10585,N_10183,N_10087);
and U10586 (N_10586,N_10378,N_10239);
xor U10587 (N_10587,N_10463,N_10212);
or U10588 (N_10588,N_10175,N_10154);
nand U10589 (N_10589,N_10100,N_10278);
and U10590 (N_10590,N_10073,N_10128);
xor U10591 (N_10591,N_10103,N_10451);
or U10592 (N_10592,N_10437,N_10076);
nand U10593 (N_10593,N_10400,N_10084);
nand U10594 (N_10594,N_10305,N_10095);
or U10595 (N_10595,N_10293,N_10097);
xor U10596 (N_10596,N_10287,N_10091);
nand U10597 (N_10597,N_10471,N_10395);
or U10598 (N_10598,N_10105,N_10050);
or U10599 (N_10599,N_10168,N_10391);
and U10600 (N_10600,N_10335,N_10343);
or U10601 (N_10601,N_10053,N_10467);
nand U10602 (N_10602,N_10386,N_10267);
xor U10603 (N_10603,N_10221,N_10179);
and U10604 (N_10604,N_10470,N_10123);
and U10605 (N_10605,N_10188,N_10196);
and U10606 (N_10606,N_10152,N_10409);
nor U10607 (N_10607,N_10469,N_10233);
and U10608 (N_10608,N_10014,N_10253);
nor U10609 (N_10609,N_10126,N_10093);
and U10610 (N_10610,N_10118,N_10042);
and U10611 (N_10611,N_10207,N_10134);
nor U10612 (N_10612,N_10415,N_10120);
nand U10613 (N_10613,N_10122,N_10447);
xor U10614 (N_10614,N_10010,N_10159);
or U10615 (N_10615,N_10299,N_10235);
nand U10616 (N_10616,N_10363,N_10319);
and U10617 (N_10617,N_10458,N_10261);
nor U10618 (N_10618,N_10382,N_10191);
or U10619 (N_10619,N_10364,N_10199);
nand U10620 (N_10620,N_10282,N_10421);
and U10621 (N_10621,N_10474,N_10383);
or U10622 (N_10622,N_10156,N_10277);
and U10623 (N_10623,N_10368,N_10237);
nor U10624 (N_10624,N_10001,N_10370);
and U10625 (N_10625,N_10490,N_10227);
and U10626 (N_10626,N_10046,N_10274);
nor U10627 (N_10627,N_10346,N_10301);
nor U10628 (N_10628,N_10265,N_10028);
xnor U10629 (N_10629,N_10460,N_10452);
and U10630 (N_10630,N_10389,N_10044);
nand U10631 (N_10631,N_10362,N_10192);
nand U10632 (N_10632,N_10204,N_10483);
nand U10633 (N_10633,N_10424,N_10388);
or U10634 (N_10634,N_10057,N_10456);
and U10635 (N_10635,N_10387,N_10385);
xnor U10636 (N_10636,N_10425,N_10482);
or U10637 (N_10637,N_10242,N_10485);
nand U10638 (N_10638,N_10422,N_10170);
and U10639 (N_10639,N_10141,N_10255);
nor U10640 (N_10640,N_10480,N_10040);
or U10641 (N_10641,N_10063,N_10206);
or U10642 (N_10642,N_10167,N_10027);
nand U10643 (N_10643,N_10219,N_10037);
nand U10644 (N_10644,N_10441,N_10443);
xor U10645 (N_10645,N_10280,N_10182);
xnor U10646 (N_10646,N_10011,N_10116);
xnor U10647 (N_10647,N_10361,N_10445);
nand U10648 (N_10648,N_10220,N_10374);
and U10649 (N_10649,N_10184,N_10074);
or U10650 (N_10650,N_10427,N_10043);
nand U10651 (N_10651,N_10405,N_10127);
or U10652 (N_10652,N_10402,N_10081);
or U10653 (N_10653,N_10289,N_10321);
xnor U10654 (N_10654,N_10489,N_10142);
or U10655 (N_10655,N_10110,N_10403);
nor U10656 (N_10656,N_10355,N_10418);
xnor U10657 (N_10657,N_10324,N_10244);
or U10658 (N_10658,N_10145,N_10135);
nor U10659 (N_10659,N_10048,N_10108);
and U10660 (N_10660,N_10281,N_10303);
or U10661 (N_10661,N_10325,N_10131);
and U10662 (N_10662,N_10208,N_10366);
nand U10663 (N_10663,N_10439,N_10353);
nor U10664 (N_10664,N_10138,N_10407);
nand U10665 (N_10665,N_10144,N_10334);
nand U10666 (N_10666,N_10397,N_10375);
nor U10667 (N_10667,N_10438,N_10349);
and U10668 (N_10668,N_10234,N_10356);
nand U10669 (N_10669,N_10320,N_10205);
and U10670 (N_10670,N_10304,N_10413);
nand U10671 (N_10671,N_10003,N_10351);
and U10672 (N_10672,N_10039,N_10203);
nand U10673 (N_10673,N_10036,N_10109);
or U10674 (N_10674,N_10246,N_10005);
or U10675 (N_10675,N_10329,N_10059);
nand U10676 (N_10676,N_10292,N_10312);
and U10677 (N_10677,N_10163,N_10295);
nand U10678 (N_10678,N_10012,N_10273);
and U10679 (N_10679,N_10106,N_10459);
nor U10680 (N_10680,N_10399,N_10369);
and U10681 (N_10681,N_10213,N_10006);
or U10682 (N_10682,N_10248,N_10069);
nand U10683 (N_10683,N_10426,N_10194);
nand U10684 (N_10684,N_10294,N_10302);
nor U10685 (N_10685,N_10004,N_10481);
or U10686 (N_10686,N_10071,N_10263);
and U10687 (N_10687,N_10176,N_10252);
and U10688 (N_10688,N_10225,N_10008);
and U10689 (N_10689,N_10058,N_10379);
nor U10690 (N_10690,N_10249,N_10226);
or U10691 (N_10691,N_10371,N_10177);
nor U10692 (N_10692,N_10229,N_10373);
nand U10693 (N_10693,N_10085,N_10245);
xor U10694 (N_10694,N_10065,N_10486);
or U10695 (N_10695,N_10376,N_10216);
xor U10696 (N_10696,N_10062,N_10256);
nand U10697 (N_10697,N_10384,N_10307);
nor U10698 (N_10698,N_10099,N_10052);
nand U10699 (N_10699,N_10406,N_10496);
or U10700 (N_10700,N_10297,N_10264);
nor U10701 (N_10701,N_10313,N_10352);
or U10702 (N_10702,N_10241,N_10338);
and U10703 (N_10703,N_10288,N_10466);
nand U10704 (N_10704,N_10254,N_10392);
nor U10705 (N_10705,N_10015,N_10479);
nand U10706 (N_10706,N_10117,N_10096);
and U10707 (N_10707,N_10240,N_10420);
or U10708 (N_10708,N_10380,N_10038);
nand U10709 (N_10709,N_10172,N_10270);
or U10710 (N_10710,N_10316,N_10396);
and U10711 (N_10711,N_10055,N_10075);
nand U10712 (N_10712,N_10173,N_10492);
nor U10713 (N_10713,N_10331,N_10102);
xnor U10714 (N_10714,N_10412,N_10432);
nor U10715 (N_10715,N_10047,N_10431);
and U10716 (N_10716,N_10092,N_10401);
nor U10717 (N_10717,N_10440,N_10472);
xor U10718 (N_10718,N_10089,N_10049);
nand U10719 (N_10719,N_10022,N_10266);
or U10720 (N_10720,N_10169,N_10171);
nor U10721 (N_10721,N_10147,N_10308);
nand U10722 (N_10722,N_10286,N_10284);
nor U10723 (N_10723,N_10064,N_10088);
nor U10724 (N_10724,N_10223,N_10487);
nor U10725 (N_10725,N_10023,N_10476);
nand U10726 (N_10726,N_10094,N_10341);
nand U10727 (N_10727,N_10114,N_10133);
or U10728 (N_10728,N_10262,N_10025);
and U10729 (N_10729,N_10408,N_10238);
nand U10730 (N_10730,N_10217,N_10268);
or U10731 (N_10731,N_10340,N_10009);
or U10732 (N_10732,N_10296,N_10410);
or U10733 (N_10733,N_10178,N_10347);
or U10734 (N_10734,N_10166,N_10337);
or U10735 (N_10735,N_10495,N_10018);
nor U10736 (N_10736,N_10189,N_10446);
and U10737 (N_10737,N_10045,N_10067);
nand U10738 (N_10738,N_10160,N_10464);
or U10739 (N_10739,N_10151,N_10283);
xnor U10740 (N_10740,N_10372,N_10115);
nor U10741 (N_10741,N_10013,N_10111);
or U10742 (N_10742,N_10359,N_10247);
nand U10743 (N_10743,N_10021,N_10119);
nand U10744 (N_10744,N_10051,N_10232);
and U10745 (N_10745,N_10314,N_10417);
xnor U10746 (N_10746,N_10072,N_10300);
nand U10747 (N_10747,N_10185,N_10155);
and U10748 (N_10748,N_10080,N_10411);
or U10749 (N_10749,N_10484,N_10498);
or U10750 (N_10750,N_10478,N_10042);
nor U10751 (N_10751,N_10294,N_10387);
or U10752 (N_10752,N_10268,N_10424);
or U10753 (N_10753,N_10319,N_10445);
xor U10754 (N_10754,N_10174,N_10183);
or U10755 (N_10755,N_10429,N_10035);
nor U10756 (N_10756,N_10171,N_10218);
or U10757 (N_10757,N_10088,N_10198);
and U10758 (N_10758,N_10196,N_10332);
or U10759 (N_10759,N_10472,N_10147);
nor U10760 (N_10760,N_10291,N_10161);
or U10761 (N_10761,N_10497,N_10136);
nor U10762 (N_10762,N_10495,N_10117);
nor U10763 (N_10763,N_10460,N_10030);
or U10764 (N_10764,N_10447,N_10487);
or U10765 (N_10765,N_10217,N_10375);
or U10766 (N_10766,N_10438,N_10324);
nor U10767 (N_10767,N_10267,N_10217);
xnor U10768 (N_10768,N_10457,N_10180);
or U10769 (N_10769,N_10150,N_10185);
or U10770 (N_10770,N_10473,N_10186);
nand U10771 (N_10771,N_10247,N_10442);
or U10772 (N_10772,N_10430,N_10397);
or U10773 (N_10773,N_10095,N_10296);
nor U10774 (N_10774,N_10312,N_10330);
nor U10775 (N_10775,N_10440,N_10253);
nand U10776 (N_10776,N_10361,N_10140);
nand U10777 (N_10777,N_10410,N_10475);
nand U10778 (N_10778,N_10002,N_10297);
or U10779 (N_10779,N_10239,N_10411);
nor U10780 (N_10780,N_10310,N_10086);
or U10781 (N_10781,N_10148,N_10053);
or U10782 (N_10782,N_10372,N_10315);
or U10783 (N_10783,N_10480,N_10361);
nand U10784 (N_10784,N_10341,N_10150);
nor U10785 (N_10785,N_10468,N_10106);
nand U10786 (N_10786,N_10467,N_10002);
or U10787 (N_10787,N_10494,N_10076);
xor U10788 (N_10788,N_10475,N_10483);
xnor U10789 (N_10789,N_10378,N_10026);
and U10790 (N_10790,N_10134,N_10230);
nand U10791 (N_10791,N_10242,N_10225);
or U10792 (N_10792,N_10483,N_10255);
xnor U10793 (N_10793,N_10125,N_10092);
or U10794 (N_10794,N_10174,N_10346);
or U10795 (N_10795,N_10100,N_10383);
and U10796 (N_10796,N_10365,N_10059);
or U10797 (N_10797,N_10370,N_10406);
and U10798 (N_10798,N_10151,N_10115);
nand U10799 (N_10799,N_10178,N_10227);
or U10800 (N_10800,N_10161,N_10426);
and U10801 (N_10801,N_10397,N_10187);
nor U10802 (N_10802,N_10003,N_10454);
and U10803 (N_10803,N_10357,N_10386);
nor U10804 (N_10804,N_10219,N_10005);
nand U10805 (N_10805,N_10178,N_10344);
nand U10806 (N_10806,N_10493,N_10131);
or U10807 (N_10807,N_10276,N_10230);
and U10808 (N_10808,N_10204,N_10145);
nor U10809 (N_10809,N_10484,N_10050);
or U10810 (N_10810,N_10347,N_10018);
or U10811 (N_10811,N_10171,N_10325);
nand U10812 (N_10812,N_10133,N_10102);
nor U10813 (N_10813,N_10383,N_10115);
or U10814 (N_10814,N_10000,N_10291);
nand U10815 (N_10815,N_10451,N_10196);
and U10816 (N_10816,N_10007,N_10145);
xor U10817 (N_10817,N_10221,N_10426);
and U10818 (N_10818,N_10308,N_10172);
nor U10819 (N_10819,N_10360,N_10159);
or U10820 (N_10820,N_10130,N_10460);
or U10821 (N_10821,N_10463,N_10291);
and U10822 (N_10822,N_10374,N_10237);
nor U10823 (N_10823,N_10199,N_10065);
or U10824 (N_10824,N_10311,N_10257);
or U10825 (N_10825,N_10439,N_10051);
and U10826 (N_10826,N_10457,N_10177);
nand U10827 (N_10827,N_10148,N_10301);
and U10828 (N_10828,N_10062,N_10477);
and U10829 (N_10829,N_10065,N_10346);
or U10830 (N_10830,N_10360,N_10213);
and U10831 (N_10831,N_10078,N_10451);
or U10832 (N_10832,N_10441,N_10356);
or U10833 (N_10833,N_10444,N_10458);
and U10834 (N_10834,N_10409,N_10314);
nand U10835 (N_10835,N_10097,N_10353);
or U10836 (N_10836,N_10165,N_10222);
xor U10837 (N_10837,N_10037,N_10281);
and U10838 (N_10838,N_10127,N_10276);
or U10839 (N_10839,N_10499,N_10393);
nor U10840 (N_10840,N_10236,N_10151);
nor U10841 (N_10841,N_10262,N_10247);
or U10842 (N_10842,N_10363,N_10311);
and U10843 (N_10843,N_10168,N_10027);
or U10844 (N_10844,N_10315,N_10032);
nand U10845 (N_10845,N_10339,N_10462);
or U10846 (N_10846,N_10432,N_10440);
or U10847 (N_10847,N_10217,N_10180);
nand U10848 (N_10848,N_10005,N_10153);
xnor U10849 (N_10849,N_10398,N_10301);
and U10850 (N_10850,N_10450,N_10412);
nand U10851 (N_10851,N_10011,N_10234);
nor U10852 (N_10852,N_10148,N_10137);
xnor U10853 (N_10853,N_10115,N_10459);
or U10854 (N_10854,N_10122,N_10256);
nand U10855 (N_10855,N_10419,N_10432);
and U10856 (N_10856,N_10180,N_10161);
and U10857 (N_10857,N_10476,N_10489);
nor U10858 (N_10858,N_10368,N_10119);
or U10859 (N_10859,N_10430,N_10187);
nor U10860 (N_10860,N_10270,N_10356);
nor U10861 (N_10861,N_10089,N_10401);
and U10862 (N_10862,N_10010,N_10076);
nor U10863 (N_10863,N_10343,N_10416);
or U10864 (N_10864,N_10299,N_10002);
nor U10865 (N_10865,N_10141,N_10360);
nand U10866 (N_10866,N_10014,N_10064);
and U10867 (N_10867,N_10332,N_10075);
xnor U10868 (N_10868,N_10199,N_10333);
nor U10869 (N_10869,N_10098,N_10473);
xor U10870 (N_10870,N_10292,N_10085);
nor U10871 (N_10871,N_10351,N_10274);
nor U10872 (N_10872,N_10406,N_10492);
or U10873 (N_10873,N_10438,N_10047);
nor U10874 (N_10874,N_10040,N_10046);
nor U10875 (N_10875,N_10451,N_10228);
or U10876 (N_10876,N_10211,N_10093);
or U10877 (N_10877,N_10156,N_10118);
nand U10878 (N_10878,N_10080,N_10040);
nand U10879 (N_10879,N_10303,N_10112);
and U10880 (N_10880,N_10464,N_10473);
and U10881 (N_10881,N_10260,N_10131);
and U10882 (N_10882,N_10095,N_10082);
nand U10883 (N_10883,N_10408,N_10276);
and U10884 (N_10884,N_10224,N_10214);
or U10885 (N_10885,N_10396,N_10249);
and U10886 (N_10886,N_10160,N_10444);
xor U10887 (N_10887,N_10354,N_10346);
and U10888 (N_10888,N_10195,N_10256);
and U10889 (N_10889,N_10464,N_10262);
nor U10890 (N_10890,N_10251,N_10380);
or U10891 (N_10891,N_10263,N_10451);
and U10892 (N_10892,N_10472,N_10032);
and U10893 (N_10893,N_10321,N_10435);
nand U10894 (N_10894,N_10065,N_10144);
nand U10895 (N_10895,N_10154,N_10052);
nand U10896 (N_10896,N_10222,N_10064);
or U10897 (N_10897,N_10058,N_10334);
nand U10898 (N_10898,N_10360,N_10150);
nand U10899 (N_10899,N_10004,N_10346);
nand U10900 (N_10900,N_10391,N_10486);
nor U10901 (N_10901,N_10429,N_10348);
nor U10902 (N_10902,N_10041,N_10158);
nand U10903 (N_10903,N_10074,N_10094);
and U10904 (N_10904,N_10053,N_10213);
nor U10905 (N_10905,N_10250,N_10488);
nand U10906 (N_10906,N_10194,N_10384);
nor U10907 (N_10907,N_10403,N_10332);
nor U10908 (N_10908,N_10398,N_10302);
xor U10909 (N_10909,N_10226,N_10106);
nor U10910 (N_10910,N_10154,N_10483);
or U10911 (N_10911,N_10245,N_10110);
or U10912 (N_10912,N_10456,N_10087);
and U10913 (N_10913,N_10380,N_10382);
nor U10914 (N_10914,N_10391,N_10451);
nor U10915 (N_10915,N_10375,N_10314);
nor U10916 (N_10916,N_10171,N_10334);
and U10917 (N_10917,N_10286,N_10370);
or U10918 (N_10918,N_10220,N_10379);
nor U10919 (N_10919,N_10096,N_10075);
and U10920 (N_10920,N_10155,N_10031);
or U10921 (N_10921,N_10419,N_10173);
or U10922 (N_10922,N_10374,N_10142);
xor U10923 (N_10923,N_10418,N_10285);
nor U10924 (N_10924,N_10352,N_10463);
nor U10925 (N_10925,N_10420,N_10020);
or U10926 (N_10926,N_10162,N_10426);
nand U10927 (N_10927,N_10231,N_10046);
nor U10928 (N_10928,N_10007,N_10026);
nor U10929 (N_10929,N_10493,N_10027);
or U10930 (N_10930,N_10310,N_10043);
nand U10931 (N_10931,N_10292,N_10205);
or U10932 (N_10932,N_10192,N_10396);
and U10933 (N_10933,N_10288,N_10348);
or U10934 (N_10934,N_10470,N_10405);
nor U10935 (N_10935,N_10126,N_10350);
nor U10936 (N_10936,N_10292,N_10157);
nand U10937 (N_10937,N_10001,N_10368);
or U10938 (N_10938,N_10201,N_10227);
nor U10939 (N_10939,N_10186,N_10205);
or U10940 (N_10940,N_10423,N_10135);
nor U10941 (N_10941,N_10177,N_10042);
and U10942 (N_10942,N_10216,N_10300);
or U10943 (N_10943,N_10286,N_10275);
and U10944 (N_10944,N_10175,N_10384);
nor U10945 (N_10945,N_10125,N_10123);
or U10946 (N_10946,N_10423,N_10407);
and U10947 (N_10947,N_10037,N_10430);
or U10948 (N_10948,N_10352,N_10319);
nor U10949 (N_10949,N_10492,N_10360);
nand U10950 (N_10950,N_10281,N_10341);
nor U10951 (N_10951,N_10182,N_10413);
or U10952 (N_10952,N_10272,N_10063);
nand U10953 (N_10953,N_10011,N_10127);
and U10954 (N_10954,N_10013,N_10098);
xor U10955 (N_10955,N_10235,N_10485);
nor U10956 (N_10956,N_10243,N_10422);
xnor U10957 (N_10957,N_10074,N_10251);
and U10958 (N_10958,N_10141,N_10393);
or U10959 (N_10959,N_10101,N_10035);
nand U10960 (N_10960,N_10020,N_10150);
nand U10961 (N_10961,N_10084,N_10010);
and U10962 (N_10962,N_10145,N_10231);
nor U10963 (N_10963,N_10165,N_10423);
nand U10964 (N_10964,N_10085,N_10179);
or U10965 (N_10965,N_10170,N_10417);
nor U10966 (N_10966,N_10404,N_10418);
nor U10967 (N_10967,N_10069,N_10475);
nand U10968 (N_10968,N_10156,N_10248);
nor U10969 (N_10969,N_10387,N_10446);
nand U10970 (N_10970,N_10479,N_10220);
nor U10971 (N_10971,N_10359,N_10123);
nor U10972 (N_10972,N_10467,N_10184);
and U10973 (N_10973,N_10055,N_10100);
nand U10974 (N_10974,N_10333,N_10216);
nor U10975 (N_10975,N_10288,N_10307);
nand U10976 (N_10976,N_10145,N_10015);
or U10977 (N_10977,N_10440,N_10129);
nand U10978 (N_10978,N_10383,N_10085);
nor U10979 (N_10979,N_10164,N_10100);
or U10980 (N_10980,N_10244,N_10322);
and U10981 (N_10981,N_10087,N_10013);
nand U10982 (N_10982,N_10013,N_10017);
xor U10983 (N_10983,N_10111,N_10131);
or U10984 (N_10984,N_10368,N_10272);
or U10985 (N_10985,N_10281,N_10147);
or U10986 (N_10986,N_10063,N_10122);
and U10987 (N_10987,N_10119,N_10213);
and U10988 (N_10988,N_10086,N_10334);
xor U10989 (N_10989,N_10377,N_10417);
nor U10990 (N_10990,N_10240,N_10490);
nand U10991 (N_10991,N_10154,N_10149);
nor U10992 (N_10992,N_10319,N_10084);
or U10993 (N_10993,N_10105,N_10143);
nand U10994 (N_10994,N_10437,N_10180);
nor U10995 (N_10995,N_10452,N_10419);
xor U10996 (N_10996,N_10368,N_10483);
and U10997 (N_10997,N_10065,N_10347);
or U10998 (N_10998,N_10265,N_10250);
and U10999 (N_10999,N_10191,N_10047);
or U11000 (N_11000,N_10713,N_10564);
or U11001 (N_11001,N_10531,N_10605);
and U11002 (N_11002,N_10970,N_10636);
nor U11003 (N_11003,N_10637,N_10642);
or U11004 (N_11004,N_10911,N_10826);
or U11005 (N_11005,N_10517,N_10542);
nor U11006 (N_11006,N_10701,N_10891);
xnor U11007 (N_11007,N_10855,N_10766);
nand U11008 (N_11008,N_10723,N_10833);
nor U11009 (N_11009,N_10575,N_10880);
and U11010 (N_11010,N_10850,N_10789);
nand U11011 (N_11011,N_10870,N_10569);
nand U11012 (N_11012,N_10595,N_10620);
or U11013 (N_11013,N_10980,N_10960);
and U11014 (N_11014,N_10614,N_10594);
nor U11015 (N_11015,N_10600,N_10705);
nor U11016 (N_11016,N_10873,N_10721);
or U11017 (N_11017,N_10938,N_10793);
nand U11018 (N_11018,N_10975,N_10769);
and U11019 (N_11019,N_10607,N_10592);
nand U11020 (N_11020,N_10673,N_10887);
nand U11021 (N_11021,N_10651,N_10667);
xor U11022 (N_11022,N_10708,N_10871);
nor U11023 (N_11023,N_10553,N_10982);
or U11024 (N_11024,N_10953,N_10612);
nand U11025 (N_11025,N_10881,N_10545);
or U11026 (N_11026,N_10778,N_10699);
nand U11027 (N_11027,N_10583,N_10886);
and U11028 (N_11028,N_10951,N_10985);
xnor U11029 (N_11029,N_10693,N_10958);
and U11030 (N_11030,N_10889,N_10779);
nand U11031 (N_11031,N_10906,N_10918);
or U11032 (N_11032,N_10734,N_10525);
nand U11033 (N_11033,N_10901,N_10824);
nor U11034 (N_11034,N_10967,N_10613);
nor U11035 (N_11035,N_10610,N_10659);
and U11036 (N_11036,N_10512,N_10672);
or U11037 (N_11037,N_10758,N_10502);
or U11038 (N_11038,N_10956,N_10922);
nand U11039 (N_11039,N_10908,N_10926);
or U11040 (N_11040,N_10562,N_10859);
xor U11041 (N_11041,N_10581,N_10747);
xnor U11042 (N_11042,N_10897,N_10552);
or U11043 (N_11043,N_10681,N_10803);
xor U11044 (N_11044,N_10930,N_10624);
nand U11045 (N_11045,N_10559,N_10692);
or U11046 (N_11046,N_10959,N_10998);
and U11047 (N_11047,N_10907,N_10650);
nor U11048 (N_11048,N_10913,N_10706);
nand U11049 (N_11049,N_10749,N_10832);
xor U11050 (N_11050,N_10523,N_10626);
xnor U11051 (N_11051,N_10878,N_10720);
nand U11052 (N_11052,N_10671,N_10649);
nor U11053 (N_11053,N_10729,N_10606);
nor U11054 (N_11054,N_10952,N_10932);
or U11055 (N_11055,N_10971,N_10522);
or U11056 (N_11056,N_10972,N_10900);
and U11057 (N_11057,N_10634,N_10576);
xor U11058 (N_11058,N_10896,N_10752);
and U11059 (N_11059,N_10532,N_10568);
and U11060 (N_11060,N_10947,N_10806);
or U11061 (N_11061,N_10735,N_10822);
and U11062 (N_11062,N_10656,N_10519);
nor U11063 (N_11063,N_10820,N_10928);
xor U11064 (N_11064,N_10995,N_10578);
nor U11065 (N_11065,N_10988,N_10515);
nor U11066 (N_11066,N_10917,N_10762);
nand U11067 (N_11067,N_10551,N_10739);
nand U11068 (N_11068,N_10899,N_10895);
nand U11069 (N_11069,N_10848,N_10537);
nor U11070 (N_11070,N_10776,N_10661);
nand U11071 (N_11071,N_10579,N_10787);
nor U11072 (N_11072,N_10834,N_10535);
nor U11073 (N_11073,N_10984,N_10567);
and U11074 (N_11074,N_10709,N_10775);
and U11075 (N_11075,N_10697,N_10548);
and U11076 (N_11076,N_10664,N_10527);
or U11077 (N_11077,N_10738,N_10754);
nand U11078 (N_11078,N_10539,N_10916);
and U11079 (N_11079,N_10874,N_10753);
or U11080 (N_11080,N_10811,N_10828);
xnor U11081 (N_11081,N_10827,N_10601);
nor U11082 (N_11082,N_10732,N_10768);
and U11083 (N_11083,N_10763,N_10508);
and U11084 (N_11084,N_10915,N_10630);
nor U11085 (N_11085,N_10815,N_10597);
xor U11086 (N_11086,N_10587,N_10838);
and U11087 (N_11087,N_10898,N_10751);
and U11088 (N_11088,N_10547,N_10509);
nand U11089 (N_11089,N_10783,N_10929);
or U11090 (N_11090,N_10686,N_10726);
and U11091 (N_11091,N_10676,N_10872);
nand U11092 (N_11092,N_10658,N_10809);
nand U11093 (N_11093,N_10611,N_10879);
nor U11094 (N_11094,N_10847,N_10841);
nand U11095 (N_11095,N_10544,N_10555);
and U11096 (N_11096,N_10866,N_10863);
and U11097 (N_11097,N_10882,N_10640);
nor U11098 (N_11098,N_10849,N_10703);
and U11099 (N_11099,N_10528,N_10730);
nand U11100 (N_11100,N_10641,N_10668);
nand U11101 (N_11101,N_10615,N_10644);
and U11102 (N_11102,N_10860,N_10976);
and U11103 (N_11103,N_10633,N_10944);
nand U11104 (N_11104,N_10660,N_10556);
and U11105 (N_11105,N_10890,N_10629);
and U11106 (N_11106,N_10510,N_10830);
nand U11107 (N_11107,N_10797,N_10513);
nor U11108 (N_11108,N_10816,N_10566);
and U11109 (N_11109,N_10961,N_10987);
or U11110 (N_11110,N_10883,N_10999);
nor U11111 (N_11111,N_10835,N_10782);
xor U11112 (N_11112,N_10557,N_10974);
nand U11113 (N_11113,N_10694,N_10675);
or U11114 (N_11114,N_10757,N_10840);
or U11115 (N_11115,N_10590,N_10585);
or U11116 (N_11116,N_10867,N_10790);
nor U11117 (N_11117,N_10875,N_10647);
nand U11118 (N_11118,N_10563,N_10571);
and U11119 (N_11119,N_10942,N_10925);
nand U11120 (N_11120,N_10996,N_10618);
nor U11121 (N_11121,N_10819,N_10679);
and U11122 (N_11122,N_10717,N_10698);
nor U11123 (N_11123,N_10628,N_10989);
and U11124 (N_11124,N_10623,N_10934);
or U11125 (N_11125,N_10530,N_10565);
nor U11126 (N_11126,N_10700,N_10716);
and U11127 (N_11127,N_10981,N_10791);
or U11128 (N_11128,N_10851,N_10943);
xor U11129 (N_11129,N_10941,N_10977);
nand U11130 (N_11130,N_10737,N_10818);
and U11131 (N_11131,N_10696,N_10731);
or U11132 (N_11132,N_10514,N_10712);
or U11133 (N_11133,N_10631,N_10584);
and U11134 (N_11134,N_10598,N_10529);
nand U11135 (N_11135,N_10654,N_10923);
or U11136 (N_11136,N_10858,N_10829);
nand U11137 (N_11137,N_10939,N_10736);
nor U11138 (N_11138,N_10733,N_10572);
nand U11139 (N_11139,N_10946,N_10655);
nor U11140 (N_11140,N_10677,N_10994);
or U11141 (N_11141,N_10516,N_10920);
and U11142 (N_11142,N_10505,N_10639);
and U11143 (N_11143,N_10670,N_10558);
nor U11144 (N_11144,N_10885,N_10905);
and U11145 (N_11145,N_10741,N_10662);
nand U11146 (N_11146,N_10540,N_10596);
and U11147 (N_11147,N_10543,N_10893);
or U11148 (N_11148,N_10921,N_10504);
nor U11149 (N_11149,N_10798,N_10714);
xnor U11150 (N_11150,N_10936,N_10894);
xnor U11151 (N_11151,N_10854,N_10799);
nand U11152 (N_11152,N_10876,N_10715);
or U11153 (N_11153,N_10627,N_10501);
nor U11154 (N_11154,N_10777,N_10805);
and U11155 (N_11155,N_10781,N_10550);
or U11156 (N_11156,N_10533,N_10538);
nand U11157 (N_11157,N_10743,N_10807);
nor U11158 (N_11158,N_10765,N_10570);
nand U11159 (N_11159,N_10617,N_10760);
nand U11160 (N_11160,N_10520,N_10742);
or U11161 (N_11161,N_10902,N_10804);
nor U11162 (N_11162,N_10688,N_10521);
nand U11163 (N_11163,N_10622,N_10912);
or U11164 (N_11164,N_10560,N_10586);
xor U11165 (N_11165,N_10577,N_10648);
xor U11166 (N_11166,N_10524,N_10674);
and U11167 (N_11167,N_10914,N_10591);
nand U11168 (N_11168,N_10582,N_10711);
and U11169 (N_11169,N_10653,N_10856);
xor U11170 (N_11170,N_10549,N_10964);
or U11171 (N_11171,N_10842,N_10904);
xor U11172 (N_11172,N_10574,N_10831);
nor U11173 (N_11173,N_10945,N_10969);
or U11174 (N_11174,N_10621,N_10632);
or U11175 (N_11175,N_10526,N_10868);
nor U11176 (N_11176,N_10643,N_10973);
or U11177 (N_11177,N_10746,N_10580);
or U11178 (N_11178,N_10852,N_10966);
nand U11179 (N_11179,N_10652,N_10604);
nor U11180 (N_11180,N_10599,N_10690);
and U11181 (N_11181,N_10800,N_10718);
nor U11182 (N_11182,N_10707,N_10684);
nor U11183 (N_11183,N_10955,N_10808);
xor U11184 (N_11184,N_10761,N_10755);
nand U11185 (N_11185,N_10957,N_10728);
and U11186 (N_11186,N_10845,N_10744);
nand U11187 (N_11187,N_10810,N_10919);
nand U11188 (N_11188,N_10954,N_10986);
or U11189 (N_11189,N_10602,N_10722);
nand U11190 (N_11190,N_10619,N_10680);
or U11191 (N_11191,N_10993,N_10903);
xor U11192 (N_11192,N_10862,N_10719);
or U11193 (N_11193,N_10979,N_10573);
nand U11194 (N_11194,N_10853,N_10931);
nand U11195 (N_11195,N_10518,N_10927);
nor U11196 (N_11196,N_10812,N_10949);
or U11197 (N_11197,N_10638,N_10704);
or U11198 (N_11198,N_10821,N_10937);
or U11199 (N_11199,N_10865,N_10978);
nand U11200 (N_11200,N_10546,N_10666);
and U11201 (N_11201,N_10817,N_10635);
nand U11202 (N_11202,N_10503,N_10933);
and U11203 (N_11203,N_10935,N_10770);
nand U11204 (N_11204,N_10507,N_10593);
nand U11205 (N_11205,N_10691,N_10784);
xnor U11206 (N_11206,N_10843,N_10864);
and U11207 (N_11207,N_10685,N_10780);
and U11208 (N_11208,N_10861,N_10813);
nor U11209 (N_11209,N_10963,N_10687);
nor U11210 (N_11210,N_10796,N_10801);
nand U11211 (N_11211,N_10561,N_10663);
xnor U11212 (N_11212,N_10702,N_10603);
nor U11213 (N_11213,N_10657,N_10825);
nand U11214 (N_11214,N_10990,N_10740);
and U11215 (N_11215,N_10892,N_10534);
xnor U11216 (N_11216,N_10727,N_10506);
nand U11217 (N_11217,N_10997,N_10725);
nand U11218 (N_11218,N_10962,N_10645);
or U11219 (N_11219,N_10837,N_10788);
nor U11220 (N_11220,N_10759,N_10609);
or U11221 (N_11221,N_10771,N_10802);
nor U11222 (N_11222,N_10772,N_10625);
and U11223 (N_11223,N_10869,N_10616);
or U11224 (N_11224,N_10750,N_10724);
xor U11225 (N_11225,N_10589,N_10745);
and U11226 (N_11226,N_10948,N_10511);
nor U11227 (N_11227,N_10554,N_10500);
nand U11228 (N_11228,N_10968,N_10940);
or U11229 (N_11229,N_10924,N_10669);
or U11230 (N_11230,N_10541,N_10665);
and U11231 (N_11231,N_10785,N_10682);
xor U11232 (N_11232,N_10764,N_10823);
nand U11233 (N_11233,N_10767,N_10857);
nor U11234 (N_11234,N_10608,N_10646);
and U11235 (N_11235,N_10992,N_10588);
xnor U11236 (N_11236,N_10689,N_10991);
nor U11237 (N_11237,N_10536,N_10877);
or U11238 (N_11238,N_10794,N_10909);
nor U11239 (N_11239,N_10888,N_10773);
or U11240 (N_11240,N_10756,N_10683);
and U11241 (N_11241,N_10795,N_10846);
and U11242 (N_11242,N_10678,N_10950);
nand U11243 (N_11243,N_10844,N_10748);
nor U11244 (N_11244,N_10710,N_10792);
or U11245 (N_11245,N_10839,N_10695);
nor U11246 (N_11246,N_10786,N_10774);
nor U11247 (N_11247,N_10884,N_10983);
nand U11248 (N_11248,N_10965,N_10836);
nor U11249 (N_11249,N_10910,N_10814);
nand U11250 (N_11250,N_10986,N_10562);
or U11251 (N_11251,N_10896,N_10894);
nor U11252 (N_11252,N_10783,N_10807);
or U11253 (N_11253,N_10517,N_10931);
nand U11254 (N_11254,N_10612,N_10879);
xor U11255 (N_11255,N_10618,N_10984);
nor U11256 (N_11256,N_10615,N_10617);
nand U11257 (N_11257,N_10730,N_10510);
xnor U11258 (N_11258,N_10997,N_10833);
nand U11259 (N_11259,N_10677,N_10515);
and U11260 (N_11260,N_10998,N_10834);
and U11261 (N_11261,N_10829,N_10653);
nand U11262 (N_11262,N_10558,N_10766);
nand U11263 (N_11263,N_10799,N_10979);
nand U11264 (N_11264,N_10523,N_10517);
xnor U11265 (N_11265,N_10584,N_10604);
nand U11266 (N_11266,N_10617,N_10953);
and U11267 (N_11267,N_10543,N_10971);
or U11268 (N_11268,N_10551,N_10560);
or U11269 (N_11269,N_10755,N_10956);
or U11270 (N_11270,N_10942,N_10845);
nand U11271 (N_11271,N_10581,N_10996);
or U11272 (N_11272,N_10513,N_10983);
nor U11273 (N_11273,N_10857,N_10663);
or U11274 (N_11274,N_10681,N_10669);
nor U11275 (N_11275,N_10737,N_10655);
nand U11276 (N_11276,N_10646,N_10580);
nor U11277 (N_11277,N_10707,N_10546);
nand U11278 (N_11278,N_10924,N_10876);
xor U11279 (N_11279,N_10600,N_10759);
and U11280 (N_11280,N_10574,N_10928);
nand U11281 (N_11281,N_10611,N_10644);
or U11282 (N_11282,N_10643,N_10883);
and U11283 (N_11283,N_10765,N_10736);
nor U11284 (N_11284,N_10669,N_10971);
nor U11285 (N_11285,N_10786,N_10936);
and U11286 (N_11286,N_10772,N_10540);
nor U11287 (N_11287,N_10527,N_10836);
nor U11288 (N_11288,N_10670,N_10763);
nand U11289 (N_11289,N_10775,N_10873);
or U11290 (N_11290,N_10942,N_10758);
or U11291 (N_11291,N_10796,N_10585);
nor U11292 (N_11292,N_10846,N_10504);
or U11293 (N_11293,N_10518,N_10800);
and U11294 (N_11294,N_10608,N_10676);
nor U11295 (N_11295,N_10760,N_10766);
and U11296 (N_11296,N_10840,N_10853);
nand U11297 (N_11297,N_10721,N_10576);
or U11298 (N_11298,N_10620,N_10851);
or U11299 (N_11299,N_10937,N_10851);
nand U11300 (N_11300,N_10841,N_10633);
nor U11301 (N_11301,N_10648,N_10820);
nand U11302 (N_11302,N_10989,N_10945);
nand U11303 (N_11303,N_10832,N_10614);
xnor U11304 (N_11304,N_10536,N_10713);
xnor U11305 (N_11305,N_10911,N_10795);
nand U11306 (N_11306,N_10913,N_10701);
or U11307 (N_11307,N_10866,N_10525);
nand U11308 (N_11308,N_10519,N_10954);
nand U11309 (N_11309,N_10722,N_10801);
xor U11310 (N_11310,N_10679,N_10997);
and U11311 (N_11311,N_10791,N_10992);
and U11312 (N_11312,N_10969,N_10536);
xnor U11313 (N_11313,N_10900,N_10641);
or U11314 (N_11314,N_10577,N_10726);
or U11315 (N_11315,N_10560,N_10512);
nor U11316 (N_11316,N_10873,N_10817);
nand U11317 (N_11317,N_10770,N_10998);
and U11318 (N_11318,N_10935,N_10910);
xnor U11319 (N_11319,N_10788,N_10832);
or U11320 (N_11320,N_10976,N_10710);
or U11321 (N_11321,N_10638,N_10775);
and U11322 (N_11322,N_10973,N_10935);
and U11323 (N_11323,N_10501,N_10697);
and U11324 (N_11324,N_10976,N_10729);
nor U11325 (N_11325,N_10987,N_10878);
xnor U11326 (N_11326,N_10901,N_10727);
and U11327 (N_11327,N_10662,N_10962);
nand U11328 (N_11328,N_10862,N_10598);
nor U11329 (N_11329,N_10973,N_10772);
nor U11330 (N_11330,N_10618,N_10919);
and U11331 (N_11331,N_10694,N_10531);
nor U11332 (N_11332,N_10961,N_10744);
nor U11333 (N_11333,N_10970,N_10736);
nor U11334 (N_11334,N_10688,N_10728);
nor U11335 (N_11335,N_10504,N_10757);
and U11336 (N_11336,N_10695,N_10676);
and U11337 (N_11337,N_10897,N_10711);
nor U11338 (N_11338,N_10608,N_10616);
nand U11339 (N_11339,N_10940,N_10990);
nand U11340 (N_11340,N_10813,N_10735);
and U11341 (N_11341,N_10528,N_10716);
nand U11342 (N_11342,N_10546,N_10968);
or U11343 (N_11343,N_10537,N_10776);
or U11344 (N_11344,N_10818,N_10794);
nand U11345 (N_11345,N_10697,N_10884);
or U11346 (N_11346,N_10967,N_10522);
nor U11347 (N_11347,N_10856,N_10718);
nor U11348 (N_11348,N_10739,N_10620);
or U11349 (N_11349,N_10769,N_10632);
and U11350 (N_11350,N_10843,N_10636);
nand U11351 (N_11351,N_10667,N_10873);
or U11352 (N_11352,N_10872,N_10825);
nand U11353 (N_11353,N_10707,N_10919);
nor U11354 (N_11354,N_10970,N_10979);
and U11355 (N_11355,N_10574,N_10625);
nor U11356 (N_11356,N_10875,N_10969);
nor U11357 (N_11357,N_10809,N_10939);
nor U11358 (N_11358,N_10843,N_10955);
nand U11359 (N_11359,N_10967,N_10536);
nand U11360 (N_11360,N_10898,N_10593);
or U11361 (N_11361,N_10656,N_10977);
and U11362 (N_11362,N_10507,N_10554);
and U11363 (N_11363,N_10574,N_10705);
xor U11364 (N_11364,N_10877,N_10874);
nand U11365 (N_11365,N_10676,N_10956);
or U11366 (N_11366,N_10630,N_10883);
xor U11367 (N_11367,N_10985,N_10757);
nor U11368 (N_11368,N_10616,N_10818);
nor U11369 (N_11369,N_10975,N_10997);
xor U11370 (N_11370,N_10554,N_10521);
nor U11371 (N_11371,N_10836,N_10668);
or U11372 (N_11372,N_10901,N_10647);
or U11373 (N_11373,N_10774,N_10900);
and U11374 (N_11374,N_10802,N_10595);
nand U11375 (N_11375,N_10819,N_10587);
nand U11376 (N_11376,N_10615,N_10833);
and U11377 (N_11377,N_10660,N_10851);
nor U11378 (N_11378,N_10618,N_10875);
nand U11379 (N_11379,N_10757,N_10576);
or U11380 (N_11380,N_10707,N_10799);
and U11381 (N_11381,N_10805,N_10641);
xnor U11382 (N_11382,N_10713,N_10833);
and U11383 (N_11383,N_10693,N_10611);
and U11384 (N_11384,N_10928,N_10747);
nor U11385 (N_11385,N_10529,N_10753);
nor U11386 (N_11386,N_10584,N_10505);
nand U11387 (N_11387,N_10703,N_10612);
and U11388 (N_11388,N_10677,N_10801);
nand U11389 (N_11389,N_10728,N_10934);
or U11390 (N_11390,N_10748,N_10531);
and U11391 (N_11391,N_10574,N_10950);
nor U11392 (N_11392,N_10599,N_10664);
or U11393 (N_11393,N_10935,N_10957);
or U11394 (N_11394,N_10746,N_10882);
nor U11395 (N_11395,N_10513,N_10536);
xnor U11396 (N_11396,N_10952,N_10568);
nor U11397 (N_11397,N_10645,N_10765);
xnor U11398 (N_11398,N_10858,N_10568);
or U11399 (N_11399,N_10945,N_10909);
nand U11400 (N_11400,N_10988,N_10616);
or U11401 (N_11401,N_10801,N_10657);
xor U11402 (N_11402,N_10835,N_10697);
or U11403 (N_11403,N_10691,N_10667);
and U11404 (N_11404,N_10982,N_10990);
and U11405 (N_11405,N_10848,N_10963);
nor U11406 (N_11406,N_10660,N_10857);
nor U11407 (N_11407,N_10710,N_10608);
nand U11408 (N_11408,N_10584,N_10962);
and U11409 (N_11409,N_10646,N_10633);
nor U11410 (N_11410,N_10660,N_10582);
and U11411 (N_11411,N_10888,N_10768);
and U11412 (N_11412,N_10508,N_10826);
nand U11413 (N_11413,N_10612,N_10670);
nor U11414 (N_11414,N_10748,N_10609);
nand U11415 (N_11415,N_10713,N_10732);
nor U11416 (N_11416,N_10514,N_10945);
nor U11417 (N_11417,N_10809,N_10965);
or U11418 (N_11418,N_10907,N_10897);
or U11419 (N_11419,N_10608,N_10546);
nand U11420 (N_11420,N_10742,N_10668);
or U11421 (N_11421,N_10636,N_10959);
nand U11422 (N_11422,N_10699,N_10845);
and U11423 (N_11423,N_10744,N_10653);
and U11424 (N_11424,N_10715,N_10891);
nand U11425 (N_11425,N_10998,N_10779);
and U11426 (N_11426,N_10903,N_10610);
and U11427 (N_11427,N_10593,N_10554);
nand U11428 (N_11428,N_10586,N_10519);
or U11429 (N_11429,N_10729,N_10538);
nor U11430 (N_11430,N_10875,N_10616);
and U11431 (N_11431,N_10917,N_10954);
or U11432 (N_11432,N_10621,N_10592);
xnor U11433 (N_11433,N_10503,N_10798);
or U11434 (N_11434,N_10675,N_10941);
and U11435 (N_11435,N_10795,N_10885);
and U11436 (N_11436,N_10625,N_10872);
nor U11437 (N_11437,N_10969,N_10696);
and U11438 (N_11438,N_10658,N_10828);
nand U11439 (N_11439,N_10520,N_10923);
xor U11440 (N_11440,N_10922,N_10677);
nor U11441 (N_11441,N_10968,N_10841);
xor U11442 (N_11442,N_10774,N_10687);
nand U11443 (N_11443,N_10676,N_10611);
or U11444 (N_11444,N_10975,N_10569);
xor U11445 (N_11445,N_10970,N_10748);
nand U11446 (N_11446,N_10676,N_10961);
xor U11447 (N_11447,N_10611,N_10510);
nand U11448 (N_11448,N_10772,N_10618);
or U11449 (N_11449,N_10627,N_10902);
nor U11450 (N_11450,N_10916,N_10711);
and U11451 (N_11451,N_10968,N_10649);
and U11452 (N_11452,N_10680,N_10905);
nand U11453 (N_11453,N_10524,N_10542);
xor U11454 (N_11454,N_10946,N_10889);
and U11455 (N_11455,N_10580,N_10620);
and U11456 (N_11456,N_10960,N_10669);
or U11457 (N_11457,N_10813,N_10603);
nor U11458 (N_11458,N_10981,N_10919);
nand U11459 (N_11459,N_10919,N_10717);
xor U11460 (N_11460,N_10946,N_10973);
xnor U11461 (N_11461,N_10924,N_10668);
and U11462 (N_11462,N_10986,N_10951);
and U11463 (N_11463,N_10749,N_10707);
nand U11464 (N_11464,N_10980,N_10629);
nand U11465 (N_11465,N_10726,N_10893);
nand U11466 (N_11466,N_10742,N_10984);
and U11467 (N_11467,N_10555,N_10696);
and U11468 (N_11468,N_10828,N_10765);
nor U11469 (N_11469,N_10932,N_10934);
nor U11470 (N_11470,N_10976,N_10784);
nand U11471 (N_11471,N_10647,N_10827);
nand U11472 (N_11472,N_10968,N_10954);
and U11473 (N_11473,N_10516,N_10812);
or U11474 (N_11474,N_10550,N_10966);
or U11475 (N_11475,N_10592,N_10844);
and U11476 (N_11476,N_10609,N_10574);
nand U11477 (N_11477,N_10523,N_10899);
nor U11478 (N_11478,N_10822,N_10759);
or U11479 (N_11479,N_10794,N_10569);
nand U11480 (N_11480,N_10740,N_10668);
or U11481 (N_11481,N_10620,N_10551);
nor U11482 (N_11482,N_10750,N_10530);
and U11483 (N_11483,N_10921,N_10519);
nand U11484 (N_11484,N_10682,N_10536);
or U11485 (N_11485,N_10958,N_10892);
xnor U11486 (N_11486,N_10879,N_10644);
nand U11487 (N_11487,N_10582,N_10806);
and U11488 (N_11488,N_10506,N_10504);
nand U11489 (N_11489,N_10992,N_10950);
nand U11490 (N_11490,N_10795,N_10609);
and U11491 (N_11491,N_10865,N_10862);
and U11492 (N_11492,N_10605,N_10791);
nor U11493 (N_11493,N_10645,N_10874);
nor U11494 (N_11494,N_10569,N_10866);
and U11495 (N_11495,N_10557,N_10682);
xor U11496 (N_11496,N_10869,N_10506);
or U11497 (N_11497,N_10596,N_10615);
xor U11498 (N_11498,N_10581,N_10734);
nor U11499 (N_11499,N_10746,N_10536);
and U11500 (N_11500,N_11341,N_11217);
nand U11501 (N_11501,N_11134,N_11022);
or U11502 (N_11502,N_11192,N_11233);
xnor U11503 (N_11503,N_11422,N_11026);
nor U11504 (N_11504,N_11468,N_11411);
nor U11505 (N_11505,N_11149,N_11014);
and U11506 (N_11506,N_11486,N_11060);
nor U11507 (N_11507,N_11450,N_11360);
and U11508 (N_11508,N_11075,N_11056);
or U11509 (N_11509,N_11396,N_11320);
nor U11510 (N_11510,N_11105,N_11040);
nor U11511 (N_11511,N_11372,N_11123);
xor U11512 (N_11512,N_11065,N_11498);
or U11513 (N_11513,N_11374,N_11323);
nor U11514 (N_11514,N_11171,N_11034);
nand U11515 (N_11515,N_11475,N_11096);
nor U11516 (N_11516,N_11263,N_11283);
xor U11517 (N_11517,N_11470,N_11358);
xor U11518 (N_11518,N_11435,N_11172);
and U11519 (N_11519,N_11159,N_11241);
nand U11520 (N_11520,N_11010,N_11295);
or U11521 (N_11521,N_11209,N_11155);
or U11522 (N_11522,N_11478,N_11292);
nand U11523 (N_11523,N_11116,N_11080);
and U11524 (N_11524,N_11156,N_11385);
nor U11525 (N_11525,N_11113,N_11214);
and U11526 (N_11526,N_11011,N_11425);
and U11527 (N_11527,N_11184,N_11180);
or U11528 (N_11528,N_11273,N_11165);
and U11529 (N_11529,N_11313,N_11198);
nand U11530 (N_11530,N_11490,N_11030);
and U11531 (N_11531,N_11083,N_11294);
nand U11532 (N_11532,N_11025,N_11434);
or U11533 (N_11533,N_11104,N_11371);
and U11534 (N_11534,N_11079,N_11230);
nor U11535 (N_11535,N_11463,N_11117);
and U11536 (N_11536,N_11076,N_11272);
and U11537 (N_11537,N_11431,N_11467);
nor U11538 (N_11538,N_11074,N_11436);
xor U11539 (N_11539,N_11400,N_11329);
or U11540 (N_11540,N_11170,N_11349);
xor U11541 (N_11541,N_11328,N_11191);
xor U11542 (N_11542,N_11419,N_11195);
nand U11543 (N_11543,N_11148,N_11231);
or U11544 (N_11544,N_11046,N_11342);
nor U11545 (N_11545,N_11441,N_11461);
and U11546 (N_11546,N_11222,N_11049);
nor U11547 (N_11547,N_11078,N_11162);
or U11548 (N_11548,N_11340,N_11006);
and U11549 (N_11549,N_11359,N_11289);
or U11550 (N_11550,N_11160,N_11062);
and U11551 (N_11551,N_11377,N_11090);
and U11552 (N_11552,N_11388,N_11373);
nor U11553 (N_11553,N_11166,N_11050);
or U11554 (N_11554,N_11392,N_11316);
nand U11555 (N_11555,N_11041,N_11386);
xor U11556 (N_11556,N_11446,N_11364);
and U11557 (N_11557,N_11367,N_11311);
or U11558 (N_11558,N_11315,N_11399);
nor U11559 (N_11559,N_11382,N_11103);
nor U11560 (N_11560,N_11420,N_11137);
nand U11561 (N_11561,N_11319,N_11484);
nor U11562 (N_11562,N_11139,N_11335);
and U11563 (N_11563,N_11063,N_11228);
and U11564 (N_11564,N_11218,N_11179);
and U11565 (N_11565,N_11347,N_11406);
xnor U11566 (N_11566,N_11143,N_11205);
xnor U11567 (N_11567,N_11269,N_11442);
and U11568 (N_11568,N_11144,N_11314);
nand U11569 (N_11569,N_11380,N_11092);
and U11570 (N_11570,N_11458,N_11408);
nand U11571 (N_11571,N_11097,N_11176);
and U11572 (N_11572,N_11015,N_11309);
nor U11573 (N_11573,N_11476,N_11128);
or U11574 (N_11574,N_11194,N_11356);
or U11575 (N_11575,N_11477,N_11394);
nand U11576 (N_11576,N_11448,N_11276);
nor U11577 (N_11577,N_11208,N_11426);
nor U11578 (N_11578,N_11039,N_11136);
and U11579 (N_11579,N_11338,N_11460);
nor U11580 (N_11580,N_11256,N_11120);
and U11581 (N_11581,N_11462,N_11277);
nor U11582 (N_11582,N_11317,N_11278);
nand U11583 (N_11583,N_11140,N_11099);
and U11584 (N_11584,N_11413,N_11142);
nand U11585 (N_11585,N_11138,N_11037);
or U11586 (N_11586,N_11302,N_11032);
or U11587 (N_11587,N_11479,N_11398);
and U11588 (N_11588,N_11487,N_11250);
and U11589 (N_11589,N_11405,N_11107);
xor U11590 (N_11590,N_11109,N_11387);
or U11591 (N_11591,N_11196,N_11084);
nor U11592 (N_11592,N_11404,N_11370);
and U11593 (N_11593,N_11366,N_11121);
or U11594 (N_11594,N_11471,N_11178);
nand U11595 (N_11595,N_11438,N_11293);
nor U11596 (N_11596,N_11362,N_11281);
and U11597 (N_11597,N_11058,N_11001);
nor U11598 (N_11598,N_11326,N_11238);
nor U11599 (N_11599,N_11457,N_11251);
or U11600 (N_11600,N_11332,N_11239);
or U11601 (N_11601,N_11031,N_11213);
and U11602 (N_11602,N_11449,N_11101);
nor U11603 (N_11603,N_11012,N_11375);
or U11604 (N_11604,N_11211,N_11111);
nand U11605 (N_11605,N_11363,N_11181);
nand U11606 (N_11606,N_11355,N_11150);
and U11607 (N_11607,N_11072,N_11053);
or U11608 (N_11608,N_11445,N_11403);
nor U11609 (N_11609,N_11091,N_11082);
or U11610 (N_11610,N_11029,N_11282);
nand U11611 (N_11611,N_11287,N_11253);
nand U11612 (N_11612,N_11390,N_11352);
nor U11613 (N_11613,N_11068,N_11330);
or U11614 (N_11614,N_11182,N_11093);
or U11615 (N_11615,N_11303,N_11249);
and U11616 (N_11616,N_11237,N_11197);
xnor U11617 (N_11617,N_11254,N_11496);
nor U11618 (N_11618,N_11019,N_11110);
nand U11619 (N_11619,N_11301,N_11207);
nand U11620 (N_11620,N_11126,N_11094);
nand U11621 (N_11621,N_11260,N_11480);
nor U11622 (N_11622,N_11004,N_11409);
xnor U11623 (N_11623,N_11225,N_11410);
xnor U11624 (N_11624,N_11221,N_11059);
xnor U11625 (N_11625,N_11146,N_11378);
or U11626 (N_11626,N_11005,N_11051);
xnor U11627 (N_11627,N_11236,N_11061);
and U11628 (N_11628,N_11047,N_11333);
and U11629 (N_11629,N_11334,N_11152);
and U11630 (N_11630,N_11044,N_11033);
nor U11631 (N_11631,N_11354,N_11379);
and U11632 (N_11632,N_11186,N_11299);
nor U11633 (N_11633,N_11023,N_11415);
xor U11634 (N_11634,N_11244,N_11325);
nand U11635 (N_11635,N_11455,N_11492);
nand U11636 (N_11636,N_11202,N_11451);
nand U11637 (N_11637,N_11234,N_11259);
and U11638 (N_11638,N_11008,N_11397);
nand U11639 (N_11639,N_11173,N_11433);
xor U11640 (N_11640,N_11391,N_11161);
nor U11641 (N_11641,N_11108,N_11339);
and U11642 (N_11642,N_11444,N_11028);
and U11643 (N_11643,N_11145,N_11350);
and U11644 (N_11644,N_11306,N_11361);
nor U11645 (N_11645,N_11465,N_11077);
and U11646 (N_11646,N_11147,N_11066);
nand U11647 (N_11647,N_11285,N_11428);
nand U11648 (N_11648,N_11045,N_11100);
or U11649 (N_11649,N_11255,N_11418);
or U11650 (N_11650,N_11157,N_11190);
nor U11651 (N_11651,N_11485,N_11219);
and U11652 (N_11652,N_11112,N_11308);
nor U11653 (N_11653,N_11095,N_11336);
nand U11654 (N_11654,N_11497,N_11327);
and U11655 (N_11655,N_11067,N_11412);
xnor U11656 (N_11656,N_11464,N_11232);
nor U11657 (N_11657,N_11235,N_11473);
nor U11658 (N_11658,N_11312,N_11102);
nand U11659 (N_11659,N_11003,N_11261);
and U11660 (N_11660,N_11027,N_11452);
nor U11661 (N_11661,N_11383,N_11226);
and U11662 (N_11662,N_11401,N_11018);
and U11663 (N_11663,N_11424,N_11453);
and U11664 (N_11664,N_11267,N_11245);
and U11665 (N_11665,N_11296,N_11286);
and U11666 (N_11666,N_11118,N_11384);
or U11667 (N_11667,N_11279,N_11472);
nand U11668 (N_11668,N_11017,N_11215);
or U11669 (N_11669,N_11071,N_11429);
xor U11670 (N_11670,N_11073,N_11151);
nand U11671 (N_11671,N_11224,N_11439);
nor U11672 (N_11672,N_11106,N_11430);
and U11673 (N_11673,N_11290,N_11368);
nand U11674 (N_11674,N_11020,N_11081);
and U11675 (N_11675,N_11085,N_11130);
nand U11676 (N_11676,N_11013,N_11203);
and U11677 (N_11677,N_11357,N_11036);
nand U11678 (N_11678,N_11199,N_11459);
nand U11679 (N_11679,N_11216,N_11432);
and U11680 (N_11680,N_11125,N_11177);
and U11681 (N_11681,N_11242,N_11114);
xnor U11682 (N_11682,N_11483,N_11491);
nand U11683 (N_11683,N_11495,N_11115);
xor U11684 (N_11684,N_11185,N_11164);
nor U11685 (N_11685,N_11423,N_11174);
nand U11686 (N_11686,N_11275,N_11042);
nand U11687 (N_11687,N_11069,N_11421);
nand U11688 (N_11688,N_11169,N_11009);
and U11689 (N_11689,N_11129,N_11322);
or U11690 (N_11690,N_11206,N_11007);
nand U11691 (N_11691,N_11381,N_11324);
xnor U11692 (N_11692,N_11456,N_11482);
nand U11693 (N_11693,N_11154,N_11098);
nand U11694 (N_11694,N_11141,N_11346);
nand U11695 (N_11695,N_11353,N_11124);
nand U11696 (N_11696,N_11167,N_11437);
xnor U11697 (N_11697,N_11133,N_11135);
nor U11698 (N_11698,N_11201,N_11300);
and U11699 (N_11699,N_11447,N_11048);
xor U11700 (N_11700,N_11344,N_11493);
and U11701 (N_11701,N_11297,N_11489);
and U11702 (N_11702,N_11305,N_11229);
or U11703 (N_11703,N_11021,N_11168);
nand U11704 (N_11704,N_11089,N_11481);
nor U11705 (N_11705,N_11365,N_11054);
or U11706 (N_11706,N_11488,N_11038);
or U11707 (N_11707,N_11345,N_11220);
and U11708 (N_11708,N_11088,N_11466);
or U11709 (N_11709,N_11270,N_11331);
and U11710 (N_11710,N_11227,N_11402);
and U11711 (N_11711,N_11262,N_11271);
and U11712 (N_11712,N_11369,N_11087);
and U11713 (N_11713,N_11064,N_11193);
nand U11714 (N_11714,N_11247,N_11189);
and U11715 (N_11715,N_11127,N_11240);
and U11716 (N_11716,N_11389,N_11416);
or U11717 (N_11717,N_11298,N_11210);
xnor U11718 (N_11718,N_11187,N_11417);
or U11719 (N_11719,N_11153,N_11284);
and U11720 (N_11720,N_11122,N_11307);
and U11721 (N_11721,N_11223,N_11348);
nand U11722 (N_11722,N_11000,N_11016);
nor U11723 (N_11723,N_11035,N_11343);
and U11724 (N_11724,N_11070,N_11002);
or U11725 (N_11725,N_11337,N_11119);
nand U11726 (N_11726,N_11183,N_11393);
nor U11727 (N_11727,N_11057,N_11440);
and U11728 (N_11728,N_11469,N_11248);
and U11729 (N_11729,N_11266,N_11132);
or U11730 (N_11730,N_11055,N_11246);
nand U11731 (N_11731,N_11376,N_11280);
xor U11732 (N_11732,N_11257,N_11321);
or U11733 (N_11733,N_11395,N_11158);
nor U11734 (N_11734,N_11274,N_11443);
nor U11735 (N_11735,N_11204,N_11264);
nand U11736 (N_11736,N_11310,N_11494);
and U11737 (N_11737,N_11052,N_11318);
nand U11738 (N_11738,N_11407,N_11258);
or U11739 (N_11739,N_11288,N_11454);
or U11740 (N_11740,N_11265,N_11304);
nor U11741 (N_11741,N_11427,N_11131);
nand U11742 (N_11742,N_11043,N_11351);
nand U11743 (N_11743,N_11291,N_11243);
or U11744 (N_11744,N_11499,N_11474);
or U11745 (N_11745,N_11252,N_11200);
nor U11746 (N_11746,N_11175,N_11268);
nor U11747 (N_11747,N_11212,N_11414);
nand U11748 (N_11748,N_11086,N_11188);
or U11749 (N_11749,N_11163,N_11024);
nor U11750 (N_11750,N_11464,N_11419);
or U11751 (N_11751,N_11035,N_11246);
or U11752 (N_11752,N_11403,N_11418);
or U11753 (N_11753,N_11140,N_11247);
nor U11754 (N_11754,N_11066,N_11371);
or U11755 (N_11755,N_11266,N_11211);
nor U11756 (N_11756,N_11416,N_11210);
nand U11757 (N_11757,N_11354,N_11453);
or U11758 (N_11758,N_11370,N_11068);
xnor U11759 (N_11759,N_11248,N_11014);
xnor U11760 (N_11760,N_11365,N_11237);
and U11761 (N_11761,N_11333,N_11220);
and U11762 (N_11762,N_11155,N_11110);
nand U11763 (N_11763,N_11233,N_11097);
and U11764 (N_11764,N_11318,N_11195);
nand U11765 (N_11765,N_11126,N_11230);
xnor U11766 (N_11766,N_11061,N_11112);
nor U11767 (N_11767,N_11115,N_11467);
or U11768 (N_11768,N_11428,N_11331);
or U11769 (N_11769,N_11418,N_11484);
nand U11770 (N_11770,N_11179,N_11120);
or U11771 (N_11771,N_11312,N_11430);
and U11772 (N_11772,N_11014,N_11302);
nand U11773 (N_11773,N_11351,N_11465);
or U11774 (N_11774,N_11336,N_11349);
or U11775 (N_11775,N_11323,N_11183);
nand U11776 (N_11776,N_11490,N_11463);
nand U11777 (N_11777,N_11263,N_11308);
nor U11778 (N_11778,N_11428,N_11163);
nor U11779 (N_11779,N_11150,N_11179);
nand U11780 (N_11780,N_11077,N_11394);
or U11781 (N_11781,N_11226,N_11025);
and U11782 (N_11782,N_11417,N_11256);
or U11783 (N_11783,N_11136,N_11258);
and U11784 (N_11784,N_11465,N_11386);
nor U11785 (N_11785,N_11027,N_11182);
xnor U11786 (N_11786,N_11372,N_11386);
nor U11787 (N_11787,N_11085,N_11499);
or U11788 (N_11788,N_11295,N_11382);
xor U11789 (N_11789,N_11040,N_11176);
nor U11790 (N_11790,N_11157,N_11346);
nand U11791 (N_11791,N_11039,N_11057);
or U11792 (N_11792,N_11406,N_11455);
nor U11793 (N_11793,N_11411,N_11313);
nor U11794 (N_11794,N_11482,N_11072);
nand U11795 (N_11795,N_11028,N_11154);
nand U11796 (N_11796,N_11217,N_11058);
nand U11797 (N_11797,N_11329,N_11252);
nand U11798 (N_11798,N_11075,N_11445);
and U11799 (N_11799,N_11232,N_11363);
nor U11800 (N_11800,N_11388,N_11113);
or U11801 (N_11801,N_11027,N_11358);
and U11802 (N_11802,N_11067,N_11478);
nand U11803 (N_11803,N_11136,N_11486);
nor U11804 (N_11804,N_11054,N_11000);
nand U11805 (N_11805,N_11317,N_11445);
nand U11806 (N_11806,N_11492,N_11434);
and U11807 (N_11807,N_11101,N_11302);
xor U11808 (N_11808,N_11320,N_11257);
and U11809 (N_11809,N_11033,N_11102);
and U11810 (N_11810,N_11210,N_11455);
nand U11811 (N_11811,N_11346,N_11382);
or U11812 (N_11812,N_11313,N_11213);
nand U11813 (N_11813,N_11448,N_11457);
nand U11814 (N_11814,N_11276,N_11489);
xor U11815 (N_11815,N_11002,N_11498);
or U11816 (N_11816,N_11340,N_11096);
and U11817 (N_11817,N_11480,N_11376);
nor U11818 (N_11818,N_11077,N_11416);
nor U11819 (N_11819,N_11283,N_11082);
and U11820 (N_11820,N_11089,N_11451);
nand U11821 (N_11821,N_11490,N_11248);
or U11822 (N_11822,N_11434,N_11258);
nor U11823 (N_11823,N_11061,N_11200);
or U11824 (N_11824,N_11129,N_11133);
and U11825 (N_11825,N_11309,N_11294);
and U11826 (N_11826,N_11492,N_11488);
nand U11827 (N_11827,N_11335,N_11237);
and U11828 (N_11828,N_11270,N_11076);
and U11829 (N_11829,N_11171,N_11120);
nand U11830 (N_11830,N_11066,N_11133);
xnor U11831 (N_11831,N_11445,N_11216);
nor U11832 (N_11832,N_11235,N_11049);
nor U11833 (N_11833,N_11392,N_11478);
and U11834 (N_11834,N_11257,N_11389);
nand U11835 (N_11835,N_11113,N_11019);
xor U11836 (N_11836,N_11161,N_11002);
nand U11837 (N_11837,N_11004,N_11131);
or U11838 (N_11838,N_11188,N_11384);
xor U11839 (N_11839,N_11050,N_11192);
and U11840 (N_11840,N_11156,N_11242);
and U11841 (N_11841,N_11270,N_11151);
nor U11842 (N_11842,N_11420,N_11302);
or U11843 (N_11843,N_11143,N_11237);
xnor U11844 (N_11844,N_11438,N_11367);
nand U11845 (N_11845,N_11389,N_11273);
or U11846 (N_11846,N_11302,N_11308);
nor U11847 (N_11847,N_11086,N_11295);
or U11848 (N_11848,N_11288,N_11134);
nor U11849 (N_11849,N_11494,N_11248);
xor U11850 (N_11850,N_11179,N_11450);
xnor U11851 (N_11851,N_11113,N_11325);
and U11852 (N_11852,N_11245,N_11214);
and U11853 (N_11853,N_11421,N_11144);
nor U11854 (N_11854,N_11233,N_11209);
nand U11855 (N_11855,N_11042,N_11170);
nor U11856 (N_11856,N_11272,N_11139);
or U11857 (N_11857,N_11306,N_11215);
or U11858 (N_11858,N_11141,N_11296);
nand U11859 (N_11859,N_11293,N_11174);
nand U11860 (N_11860,N_11440,N_11050);
nor U11861 (N_11861,N_11227,N_11094);
and U11862 (N_11862,N_11416,N_11206);
and U11863 (N_11863,N_11455,N_11247);
or U11864 (N_11864,N_11306,N_11496);
or U11865 (N_11865,N_11166,N_11099);
xor U11866 (N_11866,N_11051,N_11266);
or U11867 (N_11867,N_11123,N_11244);
or U11868 (N_11868,N_11188,N_11228);
nor U11869 (N_11869,N_11080,N_11197);
nand U11870 (N_11870,N_11128,N_11277);
and U11871 (N_11871,N_11232,N_11372);
nand U11872 (N_11872,N_11239,N_11082);
xnor U11873 (N_11873,N_11026,N_11404);
nand U11874 (N_11874,N_11076,N_11155);
nor U11875 (N_11875,N_11224,N_11388);
xor U11876 (N_11876,N_11206,N_11303);
and U11877 (N_11877,N_11047,N_11135);
nand U11878 (N_11878,N_11110,N_11325);
nor U11879 (N_11879,N_11239,N_11039);
and U11880 (N_11880,N_11380,N_11483);
nand U11881 (N_11881,N_11473,N_11022);
and U11882 (N_11882,N_11046,N_11471);
and U11883 (N_11883,N_11304,N_11498);
or U11884 (N_11884,N_11425,N_11488);
and U11885 (N_11885,N_11408,N_11184);
and U11886 (N_11886,N_11262,N_11291);
nor U11887 (N_11887,N_11292,N_11015);
nand U11888 (N_11888,N_11376,N_11195);
or U11889 (N_11889,N_11012,N_11276);
and U11890 (N_11890,N_11472,N_11280);
xor U11891 (N_11891,N_11002,N_11244);
or U11892 (N_11892,N_11371,N_11033);
or U11893 (N_11893,N_11035,N_11445);
nand U11894 (N_11894,N_11327,N_11464);
nor U11895 (N_11895,N_11137,N_11063);
xnor U11896 (N_11896,N_11234,N_11427);
or U11897 (N_11897,N_11470,N_11220);
nor U11898 (N_11898,N_11499,N_11058);
nor U11899 (N_11899,N_11388,N_11147);
or U11900 (N_11900,N_11491,N_11286);
or U11901 (N_11901,N_11022,N_11140);
or U11902 (N_11902,N_11207,N_11124);
nor U11903 (N_11903,N_11139,N_11365);
xnor U11904 (N_11904,N_11210,N_11321);
nor U11905 (N_11905,N_11045,N_11231);
or U11906 (N_11906,N_11113,N_11184);
nor U11907 (N_11907,N_11122,N_11322);
nor U11908 (N_11908,N_11469,N_11368);
and U11909 (N_11909,N_11453,N_11438);
nor U11910 (N_11910,N_11054,N_11131);
nor U11911 (N_11911,N_11461,N_11446);
nor U11912 (N_11912,N_11330,N_11308);
nand U11913 (N_11913,N_11236,N_11093);
nor U11914 (N_11914,N_11367,N_11074);
nand U11915 (N_11915,N_11148,N_11373);
or U11916 (N_11916,N_11276,N_11210);
or U11917 (N_11917,N_11188,N_11455);
xnor U11918 (N_11918,N_11206,N_11194);
nor U11919 (N_11919,N_11213,N_11062);
or U11920 (N_11920,N_11417,N_11137);
or U11921 (N_11921,N_11358,N_11029);
nand U11922 (N_11922,N_11456,N_11037);
and U11923 (N_11923,N_11245,N_11394);
nand U11924 (N_11924,N_11209,N_11361);
and U11925 (N_11925,N_11164,N_11445);
and U11926 (N_11926,N_11189,N_11391);
nand U11927 (N_11927,N_11331,N_11351);
nand U11928 (N_11928,N_11363,N_11142);
nand U11929 (N_11929,N_11252,N_11237);
xor U11930 (N_11930,N_11073,N_11497);
nor U11931 (N_11931,N_11073,N_11400);
nand U11932 (N_11932,N_11320,N_11280);
nand U11933 (N_11933,N_11282,N_11043);
nand U11934 (N_11934,N_11169,N_11016);
nor U11935 (N_11935,N_11083,N_11494);
or U11936 (N_11936,N_11426,N_11119);
or U11937 (N_11937,N_11030,N_11405);
nand U11938 (N_11938,N_11106,N_11181);
nand U11939 (N_11939,N_11124,N_11364);
xor U11940 (N_11940,N_11218,N_11192);
nor U11941 (N_11941,N_11191,N_11318);
and U11942 (N_11942,N_11322,N_11029);
or U11943 (N_11943,N_11031,N_11101);
or U11944 (N_11944,N_11156,N_11205);
or U11945 (N_11945,N_11212,N_11388);
and U11946 (N_11946,N_11259,N_11176);
and U11947 (N_11947,N_11344,N_11282);
and U11948 (N_11948,N_11374,N_11411);
nor U11949 (N_11949,N_11107,N_11149);
or U11950 (N_11950,N_11191,N_11177);
and U11951 (N_11951,N_11480,N_11354);
nor U11952 (N_11952,N_11349,N_11175);
xnor U11953 (N_11953,N_11449,N_11334);
and U11954 (N_11954,N_11418,N_11440);
nor U11955 (N_11955,N_11386,N_11188);
and U11956 (N_11956,N_11426,N_11043);
xnor U11957 (N_11957,N_11226,N_11242);
and U11958 (N_11958,N_11376,N_11401);
or U11959 (N_11959,N_11491,N_11369);
xnor U11960 (N_11960,N_11182,N_11116);
nand U11961 (N_11961,N_11168,N_11087);
and U11962 (N_11962,N_11439,N_11377);
nor U11963 (N_11963,N_11203,N_11070);
and U11964 (N_11964,N_11431,N_11432);
or U11965 (N_11965,N_11264,N_11352);
xor U11966 (N_11966,N_11085,N_11334);
or U11967 (N_11967,N_11304,N_11475);
nand U11968 (N_11968,N_11422,N_11389);
or U11969 (N_11969,N_11440,N_11151);
nor U11970 (N_11970,N_11258,N_11155);
xnor U11971 (N_11971,N_11095,N_11492);
xnor U11972 (N_11972,N_11086,N_11423);
xor U11973 (N_11973,N_11164,N_11491);
nand U11974 (N_11974,N_11488,N_11415);
nor U11975 (N_11975,N_11364,N_11309);
nand U11976 (N_11976,N_11420,N_11177);
or U11977 (N_11977,N_11360,N_11393);
or U11978 (N_11978,N_11262,N_11171);
xnor U11979 (N_11979,N_11004,N_11143);
nor U11980 (N_11980,N_11066,N_11071);
or U11981 (N_11981,N_11111,N_11386);
or U11982 (N_11982,N_11298,N_11126);
and U11983 (N_11983,N_11278,N_11087);
nor U11984 (N_11984,N_11217,N_11380);
xnor U11985 (N_11985,N_11109,N_11191);
nor U11986 (N_11986,N_11376,N_11083);
nor U11987 (N_11987,N_11173,N_11003);
nand U11988 (N_11988,N_11039,N_11263);
and U11989 (N_11989,N_11014,N_11112);
or U11990 (N_11990,N_11460,N_11456);
nor U11991 (N_11991,N_11114,N_11375);
or U11992 (N_11992,N_11229,N_11338);
and U11993 (N_11993,N_11141,N_11270);
or U11994 (N_11994,N_11140,N_11137);
nor U11995 (N_11995,N_11490,N_11185);
nor U11996 (N_11996,N_11344,N_11399);
or U11997 (N_11997,N_11094,N_11080);
and U11998 (N_11998,N_11150,N_11433);
xor U11999 (N_11999,N_11467,N_11311);
and U12000 (N_12000,N_11605,N_11717);
or U12001 (N_12001,N_11847,N_11972);
nand U12002 (N_12002,N_11640,N_11657);
and U12003 (N_12003,N_11689,N_11625);
nor U12004 (N_12004,N_11834,N_11587);
xnor U12005 (N_12005,N_11726,N_11903);
nor U12006 (N_12006,N_11861,N_11886);
and U12007 (N_12007,N_11993,N_11788);
nand U12008 (N_12008,N_11533,N_11629);
nor U12009 (N_12009,N_11645,N_11994);
nor U12010 (N_12010,N_11518,N_11647);
xor U12011 (N_12011,N_11781,N_11548);
xnor U12012 (N_12012,N_11929,N_11749);
nand U12013 (N_12013,N_11792,N_11732);
and U12014 (N_12014,N_11948,N_11571);
or U12015 (N_12015,N_11527,N_11983);
nand U12016 (N_12016,N_11683,N_11826);
and U12017 (N_12017,N_11727,N_11711);
nand U12018 (N_12018,N_11900,N_11980);
nand U12019 (N_12019,N_11982,N_11679);
and U12020 (N_12020,N_11573,N_11901);
or U12021 (N_12021,N_11643,N_11989);
nor U12022 (N_12022,N_11752,N_11957);
nand U12023 (N_12023,N_11654,N_11878);
nand U12024 (N_12024,N_11646,N_11699);
nor U12025 (N_12025,N_11927,N_11707);
nand U12026 (N_12026,N_11672,N_11904);
nor U12027 (N_12027,N_11695,N_11822);
and U12028 (N_12028,N_11636,N_11537);
nor U12029 (N_12029,N_11873,N_11540);
or U12030 (N_12030,N_11738,N_11649);
nor U12031 (N_12031,N_11524,N_11608);
xor U12032 (N_12032,N_11794,N_11896);
and U12033 (N_12033,N_11568,N_11569);
and U12034 (N_12034,N_11913,N_11741);
nand U12035 (N_12035,N_11889,N_11668);
nor U12036 (N_12036,N_11682,N_11962);
and U12037 (N_12037,N_11611,N_11633);
and U12038 (N_12038,N_11631,N_11714);
or U12039 (N_12039,N_11501,N_11881);
nor U12040 (N_12040,N_11566,N_11539);
nand U12041 (N_12041,N_11620,N_11733);
nand U12042 (N_12042,N_11685,N_11941);
and U12043 (N_12043,N_11502,N_11567);
nand U12044 (N_12044,N_11536,N_11688);
nor U12045 (N_12045,N_11856,N_11940);
xnor U12046 (N_12046,N_11543,N_11520);
nor U12047 (N_12047,N_11867,N_11894);
and U12048 (N_12048,N_11858,N_11996);
nand U12049 (N_12049,N_11746,N_11791);
nand U12050 (N_12050,N_11849,N_11736);
and U12051 (N_12051,N_11810,N_11598);
or U12052 (N_12052,N_11594,N_11698);
nand U12053 (N_12053,N_11825,N_11635);
and U12054 (N_12054,N_11658,N_11584);
and U12055 (N_12055,N_11512,N_11556);
and U12056 (N_12056,N_11574,N_11593);
nand U12057 (N_12057,N_11776,N_11987);
nand U12058 (N_12058,N_11868,N_11859);
nor U12059 (N_12059,N_11938,N_11802);
and U12060 (N_12060,N_11945,N_11525);
or U12061 (N_12061,N_11848,N_11846);
nand U12062 (N_12062,N_11747,N_11554);
or U12063 (N_12063,N_11837,N_11534);
xnor U12064 (N_12064,N_11780,N_11514);
nor U12065 (N_12065,N_11552,N_11515);
nor U12066 (N_12066,N_11816,N_11753);
nand U12067 (N_12067,N_11844,N_11511);
and U12068 (N_12068,N_11519,N_11952);
xnor U12069 (N_12069,N_11935,N_11710);
nor U12070 (N_12070,N_11516,N_11558);
and U12071 (N_12071,N_11866,N_11796);
nand U12072 (N_12072,N_11882,N_11731);
nand U12073 (N_12073,N_11914,N_11995);
nor U12074 (N_12074,N_11509,N_11755);
nand U12075 (N_12075,N_11925,N_11529);
nand U12076 (N_12076,N_11665,N_11966);
and U12077 (N_12077,N_11544,N_11575);
and U12078 (N_12078,N_11977,N_11662);
and U12079 (N_12079,N_11988,N_11637);
nor U12080 (N_12080,N_11729,N_11870);
and U12081 (N_12081,N_11939,N_11691);
nor U12082 (N_12082,N_11703,N_11949);
or U12083 (N_12083,N_11853,N_11845);
or U12084 (N_12084,N_11559,N_11560);
nor U12085 (N_12085,N_11902,N_11852);
xor U12086 (N_12086,N_11545,N_11863);
or U12087 (N_12087,N_11652,N_11697);
nor U12088 (N_12088,N_11804,N_11801);
or U12089 (N_12089,N_11706,N_11911);
or U12090 (N_12090,N_11924,N_11542);
and U12091 (N_12091,N_11674,N_11807);
or U12092 (N_12092,N_11581,N_11784);
or U12093 (N_12093,N_11819,N_11622);
nand U12094 (N_12094,N_11775,N_11772);
nand U12095 (N_12095,N_11920,N_11538);
and U12096 (N_12096,N_11626,N_11716);
nor U12097 (N_12097,N_11954,N_11670);
or U12098 (N_12098,N_11678,N_11898);
and U12099 (N_12099,N_11639,N_11730);
nand U12100 (N_12100,N_11609,N_11553);
nor U12101 (N_12101,N_11708,N_11592);
nor U12102 (N_12102,N_11963,N_11618);
nand U12103 (N_12103,N_11958,N_11748);
and U12104 (N_12104,N_11992,N_11743);
nand U12105 (N_12105,N_11589,N_11523);
nand U12106 (N_12106,N_11661,N_11500);
or U12107 (N_12107,N_11583,N_11890);
and U12108 (N_12108,N_11923,N_11719);
nand U12109 (N_12109,N_11803,N_11532);
xnor U12110 (N_12110,N_11517,N_11813);
nor U12111 (N_12111,N_11969,N_11561);
nand U12112 (N_12112,N_11831,N_11506);
nor U12113 (N_12113,N_11709,N_11968);
and U12114 (N_12114,N_11758,N_11754);
and U12115 (N_12115,N_11756,N_11806);
xor U12116 (N_12116,N_11829,N_11999);
or U12117 (N_12117,N_11768,N_11528);
nand U12118 (N_12118,N_11812,N_11634);
and U12119 (N_12119,N_11943,N_11879);
and U12120 (N_12120,N_11942,N_11783);
and U12121 (N_12121,N_11503,N_11586);
nand U12122 (N_12122,N_11650,N_11880);
nand U12123 (N_12123,N_11641,N_11808);
or U12124 (N_12124,N_11744,N_11971);
and U12125 (N_12125,N_11786,N_11951);
nor U12126 (N_12126,N_11693,N_11839);
nor U12127 (N_12127,N_11505,N_11814);
and U12128 (N_12128,N_11888,N_11700);
xnor U12129 (N_12129,N_11681,N_11600);
or U12130 (N_12130,N_11734,N_11843);
nor U12131 (N_12131,N_11774,N_11793);
nand U12132 (N_12132,N_11976,N_11887);
nand U12133 (N_12133,N_11818,N_11891);
or U12134 (N_12134,N_11798,N_11603);
nand U12135 (N_12135,N_11615,N_11895);
nor U12136 (N_12136,N_11919,N_11797);
nor U12137 (N_12137,N_11964,N_11671);
nor U12138 (N_12138,N_11928,N_11563);
nor U12139 (N_12139,N_11875,N_11860);
or U12140 (N_12140,N_11884,N_11953);
nor U12141 (N_12141,N_11740,N_11735);
nand U12142 (N_12142,N_11667,N_11893);
xor U12143 (N_12143,N_11701,N_11908);
nand U12144 (N_12144,N_11659,N_11677);
nor U12145 (N_12145,N_11690,N_11918);
and U12146 (N_12146,N_11530,N_11613);
and U12147 (N_12147,N_11765,N_11759);
or U12148 (N_12148,N_11842,N_11916);
nor U12149 (N_12149,N_11504,N_11767);
xor U12150 (N_12150,N_11850,N_11909);
and U12151 (N_12151,N_11771,N_11551);
nor U12152 (N_12152,N_11607,N_11612);
or U12153 (N_12153,N_11686,N_11932);
nor U12154 (N_12154,N_11604,N_11946);
nand U12155 (N_12155,N_11931,N_11974);
xnor U12156 (N_12156,N_11648,N_11624);
nor U12157 (N_12157,N_11936,N_11838);
nand U12158 (N_12158,N_11621,N_11669);
and U12159 (N_12159,N_11811,N_11751);
and U12160 (N_12160,N_11915,N_11981);
nand U12161 (N_12161,N_11800,N_11694);
or U12162 (N_12162,N_11926,N_11725);
or U12163 (N_12163,N_11809,N_11617);
or U12164 (N_12164,N_11950,N_11777);
xor U12165 (N_12165,N_11984,N_11773);
nand U12166 (N_12166,N_11864,N_11597);
and U12167 (N_12167,N_11585,N_11795);
or U12168 (N_12168,N_11912,N_11778);
and U12169 (N_12169,N_11985,N_11599);
or U12170 (N_12170,N_11578,N_11959);
or U12171 (N_12171,N_11970,N_11750);
nand U12172 (N_12172,N_11821,N_11872);
or U12173 (N_12173,N_11610,N_11947);
xor U12174 (N_12174,N_11590,N_11728);
nor U12175 (N_12175,N_11680,N_11905);
nor U12176 (N_12176,N_11664,N_11978);
nor U12177 (N_12177,N_11854,N_11836);
nand U12178 (N_12178,N_11865,N_11785);
nor U12179 (N_12179,N_11564,N_11973);
nand U12180 (N_12180,N_11975,N_11840);
and U12181 (N_12181,N_11656,N_11582);
nand U12182 (N_12182,N_11990,N_11546);
and U12183 (N_12183,N_11715,N_11522);
and U12184 (N_12184,N_11883,N_11828);
nand U12185 (N_12185,N_11991,N_11614);
nand U12186 (N_12186,N_11820,N_11874);
and U12187 (N_12187,N_11830,N_11997);
and U12188 (N_12188,N_11550,N_11742);
nor U12189 (N_12189,N_11580,N_11787);
nand U12190 (N_12190,N_11565,N_11857);
xnor U12191 (N_12191,N_11722,N_11760);
and U12192 (N_12192,N_11570,N_11979);
and U12193 (N_12193,N_11702,N_11547);
and U12194 (N_12194,N_11906,N_11944);
and U12195 (N_12195,N_11630,N_11644);
or U12196 (N_12196,N_11696,N_11956);
nor U12197 (N_12197,N_11934,N_11892);
and U12198 (N_12198,N_11718,N_11531);
or U12199 (N_12199,N_11619,N_11724);
or U12200 (N_12200,N_11799,N_11805);
nor U12201 (N_12201,N_11562,N_11965);
and U12202 (N_12202,N_11745,N_11782);
or U12203 (N_12203,N_11595,N_11660);
or U12204 (N_12204,N_11832,N_11541);
and U12205 (N_12205,N_11922,N_11930);
nand U12206 (N_12206,N_11897,N_11507);
nor U12207 (N_12207,N_11576,N_11655);
nand U12208 (N_12208,N_11663,N_11642);
and U12209 (N_12209,N_11602,N_11549);
xnor U12210 (N_12210,N_11723,N_11871);
nand U12211 (N_12211,N_11521,N_11967);
nor U12212 (N_12212,N_11998,N_11651);
and U12213 (N_12213,N_11855,N_11579);
or U12214 (N_12214,N_11557,N_11508);
nor U12215 (N_12215,N_11627,N_11596);
or U12216 (N_12216,N_11713,N_11591);
nand U12217 (N_12217,N_11632,N_11721);
nand U12218 (N_12218,N_11986,N_11769);
xor U12219 (N_12219,N_11705,N_11789);
or U12220 (N_12220,N_11790,N_11666);
nor U12221 (N_12221,N_11510,N_11577);
nand U12222 (N_12222,N_11739,N_11910);
nor U12223 (N_12223,N_11638,N_11763);
or U12224 (N_12224,N_11766,N_11676);
nor U12225 (N_12225,N_11817,N_11684);
and U12226 (N_12226,N_11779,N_11606);
and U12227 (N_12227,N_11628,N_11572);
and U12228 (N_12228,N_11555,N_11653);
or U12229 (N_12229,N_11757,N_11827);
and U12230 (N_12230,N_11762,N_11526);
and U12231 (N_12231,N_11824,N_11835);
xnor U12232 (N_12232,N_11960,N_11933);
and U12233 (N_12233,N_11877,N_11961);
nand U12234 (N_12234,N_11673,N_11841);
or U12235 (N_12235,N_11917,N_11535);
nand U12236 (N_12236,N_11869,N_11588);
nand U12237 (N_12237,N_11761,N_11823);
and U12238 (N_12238,N_11955,N_11770);
and U12239 (N_12239,N_11899,N_11712);
nand U12240 (N_12240,N_11737,N_11876);
xnor U12241 (N_12241,N_11937,N_11513);
and U12242 (N_12242,N_11623,N_11851);
nor U12243 (N_12243,N_11601,N_11885);
nand U12244 (N_12244,N_11675,N_11862);
nand U12245 (N_12245,N_11692,N_11921);
xor U12246 (N_12246,N_11815,N_11616);
and U12247 (N_12247,N_11687,N_11720);
nand U12248 (N_12248,N_11764,N_11833);
nor U12249 (N_12249,N_11704,N_11907);
and U12250 (N_12250,N_11877,N_11739);
nand U12251 (N_12251,N_11625,N_11500);
nor U12252 (N_12252,N_11946,N_11997);
xnor U12253 (N_12253,N_11933,N_11874);
or U12254 (N_12254,N_11707,N_11564);
nor U12255 (N_12255,N_11816,N_11756);
xor U12256 (N_12256,N_11707,N_11922);
nand U12257 (N_12257,N_11904,N_11853);
or U12258 (N_12258,N_11592,N_11680);
and U12259 (N_12259,N_11770,N_11713);
or U12260 (N_12260,N_11910,N_11737);
nor U12261 (N_12261,N_11753,N_11955);
or U12262 (N_12262,N_11794,N_11817);
and U12263 (N_12263,N_11775,N_11904);
and U12264 (N_12264,N_11551,N_11773);
nor U12265 (N_12265,N_11620,N_11990);
nand U12266 (N_12266,N_11573,N_11704);
and U12267 (N_12267,N_11912,N_11938);
xnor U12268 (N_12268,N_11604,N_11972);
or U12269 (N_12269,N_11998,N_11537);
nor U12270 (N_12270,N_11543,N_11662);
or U12271 (N_12271,N_11777,N_11656);
nor U12272 (N_12272,N_11922,N_11556);
or U12273 (N_12273,N_11862,N_11520);
and U12274 (N_12274,N_11948,N_11859);
nor U12275 (N_12275,N_11712,N_11736);
or U12276 (N_12276,N_11621,N_11950);
nand U12277 (N_12277,N_11797,N_11847);
and U12278 (N_12278,N_11586,N_11530);
and U12279 (N_12279,N_11567,N_11771);
nand U12280 (N_12280,N_11921,N_11669);
and U12281 (N_12281,N_11933,N_11720);
nand U12282 (N_12282,N_11598,N_11932);
and U12283 (N_12283,N_11681,N_11863);
nor U12284 (N_12284,N_11872,N_11589);
nor U12285 (N_12285,N_11618,N_11635);
nor U12286 (N_12286,N_11548,N_11558);
and U12287 (N_12287,N_11780,N_11848);
or U12288 (N_12288,N_11978,N_11750);
nand U12289 (N_12289,N_11642,N_11680);
xor U12290 (N_12290,N_11533,N_11939);
and U12291 (N_12291,N_11516,N_11853);
and U12292 (N_12292,N_11776,N_11683);
and U12293 (N_12293,N_11776,N_11656);
or U12294 (N_12294,N_11797,N_11964);
and U12295 (N_12295,N_11889,N_11671);
nor U12296 (N_12296,N_11913,N_11702);
or U12297 (N_12297,N_11796,N_11934);
and U12298 (N_12298,N_11709,N_11680);
and U12299 (N_12299,N_11682,N_11663);
or U12300 (N_12300,N_11647,N_11626);
and U12301 (N_12301,N_11570,N_11958);
and U12302 (N_12302,N_11595,N_11886);
nor U12303 (N_12303,N_11818,N_11741);
nor U12304 (N_12304,N_11659,N_11662);
and U12305 (N_12305,N_11863,N_11964);
or U12306 (N_12306,N_11569,N_11616);
and U12307 (N_12307,N_11669,N_11648);
nor U12308 (N_12308,N_11669,N_11545);
nor U12309 (N_12309,N_11986,N_11540);
nand U12310 (N_12310,N_11563,N_11689);
and U12311 (N_12311,N_11649,N_11810);
nand U12312 (N_12312,N_11580,N_11508);
nand U12313 (N_12313,N_11647,N_11854);
nand U12314 (N_12314,N_11697,N_11682);
nor U12315 (N_12315,N_11760,N_11781);
nor U12316 (N_12316,N_11503,N_11838);
or U12317 (N_12317,N_11711,N_11607);
nor U12318 (N_12318,N_11796,N_11932);
nor U12319 (N_12319,N_11607,N_11795);
nor U12320 (N_12320,N_11543,N_11731);
nor U12321 (N_12321,N_11831,N_11924);
or U12322 (N_12322,N_11508,N_11958);
nand U12323 (N_12323,N_11984,N_11772);
nor U12324 (N_12324,N_11628,N_11821);
xor U12325 (N_12325,N_11982,N_11943);
nor U12326 (N_12326,N_11601,N_11609);
or U12327 (N_12327,N_11604,N_11822);
nor U12328 (N_12328,N_11674,N_11797);
xnor U12329 (N_12329,N_11650,N_11860);
nand U12330 (N_12330,N_11574,N_11898);
or U12331 (N_12331,N_11638,N_11507);
nand U12332 (N_12332,N_11721,N_11999);
and U12333 (N_12333,N_11778,N_11532);
nor U12334 (N_12334,N_11922,N_11696);
nand U12335 (N_12335,N_11747,N_11895);
xnor U12336 (N_12336,N_11937,N_11918);
nor U12337 (N_12337,N_11656,N_11510);
and U12338 (N_12338,N_11558,N_11732);
and U12339 (N_12339,N_11944,N_11752);
or U12340 (N_12340,N_11762,N_11695);
and U12341 (N_12341,N_11662,N_11557);
and U12342 (N_12342,N_11880,N_11548);
nand U12343 (N_12343,N_11966,N_11931);
nand U12344 (N_12344,N_11845,N_11557);
or U12345 (N_12345,N_11791,N_11803);
or U12346 (N_12346,N_11775,N_11728);
nor U12347 (N_12347,N_11659,N_11897);
and U12348 (N_12348,N_11635,N_11990);
nand U12349 (N_12349,N_11740,N_11889);
nand U12350 (N_12350,N_11761,N_11616);
or U12351 (N_12351,N_11710,N_11552);
xor U12352 (N_12352,N_11837,N_11894);
nor U12353 (N_12353,N_11852,N_11574);
or U12354 (N_12354,N_11612,N_11864);
nand U12355 (N_12355,N_11704,N_11979);
nor U12356 (N_12356,N_11838,N_11771);
and U12357 (N_12357,N_11813,N_11685);
nand U12358 (N_12358,N_11524,N_11881);
or U12359 (N_12359,N_11689,N_11642);
or U12360 (N_12360,N_11568,N_11616);
nand U12361 (N_12361,N_11509,N_11934);
nand U12362 (N_12362,N_11875,N_11846);
and U12363 (N_12363,N_11649,N_11971);
nand U12364 (N_12364,N_11849,N_11879);
or U12365 (N_12365,N_11562,N_11929);
nand U12366 (N_12366,N_11672,N_11845);
or U12367 (N_12367,N_11639,N_11562);
xnor U12368 (N_12368,N_11537,N_11770);
nand U12369 (N_12369,N_11724,N_11972);
nand U12370 (N_12370,N_11895,N_11874);
nor U12371 (N_12371,N_11769,N_11770);
xnor U12372 (N_12372,N_11522,N_11717);
nand U12373 (N_12373,N_11567,N_11639);
or U12374 (N_12374,N_11604,N_11580);
and U12375 (N_12375,N_11549,N_11937);
or U12376 (N_12376,N_11949,N_11895);
nor U12377 (N_12377,N_11922,N_11749);
xnor U12378 (N_12378,N_11601,N_11673);
and U12379 (N_12379,N_11775,N_11666);
or U12380 (N_12380,N_11602,N_11619);
or U12381 (N_12381,N_11771,N_11910);
and U12382 (N_12382,N_11879,N_11877);
nor U12383 (N_12383,N_11828,N_11518);
and U12384 (N_12384,N_11964,N_11672);
nor U12385 (N_12385,N_11928,N_11938);
and U12386 (N_12386,N_11894,N_11977);
or U12387 (N_12387,N_11773,N_11768);
and U12388 (N_12388,N_11680,N_11771);
nor U12389 (N_12389,N_11503,N_11650);
or U12390 (N_12390,N_11910,N_11717);
xor U12391 (N_12391,N_11706,N_11680);
and U12392 (N_12392,N_11671,N_11771);
nand U12393 (N_12393,N_11661,N_11583);
or U12394 (N_12394,N_11781,N_11801);
nor U12395 (N_12395,N_11562,N_11973);
xor U12396 (N_12396,N_11547,N_11704);
nor U12397 (N_12397,N_11734,N_11502);
and U12398 (N_12398,N_11862,N_11591);
nand U12399 (N_12399,N_11622,N_11579);
and U12400 (N_12400,N_11860,N_11611);
or U12401 (N_12401,N_11824,N_11725);
nor U12402 (N_12402,N_11979,N_11536);
or U12403 (N_12403,N_11799,N_11631);
or U12404 (N_12404,N_11550,N_11799);
nor U12405 (N_12405,N_11798,N_11749);
and U12406 (N_12406,N_11929,N_11735);
nor U12407 (N_12407,N_11687,N_11509);
or U12408 (N_12408,N_11939,N_11864);
and U12409 (N_12409,N_11876,N_11889);
and U12410 (N_12410,N_11992,N_11996);
or U12411 (N_12411,N_11977,N_11860);
xnor U12412 (N_12412,N_11763,N_11900);
or U12413 (N_12413,N_11819,N_11743);
nor U12414 (N_12414,N_11544,N_11976);
and U12415 (N_12415,N_11931,N_11547);
and U12416 (N_12416,N_11571,N_11686);
xnor U12417 (N_12417,N_11637,N_11805);
xnor U12418 (N_12418,N_11584,N_11890);
nand U12419 (N_12419,N_11628,N_11985);
nand U12420 (N_12420,N_11503,N_11754);
or U12421 (N_12421,N_11717,N_11822);
nor U12422 (N_12422,N_11853,N_11767);
and U12423 (N_12423,N_11940,N_11695);
and U12424 (N_12424,N_11841,N_11867);
nor U12425 (N_12425,N_11999,N_11757);
xor U12426 (N_12426,N_11824,N_11841);
and U12427 (N_12427,N_11857,N_11815);
nand U12428 (N_12428,N_11869,N_11554);
nor U12429 (N_12429,N_11710,N_11648);
nor U12430 (N_12430,N_11759,N_11988);
and U12431 (N_12431,N_11747,N_11969);
or U12432 (N_12432,N_11502,N_11537);
nor U12433 (N_12433,N_11818,N_11880);
or U12434 (N_12434,N_11573,N_11763);
nor U12435 (N_12435,N_11647,N_11932);
or U12436 (N_12436,N_11669,N_11580);
nor U12437 (N_12437,N_11567,N_11995);
or U12438 (N_12438,N_11836,N_11620);
nor U12439 (N_12439,N_11800,N_11635);
nand U12440 (N_12440,N_11783,N_11993);
nor U12441 (N_12441,N_11835,N_11854);
and U12442 (N_12442,N_11735,N_11977);
and U12443 (N_12443,N_11898,N_11886);
or U12444 (N_12444,N_11541,N_11947);
or U12445 (N_12445,N_11707,N_11611);
or U12446 (N_12446,N_11941,N_11936);
nor U12447 (N_12447,N_11562,N_11803);
nand U12448 (N_12448,N_11723,N_11669);
nor U12449 (N_12449,N_11636,N_11639);
or U12450 (N_12450,N_11821,N_11858);
and U12451 (N_12451,N_11911,N_11883);
nand U12452 (N_12452,N_11739,N_11505);
and U12453 (N_12453,N_11839,N_11989);
and U12454 (N_12454,N_11518,N_11559);
or U12455 (N_12455,N_11851,N_11982);
and U12456 (N_12456,N_11904,N_11956);
and U12457 (N_12457,N_11699,N_11524);
nor U12458 (N_12458,N_11805,N_11851);
nand U12459 (N_12459,N_11746,N_11824);
nand U12460 (N_12460,N_11768,N_11592);
and U12461 (N_12461,N_11909,N_11977);
or U12462 (N_12462,N_11784,N_11978);
xnor U12463 (N_12463,N_11571,N_11608);
xnor U12464 (N_12464,N_11775,N_11515);
xnor U12465 (N_12465,N_11561,N_11828);
nor U12466 (N_12466,N_11800,N_11861);
or U12467 (N_12467,N_11833,N_11955);
nand U12468 (N_12468,N_11965,N_11946);
and U12469 (N_12469,N_11918,N_11879);
nand U12470 (N_12470,N_11910,N_11842);
or U12471 (N_12471,N_11849,N_11949);
or U12472 (N_12472,N_11926,N_11617);
nand U12473 (N_12473,N_11696,N_11907);
or U12474 (N_12474,N_11713,N_11718);
or U12475 (N_12475,N_11845,N_11844);
nand U12476 (N_12476,N_11538,N_11702);
nand U12477 (N_12477,N_11566,N_11973);
or U12478 (N_12478,N_11611,N_11709);
or U12479 (N_12479,N_11544,N_11506);
nand U12480 (N_12480,N_11933,N_11576);
or U12481 (N_12481,N_11951,N_11701);
nand U12482 (N_12482,N_11580,N_11664);
nand U12483 (N_12483,N_11655,N_11926);
xnor U12484 (N_12484,N_11677,N_11631);
nor U12485 (N_12485,N_11633,N_11504);
nand U12486 (N_12486,N_11816,N_11815);
nor U12487 (N_12487,N_11787,N_11683);
and U12488 (N_12488,N_11826,N_11843);
or U12489 (N_12489,N_11640,N_11771);
nand U12490 (N_12490,N_11957,N_11871);
and U12491 (N_12491,N_11742,N_11669);
xnor U12492 (N_12492,N_11917,N_11756);
nor U12493 (N_12493,N_11760,N_11963);
and U12494 (N_12494,N_11582,N_11513);
nor U12495 (N_12495,N_11540,N_11936);
xnor U12496 (N_12496,N_11511,N_11912);
nand U12497 (N_12497,N_11856,N_11746);
nor U12498 (N_12498,N_11731,N_11845);
and U12499 (N_12499,N_11824,N_11994);
and U12500 (N_12500,N_12073,N_12384);
nand U12501 (N_12501,N_12252,N_12458);
nand U12502 (N_12502,N_12326,N_12291);
nand U12503 (N_12503,N_12297,N_12159);
nand U12504 (N_12504,N_12399,N_12242);
nand U12505 (N_12505,N_12048,N_12164);
and U12506 (N_12506,N_12107,N_12112);
xnor U12507 (N_12507,N_12488,N_12121);
xnor U12508 (N_12508,N_12306,N_12434);
nand U12509 (N_12509,N_12483,N_12081);
xnor U12510 (N_12510,N_12096,N_12018);
nand U12511 (N_12511,N_12473,N_12254);
nor U12512 (N_12512,N_12077,N_12286);
nand U12513 (N_12513,N_12479,N_12221);
xor U12514 (N_12514,N_12336,N_12064);
xnor U12515 (N_12515,N_12255,N_12114);
and U12516 (N_12516,N_12367,N_12403);
or U12517 (N_12517,N_12176,N_12448);
nor U12518 (N_12518,N_12147,N_12020);
xnor U12519 (N_12519,N_12142,N_12146);
or U12520 (N_12520,N_12237,N_12000);
or U12521 (N_12521,N_12318,N_12080);
or U12522 (N_12522,N_12315,N_12132);
nor U12523 (N_12523,N_12011,N_12395);
nand U12524 (N_12524,N_12420,N_12332);
nand U12525 (N_12525,N_12365,N_12006);
xnor U12526 (N_12526,N_12225,N_12460);
and U12527 (N_12527,N_12193,N_12102);
or U12528 (N_12528,N_12314,N_12369);
nand U12529 (N_12529,N_12490,N_12359);
and U12530 (N_12530,N_12465,N_12281);
nand U12531 (N_12531,N_12117,N_12498);
and U12532 (N_12532,N_12189,N_12247);
xnor U12533 (N_12533,N_12099,N_12249);
nand U12534 (N_12534,N_12026,N_12425);
and U12535 (N_12535,N_12098,N_12442);
or U12536 (N_12536,N_12285,N_12139);
or U12537 (N_12537,N_12371,N_12033);
nand U12538 (N_12538,N_12497,N_12426);
nand U12539 (N_12539,N_12309,N_12109);
and U12540 (N_12540,N_12432,N_12041);
nand U12541 (N_12541,N_12447,N_12428);
and U12542 (N_12542,N_12331,N_12317);
or U12543 (N_12543,N_12400,N_12195);
or U12544 (N_12544,N_12040,N_12450);
nor U12545 (N_12545,N_12330,N_12036);
and U12546 (N_12546,N_12191,N_12017);
nand U12547 (N_12547,N_12269,N_12272);
and U12548 (N_12548,N_12230,N_12149);
nand U12549 (N_12549,N_12407,N_12050);
nand U12550 (N_12550,N_12224,N_12072);
nor U12551 (N_12551,N_12101,N_12328);
nand U12552 (N_12552,N_12235,N_12423);
and U12553 (N_12553,N_12268,N_12324);
and U12554 (N_12554,N_12484,N_12223);
nand U12555 (N_12555,N_12319,N_12051);
or U12556 (N_12556,N_12244,N_12311);
or U12557 (N_12557,N_12207,N_12105);
xnor U12558 (N_12558,N_12476,N_12203);
and U12559 (N_12559,N_12469,N_12499);
nor U12560 (N_12560,N_12023,N_12370);
and U12561 (N_12561,N_12045,N_12402);
nand U12562 (N_12562,N_12008,N_12486);
nand U12563 (N_12563,N_12382,N_12313);
nand U12564 (N_12564,N_12405,N_12350);
xnor U12565 (N_12565,N_12438,N_12414);
and U12566 (N_12566,N_12019,N_12219);
nor U12567 (N_12567,N_12456,N_12113);
nor U12568 (N_12568,N_12358,N_12322);
and U12569 (N_12569,N_12002,N_12089);
nand U12570 (N_12570,N_12094,N_12321);
and U12571 (N_12571,N_12063,N_12192);
or U12572 (N_12572,N_12393,N_12348);
nand U12573 (N_12573,N_12119,N_12377);
xor U12574 (N_12574,N_12152,N_12014);
and U12575 (N_12575,N_12129,N_12341);
nand U12576 (N_12576,N_12214,N_12282);
nor U12577 (N_12577,N_12446,N_12211);
xnor U12578 (N_12578,N_12179,N_12386);
or U12579 (N_12579,N_12238,N_12250);
nor U12580 (N_12580,N_12210,N_12168);
nor U12581 (N_12581,N_12131,N_12108);
or U12582 (N_12582,N_12294,N_12482);
nand U12583 (N_12583,N_12299,N_12441);
nor U12584 (N_12584,N_12376,N_12001);
nand U12585 (N_12585,N_12177,N_12277);
xnor U12586 (N_12586,N_12346,N_12429);
or U12587 (N_12587,N_12273,N_12069);
or U12588 (N_12588,N_12271,N_12160);
nand U12589 (N_12589,N_12337,N_12290);
nor U12590 (N_12590,N_12355,N_12354);
or U12591 (N_12591,N_12178,N_12095);
nor U12592 (N_12592,N_12188,N_12245);
or U12593 (N_12593,N_12270,N_12467);
nor U12594 (N_12594,N_12103,N_12031);
xnor U12595 (N_12595,N_12265,N_12340);
or U12596 (N_12596,N_12039,N_12136);
nand U12597 (N_12597,N_12278,N_12258);
nand U12598 (N_12598,N_12363,N_12165);
nor U12599 (N_12599,N_12366,N_12161);
or U12600 (N_12600,N_12431,N_12236);
nor U12601 (N_12601,N_12260,N_12130);
and U12602 (N_12602,N_12185,N_12391);
or U12603 (N_12603,N_12397,N_12086);
and U12604 (N_12604,N_12406,N_12443);
nand U12605 (N_12605,N_12323,N_12227);
or U12606 (N_12606,N_12216,N_12228);
xnor U12607 (N_12607,N_12015,N_12459);
nor U12608 (N_12608,N_12209,N_12030);
or U12609 (N_12609,N_12283,N_12175);
or U12610 (N_12610,N_12424,N_12356);
nor U12611 (N_12611,N_12170,N_12204);
nor U12612 (N_12612,N_12333,N_12196);
and U12613 (N_12613,N_12257,N_12025);
or U12614 (N_12614,N_12464,N_12375);
nor U12615 (N_12615,N_12259,N_12055);
nand U12616 (N_12616,N_12347,N_12118);
nor U12617 (N_12617,N_12436,N_12262);
or U12618 (N_12618,N_12231,N_12280);
xor U12619 (N_12619,N_12120,N_12145);
and U12620 (N_12620,N_12419,N_12357);
nand U12621 (N_12621,N_12032,N_12368);
or U12622 (N_12622,N_12300,N_12218);
xor U12623 (N_12623,N_12302,N_12275);
xnor U12624 (N_12624,N_12292,N_12415);
or U12625 (N_12625,N_12016,N_12056);
nor U12626 (N_12626,N_12213,N_12220);
xor U12627 (N_12627,N_12453,N_12138);
xor U12628 (N_12628,N_12116,N_12061);
or U12629 (N_12629,N_12480,N_12493);
and U12630 (N_12630,N_12455,N_12110);
nand U12631 (N_12631,N_12457,N_12345);
and U12632 (N_12632,N_12007,N_12401);
or U12633 (N_12633,N_12229,N_12416);
or U12634 (N_12634,N_12339,N_12035);
or U12635 (N_12635,N_12334,N_12353);
and U12636 (N_12636,N_12287,N_12241);
nand U12637 (N_12637,N_12010,N_12215);
and U12638 (N_12638,N_12123,N_12233);
and U12639 (N_12639,N_12454,N_12304);
and U12640 (N_12640,N_12070,N_12044);
nand U12641 (N_12641,N_12157,N_12279);
xnor U12642 (N_12642,N_12404,N_12274);
or U12643 (N_12643,N_12184,N_12494);
nor U12644 (N_12644,N_12390,N_12090);
or U12645 (N_12645,N_12474,N_12325);
nand U12646 (N_12646,N_12174,N_12451);
nor U12647 (N_12647,N_12388,N_12135);
and U12648 (N_12648,N_12127,N_12009);
nor U12649 (N_12649,N_12289,N_12182);
or U12650 (N_12650,N_12128,N_12083);
and U12651 (N_12651,N_12343,N_12091);
xnor U12652 (N_12652,N_12153,N_12351);
and U12653 (N_12653,N_12320,N_12173);
nand U12654 (N_12654,N_12166,N_12288);
or U12655 (N_12655,N_12046,N_12037);
nor U12656 (N_12656,N_12349,N_12410);
nand U12657 (N_12657,N_12004,N_12124);
nand U12658 (N_12658,N_12155,N_12487);
nand U12659 (N_12659,N_12034,N_12059);
xor U12660 (N_12660,N_12243,N_12167);
nand U12661 (N_12661,N_12085,N_12012);
nor U12662 (N_12662,N_12200,N_12158);
and U12663 (N_12663,N_12327,N_12435);
and U12664 (N_12664,N_12125,N_12115);
nor U12665 (N_12665,N_12495,N_12389);
or U12666 (N_12666,N_12372,N_12162);
nand U12667 (N_12667,N_12133,N_12104);
and U12668 (N_12668,N_12137,N_12013);
nand U12669 (N_12669,N_12226,N_12197);
xor U12670 (N_12670,N_12043,N_12444);
and U12671 (N_12671,N_12088,N_12276);
and U12672 (N_12672,N_12169,N_12461);
or U12673 (N_12673,N_12201,N_12383);
and U12674 (N_12674,N_12413,N_12100);
xnor U12675 (N_12675,N_12251,N_12392);
nor U12676 (N_12676,N_12471,N_12364);
nor U12677 (N_12677,N_12478,N_12163);
and U12678 (N_12678,N_12409,N_12361);
and U12679 (N_12679,N_12298,N_12148);
or U12680 (N_12680,N_12053,N_12187);
nand U12681 (N_12681,N_12057,N_12418);
nor U12682 (N_12682,N_12047,N_12154);
xnor U12683 (N_12683,N_12212,N_12335);
nor U12684 (N_12684,N_12344,N_12144);
and U12685 (N_12685,N_12087,N_12097);
nand U12686 (N_12686,N_12303,N_12232);
xor U12687 (N_12687,N_12060,N_12068);
nand U12688 (N_12688,N_12411,N_12111);
or U12689 (N_12689,N_12208,N_12199);
or U12690 (N_12690,N_12263,N_12362);
and U12691 (N_12691,N_12295,N_12234);
nor U12692 (N_12692,N_12470,N_12305);
xor U12693 (N_12693,N_12076,N_12477);
or U12694 (N_12694,N_12445,N_12449);
nand U12695 (N_12695,N_12217,N_12452);
nor U12696 (N_12696,N_12143,N_12038);
nor U12697 (N_12697,N_12052,N_12338);
nand U12698 (N_12698,N_12183,N_12062);
and U12699 (N_12699,N_12472,N_12082);
nor U12700 (N_12700,N_12222,N_12181);
nand U12701 (N_12701,N_12394,N_12439);
xor U12702 (N_12702,N_12342,N_12190);
nand U12703 (N_12703,N_12027,N_12239);
nor U12704 (N_12704,N_12022,N_12024);
nor U12705 (N_12705,N_12316,N_12466);
or U12706 (N_12706,N_12079,N_12058);
and U12707 (N_12707,N_12408,N_12180);
or U12708 (N_12708,N_12092,N_12093);
and U12709 (N_12709,N_12156,N_12475);
nand U12710 (N_12710,N_12374,N_12003);
and U12711 (N_12711,N_12310,N_12150);
nor U12712 (N_12712,N_12385,N_12054);
and U12713 (N_12713,N_12496,N_12378);
xnor U12714 (N_12714,N_12122,N_12489);
and U12715 (N_12715,N_12381,N_12248);
nor U12716 (N_12716,N_12186,N_12106);
and U12717 (N_12717,N_12421,N_12067);
and U12718 (N_12718,N_12194,N_12440);
nor U12719 (N_12719,N_12261,N_12065);
nand U12720 (N_12720,N_12387,N_12240);
xor U12721 (N_12721,N_12134,N_12430);
nor U12722 (N_12722,N_12312,N_12049);
nand U12723 (N_12723,N_12066,N_12246);
nand U12724 (N_12724,N_12028,N_12264);
and U12725 (N_12725,N_12396,N_12266);
and U12726 (N_12726,N_12029,N_12485);
nand U12727 (N_12727,N_12427,N_12198);
xor U12728 (N_12728,N_12206,N_12492);
or U12729 (N_12729,N_12463,N_12141);
or U12730 (N_12730,N_12284,N_12267);
nand U12731 (N_12731,N_12462,N_12352);
nor U12732 (N_12732,N_12433,N_12308);
nor U12733 (N_12733,N_12296,N_12084);
and U12734 (N_12734,N_12373,N_12005);
or U12735 (N_12735,N_12075,N_12437);
nor U12736 (N_12736,N_12253,N_12071);
and U12737 (N_12737,N_12293,N_12379);
nand U12738 (N_12738,N_12380,N_12202);
xor U12739 (N_12739,N_12205,N_12172);
and U12740 (N_12740,N_12074,N_12301);
xnor U12741 (N_12741,N_12021,N_12398);
nand U12742 (N_12742,N_12491,N_12417);
and U12743 (N_12743,N_12481,N_12307);
and U12744 (N_12744,N_12078,N_12412);
nand U12745 (N_12745,N_12256,N_12468);
nor U12746 (N_12746,N_12126,N_12329);
nand U12747 (N_12747,N_12140,N_12422);
nor U12748 (N_12748,N_12042,N_12171);
nand U12749 (N_12749,N_12360,N_12151);
nand U12750 (N_12750,N_12348,N_12163);
or U12751 (N_12751,N_12379,N_12345);
and U12752 (N_12752,N_12104,N_12130);
nand U12753 (N_12753,N_12005,N_12315);
or U12754 (N_12754,N_12497,N_12200);
or U12755 (N_12755,N_12492,N_12191);
nor U12756 (N_12756,N_12165,N_12392);
and U12757 (N_12757,N_12371,N_12456);
nor U12758 (N_12758,N_12134,N_12270);
or U12759 (N_12759,N_12426,N_12072);
nand U12760 (N_12760,N_12406,N_12432);
and U12761 (N_12761,N_12397,N_12220);
nand U12762 (N_12762,N_12438,N_12419);
and U12763 (N_12763,N_12257,N_12273);
nand U12764 (N_12764,N_12308,N_12201);
or U12765 (N_12765,N_12040,N_12485);
xnor U12766 (N_12766,N_12088,N_12474);
nand U12767 (N_12767,N_12110,N_12286);
nand U12768 (N_12768,N_12083,N_12427);
or U12769 (N_12769,N_12367,N_12158);
and U12770 (N_12770,N_12071,N_12399);
nor U12771 (N_12771,N_12449,N_12175);
and U12772 (N_12772,N_12008,N_12389);
nor U12773 (N_12773,N_12410,N_12228);
or U12774 (N_12774,N_12318,N_12453);
xnor U12775 (N_12775,N_12105,N_12300);
or U12776 (N_12776,N_12177,N_12094);
nand U12777 (N_12777,N_12099,N_12208);
xor U12778 (N_12778,N_12473,N_12422);
or U12779 (N_12779,N_12058,N_12283);
and U12780 (N_12780,N_12492,N_12483);
nand U12781 (N_12781,N_12276,N_12483);
nor U12782 (N_12782,N_12350,N_12263);
xnor U12783 (N_12783,N_12147,N_12148);
nor U12784 (N_12784,N_12327,N_12310);
nor U12785 (N_12785,N_12224,N_12478);
xor U12786 (N_12786,N_12138,N_12047);
nand U12787 (N_12787,N_12280,N_12288);
nor U12788 (N_12788,N_12214,N_12457);
or U12789 (N_12789,N_12477,N_12250);
nand U12790 (N_12790,N_12241,N_12389);
and U12791 (N_12791,N_12489,N_12373);
nor U12792 (N_12792,N_12351,N_12310);
or U12793 (N_12793,N_12349,N_12126);
xnor U12794 (N_12794,N_12495,N_12493);
or U12795 (N_12795,N_12065,N_12306);
xor U12796 (N_12796,N_12172,N_12306);
or U12797 (N_12797,N_12299,N_12294);
or U12798 (N_12798,N_12013,N_12316);
nand U12799 (N_12799,N_12206,N_12273);
and U12800 (N_12800,N_12451,N_12176);
nand U12801 (N_12801,N_12441,N_12058);
or U12802 (N_12802,N_12336,N_12072);
nand U12803 (N_12803,N_12081,N_12198);
and U12804 (N_12804,N_12339,N_12491);
nor U12805 (N_12805,N_12165,N_12260);
xnor U12806 (N_12806,N_12032,N_12088);
xor U12807 (N_12807,N_12465,N_12072);
nor U12808 (N_12808,N_12087,N_12305);
or U12809 (N_12809,N_12341,N_12396);
and U12810 (N_12810,N_12277,N_12185);
nand U12811 (N_12811,N_12076,N_12087);
or U12812 (N_12812,N_12170,N_12173);
nand U12813 (N_12813,N_12303,N_12226);
xnor U12814 (N_12814,N_12273,N_12339);
nand U12815 (N_12815,N_12169,N_12130);
nor U12816 (N_12816,N_12401,N_12186);
and U12817 (N_12817,N_12310,N_12000);
nor U12818 (N_12818,N_12304,N_12147);
and U12819 (N_12819,N_12259,N_12146);
or U12820 (N_12820,N_12459,N_12390);
or U12821 (N_12821,N_12171,N_12352);
xor U12822 (N_12822,N_12290,N_12196);
and U12823 (N_12823,N_12219,N_12233);
or U12824 (N_12824,N_12132,N_12083);
and U12825 (N_12825,N_12048,N_12073);
and U12826 (N_12826,N_12359,N_12434);
nor U12827 (N_12827,N_12427,N_12495);
and U12828 (N_12828,N_12458,N_12229);
xnor U12829 (N_12829,N_12055,N_12296);
nor U12830 (N_12830,N_12272,N_12115);
nor U12831 (N_12831,N_12155,N_12457);
nor U12832 (N_12832,N_12004,N_12169);
and U12833 (N_12833,N_12443,N_12000);
nor U12834 (N_12834,N_12355,N_12332);
nor U12835 (N_12835,N_12092,N_12244);
or U12836 (N_12836,N_12301,N_12479);
or U12837 (N_12837,N_12318,N_12361);
and U12838 (N_12838,N_12490,N_12340);
or U12839 (N_12839,N_12074,N_12110);
nor U12840 (N_12840,N_12003,N_12362);
nor U12841 (N_12841,N_12150,N_12193);
or U12842 (N_12842,N_12427,N_12139);
or U12843 (N_12843,N_12183,N_12013);
or U12844 (N_12844,N_12181,N_12416);
and U12845 (N_12845,N_12202,N_12119);
or U12846 (N_12846,N_12071,N_12417);
xor U12847 (N_12847,N_12476,N_12202);
nor U12848 (N_12848,N_12468,N_12465);
nand U12849 (N_12849,N_12151,N_12029);
xnor U12850 (N_12850,N_12183,N_12412);
or U12851 (N_12851,N_12331,N_12080);
nand U12852 (N_12852,N_12223,N_12042);
and U12853 (N_12853,N_12031,N_12105);
nor U12854 (N_12854,N_12064,N_12102);
xor U12855 (N_12855,N_12271,N_12365);
and U12856 (N_12856,N_12140,N_12284);
nor U12857 (N_12857,N_12463,N_12075);
nor U12858 (N_12858,N_12253,N_12148);
nand U12859 (N_12859,N_12145,N_12187);
and U12860 (N_12860,N_12277,N_12391);
nor U12861 (N_12861,N_12383,N_12040);
nand U12862 (N_12862,N_12286,N_12118);
xnor U12863 (N_12863,N_12372,N_12164);
nand U12864 (N_12864,N_12011,N_12137);
nor U12865 (N_12865,N_12175,N_12406);
or U12866 (N_12866,N_12221,N_12209);
xnor U12867 (N_12867,N_12099,N_12400);
and U12868 (N_12868,N_12098,N_12154);
nand U12869 (N_12869,N_12046,N_12377);
nand U12870 (N_12870,N_12158,N_12061);
nor U12871 (N_12871,N_12399,N_12332);
or U12872 (N_12872,N_12145,N_12189);
nand U12873 (N_12873,N_12042,N_12496);
nand U12874 (N_12874,N_12160,N_12212);
and U12875 (N_12875,N_12096,N_12278);
and U12876 (N_12876,N_12278,N_12450);
nand U12877 (N_12877,N_12015,N_12142);
xor U12878 (N_12878,N_12052,N_12263);
and U12879 (N_12879,N_12412,N_12205);
nand U12880 (N_12880,N_12252,N_12124);
or U12881 (N_12881,N_12200,N_12206);
and U12882 (N_12882,N_12412,N_12426);
nor U12883 (N_12883,N_12376,N_12021);
nor U12884 (N_12884,N_12222,N_12164);
nand U12885 (N_12885,N_12181,N_12170);
nand U12886 (N_12886,N_12463,N_12104);
xor U12887 (N_12887,N_12059,N_12008);
nand U12888 (N_12888,N_12334,N_12406);
nand U12889 (N_12889,N_12479,N_12385);
nand U12890 (N_12890,N_12320,N_12499);
and U12891 (N_12891,N_12154,N_12478);
nor U12892 (N_12892,N_12100,N_12000);
or U12893 (N_12893,N_12426,N_12268);
nand U12894 (N_12894,N_12438,N_12096);
or U12895 (N_12895,N_12377,N_12147);
and U12896 (N_12896,N_12045,N_12009);
nand U12897 (N_12897,N_12397,N_12317);
and U12898 (N_12898,N_12223,N_12152);
or U12899 (N_12899,N_12090,N_12034);
xnor U12900 (N_12900,N_12431,N_12393);
and U12901 (N_12901,N_12392,N_12400);
nor U12902 (N_12902,N_12202,N_12251);
nor U12903 (N_12903,N_12415,N_12386);
nand U12904 (N_12904,N_12245,N_12425);
nand U12905 (N_12905,N_12348,N_12478);
nor U12906 (N_12906,N_12269,N_12048);
nand U12907 (N_12907,N_12197,N_12158);
and U12908 (N_12908,N_12297,N_12203);
nand U12909 (N_12909,N_12251,N_12278);
nor U12910 (N_12910,N_12281,N_12229);
and U12911 (N_12911,N_12316,N_12173);
and U12912 (N_12912,N_12494,N_12424);
nor U12913 (N_12913,N_12350,N_12437);
and U12914 (N_12914,N_12314,N_12417);
or U12915 (N_12915,N_12028,N_12399);
or U12916 (N_12916,N_12371,N_12376);
or U12917 (N_12917,N_12488,N_12339);
nand U12918 (N_12918,N_12036,N_12144);
and U12919 (N_12919,N_12167,N_12394);
nor U12920 (N_12920,N_12210,N_12243);
xnor U12921 (N_12921,N_12108,N_12416);
nand U12922 (N_12922,N_12348,N_12411);
and U12923 (N_12923,N_12196,N_12485);
or U12924 (N_12924,N_12100,N_12441);
nor U12925 (N_12925,N_12048,N_12034);
nand U12926 (N_12926,N_12136,N_12246);
xor U12927 (N_12927,N_12441,N_12331);
nand U12928 (N_12928,N_12276,N_12292);
or U12929 (N_12929,N_12159,N_12016);
and U12930 (N_12930,N_12466,N_12374);
and U12931 (N_12931,N_12108,N_12035);
or U12932 (N_12932,N_12124,N_12370);
nor U12933 (N_12933,N_12252,N_12130);
nand U12934 (N_12934,N_12302,N_12001);
and U12935 (N_12935,N_12029,N_12068);
nand U12936 (N_12936,N_12230,N_12423);
and U12937 (N_12937,N_12012,N_12350);
nand U12938 (N_12938,N_12170,N_12389);
or U12939 (N_12939,N_12357,N_12326);
xnor U12940 (N_12940,N_12165,N_12021);
nand U12941 (N_12941,N_12164,N_12474);
nand U12942 (N_12942,N_12345,N_12210);
nand U12943 (N_12943,N_12265,N_12037);
nand U12944 (N_12944,N_12380,N_12361);
nor U12945 (N_12945,N_12249,N_12013);
nor U12946 (N_12946,N_12485,N_12137);
nor U12947 (N_12947,N_12160,N_12386);
and U12948 (N_12948,N_12209,N_12381);
nor U12949 (N_12949,N_12158,N_12201);
nor U12950 (N_12950,N_12176,N_12497);
or U12951 (N_12951,N_12228,N_12096);
or U12952 (N_12952,N_12343,N_12371);
or U12953 (N_12953,N_12486,N_12469);
nor U12954 (N_12954,N_12326,N_12320);
and U12955 (N_12955,N_12286,N_12001);
and U12956 (N_12956,N_12280,N_12159);
xor U12957 (N_12957,N_12011,N_12066);
nand U12958 (N_12958,N_12344,N_12480);
nor U12959 (N_12959,N_12399,N_12361);
or U12960 (N_12960,N_12345,N_12056);
nand U12961 (N_12961,N_12074,N_12313);
nand U12962 (N_12962,N_12179,N_12035);
nor U12963 (N_12963,N_12035,N_12323);
and U12964 (N_12964,N_12425,N_12055);
nor U12965 (N_12965,N_12392,N_12094);
and U12966 (N_12966,N_12227,N_12382);
xnor U12967 (N_12967,N_12329,N_12286);
nand U12968 (N_12968,N_12274,N_12120);
nor U12969 (N_12969,N_12436,N_12160);
xnor U12970 (N_12970,N_12143,N_12460);
nand U12971 (N_12971,N_12037,N_12380);
nor U12972 (N_12972,N_12232,N_12448);
and U12973 (N_12973,N_12345,N_12018);
nor U12974 (N_12974,N_12129,N_12465);
nand U12975 (N_12975,N_12391,N_12360);
and U12976 (N_12976,N_12450,N_12358);
xnor U12977 (N_12977,N_12106,N_12064);
nor U12978 (N_12978,N_12464,N_12177);
nand U12979 (N_12979,N_12044,N_12272);
nor U12980 (N_12980,N_12131,N_12165);
or U12981 (N_12981,N_12307,N_12319);
nand U12982 (N_12982,N_12031,N_12011);
nor U12983 (N_12983,N_12223,N_12176);
or U12984 (N_12984,N_12479,N_12001);
or U12985 (N_12985,N_12396,N_12216);
or U12986 (N_12986,N_12333,N_12167);
nor U12987 (N_12987,N_12104,N_12187);
nand U12988 (N_12988,N_12196,N_12232);
nor U12989 (N_12989,N_12215,N_12038);
and U12990 (N_12990,N_12045,N_12099);
nor U12991 (N_12991,N_12465,N_12178);
and U12992 (N_12992,N_12159,N_12183);
nor U12993 (N_12993,N_12202,N_12099);
nand U12994 (N_12994,N_12018,N_12427);
nor U12995 (N_12995,N_12485,N_12450);
nor U12996 (N_12996,N_12331,N_12354);
or U12997 (N_12997,N_12219,N_12366);
nor U12998 (N_12998,N_12319,N_12035);
nand U12999 (N_12999,N_12154,N_12254);
or U13000 (N_13000,N_12956,N_12853);
and U13001 (N_13001,N_12898,N_12864);
and U13002 (N_13002,N_12984,N_12510);
or U13003 (N_13003,N_12993,N_12845);
nor U13004 (N_13004,N_12810,N_12971);
nor U13005 (N_13005,N_12721,N_12531);
and U13006 (N_13006,N_12896,N_12715);
and U13007 (N_13007,N_12661,N_12940);
nor U13008 (N_13008,N_12842,N_12932);
and U13009 (N_13009,N_12995,N_12773);
or U13010 (N_13010,N_12994,N_12950);
and U13011 (N_13011,N_12849,N_12569);
and U13012 (N_13012,N_12835,N_12673);
and U13013 (N_13013,N_12635,N_12809);
nand U13014 (N_13014,N_12726,N_12762);
nand U13015 (N_13015,N_12527,N_12825);
nor U13016 (N_13016,N_12897,N_12657);
and U13017 (N_13017,N_12700,N_12929);
nor U13018 (N_13018,N_12627,N_12866);
and U13019 (N_13019,N_12970,N_12823);
and U13020 (N_13020,N_12681,N_12728);
or U13021 (N_13021,N_12784,N_12822);
and U13022 (N_13022,N_12892,N_12840);
nor U13023 (N_13023,N_12588,N_12814);
or U13024 (N_13024,N_12985,N_12554);
nor U13025 (N_13025,N_12795,N_12989);
and U13026 (N_13026,N_12912,N_12576);
nor U13027 (N_13027,N_12933,N_12557);
and U13028 (N_13028,N_12677,N_12858);
or U13029 (N_13029,N_12511,N_12747);
nand U13030 (N_13030,N_12753,N_12599);
nor U13031 (N_13031,N_12804,N_12911);
and U13032 (N_13032,N_12902,N_12582);
or U13033 (N_13033,N_12713,N_12552);
nor U13034 (N_13034,N_12818,N_12678);
or U13035 (N_13035,N_12546,N_12913);
nand U13036 (N_13036,N_12847,N_12811);
or U13037 (N_13037,N_12596,N_12951);
and U13038 (N_13038,N_12748,N_12626);
nand U13039 (N_13039,N_12957,N_12535);
and U13040 (N_13040,N_12901,N_12570);
nor U13041 (N_13041,N_12834,N_12996);
and U13042 (N_13042,N_12883,N_12863);
nand U13043 (N_13043,N_12642,N_12826);
nand U13044 (N_13044,N_12653,N_12509);
and U13045 (N_13045,N_12832,N_12530);
nand U13046 (N_13046,N_12663,N_12614);
nor U13047 (N_13047,N_12972,N_12595);
and U13048 (N_13048,N_12587,N_12766);
nand U13049 (N_13049,N_12791,N_12899);
nand U13050 (N_13050,N_12960,N_12656);
nand U13051 (N_13051,N_12550,N_12556);
nor U13052 (N_13052,N_12904,N_12613);
nor U13053 (N_13053,N_12575,N_12819);
nor U13054 (N_13054,N_12860,N_12645);
or U13055 (N_13055,N_12705,N_12695);
nor U13056 (N_13056,N_12871,N_12954);
or U13057 (N_13057,N_12732,N_12693);
or U13058 (N_13058,N_12651,N_12636);
xnor U13059 (N_13059,N_12601,N_12760);
xor U13060 (N_13060,N_12615,N_12749);
and U13061 (N_13061,N_12696,N_12820);
and U13062 (N_13062,N_12606,N_12914);
or U13063 (N_13063,N_12944,N_12528);
or U13064 (N_13064,N_12500,N_12772);
and U13065 (N_13065,N_12514,N_12729);
and U13066 (N_13066,N_12837,N_12859);
xor U13067 (N_13067,N_12807,N_12674);
nand U13068 (N_13068,N_12505,N_12916);
nor U13069 (N_13069,N_12720,N_12768);
nor U13070 (N_13070,N_12709,N_12649);
nand U13071 (N_13071,N_12537,N_12888);
nor U13072 (N_13072,N_12752,N_12694);
nor U13073 (N_13073,N_12880,N_12644);
nor U13074 (N_13074,N_12544,N_12746);
nor U13075 (N_13075,N_12629,N_12586);
nand U13076 (N_13076,N_12563,N_12955);
nand U13077 (N_13077,N_12517,N_12981);
nor U13078 (N_13078,N_12943,N_12787);
xnor U13079 (N_13079,N_12654,N_12877);
or U13080 (N_13080,N_12839,N_12502);
nor U13081 (N_13081,N_12919,N_12549);
nor U13082 (N_13082,N_12688,N_12579);
nand U13083 (N_13083,N_12692,N_12610);
or U13084 (N_13084,N_12506,N_12738);
nor U13085 (N_13085,N_12703,N_12854);
and U13086 (N_13086,N_12894,N_12761);
nand U13087 (N_13087,N_12706,N_12755);
nand U13088 (N_13088,N_12684,N_12648);
nand U13089 (N_13089,N_12875,N_12609);
nand U13090 (N_13090,N_12934,N_12948);
or U13091 (N_13091,N_12691,N_12812);
and U13092 (N_13092,N_12597,N_12959);
nor U13093 (N_13093,N_12638,N_12515);
nor U13094 (N_13094,N_12930,N_12872);
nor U13095 (N_13095,N_12607,N_12660);
nand U13096 (N_13096,N_12725,N_12764);
nor U13097 (N_13097,N_12740,N_12909);
nor U13098 (N_13098,N_12589,N_12824);
and U13099 (N_13099,N_12625,N_12986);
nand U13100 (N_13100,N_12618,N_12590);
and U13101 (N_13101,N_12813,N_12992);
xnor U13102 (N_13102,N_12593,N_12920);
nand U13103 (N_13103,N_12861,N_12758);
nand U13104 (N_13104,N_12591,N_12953);
and U13105 (N_13105,N_12857,N_12947);
or U13106 (N_13106,N_12975,N_12621);
nand U13107 (N_13107,N_12757,N_12682);
nand U13108 (N_13108,N_12829,N_12543);
nor U13109 (N_13109,N_12698,N_12503);
nand U13110 (N_13110,N_12927,N_12577);
nand U13111 (N_13111,N_12988,N_12868);
and U13112 (N_13112,N_12658,N_12905);
nor U13113 (N_13113,N_12873,N_12850);
nand U13114 (N_13114,N_12977,N_12906);
nor U13115 (N_13115,N_12745,N_12718);
xor U13116 (N_13116,N_12910,N_12655);
and U13117 (N_13117,N_12798,N_12632);
nand U13118 (N_13118,N_12806,N_12961);
or U13119 (N_13119,N_12997,N_12548);
nand U13120 (N_13120,N_12519,N_12903);
and U13121 (N_13121,N_12717,N_12782);
and U13122 (N_13122,N_12701,N_12641);
nand U13123 (N_13123,N_12803,N_12634);
or U13124 (N_13124,N_12887,N_12687);
and U13125 (N_13125,N_12767,N_12821);
or U13126 (N_13126,N_12611,N_12838);
nand U13127 (N_13127,N_12884,N_12652);
nor U13128 (N_13128,N_12939,N_12707);
or U13129 (N_13129,N_12763,N_12774);
and U13130 (N_13130,N_12533,N_12900);
and U13131 (N_13131,N_12800,N_12616);
and U13132 (N_13132,N_12802,N_12742);
nand U13133 (N_13133,N_12846,N_12699);
xnor U13134 (N_13134,N_12796,N_12793);
or U13135 (N_13135,N_12555,N_12572);
or U13136 (N_13136,N_12893,N_12672);
or U13137 (N_13137,N_12917,N_12612);
nand U13138 (N_13138,N_12662,N_12711);
or U13139 (N_13139,N_12743,N_12565);
and U13140 (N_13140,N_12668,N_12578);
xor U13141 (N_13141,N_12622,N_12551);
nand U13142 (N_13142,N_12778,N_12559);
and U13143 (N_13143,N_12862,N_12553);
or U13144 (N_13144,N_12815,N_12744);
nand U13145 (N_13145,N_12870,N_12750);
and U13146 (N_13146,N_12967,N_12723);
nor U13147 (N_13147,N_12998,N_12731);
nand U13148 (N_13148,N_12922,N_12666);
or U13149 (N_13149,N_12639,N_12908);
nand U13150 (N_13150,N_12968,N_12801);
nand U13151 (N_13151,N_12874,N_12816);
or U13152 (N_13152,N_12714,N_12524);
nor U13153 (N_13153,N_12679,N_12925);
and U13154 (N_13154,N_12501,N_12879);
nor U13155 (N_13155,N_12584,N_12776);
nor U13156 (N_13156,N_12958,N_12560);
or U13157 (N_13157,N_12878,N_12671);
or U13158 (N_13158,N_12617,N_12504);
nand U13159 (N_13159,N_12799,N_12538);
nand U13160 (N_13160,N_12710,N_12737);
and U13161 (N_13161,N_12921,N_12759);
and U13162 (N_13162,N_12885,N_12828);
nand U13163 (N_13163,N_12805,N_12980);
nor U13164 (N_13164,N_12526,N_12852);
nand U13165 (N_13165,N_12667,N_12686);
or U13166 (N_13166,N_12628,N_12562);
or U13167 (N_13167,N_12963,N_12594);
or U13168 (N_13168,N_12508,N_12937);
xnor U13169 (N_13169,N_12574,N_12520);
nand U13170 (N_13170,N_12727,N_12633);
nor U13171 (N_13171,N_12895,N_12869);
nand U13172 (N_13172,N_12876,N_12891);
or U13173 (N_13173,N_12935,N_12716);
nand U13174 (N_13174,N_12754,N_12689);
or U13175 (N_13175,N_12928,N_12534);
and U13176 (N_13176,N_12771,N_12739);
nand U13177 (N_13177,N_12830,N_12571);
nand U13178 (N_13178,N_12797,N_12881);
and U13179 (N_13179,N_12915,N_12702);
nand U13180 (N_13180,N_12507,N_12529);
nand U13181 (N_13181,N_12790,N_12525);
and U13182 (N_13182,N_12608,N_12545);
xnor U13183 (N_13183,N_12558,N_12532);
and U13184 (N_13184,N_12604,N_12598);
xor U13185 (N_13185,N_12786,N_12640);
nor U13186 (N_13186,N_12844,N_12965);
or U13187 (N_13187,N_12808,N_12521);
nand U13188 (N_13188,N_12733,N_12769);
xor U13189 (N_13189,N_12573,N_12775);
xnor U13190 (N_13190,N_12924,N_12991);
nor U13191 (N_13191,N_12938,N_12974);
or U13192 (N_13192,N_12539,N_12650);
nor U13193 (N_13193,N_12882,N_12647);
xor U13194 (N_13194,N_12949,N_12827);
nand U13195 (N_13195,N_12973,N_12966);
nand U13196 (N_13196,N_12907,N_12785);
or U13197 (N_13197,N_12741,N_12789);
or U13198 (N_13198,N_12724,N_12946);
and U13199 (N_13199,N_12522,N_12600);
and U13200 (N_13200,N_12665,N_12603);
nand U13201 (N_13201,N_12890,N_12683);
and U13202 (N_13202,N_12719,N_12983);
and U13203 (N_13203,N_12936,N_12630);
and U13204 (N_13204,N_12585,N_12926);
and U13205 (N_13205,N_12540,N_12777);
or U13206 (N_13206,N_12841,N_12792);
nor U13207 (N_13207,N_12856,N_12918);
and U13208 (N_13208,N_12978,N_12583);
nor U13209 (N_13209,N_12547,N_12962);
or U13210 (N_13210,N_12664,N_12886);
and U13211 (N_13211,N_12999,N_12708);
nand U13212 (N_13212,N_12736,N_12561);
nor U13213 (N_13213,N_12923,N_12541);
xor U13214 (N_13214,N_12602,N_12851);
xor U13215 (N_13215,N_12867,N_12865);
or U13216 (N_13216,N_12942,N_12513);
or U13217 (N_13217,N_12964,N_12735);
xnor U13218 (N_13218,N_12567,N_12976);
nor U13219 (N_13219,N_12623,N_12889);
nor U13220 (N_13220,N_12685,N_12581);
and U13221 (N_13221,N_12669,N_12512);
and U13222 (N_13222,N_12783,N_12605);
nor U13223 (N_13223,N_12518,N_12643);
nand U13224 (N_13224,N_12779,N_12848);
and U13225 (N_13225,N_12765,N_12979);
nor U13226 (N_13226,N_12734,N_12697);
nor U13227 (N_13227,N_12945,N_12676);
nand U13228 (N_13228,N_12969,N_12751);
and U13229 (N_13229,N_12794,N_12941);
nor U13230 (N_13230,N_12592,N_12990);
or U13231 (N_13231,N_12624,N_12952);
or U13232 (N_13232,N_12712,N_12542);
and U13233 (N_13233,N_12982,N_12670);
nor U13234 (N_13234,N_12780,N_12931);
and U13235 (N_13235,N_12987,N_12580);
or U13236 (N_13236,N_12730,N_12855);
nor U13237 (N_13237,N_12566,N_12680);
or U13238 (N_13238,N_12843,N_12631);
nor U13239 (N_13239,N_12833,N_12564);
nor U13240 (N_13240,N_12781,N_12536);
nor U13241 (N_13241,N_12637,N_12722);
or U13242 (N_13242,N_12620,N_12516);
nand U13243 (N_13243,N_12770,N_12646);
nor U13244 (N_13244,N_12831,N_12619);
xnor U13245 (N_13245,N_12523,N_12704);
nand U13246 (N_13246,N_12659,N_12788);
nand U13247 (N_13247,N_12675,N_12836);
nand U13248 (N_13248,N_12756,N_12690);
xnor U13249 (N_13249,N_12568,N_12817);
and U13250 (N_13250,N_12575,N_12718);
or U13251 (N_13251,N_12535,N_12784);
or U13252 (N_13252,N_12817,N_12892);
nor U13253 (N_13253,N_12935,N_12888);
nor U13254 (N_13254,N_12527,N_12839);
nor U13255 (N_13255,N_12775,N_12897);
or U13256 (N_13256,N_12834,N_12946);
nand U13257 (N_13257,N_12749,N_12535);
and U13258 (N_13258,N_12924,N_12961);
or U13259 (N_13259,N_12681,N_12869);
or U13260 (N_13260,N_12890,N_12922);
nor U13261 (N_13261,N_12778,N_12714);
and U13262 (N_13262,N_12991,N_12632);
nand U13263 (N_13263,N_12894,N_12925);
nor U13264 (N_13264,N_12811,N_12967);
or U13265 (N_13265,N_12920,N_12600);
nor U13266 (N_13266,N_12567,N_12750);
or U13267 (N_13267,N_12620,N_12590);
or U13268 (N_13268,N_12624,N_12856);
nor U13269 (N_13269,N_12542,N_12554);
xor U13270 (N_13270,N_12667,N_12602);
and U13271 (N_13271,N_12671,N_12623);
xor U13272 (N_13272,N_12980,N_12922);
or U13273 (N_13273,N_12757,N_12768);
or U13274 (N_13274,N_12701,N_12611);
nand U13275 (N_13275,N_12960,N_12702);
nand U13276 (N_13276,N_12528,N_12508);
nor U13277 (N_13277,N_12997,N_12916);
nand U13278 (N_13278,N_12948,N_12802);
and U13279 (N_13279,N_12582,N_12508);
nor U13280 (N_13280,N_12846,N_12648);
nand U13281 (N_13281,N_12616,N_12946);
xnor U13282 (N_13282,N_12592,N_12651);
nor U13283 (N_13283,N_12638,N_12695);
and U13284 (N_13284,N_12577,N_12635);
nor U13285 (N_13285,N_12743,N_12768);
or U13286 (N_13286,N_12702,N_12861);
and U13287 (N_13287,N_12909,N_12906);
nor U13288 (N_13288,N_12700,N_12879);
and U13289 (N_13289,N_12546,N_12554);
nor U13290 (N_13290,N_12722,N_12752);
nor U13291 (N_13291,N_12889,N_12684);
nor U13292 (N_13292,N_12819,N_12581);
and U13293 (N_13293,N_12549,N_12826);
and U13294 (N_13294,N_12593,N_12628);
nand U13295 (N_13295,N_12610,N_12650);
or U13296 (N_13296,N_12928,N_12593);
nand U13297 (N_13297,N_12942,N_12777);
nor U13298 (N_13298,N_12879,N_12852);
nand U13299 (N_13299,N_12597,N_12591);
xor U13300 (N_13300,N_12937,N_12974);
or U13301 (N_13301,N_12589,N_12892);
nand U13302 (N_13302,N_12566,N_12535);
xnor U13303 (N_13303,N_12783,N_12501);
nor U13304 (N_13304,N_12943,N_12573);
xor U13305 (N_13305,N_12814,N_12839);
nand U13306 (N_13306,N_12542,N_12586);
and U13307 (N_13307,N_12853,N_12757);
or U13308 (N_13308,N_12807,N_12679);
nand U13309 (N_13309,N_12958,N_12936);
or U13310 (N_13310,N_12847,N_12708);
nor U13311 (N_13311,N_12860,N_12900);
and U13312 (N_13312,N_12703,N_12887);
or U13313 (N_13313,N_12745,N_12689);
nor U13314 (N_13314,N_12893,N_12886);
and U13315 (N_13315,N_12791,N_12933);
and U13316 (N_13316,N_12665,N_12856);
or U13317 (N_13317,N_12858,N_12981);
or U13318 (N_13318,N_12869,N_12650);
nor U13319 (N_13319,N_12828,N_12938);
or U13320 (N_13320,N_12756,N_12729);
or U13321 (N_13321,N_12781,N_12660);
nand U13322 (N_13322,N_12744,N_12938);
nand U13323 (N_13323,N_12597,N_12525);
and U13324 (N_13324,N_12715,N_12500);
and U13325 (N_13325,N_12696,N_12731);
and U13326 (N_13326,N_12691,N_12765);
nand U13327 (N_13327,N_12838,N_12617);
or U13328 (N_13328,N_12585,N_12821);
and U13329 (N_13329,N_12669,N_12536);
nor U13330 (N_13330,N_12841,N_12965);
and U13331 (N_13331,N_12642,N_12599);
xor U13332 (N_13332,N_12919,N_12636);
xor U13333 (N_13333,N_12540,N_12562);
xor U13334 (N_13334,N_12993,N_12851);
nand U13335 (N_13335,N_12745,N_12602);
nor U13336 (N_13336,N_12571,N_12652);
nor U13337 (N_13337,N_12531,N_12554);
nand U13338 (N_13338,N_12764,N_12636);
nor U13339 (N_13339,N_12654,N_12759);
nor U13340 (N_13340,N_12757,N_12664);
and U13341 (N_13341,N_12613,N_12544);
or U13342 (N_13342,N_12612,N_12854);
or U13343 (N_13343,N_12621,N_12855);
xnor U13344 (N_13344,N_12782,N_12725);
nand U13345 (N_13345,N_12802,N_12970);
or U13346 (N_13346,N_12861,N_12723);
or U13347 (N_13347,N_12612,N_12564);
nand U13348 (N_13348,N_12947,N_12867);
nor U13349 (N_13349,N_12585,N_12877);
and U13350 (N_13350,N_12979,N_12961);
nand U13351 (N_13351,N_12889,N_12768);
nand U13352 (N_13352,N_12633,N_12566);
or U13353 (N_13353,N_12507,N_12968);
and U13354 (N_13354,N_12548,N_12658);
nor U13355 (N_13355,N_12527,N_12974);
nand U13356 (N_13356,N_12574,N_12649);
nor U13357 (N_13357,N_12902,N_12799);
or U13358 (N_13358,N_12624,N_12918);
nand U13359 (N_13359,N_12821,N_12689);
nand U13360 (N_13360,N_12813,N_12723);
nand U13361 (N_13361,N_12951,N_12572);
nand U13362 (N_13362,N_12951,N_12536);
xor U13363 (N_13363,N_12546,N_12744);
and U13364 (N_13364,N_12786,N_12730);
nor U13365 (N_13365,N_12877,N_12567);
nand U13366 (N_13366,N_12739,N_12673);
nor U13367 (N_13367,N_12542,N_12765);
or U13368 (N_13368,N_12811,N_12797);
or U13369 (N_13369,N_12852,N_12521);
nand U13370 (N_13370,N_12571,N_12836);
or U13371 (N_13371,N_12703,N_12967);
nand U13372 (N_13372,N_12888,N_12908);
nor U13373 (N_13373,N_12713,N_12602);
nor U13374 (N_13374,N_12805,N_12729);
or U13375 (N_13375,N_12720,N_12667);
nor U13376 (N_13376,N_12824,N_12541);
or U13377 (N_13377,N_12686,N_12614);
or U13378 (N_13378,N_12554,N_12708);
or U13379 (N_13379,N_12977,N_12929);
and U13380 (N_13380,N_12746,N_12639);
xor U13381 (N_13381,N_12775,N_12765);
or U13382 (N_13382,N_12984,N_12635);
nand U13383 (N_13383,N_12697,N_12696);
nand U13384 (N_13384,N_12708,N_12537);
nand U13385 (N_13385,N_12509,N_12731);
xnor U13386 (N_13386,N_12971,N_12581);
nor U13387 (N_13387,N_12781,N_12789);
and U13388 (N_13388,N_12519,N_12503);
nand U13389 (N_13389,N_12658,N_12545);
nor U13390 (N_13390,N_12770,N_12573);
nor U13391 (N_13391,N_12783,N_12928);
nand U13392 (N_13392,N_12718,N_12720);
nand U13393 (N_13393,N_12688,N_12593);
or U13394 (N_13394,N_12623,N_12532);
nor U13395 (N_13395,N_12640,N_12857);
nand U13396 (N_13396,N_12655,N_12786);
or U13397 (N_13397,N_12798,N_12606);
nand U13398 (N_13398,N_12645,N_12599);
nor U13399 (N_13399,N_12581,N_12959);
and U13400 (N_13400,N_12669,N_12561);
nor U13401 (N_13401,N_12829,N_12564);
and U13402 (N_13402,N_12925,N_12840);
and U13403 (N_13403,N_12576,N_12995);
or U13404 (N_13404,N_12508,N_12642);
and U13405 (N_13405,N_12857,N_12686);
or U13406 (N_13406,N_12624,N_12717);
or U13407 (N_13407,N_12572,N_12734);
and U13408 (N_13408,N_12725,N_12998);
or U13409 (N_13409,N_12646,N_12709);
and U13410 (N_13410,N_12703,N_12874);
and U13411 (N_13411,N_12986,N_12607);
nand U13412 (N_13412,N_12531,N_12678);
and U13413 (N_13413,N_12664,N_12936);
or U13414 (N_13414,N_12533,N_12615);
nand U13415 (N_13415,N_12531,N_12793);
and U13416 (N_13416,N_12795,N_12620);
or U13417 (N_13417,N_12635,N_12792);
xor U13418 (N_13418,N_12972,N_12877);
nor U13419 (N_13419,N_12702,N_12907);
or U13420 (N_13420,N_12786,N_12753);
nand U13421 (N_13421,N_12532,N_12757);
or U13422 (N_13422,N_12587,N_12698);
nand U13423 (N_13423,N_12738,N_12996);
nand U13424 (N_13424,N_12676,N_12511);
or U13425 (N_13425,N_12586,N_12521);
or U13426 (N_13426,N_12841,N_12519);
xnor U13427 (N_13427,N_12854,N_12984);
or U13428 (N_13428,N_12745,N_12800);
nand U13429 (N_13429,N_12527,N_12666);
nand U13430 (N_13430,N_12643,N_12624);
or U13431 (N_13431,N_12963,N_12972);
nor U13432 (N_13432,N_12970,N_12503);
and U13433 (N_13433,N_12595,N_12728);
or U13434 (N_13434,N_12947,N_12729);
and U13435 (N_13435,N_12522,N_12782);
and U13436 (N_13436,N_12660,N_12871);
or U13437 (N_13437,N_12748,N_12553);
xnor U13438 (N_13438,N_12626,N_12534);
nand U13439 (N_13439,N_12969,N_12821);
and U13440 (N_13440,N_12805,N_12564);
nor U13441 (N_13441,N_12607,N_12834);
nand U13442 (N_13442,N_12519,N_12862);
nor U13443 (N_13443,N_12665,N_12606);
or U13444 (N_13444,N_12663,N_12931);
xnor U13445 (N_13445,N_12616,N_12961);
nor U13446 (N_13446,N_12806,N_12843);
nor U13447 (N_13447,N_12822,N_12624);
nand U13448 (N_13448,N_12886,N_12716);
and U13449 (N_13449,N_12851,N_12633);
and U13450 (N_13450,N_12787,N_12922);
nand U13451 (N_13451,N_12935,N_12832);
or U13452 (N_13452,N_12827,N_12639);
or U13453 (N_13453,N_12572,N_12875);
nor U13454 (N_13454,N_12965,N_12591);
or U13455 (N_13455,N_12626,N_12793);
nand U13456 (N_13456,N_12617,N_12702);
and U13457 (N_13457,N_12733,N_12920);
xnor U13458 (N_13458,N_12506,N_12588);
nor U13459 (N_13459,N_12776,N_12912);
nor U13460 (N_13460,N_12629,N_12503);
or U13461 (N_13461,N_12828,N_12878);
xor U13462 (N_13462,N_12929,N_12850);
xnor U13463 (N_13463,N_12506,N_12904);
and U13464 (N_13464,N_12765,N_12706);
nand U13465 (N_13465,N_12664,N_12580);
nand U13466 (N_13466,N_12876,N_12895);
and U13467 (N_13467,N_12578,N_12538);
nand U13468 (N_13468,N_12859,N_12570);
xnor U13469 (N_13469,N_12912,N_12902);
nand U13470 (N_13470,N_12784,N_12649);
or U13471 (N_13471,N_12549,N_12532);
nand U13472 (N_13472,N_12588,N_12968);
nor U13473 (N_13473,N_12856,N_12800);
or U13474 (N_13474,N_12826,N_12878);
nand U13475 (N_13475,N_12802,N_12880);
or U13476 (N_13476,N_12630,N_12642);
nor U13477 (N_13477,N_12976,N_12933);
nor U13478 (N_13478,N_12784,N_12960);
nand U13479 (N_13479,N_12770,N_12517);
or U13480 (N_13480,N_12940,N_12748);
xor U13481 (N_13481,N_12847,N_12531);
and U13482 (N_13482,N_12699,N_12684);
nand U13483 (N_13483,N_12673,N_12607);
nor U13484 (N_13484,N_12661,N_12910);
or U13485 (N_13485,N_12705,N_12902);
nand U13486 (N_13486,N_12513,N_12922);
nor U13487 (N_13487,N_12977,N_12878);
xnor U13488 (N_13488,N_12629,N_12670);
nand U13489 (N_13489,N_12830,N_12740);
or U13490 (N_13490,N_12741,N_12949);
and U13491 (N_13491,N_12997,N_12570);
xnor U13492 (N_13492,N_12642,N_12533);
nor U13493 (N_13493,N_12928,N_12753);
and U13494 (N_13494,N_12548,N_12999);
or U13495 (N_13495,N_12503,N_12596);
nor U13496 (N_13496,N_12982,N_12695);
and U13497 (N_13497,N_12662,N_12843);
nor U13498 (N_13498,N_12861,N_12590);
or U13499 (N_13499,N_12790,N_12820);
nand U13500 (N_13500,N_13044,N_13447);
nor U13501 (N_13501,N_13056,N_13104);
nor U13502 (N_13502,N_13188,N_13074);
and U13503 (N_13503,N_13351,N_13361);
nor U13504 (N_13504,N_13296,N_13103);
xnor U13505 (N_13505,N_13384,N_13292);
and U13506 (N_13506,N_13346,N_13010);
xor U13507 (N_13507,N_13211,N_13113);
xnor U13508 (N_13508,N_13082,N_13124);
and U13509 (N_13509,N_13043,N_13100);
nand U13510 (N_13510,N_13073,N_13328);
or U13511 (N_13511,N_13051,N_13020);
and U13512 (N_13512,N_13248,N_13404);
xnor U13513 (N_13513,N_13241,N_13161);
or U13514 (N_13514,N_13414,N_13255);
nor U13515 (N_13515,N_13290,N_13186);
and U13516 (N_13516,N_13151,N_13135);
xnor U13517 (N_13517,N_13326,N_13352);
and U13518 (N_13518,N_13286,N_13230);
nor U13519 (N_13519,N_13412,N_13087);
nor U13520 (N_13520,N_13358,N_13386);
nand U13521 (N_13521,N_13185,N_13236);
or U13522 (N_13522,N_13072,N_13029);
and U13523 (N_13523,N_13396,N_13267);
nor U13524 (N_13524,N_13432,N_13116);
nand U13525 (N_13525,N_13148,N_13042);
xnor U13526 (N_13526,N_13395,N_13167);
or U13527 (N_13527,N_13075,N_13122);
nor U13528 (N_13528,N_13277,N_13354);
nand U13529 (N_13529,N_13329,N_13257);
nor U13530 (N_13530,N_13478,N_13136);
and U13531 (N_13531,N_13260,N_13454);
nand U13532 (N_13532,N_13298,N_13037);
or U13533 (N_13533,N_13221,N_13471);
and U13534 (N_13534,N_13439,N_13345);
nand U13535 (N_13535,N_13280,N_13455);
xnor U13536 (N_13536,N_13005,N_13464);
nand U13537 (N_13537,N_13394,N_13406);
nand U13538 (N_13538,N_13275,N_13215);
nand U13539 (N_13539,N_13348,N_13141);
or U13540 (N_13540,N_13233,N_13262);
nor U13541 (N_13541,N_13397,N_13118);
and U13542 (N_13542,N_13295,N_13381);
nand U13543 (N_13543,N_13300,N_13039);
or U13544 (N_13544,N_13067,N_13001);
nor U13545 (N_13545,N_13026,N_13476);
and U13546 (N_13546,N_13377,N_13283);
or U13547 (N_13547,N_13134,N_13330);
xnor U13548 (N_13548,N_13047,N_13227);
nand U13549 (N_13549,N_13387,N_13291);
and U13550 (N_13550,N_13390,N_13278);
xnor U13551 (N_13551,N_13419,N_13425);
nor U13552 (N_13552,N_13190,N_13007);
or U13553 (N_13553,N_13049,N_13362);
and U13554 (N_13554,N_13132,N_13054);
nor U13555 (N_13555,N_13468,N_13111);
and U13556 (N_13556,N_13149,N_13484);
or U13557 (N_13557,N_13415,N_13340);
and U13558 (N_13558,N_13324,N_13426);
nor U13559 (N_13559,N_13120,N_13091);
nand U13560 (N_13560,N_13318,N_13006);
nand U13561 (N_13561,N_13423,N_13025);
and U13562 (N_13562,N_13206,N_13433);
and U13563 (N_13563,N_13107,N_13309);
nand U13564 (N_13564,N_13287,N_13453);
or U13565 (N_13565,N_13182,N_13334);
and U13566 (N_13566,N_13181,N_13071);
or U13567 (N_13567,N_13461,N_13179);
and U13568 (N_13568,N_13360,N_13108);
and U13569 (N_13569,N_13028,N_13140);
xor U13570 (N_13570,N_13163,N_13229);
nand U13571 (N_13571,N_13040,N_13194);
nand U13572 (N_13572,N_13031,N_13207);
or U13573 (N_13573,N_13168,N_13199);
and U13574 (N_13574,N_13183,N_13413);
nand U13575 (N_13575,N_13143,N_13203);
nor U13576 (N_13576,N_13490,N_13033);
and U13577 (N_13577,N_13019,N_13322);
or U13578 (N_13578,N_13353,N_13232);
and U13579 (N_13579,N_13373,N_13385);
and U13580 (N_13580,N_13105,N_13422);
nor U13581 (N_13581,N_13234,N_13223);
nor U13582 (N_13582,N_13115,N_13050);
nand U13583 (N_13583,N_13024,N_13416);
nor U13584 (N_13584,N_13349,N_13251);
nand U13585 (N_13585,N_13237,N_13224);
and U13586 (N_13586,N_13057,N_13070);
and U13587 (N_13587,N_13448,N_13121);
or U13588 (N_13588,N_13469,N_13269);
or U13589 (N_13589,N_13150,N_13171);
nor U13590 (N_13590,N_13158,N_13479);
xor U13591 (N_13591,N_13052,N_13058);
xnor U13592 (N_13592,N_13127,N_13356);
nor U13593 (N_13593,N_13123,N_13247);
or U13594 (N_13594,N_13420,N_13243);
nor U13595 (N_13595,N_13027,N_13078);
and U13596 (N_13596,N_13392,N_13137);
nor U13597 (N_13597,N_13271,N_13041);
nor U13598 (N_13598,N_13289,N_13125);
nand U13599 (N_13599,N_13443,N_13202);
nor U13600 (N_13600,N_13409,N_13189);
and U13601 (N_13601,N_13193,N_13098);
xor U13602 (N_13602,N_13055,N_13184);
nor U13603 (N_13603,N_13284,N_13252);
or U13604 (N_13604,N_13485,N_13378);
and U13605 (N_13605,N_13048,N_13177);
and U13606 (N_13606,N_13314,N_13012);
xnor U13607 (N_13607,N_13210,N_13101);
or U13608 (N_13608,N_13282,N_13154);
nand U13609 (N_13609,N_13458,N_13198);
nand U13610 (N_13610,N_13475,N_13259);
nor U13611 (N_13611,N_13160,N_13117);
or U13612 (N_13612,N_13011,N_13402);
and U13613 (N_13613,N_13445,N_13365);
and U13614 (N_13614,N_13465,N_13488);
xor U13615 (N_13615,N_13312,N_13467);
xnor U13616 (N_13616,N_13305,N_13045);
nor U13617 (N_13617,N_13128,N_13003);
nand U13618 (N_13618,N_13153,N_13350);
nor U13619 (N_13619,N_13090,N_13470);
nor U13620 (N_13620,N_13380,N_13421);
nor U13621 (N_13621,N_13327,N_13133);
or U13622 (N_13622,N_13359,N_13155);
nand U13623 (N_13623,N_13452,N_13459);
nor U13624 (N_13624,N_13323,N_13431);
and U13625 (N_13625,N_13480,N_13173);
or U13626 (N_13626,N_13268,N_13279);
nand U13627 (N_13627,N_13482,N_13273);
nand U13628 (N_13628,N_13144,N_13253);
nand U13629 (N_13629,N_13444,N_13457);
or U13630 (N_13630,N_13331,N_13030);
nand U13631 (N_13631,N_13428,N_13401);
nor U13632 (N_13632,N_13261,N_13342);
or U13633 (N_13633,N_13368,N_13213);
xnor U13634 (N_13634,N_13367,N_13242);
nor U13635 (N_13635,N_13473,N_13493);
or U13636 (N_13636,N_13097,N_13214);
nor U13637 (N_13637,N_13336,N_13366);
nor U13638 (N_13638,N_13440,N_13483);
or U13639 (N_13639,N_13317,N_13166);
nor U13640 (N_13640,N_13313,N_13274);
or U13641 (N_13641,N_13009,N_13270);
or U13642 (N_13642,N_13217,N_13263);
or U13643 (N_13643,N_13303,N_13212);
and U13644 (N_13644,N_13341,N_13398);
xor U13645 (N_13645,N_13172,N_13302);
xor U13646 (N_13646,N_13169,N_13079);
nand U13647 (N_13647,N_13200,N_13126);
and U13648 (N_13648,N_13235,N_13335);
nor U13649 (N_13649,N_13410,N_13060);
and U13650 (N_13650,N_13288,N_13363);
nand U13651 (N_13651,N_13487,N_13429);
or U13652 (N_13652,N_13094,N_13441);
xor U13653 (N_13653,N_13021,N_13080);
or U13654 (N_13654,N_13102,N_13192);
xnor U13655 (N_13655,N_13038,N_13245);
nor U13656 (N_13656,N_13228,N_13156);
or U13657 (N_13657,N_13088,N_13494);
or U13658 (N_13658,N_13053,N_13311);
nor U13659 (N_13659,N_13338,N_13017);
nand U13660 (N_13660,N_13489,N_13015);
and U13661 (N_13661,N_13205,N_13472);
xnor U13662 (N_13662,N_13265,N_13405);
nand U13663 (N_13663,N_13370,N_13254);
nand U13664 (N_13664,N_13063,N_13089);
nand U13665 (N_13665,N_13272,N_13427);
nor U13666 (N_13666,N_13164,N_13065);
nor U13667 (N_13667,N_13142,N_13191);
and U13668 (N_13668,N_13109,N_13276);
and U13669 (N_13669,N_13092,N_13357);
nor U13670 (N_13670,N_13096,N_13308);
and U13671 (N_13671,N_13486,N_13449);
nand U13672 (N_13672,N_13138,N_13446);
or U13673 (N_13673,N_13400,N_13437);
nand U13674 (N_13674,N_13204,N_13481);
nand U13675 (N_13675,N_13337,N_13294);
and U13676 (N_13676,N_13399,N_13496);
and U13677 (N_13677,N_13208,N_13320);
and U13678 (N_13678,N_13466,N_13152);
or U13679 (N_13679,N_13477,N_13339);
nand U13680 (N_13680,N_13299,N_13046);
nor U13681 (N_13681,N_13258,N_13244);
nor U13682 (N_13682,N_13495,N_13371);
nor U13683 (N_13683,N_13424,N_13411);
and U13684 (N_13684,N_13474,N_13226);
or U13685 (N_13685,N_13036,N_13139);
nor U13686 (N_13686,N_13306,N_13375);
nand U13687 (N_13687,N_13246,N_13225);
and U13688 (N_13688,N_13376,N_13013);
and U13689 (N_13689,N_13165,N_13333);
nor U13690 (N_13690,N_13408,N_13238);
or U13691 (N_13691,N_13417,N_13383);
and U13692 (N_13692,N_13372,N_13130);
or U13693 (N_13693,N_13114,N_13180);
and U13694 (N_13694,N_13491,N_13403);
nor U13695 (N_13695,N_13316,N_13176);
or U13696 (N_13696,N_13456,N_13374);
and U13697 (N_13697,N_13321,N_13435);
and U13698 (N_13698,N_13068,N_13196);
or U13699 (N_13699,N_13129,N_13451);
and U13700 (N_13700,N_13066,N_13146);
nand U13701 (N_13701,N_13218,N_13095);
nor U13702 (N_13702,N_13388,N_13059);
or U13703 (N_13703,N_13219,N_13112);
and U13704 (N_13704,N_13239,N_13178);
xnor U13705 (N_13705,N_13016,N_13174);
nand U13706 (N_13706,N_13281,N_13285);
and U13707 (N_13707,N_13389,N_13022);
nor U13708 (N_13708,N_13018,N_13145);
and U13709 (N_13709,N_13023,N_13093);
or U13710 (N_13710,N_13430,N_13301);
and U13711 (N_13711,N_13081,N_13304);
nand U13712 (N_13712,N_13442,N_13460);
or U13713 (N_13713,N_13170,N_13499);
and U13714 (N_13714,N_13084,N_13434);
or U13715 (N_13715,N_13250,N_13034);
and U13716 (N_13716,N_13110,N_13369);
xnor U13717 (N_13717,N_13462,N_13195);
and U13718 (N_13718,N_13187,N_13492);
xor U13719 (N_13719,N_13256,N_13249);
or U13720 (N_13720,N_13355,N_13436);
nor U13721 (N_13721,N_13197,N_13438);
nand U13722 (N_13722,N_13099,N_13014);
nand U13723 (N_13723,N_13216,N_13119);
and U13724 (N_13724,N_13004,N_13498);
nor U13725 (N_13725,N_13220,N_13077);
nand U13726 (N_13726,N_13106,N_13083);
nand U13727 (N_13727,N_13008,N_13000);
or U13728 (N_13728,N_13407,N_13032);
xnor U13729 (N_13729,N_13450,N_13061);
nor U13730 (N_13730,N_13393,N_13315);
nor U13731 (N_13731,N_13307,N_13085);
and U13732 (N_13732,N_13266,N_13344);
nor U13733 (N_13733,N_13240,N_13347);
or U13734 (N_13734,N_13343,N_13201);
xor U13735 (N_13735,N_13497,N_13382);
or U13736 (N_13736,N_13086,N_13131);
or U13737 (N_13737,N_13293,N_13159);
nor U13738 (N_13738,N_13147,N_13222);
or U13739 (N_13739,N_13064,N_13325);
nand U13740 (N_13740,N_13076,N_13175);
xnor U13741 (N_13741,N_13264,N_13319);
and U13742 (N_13742,N_13379,N_13002);
and U13743 (N_13743,N_13162,N_13463);
nand U13744 (N_13744,N_13332,N_13297);
and U13745 (N_13745,N_13391,N_13310);
or U13746 (N_13746,N_13035,N_13364);
and U13747 (N_13747,N_13418,N_13209);
nor U13748 (N_13748,N_13069,N_13231);
nand U13749 (N_13749,N_13157,N_13062);
nor U13750 (N_13750,N_13037,N_13352);
nor U13751 (N_13751,N_13374,N_13385);
nand U13752 (N_13752,N_13290,N_13434);
nor U13753 (N_13753,N_13473,N_13141);
nor U13754 (N_13754,N_13063,N_13111);
nand U13755 (N_13755,N_13190,N_13239);
nor U13756 (N_13756,N_13471,N_13159);
and U13757 (N_13757,N_13170,N_13274);
or U13758 (N_13758,N_13093,N_13459);
nand U13759 (N_13759,N_13469,N_13163);
nand U13760 (N_13760,N_13085,N_13324);
and U13761 (N_13761,N_13249,N_13344);
nand U13762 (N_13762,N_13215,N_13045);
and U13763 (N_13763,N_13364,N_13219);
or U13764 (N_13764,N_13444,N_13371);
or U13765 (N_13765,N_13130,N_13371);
and U13766 (N_13766,N_13196,N_13463);
and U13767 (N_13767,N_13086,N_13025);
and U13768 (N_13768,N_13218,N_13190);
or U13769 (N_13769,N_13320,N_13278);
nor U13770 (N_13770,N_13297,N_13432);
or U13771 (N_13771,N_13077,N_13168);
and U13772 (N_13772,N_13140,N_13224);
and U13773 (N_13773,N_13357,N_13384);
nor U13774 (N_13774,N_13344,N_13454);
nor U13775 (N_13775,N_13449,N_13100);
xnor U13776 (N_13776,N_13162,N_13354);
and U13777 (N_13777,N_13346,N_13077);
nand U13778 (N_13778,N_13340,N_13146);
nor U13779 (N_13779,N_13063,N_13221);
nand U13780 (N_13780,N_13221,N_13034);
and U13781 (N_13781,N_13140,N_13189);
nor U13782 (N_13782,N_13191,N_13001);
nand U13783 (N_13783,N_13182,N_13405);
nor U13784 (N_13784,N_13098,N_13071);
nor U13785 (N_13785,N_13077,N_13405);
nor U13786 (N_13786,N_13050,N_13432);
nand U13787 (N_13787,N_13430,N_13292);
nor U13788 (N_13788,N_13166,N_13059);
or U13789 (N_13789,N_13254,N_13185);
xnor U13790 (N_13790,N_13097,N_13127);
and U13791 (N_13791,N_13220,N_13430);
or U13792 (N_13792,N_13038,N_13280);
nand U13793 (N_13793,N_13352,N_13012);
and U13794 (N_13794,N_13214,N_13125);
xor U13795 (N_13795,N_13242,N_13070);
and U13796 (N_13796,N_13011,N_13115);
nand U13797 (N_13797,N_13029,N_13404);
xnor U13798 (N_13798,N_13385,N_13372);
xor U13799 (N_13799,N_13241,N_13210);
nor U13800 (N_13800,N_13405,N_13129);
or U13801 (N_13801,N_13235,N_13298);
nand U13802 (N_13802,N_13287,N_13250);
and U13803 (N_13803,N_13325,N_13367);
nand U13804 (N_13804,N_13029,N_13001);
or U13805 (N_13805,N_13012,N_13360);
and U13806 (N_13806,N_13248,N_13408);
or U13807 (N_13807,N_13313,N_13496);
nand U13808 (N_13808,N_13134,N_13221);
or U13809 (N_13809,N_13246,N_13232);
nor U13810 (N_13810,N_13336,N_13337);
and U13811 (N_13811,N_13466,N_13267);
nor U13812 (N_13812,N_13187,N_13384);
and U13813 (N_13813,N_13434,N_13028);
nand U13814 (N_13814,N_13063,N_13422);
or U13815 (N_13815,N_13288,N_13007);
and U13816 (N_13816,N_13459,N_13020);
nand U13817 (N_13817,N_13262,N_13263);
nor U13818 (N_13818,N_13457,N_13118);
and U13819 (N_13819,N_13286,N_13052);
xor U13820 (N_13820,N_13200,N_13451);
and U13821 (N_13821,N_13280,N_13124);
nand U13822 (N_13822,N_13108,N_13300);
nand U13823 (N_13823,N_13498,N_13435);
and U13824 (N_13824,N_13499,N_13359);
or U13825 (N_13825,N_13412,N_13437);
nand U13826 (N_13826,N_13011,N_13029);
nor U13827 (N_13827,N_13236,N_13471);
nand U13828 (N_13828,N_13324,N_13298);
or U13829 (N_13829,N_13435,N_13006);
xor U13830 (N_13830,N_13389,N_13153);
nor U13831 (N_13831,N_13152,N_13463);
nand U13832 (N_13832,N_13010,N_13147);
nor U13833 (N_13833,N_13117,N_13071);
and U13834 (N_13834,N_13328,N_13403);
or U13835 (N_13835,N_13300,N_13336);
nor U13836 (N_13836,N_13302,N_13171);
or U13837 (N_13837,N_13200,N_13374);
or U13838 (N_13838,N_13117,N_13037);
or U13839 (N_13839,N_13179,N_13013);
xor U13840 (N_13840,N_13258,N_13343);
and U13841 (N_13841,N_13471,N_13197);
nand U13842 (N_13842,N_13285,N_13044);
nor U13843 (N_13843,N_13331,N_13330);
nand U13844 (N_13844,N_13218,N_13440);
nor U13845 (N_13845,N_13057,N_13477);
xnor U13846 (N_13846,N_13351,N_13349);
nand U13847 (N_13847,N_13450,N_13104);
or U13848 (N_13848,N_13002,N_13237);
nand U13849 (N_13849,N_13033,N_13488);
nor U13850 (N_13850,N_13405,N_13014);
nand U13851 (N_13851,N_13396,N_13268);
and U13852 (N_13852,N_13395,N_13354);
and U13853 (N_13853,N_13441,N_13097);
and U13854 (N_13854,N_13409,N_13165);
and U13855 (N_13855,N_13423,N_13217);
or U13856 (N_13856,N_13361,N_13365);
nor U13857 (N_13857,N_13015,N_13499);
and U13858 (N_13858,N_13397,N_13041);
nor U13859 (N_13859,N_13426,N_13177);
nor U13860 (N_13860,N_13445,N_13101);
nor U13861 (N_13861,N_13011,N_13361);
or U13862 (N_13862,N_13349,N_13354);
and U13863 (N_13863,N_13084,N_13037);
xnor U13864 (N_13864,N_13374,N_13355);
nor U13865 (N_13865,N_13020,N_13436);
nand U13866 (N_13866,N_13032,N_13300);
or U13867 (N_13867,N_13199,N_13126);
xnor U13868 (N_13868,N_13104,N_13044);
nor U13869 (N_13869,N_13001,N_13136);
nand U13870 (N_13870,N_13409,N_13153);
nand U13871 (N_13871,N_13032,N_13235);
or U13872 (N_13872,N_13488,N_13227);
nand U13873 (N_13873,N_13409,N_13201);
nor U13874 (N_13874,N_13464,N_13048);
or U13875 (N_13875,N_13007,N_13151);
and U13876 (N_13876,N_13240,N_13219);
or U13877 (N_13877,N_13235,N_13213);
nor U13878 (N_13878,N_13252,N_13416);
nand U13879 (N_13879,N_13454,N_13077);
nand U13880 (N_13880,N_13398,N_13090);
or U13881 (N_13881,N_13381,N_13402);
nor U13882 (N_13882,N_13370,N_13313);
and U13883 (N_13883,N_13086,N_13264);
nor U13884 (N_13884,N_13143,N_13389);
and U13885 (N_13885,N_13055,N_13316);
nand U13886 (N_13886,N_13368,N_13420);
and U13887 (N_13887,N_13234,N_13153);
and U13888 (N_13888,N_13321,N_13028);
nor U13889 (N_13889,N_13481,N_13440);
nor U13890 (N_13890,N_13298,N_13188);
nand U13891 (N_13891,N_13382,N_13402);
and U13892 (N_13892,N_13195,N_13232);
and U13893 (N_13893,N_13080,N_13124);
nor U13894 (N_13894,N_13110,N_13004);
xor U13895 (N_13895,N_13479,N_13126);
nand U13896 (N_13896,N_13237,N_13154);
nand U13897 (N_13897,N_13034,N_13117);
nand U13898 (N_13898,N_13446,N_13367);
and U13899 (N_13899,N_13116,N_13490);
xor U13900 (N_13900,N_13437,N_13391);
nand U13901 (N_13901,N_13121,N_13317);
xor U13902 (N_13902,N_13348,N_13219);
nand U13903 (N_13903,N_13086,N_13318);
or U13904 (N_13904,N_13322,N_13084);
or U13905 (N_13905,N_13422,N_13019);
nand U13906 (N_13906,N_13485,N_13406);
nand U13907 (N_13907,N_13172,N_13459);
and U13908 (N_13908,N_13160,N_13312);
xor U13909 (N_13909,N_13041,N_13455);
and U13910 (N_13910,N_13418,N_13260);
or U13911 (N_13911,N_13272,N_13218);
nor U13912 (N_13912,N_13430,N_13205);
nor U13913 (N_13913,N_13423,N_13268);
nor U13914 (N_13914,N_13084,N_13047);
or U13915 (N_13915,N_13447,N_13421);
nor U13916 (N_13916,N_13233,N_13212);
nor U13917 (N_13917,N_13055,N_13336);
or U13918 (N_13918,N_13484,N_13071);
nand U13919 (N_13919,N_13482,N_13371);
and U13920 (N_13920,N_13024,N_13088);
nand U13921 (N_13921,N_13433,N_13306);
or U13922 (N_13922,N_13354,N_13418);
and U13923 (N_13923,N_13465,N_13280);
and U13924 (N_13924,N_13124,N_13285);
nand U13925 (N_13925,N_13044,N_13020);
xnor U13926 (N_13926,N_13072,N_13452);
or U13927 (N_13927,N_13082,N_13192);
nor U13928 (N_13928,N_13353,N_13082);
xor U13929 (N_13929,N_13311,N_13494);
nor U13930 (N_13930,N_13202,N_13216);
nand U13931 (N_13931,N_13080,N_13461);
and U13932 (N_13932,N_13205,N_13320);
nand U13933 (N_13933,N_13057,N_13196);
xor U13934 (N_13934,N_13011,N_13420);
nand U13935 (N_13935,N_13377,N_13290);
nand U13936 (N_13936,N_13064,N_13357);
or U13937 (N_13937,N_13026,N_13042);
nor U13938 (N_13938,N_13289,N_13187);
nand U13939 (N_13939,N_13499,N_13013);
and U13940 (N_13940,N_13379,N_13331);
nor U13941 (N_13941,N_13478,N_13342);
nand U13942 (N_13942,N_13274,N_13216);
nand U13943 (N_13943,N_13291,N_13258);
and U13944 (N_13944,N_13279,N_13073);
and U13945 (N_13945,N_13337,N_13008);
and U13946 (N_13946,N_13321,N_13042);
and U13947 (N_13947,N_13295,N_13393);
and U13948 (N_13948,N_13157,N_13219);
nor U13949 (N_13949,N_13408,N_13001);
nand U13950 (N_13950,N_13161,N_13352);
nand U13951 (N_13951,N_13228,N_13012);
nand U13952 (N_13952,N_13157,N_13355);
and U13953 (N_13953,N_13016,N_13341);
xor U13954 (N_13954,N_13392,N_13482);
nand U13955 (N_13955,N_13291,N_13158);
nand U13956 (N_13956,N_13364,N_13187);
nor U13957 (N_13957,N_13451,N_13403);
nor U13958 (N_13958,N_13171,N_13223);
nor U13959 (N_13959,N_13322,N_13364);
nand U13960 (N_13960,N_13348,N_13385);
xor U13961 (N_13961,N_13265,N_13234);
or U13962 (N_13962,N_13335,N_13406);
or U13963 (N_13963,N_13381,N_13468);
nor U13964 (N_13964,N_13317,N_13355);
or U13965 (N_13965,N_13460,N_13335);
or U13966 (N_13966,N_13156,N_13393);
and U13967 (N_13967,N_13359,N_13137);
nor U13968 (N_13968,N_13318,N_13140);
and U13969 (N_13969,N_13166,N_13301);
nor U13970 (N_13970,N_13465,N_13037);
nand U13971 (N_13971,N_13288,N_13021);
and U13972 (N_13972,N_13410,N_13201);
or U13973 (N_13973,N_13216,N_13222);
xnor U13974 (N_13974,N_13057,N_13420);
nor U13975 (N_13975,N_13269,N_13211);
or U13976 (N_13976,N_13231,N_13235);
nor U13977 (N_13977,N_13101,N_13369);
nand U13978 (N_13978,N_13478,N_13430);
or U13979 (N_13979,N_13370,N_13448);
or U13980 (N_13980,N_13492,N_13226);
and U13981 (N_13981,N_13474,N_13104);
or U13982 (N_13982,N_13084,N_13122);
or U13983 (N_13983,N_13351,N_13299);
nand U13984 (N_13984,N_13273,N_13246);
or U13985 (N_13985,N_13267,N_13132);
nor U13986 (N_13986,N_13311,N_13466);
or U13987 (N_13987,N_13043,N_13129);
nand U13988 (N_13988,N_13464,N_13074);
and U13989 (N_13989,N_13366,N_13300);
nand U13990 (N_13990,N_13130,N_13233);
nand U13991 (N_13991,N_13187,N_13407);
or U13992 (N_13992,N_13222,N_13405);
and U13993 (N_13993,N_13092,N_13457);
or U13994 (N_13994,N_13162,N_13192);
nor U13995 (N_13995,N_13029,N_13295);
nor U13996 (N_13996,N_13451,N_13182);
or U13997 (N_13997,N_13461,N_13392);
xor U13998 (N_13998,N_13100,N_13444);
and U13999 (N_13999,N_13211,N_13383);
or U14000 (N_14000,N_13777,N_13856);
or U14001 (N_14001,N_13647,N_13829);
and U14002 (N_14002,N_13764,N_13742);
nand U14003 (N_14003,N_13760,N_13666);
nand U14004 (N_14004,N_13553,N_13757);
nor U14005 (N_14005,N_13565,N_13785);
and U14006 (N_14006,N_13986,N_13802);
or U14007 (N_14007,N_13720,N_13899);
xnor U14008 (N_14008,N_13937,N_13705);
or U14009 (N_14009,N_13660,N_13828);
nor U14010 (N_14010,N_13509,N_13637);
xnor U14011 (N_14011,N_13722,N_13741);
or U14012 (N_14012,N_13568,N_13857);
and U14013 (N_14013,N_13896,N_13706);
or U14014 (N_14014,N_13795,N_13580);
or U14015 (N_14015,N_13906,N_13767);
and U14016 (N_14016,N_13863,N_13933);
or U14017 (N_14017,N_13999,N_13745);
or U14018 (N_14018,N_13578,N_13679);
and U14019 (N_14019,N_13729,N_13934);
nand U14020 (N_14020,N_13938,N_13738);
or U14021 (N_14021,N_13880,N_13608);
and U14022 (N_14022,N_13525,N_13836);
nor U14023 (N_14023,N_13981,N_13617);
and U14024 (N_14024,N_13844,N_13708);
or U14025 (N_14025,N_13774,N_13547);
nand U14026 (N_14026,N_13710,N_13854);
nor U14027 (N_14027,N_13630,N_13895);
nor U14028 (N_14028,N_13675,N_13588);
nor U14029 (N_14029,N_13585,N_13668);
or U14030 (N_14030,N_13589,N_13945);
nand U14031 (N_14031,N_13766,N_13761);
or U14032 (N_14032,N_13622,N_13826);
nand U14033 (N_14033,N_13544,N_13909);
or U14034 (N_14034,N_13918,N_13871);
nor U14035 (N_14035,N_13897,N_13733);
nand U14036 (N_14036,N_13979,N_13626);
nor U14037 (N_14037,N_13614,N_13878);
or U14038 (N_14038,N_13845,N_13859);
nor U14039 (N_14039,N_13935,N_13962);
and U14040 (N_14040,N_13913,N_13646);
or U14041 (N_14041,N_13638,N_13961);
and U14042 (N_14042,N_13590,N_13743);
nand U14043 (N_14043,N_13873,N_13567);
nor U14044 (N_14044,N_13876,N_13649);
nand U14045 (N_14045,N_13592,N_13692);
nand U14046 (N_14046,N_13855,N_13701);
or U14047 (N_14047,N_13877,N_13858);
xor U14048 (N_14048,N_13573,N_13519);
or U14049 (N_14049,N_13950,N_13967);
xnor U14050 (N_14050,N_13786,N_13531);
and U14051 (N_14051,N_13542,N_13618);
nor U14052 (N_14052,N_13992,N_13921);
or U14053 (N_14053,N_13684,N_13534);
and U14054 (N_14054,N_13651,N_13699);
nor U14055 (N_14055,N_13557,N_13794);
and U14056 (N_14056,N_13540,N_13968);
xnor U14057 (N_14057,N_13615,N_13515);
nor U14058 (N_14058,N_13511,N_13672);
or U14059 (N_14059,N_13572,N_13922);
and U14060 (N_14060,N_13719,N_13521);
or U14061 (N_14061,N_13532,N_13582);
nor U14062 (N_14062,N_13984,N_13656);
nor U14063 (N_14063,N_13955,N_13690);
or U14064 (N_14064,N_13972,N_13975);
nand U14065 (N_14065,N_13814,N_13905);
nor U14066 (N_14066,N_13714,N_13529);
and U14067 (N_14067,N_13587,N_13505);
nand U14068 (N_14068,N_13610,N_13591);
nand U14069 (N_14069,N_13611,N_13623);
nand U14070 (N_14070,N_13885,N_13987);
or U14071 (N_14071,N_13792,N_13954);
xor U14072 (N_14072,N_13550,N_13537);
xor U14073 (N_14073,N_13797,N_13980);
xnor U14074 (N_14074,N_13601,N_13867);
or U14075 (N_14075,N_13793,N_13772);
xor U14076 (N_14076,N_13998,N_13847);
and U14077 (N_14077,N_13700,N_13953);
and U14078 (N_14078,N_13951,N_13846);
nand U14079 (N_14079,N_13809,N_13508);
nand U14080 (N_14080,N_13883,N_13513);
nor U14081 (N_14081,N_13518,N_13890);
and U14082 (N_14082,N_13501,N_13594);
or U14083 (N_14083,N_13503,N_13816);
and U14084 (N_14084,N_13898,N_13801);
nand U14085 (N_14085,N_13579,N_13747);
or U14086 (N_14086,N_13755,N_13609);
nor U14087 (N_14087,N_13778,N_13969);
or U14088 (N_14088,N_13527,N_13657);
nand U14089 (N_14089,N_13990,N_13832);
and U14090 (N_14090,N_13596,N_13759);
nand U14091 (N_14091,N_13948,N_13841);
nand U14092 (N_14092,N_13732,N_13808);
nor U14093 (N_14093,N_13686,N_13650);
and U14094 (N_14094,N_13944,N_13908);
or U14095 (N_14095,N_13824,N_13868);
nor U14096 (N_14096,N_13512,N_13667);
nor U14097 (N_14097,N_13533,N_13754);
xor U14098 (N_14098,N_13973,N_13887);
or U14099 (N_14099,N_13516,N_13976);
or U14100 (N_14100,N_13932,N_13566);
or U14101 (N_14101,N_13718,N_13558);
xnor U14102 (N_14102,N_13703,N_13555);
and U14103 (N_14103,N_13655,N_13597);
nand U14104 (N_14104,N_13691,N_13731);
or U14105 (N_14105,N_13715,N_13886);
nand U14106 (N_14106,N_13506,N_13983);
and U14107 (N_14107,N_13966,N_13612);
and U14108 (N_14108,N_13977,N_13765);
and U14109 (N_14109,N_13561,N_13571);
nor U14110 (N_14110,N_13843,N_13923);
and U14111 (N_14111,N_13734,N_13861);
nand U14112 (N_14112,N_13822,N_13598);
and U14113 (N_14113,N_13924,N_13996);
or U14114 (N_14114,N_13600,N_13864);
nor U14115 (N_14115,N_13919,N_13834);
nor U14116 (N_14116,N_13744,N_13997);
nand U14117 (N_14117,N_13978,N_13952);
nand U14118 (N_14118,N_13548,N_13763);
and U14119 (N_14119,N_13685,N_13891);
and U14120 (N_14120,N_13904,N_13881);
or U14121 (N_14121,N_13627,N_13842);
nor U14122 (N_14122,N_13549,N_13709);
or U14123 (N_14123,N_13963,N_13974);
nand U14124 (N_14124,N_13912,N_13697);
or U14125 (N_14125,N_13957,N_13749);
and U14126 (N_14126,N_13993,N_13640);
nand U14127 (N_14127,N_13889,N_13903);
or U14128 (N_14128,N_13599,N_13639);
nand U14129 (N_14129,N_13631,N_13752);
nor U14130 (N_14130,N_13524,N_13835);
and U14131 (N_14131,N_13804,N_13581);
and U14132 (N_14132,N_13791,N_13616);
nand U14133 (N_14133,N_13546,N_13798);
nor U14134 (N_14134,N_13652,N_13702);
nor U14135 (N_14135,N_13676,N_13624);
and U14136 (N_14136,N_13874,N_13815);
and U14137 (N_14137,N_13860,N_13964);
nor U14138 (N_14138,N_13504,N_13787);
nor U14139 (N_14139,N_13807,N_13959);
nand U14140 (N_14140,N_13717,N_13607);
xor U14141 (N_14141,N_13569,N_13852);
or U14142 (N_14142,N_13751,N_13730);
nor U14143 (N_14143,N_13748,N_13989);
nand U14144 (N_14144,N_13879,N_13539);
nand U14145 (N_14145,N_13910,N_13570);
nand U14146 (N_14146,N_13613,N_13817);
and U14147 (N_14147,N_13696,N_13551);
or U14148 (N_14148,N_13872,N_13949);
or U14149 (N_14149,N_13773,N_13894);
nor U14150 (N_14150,N_13595,N_13819);
nor U14151 (N_14151,N_13769,N_13812);
and U14152 (N_14152,N_13716,N_13888);
nand U14153 (N_14153,N_13866,N_13528);
nand U14154 (N_14154,N_13522,N_13543);
nor U14155 (N_14155,N_13633,N_13634);
and U14156 (N_14156,N_13711,N_13625);
or U14157 (N_14157,N_13689,N_13712);
and U14158 (N_14158,N_13849,N_13507);
or U14159 (N_14159,N_13870,N_13960);
or U14160 (N_14160,N_13982,N_13830);
or U14161 (N_14161,N_13673,N_13810);
or U14162 (N_14162,N_13917,N_13771);
nor U14163 (N_14163,N_13662,N_13784);
and U14164 (N_14164,N_13707,N_13768);
and U14165 (N_14165,N_13510,N_13929);
nor U14166 (N_14166,N_13928,N_13671);
and U14167 (N_14167,N_13915,N_13838);
or U14168 (N_14168,N_13837,N_13688);
and U14169 (N_14169,N_13818,N_13682);
and U14170 (N_14170,N_13704,N_13593);
or U14171 (N_14171,N_13602,N_13931);
and U14172 (N_14172,N_13514,N_13994);
nor U14173 (N_14173,N_13827,N_13869);
or U14174 (N_14174,N_13723,N_13674);
nand U14175 (N_14175,N_13781,N_13942);
nor U14176 (N_14176,N_13681,N_13645);
nor U14177 (N_14177,N_13737,N_13806);
nand U14178 (N_14178,N_13940,N_13517);
xnor U14179 (N_14179,N_13776,N_13805);
or U14180 (N_14180,N_13677,N_13939);
xnor U14181 (N_14181,N_13821,N_13713);
or U14182 (N_14182,N_13750,N_13739);
or U14183 (N_14183,N_13621,N_13853);
and U14184 (N_14184,N_13619,N_13559);
nor U14185 (N_14185,N_13520,N_13564);
nor U14186 (N_14186,N_13831,N_13694);
xor U14187 (N_14187,N_13523,N_13995);
nand U14188 (N_14188,N_13563,N_13925);
nor U14189 (N_14189,N_13862,N_13728);
nor U14190 (N_14190,N_13991,N_13892);
nor U14191 (N_14191,N_13965,N_13556);
xnor U14192 (N_14192,N_13800,N_13782);
nor U14193 (N_14193,N_13893,N_13687);
xor U14194 (N_14194,N_13670,N_13648);
nand U14195 (N_14195,N_13985,N_13916);
nor U14196 (N_14196,N_13902,N_13783);
nand U14197 (N_14197,N_13721,N_13538);
nand U14198 (N_14198,N_13663,N_13927);
or U14199 (N_14199,N_13988,N_13636);
or U14200 (N_14200,N_13605,N_13698);
or U14201 (N_14201,N_13583,N_13604);
nand U14202 (N_14202,N_13628,N_13606);
nand U14203 (N_14203,N_13669,N_13574);
xor U14204 (N_14204,N_13775,N_13920);
or U14205 (N_14205,N_13643,N_13536);
nand U14206 (N_14206,N_13658,N_13803);
nand U14207 (N_14207,N_13644,N_13552);
nor U14208 (N_14208,N_13735,N_13840);
and U14209 (N_14209,N_13825,N_13926);
xnor U14210 (N_14210,N_13661,N_13653);
nand U14211 (N_14211,N_13884,N_13839);
or U14212 (N_14212,N_13641,N_13820);
and U14213 (N_14213,N_13746,N_13577);
nor U14214 (N_14214,N_13535,N_13813);
nand U14215 (N_14215,N_13789,N_13758);
or U14216 (N_14216,N_13753,N_13725);
nand U14217 (N_14217,N_13654,N_13848);
nor U14218 (N_14218,N_13500,N_13882);
and U14219 (N_14219,N_13545,N_13664);
nand U14220 (N_14220,N_13788,N_13823);
nand U14221 (N_14221,N_13683,N_13680);
xor U14222 (N_14222,N_13900,N_13629);
xnor U14223 (N_14223,N_13620,N_13541);
nor U14224 (N_14224,N_13770,N_13736);
nand U14225 (N_14225,N_13554,N_13956);
nor U14226 (N_14226,N_13941,N_13875);
and U14227 (N_14227,N_13901,N_13811);
and U14228 (N_14228,N_13632,N_13865);
nand U14229 (N_14229,N_13851,N_13693);
nor U14230 (N_14230,N_13946,N_13796);
nand U14231 (N_14231,N_13943,N_13576);
and U14232 (N_14232,N_13726,N_13678);
nand U14233 (N_14233,N_13586,N_13659);
nand U14234 (N_14234,N_13850,N_13575);
nand U14235 (N_14235,N_13936,N_13780);
nor U14236 (N_14236,N_13560,N_13724);
and U14237 (N_14237,N_13970,N_13584);
nor U14238 (N_14238,N_13502,N_13914);
or U14239 (N_14239,N_13790,N_13695);
or U14240 (N_14240,N_13642,N_13762);
nor U14241 (N_14241,N_13833,N_13911);
or U14242 (N_14242,N_13740,N_13727);
or U14243 (N_14243,N_13603,N_13799);
or U14244 (N_14244,N_13930,N_13526);
and U14245 (N_14245,N_13907,N_13947);
or U14246 (N_14246,N_13971,N_13562);
and U14247 (N_14247,N_13779,N_13756);
nand U14248 (N_14248,N_13635,N_13958);
nor U14249 (N_14249,N_13665,N_13530);
nand U14250 (N_14250,N_13930,N_13824);
nor U14251 (N_14251,N_13860,N_13545);
nand U14252 (N_14252,N_13831,N_13997);
nor U14253 (N_14253,N_13606,N_13709);
nor U14254 (N_14254,N_13583,N_13597);
or U14255 (N_14255,N_13811,N_13569);
nor U14256 (N_14256,N_13819,N_13949);
nor U14257 (N_14257,N_13526,N_13568);
and U14258 (N_14258,N_13912,N_13699);
nand U14259 (N_14259,N_13807,N_13871);
and U14260 (N_14260,N_13568,N_13749);
xor U14261 (N_14261,N_13611,N_13698);
nor U14262 (N_14262,N_13714,N_13643);
nor U14263 (N_14263,N_13598,N_13791);
or U14264 (N_14264,N_13549,N_13962);
and U14265 (N_14265,N_13853,N_13644);
nor U14266 (N_14266,N_13527,N_13991);
and U14267 (N_14267,N_13669,N_13809);
and U14268 (N_14268,N_13760,N_13989);
nand U14269 (N_14269,N_13768,N_13751);
and U14270 (N_14270,N_13730,N_13674);
or U14271 (N_14271,N_13681,N_13864);
xor U14272 (N_14272,N_13558,N_13680);
and U14273 (N_14273,N_13828,N_13801);
nor U14274 (N_14274,N_13594,N_13615);
nor U14275 (N_14275,N_13731,N_13689);
and U14276 (N_14276,N_13516,N_13562);
nand U14277 (N_14277,N_13599,N_13576);
xor U14278 (N_14278,N_13911,N_13596);
or U14279 (N_14279,N_13503,N_13945);
and U14280 (N_14280,N_13863,N_13914);
nor U14281 (N_14281,N_13654,N_13709);
nand U14282 (N_14282,N_13748,N_13661);
nor U14283 (N_14283,N_13941,N_13980);
nor U14284 (N_14284,N_13909,N_13570);
or U14285 (N_14285,N_13997,N_13651);
nor U14286 (N_14286,N_13631,N_13962);
nor U14287 (N_14287,N_13775,N_13602);
nor U14288 (N_14288,N_13754,N_13882);
nand U14289 (N_14289,N_13904,N_13667);
or U14290 (N_14290,N_13832,N_13530);
and U14291 (N_14291,N_13617,N_13792);
nor U14292 (N_14292,N_13652,N_13574);
nand U14293 (N_14293,N_13592,N_13992);
and U14294 (N_14294,N_13971,N_13657);
nand U14295 (N_14295,N_13624,N_13882);
nor U14296 (N_14296,N_13503,N_13756);
nand U14297 (N_14297,N_13513,N_13681);
or U14298 (N_14298,N_13742,N_13848);
nand U14299 (N_14299,N_13914,N_13930);
and U14300 (N_14300,N_13836,N_13756);
xor U14301 (N_14301,N_13824,N_13760);
nor U14302 (N_14302,N_13928,N_13582);
nand U14303 (N_14303,N_13713,N_13621);
and U14304 (N_14304,N_13881,N_13850);
nor U14305 (N_14305,N_13540,N_13800);
or U14306 (N_14306,N_13703,N_13562);
or U14307 (N_14307,N_13795,N_13978);
nand U14308 (N_14308,N_13646,N_13912);
or U14309 (N_14309,N_13973,N_13847);
and U14310 (N_14310,N_13761,N_13660);
nor U14311 (N_14311,N_13844,N_13531);
nor U14312 (N_14312,N_13671,N_13921);
and U14313 (N_14313,N_13636,N_13678);
or U14314 (N_14314,N_13872,N_13833);
xnor U14315 (N_14315,N_13562,N_13796);
nor U14316 (N_14316,N_13976,N_13699);
nor U14317 (N_14317,N_13772,N_13663);
nor U14318 (N_14318,N_13973,N_13786);
nand U14319 (N_14319,N_13973,N_13597);
and U14320 (N_14320,N_13502,N_13606);
or U14321 (N_14321,N_13684,N_13832);
nor U14322 (N_14322,N_13540,N_13715);
nor U14323 (N_14323,N_13592,N_13544);
nand U14324 (N_14324,N_13917,N_13755);
nand U14325 (N_14325,N_13751,N_13876);
and U14326 (N_14326,N_13892,N_13511);
xnor U14327 (N_14327,N_13933,N_13864);
nand U14328 (N_14328,N_13696,N_13929);
and U14329 (N_14329,N_13948,N_13975);
nand U14330 (N_14330,N_13900,N_13866);
or U14331 (N_14331,N_13950,N_13678);
xor U14332 (N_14332,N_13921,N_13633);
or U14333 (N_14333,N_13609,N_13546);
nand U14334 (N_14334,N_13815,N_13645);
or U14335 (N_14335,N_13938,N_13838);
and U14336 (N_14336,N_13643,N_13646);
nor U14337 (N_14337,N_13931,N_13588);
or U14338 (N_14338,N_13710,N_13513);
nand U14339 (N_14339,N_13918,N_13630);
and U14340 (N_14340,N_13664,N_13919);
nand U14341 (N_14341,N_13595,N_13524);
and U14342 (N_14342,N_13964,N_13710);
and U14343 (N_14343,N_13789,N_13946);
nand U14344 (N_14344,N_13768,N_13611);
nand U14345 (N_14345,N_13900,N_13715);
nor U14346 (N_14346,N_13682,N_13586);
xor U14347 (N_14347,N_13988,N_13983);
and U14348 (N_14348,N_13536,N_13773);
nand U14349 (N_14349,N_13552,N_13861);
and U14350 (N_14350,N_13959,N_13798);
and U14351 (N_14351,N_13924,N_13720);
nor U14352 (N_14352,N_13819,N_13549);
nor U14353 (N_14353,N_13930,N_13631);
or U14354 (N_14354,N_13867,N_13880);
and U14355 (N_14355,N_13739,N_13782);
nand U14356 (N_14356,N_13815,N_13871);
xnor U14357 (N_14357,N_13789,N_13726);
xnor U14358 (N_14358,N_13937,N_13671);
nor U14359 (N_14359,N_13959,N_13861);
and U14360 (N_14360,N_13688,N_13619);
xnor U14361 (N_14361,N_13678,N_13550);
nand U14362 (N_14362,N_13969,N_13691);
nor U14363 (N_14363,N_13787,N_13507);
or U14364 (N_14364,N_13768,N_13565);
xnor U14365 (N_14365,N_13529,N_13841);
and U14366 (N_14366,N_13786,N_13673);
nand U14367 (N_14367,N_13794,N_13879);
nand U14368 (N_14368,N_13826,N_13805);
nor U14369 (N_14369,N_13829,N_13826);
or U14370 (N_14370,N_13768,N_13998);
nand U14371 (N_14371,N_13674,N_13529);
nand U14372 (N_14372,N_13709,N_13991);
or U14373 (N_14373,N_13526,N_13703);
and U14374 (N_14374,N_13949,N_13531);
or U14375 (N_14375,N_13976,N_13778);
xnor U14376 (N_14376,N_13887,N_13565);
nor U14377 (N_14377,N_13505,N_13889);
nor U14378 (N_14378,N_13716,N_13624);
and U14379 (N_14379,N_13866,N_13815);
nand U14380 (N_14380,N_13534,N_13735);
and U14381 (N_14381,N_13885,N_13973);
or U14382 (N_14382,N_13867,N_13617);
and U14383 (N_14383,N_13808,N_13962);
nand U14384 (N_14384,N_13705,N_13538);
or U14385 (N_14385,N_13747,N_13613);
nand U14386 (N_14386,N_13880,N_13574);
nor U14387 (N_14387,N_13671,N_13578);
nand U14388 (N_14388,N_13837,N_13730);
or U14389 (N_14389,N_13582,N_13631);
nor U14390 (N_14390,N_13627,N_13883);
or U14391 (N_14391,N_13621,N_13953);
or U14392 (N_14392,N_13966,N_13741);
nand U14393 (N_14393,N_13542,N_13597);
and U14394 (N_14394,N_13621,N_13973);
nand U14395 (N_14395,N_13797,N_13605);
and U14396 (N_14396,N_13852,N_13553);
or U14397 (N_14397,N_13573,N_13693);
nand U14398 (N_14398,N_13525,N_13568);
nor U14399 (N_14399,N_13906,N_13534);
and U14400 (N_14400,N_13940,N_13858);
or U14401 (N_14401,N_13591,N_13986);
nor U14402 (N_14402,N_13948,N_13984);
nand U14403 (N_14403,N_13873,N_13539);
and U14404 (N_14404,N_13742,N_13535);
xor U14405 (N_14405,N_13561,N_13917);
or U14406 (N_14406,N_13849,N_13639);
nand U14407 (N_14407,N_13747,N_13639);
nor U14408 (N_14408,N_13614,N_13697);
or U14409 (N_14409,N_13944,N_13771);
and U14410 (N_14410,N_13781,N_13769);
or U14411 (N_14411,N_13904,N_13575);
nand U14412 (N_14412,N_13679,N_13777);
nor U14413 (N_14413,N_13588,N_13821);
and U14414 (N_14414,N_13621,N_13826);
nor U14415 (N_14415,N_13613,N_13617);
nand U14416 (N_14416,N_13556,N_13558);
nor U14417 (N_14417,N_13756,N_13516);
and U14418 (N_14418,N_13885,N_13994);
or U14419 (N_14419,N_13624,N_13514);
nor U14420 (N_14420,N_13907,N_13890);
and U14421 (N_14421,N_13670,N_13964);
nor U14422 (N_14422,N_13643,N_13742);
or U14423 (N_14423,N_13782,N_13533);
nand U14424 (N_14424,N_13521,N_13535);
nand U14425 (N_14425,N_13509,N_13844);
nand U14426 (N_14426,N_13818,N_13524);
and U14427 (N_14427,N_13532,N_13955);
and U14428 (N_14428,N_13828,N_13887);
nor U14429 (N_14429,N_13576,N_13543);
or U14430 (N_14430,N_13567,N_13915);
and U14431 (N_14431,N_13652,N_13618);
nand U14432 (N_14432,N_13585,N_13721);
or U14433 (N_14433,N_13953,N_13607);
and U14434 (N_14434,N_13608,N_13999);
and U14435 (N_14435,N_13666,N_13926);
or U14436 (N_14436,N_13668,N_13705);
nor U14437 (N_14437,N_13984,N_13844);
and U14438 (N_14438,N_13627,N_13833);
nand U14439 (N_14439,N_13877,N_13730);
or U14440 (N_14440,N_13970,N_13837);
nor U14441 (N_14441,N_13503,N_13780);
or U14442 (N_14442,N_13766,N_13838);
or U14443 (N_14443,N_13982,N_13841);
or U14444 (N_14444,N_13828,N_13861);
and U14445 (N_14445,N_13637,N_13784);
nand U14446 (N_14446,N_13523,N_13839);
xor U14447 (N_14447,N_13564,N_13765);
nand U14448 (N_14448,N_13910,N_13759);
and U14449 (N_14449,N_13511,N_13853);
or U14450 (N_14450,N_13749,N_13757);
and U14451 (N_14451,N_13794,N_13509);
xnor U14452 (N_14452,N_13867,N_13500);
nor U14453 (N_14453,N_13974,N_13835);
or U14454 (N_14454,N_13937,N_13616);
nand U14455 (N_14455,N_13911,N_13840);
nand U14456 (N_14456,N_13623,N_13505);
nand U14457 (N_14457,N_13646,N_13677);
and U14458 (N_14458,N_13857,N_13973);
or U14459 (N_14459,N_13898,N_13906);
xnor U14460 (N_14460,N_13778,N_13612);
or U14461 (N_14461,N_13941,N_13862);
nand U14462 (N_14462,N_13794,N_13715);
or U14463 (N_14463,N_13523,N_13585);
nand U14464 (N_14464,N_13861,N_13772);
and U14465 (N_14465,N_13845,N_13783);
or U14466 (N_14466,N_13577,N_13749);
nand U14467 (N_14467,N_13871,N_13597);
xnor U14468 (N_14468,N_13598,N_13568);
nand U14469 (N_14469,N_13576,N_13911);
nor U14470 (N_14470,N_13963,N_13720);
or U14471 (N_14471,N_13739,N_13942);
nor U14472 (N_14472,N_13846,N_13705);
and U14473 (N_14473,N_13801,N_13577);
nor U14474 (N_14474,N_13502,N_13508);
nor U14475 (N_14475,N_13880,N_13809);
nand U14476 (N_14476,N_13589,N_13775);
or U14477 (N_14477,N_13703,N_13505);
xnor U14478 (N_14478,N_13594,N_13931);
and U14479 (N_14479,N_13647,N_13783);
nand U14480 (N_14480,N_13668,N_13819);
nand U14481 (N_14481,N_13674,N_13938);
xor U14482 (N_14482,N_13936,N_13980);
or U14483 (N_14483,N_13993,N_13560);
xnor U14484 (N_14484,N_13691,N_13902);
nand U14485 (N_14485,N_13635,N_13819);
or U14486 (N_14486,N_13935,N_13528);
nand U14487 (N_14487,N_13824,N_13570);
nand U14488 (N_14488,N_13734,N_13664);
nand U14489 (N_14489,N_13930,N_13565);
nor U14490 (N_14490,N_13979,N_13782);
nand U14491 (N_14491,N_13740,N_13615);
nor U14492 (N_14492,N_13670,N_13868);
nor U14493 (N_14493,N_13714,N_13718);
nand U14494 (N_14494,N_13664,N_13746);
or U14495 (N_14495,N_13554,N_13582);
nor U14496 (N_14496,N_13689,N_13870);
nand U14497 (N_14497,N_13887,N_13538);
nor U14498 (N_14498,N_13834,N_13669);
or U14499 (N_14499,N_13856,N_13548);
xor U14500 (N_14500,N_14140,N_14004);
nor U14501 (N_14501,N_14229,N_14189);
nand U14502 (N_14502,N_14454,N_14069);
nor U14503 (N_14503,N_14318,N_14343);
and U14504 (N_14504,N_14136,N_14224);
xnor U14505 (N_14505,N_14392,N_14449);
nor U14506 (N_14506,N_14247,N_14349);
nand U14507 (N_14507,N_14493,N_14071);
or U14508 (N_14508,N_14096,N_14179);
nor U14509 (N_14509,N_14296,N_14066);
or U14510 (N_14510,N_14172,N_14329);
nand U14511 (N_14511,N_14499,N_14466);
or U14512 (N_14512,N_14150,N_14193);
nand U14513 (N_14513,N_14480,N_14129);
or U14514 (N_14514,N_14464,N_14366);
nor U14515 (N_14515,N_14294,N_14323);
nor U14516 (N_14516,N_14341,N_14031);
nand U14517 (N_14517,N_14227,N_14041);
nand U14518 (N_14518,N_14173,N_14158);
and U14519 (N_14519,N_14133,N_14080);
or U14520 (N_14520,N_14235,N_14197);
nand U14521 (N_14521,N_14035,N_14346);
or U14522 (N_14522,N_14107,N_14125);
nand U14523 (N_14523,N_14397,N_14216);
nand U14524 (N_14524,N_14435,N_14274);
nor U14525 (N_14525,N_14325,N_14087);
nor U14526 (N_14526,N_14228,N_14255);
and U14527 (N_14527,N_14220,N_14057);
nand U14528 (N_14528,N_14091,N_14286);
nor U14529 (N_14529,N_14109,N_14036);
nor U14530 (N_14530,N_14385,N_14012);
nor U14531 (N_14531,N_14440,N_14411);
or U14532 (N_14532,N_14095,N_14160);
nand U14533 (N_14533,N_14259,N_14317);
nand U14534 (N_14534,N_14132,N_14092);
or U14535 (N_14535,N_14357,N_14446);
nand U14536 (N_14536,N_14056,N_14340);
nand U14537 (N_14537,N_14462,N_14332);
or U14538 (N_14538,N_14008,N_14492);
or U14539 (N_14539,N_14477,N_14321);
nand U14540 (N_14540,N_14037,N_14076);
nand U14541 (N_14541,N_14430,N_14350);
xor U14542 (N_14542,N_14042,N_14134);
nor U14543 (N_14543,N_14073,N_14040);
nand U14544 (N_14544,N_14112,N_14362);
nand U14545 (N_14545,N_14258,N_14077);
nand U14546 (N_14546,N_14272,N_14243);
nand U14547 (N_14547,N_14183,N_14469);
or U14548 (N_14548,N_14484,N_14100);
nor U14549 (N_14549,N_14423,N_14382);
and U14550 (N_14550,N_14265,N_14260);
and U14551 (N_14551,N_14312,N_14088);
nand U14552 (N_14552,N_14097,N_14471);
xor U14553 (N_14553,N_14305,N_14441);
nor U14554 (N_14554,N_14117,N_14068);
and U14555 (N_14555,N_14297,N_14245);
nor U14556 (N_14556,N_14447,N_14428);
nor U14557 (N_14557,N_14303,N_14249);
nor U14558 (N_14558,N_14452,N_14386);
nor U14559 (N_14559,N_14439,N_14310);
nand U14560 (N_14560,N_14413,N_14206);
nor U14561 (N_14561,N_14010,N_14024);
or U14562 (N_14562,N_14239,N_14082);
and U14563 (N_14563,N_14060,N_14052);
nand U14564 (N_14564,N_14328,N_14148);
nor U14565 (N_14565,N_14370,N_14019);
or U14566 (N_14566,N_14487,N_14049);
nand U14567 (N_14567,N_14364,N_14293);
nor U14568 (N_14568,N_14236,N_14013);
nor U14569 (N_14569,N_14048,N_14157);
nor U14570 (N_14570,N_14391,N_14098);
nand U14571 (N_14571,N_14496,N_14075);
nor U14572 (N_14572,N_14495,N_14029);
nand U14573 (N_14573,N_14166,N_14139);
xor U14574 (N_14574,N_14225,N_14395);
nand U14575 (N_14575,N_14127,N_14375);
nor U14576 (N_14576,N_14345,N_14147);
nor U14577 (N_14577,N_14211,N_14400);
or U14578 (N_14578,N_14209,N_14408);
nor U14579 (N_14579,N_14241,N_14009);
nand U14580 (N_14580,N_14256,N_14105);
or U14581 (N_14581,N_14353,N_14111);
or U14582 (N_14582,N_14420,N_14106);
and U14583 (N_14583,N_14307,N_14352);
or U14584 (N_14584,N_14055,N_14473);
or U14585 (N_14585,N_14421,N_14034);
nor U14586 (N_14586,N_14017,N_14360);
nor U14587 (N_14587,N_14119,N_14007);
and U14588 (N_14588,N_14410,N_14185);
nand U14589 (N_14589,N_14336,N_14254);
or U14590 (N_14590,N_14058,N_14394);
nand U14591 (N_14591,N_14291,N_14289);
nor U14592 (N_14592,N_14015,N_14269);
nand U14593 (N_14593,N_14151,N_14084);
and U14594 (N_14594,N_14188,N_14374);
and U14595 (N_14595,N_14416,N_14371);
nor U14596 (N_14596,N_14306,N_14481);
and U14597 (N_14597,N_14231,N_14458);
or U14598 (N_14598,N_14347,N_14018);
and U14599 (N_14599,N_14486,N_14402);
nor U14600 (N_14600,N_14497,N_14202);
nand U14601 (N_14601,N_14383,N_14445);
or U14602 (N_14602,N_14155,N_14456);
nand U14603 (N_14603,N_14381,N_14461);
nand U14604 (N_14604,N_14152,N_14417);
nor U14605 (N_14605,N_14176,N_14472);
and U14606 (N_14606,N_14368,N_14090);
nor U14607 (N_14607,N_14064,N_14443);
nand U14608 (N_14608,N_14200,N_14372);
nor U14609 (N_14609,N_14271,N_14014);
or U14610 (N_14610,N_14288,N_14468);
or U14611 (N_14611,N_14062,N_14169);
or U14612 (N_14612,N_14177,N_14161);
and U14613 (N_14613,N_14072,N_14223);
xnor U14614 (N_14614,N_14070,N_14240);
or U14615 (N_14615,N_14108,N_14438);
nand U14616 (N_14616,N_14354,N_14337);
nand U14617 (N_14617,N_14181,N_14415);
nand U14618 (N_14618,N_14118,N_14167);
xor U14619 (N_14619,N_14054,N_14032);
nor U14620 (N_14620,N_14050,N_14210);
and U14621 (N_14621,N_14011,N_14482);
nor U14622 (N_14622,N_14026,N_14268);
nand U14623 (N_14623,N_14373,N_14083);
nand U14624 (N_14624,N_14102,N_14283);
or U14625 (N_14625,N_14067,N_14038);
xor U14626 (N_14626,N_14006,N_14237);
and U14627 (N_14627,N_14455,N_14074);
xnor U14628 (N_14628,N_14021,N_14030);
nand U14629 (N_14629,N_14101,N_14367);
nor U14630 (N_14630,N_14355,N_14401);
and U14631 (N_14631,N_14207,N_14463);
nand U14632 (N_14632,N_14356,N_14184);
and U14633 (N_14633,N_14485,N_14379);
nand U14634 (N_14634,N_14406,N_14339);
nand U14635 (N_14635,N_14154,N_14190);
and U14636 (N_14636,N_14145,N_14027);
nor U14637 (N_14637,N_14278,N_14182);
xnor U14638 (N_14638,N_14214,N_14094);
xnor U14639 (N_14639,N_14232,N_14348);
or U14640 (N_14640,N_14427,N_14396);
nand U14641 (N_14641,N_14412,N_14047);
and U14642 (N_14642,N_14114,N_14033);
and U14643 (N_14643,N_14479,N_14436);
or U14644 (N_14644,N_14279,N_14489);
nor U14645 (N_14645,N_14180,N_14314);
nor U14646 (N_14646,N_14437,N_14028);
nor U14647 (N_14647,N_14065,N_14465);
nor U14648 (N_14648,N_14208,N_14344);
nand U14649 (N_14649,N_14308,N_14144);
nand U14650 (N_14650,N_14213,N_14282);
or U14651 (N_14651,N_14230,N_14322);
xnor U14652 (N_14652,N_14005,N_14351);
nor U14653 (N_14653,N_14311,N_14078);
nor U14654 (N_14654,N_14498,N_14266);
nand U14655 (N_14655,N_14262,N_14426);
nand U14656 (N_14656,N_14378,N_14363);
nor U14657 (N_14657,N_14261,N_14126);
xnor U14658 (N_14658,N_14331,N_14389);
or U14659 (N_14659,N_14298,N_14292);
xor U14660 (N_14660,N_14043,N_14153);
nor U14661 (N_14661,N_14377,N_14121);
and U14662 (N_14662,N_14104,N_14342);
or U14663 (N_14663,N_14002,N_14196);
nor U14664 (N_14664,N_14238,N_14467);
xnor U14665 (N_14665,N_14277,N_14316);
and U14666 (N_14666,N_14165,N_14120);
nor U14667 (N_14667,N_14398,N_14163);
and U14668 (N_14668,N_14276,N_14061);
nor U14669 (N_14669,N_14187,N_14085);
nor U14670 (N_14670,N_14405,N_14334);
and U14671 (N_14671,N_14434,N_14474);
nor U14672 (N_14672,N_14309,N_14201);
xor U14673 (N_14673,N_14414,N_14319);
xor U14674 (N_14674,N_14124,N_14403);
or U14675 (N_14675,N_14257,N_14001);
nand U14676 (N_14676,N_14450,N_14020);
and U14677 (N_14677,N_14330,N_14324);
xor U14678 (N_14678,N_14142,N_14444);
or U14679 (N_14679,N_14267,N_14460);
and U14680 (N_14680,N_14453,N_14099);
nor U14681 (N_14681,N_14217,N_14023);
nor U14682 (N_14682,N_14159,N_14470);
and U14683 (N_14683,N_14053,N_14300);
nor U14684 (N_14684,N_14016,N_14320);
nand U14685 (N_14685,N_14284,N_14263);
nor U14686 (N_14686,N_14476,N_14404);
and U14687 (N_14687,N_14326,N_14361);
and U14688 (N_14688,N_14252,N_14204);
nor U14689 (N_14689,N_14081,N_14250);
and U14690 (N_14690,N_14433,N_14162);
and U14691 (N_14691,N_14335,N_14365);
or U14692 (N_14692,N_14103,N_14304);
and U14693 (N_14693,N_14149,N_14483);
and U14694 (N_14694,N_14138,N_14115);
nand U14695 (N_14695,N_14222,N_14244);
and U14696 (N_14696,N_14275,N_14424);
and U14697 (N_14697,N_14143,N_14390);
nor U14698 (N_14698,N_14422,N_14141);
nor U14699 (N_14699,N_14137,N_14253);
and U14700 (N_14700,N_14295,N_14234);
nand U14701 (N_14701,N_14171,N_14419);
nand U14702 (N_14702,N_14384,N_14388);
or U14703 (N_14703,N_14429,N_14299);
nand U14704 (N_14704,N_14000,N_14191);
and U14705 (N_14705,N_14186,N_14110);
nor U14706 (N_14706,N_14387,N_14358);
and U14707 (N_14707,N_14301,N_14475);
nand U14708 (N_14708,N_14174,N_14490);
nand U14709 (N_14709,N_14369,N_14393);
or U14710 (N_14710,N_14130,N_14315);
nor U14711 (N_14711,N_14407,N_14233);
or U14712 (N_14712,N_14025,N_14451);
nor U14713 (N_14713,N_14116,N_14168);
nand U14714 (N_14714,N_14156,N_14242);
nor U14715 (N_14715,N_14199,N_14290);
nand U14716 (N_14716,N_14063,N_14113);
or U14717 (N_14717,N_14376,N_14425);
nand U14718 (N_14718,N_14146,N_14205);
and U14719 (N_14719,N_14448,N_14059);
and U14720 (N_14720,N_14089,N_14226);
and U14721 (N_14721,N_14003,N_14248);
or U14722 (N_14722,N_14022,N_14302);
nor U14723 (N_14723,N_14409,N_14442);
and U14724 (N_14724,N_14285,N_14270);
nor U14725 (N_14725,N_14218,N_14093);
or U14726 (N_14726,N_14123,N_14246);
or U14727 (N_14727,N_14164,N_14046);
nand U14728 (N_14728,N_14086,N_14215);
and U14729 (N_14729,N_14135,N_14051);
nand U14730 (N_14730,N_14194,N_14264);
nand U14731 (N_14731,N_14192,N_14431);
nor U14732 (N_14732,N_14457,N_14494);
nand U14733 (N_14733,N_14195,N_14380);
nand U14734 (N_14734,N_14039,N_14170);
nor U14735 (N_14735,N_14399,N_14432);
or U14736 (N_14736,N_14338,N_14491);
and U14737 (N_14737,N_14221,N_14203);
xnor U14738 (N_14738,N_14418,N_14251);
nand U14739 (N_14739,N_14327,N_14198);
nand U14740 (N_14740,N_14273,N_14175);
nand U14741 (N_14741,N_14131,N_14313);
nor U14742 (N_14742,N_14044,N_14333);
nor U14743 (N_14743,N_14359,N_14178);
nand U14744 (N_14744,N_14122,N_14219);
nor U14745 (N_14745,N_14212,N_14287);
or U14746 (N_14746,N_14488,N_14459);
nand U14747 (N_14747,N_14045,N_14280);
nor U14748 (N_14748,N_14128,N_14478);
nor U14749 (N_14749,N_14281,N_14079);
or U14750 (N_14750,N_14328,N_14234);
nand U14751 (N_14751,N_14025,N_14448);
and U14752 (N_14752,N_14026,N_14167);
or U14753 (N_14753,N_14466,N_14032);
nand U14754 (N_14754,N_14088,N_14452);
nand U14755 (N_14755,N_14306,N_14022);
and U14756 (N_14756,N_14039,N_14210);
nand U14757 (N_14757,N_14116,N_14414);
and U14758 (N_14758,N_14089,N_14352);
and U14759 (N_14759,N_14363,N_14016);
and U14760 (N_14760,N_14404,N_14199);
and U14761 (N_14761,N_14411,N_14450);
and U14762 (N_14762,N_14464,N_14262);
nand U14763 (N_14763,N_14092,N_14309);
or U14764 (N_14764,N_14041,N_14098);
nor U14765 (N_14765,N_14335,N_14192);
and U14766 (N_14766,N_14467,N_14385);
and U14767 (N_14767,N_14322,N_14056);
and U14768 (N_14768,N_14113,N_14389);
nand U14769 (N_14769,N_14390,N_14113);
nor U14770 (N_14770,N_14341,N_14318);
nor U14771 (N_14771,N_14050,N_14390);
nand U14772 (N_14772,N_14056,N_14488);
or U14773 (N_14773,N_14487,N_14161);
or U14774 (N_14774,N_14459,N_14165);
or U14775 (N_14775,N_14444,N_14400);
nand U14776 (N_14776,N_14282,N_14352);
nor U14777 (N_14777,N_14059,N_14230);
nor U14778 (N_14778,N_14120,N_14247);
and U14779 (N_14779,N_14463,N_14363);
nand U14780 (N_14780,N_14353,N_14462);
nor U14781 (N_14781,N_14413,N_14272);
and U14782 (N_14782,N_14009,N_14278);
nand U14783 (N_14783,N_14494,N_14304);
nand U14784 (N_14784,N_14306,N_14277);
xor U14785 (N_14785,N_14061,N_14389);
nand U14786 (N_14786,N_14285,N_14325);
and U14787 (N_14787,N_14161,N_14398);
or U14788 (N_14788,N_14474,N_14059);
nor U14789 (N_14789,N_14261,N_14487);
xor U14790 (N_14790,N_14283,N_14267);
and U14791 (N_14791,N_14201,N_14244);
xnor U14792 (N_14792,N_14457,N_14263);
nor U14793 (N_14793,N_14288,N_14004);
nand U14794 (N_14794,N_14237,N_14423);
nor U14795 (N_14795,N_14035,N_14003);
and U14796 (N_14796,N_14089,N_14080);
or U14797 (N_14797,N_14451,N_14215);
xor U14798 (N_14798,N_14117,N_14451);
and U14799 (N_14799,N_14350,N_14138);
or U14800 (N_14800,N_14429,N_14018);
or U14801 (N_14801,N_14279,N_14177);
nor U14802 (N_14802,N_14360,N_14139);
and U14803 (N_14803,N_14468,N_14414);
and U14804 (N_14804,N_14277,N_14254);
nand U14805 (N_14805,N_14485,N_14068);
or U14806 (N_14806,N_14397,N_14264);
and U14807 (N_14807,N_14370,N_14018);
and U14808 (N_14808,N_14383,N_14182);
or U14809 (N_14809,N_14317,N_14088);
xnor U14810 (N_14810,N_14132,N_14334);
nand U14811 (N_14811,N_14250,N_14319);
nor U14812 (N_14812,N_14453,N_14032);
nand U14813 (N_14813,N_14084,N_14397);
and U14814 (N_14814,N_14357,N_14444);
or U14815 (N_14815,N_14299,N_14231);
and U14816 (N_14816,N_14133,N_14333);
xnor U14817 (N_14817,N_14137,N_14153);
and U14818 (N_14818,N_14381,N_14412);
nand U14819 (N_14819,N_14031,N_14049);
and U14820 (N_14820,N_14236,N_14366);
xnor U14821 (N_14821,N_14370,N_14471);
nand U14822 (N_14822,N_14359,N_14434);
and U14823 (N_14823,N_14474,N_14177);
nor U14824 (N_14824,N_14172,N_14237);
nor U14825 (N_14825,N_14076,N_14265);
xor U14826 (N_14826,N_14480,N_14264);
nand U14827 (N_14827,N_14395,N_14319);
or U14828 (N_14828,N_14360,N_14019);
or U14829 (N_14829,N_14096,N_14435);
and U14830 (N_14830,N_14042,N_14285);
or U14831 (N_14831,N_14412,N_14468);
or U14832 (N_14832,N_14057,N_14160);
nor U14833 (N_14833,N_14036,N_14362);
nand U14834 (N_14834,N_14476,N_14346);
and U14835 (N_14835,N_14251,N_14480);
nor U14836 (N_14836,N_14124,N_14244);
or U14837 (N_14837,N_14174,N_14463);
nor U14838 (N_14838,N_14161,N_14425);
xnor U14839 (N_14839,N_14471,N_14010);
nand U14840 (N_14840,N_14380,N_14498);
nor U14841 (N_14841,N_14084,N_14018);
or U14842 (N_14842,N_14117,N_14181);
nand U14843 (N_14843,N_14383,N_14422);
and U14844 (N_14844,N_14171,N_14255);
and U14845 (N_14845,N_14142,N_14025);
nand U14846 (N_14846,N_14362,N_14428);
nor U14847 (N_14847,N_14405,N_14486);
nand U14848 (N_14848,N_14020,N_14416);
and U14849 (N_14849,N_14324,N_14150);
nand U14850 (N_14850,N_14387,N_14154);
nor U14851 (N_14851,N_14072,N_14413);
and U14852 (N_14852,N_14352,N_14130);
xnor U14853 (N_14853,N_14174,N_14370);
nor U14854 (N_14854,N_14022,N_14102);
nand U14855 (N_14855,N_14242,N_14107);
nand U14856 (N_14856,N_14181,N_14080);
nand U14857 (N_14857,N_14189,N_14170);
nor U14858 (N_14858,N_14141,N_14240);
nor U14859 (N_14859,N_14081,N_14130);
nand U14860 (N_14860,N_14241,N_14323);
nand U14861 (N_14861,N_14400,N_14419);
and U14862 (N_14862,N_14487,N_14162);
and U14863 (N_14863,N_14000,N_14204);
or U14864 (N_14864,N_14036,N_14275);
nor U14865 (N_14865,N_14459,N_14387);
or U14866 (N_14866,N_14128,N_14234);
and U14867 (N_14867,N_14095,N_14437);
xnor U14868 (N_14868,N_14083,N_14432);
and U14869 (N_14869,N_14241,N_14352);
xnor U14870 (N_14870,N_14318,N_14388);
nand U14871 (N_14871,N_14240,N_14463);
and U14872 (N_14872,N_14233,N_14149);
xnor U14873 (N_14873,N_14408,N_14059);
nand U14874 (N_14874,N_14106,N_14389);
nand U14875 (N_14875,N_14211,N_14248);
nand U14876 (N_14876,N_14374,N_14468);
nor U14877 (N_14877,N_14223,N_14346);
xnor U14878 (N_14878,N_14150,N_14034);
or U14879 (N_14879,N_14074,N_14389);
and U14880 (N_14880,N_14094,N_14480);
nand U14881 (N_14881,N_14485,N_14482);
nor U14882 (N_14882,N_14048,N_14011);
nand U14883 (N_14883,N_14347,N_14349);
xor U14884 (N_14884,N_14487,N_14094);
or U14885 (N_14885,N_14225,N_14373);
or U14886 (N_14886,N_14361,N_14227);
xnor U14887 (N_14887,N_14274,N_14250);
nand U14888 (N_14888,N_14382,N_14002);
nor U14889 (N_14889,N_14028,N_14160);
nand U14890 (N_14890,N_14193,N_14122);
or U14891 (N_14891,N_14098,N_14387);
and U14892 (N_14892,N_14470,N_14151);
nor U14893 (N_14893,N_14191,N_14114);
nor U14894 (N_14894,N_14303,N_14461);
and U14895 (N_14895,N_14284,N_14479);
and U14896 (N_14896,N_14213,N_14058);
nand U14897 (N_14897,N_14385,N_14396);
nand U14898 (N_14898,N_14327,N_14178);
xor U14899 (N_14899,N_14098,N_14094);
nor U14900 (N_14900,N_14038,N_14449);
nand U14901 (N_14901,N_14406,N_14372);
nand U14902 (N_14902,N_14090,N_14097);
nor U14903 (N_14903,N_14234,N_14453);
and U14904 (N_14904,N_14453,N_14012);
nor U14905 (N_14905,N_14229,N_14018);
xnor U14906 (N_14906,N_14176,N_14248);
nand U14907 (N_14907,N_14440,N_14170);
nand U14908 (N_14908,N_14448,N_14034);
nor U14909 (N_14909,N_14229,N_14370);
nand U14910 (N_14910,N_14382,N_14260);
nand U14911 (N_14911,N_14191,N_14083);
nor U14912 (N_14912,N_14112,N_14376);
nor U14913 (N_14913,N_14042,N_14122);
or U14914 (N_14914,N_14215,N_14261);
xnor U14915 (N_14915,N_14283,N_14133);
nor U14916 (N_14916,N_14113,N_14297);
and U14917 (N_14917,N_14262,N_14396);
or U14918 (N_14918,N_14387,N_14399);
nor U14919 (N_14919,N_14441,N_14425);
or U14920 (N_14920,N_14485,N_14124);
or U14921 (N_14921,N_14332,N_14369);
and U14922 (N_14922,N_14305,N_14121);
nor U14923 (N_14923,N_14298,N_14200);
nand U14924 (N_14924,N_14309,N_14492);
and U14925 (N_14925,N_14136,N_14326);
nor U14926 (N_14926,N_14390,N_14299);
nor U14927 (N_14927,N_14339,N_14425);
and U14928 (N_14928,N_14367,N_14075);
and U14929 (N_14929,N_14379,N_14027);
and U14930 (N_14930,N_14238,N_14396);
and U14931 (N_14931,N_14203,N_14151);
nor U14932 (N_14932,N_14436,N_14409);
and U14933 (N_14933,N_14409,N_14016);
and U14934 (N_14934,N_14447,N_14365);
or U14935 (N_14935,N_14148,N_14417);
or U14936 (N_14936,N_14012,N_14469);
or U14937 (N_14937,N_14019,N_14090);
nor U14938 (N_14938,N_14093,N_14083);
and U14939 (N_14939,N_14306,N_14312);
nand U14940 (N_14940,N_14439,N_14019);
and U14941 (N_14941,N_14083,N_14171);
and U14942 (N_14942,N_14351,N_14460);
or U14943 (N_14943,N_14182,N_14129);
or U14944 (N_14944,N_14093,N_14390);
nand U14945 (N_14945,N_14205,N_14045);
nor U14946 (N_14946,N_14410,N_14443);
nor U14947 (N_14947,N_14465,N_14025);
nor U14948 (N_14948,N_14200,N_14137);
and U14949 (N_14949,N_14112,N_14281);
xnor U14950 (N_14950,N_14085,N_14342);
or U14951 (N_14951,N_14049,N_14011);
nand U14952 (N_14952,N_14483,N_14188);
nor U14953 (N_14953,N_14331,N_14339);
xnor U14954 (N_14954,N_14207,N_14149);
and U14955 (N_14955,N_14092,N_14293);
nor U14956 (N_14956,N_14261,N_14285);
or U14957 (N_14957,N_14275,N_14209);
xor U14958 (N_14958,N_14243,N_14349);
nand U14959 (N_14959,N_14249,N_14133);
nor U14960 (N_14960,N_14154,N_14102);
nand U14961 (N_14961,N_14461,N_14252);
xnor U14962 (N_14962,N_14313,N_14470);
nor U14963 (N_14963,N_14437,N_14401);
nand U14964 (N_14964,N_14157,N_14273);
nor U14965 (N_14965,N_14149,N_14263);
or U14966 (N_14966,N_14436,N_14235);
and U14967 (N_14967,N_14458,N_14036);
and U14968 (N_14968,N_14457,N_14247);
and U14969 (N_14969,N_14438,N_14483);
xnor U14970 (N_14970,N_14351,N_14210);
xnor U14971 (N_14971,N_14003,N_14055);
nand U14972 (N_14972,N_14283,N_14461);
nand U14973 (N_14973,N_14439,N_14054);
nor U14974 (N_14974,N_14316,N_14060);
xnor U14975 (N_14975,N_14285,N_14363);
nand U14976 (N_14976,N_14269,N_14283);
nor U14977 (N_14977,N_14188,N_14088);
xor U14978 (N_14978,N_14335,N_14228);
nor U14979 (N_14979,N_14248,N_14305);
nor U14980 (N_14980,N_14233,N_14142);
and U14981 (N_14981,N_14295,N_14290);
xnor U14982 (N_14982,N_14211,N_14040);
and U14983 (N_14983,N_14350,N_14036);
xor U14984 (N_14984,N_14196,N_14013);
and U14985 (N_14985,N_14413,N_14280);
xor U14986 (N_14986,N_14170,N_14175);
nand U14987 (N_14987,N_14153,N_14470);
and U14988 (N_14988,N_14045,N_14484);
or U14989 (N_14989,N_14040,N_14309);
and U14990 (N_14990,N_14242,N_14389);
or U14991 (N_14991,N_14226,N_14103);
and U14992 (N_14992,N_14211,N_14302);
xnor U14993 (N_14993,N_14325,N_14337);
nor U14994 (N_14994,N_14367,N_14496);
nand U14995 (N_14995,N_14459,N_14480);
xnor U14996 (N_14996,N_14064,N_14097);
and U14997 (N_14997,N_14188,N_14209);
nand U14998 (N_14998,N_14042,N_14224);
xor U14999 (N_14999,N_14157,N_14165);
or U15000 (N_15000,N_14709,N_14807);
nor U15001 (N_15001,N_14936,N_14684);
nor U15002 (N_15002,N_14802,N_14842);
nand U15003 (N_15003,N_14710,N_14954);
and U15004 (N_15004,N_14873,N_14849);
nand U15005 (N_15005,N_14883,N_14526);
or U15006 (N_15006,N_14516,N_14626);
nor U15007 (N_15007,N_14756,N_14539);
and U15008 (N_15008,N_14544,N_14971);
and U15009 (N_15009,N_14831,N_14644);
nor U15010 (N_15010,N_14941,N_14905);
nor U15011 (N_15011,N_14512,N_14530);
nor U15012 (N_15012,N_14517,N_14976);
and U15013 (N_15013,N_14725,N_14909);
nand U15014 (N_15014,N_14755,N_14546);
nand U15015 (N_15015,N_14576,N_14639);
nor U15016 (N_15016,N_14803,N_14574);
or U15017 (N_15017,N_14538,N_14955);
xnor U15018 (N_15018,N_14750,N_14534);
or U15019 (N_15019,N_14880,N_14540);
xor U15020 (N_15020,N_14808,N_14996);
nand U15021 (N_15021,N_14821,N_14901);
and U15022 (N_15022,N_14765,N_14874);
nor U15023 (N_15023,N_14839,N_14716);
nor U15024 (N_15024,N_14903,N_14701);
nor U15025 (N_15025,N_14810,N_14548);
xnor U15026 (N_15026,N_14916,N_14693);
and U15027 (N_15027,N_14653,N_14929);
nand U15028 (N_15028,N_14742,N_14588);
or U15029 (N_15029,N_14781,N_14603);
or U15030 (N_15030,N_14950,N_14897);
or U15031 (N_15031,N_14993,N_14793);
xor U15032 (N_15032,N_14975,N_14577);
nand U15033 (N_15033,N_14847,N_14659);
xnor U15034 (N_15034,N_14749,N_14583);
or U15035 (N_15035,N_14715,N_14999);
nand U15036 (N_15036,N_14629,N_14942);
or U15037 (N_15037,N_14650,N_14678);
nor U15038 (N_15038,N_14616,N_14879);
or U15039 (N_15039,N_14994,N_14806);
nor U15040 (N_15040,N_14663,N_14966);
nand U15041 (N_15041,N_14763,N_14830);
or U15042 (N_15042,N_14665,N_14523);
nand U15043 (N_15043,N_14875,N_14786);
nor U15044 (N_15044,N_14995,N_14894);
nor U15045 (N_15045,N_14753,N_14984);
or U15046 (N_15046,N_14664,N_14537);
or U15047 (N_15047,N_14513,N_14835);
and U15048 (N_15048,N_14852,N_14918);
and U15049 (N_15049,N_14885,N_14989);
or U15050 (N_15050,N_14913,N_14974);
or U15051 (N_15051,N_14933,N_14967);
and U15052 (N_15052,N_14784,N_14570);
and U15053 (N_15053,N_14637,N_14815);
nand U15054 (N_15054,N_14535,N_14549);
nand U15055 (N_15055,N_14791,N_14820);
or U15056 (N_15056,N_14651,N_14553);
nor U15057 (N_15057,N_14602,N_14811);
nor U15058 (N_15058,N_14600,N_14719);
nor U15059 (N_15059,N_14944,N_14589);
nor U15060 (N_15060,N_14970,N_14630);
nor U15061 (N_15061,N_14527,N_14634);
xor U15062 (N_15062,N_14814,N_14587);
nand U15063 (N_15063,N_14851,N_14677);
nor U15064 (N_15064,N_14698,N_14843);
or U15065 (N_15065,N_14782,N_14552);
nand U15066 (N_15066,N_14785,N_14558);
or U15067 (N_15067,N_14819,N_14985);
nor U15068 (N_15068,N_14920,N_14826);
nand U15069 (N_15069,N_14979,N_14703);
or U15070 (N_15070,N_14674,N_14518);
or U15071 (N_15071,N_14987,N_14620);
or U15072 (N_15072,N_14809,N_14829);
and U15073 (N_15073,N_14688,N_14992);
xnor U15074 (N_15074,N_14866,N_14870);
nand U15075 (N_15075,N_14998,N_14708);
and U15076 (N_15076,N_14640,N_14772);
or U15077 (N_15077,N_14566,N_14717);
and U15078 (N_15078,N_14726,N_14615);
and U15079 (N_15079,N_14585,N_14804);
nand U15080 (N_15080,N_14670,N_14595);
nor U15081 (N_15081,N_14692,N_14956);
or U15082 (N_15082,N_14813,N_14667);
or U15083 (N_15083,N_14505,N_14612);
nor U15084 (N_15084,N_14965,N_14982);
xor U15085 (N_15085,N_14748,N_14925);
or U15086 (N_15086,N_14766,N_14572);
or U15087 (N_15087,N_14529,N_14652);
nor U15088 (N_15088,N_14571,N_14949);
and U15089 (N_15089,N_14641,N_14649);
and U15090 (N_15090,N_14628,N_14617);
xor U15091 (N_15091,N_14788,N_14760);
or U15092 (N_15092,N_14931,N_14777);
nor U15093 (N_15093,N_14606,N_14877);
nand U15094 (N_15094,N_14502,N_14896);
xor U15095 (N_15095,N_14927,N_14705);
nor U15096 (N_15096,N_14978,N_14579);
nor U15097 (N_15097,N_14799,N_14754);
or U15098 (N_15098,N_14739,N_14864);
xor U15099 (N_15099,N_14697,N_14919);
nand U15100 (N_15100,N_14578,N_14945);
nor U15101 (N_15101,N_14694,N_14997);
and U15102 (N_15102,N_14671,N_14594);
xor U15103 (N_15103,N_14632,N_14733);
nor U15104 (N_15104,N_14898,N_14951);
and U15105 (N_15105,N_14771,N_14604);
or U15106 (N_15106,N_14895,N_14867);
or U15107 (N_15107,N_14946,N_14661);
and U15108 (N_15108,N_14768,N_14557);
nand U15109 (N_15109,N_14747,N_14769);
nor U15110 (N_15110,N_14887,N_14536);
and U15111 (N_15111,N_14961,N_14668);
or U15112 (N_15112,N_14882,N_14625);
xnor U15113 (N_15113,N_14657,N_14565);
or U15114 (N_15114,N_14834,N_14775);
and U15115 (N_15115,N_14704,N_14861);
and U15116 (N_15116,N_14857,N_14972);
or U15117 (N_15117,N_14500,N_14921);
nor U15118 (N_15118,N_14690,N_14547);
xor U15119 (N_15119,N_14900,N_14506);
xnor U15120 (N_15120,N_14618,N_14860);
xnor U15121 (N_15121,N_14679,N_14609);
nand U15122 (N_15122,N_14714,N_14761);
or U15123 (N_15123,N_14582,N_14743);
nor U15124 (N_15124,N_14988,N_14736);
and U15125 (N_15125,N_14990,N_14531);
nor U15126 (N_15126,N_14683,N_14627);
or U15127 (N_15127,N_14605,N_14554);
and U15128 (N_15128,N_14947,N_14737);
nand U15129 (N_15129,N_14828,N_14573);
nand U15130 (N_15130,N_14818,N_14685);
nand U15131 (N_15131,N_14669,N_14621);
and U15132 (N_15132,N_14568,N_14586);
and U15133 (N_15133,N_14699,N_14796);
and U15134 (N_15134,N_14840,N_14855);
nor U15135 (N_15135,N_14859,N_14837);
and U15136 (N_15136,N_14924,N_14889);
and U15137 (N_15137,N_14752,N_14555);
nand U15138 (N_15138,N_14778,N_14613);
nand U15139 (N_15139,N_14937,N_14524);
and U15140 (N_15140,N_14886,N_14610);
or U15141 (N_15141,N_14938,N_14700);
nand U15142 (N_15142,N_14655,N_14926);
nor U15143 (N_15143,N_14686,N_14917);
or U15144 (N_15144,N_14758,N_14624);
and U15145 (N_15145,N_14598,N_14790);
nand U15146 (N_15146,N_14608,N_14767);
nor U15147 (N_15147,N_14977,N_14729);
nand U15148 (N_15148,N_14648,N_14510);
nand U15149 (N_15149,N_14824,N_14521);
nand U15150 (N_15150,N_14596,N_14783);
nor U15151 (N_15151,N_14968,N_14731);
nand U15152 (N_15152,N_14948,N_14520);
nand U15153 (N_15153,N_14904,N_14593);
and U15154 (N_15154,N_14564,N_14541);
nor U15155 (N_15155,N_14706,N_14718);
or U15156 (N_15156,N_14822,N_14935);
or U15157 (N_15157,N_14862,N_14680);
nor U15158 (N_15158,N_14922,N_14890);
nand U15159 (N_15159,N_14892,N_14939);
nor U15160 (N_15160,N_14720,N_14884);
nor U15161 (N_15161,N_14673,N_14812);
nor U15162 (N_15162,N_14681,N_14780);
nand U15163 (N_15163,N_14893,N_14881);
and U15164 (N_15164,N_14846,N_14832);
or U15165 (N_15165,N_14508,N_14740);
and U15166 (N_15166,N_14962,N_14592);
and U15167 (N_15167,N_14848,N_14580);
and U15168 (N_15168,N_14635,N_14519);
nand U15169 (N_15169,N_14643,N_14601);
xnor U15170 (N_15170,N_14854,N_14953);
xnor U15171 (N_15171,N_14713,N_14636);
nor U15172 (N_15172,N_14528,N_14741);
nand U15173 (N_15173,N_14872,N_14853);
nand U15174 (N_15174,N_14646,N_14991);
or U15175 (N_15175,N_14934,N_14823);
xnor U15176 (N_15176,N_14732,N_14730);
nor U15177 (N_15177,N_14559,N_14660);
nand U15178 (N_15178,N_14562,N_14908);
or U15179 (N_15179,N_14721,N_14759);
or U15180 (N_15180,N_14631,N_14711);
xor U15181 (N_15181,N_14675,N_14682);
nor U15182 (N_15182,N_14712,N_14622);
xor U15183 (N_15183,N_14633,N_14981);
xnor U15184 (N_15184,N_14691,N_14762);
nand U15185 (N_15185,N_14878,N_14676);
nand U15186 (N_15186,N_14638,N_14507);
or U15187 (N_15187,N_14911,N_14695);
nor U15188 (N_15188,N_14658,N_14532);
and U15189 (N_15189,N_14869,N_14983);
nor U15190 (N_15190,N_14662,N_14569);
and U15191 (N_15191,N_14827,N_14797);
nand U15192 (N_15192,N_14779,N_14910);
and U15193 (N_15193,N_14614,N_14980);
nor U15194 (N_15194,N_14522,N_14607);
and U15195 (N_15195,N_14958,N_14746);
nor U15196 (N_15196,N_14789,N_14850);
and U15197 (N_15197,N_14543,N_14656);
xnor U15198 (N_15198,N_14923,N_14932);
and U15199 (N_15199,N_14841,N_14645);
or U15200 (N_15200,N_14584,N_14551);
nor U15201 (N_15201,N_14792,N_14575);
nand U15202 (N_15202,N_14801,N_14776);
and U15203 (N_15203,N_14556,N_14542);
nand U15204 (N_15204,N_14666,N_14973);
nor U15205 (N_15205,N_14734,N_14744);
nand U15206 (N_15206,N_14914,N_14986);
nor U15207 (N_15207,N_14816,N_14647);
and U15208 (N_15208,N_14795,N_14800);
or U15209 (N_15209,N_14805,N_14928);
and U15210 (N_15210,N_14722,N_14871);
nand U15211 (N_15211,N_14906,N_14590);
or U15212 (N_15212,N_14672,N_14957);
and U15213 (N_15213,N_14623,N_14902);
xnor U15214 (N_15214,N_14764,N_14838);
nor U15215 (N_15215,N_14888,N_14591);
nor U15216 (N_15216,N_14724,N_14727);
nor U15217 (N_15217,N_14735,N_14858);
xor U15218 (N_15218,N_14868,N_14930);
xor U15219 (N_15219,N_14899,N_14833);
nor U15220 (N_15220,N_14563,N_14509);
nand U15221 (N_15221,N_14504,N_14503);
nor U15222 (N_15222,N_14787,N_14773);
nand U15223 (N_15223,N_14515,N_14774);
or U15224 (N_15224,N_14723,N_14865);
nor U15225 (N_15225,N_14738,N_14863);
or U15226 (N_15226,N_14702,N_14599);
xor U15227 (N_15227,N_14891,N_14907);
or U15228 (N_15228,N_14817,N_14952);
xor U15229 (N_15229,N_14794,N_14611);
or U15230 (N_15230,N_14561,N_14959);
nor U15231 (N_15231,N_14915,N_14689);
and U15232 (N_15232,N_14567,N_14770);
nor U15233 (N_15233,N_14696,N_14545);
nand U15234 (N_15234,N_14511,N_14745);
or U15235 (N_15235,N_14751,N_14825);
xnor U15236 (N_15236,N_14943,N_14728);
nand U15237 (N_15237,N_14525,N_14963);
or U15238 (N_15238,N_14960,N_14581);
xnor U15239 (N_15239,N_14844,N_14687);
nand U15240 (N_15240,N_14798,N_14856);
and U15241 (N_15241,N_14501,N_14560);
nor U15242 (N_15242,N_14619,N_14757);
and U15243 (N_15243,N_14964,N_14876);
nor U15244 (N_15244,N_14940,N_14597);
or U15245 (N_15245,N_14533,N_14642);
or U15246 (N_15246,N_14845,N_14836);
or U15247 (N_15247,N_14550,N_14654);
nand U15248 (N_15248,N_14912,N_14707);
nand U15249 (N_15249,N_14969,N_14514);
nor U15250 (N_15250,N_14980,N_14679);
xor U15251 (N_15251,N_14626,N_14660);
or U15252 (N_15252,N_14762,N_14579);
or U15253 (N_15253,N_14708,N_14837);
or U15254 (N_15254,N_14539,N_14929);
nand U15255 (N_15255,N_14658,N_14526);
nor U15256 (N_15256,N_14505,N_14693);
nor U15257 (N_15257,N_14906,N_14993);
xnor U15258 (N_15258,N_14874,N_14831);
and U15259 (N_15259,N_14990,N_14932);
nand U15260 (N_15260,N_14602,N_14537);
nor U15261 (N_15261,N_14620,N_14729);
and U15262 (N_15262,N_14917,N_14573);
or U15263 (N_15263,N_14772,N_14984);
nor U15264 (N_15264,N_14790,N_14764);
nor U15265 (N_15265,N_14534,N_14546);
nor U15266 (N_15266,N_14971,N_14564);
nand U15267 (N_15267,N_14758,N_14788);
nand U15268 (N_15268,N_14878,N_14983);
and U15269 (N_15269,N_14794,N_14663);
or U15270 (N_15270,N_14587,N_14566);
and U15271 (N_15271,N_14842,N_14631);
nand U15272 (N_15272,N_14826,N_14659);
nor U15273 (N_15273,N_14765,N_14808);
and U15274 (N_15274,N_14933,N_14591);
nand U15275 (N_15275,N_14915,N_14803);
and U15276 (N_15276,N_14852,N_14571);
nor U15277 (N_15277,N_14960,N_14871);
and U15278 (N_15278,N_14560,N_14547);
and U15279 (N_15279,N_14730,N_14821);
and U15280 (N_15280,N_14950,N_14694);
nand U15281 (N_15281,N_14754,N_14563);
and U15282 (N_15282,N_14865,N_14661);
or U15283 (N_15283,N_14911,N_14563);
or U15284 (N_15284,N_14565,N_14639);
nand U15285 (N_15285,N_14570,N_14659);
or U15286 (N_15286,N_14942,N_14865);
or U15287 (N_15287,N_14708,N_14535);
and U15288 (N_15288,N_14553,N_14693);
nor U15289 (N_15289,N_14738,N_14818);
nor U15290 (N_15290,N_14629,N_14864);
and U15291 (N_15291,N_14596,N_14910);
nor U15292 (N_15292,N_14848,N_14559);
nand U15293 (N_15293,N_14831,N_14903);
or U15294 (N_15294,N_14512,N_14920);
and U15295 (N_15295,N_14908,N_14891);
nor U15296 (N_15296,N_14865,N_14607);
xnor U15297 (N_15297,N_14858,N_14659);
or U15298 (N_15298,N_14807,N_14777);
nand U15299 (N_15299,N_14803,N_14788);
or U15300 (N_15300,N_14668,N_14886);
nor U15301 (N_15301,N_14577,N_14867);
nand U15302 (N_15302,N_14659,N_14818);
xor U15303 (N_15303,N_14917,N_14912);
or U15304 (N_15304,N_14649,N_14916);
xnor U15305 (N_15305,N_14536,N_14784);
or U15306 (N_15306,N_14980,N_14933);
and U15307 (N_15307,N_14681,N_14862);
xor U15308 (N_15308,N_14633,N_14510);
nor U15309 (N_15309,N_14898,N_14892);
or U15310 (N_15310,N_14590,N_14904);
nor U15311 (N_15311,N_14830,N_14962);
xor U15312 (N_15312,N_14996,N_14639);
xor U15313 (N_15313,N_14781,N_14783);
xor U15314 (N_15314,N_14693,N_14739);
nand U15315 (N_15315,N_14985,N_14970);
nand U15316 (N_15316,N_14573,N_14663);
nor U15317 (N_15317,N_14673,N_14771);
and U15318 (N_15318,N_14571,N_14837);
nor U15319 (N_15319,N_14866,N_14683);
nor U15320 (N_15320,N_14986,N_14996);
and U15321 (N_15321,N_14822,N_14732);
and U15322 (N_15322,N_14864,N_14808);
xor U15323 (N_15323,N_14546,N_14745);
nand U15324 (N_15324,N_14801,N_14846);
or U15325 (N_15325,N_14623,N_14934);
nand U15326 (N_15326,N_14847,N_14908);
or U15327 (N_15327,N_14767,N_14864);
or U15328 (N_15328,N_14784,N_14608);
nand U15329 (N_15329,N_14885,N_14695);
or U15330 (N_15330,N_14728,N_14869);
nand U15331 (N_15331,N_14504,N_14787);
nor U15332 (N_15332,N_14933,N_14527);
nand U15333 (N_15333,N_14661,N_14739);
and U15334 (N_15334,N_14855,N_14992);
nor U15335 (N_15335,N_14807,N_14577);
and U15336 (N_15336,N_14590,N_14992);
or U15337 (N_15337,N_14654,N_14755);
or U15338 (N_15338,N_14610,N_14918);
nand U15339 (N_15339,N_14637,N_14850);
and U15340 (N_15340,N_14834,N_14835);
nor U15341 (N_15341,N_14674,N_14952);
nor U15342 (N_15342,N_14927,N_14679);
nor U15343 (N_15343,N_14556,N_14897);
nor U15344 (N_15344,N_14795,N_14888);
or U15345 (N_15345,N_14632,N_14947);
nand U15346 (N_15346,N_14574,N_14757);
or U15347 (N_15347,N_14900,N_14867);
nor U15348 (N_15348,N_14617,N_14637);
nand U15349 (N_15349,N_14951,N_14562);
or U15350 (N_15350,N_14714,N_14751);
and U15351 (N_15351,N_14793,N_14910);
nand U15352 (N_15352,N_14689,N_14840);
xor U15353 (N_15353,N_14715,N_14777);
nor U15354 (N_15354,N_14637,N_14724);
nand U15355 (N_15355,N_14881,N_14590);
nor U15356 (N_15356,N_14935,N_14552);
or U15357 (N_15357,N_14922,N_14955);
or U15358 (N_15358,N_14704,N_14889);
xnor U15359 (N_15359,N_14929,N_14788);
or U15360 (N_15360,N_14855,N_14665);
nand U15361 (N_15361,N_14886,N_14767);
and U15362 (N_15362,N_14823,N_14871);
nor U15363 (N_15363,N_14855,N_14614);
or U15364 (N_15364,N_14816,N_14545);
or U15365 (N_15365,N_14502,N_14977);
nor U15366 (N_15366,N_14759,N_14653);
or U15367 (N_15367,N_14919,N_14951);
nand U15368 (N_15368,N_14733,N_14661);
nor U15369 (N_15369,N_14672,N_14500);
or U15370 (N_15370,N_14769,N_14586);
or U15371 (N_15371,N_14741,N_14973);
xnor U15372 (N_15372,N_14647,N_14704);
nor U15373 (N_15373,N_14678,N_14887);
nor U15374 (N_15374,N_14640,N_14957);
nor U15375 (N_15375,N_14522,N_14739);
nand U15376 (N_15376,N_14770,N_14879);
nor U15377 (N_15377,N_14774,N_14721);
xnor U15378 (N_15378,N_14522,N_14985);
nor U15379 (N_15379,N_14592,N_14753);
nand U15380 (N_15380,N_14794,N_14688);
nor U15381 (N_15381,N_14779,N_14625);
and U15382 (N_15382,N_14603,N_14759);
xnor U15383 (N_15383,N_14732,N_14984);
nor U15384 (N_15384,N_14508,N_14645);
and U15385 (N_15385,N_14920,N_14679);
xor U15386 (N_15386,N_14974,N_14687);
and U15387 (N_15387,N_14739,N_14882);
nor U15388 (N_15388,N_14835,N_14547);
nand U15389 (N_15389,N_14899,N_14589);
or U15390 (N_15390,N_14949,N_14576);
nor U15391 (N_15391,N_14845,N_14784);
nand U15392 (N_15392,N_14653,N_14526);
nor U15393 (N_15393,N_14615,N_14908);
xnor U15394 (N_15394,N_14524,N_14837);
nand U15395 (N_15395,N_14873,N_14708);
or U15396 (N_15396,N_14632,N_14953);
nor U15397 (N_15397,N_14800,N_14841);
and U15398 (N_15398,N_14516,N_14610);
or U15399 (N_15399,N_14679,N_14651);
nand U15400 (N_15400,N_14595,N_14905);
or U15401 (N_15401,N_14565,N_14684);
nand U15402 (N_15402,N_14997,N_14846);
nor U15403 (N_15403,N_14828,N_14654);
or U15404 (N_15404,N_14534,N_14762);
and U15405 (N_15405,N_14849,N_14705);
and U15406 (N_15406,N_14929,N_14541);
nor U15407 (N_15407,N_14665,N_14619);
nor U15408 (N_15408,N_14799,N_14715);
or U15409 (N_15409,N_14509,N_14816);
and U15410 (N_15410,N_14508,N_14572);
and U15411 (N_15411,N_14724,N_14765);
or U15412 (N_15412,N_14945,N_14682);
or U15413 (N_15413,N_14654,N_14783);
or U15414 (N_15414,N_14900,N_14698);
and U15415 (N_15415,N_14614,N_14997);
and U15416 (N_15416,N_14971,N_14947);
and U15417 (N_15417,N_14522,N_14986);
nor U15418 (N_15418,N_14987,N_14627);
nor U15419 (N_15419,N_14726,N_14952);
and U15420 (N_15420,N_14578,N_14893);
nand U15421 (N_15421,N_14898,N_14689);
and U15422 (N_15422,N_14848,N_14516);
nand U15423 (N_15423,N_14636,N_14600);
nor U15424 (N_15424,N_14852,N_14862);
and U15425 (N_15425,N_14687,N_14954);
and U15426 (N_15426,N_14908,N_14716);
xnor U15427 (N_15427,N_14511,N_14517);
nand U15428 (N_15428,N_14604,N_14846);
or U15429 (N_15429,N_14602,N_14642);
and U15430 (N_15430,N_14670,N_14652);
nor U15431 (N_15431,N_14676,N_14506);
nand U15432 (N_15432,N_14620,N_14562);
and U15433 (N_15433,N_14524,N_14662);
and U15434 (N_15434,N_14572,N_14949);
or U15435 (N_15435,N_14615,N_14628);
nand U15436 (N_15436,N_14541,N_14933);
or U15437 (N_15437,N_14511,N_14733);
nand U15438 (N_15438,N_14790,N_14736);
and U15439 (N_15439,N_14538,N_14621);
or U15440 (N_15440,N_14963,N_14704);
and U15441 (N_15441,N_14561,N_14963);
nor U15442 (N_15442,N_14516,N_14951);
xor U15443 (N_15443,N_14782,N_14746);
or U15444 (N_15444,N_14596,N_14929);
and U15445 (N_15445,N_14751,N_14589);
xor U15446 (N_15446,N_14825,N_14779);
nor U15447 (N_15447,N_14768,N_14719);
nand U15448 (N_15448,N_14725,N_14531);
or U15449 (N_15449,N_14918,N_14682);
nand U15450 (N_15450,N_14618,N_14782);
nor U15451 (N_15451,N_14500,N_14536);
nor U15452 (N_15452,N_14504,N_14719);
nand U15453 (N_15453,N_14756,N_14961);
xor U15454 (N_15454,N_14835,N_14943);
nand U15455 (N_15455,N_14633,N_14870);
or U15456 (N_15456,N_14688,N_14633);
nor U15457 (N_15457,N_14536,N_14693);
and U15458 (N_15458,N_14804,N_14701);
nand U15459 (N_15459,N_14986,N_14913);
or U15460 (N_15460,N_14934,N_14581);
nand U15461 (N_15461,N_14582,N_14758);
or U15462 (N_15462,N_14669,N_14918);
or U15463 (N_15463,N_14833,N_14738);
or U15464 (N_15464,N_14670,N_14863);
xnor U15465 (N_15465,N_14603,N_14818);
xor U15466 (N_15466,N_14663,N_14571);
or U15467 (N_15467,N_14822,N_14569);
nor U15468 (N_15468,N_14570,N_14662);
and U15469 (N_15469,N_14512,N_14564);
or U15470 (N_15470,N_14990,N_14633);
nand U15471 (N_15471,N_14633,N_14619);
and U15472 (N_15472,N_14549,N_14560);
nand U15473 (N_15473,N_14799,N_14622);
or U15474 (N_15474,N_14654,N_14728);
and U15475 (N_15475,N_14879,N_14564);
xor U15476 (N_15476,N_14668,N_14816);
nor U15477 (N_15477,N_14975,N_14898);
or U15478 (N_15478,N_14961,N_14595);
or U15479 (N_15479,N_14845,N_14571);
nor U15480 (N_15480,N_14690,N_14884);
or U15481 (N_15481,N_14733,N_14639);
and U15482 (N_15482,N_14693,N_14948);
nand U15483 (N_15483,N_14921,N_14911);
xnor U15484 (N_15484,N_14710,N_14526);
xor U15485 (N_15485,N_14898,N_14927);
nand U15486 (N_15486,N_14904,N_14504);
xnor U15487 (N_15487,N_14941,N_14922);
and U15488 (N_15488,N_14986,N_14877);
nand U15489 (N_15489,N_14837,N_14990);
nor U15490 (N_15490,N_14940,N_14611);
and U15491 (N_15491,N_14549,N_14804);
and U15492 (N_15492,N_14694,N_14568);
nor U15493 (N_15493,N_14939,N_14864);
and U15494 (N_15494,N_14635,N_14910);
xnor U15495 (N_15495,N_14901,N_14717);
or U15496 (N_15496,N_14757,N_14914);
nand U15497 (N_15497,N_14604,N_14991);
and U15498 (N_15498,N_14527,N_14848);
nor U15499 (N_15499,N_14500,N_14519);
nor U15500 (N_15500,N_15322,N_15461);
and U15501 (N_15501,N_15009,N_15042);
nor U15502 (N_15502,N_15310,N_15220);
nor U15503 (N_15503,N_15185,N_15339);
and U15504 (N_15504,N_15386,N_15488);
nor U15505 (N_15505,N_15482,N_15391);
or U15506 (N_15506,N_15279,N_15382);
or U15507 (N_15507,N_15441,N_15135);
or U15508 (N_15508,N_15173,N_15206);
and U15509 (N_15509,N_15238,N_15025);
nor U15510 (N_15510,N_15224,N_15203);
xor U15511 (N_15511,N_15127,N_15290);
nor U15512 (N_15512,N_15214,N_15332);
and U15513 (N_15513,N_15340,N_15007);
or U15514 (N_15514,N_15186,N_15342);
nand U15515 (N_15515,N_15284,N_15478);
nor U15516 (N_15516,N_15176,N_15160);
and U15517 (N_15517,N_15018,N_15414);
nand U15518 (N_15518,N_15493,N_15169);
nor U15519 (N_15519,N_15205,N_15247);
nand U15520 (N_15520,N_15435,N_15336);
nor U15521 (N_15521,N_15243,N_15014);
nor U15522 (N_15522,N_15302,N_15081);
and U15523 (N_15523,N_15005,N_15193);
xor U15524 (N_15524,N_15099,N_15418);
nand U15525 (N_15525,N_15385,N_15432);
and U15526 (N_15526,N_15459,N_15352);
nand U15527 (N_15527,N_15106,N_15469);
or U15528 (N_15528,N_15394,N_15375);
or U15529 (N_15529,N_15032,N_15334);
and U15530 (N_15530,N_15345,N_15240);
nand U15531 (N_15531,N_15314,N_15098);
and U15532 (N_15532,N_15162,N_15323);
nor U15533 (N_15533,N_15113,N_15150);
or U15534 (N_15534,N_15016,N_15415);
or U15535 (N_15535,N_15120,N_15215);
or U15536 (N_15536,N_15367,N_15008);
nor U15537 (N_15537,N_15174,N_15430);
or U15538 (N_15538,N_15064,N_15245);
nand U15539 (N_15539,N_15115,N_15295);
or U15540 (N_15540,N_15209,N_15420);
nand U15541 (N_15541,N_15273,N_15464);
nor U15542 (N_15542,N_15318,N_15251);
and U15543 (N_15543,N_15211,N_15147);
and U15544 (N_15544,N_15440,N_15368);
nand U15545 (N_15545,N_15297,N_15024);
or U15546 (N_15546,N_15242,N_15082);
or U15547 (N_15547,N_15110,N_15033);
or U15548 (N_15548,N_15476,N_15254);
nor U15549 (N_15549,N_15274,N_15192);
or U15550 (N_15550,N_15156,N_15483);
or U15551 (N_15551,N_15378,N_15079);
nor U15552 (N_15552,N_15264,N_15012);
xor U15553 (N_15553,N_15196,N_15383);
and U15554 (N_15554,N_15261,N_15445);
or U15555 (N_15555,N_15299,N_15117);
nand U15556 (N_15556,N_15002,N_15104);
nor U15557 (N_15557,N_15419,N_15125);
and U15558 (N_15558,N_15460,N_15021);
nor U15559 (N_15559,N_15294,N_15085);
or U15560 (N_15560,N_15409,N_15423);
or U15561 (N_15561,N_15275,N_15103);
nor U15562 (N_15562,N_15475,N_15286);
or U15563 (N_15563,N_15281,N_15132);
nand U15564 (N_15564,N_15401,N_15210);
and U15565 (N_15565,N_15232,N_15112);
nand U15566 (N_15566,N_15278,N_15397);
or U15567 (N_15567,N_15496,N_15041);
or U15568 (N_15568,N_15031,N_15320);
and U15569 (N_15569,N_15481,N_15234);
nand U15570 (N_15570,N_15265,N_15096);
or U15571 (N_15571,N_15017,N_15027);
nor U15572 (N_15572,N_15470,N_15260);
or U15573 (N_15573,N_15425,N_15355);
nor U15574 (N_15574,N_15022,N_15305);
or U15575 (N_15575,N_15485,N_15035);
xor U15576 (N_15576,N_15263,N_15202);
nor U15577 (N_15577,N_15097,N_15237);
or U15578 (N_15578,N_15114,N_15328);
and U15579 (N_15579,N_15093,N_15387);
or U15580 (N_15580,N_15226,N_15457);
or U15581 (N_15581,N_15412,N_15066);
or U15582 (N_15582,N_15129,N_15253);
or U15583 (N_15583,N_15123,N_15316);
and U15584 (N_15584,N_15163,N_15487);
xor U15585 (N_15585,N_15402,N_15139);
nand U15586 (N_15586,N_15410,N_15088);
or U15587 (N_15587,N_15450,N_15443);
nor U15588 (N_15588,N_15241,N_15142);
nand U15589 (N_15589,N_15447,N_15134);
xor U15590 (N_15590,N_15231,N_15276);
and U15591 (N_15591,N_15213,N_15061);
or U15592 (N_15592,N_15236,N_15317);
nor U15593 (N_15593,N_15092,N_15019);
xor U15594 (N_15594,N_15000,N_15140);
nor U15595 (N_15595,N_15189,N_15034);
nand U15596 (N_15596,N_15072,N_15172);
nand U15597 (N_15597,N_15298,N_15122);
or U15598 (N_15598,N_15063,N_15369);
nand U15599 (N_15599,N_15379,N_15486);
nor U15600 (N_15600,N_15148,N_15494);
and U15601 (N_15601,N_15056,N_15288);
nor U15602 (N_15602,N_15146,N_15168);
and U15603 (N_15603,N_15145,N_15116);
or U15604 (N_15604,N_15083,N_15325);
or U15605 (N_15605,N_15393,N_15131);
and U15606 (N_15606,N_15304,N_15078);
and U15607 (N_15607,N_15407,N_15060);
nor U15608 (N_15608,N_15144,N_15257);
nor U15609 (N_15609,N_15400,N_15178);
nor U15610 (N_15610,N_15405,N_15490);
nand U15611 (N_15611,N_15433,N_15427);
nand U15612 (N_15612,N_15121,N_15474);
or U15613 (N_15613,N_15084,N_15171);
xnor U15614 (N_15614,N_15353,N_15453);
nand U15615 (N_15615,N_15479,N_15499);
and U15616 (N_15616,N_15216,N_15349);
nand U15617 (N_15617,N_15293,N_15262);
nor U15618 (N_15618,N_15439,N_15181);
nand U15619 (N_15619,N_15180,N_15444);
and U15620 (N_15620,N_15200,N_15244);
or U15621 (N_15621,N_15381,N_15292);
nand U15622 (N_15622,N_15363,N_15086);
or U15623 (N_15623,N_15046,N_15313);
and U15624 (N_15624,N_15187,N_15119);
nor U15625 (N_15625,N_15319,N_15102);
or U15626 (N_15626,N_15158,N_15337);
xor U15627 (N_15627,N_15100,N_15309);
or U15628 (N_15628,N_15473,N_15184);
nor U15629 (N_15629,N_15437,N_15164);
nor U15630 (N_15630,N_15347,N_15311);
nand U15631 (N_15631,N_15073,N_15133);
and U15632 (N_15632,N_15175,N_15235);
nor U15633 (N_15633,N_15404,N_15068);
nor U15634 (N_15634,N_15182,N_15333);
nand U15635 (N_15635,N_15417,N_15455);
or U15636 (N_15636,N_15268,N_15364);
nor U15637 (N_15637,N_15348,N_15159);
or U15638 (N_15638,N_15495,N_15076);
nor U15639 (N_15639,N_15312,N_15011);
nor U15640 (N_15640,N_15390,N_15054);
xor U15641 (N_15641,N_15207,N_15472);
or U15642 (N_15642,N_15366,N_15300);
and U15643 (N_15643,N_15108,N_15201);
and U15644 (N_15644,N_15036,N_15259);
and U15645 (N_15645,N_15413,N_15198);
and U15646 (N_15646,N_15357,N_15388);
or U15647 (N_15647,N_15395,N_15406);
nand U15648 (N_15648,N_15468,N_15408);
nor U15649 (N_15649,N_15343,N_15266);
nor U15650 (N_15650,N_15255,N_15030);
nand U15651 (N_15651,N_15167,N_15227);
nand U15652 (N_15652,N_15095,N_15285);
and U15653 (N_15653,N_15372,N_15059);
and U15654 (N_15654,N_15087,N_15258);
nand U15655 (N_15655,N_15448,N_15296);
nor U15656 (N_15656,N_15471,N_15043);
xor U15657 (N_15657,N_15212,N_15277);
or U15658 (N_15658,N_15351,N_15438);
or U15659 (N_15659,N_15049,N_15015);
and U15660 (N_15660,N_15228,N_15452);
and U15661 (N_15661,N_15126,N_15111);
or U15662 (N_15662,N_15052,N_15089);
and U15663 (N_15663,N_15177,N_15331);
nand U15664 (N_15664,N_15329,N_15197);
or U15665 (N_15665,N_15341,N_15436);
or U15666 (N_15666,N_15023,N_15006);
and U15667 (N_15667,N_15359,N_15491);
or U15668 (N_15668,N_15053,N_15327);
and U15669 (N_15669,N_15190,N_15039);
nand U15670 (N_15670,N_15465,N_15107);
or U15671 (N_15671,N_15149,N_15128);
nand U15672 (N_15672,N_15045,N_15396);
nor U15673 (N_15673,N_15303,N_15280);
and U15674 (N_15674,N_15252,N_15020);
nor U15675 (N_15675,N_15071,N_15040);
or U15676 (N_15676,N_15358,N_15239);
and U15677 (N_15677,N_15467,N_15058);
xnor U15678 (N_15678,N_15466,N_15246);
nor U15679 (N_15679,N_15048,N_15118);
or U15680 (N_15680,N_15399,N_15248);
nor U15681 (N_15681,N_15271,N_15335);
nor U15682 (N_15682,N_15194,N_15074);
nand U15683 (N_15683,N_15219,N_15130);
xor U15684 (N_15684,N_15289,N_15165);
and U15685 (N_15685,N_15250,N_15094);
xor U15686 (N_15686,N_15230,N_15057);
nand U15687 (N_15687,N_15301,N_15380);
or U15688 (N_15688,N_15428,N_15223);
and U15689 (N_15689,N_15191,N_15003);
nand U15690 (N_15690,N_15055,N_15101);
or U15691 (N_15691,N_15195,N_15037);
and U15692 (N_15692,N_15324,N_15492);
nor U15693 (N_15693,N_15456,N_15384);
or U15694 (N_15694,N_15065,N_15075);
nor U15695 (N_15695,N_15429,N_15070);
and U15696 (N_15696,N_15137,N_15221);
or U15697 (N_15697,N_15321,N_15365);
and U15698 (N_15698,N_15421,N_15308);
or U15699 (N_15699,N_15291,N_15426);
nor U15700 (N_15700,N_15013,N_15267);
or U15701 (N_15701,N_15346,N_15287);
or U15702 (N_15702,N_15424,N_15344);
nand U15703 (N_15703,N_15141,N_15218);
and U15704 (N_15704,N_15480,N_15138);
nand U15705 (N_15705,N_15477,N_15051);
and U15706 (N_15706,N_15179,N_15204);
or U15707 (N_15707,N_15155,N_15062);
and U15708 (N_15708,N_15451,N_15028);
or U15709 (N_15709,N_15411,N_15449);
or U15710 (N_15710,N_15222,N_15090);
or U15711 (N_15711,N_15249,N_15356);
or U15712 (N_15712,N_15484,N_15124);
nand U15713 (N_15713,N_15029,N_15403);
nor U15714 (N_15714,N_15136,N_15462);
nor U15715 (N_15715,N_15069,N_15446);
or U15716 (N_15716,N_15001,N_15498);
nand U15717 (N_15717,N_15272,N_15422);
nor U15718 (N_15718,N_15360,N_15256);
and U15719 (N_15719,N_15389,N_15038);
nor U15720 (N_15720,N_15166,N_15199);
nor U15721 (N_15721,N_15004,N_15229);
and U15722 (N_15722,N_15463,N_15361);
and U15723 (N_15723,N_15354,N_15315);
or U15724 (N_15724,N_15362,N_15307);
xnor U15725 (N_15725,N_15183,N_15010);
nor U15726 (N_15726,N_15282,N_15371);
and U15727 (N_15727,N_15374,N_15283);
or U15728 (N_15728,N_15170,N_15269);
nand U15729 (N_15729,N_15152,N_15326);
nor U15730 (N_15730,N_15044,N_15161);
and U15731 (N_15731,N_15208,N_15050);
nor U15732 (N_15732,N_15233,N_15306);
and U15733 (N_15733,N_15047,N_15143);
nor U15734 (N_15734,N_15338,N_15077);
or U15735 (N_15735,N_15091,N_15416);
nor U15736 (N_15736,N_15151,N_15442);
or U15737 (N_15737,N_15080,N_15392);
nand U15738 (N_15738,N_15225,N_15377);
or U15739 (N_15739,N_15105,N_15026);
and U15740 (N_15740,N_15434,N_15067);
or U15741 (N_15741,N_15497,N_15350);
or U15742 (N_15742,N_15217,N_15370);
xnor U15743 (N_15743,N_15157,N_15373);
nand U15744 (N_15744,N_15188,N_15153);
or U15745 (N_15745,N_15454,N_15109);
and U15746 (N_15746,N_15154,N_15376);
nor U15747 (N_15747,N_15330,N_15458);
nand U15748 (N_15748,N_15431,N_15270);
or U15749 (N_15749,N_15398,N_15489);
xnor U15750 (N_15750,N_15465,N_15168);
xor U15751 (N_15751,N_15224,N_15118);
and U15752 (N_15752,N_15058,N_15149);
and U15753 (N_15753,N_15481,N_15457);
and U15754 (N_15754,N_15301,N_15402);
and U15755 (N_15755,N_15456,N_15057);
and U15756 (N_15756,N_15200,N_15000);
nor U15757 (N_15757,N_15437,N_15249);
and U15758 (N_15758,N_15283,N_15345);
nand U15759 (N_15759,N_15309,N_15450);
or U15760 (N_15760,N_15207,N_15125);
nand U15761 (N_15761,N_15112,N_15225);
xor U15762 (N_15762,N_15121,N_15302);
or U15763 (N_15763,N_15404,N_15055);
nor U15764 (N_15764,N_15002,N_15033);
xnor U15765 (N_15765,N_15262,N_15069);
and U15766 (N_15766,N_15219,N_15076);
nand U15767 (N_15767,N_15306,N_15341);
and U15768 (N_15768,N_15248,N_15485);
xnor U15769 (N_15769,N_15074,N_15126);
nand U15770 (N_15770,N_15164,N_15270);
and U15771 (N_15771,N_15267,N_15271);
nand U15772 (N_15772,N_15229,N_15205);
nor U15773 (N_15773,N_15249,N_15483);
or U15774 (N_15774,N_15214,N_15468);
or U15775 (N_15775,N_15346,N_15245);
and U15776 (N_15776,N_15361,N_15062);
nor U15777 (N_15777,N_15386,N_15450);
or U15778 (N_15778,N_15018,N_15361);
and U15779 (N_15779,N_15221,N_15413);
nor U15780 (N_15780,N_15153,N_15029);
xnor U15781 (N_15781,N_15214,N_15261);
or U15782 (N_15782,N_15170,N_15303);
and U15783 (N_15783,N_15327,N_15005);
or U15784 (N_15784,N_15040,N_15449);
and U15785 (N_15785,N_15065,N_15132);
nor U15786 (N_15786,N_15323,N_15196);
and U15787 (N_15787,N_15157,N_15037);
and U15788 (N_15788,N_15212,N_15388);
xnor U15789 (N_15789,N_15146,N_15119);
nand U15790 (N_15790,N_15386,N_15373);
or U15791 (N_15791,N_15373,N_15351);
nand U15792 (N_15792,N_15172,N_15348);
nand U15793 (N_15793,N_15153,N_15241);
xor U15794 (N_15794,N_15092,N_15142);
nor U15795 (N_15795,N_15373,N_15394);
xnor U15796 (N_15796,N_15064,N_15417);
nand U15797 (N_15797,N_15081,N_15101);
xor U15798 (N_15798,N_15220,N_15438);
or U15799 (N_15799,N_15411,N_15210);
nand U15800 (N_15800,N_15022,N_15255);
nand U15801 (N_15801,N_15238,N_15090);
nor U15802 (N_15802,N_15108,N_15377);
nor U15803 (N_15803,N_15486,N_15193);
nand U15804 (N_15804,N_15122,N_15417);
and U15805 (N_15805,N_15324,N_15084);
nand U15806 (N_15806,N_15023,N_15027);
nor U15807 (N_15807,N_15107,N_15283);
nand U15808 (N_15808,N_15410,N_15091);
xnor U15809 (N_15809,N_15286,N_15109);
or U15810 (N_15810,N_15022,N_15021);
nand U15811 (N_15811,N_15380,N_15006);
or U15812 (N_15812,N_15479,N_15204);
and U15813 (N_15813,N_15078,N_15212);
and U15814 (N_15814,N_15129,N_15073);
xor U15815 (N_15815,N_15180,N_15405);
or U15816 (N_15816,N_15248,N_15064);
nand U15817 (N_15817,N_15179,N_15252);
or U15818 (N_15818,N_15428,N_15347);
or U15819 (N_15819,N_15323,N_15329);
nor U15820 (N_15820,N_15075,N_15433);
nand U15821 (N_15821,N_15123,N_15314);
and U15822 (N_15822,N_15283,N_15258);
and U15823 (N_15823,N_15474,N_15381);
xnor U15824 (N_15824,N_15255,N_15050);
and U15825 (N_15825,N_15296,N_15031);
or U15826 (N_15826,N_15468,N_15389);
nand U15827 (N_15827,N_15315,N_15383);
and U15828 (N_15828,N_15244,N_15164);
and U15829 (N_15829,N_15198,N_15437);
nand U15830 (N_15830,N_15432,N_15439);
nor U15831 (N_15831,N_15026,N_15431);
nor U15832 (N_15832,N_15143,N_15263);
and U15833 (N_15833,N_15436,N_15217);
and U15834 (N_15834,N_15099,N_15073);
or U15835 (N_15835,N_15097,N_15431);
or U15836 (N_15836,N_15159,N_15381);
or U15837 (N_15837,N_15183,N_15144);
nor U15838 (N_15838,N_15242,N_15321);
or U15839 (N_15839,N_15087,N_15014);
xor U15840 (N_15840,N_15329,N_15136);
or U15841 (N_15841,N_15024,N_15218);
and U15842 (N_15842,N_15417,N_15121);
or U15843 (N_15843,N_15402,N_15094);
nor U15844 (N_15844,N_15016,N_15434);
or U15845 (N_15845,N_15086,N_15183);
and U15846 (N_15846,N_15475,N_15441);
nor U15847 (N_15847,N_15452,N_15188);
nor U15848 (N_15848,N_15045,N_15069);
nor U15849 (N_15849,N_15383,N_15292);
nor U15850 (N_15850,N_15287,N_15102);
or U15851 (N_15851,N_15309,N_15102);
nand U15852 (N_15852,N_15324,N_15147);
and U15853 (N_15853,N_15460,N_15097);
nand U15854 (N_15854,N_15004,N_15198);
nor U15855 (N_15855,N_15396,N_15439);
or U15856 (N_15856,N_15047,N_15151);
nor U15857 (N_15857,N_15157,N_15366);
xnor U15858 (N_15858,N_15179,N_15362);
nor U15859 (N_15859,N_15155,N_15070);
xor U15860 (N_15860,N_15020,N_15094);
nor U15861 (N_15861,N_15450,N_15422);
nor U15862 (N_15862,N_15171,N_15159);
nand U15863 (N_15863,N_15250,N_15200);
and U15864 (N_15864,N_15415,N_15370);
nor U15865 (N_15865,N_15173,N_15002);
nor U15866 (N_15866,N_15426,N_15395);
and U15867 (N_15867,N_15128,N_15495);
nand U15868 (N_15868,N_15206,N_15430);
nand U15869 (N_15869,N_15348,N_15408);
and U15870 (N_15870,N_15477,N_15458);
and U15871 (N_15871,N_15078,N_15342);
nor U15872 (N_15872,N_15340,N_15283);
nor U15873 (N_15873,N_15142,N_15030);
and U15874 (N_15874,N_15314,N_15011);
and U15875 (N_15875,N_15199,N_15327);
nand U15876 (N_15876,N_15084,N_15169);
nor U15877 (N_15877,N_15290,N_15499);
and U15878 (N_15878,N_15473,N_15064);
nor U15879 (N_15879,N_15027,N_15308);
nor U15880 (N_15880,N_15438,N_15122);
nor U15881 (N_15881,N_15003,N_15065);
xnor U15882 (N_15882,N_15083,N_15223);
or U15883 (N_15883,N_15383,N_15102);
and U15884 (N_15884,N_15295,N_15476);
and U15885 (N_15885,N_15184,N_15369);
and U15886 (N_15886,N_15337,N_15332);
or U15887 (N_15887,N_15309,N_15320);
nand U15888 (N_15888,N_15242,N_15149);
or U15889 (N_15889,N_15393,N_15218);
or U15890 (N_15890,N_15110,N_15208);
nor U15891 (N_15891,N_15169,N_15285);
nand U15892 (N_15892,N_15256,N_15222);
and U15893 (N_15893,N_15021,N_15493);
and U15894 (N_15894,N_15040,N_15429);
or U15895 (N_15895,N_15411,N_15289);
nor U15896 (N_15896,N_15304,N_15172);
or U15897 (N_15897,N_15140,N_15219);
and U15898 (N_15898,N_15259,N_15212);
nand U15899 (N_15899,N_15010,N_15384);
nand U15900 (N_15900,N_15082,N_15399);
or U15901 (N_15901,N_15143,N_15430);
nor U15902 (N_15902,N_15419,N_15488);
xnor U15903 (N_15903,N_15006,N_15037);
or U15904 (N_15904,N_15189,N_15434);
nor U15905 (N_15905,N_15231,N_15122);
nand U15906 (N_15906,N_15072,N_15343);
or U15907 (N_15907,N_15490,N_15301);
nor U15908 (N_15908,N_15276,N_15202);
xnor U15909 (N_15909,N_15326,N_15489);
and U15910 (N_15910,N_15434,N_15301);
and U15911 (N_15911,N_15332,N_15341);
or U15912 (N_15912,N_15303,N_15068);
nand U15913 (N_15913,N_15008,N_15168);
or U15914 (N_15914,N_15458,N_15074);
xnor U15915 (N_15915,N_15335,N_15414);
or U15916 (N_15916,N_15402,N_15193);
or U15917 (N_15917,N_15344,N_15026);
nor U15918 (N_15918,N_15321,N_15233);
nor U15919 (N_15919,N_15087,N_15312);
or U15920 (N_15920,N_15095,N_15308);
nor U15921 (N_15921,N_15229,N_15426);
nand U15922 (N_15922,N_15381,N_15123);
xor U15923 (N_15923,N_15386,N_15401);
nor U15924 (N_15924,N_15380,N_15113);
and U15925 (N_15925,N_15081,N_15221);
xor U15926 (N_15926,N_15082,N_15318);
or U15927 (N_15927,N_15437,N_15351);
nor U15928 (N_15928,N_15271,N_15077);
nor U15929 (N_15929,N_15075,N_15012);
nand U15930 (N_15930,N_15484,N_15299);
nor U15931 (N_15931,N_15494,N_15379);
and U15932 (N_15932,N_15002,N_15469);
and U15933 (N_15933,N_15137,N_15444);
and U15934 (N_15934,N_15011,N_15125);
nand U15935 (N_15935,N_15145,N_15067);
or U15936 (N_15936,N_15088,N_15136);
nor U15937 (N_15937,N_15494,N_15370);
or U15938 (N_15938,N_15096,N_15451);
and U15939 (N_15939,N_15120,N_15145);
nand U15940 (N_15940,N_15109,N_15063);
nand U15941 (N_15941,N_15017,N_15471);
nor U15942 (N_15942,N_15403,N_15239);
nand U15943 (N_15943,N_15120,N_15406);
xnor U15944 (N_15944,N_15279,N_15324);
or U15945 (N_15945,N_15359,N_15047);
or U15946 (N_15946,N_15027,N_15388);
nand U15947 (N_15947,N_15477,N_15267);
xnor U15948 (N_15948,N_15001,N_15206);
and U15949 (N_15949,N_15325,N_15128);
nand U15950 (N_15950,N_15401,N_15374);
and U15951 (N_15951,N_15243,N_15030);
nor U15952 (N_15952,N_15423,N_15217);
nand U15953 (N_15953,N_15266,N_15469);
and U15954 (N_15954,N_15340,N_15304);
and U15955 (N_15955,N_15175,N_15009);
nand U15956 (N_15956,N_15098,N_15374);
nor U15957 (N_15957,N_15357,N_15186);
or U15958 (N_15958,N_15442,N_15088);
or U15959 (N_15959,N_15048,N_15039);
or U15960 (N_15960,N_15486,N_15257);
nor U15961 (N_15961,N_15088,N_15048);
and U15962 (N_15962,N_15182,N_15216);
and U15963 (N_15963,N_15218,N_15023);
nand U15964 (N_15964,N_15063,N_15320);
nor U15965 (N_15965,N_15100,N_15336);
nand U15966 (N_15966,N_15452,N_15374);
nand U15967 (N_15967,N_15455,N_15406);
and U15968 (N_15968,N_15349,N_15243);
and U15969 (N_15969,N_15472,N_15160);
or U15970 (N_15970,N_15206,N_15340);
and U15971 (N_15971,N_15494,N_15159);
and U15972 (N_15972,N_15252,N_15084);
or U15973 (N_15973,N_15052,N_15062);
or U15974 (N_15974,N_15097,N_15023);
or U15975 (N_15975,N_15000,N_15085);
and U15976 (N_15976,N_15443,N_15185);
and U15977 (N_15977,N_15272,N_15346);
nand U15978 (N_15978,N_15226,N_15442);
xor U15979 (N_15979,N_15101,N_15162);
and U15980 (N_15980,N_15054,N_15186);
or U15981 (N_15981,N_15448,N_15415);
and U15982 (N_15982,N_15362,N_15133);
or U15983 (N_15983,N_15379,N_15384);
xnor U15984 (N_15984,N_15196,N_15303);
xor U15985 (N_15985,N_15314,N_15231);
and U15986 (N_15986,N_15086,N_15356);
and U15987 (N_15987,N_15183,N_15039);
nor U15988 (N_15988,N_15398,N_15112);
nand U15989 (N_15989,N_15065,N_15396);
and U15990 (N_15990,N_15080,N_15177);
or U15991 (N_15991,N_15067,N_15499);
nor U15992 (N_15992,N_15443,N_15026);
nand U15993 (N_15993,N_15360,N_15339);
or U15994 (N_15994,N_15236,N_15011);
or U15995 (N_15995,N_15226,N_15256);
nor U15996 (N_15996,N_15463,N_15115);
or U15997 (N_15997,N_15050,N_15298);
xor U15998 (N_15998,N_15185,N_15043);
or U15999 (N_15999,N_15397,N_15497);
or U16000 (N_16000,N_15697,N_15720);
and U16001 (N_16001,N_15640,N_15791);
and U16002 (N_16002,N_15989,N_15570);
and U16003 (N_16003,N_15765,N_15584);
nand U16004 (N_16004,N_15810,N_15968);
and U16005 (N_16005,N_15838,N_15926);
nand U16006 (N_16006,N_15759,N_15598);
and U16007 (N_16007,N_15876,N_15757);
or U16008 (N_16008,N_15731,N_15800);
or U16009 (N_16009,N_15885,N_15874);
xnor U16010 (N_16010,N_15955,N_15820);
nor U16011 (N_16011,N_15949,N_15884);
and U16012 (N_16012,N_15725,N_15933);
or U16013 (N_16013,N_15695,N_15612);
nor U16014 (N_16014,N_15806,N_15663);
or U16015 (N_16015,N_15661,N_15898);
nand U16016 (N_16016,N_15622,N_15694);
and U16017 (N_16017,N_15659,N_15973);
nor U16018 (N_16018,N_15650,N_15672);
nand U16019 (N_16019,N_15771,N_15678);
xor U16020 (N_16020,N_15586,N_15675);
and U16021 (N_16021,N_15630,N_15578);
or U16022 (N_16022,N_15875,N_15600);
or U16023 (N_16023,N_15547,N_15819);
nand U16024 (N_16024,N_15631,N_15729);
and U16025 (N_16025,N_15770,N_15544);
or U16026 (N_16026,N_15746,N_15660);
or U16027 (N_16027,N_15868,N_15902);
xnor U16028 (N_16028,N_15957,N_15548);
nor U16029 (N_16029,N_15644,N_15888);
nand U16030 (N_16030,N_15946,N_15512);
nor U16031 (N_16031,N_15684,N_15528);
and U16032 (N_16032,N_15818,N_15680);
nand U16033 (N_16033,N_15763,N_15747);
and U16034 (N_16034,N_15950,N_15550);
and U16035 (N_16035,N_15718,N_15906);
or U16036 (N_16036,N_15863,N_15614);
nand U16037 (N_16037,N_15561,N_15596);
nor U16038 (N_16038,N_15951,N_15877);
nand U16039 (N_16039,N_15904,N_15538);
nor U16040 (N_16040,N_15750,N_15710);
or U16041 (N_16041,N_15626,N_15722);
nand U16042 (N_16042,N_15577,N_15628);
nor U16043 (N_16043,N_15505,N_15674);
and U16044 (N_16044,N_15590,N_15603);
nor U16045 (N_16045,N_15593,N_15517);
nand U16046 (N_16046,N_15783,N_15691);
and U16047 (N_16047,N_15769,N_15959);
nor U16048 (N_16048,N_15567,N_15982);
nand U16049 (N_16049,N_15647,N_15639);
nand U16050 (N_16050,N_15671,N_15627);
and U16051 (N_16051,N_15866,N_15589);
nand U16052 (N_16052,N_15900,N_15733);
nand U16053 (N_16053,N_15635,N_15536);
nor U16054 (N_16054,N_15696,N_15778);
and U16055 (N_16055,N_15713,N_15616);
or U16056 (N_16056,N_15918,N_15814);
or U16057 (N_16057,N_15840,N_15782);
and U16058 (N_16058,N_15935,N_15604);
nor U16059 (N_16059,N_15607,N_15541);
nand U16060 (N_16060,N_15502,N_15751);
nor U16061 (N_16061,N_15523,N_15862);
or U16062 (N_16062,N_15673,N_15821);
xnor U16063 (N_16063,N_15668,N_15998);
or U16064 (N_16064,N_15855,N_15905);
nand U16065 (N_16065,N_15909,N_15851);
nor U16066 (N_16066,N_15755,N_15756);
nand U16067 (N_16067,N_15859,N_15934);
and U16068 (N_16068,N_15901,N_15585);
nor U16069 (N_16069,N_15915,N_15619);
xnor U16070 (N_16070,N_15845,N_15999);
and U16071 (N_16071,N_15768,N_15583);
nor U16072 (N_16072,N_15519,N_15752);
nand U16073 (N_16073,N_15568,N_15521);
xnor U16074 (N_16074,N_15858,N_15636);
and U16075 (N_16075,N_15942,N_15686);
nand U16076 (N_16076,N_15848,N_15913);
or U16077 (N_16077,N_15709,N_15816);
nand U16078 (N_16078,N_15534,N_15588);
and U16079 (N_16079,N_15560,N_15625);
nand U16080 (N_16080,N_15843,N_15923);
nor U16081 (N_16081,N_15667,N_15856);
and U16082 (N_16082,N_15500,N_15665);
xnor U16083 (N_16083,N_15551,N_15727);
nand U16084 (N_16084,N_15634,N_15824);
nand U16085 (N_16085,N_15565,N_15784);
nand U16086 (N_16086,N_15854,N_15846);
nand U16087 (N_16087,N_15895,N_15837);
nor U16088 (N_16088,N_15948,N_15569);
xnor U16089 (N_16089,N_15655,N_15704);
nand U16090 (N_16090,N_15700,N_15742);
and U16091 (N_16091,N_15822,N_15737);
and U16092 (N_16092,N_15886,N_15741);
or U16093 (N_16093,N_15878,N_15676);
nand U16094 (N_16094,N_15992,N_15508);
and U16095 (N_16095,N_15947,N_15723);
or U16096 (N_16096,N_15797,N_15597);
xnor U16097 (N_16097,N_15896,N_15652);
and U16098 (N_16098,N_15830,N_15869);
nor U16099 (N_16099,N_15795,N_15566);
nand U16100 (N_16100,N_15621,N_15562);
nor U16101 (N_16101,N_15609,N_15681);
xnor U16102 (N_16102,N_15773,N_15610);
or U16103 (N_16103,N_15707,N_15531);
or U16104 (N_16104,N_15775,N_15572);
or U16105 (N_16105,N_15618,N_15910);
or U16106 (N_16106,N_15847,N_15699);
or U16107 (N_16107,N_15711,N_15839);
or U16108 (N_16108,N_15601,N_15556);
and U16109 (N_16109,N_15542,N_15903);
or U16110 (N_16110,N_15907,N_15921);
nor U16111 (N_16111,N_15804,N_15932);
and U16112 (N_16112,N_15996,N_15664);
nor U16113 (N_16113,N_15997,N_15766);
nand U16114 (N_16114,N_15730,N_15891);
xor U16115 (N_16115,N_15811,N_15842);
nand U16116 (N_16116,N_15549,N_15624);
xor U16117 (N_16117,N_15779,N_15981);
and U16118 (N_16118,N_15507,N_15687);
nor U16119 (N_16119,N_15645,N_15844);
nand U16120 (N_16120,N_15501,N_15753);
nand U16121 (N_16121,N_15887,N_15834);
nor U16122 (N_16122,N_15809,N_15958);
nor U16123 (N_16123,N_15794,N_15726);
nand U16124 (N_16124,N_15688,N_15703);
nand U16125 (N_16125,N_15605,N_15827);
nand U16126 (N_16126,N_15657,N_15860);
nor U16127 (N_16127,N_15653,N_15835);
nor U16128 (N_16128,N_15579,N_15965);
nor U16129 (N_16129,N_15513,N_15881);
nand U16130 (N_16130,N_15914,N_15836);
nand U16131 (N_16131,N_15801,N_15826);
or U16132 (N_16132,N_15682,N_15582);
and U16133 (N_16133,N_15788,N_15789);
and U16134 (N_16134,N_15944,N_15745);
or U16135 (N_16135,N_15798,N_15931);
and U16136 (N_16136,N_15698,N_15980);
nand U16137 (N_16137,N_15899,N_15606);
nor U16138 (N_16138,N_15764,N_15829);
nor U16139 (N_16139,N_15977,N_15833);
nor U16140 (N_16140,N_15558,N_15587);
or U16141 (N_16141,N_15917,N_15685);
or U16142 (N_16142,N_15518,N_15516);
nand U16143 (N_16143,N_15633,N_15506);
or U16144 (N_16144,N_15754,N_15744);
nand U16145 (N_16145,N_15649,N_15889);
nor U16146 (N_16146,N_15939,N_15890);
nand U16147 (N_16147,N_15740,N_15928);
nor U16148 (N_16148,N_15530,N_15792);
and U16149 (N_16149,N_15529,N_15545);
or U16150 (N_16150,N_15849,N_15805);
nand U16151 (N_16151,N_15808,N_15969);
or U16152 (N_16152,N_15785,N_15962);
nor U16153 (N_16153,N_15922,N_15748);
nand U16154 (N_16154,N_15552,N_15790);
xnor U16155 (N_16155,N_15520,N_15592);
xnor U16156 (N_16156,N_15613,N_15813);
nor U16157 (N_16157,N_15924,N_15632);
and U16158 (N_16158,N_15728,N_15594);
nand U16159 (N_16159,N_15930,N_15739);
nand U16160 (N_16160,N_15706,N_15925);
or U16161 (N_16161,N_15679,N_15546);
nor U16162 (N_16162,N_15514,N_15774);
and U16163 (N_16163,N_15972,N_15736);
and U16164 (N_16164,N_15908,N_15692);
nor U16165 (N_16165,N_15503,N_15537);
nand U16166 (N_16166,N_15581,N_15850);
nand U16167 (N_16167,N_15526,N_15873);
or U16168 (N_16168,N_15662,N_15882);
nor U16169 (N_16169,N_15823,N_15963);
nor U16170 (N_16170,N_15853,N_15749);
or U16171 (N_16171,N_15995,N_15654);
nand U16172 (N_16172,N_15870,N_15988);
nor U16173 (N_16173,N_15984,N_15786);
and U16174 (N_16174,N_15825,N_15976);
nor U16175 (N_16175,N_15971,N_15724);
nor U16176 (N_16176,N_15608,N_15919);
nor U16177 (N_16177,N_15832,N_15979);
or U16178 (N_16178,N_15535,N_15761);
nor U16179 (N_16179,N_15555,N_15815);
nand U16180 (N_16180,N_15894,N_15575);
nand U16181 (N_16181,N_15689,N_15702);
nor U16182 (N_16182,N_15641,N_15945);
xor U16183 (N_16183,N_15807,N_15677);
nor U16184 (N_16184,N_15719,N_15865);
xor U16185 (N_16185,N_15638,N_15554);
or U16186 (N_16186,N_15817,N_15666);
or U16187 (N_16187,N_15532,N_15576);
nor U16188 (N_16188,N_15892,N_15717);
xor U16189 (N_16189,N_15956,N_15690);
nor U16190 (N_16190,N_15802,N_15620);
and U16191 (N_16191,N_15966,N_15880);
nand U16192 (N_16192,N_15777,N_15857);
nand U16193 (N_16193,N_15812,N_15705);
or U16194 (N_16194,N_15656,N_15611);
nand U16195 (N_16195,N_15615,N_15602);
nand U16196 (N_16196,N_15658,N_15781);
nand U16197 (N_16197,N_15940,N_15841);
nor U16198 (N_16198,N_15954,N_15573);
and U16199 (N_16199,N_15623,N_15767);
nand U16200 (N_16200,N_15993,N_15522);
or U16201 (N_16201,N_15643,N_15511);
and U16202 (N_16202,N_15964,N_15539);
or U16203 (N_16203,N_15960,N_15952);
and U16204 (N_16204,N_15793,N_15911);
and U16205 (N_16205,N_15540,N_15986);
or U16206 (N_16206,N_15617,N_15937);
nor U16207 (N_16207,N_15864,N_15912);
or U16208 (N_16208,N_15599,N_15929);
nor U16209 (N_16209,N_15629,N_15524);
and U16210 (N_16210,N_15714,N_15708);
xnor U16211 (N_16211,N_15559,N_15637);
and U16212 (N_16212,N_15543,N_15734);
nor U16213 (N_16213,N_15515,N_15743);
or U16214 (N_16214,N_15927,N_15852);
and U16215 (N_16215,N_15796,N_15985);
or U16216 (N_16216,N_15871,N_15760);
or U16217 (N_16217,N_15787,N_15780);
and U16218 (N_16218,N_15799,N_15510);
and U16219 (N_16219,N_15738,N_15670);
nor U16220 (N_16220,N_15776,N_15897);
nor U16221 (N_16221,N_15936,N_15701);
nand U16222 (N_16222,N_15762,N_15987);
xor U16223 (N_16223,N_15557,N_15553);
xnor U16224 (N_16224,N_15916,N_15504);
and U16225 (N_16225,N_15580,N_15967);
or U16226 (N_16226,N_15772,N_15975);
or U16227 (N_16227,N_15861,N_15893);
and U16228 (N_16228,N_15527,N_15642);
xnor U16229 (N_16229,N_15920,N_15735);
xor U16230 (N_16230,N_15564,N_15970);
or U16231 (N_16231,N_15872,N_15994);
nand U16232 (N_16232,N_15712,N_15533);
nor U16233 (N_16233,N_15646,N_15758);
nand U16234 (N_16234,N_15721,N_15883);
nor U16235 (N_16235,N_15716,N_15525);
and U16236 (N_16236,N_15651,N_15683);
or U16237 (N_16237,N_15563,N_15732);
or U16238 (N_16238,N_15693,N_15803);
xnor U16239 (N_16239,N_15983,N_15953);
and U16240 (N_16240,N_15941,N_15974);
nand U16241 (N_16241,N_15509,N_15715);
nor U16242 (N_16242,N_15867,N_15978);
or U16243 (N_16243,N_15591,N_15669);
nor U16244 (N_16244,N_15574,N_15831);
and U16245 (N_16245,N_15595,N_15828);
nor U16246 (N_16246,N_15938,N_15571);
nor U16247 (N_16247,N_15991,N_15990);
xnor U16248 (N_16248,N_15961,N_15648);
nand U16249 (N_16249,N_15879,N_15943);
xor U16250 (N_16250,N_15504,N_15518);
or U16251 (N_16251,N_15604,N_15521);
or U16252 (N_16252,N_15580,N_15939);
nor U16253 (N_16253,N_15760,N_15646);
nor U16254 (N_16254,N_15726,N_15554);
and U16255 (N_16255,N_15900,N_15667);
xnor U16256 (N_16256,N_15718,N_15537);
and U16257 (N_16257,N_15626,N_15551);
nor U16258 (N_16258,N_15591,N_15837);
or U16259 (N_16259,N_15996,N_15621);
and U16260 (N_16260,N_15869,N_15976);
xor U16261 (N_16261,N_15829,N_15754);
and U16262 (N_16262,N_15718,N_15523);
and U16263 (N_16263,N_15927,N_15920);
nor U16264 (N_16264,N_15695,N_15752);
or U16265 (N_16265,N_15708,N_15896);
nor U16266 (N_16266,N_15561,N_15696);
and U16267 (N_16267,N_15890,N_15662);
nor U16268 (N_16268,N_15504,N_15953);
or U16269 (N_16269,N_15536,N_15800);
and U16270 (N_16270,N_15500,N_15674);
nand U16271 (N_16271,N_15668,N_15878);
nand U16272 (N_16272,N_15901,N_15973);
and U16273 (N_16273,N_15509,N_15651);
nand U16274 (N_16274,N_15606,N_15962);
nand U16275 (N_16275,N_15782,N_15830);
nand U16276 (N_16276,N_15866,N_15846);
and U16277 (N_16277,N_15689,N_15886);
nand U16278 (N_16278,N_15950,N_15921);
nand U16279 (N_16279,N_15821,N_15562);
and U16280 (N_16280,N_15942,N_15595);
or U16281 (N_16281,N_15669,N_15680);
or U16282 (N_16282,N_15671,N_15710);
xnor U16283 (N_16283,N_15522,N_15680);
or U16284 (N_16284,N_15547,N_15823);
nor U16285 (N_16285,N_15598,N_15691);
or U16286 (N_16286,N_15632,N_15557);
nand U16287 (N_16287,N_15914,N_15868);
or U16288 (N_16288,N_15747,N_15979);
nor U16289 (N_16289,N_15895,N_15500);
and U16290 (N_16290,N_15561,N_15646);
nand U16291 (N_16291,N_15659,N_15796);
and U16292 (N_16292,N_15960,N_15734);
nor U16293 (N_16293,N_15916,N_15900);
nand U16294 (N_16294,N_15779,N_15679);
or U16295 (N_16295,N_15676,N_15927);
or U16296 (N_16296,N_15622,N_15534);
nand U16297 (N_16297,N_15957,N_15782);
and U16298 (N_16298,N_15962,N_15707);
or U16299 (N_16299,N_15580,N_15875);
nor U16300 (N_16300,N_15746,N_15761);
nor U16301 (N_16301,N_15728,N_15651);
nand U16302 (N_16302,N_15664,N_15742);
or U16303 (N_16303,N_15861,N_15686);
xnor U16304 (N_16304,N_15858,N_15729);
xnor U16305 (N_16305,N_15774,N_15724);
nor U16306 (N_16306,N_15760,N_15896);
xor U16307 (N_16307,N_15567,N_15972);
and U16308 (N_16308,N_15722,N_15532);
nor U16309 (N_16309,N_15508,N_15627);
nor U16310 (N_16310,N_15922,N_15764);
nor U16311 (N_16311,N_15880,N_15727);
nand U16312 (N_16312,N_15976,N_15905);
and U16313 (N_16313,N_15529,N_15845);
or U16314 (N_16314,N_15870,N_15590);
or U16315 (N_16315,N_15788,N_15974);
and U16316 (N_16316,N_15755,N_15794);
and U16317 (N_16317,N_15628,N_15845);
nor U16318 (N_16318,N_15876,N_15690);
xnor U16319 (N_16319,N_15846,N_15540);
and U16320 (N_16320,N_15919,N_15748);
nand U16321 (N_16321,N_15937,N_15780);
and U16322 (N_16322,N_15927,N_15844);
xor U16323 (N_16323,N_15789,N_15996);
xnor U16324 (N_16324,N_15872,N_15637);
or U16325 (N_16325,N_15832,N_15581);
nor U16326 (N_16326,N_15530,N_15873);
nor U16327 (N_16327,N_15962,N_15869);
and U16328 (N_16328,N_15865,N_15927);
nand U16329 (N_16329,N_15530,N_15772);
nor U16330 (N_16330,N_15841,N_15538);
or U16331 (N_16331,N_15600,N_15546);
or U16332 (N_16332,N_15865,N_15957);
nand U16333 (N_16333,N_15861,N_15521);
nor U16334 (N_16334,N_15711,N_15993);
or U16335 (N_16335,N_15624,N_15644);
nor U16336 (N_16336,N_15744,N_15632);
nor U16337 (N_16337,N_15995,N_15517);
nor U16338 (N_16338,N_15509,N_15811);
nor U16339 (N_16339,N_15747,N_15706);
or U16340 (N_16340,N_15676,N_15647);
nor U16341 (N_16341,N_15889,N_15897);
or U16342 (N_16342,N_15685,N_15752);
or U16343 (N_16343,N_15516,N_15539);
and U16344 (N_16344,N_15751,N_15819);
xnor U16345 (N_16345,N_15817,N_15808);
nand U16346 (N_16346,N_15909,N_15623);
xor U16347 (N_16347,N_15790,N_15945);
and U16348 (N_16348,N_15556,N_15796);
or U16349 (N_16349,N_15546,N_15836);
and U16350 (N_16350,N_15882,N_15679);
nand U16351 (N_16351,N_15739,N_15793);
nor U16352 (N_16352,N_15815,N_15821);
or U16353 (N_16353,N_15897,N_15501);
nor U16354 (N_16354,N_15922,N_15934);
or U16355 (N_16355,N_15968,N_15953);
or U16356 (N_16356,N_15967,N_15884);
nand U16357 (N_16357,N_15918,N_15835);
nor U16358 (N_16358,N_15684,N_15924);
xnor U16359 (N_16359,N_15888,N_15788);
nor U16360 (N_16360,N_15898,N_15914);
nor U16361 (N_16361,N_15790,N_15901);
nand U16362 (N_16362,N_15655,N_15544);
or U16363 (N_16363,N_15532,N_15583);
and U16364 (N_16364,N_15985,N_15938);
xnor U16365 (N_16365,N_15525,N_15683);
xor U16366 (N_16366,N_15829,N_15535);
or U16367 (N_16367,N_15930,N_15629);
xor U16368 (N_16368,N_15976,N_15666);
and U16369 (N_16369,N_15789,N_15962);
nand U16370 (N_16370,N_15793,N_15605);
and U16371 (N_16371,N_15558,N_15979);
nand U16372 (N_16372,N_15730,N_15665);
nand U16373 (N_16373,N_15760,N_15786);
or U16374 (N_16374,N_15507,N_15836);
nand U16375 (N_16375,N_15665,N_15650);
nor U16376 (N_16376,N_15616,N_15805);
and U16377 (N_16377,N_15999,N_15872);
or U16378 (N_16378,N_15669,N_15529);
and U16379 (N_16379,N_15620,N_15930);
nor U16380 (N_16380,N_15544,N_15986);
xor U16381 (N_16381,N_15760,N_15865);
nand U16382 (N_16382,N_15639,N_15767);
or U16383 (N_16383,N_15840,N_15510);
and U16384 (N_16384,N_15724,N_15814);
and U16385 (N_16385,N_15710,N_15640);
nor U16386 (N_16386,N_15633,N_15567);
or U16387 (N_16387,N_15867,N_15766);
or U16388 (N_16388,N_15915,N_15737);
xnor U16389 (N_16389,N_15636,N_15680);
and U16390 (N_16390,N_15845,N_15855);
or U16391 (N_16391,N_15647,N_15602);
and U16392 (N_16392,N_15603,N_15857);
and U16393 (N_16393,N_15909,N_15638);
xnor U16394 (N_16394,N_15990,N_15621);
or U16395 (N_16395,N_15944,N_15675);
nor U16396 (N_16396,N_15921,N_15653);
xor U16397 (N_16397,N_15502,N_15555);
or U16398 (N_16398,N_15897,N_15735);
nand U16399 (N_16399,N_15887,N_15976);
or U16400 (N_16400,N_15784,N_15577);
nand U16401 (N_16401,N_15585,N_15687);
nand U16402 (N_16402,N_15987,N_15800);
nand U16403 (N_16403,N_15970,N_15816);
and U16404 (N_16404,N_15754,N_15573);
nor U16405 (N_16405,N_15574,N_15747);
and U16406 (N_16406,N_15598,N_15917);
or U16407 (N_16407,N_15616,N_15929);
or U16408 (N_16408,N_15534,N_15633);
and U16409 (N_16409,N_15719,N_15589);
and U16410 (N_16410,N_15740,N_15594);
nor U16411 (N_16411,N_15783,N_15687);
and U16412 (N_16412,N_15501,N_15780);
and U16413 (N_16413,N_15608,N_15896);
xor U16414 (N_16414,N_15707,N_15862);
nor U16415 (N_16415,N_15650,N_15704);
nor U16416 (N_16416,N_15943,N_15527);
nand U16417 (N_16417,N_15965,N_15881);
and U16418 (N_16418,N_15686,N_15695);
nor U16419 (N_16419,N_15745,N_15899);
and U16420 (N_16420,N_15741,N_15939);
and U16421 (N_16421,N_15522,N_15631);
xor U16422 (N_16422,N_15842,N_15734);
nor U16423 (N_16423,N_15629,N_15980);
and U16424 (N_16424,N_15542,N_15931);
nand U16425 (N_16425,N_15705,N_15610);
xnor U16426 (N_16426,N_15532,N_15881);
and U16427 (N_16427,N_15818,N_15509);
nand U16428 (N_16428,N_15687,N_15952);
nand U16429 (N_16429,N_15874,N_15974);
nor U16430 (N_16430,N_15585,N_15642);
or U16431 (N_16431,N_15601,N_15771);
nand U16432 (N_16432,N_15567,N_15882);
and U16433 (N_16433,N_15553,N_15983);
or U16434 (N_16434,N_15780,N_15661);
or U16435 (N_16435,N_15501,N_15958);
nand U16436 (N_16436,N_15957,N_15964);
or U16437 (N_16437,N_15972,N_15520);
nor U16438 (N_16438,N_15825,N_15813);
and U16439 (N_16439,N_15621,N_15639);
nor U16440 (N_16440,N_15918,N_15886);
nor U16441 (N_16441,N_15856,N_15761);
and U16442 (N_16442,N_15969,N_15792);
or U16443 (N_16443,N_15549,N_15501);
nor U16444 (N_16444,N_15524,N_15913);
and U16445 (N_16445,N_15745,N_15947);
or U16446 (N_16446,N_15808,N_15662);
nor U16447 (N_16447,N_15783,N_15762);
nor U16448 (N_16448,N_15840,N_15591);
and U16449 (N_16449,N_15877,N_15924);
or U16450 (N_16450,N_15763,N_15946);
or U16451 (N_16451,N_15811,N_15544);
nand U16452 (N_16452,N_15532,N_15946);
or U16453 (N_16453,N_15896,N_15604);
nor U16454 (N_16454,N_15855,N_15946);
nor U16455 (N_16455,N_15870,N_15910);
nor U16456 (N_16456,N_15891,N_15525);
nor U16457 (N_16457,N_15914,N_15590);
nand U16458 (N_16458,N_15757,N_15663);
and U16459 (N_16459,N_15625,N_15677);
and U16460 (N_16460,N_15820,N_15904);
nand U16461 (N_16461,N_15599,N_15722);
nor U16462 (N_16462,N_15766,N_15869);
xnor U16463 (N_16463,N_15531,N_15803);
xor U16464 (N_16464,N_15875,N_15691);
and U16465 (N_16465,N_15715,N_15908);
or U16466 (N_16466,N_15747,N_15983);
or U16467 (N_16467,N_15890,N_15550);
nand U16468 (N_16468,N_15864,N_15596);
and U16469 (N_16469,N_15710,N_15972);
nor U16470 (N_16470,N_15660,N_15742);
or U16471 (N_16471,N_15803,N_15528);
and U16472 (N_16472,N_15908,N_15779);
and U16473 (N_16473,N_15528,N_15513);
nand U16474 (N_16474,N_15622,N_15675);
nor U16475 (N_16475,N_15865,N_15652);
nor U16476 (N_16476,N_15731,N_15717);
xor U16477 (N_16477,N_15833,N_15657);
and U16478 (N_16478,N_15839,N_15731);
and U16479 (N_16479,N_15965,N_15560);
or U16480 (N_16480,N_15753,N_15707);
nand U16481 (N_16481,N_15642,N_15669);
and U16482 (N_16482,N_15829,N_15882);
nor U16483 (N_16483,N_15641,N_15718);
or U16484 (N_16484,N_15769,N_15522);
or U16485 (N_16485,N_15779,N_15569);
nor U16486 (N_16486,N_15864,N_15739);
or U16487 (N_16487,N_15862,N_15680);
nand U16488 (N_16488,N_15978,N_15864);
or U16489 (N_16489,N_15512,N_15692);
and U16490 (N_16490,N_15828,N_15677);
xor U16491 (N_16491,N_15657,N_15512);
nand U16492 (N_16492,N_15576,N_15773);
and U16493 (N_16493,N_15964,N_15568);
nand U16494 (N_16494,N_15529,N_15607);
and U16495 (N_16495,N_15587,N_15682);
nand U16496 (N_16496,N_15635,N_15785);
and U16497 (N_16497,N_15802,N_15555);
nand U16498 (N_16498,N_15793,N_15626);
nor U16499 (N_16499,N_15770,N_15916);
nand U16500 (N_16500,N_16211,N_16230);
or U16501 (N_16501,N_16409,N_16289);
and U16502 (N_16502,N_16003,N_16036);
nand U16503 (N_16503,N_16376,N_16018);
nand U16504 (N_16504,N_16461,N_16214);
nand U16505 (N_16505,N_16467,N_16206);
or U16506 (N_16506,N_16380,N_16255);
or U16507 (N_16507,N_16382,N_16043);
or U16508 (N_16508,N_16087,N_16383);
nand U16509 (N_16509,N_16299,N_16292);
and U16510 (N_16510,N_16011,N_16294);
and U16511 (N_16511,N_16121,N_16209);
nor U16512 (N_16512,N_16095,N_16260);
or U16513 (N_16513,N_16414,N_16207);
or U16514 (N_16514,N_16009,N_16212);
or U16515 (N_16515,N_16397,N_16429);
or U16516 (N_16516,N_16188,N_16102);
nand U16517 (N_16517,N_16477,N_16218);
and U16518 (N_16518,N_16424,N_16028);
xor U16519 (N_16519,N_16071,N_16059);
nor U16520 (N_16520,N_16280,N_16172);
nand U16521 (N_16521,N_16042,N_16193);
and U16522 (N_16522,N_16189,N_16181);
nor U16523 (N_16523,N_16323,N_16040);
or U16524 (N_16524,N_16064,N_16106);
nor U16525 (N_16525,N_16030,N_16486);
and U16526 (N_16526,N_16034,N_16275);
and U16527 (N_16527,N_16041,N_16026);
or U16528 (N_16528,N_16229,N_16139);
or U16529 (N_16529,N_16201,N_16163);
xnor U16530 (N_16530,N_16145,N_16360);
and U16531 (N_16531,N_16318,N_16354);
or U16532 (N_16532,N_16476,N_16090);
nor U16533 (N_16533,N_16479,N_16012);
xor U16534 (N_16534,N_16287,N_16123);
nand U16535 (N_16535,N_16398,N_16478);
and U16536 (N_16536,N_16343,N_16438);
and U16537 (N_16537,N_16044,N_16290);
and U16538 (N_16538,N_16452,N_16325);
and U16539 (N_16539,N_16497,N_16241);
and U16540 (N_16540,N_16270,N_16352);
and U16541 (N_16541,N_16279,N_16025);
nor U16542 (N_16542,N_16413,N_16334);
and U16543 (N_16543,N_16154,N_16156);
nand U16544 (N_16544,N_16445,N_16359);
and U16545 (N_16545,N_16494,N_16308);
and U16546 (N_16546,N_16342,N_16276);
nor U16547 (N_16547,N_16311,N_16456);
or U16548 (N_16548,N_16235,N_16069);
nand U16549 (N_16549,N_16174,N_16115);
xor U16550 (N_16550,N_16305,N_16084);
and U16551 (N_16551,N_16273,N_16459);
nand U16552 (N_16552,N_16444,N_16331);
nor U16553 (N_16553,N_16132,N_16286);
or U16554 (N_16554,N_16135,N_16379);
or U16555 (N_16555,N_16387,N_16415);
or U16556 (N_16556,N_16245,N_16081);
xor U16557 (N_16557,N_16265,N_16303);
nor U16558 (N_16558,N_16021,N_16107);
and U16559 (N_16559,N_16431,N_16262);
nand U16560 (N_16560,N_16017,N_16237);
xnor U16561 (N_16561,N_16392,N_16184);
or U16562 (N_16562,N_16449,N_16243);
and U16563 (N_16563,N_16490,N_16460);
nor U16564 (N_16564,N_16264,N_16086);
or U16565 (N_16565,N_16162,N_16187);
xnor U16566 (N_16566,N_16420,N_16465);
or U16567 (N_16567,N_16313,N_16196);
nand U16568 (N_16568,N_16428,N_16105);
or U16569 (N_16569,N_16134,N_16129);
xnor U16570 (N_16570,N_16151,N_16083);
nor U16571 (N_16571,N_16089,N_16422);
and U16572 (N_16572,N_16390,N_16101);
and U16573 (N_16573,N_16402,N_16124);
or U16574 (N_16574,N_16351,N_16216);
xor U16575 (N_16575,N_16329,N_16203);
and U16576 (N_16576,N_16116,N_16246);
nor U16577 (N_16577,N_16407,N_16070);
nand U16578 (N_16578,N_16498,N_16088);
xnor U16579 (N_16579,N_16263,N_16386);
xor U16580 (N_16580,N_16073,N_16450);
or U16581 (N_16581,N_16222,N_16335);
and U16582 (N_16582,N_16148,N_16256);
nand U16583 (N_16583,N_16100,N_16253);
xor U16584 (N_16584,N_16370,N_16147);
nor U16585 (N_16585,N_16142,N_16098);
nor U16586 (N_16586,N_16330,N_16136);
nor U16587 (N_16587,N_16391,N_16179);
nand U16588 (N_16588,N_16492,N_16037);
nor U16589 (N_16589,N_16340,N_16175);
xnor U16590 (N_16590,N_16261,N_16371);
and U16591 (N_16591,N_16050,N_16168);
or U16592 (N_16592,N_16078,N_16339);
nand U16593 (N_16593,N_16117,N_16099);
or U16594 (N_16594,N_16451,N_16125);
nand U16595 (N_16595,N_16271,N_16378);
nand U16596 (N_16596,N_16297,N_16358);
nor U16597 (N_16597,N_16423,N_16144);
nor U16598 (N_16598,N_16307,N_16048);
nor U16599 (N_16599,N_16401,N_16150);
nand U16600 (N_16600,N_16249,N_16205);
or U16601 (N_16601,N_16075,N_16404);
nand U16602 (N_16602,N_16257,N_16433);
nand U16603 (N_16603,N_16067,N_16356);
xnor U16604 (N_16604,N_16227,N_16362);
nand U16605 (N_16605,N_16439,N_16074);
or U16606 (N_16606,N_16332,N_16014);
xor U16607 (N_16607,N_16137,N_16412);
and U16608 (N_16608,N_16233,N_16473);
and U16609 (N_16609,N_16155,N_16349);
or U16610 (N_16610,N_16242,N_16298);
or U16611 (N_16611,N_16295,N_16114);
nand U16612 (N_16612,N_16060,N_16062);
and U16613 (N_16613,N_16344,N_16244);
or U16614 (N_16614,N_16493,N_16015);
and U16615 (N_16615,N_16384,N_16027);
nor U16616 (N_16616,N_16023,N_16381);
and U16617 (N_16617,N_16133,N_16008);
and U16618 (N_16618,N_16177,N_16464);
nor U16619 (N_16619,N_16259,N_16058);
and U16620 (N_16620,N_16314,N_16063);
nor U16621 (N_16621,N_16369,N_16210);
nor U16622 (N_16622,N_16388,N_16056);
nor U16623 (N_16623,N_16171,N_16283);
nand U16624 (N_16624,N_16327,N_16000);
nor U16625 (N_16625,N_16110,N_16337);
nand U16626 (N_16626,N_16466,N_16010);
or U16627 (N_16627,N_16096,N_16453);
nor U16628 (N_16628,N_16143,N_16483);
xnor U16629 (N_16629,N_16239,N_16372);
or U16630 (N_16630,N_16045,N_16104);
nor U16631 (N_16631,N_16421,N_16321);
or U16632 (N_16632,N_16394,N_16302);
nor U16633 (N_16633,N_16085,N_16190);
nand U16634 (N_16634,N_16247,N_16232);
nor U16635 (N_16635,N_16068,N_16169);
and U16636 (N_16636,N_16033,N_16441);
nand U16637 (N_16637,N_16443,N_16411);
xnor U16638 (N_16638,N_16204,N_16454);
nand U16639 (N_16639,N_16251,N_16375);
nand U16640 (N_16640,N_16170,N_16317);
xnor U16641 (N_16641,N_16474,N_16426);
and U16642 (N_16642,N_16178,N_16066);
nor U16643 (N_16643,N_16248,N_16215);
xor U16644 (N_16644,N_16208,N_16319);
or U16645 (N_16645,N_16495,N_16480);
nor U16646 (N_16646,N_16430,N_16425);
nor U16647 (N_16647,N_16320,N_16268);
or U16648 (N_16648,N_16119,N_16161);
and U16649 (N_16649,N_16468,N_16140);
nand U16650 (N_16650,N_16442,N_16182);
or U16651 (N_16651,N_16019,N_16437);
or U16652 (N_16652,N_16225,N_16032);
nand U16653 (N_16653,N_16173,N_16219);
nor U16654 (N_16654,N_16291,N_16475);
and U16655 (N_16655,N_16434,N_16355);
xor U16656 (N_16656,N_16346,N_16361);
xor U16657 (N_16657,N_16158,N_16373);
nand U16658 (N_16658,N_16293,N_16304);
nor U16659 (N_16659,N_16416,N_16024);
or U16660 (N_16660,N_16228,N_16353);
or U16661 (N_16661,N_16146,N_16427);
nand U16662 (N_16662,N_16336,N_16252);
xnor U16663 (N_16663,N_16051,N_16258);
nand U16664 (N_16664,N_16231,N_16489);
or U16665 (N_16665,N_16418,N_16417);
nor U16666 (N_16666,N_16274,N_16395);
nand U16667 (N_16667,N_16213,N_16300);
and U16668 (N_16668,N_16013,N_16006);
or U16669 (N_16669,N_16191,N_16152);
nand U16670 (N_16670,N_16122,N_16192);
xnor U16671 (N_16671,N_16164,N_16345);
nand U16672 (N_16672,N_16350,N_16016);
and U16673 (N_16673,N_16315,N_16326);
xor U16674 (N_16674,N_16496,N_16223);
xor U16675 (N_16675,N_16022,N_16367);
nor U16676 (N_16676,N_16296,N_16250);
nand U16677 (N_16677,N_16254,N_16316);
and U16678 (N_16678,N_16202,N_16185);
xnor U16679 (N_16679,N_16131,N_16004);
nand U16680 (N_16680,N_16054,N_16385);
nand U16681 (N_16681,N_16167,N_16029);
and U16682 (N_16682,N_16093,N_16092);
xor U16683 (N_16683,N_16130,N_16183);
nor U16684 (N_16684,N_16138,N_16103);
and U16685 (N_16685,N_16488,N_16272);
nand U16686 (N_16686,N_16079,N_16128);
xor U16687 (N_16687,N_16111,N_16091);
and U16688 (N_16688,N_16472,N_16338);
nor U16689 (N_16689,N_16126,N_16047);
xnor U16690 (N_16690,N_16341,N_16447);
nor U16691 (N_16691,N_16240,N_16076);
or U16692 (N_16692,N_16482,N_16324);
xnor U16693 (N_16693,N_16002,N_16436);
or U16694 (N_16694,N_16234,N_16057);
nand U16695 (N_16695,N_16396,N_16469);
and U16696 (N_16696,N_16389,N_16108);
nor U16697 (N_16697,N_16288,N_16348);
or U16698 (N_16698,N_16186,N_16374);
xor U16699 (N_16699,N_16306,N_16109);
nand U16700 (N_16700,N_16127,N_16470);
and U16701 (N_16701,N_16072,N_16277);
and U16702 (N_16702,N_16403,N_16065);
xnor U16703 (N_16703,N_16357,N_16267);
or U16704 (N_16704,N_16052,N_16405);
or U16705 (N_16705,N_16097,N_16157);
nand U16706 (N_16706,N_16053,N_16408);
nand U16707 (N_16707,N_16238,N_16365);
and U16708 (N_16708,N_16094,N_16285);
nand U16709 (N_16709,N_16165,N_16195);
and U16710 (N_16710,N_16446,N_16120);
nor U16711 (N_16711,N_16406,N_16118);
xnor U16712 (N_16712,N_16322,N_16455);
and U16713 (N_16713,N_16159,N_16035);
and U16714 (N_16714,N_16347,N_16061);
nor U16715 (N_16715,N_16200,N_16199);
nor U16716 (N_16716,N_16194,N_16220);
nand U16717 (N_16717,N_16463,N_16419);
and U16718 (N_16718,N_16366,N_16221);
nor U16719 (N_16719,N_16435,N_16236);
nand U16720 (N_16720,N_16400,N_16432);
nand U16721 (N_16721,N_16471,N_16457);
or U16722 (N_16722,N_16180,N_16410);
and U16723 (N_16723,N_16007,N_16393);
nor U16724 (N_16724,N_16039,N_16364);
or U16725 (N_16725,N_16197,N_16082);
or U16726 (N_16726,N_16038,N_16266);
nand U16727 (N_16727,N_16458,N_16462);
nor U16728 (N_16728,N_16328,N_16224);
nand U16729 (N_16729,N_16284,N_16481);
or U16730 (N_16730,N_16080,N_16363);
or U16731 (N_16731,N_16020,N_16487);
nand U16732 (N_16732,N_16484,N_16440);
or U16733 (N_16733,N_16368,N_16141);
or U16734 (N_16734,N_16149,N_16160);
or U16735 (N_16735,N_16448,N_16153);
nor U16736 (N_16736,N_16217,N_16166);
xor U16737 (N_16737,N_16269,N_16399);
nand U16738 (N_16738,N_16046,N_16499);
and U16739 (N_16739,N_16001,N_16491);
nor U16740 (N_16740,N_16310,N_16198);
nand U16741 (N_16741,N_16055,N_16309);
or U16742 (N_16742,N_16485,N_16112);
nor U16743 (N_16743,N_16113,N_16312);
nor U16744 (N_16744,N_16049,N_16077);
or U16745 (N_16745,N_16377,N_16333);
nor U16746 (N_16746,N_16226,N_16005);
and U16747 (N_16747,N_16278,N_16031);
nand U16748 (N_16748,N_16301,N_16282);
or U16749 (N_16749,N_16281,N_16176);
nand U16750 (N_16750,N_16255,N_16490);
xnor U16751 (N_16751,N_16131,N_16141);
and U16752 (N_16752,N_16123,N_16029);
and U16753 (N_16753,N_16114,N_16484);
and U16754 (N_16754,N_16186,N_16477);
and U16755 (N_16755,N_16273,N_16241);
and U16756 (N_16756,N_16413,N_16080);
nand U16757 (N_16757,N_16266,N_16061);
nor U16758 (N_16758,N_16256,N_16084);
and U16759 (N_16759,N_16423,N_16186);
and U16760 (N_16760,N_16018,N_16357);
and U16761 (N_16761,N_16027,N_16024);
and U16762 (N_16762,N_16366,N_16020);
nor U16763 (N_16763,N_16335,N_16065);
nand U16764 (N_16764,N_16492,N_16439);
xor U16765 (N_16765,N_16044,N_16478);
xor U16766 (N_16766,N_16402,N_16125);
and U16767 (N_16767,N_16226,N_16178);
or U16768 (N_16768,N_16471,N_16316);
xor U16769 (N_16769,N_16380,N_16274);
or U16770 (N_16770,N_16296,N_16348);
nand U16771 (N_16771,N_16348,N_16157);
nand U16772 (N_16772,N_16450,N_16249);
and U16773 (N_16773,N_16012,N_16289);
or U16774 (N_16774,N_16414,N_16293);
xor U16775 (N_16775,N_16322,N_16274);
nor U16776 (N_16776,N_16290,N_16477);
nand U16777 (N_16777,N_16483,N_16105);
or U16778 (N_16778,N_16394,N_16447);
or U16779 (N_16779,N_16354,N_16014);
or U16780 (N_16780,N_16116,N_16335);
nor U16781 (N_16781,N_16446,N_16156);
or U16782 (N_16782,N_16331,N_16418);
or U16783 (N_16783,N_16099,N_16374);
nor U16784 (N_16784,N_16166,N_16051);
nor U16785 (N_16785,N_16424,N_16068);
or U16786 (N_16786,N_16264,N_16115);
or U16787 (N_16787,N_16003,N_16071);
or U16788 (N_16788,N_16182,N_16070);
and U16789 (N_16789,N_16400,N_16331);
nand U16790 (N_16790,N_16483,N_16079);
and U16791 (N_16791,N_16356,N_16252);
nor U16792 (N_16792,N_16450,N_16472);
nor U16793 (N_16793,N_16329,N_16443);
or U16794 (N_16794,N_16267,N_16446);
nor U16795 (N_16795,N_16397,N_16104);
nand U16796 (N_16796,N_16144,N_16017);
nand U16797 (N_16797,N_16079,N_16494);
nor U16798 (N_16798,N_16020,N_16231);
xor U16799 (N_16799,N_16121,N_16480);
or U16800 (N_16800,N_16242,N_16364);
nand U16801 (N_16801,N_16153,N_16188);
or U16802 (N_16802,N_16363,N_16071);
or U16803 (N_16803,N_16329,N_16226);
nor U16804 (N_16804,N_16491,N_16379);
xor U16805 (N_16805,N_16420,N_16240);
and U16806 (N_16806,N_16236,N_16097);
or U16807 (N_16807,N_16432,N_16061);
nand U16808 (N_16808,N_16390,N_16132);
and U16809 (N_16809,N_16083,N_16289);
and U16810 (N_16810,N_16441,N_16046);
nor U16811 (N_16811,N_16035,N_16484);
and U16812 (N_16812,N_16468,N_16100);
or U16813 (N_16813,N_16364,N_16177);
nand U16814 (N_16814,N_16079,N_16259);
nand U16815 (N_16815,N_16269,N_16198);
and U16816 (N_16816,N_16031,N_16281);
xor U16817 (N_16817,N_16060,N_16266);
and U16818 (N_16818,N_16422,N_16232);
or U16819 (N_16819,N_16131,N_16459);
nand U16820 (N_16820,N_16435,N_16023);
nand U16821 (N_16821,N_16319,N_16405);
and U16822 (N_16822,N_16308,N_16057);
nor U16823 (N_16823,N_16060,N_16282);
nor U16824 (N_16824,N_16185,N_16380);
nand U16825 (N_16825,N_16220,N_16053);
nand U16826 (N_16826,N_16010,N_16299);
nand U16827 (N_16827,N_16249,N_16018);
nand U16828 (N_16828,N_16169,N_16079);
xnor U16829 (N_16829,N_16309,N_16059);
or U16830 (N_16830,N_16480,N_16209);
nand U16831 (N_16831,N_16337,N_16152);
or U16832 (N_16832,N_16070,N_16461);
and U16833 (N_16833,N_16474,N_16047);
nand U16834 (N_16834,N_16342,N_16036);
or U16835 (N_16835,N_16413,N_16298);
xor U16836 (N_16836,N_16423,N_16115);
xnor U16837 (N_16837,N_16134,N_16436);
or U16838 (N_16838,N_16045,N_16198);
nand U16839 (N_16839,N_16190,N_16127);
xor U16840 (N_16840,N_16015,N_16404);
or U16841 (N_16841,N_16039,N_16360);
nand U16842 (N_16842,N_16156,N_16165);
or U16843 (N_16843,N_16496,N_16005);
and U16844 (N_16844,N_16301,N_16025);
and U16845 (N_16845,N_16379,N_16161);
and U16846 (N_16846,N_16217,N_16329);
nor U16847 (N_16847,N_16202,N_16407);
and U16848 (N_16848,N_16243,N_16050);
and U16849 (N_16849,N_16466,N_16196);
xnor U16850 (N_16850,N_16212,N_16473);
nor U16851 (N_16851,N_16033,N_16297);
or U16852 (N_16852,N_16106,N_16385);
nand U16853 (N_16853,N_16433,N_16436);
and U16854 (N_16854,N_16213,N_16084);
nor U16855 (N_16855,N_16026,N_16136);
nand U16856 (N_16856,N_16012,N_16107);
nand U16857 (N_16857,N_16273,N_16006);
and U16858 (N_16858,N_16268,N_16276);
and U16859 (N_16859,N_16222,N_16458);
nand U16860 (N_16860,N_16493,N_16430);
and U16861 (N_16861,N_16332,N_16126);
and U16862 (N_16862,N_16428,N_16004);
xnor U16863 (N_16863,N_16177,N_16211);
nor U16864 (N_16864,N_16167,N_16368);
or U16865 (N_16865,N_16358,N_16176);
xor U16866 (N_16866,N_16291,N_16371);
nand U16867 (N_16867,N_16421,N_16222);
and U16868 (N_16868,N_16362,N_16242);
or U16869 (N_16869,N_16191,N_16051);
or U16870 (N_16870,N_16222,N_16384);
and U16871 (N_16871,N_16224,N_16398);
nor U16872 (N_16872,N_16281,N_16036);
or U16873 (N_16873,N_16310,N_16389);
nor U16874 (N_16874,N_16201,N_16017);
xor U16875 (N_16875,N_16357,N_16036);
nor U16876 (N_16876,N_16379,N_16208);
nor U16877 (N_16877,N_16014,N_16027);
nand U16878 (N_16878,N_16468,N_16141);
xor U16879 (N_16879,N_16418,N_16442);
and U16880 (N_16880,N_16266,N_16496);
nand U16881 (N_16881,N_16136,N_16420);
nor U16882 (N_16882,N_16473,N_16097);
and U16883 (N_16883,N_16104,N_16236);
and U16884 (N_16884,N_16263,N_16428);
nand U16885 (N_16885,N_16433,N_16304);
xnor U16886 (N_16886,N_16275,N_16049);
nand U16887 (N_16887,N_16258,N_16431);
nand U16888 (N_16888,N_16168,N_16153);
or U16889 (N_16889,N_16432,N_16113);
nand U16890 (N_16890,N_16262,N_16142);
and U16891 (N_16891,N_16161,N_16496);
nor U16892 (N_16892,N_16199,N_16458);
or U16893 (N_16893,N_16264,N_16342);
or U16894 (N_16894,N_16280,N_16014);
nor U16895 (N_16895,N_16448,N_16234);
or U16896 (N_16896,N_16475,N_16231);
nor U16897 (N_16897,N_16019,N_16223);
or U16898 (N_16898,N_16422,N_16153);
nor U16899 (N_16899,N_16116,N_16185);
xor U16900 (N_16900,N_16072,N_16290);
and U16901 (N_16901,N_16020,N_16482);
nor U16902 (N_16902,N_16423,N_16400);
nand U16903 (N_16903,N_16394,N_16153);
and U16904 (N_16904,N_16068,N_16087);
and U16905 (N_16905,N_16385,N_16025);
xnor U16906 (N_16906,N_16229,N_16147);
and U16907 (N_16907,N_16464,N_16083);
and U16908 (N_16908,N_16156,N_16016);
nand U16909 (N_16909,N_16197,N_16043);
and U16910 (N_16910,N_16375,N_16302);
nor U16911 (N_16911,N_16417,N_16110);
nor U16912 (N_16912,N_16038,N_16136);
nor U16913 (N_16913,N_16117,N_16239);
nor U16914 (N_16914,N_16089,N_16429);
nor U16915 (N_16915,N_16013,N_16183);
and U16916 (N_16916,N_16230,N_16031);
and U16917 (N_16917,N_16014,N_16290);
or U16918 (N_16918,N_16188,N_16018);
xor U16919 (N_16919,N_16339,N_16242);
nor U16920 (N_16920,N_16433,N_16401);
and U16921 (N_16921,N_16069,N_16295);
and U16922 (N_16922,N_16028,N_16433);
or U16923 (N_16923,N_16395,N_16254);
and U16924 (N_16924,N_16388,N_16006);
nor U16925 (N_16925,N_16228,N_16076);
nand U16926 (N_16926,N_16199,N_16272);
or U16927 (N_16927,N_16253,N_16175);
or U16928 (N_16928,N_16130,N_16354);
nor U16929 (N_16929,N_16015,N_16127);
nor U16930 (N_16930,N_16410,N_16131);
nor U16931 (N_16931,N_16390,N_16421);
and U16932 (N_16932,N_16317,N_16184);
xnor U16933 (N_16933,N_16293,N_16428);
xor U16934 (N_16934,N_16197,N_16047);
or U16935 (N_16935,N_16011,N_16350);
nor U16936 (N_16936,N_16316,N_16449);
nand U16937 (N_16937,N_16449,N_16175);
nand U16938 (N_16938,N_16430,N_16351);
nand U16939 (N_16939,N_16076,N_16018);
or U16940 (N_16940,N_16018,N_16473);
or U16941 (N_16941,N_16211,N_16413);
nand U16942 (N_16942,N_16329,N_16286);
nand U16943 (N_16943,N_16436,N_16487);
or U16944 (N_16944,N_16156,N_16121);
xnor U16945 (N_16945,N_16370,N_16271);
or U16946 (N_16946,N_16101,N_16432);
or U16947 (N_16947,N_16376,N_16056);
or U16948 (N_16948,N_16067,N_16420);
nand U16949 (N_16949,N_16396,N_16431);
nor U16950 (N_16950,N_16451,N_16182);
nand U16951 (N_16951,N_16453,N_16374);
or U16952 (N_16952,N_16252,N_16165);
nor U16953 (N_16953,N_16036,N_16046);
nand U16954 (N_16954,N_16100,N_16296);
nor U16955 (N_16955,N_16282,N_16260);
nand U16956 (N_16956,N_16470,N_16490);
and U16957 (N_16957,N_16202,N_16168);
nor U16958 (N_16958,N_16439,N_16094);
and U16959 (N_16959,N_16165,N_16472);
or U16960 (N_16960,N_16413,N_16458);
and U16961 (N_16961,N_16377,N_16026);
or U16962 (N_16962,N_16124,N_16231);
and U16963 (N_16963,N_16222,N_16380);
nor U16964 (N_16964,N_16086,N_16451);
or U16965 (N_16965,N_16476,N_16063);
or U16966 (N_16966,N_16233,N_16400);
and U16967 (N_16967,N_16462,N_16220);
or U16968 (N_16968,N_16258,N_16459);
nor U16969 (N_16969,N_16015,N_16410);
or U16970 (N_16970,N_16340,N_16350);
nor U16971 (N_16971,N_16000,N_16011);
nor U16972 (N_16972,N_16021,N_16383);
and U16973 (N_16973,N_16096,N_16314);
or U16974 (N_16974,N_16295,N_16397);
or U16975 (N_16975,N_16264,N_16404);
nor U16976 (N_16976,N_16333,N_16082);
xor U16977 (N_16977,N_16021,N_16440);
or U16978 (N_16978,N_16123,N_16377);
nor U16979 (N_16979,N_16298,N_16403);
and U16980 (N_16980,N_16401,N_16490);
and U16981 (N_16981,N_16477,N_16380);
nand U16982 (N_16982,N_16452,N_16119);
and U16983 (N_16983,N_16438,N_16398);
or U16984 (N_16984,N_16155,N_16388);
nand U16985 (N_16985,N_16016,N_16069);
or U16986 (N_16986,N_16230,N_16274);
nand U16987 (N_16987,N_16447,N_16108);
nand U16988 (N_16988,N_16486,N_16172);
and U16989 (N_16989,N_16421,N_16468);
nand U16990 (N_16990,N_16105,N_16253);
and U16991 (N_16991,N_16113,N_16486);
nor U16992 (N_16992,N_16137,N_16303);
nand U16993 (N_16993,N_16181,N_16150);
or U16994 (N_16994,N_16394,N_16359);
and U16995 (N_16995,N_16478,N_16437);
and U16996 (N_16996,N_16305,N_16342);
nor U16997 (N_16997,N_16040,N_16032);
nor U16998 (N_16998,N_16109,N_16019);
nand U16999 (N_16999,N_16172,N_16457);
nand U17000 (N_17000,N_16641,N_16747);
and U17001 (N_17001,N_16729,N_16913);
or U17002 (N_17002,N_16652,N_16651);
and U17003 (N_17003,N_16914,N_16869);
nor U17004 (N_17004,N_16736,N_16806);
nor U17005 (N_17005,N_16676,N_16529);
nor U17006 (N_17006,N_16885,N_16799);
nand U17007 (N_17007,N_16978,N_16589);
or U17008 (N_17008,N_16707,N_16867);
xor U17009 (N_17009,N_16601,N_16740);
nor U17010 (N_17010,N_16520,N_16685);
nand U17011 (N_17011,N_16540,N_16675);
and U17012 (N_17012,N_16813,N_16743);
or U17013 (N_17013,N_16573,N_16732);
or U17014 (N_17014,N_16980,N_16817);
nand U17015 (N_17015,N_16845,N_16766);
or U17016 (N_17016,N_16622,N_16548);
or U17017 (N_17017,N_16670,N_16852);
or U17018 (N_17018,N_16557,N_16728);
xnor U17019 (N_17019,N_16882,N_16619);
nand U17020 (N_17020,N_16764,N_16769);
or U17021 (N_17021,N_16881,N_16503);
or U17022 (N_17022,N_16804,N_16849);
nand U17023 (N_17023,N_16585,N_16667);
or U17024 (N_17024,N_16955,N_16679);
xnor U17025 (N_17025,N_16860,N_16657);
nor U17026 (N_17026,N_16857,N_16789);
or U17027 (N_17027,N_16604,N_16694);
xor U17028 (N_17028,N_16504,N_16558);
nor U17029 (N_17029,N_16538,N_16579);
nand U17030 (N_17030,N_16810,N_16888);
and U17031 (N_17031,N_16526,N_16886);
or U17032 (N_17032,N_16576,N_16759);
nand U17033 (N_17033,N_16848,N_16894);
nand U17034 (N_17034,N_16976,N_16807);
nand U17035 (N_17035,N_16509,N_16981);
nand U17036 (N_17036,N_16925,N_16872);
and U17037 (N_17037,N_16835,N_16896);
or U17038 (N_17038,N_16906,N_16880);
nand U17039 (N_17039,N_16975,N_16772);
xor U17040 (N_17040,N_16803,N_16866);
or U17041 (N_17041,N_16550,N_16793);
xnor U17042 (N_17042,N_16714,N_16615);
nand U17043 (N_17043,N_16532,N_16546);
or U17044 (N_17044,N_16755,N_16663);
xnor U17045 (N_17045,N_16762,N_16571);
nor U17046 (N_17046,N_16612,N_16570);
or U17047 (N_17047,N_16842,N_16953);
nand U17048 (N_17048,N_16556,N_16752);
nand U17049 (N_17049,N_16705,N_16930);
and U17050 (N_17050,N_16654,N_16517);
and U17051 (N_17051,N_16985,N_16551);
or U17052 (N_17052,N_16902,N_16515);
or U17053 (N_17053,N_16758,N_16844);
nand U17054 (N_17054,N_16878,N_16934);
nor U17055 (N_17055,N_16767,N_16677);
nand U17056 (N_17056,N_16578,N_16837);
nand U17057 (N_17057,N_16632,N_16647);
nand U17058 (N_17058,N_16907,N_16822);
nand U17059 (N_17059,N_16527,N_16513);
xor U17060 (N_17060,N_16846,N_16782);
or U17061 (N_17061,N_16923,N_16610);
and U17062 (N_17062,N_16876,N_16502);
or U17063 (N_17063,N_16709,N_16899);
nand U17064 (N_17064,N_16725,N_16838);
or U17065 (N_17065,N_16761,N_16908);
nand U17066 (N_17066,N_16718,N_16785);
xnor U17067 (N_17067,N_16713,N_16543);
nand U17068 (N_17068,N_16653,N_16959);
and U17069 (N_17069,N_16825,N_16567);
nor U17070 (N_17070,N_16819,N_16693);
nor U17071 (N_17071,N_16832,N_16982);
nand U17072 (N_17072,N_16523,N_16587);
xor U17073 (N_17073,N_16965,N_16892);
and U17074 (N_17074,N_16895,N_16940);
nand U17075 (N_17075,N_16921,N_16927);
and U17076 (N_17076,N_16948,N_16871);
or U17077 (N_17077,N_16995,N_16569);
nand U17078 (N_17078,N_16701,N_16554);
or U17079 (N_17079,N_16583,N_16990);
nor U17080 (N_17080,N_16744,N_16912);
xor U17081 (N_17081,N_16545,N_16672);
nand U17082 (N_17082,N_16501,N_16581);
xor U17083 (N_17083,N_16691,N_16564);
or U17084 (N_17084,N_16771,N_16774);
and U17085 (N_17085,N_16915,N_16661);
nor U17086 (N_17086,N_16624,N_16608);
or U17087 (N_17087,N_16642,N_16794);
nand U17088 (N_17088,N_16814,N_16682);
nand U17089 (N_17089,N_16506,N_16633);
nor U17090 (N_17090,N_16851,N_16778);
nand U17091 (N_17091,N_16737,N_16629);
or U17092 (N_17092,N_16673,N_16577);
and U17093 (N_17093,N_16535,N_16988);
or U17094 (N_17094,N_16531,N_16731);
or U17095 (N_17095,N_16592,N_16855);
nor U17096 (N_17096,N_16820,N_16987);
nor U17097 (N_17097,N_16598,N_16645);
nand U17098 (N_17098,N_16649,N_16974);
and U17099 (N_17099,N_16710,N_16722);
nand U17100 (N_17100,N_16815,N_16984);
nand U17101 (N_17101,N_16524,N_16565);
or U17102 (N_17102,N_16611,N_16922);
or U17103 (N_17103,N_16600,N_16560);
nor U17104 (N_17104,N_16999,N_16519);
and U17105 (N_17105,N_16836,N_16516);
and U17106 (N_17106,N_16937,N_16827);
nand U17107 (N_17107,N_16536,N_16668);
nand U17108 (N_17108,N_16856,N_16893);
nand U17109 (N_17109,N_16919,N_16910);
and U17110 (N_17110,N_16897,N_16765);
nand U17111 (N_17111,N_16648,N_16802);
nand U17112 (N_17112,N_16741,N_16865);
nor U17113 (N_17113,N_16616,N_16784);
nand U17114 (N_17114,N_16760,N_16864);
or U17115 (N_17115,N_16541,N_16639);
nor U17116 (N_17116,N_16542,N_16775);
and U17117 (N_17117,N_16530,N_16644);
or U17118 (N_17118,N_16599,N_16572);
and U17119 (N_17119,N_16681,N_16883);
nor U17120 (N_17120,N_16879,N_16977);
and U17121 (N_17121,N_16783,N_16754);
and U17122 (N_17122,N_16839,N_16808);
nor U17123 (N_17123,N_16544,N_16753);
or U17124 (N_17124,N_16963,N_16858);
nand U17125 (N_17125,N_16702,N_16917);
nand U17126 (N_17126,N_16840,N_16751);
nor U17127 (N_17127,N_16946,N_16818);
and U17128 (N_17128,N_16584,N_16631);
xnor U17129 (N_17129,N_16525,N_16863);
xor U17130 (N_17130,N_16993,N_16952);
or U17131 (N_17131,N_16843,N_16684);
xnor U17132 (N_17132,N_16841,N_16549);
nand U17133 (N_17133,N_16596,N_16662);
and U17134 (N_17134,N_16949,N_16861);
and U17135 (N_17135,N_16877,N_16621);
nor U17136 (N_17136,N_16792,N_16966);
and U17137 (N_17137,N_16547,N_16826);
and U17138 (N_17138,N_16795,N_16958);
nor U17139 (N_17139,N_16593,N_16781);
or U17140 (N_17140,N_16730,N_16575);
or U17141 (N_17141,N_16669,N_16773);
nor U17142 (N_17142,N_16749,N_16680);
and U17143 (N_17143,N_16534,N_16780);
nand U17144 (N_17144,N_16687,N_16521);
or U17145 (N_17145,N_16805,N_16874);
nand U17146 (N_17146,N_16924,N_16791);
nand U17147 (N_17147,N_16986,N_16689);
and U17148 (N_17148,N_16787,N_16715);
nand U17149 (N_17149,N_16996,N_16816);
nor U17150 (N_17150,N_16582,N_16637);
nor U17151 (N_17151,N_16559,N_16994);
and U17152 (N_17152,N_16964,N_16933);
and U17153 (N_17153,N_16742,N_16979);
and U17154 (N_17154,N_16904,N_16875);
and U17155 (N_17155,N_16983,N_16954);
nand U17156 (N_17156,N_16514,N_16683);
nor U17157 (N_17157,N_16779,N_16717);
nor U17158 (N_17158,N_16505,N_16929);
nor U17159 (N_17159,N_16739,N_16539);
nor U17160 (N_17160,N_16692,N_16796);
or U17161 (N_17161,N_16870,N_16727);
or U17162 (N_17162,N_16768,N_16757);
or U17163 (N_17163,N_16628,N_16511);
nor U17164 (N_17164,N_16568,N_16738);
and U17165 (N_17165,N_16947,N_16706);
and U17166 (N_17166,N_16972,N_16969);
and U17167 (N_17167,N_16935,N_16950);
nand U17168 (N_17168,N_16603,N_16697);
nor U17169 (N_17169,N_16678,N_16973);
nand U17170 (N_17170,N_16811,N_16797);
xnor U17171 (N_17171,N_16597,N_16650);
nor U17172 (N_17172,N_16580,N_16723);
or U17173 (N_17173,N_16800,N_16625);
nor U17174 (N_17174,N_16607,N_16655);
and U17175 (N_17175,N_16850,N_16847);
nand U17176 (N_17176,N_16574,N_16735);
nor U17177 (N_17177,N_16620,N_16553);
and U17178 (N_17178,N_16627,N_16821);
or U17179 (N_17179,N_16777,N_16586);
xor U17180 (N_17180,N_16830,N_16696);
nor U17181 (N_17181,N_16756,N_16688);
nor U17182 (N_17182,N_16656,N_16928);
nand U17183 (N_17183,N_16961,N_16720);
xor U17184 (N_17184,N_16905,N_16528);
or U17185 (N_17185,N_16634,N_16831);
or U17186 (N_17186,N_16932,N_16721);
nand U17187 (N_17187,N_16674,N_16618);
nor U17188 (N_17188,N_16828,N_16834);
and U17189 (N_17189,N_16659,N_16970);
xnor U17190 (N_17190,N_16562,N_16500);
xor U17191 (N_17191,N_16991,N_16901);
or U17192 (N_17192,N_16595,N_16941);
and U17193 (N_17193,N_16809,N_16719);
or U17194 (N_17194,N_16533,N_16889);
nor U17195 (N_17195,N_16591,N_16884);
nor U17196 (N_17196,N_16555,N_16887);
nor U17197 (N_17197,N_16960,N_16911);
and U17198 (N_17198,N_16646,N_16695);
nor U17199 (N_17199,N_16638,N_16898);
nand U17200 (N_17200,N_16665,N_16660);
nor U17201 (N_17201,N_16931,N_16862);
and U17202 (N_17202,N_16951,N_16700);
nand U17203 (N_17203,N_16748,N_16643);
nand U17204 (N_17204,N_16939,N_16724);
and U17205 (N_17205,N_16686,N_16823);
nor U17206 (N_17206,N_16943,N_16926);
or U17207 (N_17207,N_16522,N_16900);
nor U17208 (N_17208,N_16868,N_16708);
or U17209 (N_17209,N_16859,N_16630);
and U17210 (N_17210,N_16690,N_16746);
xnor U17211 (N_17211,N_16635,N_16938);
or U17212 (N_17212,N_16873,N_16590);
xnor U17213 (N_17213,N_16698,N_16671);
and U17214 (N_17214,N_16606,N_16962);
and U17215 (N_17215,N_16664,N_16942);
nor U17216 (N_17216,N_16704,N_16989);
or U17217 (N_17217,N_16552,N_16786);
or U17218 (N_17218,N_16512,N_16801);
nor U17219 (N_17219,N_16602,N_16916);
nor U17220 (N_17220,N_16853,N_16566);
nand U17221 (N_17221,N_16537,N_16829);
and U17222 (N_17222,N_16518,N_16640);
nor U17223 (N_17223,N_16790,N_16711);
or U17224 (N_17224,N_16609,N_16666);
or U17225 (N_17225,N_16507,N_16594);
and U17226 (N_17226,N_16613,N_16992);
nand U17227 (N_17227,N_16776,N_16957);
and U17228 (N_17228,N_16998,N_16712);
nor U17229 (N_17229,N_16890,N_16944);
and U17230 (N_17230,N_16703,N_16903);
and U17231 (N_17231,N_16561,N_16920);
or U17232 (N_17232,N_16968,N_16909);
nand U17233 (N_17233,N_16891,N_16588);
or U17234 (N_17234,N_16563,N_16636);
nor U17235 (N_17235,N_16658,N_16854);
and U17236 (N_17236,N_16626,N_16936);
xor U17237 (N_17237,N_16918,N_16716);
and U17238 (N_17238,N_16623,N_16750);
nor U17239 (N_17239,N_16733,N_16770);
nand U17240 (N_17240,N_16734,N_16510);
and U17241 (N_17241,N_16833,N_16945);
and U17242 (N_17242,N_16812,N_16967);
xor U17243 (N_17243,N_16997,N_16824);
nor U17244 (N_17244,N_16614,N_16745);
nand U17245 (N_17245,N_16726,N_16956);
nand U17246 (N_17246,N_16605,N_16699);
xor U17247 (N_17247,N_16788,N_16798);
nand U17248 (N_17248,N_16617,N_16508);
and U17249 (N_17249,N_16971,N_16763);
xor U17250 (N_17250,N_16999,N_16761);
and U17251 (N_17251,N_16867,N_16790);
nor U17252 (N_17252,N_16959,N_16678);
and U17253 (N_17253,N_16796,N_16586);
nand U17254 (N_17254,N_16840,N_16521);
nor U17255 (N_17255,N_16968,N_16754);
or U17256 (N_17256,N_16838,N_16982);
and U17257 (N_17257,N_16528,N_16978);
xnor U17258 (N_17258,N_16659,N_16908);
and U17259 (N_17259,N_16539,N_16961);
and U17260 (N_17260,N_16755,N_16706);
and U17261 (N_17261,N_16836,N_16925);
nor U17262 (N_17262,N_16627,N_16646);
or U17263 (N_17263,N_16752,N_16522);
nand U17264 (N_17264,N_16550,N_16705);
nor U17265 (N_17265,N_16852,N_16969);
or U17266 (N_17266,N_16820,N_16723);
nand U17267 (N_17267,N_16557,N_16920);
nor U17268 (N_17268,N_16928,N_16750);
and U17269 (N_17269,N_16685,N_16548);
nand U17270 (N_17270,N_16871,N_16745);
and U17271 (N_17271,N_16768,N_16554);
and U17272 (N_17272,N_16641,N_16918);
and U17273 (N_17273,N_16528,N_16586);
or U17274 (N_17274,N_16696,N_16930);
nand U17275 (N_17275,N_16994,N_16515);
or U17276 (N_17276,N_16531,N_16793);
or U17277 (N_17277,N_16681,N_16912);
xor U17278 (N_17278,N_16505,N_16517);
nand U17279 (N_17279,N_16828,N_16522);
nor U17280 (N_17280,N_16897,N_16528);
and U17281 (N_17281,N_16598,N_16788);
nand U17282 (N_17282,N_16662,N_16840);
or U17283 (N_17283,N_16597,N_16856);
nand U17284 (N_17284,N_16911,N_16733);
and U17285 (N_17285,N_16898,N_16802);
xnor U17286 (N_17286,N_16780,N_16663);
nor U17287 (N_17287,N_16713,N_16597);
nor U17288 (N_17288,N_16592,N_16668);
nor U17289 (N_17289,N_16594,N_16945);
nor U17290 (N_17290,N_16504,N_16634);
nand U17291 (N_17291,N_16916,N_16659);
nor U17292 (N_17292,N_16905,N_16737);
or U17293 (N_17293,N_16877,N_16893);
nand U17294 (N_17294,N_16896,N_16519);
or U17295 (N_17295,N_16988,N_16503);
and U17296 (N_17296,N_16930,N_16625);
nor U17297 (N_17297,N_16622,N_16807);
or U17298 (N_17298,N_16635,N_16732);
or U17299 (N_17299,N_16821,N_16726);
nand U17300 (N_17300,N_16680,N_16730);
nor U17301 (N_17301,N_16811,N_16846);
nor U17302 (N_17302,N_16568,N_16739);
nor U17303 (N_17303,N_16817,N_16735);
nand U17304 (N_17304,N_16825,N_16585);
and U17305 (N_17305,N_16921,N_16507);
nor U17306 (N_17306,N_16579,N_16806);
or U17307 (N_17307,N_16946,N_16611);
nand U17308 (N_17308,N_16694,N_16899);
nor U17309 (N_17309,N_16746,N_16843);
and U17310 (N_17310,N_16739,N_16903);
and U17311 (N_17311,N_16550,N_16852);
and U17312 (N_17312,N_16802,N_16698);
nand U17313 (N_17313,N_16988,N_16908);
nand U17314 (N_17314,N_16704,N_16927);
xnor U17315 (N_17315,N_16804,N_16986);
nand U17316 (N_17316,N_16920,N_16961);
nand U17317 (N_17317,N_16922,N_16905);
nand U17318 (N_17318,N_16578,N_16827);
nand U17319 (N_17319,N_16787,N_16778);
xor U17320 (N_17320,N_16992,N_16961);
and U17321 (N_17321,N_16725,N_16880);
or U17322 (N_17322,N_16871,N_16914);
or U17323 (N_17323,N_16998,N_16796);
nand U17324 (N_17324,N_16725,N_16580);
nor U17325 (N_17325,N_16726,N_16755);
and U17326 (N_17326,N_16830,N_16883);
and U17327 (N_17327,N_16567,N_16874);
nand U17328 (N_17328,N_16991,N_16720);
nor U17329 (N_17329,N_16615,N_16907);
or U17330 (N_17330,N_16892,N_16796);
or U17331 (N_17331,N_16975,N_16814);
xnor U17332 (N_17332,N_16867,N_16525);
nand U17333 (N_17333,N_16634,N_16848);
or U17334 (N_17334,N_16955,N_16725);
or U17335 (N_17335,N_16980,N_16810);
xor U17336 (N_17336,N_16726,N_16773);
or U17337 (N_17337,N_16630,N_16525);
nor U17338 (N_17338,N_16592,N_16771);
and U17339 (N_17339,N_16916,N_16751);
or U17340 (N_17340,N_16544,N_16679);
or U17341 (N_17341,N_16781,N_16971);
nor U17342 (N_17342,N_16874,N_16750);
nor U17343 (N_17343,N_16618,N_16590);
and U17344 (N_17344,N_16867,N_16866);
nor U17345 (N_17345,N_16558,N_16804);
and U17346 (N_17346,N_16877,N_16534);
and U17347 (N_17347,N_16826,N_16719);
or U17348 (N_17348,N_16970,N_16617);
nand U17349 (N_17349,N_16677,N_16539);
nand U17350 (N_17350,N_16942,N_16886);
nand U17351 (N_17351,N_16982,N_16780);
nand U17352 (N_17352,N_16805,N_16865);
nand U17353 (N_17353,N_16721,N_16883);
or U17354 (N_17354,N_16920,N_16935);
and U17355 (N_17355,N_16694,N_16954);
and U17356 (N_17356,N_16940,N_16735);
and U17357 (N_17357,N_16695,N_16933);
or U17358 (N_17358,N_16696,N_16921);
nor U17359 (N_17359,N_16910,N_16819);
nor U17360 (N_17360,N_16971,N_16709);
and U17361 (N_17361,N_16548,N_16865);
nor U17362 (N_17362,N_16826,N_16592);
or U17363 (N_17363,N_16975,N_16988);
nand U17364 (N_17364,N_16507,N_16653);
nor U17365 (N_17365,N_16648,N_16905);
and U17366 (N_17366,N_16656,N_16950);
nand U17367 (N_17367,N_16521,N_16691);
xor U17368 (N_17368,N_16583,N_16898);
or U17369 (N_17369,N_16535,N_16980);
nand U17370 (N_17370,N_16806,N_16861);
or U17371 (N_17371,N_16625,N_16735);
nand U17372 (N_17372,N_16901,N_16967);
nand U17373 (N_17373,N_16652,N_16992);
nor U17374 (N_17374,N_16562,N_16704);
nand U17375 (N_17375,N_16611,N_16951);
nand U17376 (N_17376,N_16861,N_16777);
nor U17377 (N_17377,N_16717,N_16648);
nand U17378 (N_17378,N_16788,N_16986);
nand U17379 (N_17379,N_16612,N_16645);
and U17380 (N_17380,N_16914,N_16612);
or U17381 (N_17381,N_16991,N_16874);
or U17382 (N_17382,N_16514,N_16816);
or U17383 (N_17383,N_16616,N_16901);
and U17384 (N_17384,N_16713,N_16683);
nor U17385 (N_17385,N_16738,N_16587);
and U17386 (N_17386,N_16939,N_16773);
nand U17387 (N_17387,N_16764,N_16665);
or U17388 (N_17388,N_16792,N_16592);
nor U17389 (N_17389,N_16970,N_16878);
nand U17390 (N_17390,N_16975,N_16632);
nor U17391 (N_17391,N_16697,N_16785);
or U17392 (N_17392,N_16894,N_16869);
xor U17393 (N_17393,N_16695,N_16841);
xor U17394 (N_17394,N_16642,N_16670);
nor U17395 (N_17395,N_16745,N_16653);
nor U17396 (N_17396,N_16923,N_16704);
or U17397 (N_17397,N_16556,N_16954);
or U17398 (N_17398,N_16798,N_16523);
and U17399 (N_17399,N_16707,N_16960);
nand U17400 (N_17400,N_16536,N_16735);
nor U17401 (N_17401,N_16549,N_16672);
or U17402 (N_17402,N_16740,N_16987);
xnor U17403 (N_17403,N_16776,N_16609);
xor U17404 (N_17404,N_16956,N_16546);
and U17405 (N_17405,N_16616,N_16759);
and U17406 (N_17406,N_16919,N_16849);
or U17407 (N_17407,N_16567,N_16634);
and U17408 (N_17408,N_16913,N_16684);
nand U17409 (N_17409,N_16578,N_16989);
nand U17410 (N_17410,N_16519,N_16885);
nor U17411 (N_17411,N_16645,N_16509);
and U17412 (N_17412,N_16784,N_16598);
nor U17413 (N_17413,N_16615,N_16844);
nand U17414 (N_17414,N_16781,N_16908);
or U17415 (N_17415,N_16778,N_16661);
nand U17416 (N_17416,N_16530,N_16795);
xor U17417 (N_17417,N_16626,N_16625);
nand U17418 (N_17418,N_16625,N_16906);
or U17419 (N_17419,N_16912,N_16513);
and U17420 (N_17420,N_16721,N_16739);
nor U17421 (N_17421,N_16955,N_16776);
or U17422 (N_17422,N_16958,N_16735);
nor U17423 (N_17423,N_16924,N_16675);
xnor U17424 (N_17424,N_16534,N_16549);
or U17425 (N_17425,N_16750,N_16800);
and U17426 (N_17426,N_16683,N_16908);
nand U17427 (N_17427,N_16912,N_16621);
nor U17428 (N_17428,N_16724,N_16897);
nor U17429 (N_17429,N_16947,N_16874);
or U17430 (N_17430,N_16586,N_16991);
or U17431 (N_17431,N_16892,N_16766);
nor U17432 (N_17432,N_16901,N_16899);
or U17433 (N_17433,N_16994,N_16966);
xor U17434 (N_17434,N_16741,N_16702);
or U17435 (N_17435,N_16818,N_16618);
and U17436 (N_17436,N_16897,N_16868);
or U17437 (N_17437,N_16697,N_16929);
nor U17438 (N_17438,N_16514,N_16812);
nand U17439 (N_17439,N_16837,N_16555);
or U17440 (N_17440,N_16653,N_16747);
and U17441 (N_17441,N_16546,N_16581);
nand U17442 (N_17442,N_16735,N_16957);
nor U17443 (N_17443,N_16918,N_16802);
xnor U17444 (N_17444,N_16545,N_16807);
nor U17445 (N_17445,N_16781,N_16611);
and U17446 (N_17446,N_16541,N_16649);
nand U17447 (N_17447,N_16935,N_16908);
or U17448 (N_17448,N_16996,N_16719);
nand U17449 (N_17449,N_16584,N_16767);
nor U17450 (N_17450,N_16813,N_16972);
and U17451 (N_17451,N_16810,N_16795);
nand U17452 (N_17452,N_16741,N_16952);
nor U17453 (N_17453,N_16784,N_16506);
nand U17454 (N_17454,N_16981,N_16777);
or U17455 (N_17455,N_16969,N_16668);
nor U17456 (N_17456,N_16898,N_16542);
and U17457 (N_17457,N_16836,N_16743);
nor U17458 (N_17458,N_16870,N_16554);
xor U17459 (N_17459,N_16685,N_16953);
or U17460 (N_17460,N_16942,N_16547);
or U17461 (N_17461,N_16982,N_16718);
nand U17462 (N_17462,N_16523,N_16573);
nor U17463 (N_17463,N_16882,N_16764);
nor U17464 (N_17464,N_16915,N_16829);
nand U17465 (N_17465,N_16733,N_16759);
and U17466 (N_17466,N_16697,N_16849);
or U17467 (N_17467,N_16564,N_16740);
or U17468 (N_17468,N_16514,N_16718);
nand U17469 (N_17469,N_16748,N_16540);
nand U17470 (N_17470,N_16748,N_16950);
and U17471 (N_17471,N_16620,N_16909);
nand U17472 (N_17472,N_16703,N_16989);
or U17473 (N_17473,N_16890,N_16629);
nor U17474 (N_17474,N_16568,N_16653);
and U17475 (N_17475,N_16670,N_16934);
nand U17476 (N_17476,N_16830,N_16900);
and U17477 (N_17477,N_16677,N_16540);
and U17478 (N_17478,N_16985,N_16552);
nand U17479 (N_17479,N_16937,N_16808);
or U17480 (N_17480,N_16531,N_16623);
and U17481 (N_17481,N_16769,N_16743);
and U17482 (N_17482,N_16552,N_16790);
nor U17483 (N_17483,N_16776,N_16651);
nand U17484 (N_17484,N_16940,N_16687);
or U17485 (N_17485,N_16806,N_16998);
or U17486 (N_17486,N_16578,N_16943);
nand U17487 (N_17487,N_16607,N_16702);
nand U17488 (N_17488,N_16572,N_16829);
nor U17489 (N_17489,N_16772,N_16676);
and U17490 (N_17490,N_16728,N_16778);
nor U17491 (N_17491,N_16550,N_16999);
nand U17492 (N_17492,N_16837,N_16740);
or U17493 (N_17493,N_16735,N_16705);
nand U17494 (N_17494,N_16571,N_16703);
or U17495 (N_17495,N_16853,N_16647);
and U17496 (N_17496,N_16619,N_16935);
and U17497 (N_17497,N_16829,N_16860);
nor U17498 (N_17498,N_16961,N_16504);
nand U17499 (N_17499,N_16505,N_16506);
or U17500 (N_17500,N_17355,N_17468);
or U17501 (N_17501,N_17164,N_17002);
nor U17502 (N_17502,N_17000,N_17317);
xor U17503 (N_17503,N_17329,N_17190);
xor U17504 (N_17504,N_17387,N_17263);
nor U17505 (N_17505,N_17496,N_17083);
nor U17506 (N_17506,N_17349,N_17094);
or U17507 (N_17507,N_17093,N_17389);
and U17508 (N_17508,N_17417,N_17401);
and U17509 (N_17509,N_17323,N_17006);
nor U17510 (N_17510,N_17021,N_17269);
nor U17511 (N_17511,N_17178,N_17223);
and U17512 (N_17512,N_17275,N_17110);
nand U17513 (N_17513,N_17290,N_17077);
xnor U17514 (N_17514,N_17037,N_17370);
nand U17515 (N_17515,N_17489,N_17114);
and U17516 (N_17516,N_17425,N_17384);
and U17517 (N_17517,N_17038,N_17013);
and U17518 (N_17518,N_17180,N_17103);
or U17519 (N_17519,N_17377,N_17327);
nand U17520 (N_17520,N_17135,N_17342);
or U17521 (N_17521,N_17189,N_17186);
and U17522 (N_17522,N_17280,N_17367);
or U17523 (N_17523,N_17410,N_17335);
nand U17524 (N_17524,N_17391,N_17369);
and U17525 (N_17525,N_17272,N_17455);
and U17526 (N_17526,N_17497,N_17003);
and U17527 (N_17527,N_17396,N_17406);
nand U17528 (N_17528,N_17218,N_17343);
xnor U17529 (N_17529,N_17357,N_17245);
and U17530 (N_17530,N_17195,N_17145);
and U17531 (N_17531,N_17388,N_17289);
nor U17532 (N_17532,N_17208,N_17404);
nand U17533 (N_17533,N_17113,N_17437);
and U17534 (N_17534,N_17467,N_17112);
nand U17535 (N_17535,N_17028,N_17219);
nor U17536 (N_17536,N_17092,N_17395);
nor U17537 (N_17537,N_17232,N_17148);
xnor U17538 (N_17538,N_17324,N_17490);
nor U17539 (N_17539,N_17044,N_17076);
nor U17540 (N_17540,N_17360,N_17098);
xor U17541 (N_17541,N_17271,N_17282);
and U17542 (N_17542,N_17056,N_17315);
nand U17543 (N_17543,N_17196,N_17022);
and U17544 (N_17544,N_17060,N_17305);
and U17545 (N_17545,N_17328,N_17308);
nand U17546 (N_17546,N_17130,N_17411);
and U17547 (N_17547,N_17236,N_17181);
xor U17548 (N_17548,N_17316,N_17378);
and U17549 (N_17549,N_17095,N_17380);
and U17550 (N_17550,N_17122,N_17207);
nor U17551 (N_17551,N_17458,N_17477);
and U17552 (N_17552,N_17386,N_17184);
nand U17553 (N_17553,N_17452,N_17311);
and U17554 (N_17554,N_17153,N_17019);
nand U17555 (N_17555,N_17158,N_17298);
nor U17556 (N_17556,N_17366,N_17310);
and U17557 (N_17557,N_17071,N_17213);
or U17558 (N_17558,N_17233,N_17020);
or U17559 (N_17559,N_17162,N_17192);
nor U17560 (N_17560,N_17474,N_17206);
or U17561 (N_17561,N_17188,N_17149);
and U17562 (N_17562,N_17499,N_17362);
xor U17563 (N_17563,N_17125,N_17059);
or U17564 (N_17564,N_17050,N_17382);
or U17565 (N_17565,N_17246,N_17185);
and U17566 (N_17566,N_17255,N_17243);
nand U17567 (N_17567,N_17129,N_17226);
or U17568 (N_17568,N_17069,N_17108);
nand U17569 (N_17569,N_17090,N_17228);
nor U17570 (N_17570,N_17211,N_17011);
and U17571 (N_17571,N_17075,N_17447);
nor U17572 (N_17572,N_17177,N_17257);
xor U17573 (N_17573,N_17166,N_17277);
xnor U17574 (N_17574,N_17422,N_17167);
nor U17575 (N_17575,N_17091,N_17444);
nand U17576 (N_17576,N_17152,N_17194);
nand U17577 (N_17577,N_17339,N_17442);
or U17578 (N_17578,N_17459,N_17304);
nor U17579 (N_17579,N_17105,N_17402);
or U17580 (N_17580,N_17332,N_17048);
and U17581 (N_17581,N_17309,N_17081);
nand U17582 (N_17582,N_17372,N_17465);
xor U17583 (N_17583,N_17292,N_17348);
nand U17584 (N_17584,N_17276,N_17222);
or U17585 (N_17585,N_17143,N_17318);
and U17586 (N_17586,N_17104,N_17136);
or U17587 (N_17587,N_17159,N_17487);
nor U17588 (N_17588,N_17408,N_17375);
nor U17589 (N_17589,N_17086,N_17085);
or U17590 (N_17590,N_17405,N_17432);
nor U17591 (N_17591,N_17299,N_17495);
and U17592 (N_17592,N_17448,N_17397);
nor U17593 (N_17593,N_17379,N_17281);
or U17594 (N_17594,N_17144,N_17101);
and U17595 (N_17595,N_17428,N_17027);
nand U17596 (N_17596,N_17287,N_17295);
and U17597 (N_17597,N_17454,N_17041);
or U17598 (N_17598,N_17390,N_17214);
xnor U17599 (N_17599,N_17294,N_17209);
xor U17600 (N_17600,N_17365,N_17183);
or U17601 (N_17601,N_17057,N_17017);
nor U17602 (N_17602,N_17361,N_17446);
xor U17603 (N_17603,N_17313,N_17494);
nand U17604 (N_17604,N_17466,N_17260);
and U17605 (N_17605,N_17285,N_17320);
or U17606 (N_17606,N_17481,N_17248);
or U17607 (N_17607,N_17440,N_17203);
nor U17608 (N_17608,N_17321,N_17398);
nand U17609 (N_17609,N_17385,N_17413);
xnor U17610 (N_17610,N_17025,N_17119);
nor U17611 (N_17611,N_17097,N_17035);
and U17612 (N_17612,N_17023,N_17492);
and U17613 (N_17613,N_17234,N_17146);
nor U17614 (N_17614,N_17126,N_17221);
nand U17615 (N_17615,N_17151,N_17049);
nor U17616 (N_17616,N_17431,N_17066);
nand U17617 (N_17617,N_17393,N_17029);
nand U17618 (N_17618,N_17034,N_17055);
or U17619 (N_17619,N_17224,N_17168);
and U17620 (N_17620,N_17063,N_17358);
nand U17621 (N_17621,N_17302,N_17399);
or U17622 (N_17622,N_17179,N_17150);
xor U17623 (N_17623,N_17051,N_17176);
and U17624 (N_17624,N_17284,N_17251);
nand U17625 (N_17625,N_17383,N_17258);
nor U17626 (N_17626,N_17419,N_17336);
nor U17627 (N_17627,N_17249,N_17058);
and U17628 (N_17628,N_17331,N_17307);
or U17629 (N_17629,N_17430,N_17330);
nand U17630 (N_17630,N_17345,N_17244);
nand U17631 (N_17631,N_17288,N_17068);
or U17632 (N_17632,N_17102,N_17237);
and U17633 (N_17633,N_17198,N_17363);
xnor U17634 (N_17634,N_17427,N_17485);
or U17635 (N_17635,N_17476,N_17306);
or U17636 (N_17636,N_17436,N_17368);
nor U17637 (N_17637,N_17227,N_17400);
or U17638 (N_17638,N_17250,N_17479);
nand U17639 (N_17639,N_17475,N_17464);
and U17640 (N_17640,N_17087,N_17043);
or U17641 (N_17641,N_17191,N_17457);
or U17642 (N_17642,N_17210,N_17010);
xor U17643 (N_17643,N_17341,N_17078);
or U17644 (N_17644,N_17157,N_17215);
nor U17645 (N_17645,N_17337,N_17259);
and U17646 (N_17646,N_17117,N_17033);
nor U17647 (N_17647,N_17353,N_17225);
nand U17648 (N_17648,N_17433,N_17175);
and U17649 (N_17649,N_17418,N_17121);
nand U17650 (N_17650,N_17450,N_17200);
and U17651 (N_17651,N_17074,N_17173);
nor U17652 (N_17652,N_17443,N_17344);
and U17653 (N_17653,N_17351,N_17373);
and U17654 (N_17654,N_17137,N_17202);
xor U17655 (N_17655,N_17160,N_17445);
nand U17656 (N_17656,N_17325,N_17484);
nor U17657 (N_17657,N_17242,N_17291);
and U17658 (N_17658,N_17045,N_17460);
and U17659 (N_17659,N_17434,N_17127);
and U17660 (N_17660,N_17270,N_17334);
nand U17661 (N_17661,N_17201,N_17297);
nand U17662 (N_17662,N_17174,N_17120);
or U17663 (N_17663,N_17491,N_17165);
and U17664 (N_17664,N_17449,N_17403);
nor U17665 (N_17665,N_17073,N_17264);
or U17666 (N_17666,N_17123,N_17187);
or U17667 (N_17667,N_17478,N_17100);
nand U17668 (N_17668,N_17266,N_17156);
and U17669 (N_17669,N_17182,N_17412);
nand U17670 (N_17670,N_17473,N_17435);
and U17671 (N_17671,N_17065,N_17014);
nor U17672 (N_17672,N_17140,N_17079);
nand U17673 (N_17673,N_17261,N_17267);
or U17674 (N_17674,N_17018,N_17001);
or U17675 (N_17675,N_17216,N_17429);
or U17676 (N_17676,N_17482,N_17278);
and U17677 (N_17677,N_17107,N_17199);
nor U17678 (N_17678,N_17109,N_17283);
and U17679 (N_17679,N_17134,N_17352);
or U17680 (N_17680,N_17072,N_17253);
nand U17681 (N_17681,N_17133,N_17009);
and U17682 (N_17682,N_17241,N_17231);
and U17683 (N_17683,N_17338,N_17061);
nor U17684 (N_17684,N_17229,N_17024);
and U17685 (N_17685,N_17423,N_17407);
or U17686 (N_17686,N_17042,N_17131);
xor U17687 (N_17687,N_17220,N_17080);
nand U17688 (N_17688,N_17070,N_17052);
nor U17689 (N_17689,N_17374,N_17314);
nor U17690 (N_17690,N_17286,N_17064);
nand U17691 (N_17691,N_17394,N_17016);
xnor U17692 (N_17692,N_17067,N_17141);
nand U17693 (N_17693,N_17116,N_17279);
and U17694 (N_17694,N_17132,N_17171);
and U17695 (N_17695,N_17138,N_17356);
or U17696 (N_17696,N_17089,N_17273);
nand U17697 (N_17697,N_17256,N_17247);
nor U17698 (N_17698,N_17300,N_17409);
nand U17699 (N_17699,N_17359,N_17193);
or U17700 (N_17700,N_17456,N_17217);
nor U17701 (N_17701,N_17439,N_17462);
or U17702 (N_17702,N_17128,N_17205);
or U17703 (N_17703,N_17030,N_17350);
nand U17704 (N_17704,N_17461,N_17488);
nand U17705 (N_17705,N_17254,N_17470);
xor U17706 (N_17706,N_17155,N_17252);
or U17707 (N_17707,N_17340,N_17169);
and U17708 (N_17708,N_17106,N_17441);
nand U17709 (N_17709,N_17347,N_17262);
nand U17710 (N_17710,N_17376,N_17472);
nand U17711 (N_17711,N_17274,N_17139);
and U17712 (N_17712,N_17005,N_17142);
nor U17713 (N_17713,N_17015,N_17036);
nor U17714 (N_17714,N_17235,N_17031);
nand U17715 (N_17715,N_17039,N_17451);
nand U17716 (N_17716,N_17414,N_17115);
or U17717 (N_17717,N_17230,N_17172);
and U17718 (N_17718,N_17212,N_17333);
or U17719 (N_17719,N_17493,N_17040);
or U17720 (N_17720,N_17046,N_17483);
nand U17721 (N_17721,N_17381,N_17326);
xnor U17722 (N_17722,N_17240,N_17498);
nand U17723 (N_17723,N_17032,N_17319);
xor U17724 (N_17724,N_17364,N_17469);
nand U17725 (N_17725,N_17265,N_17424);
and U17726 (N_17726,N_17096,N_17296);
nor U17727 (N_17727,N_17170,N_17197);
or U17728 (N_17728,N_17415,N_17463);
and U17729 (N_17729,N_17421,N_17471);
nor U17730 (N_17730,N_17371,N_17239);
nand U17731 (N_17731,N_17293,N_17007);
nand U17732 (N_17732,N_17438,N_17161);
and U17733 (N_17733,N_17147,N_17392);
or U17734 (N_17734,N_17008,N_17099);
nor U17735 (N_17735,N_17416,N_17301);
xnor U17736 (N_17736,N_17004,N_17420);
and U17737 (N_17737,N_17053,N_17124);
or U17738 (N_17738,N_17426,N_17268);
nor U17739 (N_17739,N_17453,N_17026);
or U17740 (N_17740,N_17154,N_17322);
or U17741 (N_17741,N_17084,N_17054);
and U17742 (N_17742,N_17486,N_17062);
xor U17743 (N_17743,N_17354,N_17204);
xnor U17744 (N_17744,N_17012,N_17238);
or U17745 (N_17745,N_17346,N_17118);
nand U17746 (N_17746,N_17312,N_17088);
nand U17747 (N_17747,N_17111,N_17047);
nand U17748 (N_17748,N_17480,N_17303);
or U17749 (N_17749,N_17163,N_17082);
and U17750 (N_17750,N_17045,N_17185);
xnor U17751 (N_17751,N_17063,N_17243);
nand U17752 (N_17752,N_17063,N_17242);
and U17753 (N_17753,N_17281,N_17400);
xnor U17754 (N_17754,N_17408,N_17383);
nor U17755 (N_17755,N_17349,N_17014);
nand U17756 (N_17756,N_17172,N_17075);
or U17757 (N_17757,N_17085,N_17073);
and U17758 (N_17758,N_17242,N_17031);
or U17759 (N_17759,N_17417,N_17306);
and U17760 (N_17760,N_17095,N_17315);
xor U17761 (N_17761,N_17151,N_17129);
nor U17762 (N_17762,N_17028,N_17237);
nor U17763 (N_17763,N_17128,N_17441);
or U17764 (N_17764,N_17403,N_17434);
or U17765 (N_17765,N_17481,N_17084);
or U17766 (N_17766,N_17365,N_17054);
nor U17767 (N_17767,N_17490,N_17027);
nor U17768 (N_17768,N_17410,N_17482);
nor U17769 (N_17769,N_17215,N_17462);
nor U17770 (N_17770,N_17443,N_17090);
nor U17771 (N_17771,N_17231,N_17494);
or U17772 (N_17772,N_17481,N_17360);
xnor U17773 (N_17773,N_17367,N_17435);
and U17774 (N_17774,N_17094,N_17396);
nor U17775 (N_17775,N_17016,N_17296);
and U17776 (N_17776,N_17290,N_17098);
or U17777 (N_17777,N_17226,N_17390);
nand U17778 (N_17778,N_17265,N_17005);
or U17779 (N_17779,N_17045,N_17436);
nor U17780 (N_17780,N_17111,N_17033);
or U17781 (N_17781,N_17015,N_17139);
and U17782 (N_17782,N_17107,N_17293);
xnor U17783 (N_17783,N_17246,N_17313);
or U17784 (N_17784,N_17192,N_17318);
or U17785 (N_17785,N_17111,N_17002);
nand U17786 (N_17786,N_17047,N_17212);
or U17787 (N_17787,N_17473,N_17436);
and U17788 (N_17788,N_17438,N_17198);
xor U17789 (N_17789,N_17154,N_17180);
xnor U17790 (N_17790,N_17155,N_17053);
or U17791 (N_17791,N_17066,N_17370);
and U17792 (N_17792,N_17428,N_17268);
xnor U17793 (N_17793,N_17428,N_17351);
nand U17794 (N_17794,N_17421,N_17056);
nand U17795 (N_17795,N_17090,N_17262);
and U17796 (N_17796,N_17238,N_17425);
xnor U17797 (N_17797,N_17256,N_17102);
or U17798 (N_17798,N_17303,N_17071);
xnor U17799 (N_17799,N_17062,N_17377);
nand U17800 (N_17800,N_17282,N_17493);
nor U17801 (N_17801,N_17376,N_17124);
and U17802 (N_17802,N_17465,N_17289);
xnor U17803 (N_17803,N_17433,N_17297);
and U17804 (N_17804,N_17002,N_17385);
and U17805 (N_17805,N_17355,N_17480);
nand U17806 (N_17806,N_17134,N_17073);
and U17807 (N_17807,N_17062,N_17378);
and U17808 (N_17808,N_17385,N_17289);
or U17809 (N_17809,N_17426,N_17450);
or U17810 (N_17810,N_17151,N_17053);
xnor U17811 (N_17811,N_17159,N_17205);
and U17812 (N_17812,N_17210,N_17217);
nor U17813 (N_17813,N_17195,N_17363);
and U17814 (N_17814,N_17032,N_17475);
nor U17815 (N_17815,N_17302,N_17211);
and U17816 (N_17816,N_17410,N_17382);
or U17817 (N_17817,N_17375,N_17379);
nand U17818 (N_17818,N_17274,N_17071);
nor U17819 (N_17819,N_17112,N_17043);
or U17820 (N_17820,N_17459,N_17449);
or U17821 (N_17821,N_17314,N_17173);
nand U17822 (N_17822,N_17268,N_17228);
or U17823 (N_17823,N_17476,N_17070);
and U17824 (N_17824,N_17175,N_17248);
nand U17825 (N_17825,N_17111,N_17051);
nand U17826 (N_17826,N_17414,N_17095);
or U17827 (N_17827,N_17378,N_17073);
or U17828 (N_17828,N_17094,N_17315);
nand U17829 (N_17829,N_17101,N_17381);
nor U17830 (N_17830,N_17368,N_17090);
and U17831 (N_17831,N_17155,N_17113);
or U17832 (N_17832,N_17144,N_17054);
and U17833 (N_17833,N_17135,N_17358);
or U17834 (N_17834,N_17090,N_17175);
or U17835 (N_17835,N_17332,N_17319);
or U17836 (N_17836,N_17108,N_17287);
nand U17837 (N_17837,N_17154,N_17371);
xnor U17838 (N_17838,N_17164,N_17261);
nand U17839 (N_17839,N_17278,N_17293);
nor U17840 (N_17840,N_17207,N_17024);
or U17841 (N_17841,N_17456,N_17417);
nor U17842 (N_17842,N_17130,N_17033);
or U17843 (N_17843,N_17409,N_17411);
nor U17844 (N_17844,N_17250,N_17096);
nor U17845 (N_17845,N_17134,N_17259);
xnor U17846 (N_17846,N_17446,N_17173);
nor U17847 (N_17847,N_17174,N_17204);
or U17848 (N_17848,N_17357,N_17451);
nand U17849 (N_17849,N_17092,N_17322);
xnor U17850 (N_17850,N_17113,N_17084);
or U17851 (N_17851,N_17236,N_17322);
or U17852 (N_17852,N_17366,N_17316);
nand U17853 (N_17853,N_17280,N_17044);
nand U17854 (N_17854,N_17356,N_17477);
nand U17855 (N_17855,N_17128,N_17243);
nand U17856 (N_17856,N_17045,N_17479);
xor U17857 (N_17857,N_17017,N_17487);
nand U17858 (N_17858,N_17259,N_17145);
nor U17859 (N_17859,N_17114,N_17460);
and U17860 (N_17860,N_17385,N_17483);
and U17861 (N_17861,N_17291,N_17117);
nand U17862 (N_17862,N_17086,N_17325);
or U17863 (N_17863,N_17224,N_17146);
and U17864 (N_17864,N_17278,N_17245);
nor U17865 (N_17865,N_17475,N_17306);
or U17866 (N_17866,N_17179,N_17227);
nor U17867 (N_17867,N_17444,N_17246);
nor U17868 (N_17868,N_17041,N_17468);
or U17869 (N_17869,N_17033,N_17171);
nand U17870 (N_17870,N_17007,N_17404);
nand U17871 (N_17871,N_17051,N_17182);
nand U17872 (N_17872,N_17322,N_17226);
nor U17873 (N_17873,N_17469,N_17026);
nor U17874 (N_17874,N_17178,N_17314);
nor U17875 (N_17875,N_17341,N_17024);
xor U17876 (N_17876,N_17263,N_17310);
and U17877 (N_17877,N_17483,N_17067);
nand U17878 (N_17878,N_17224,N_17454);
and U17879 (N_17879,N_17059,N_17083);
xnor U17880 (N_17880,N_17113,N_17349);
or U17881 (N_17881,N_17272,N_17436);
or U17882 (N_17882,N_17471,N_17466);
nand U17883 (N_17883,N_17429,N_17004);
xnor U17884 (N_17884,N_17318,N_17200);
nand U17885 (N_17885,N_17214,N_17020);
or U17886 (N_17886,N_17270,N_17324);
and U17887 (N_17887,N_17470,N_17033);
or U17888 (N_17888,N_17139,N_17490);
xnor U17889 (N_17889,N_17196,N_17093);
xnor U17890 (N_17890,N_17441,N_17216);
nor U17891 (N_17891,N_17386,N_17160);
and U17892 (N_17892,N_17261,N_17302);
or U17893 (N_17893,N_17409,N_17199);
or U17894 (N_17894,N_17337,N_17414);
or U17895 (N_17895,N_17223,N_17233);
and U17896 (N_17896,N_17282,N_17170);
and U17897 (N_17897,N_17012,N_17213);
nor U17898 (N_17898,N_17318,N_17013);
and U17899 (N_17899,N_17277,N_17310);
or U17900 (N_17900,N_17134,N_17150);
and U17901 (N_17901,N_17430,N_17426);
and U17902 (N_17902,N_17007,N_17433);
nor U17903 (N_17903,N_17339,N_17114);
xnor U17904 (N_17904,N_17105,N_17179);
and U17905 (N_17905,N_17379,N_17454);
nor U17906 (N_17906,N_17261,N_17212);
or U17907 (N_17907,N_17463,N_17408);
or U17908 (N_17908,N_17054,N_17469);
nor U17909 (N_17909,N_17202,N_17345);
nor U17910 (N_17910,N_17454,N_17377);
or U17911 (N_17911,N_17006,N_17356);
nand U17912 (N_17912,N_17319,N_17091);
nor U17913 (N_17913,N_17462,N_17316);
xnor U17914 (N_17914,N_17108,N_17420);
nand U17915 (N_17915,N_17222,N_17366);
or U17916 (N_17916,N_17476,N_17048);
nand U17917 (N_17917,N_17430,N_17044);
and U17918 (N_17918,N_17226,N_17015);
nor U17919 (N_17919,N_17148,N_17373);
or U17920 (N_17920,N_17294,N_17337);
and U17921 (N_17921,N_17468,N_17392);
nand U17922 (N_17922,N_17416,N_17066);
and U17923 (N_17923,N_17077,N_17054);
or U17924 (N_17924,N_17375,N_17489);
and U17925 (N_17925,N_17022,N_17432);
or U17926 (N_17926,N_17318,N_17104);
xnor U17927 (N_17927,N_17234,N_17183);
nor U17928 (N_17928,N_17132,N_17490);
nor U17929 (N_17929,N_17073,N_17190);
xor U17930 (N_17930,N_17403,N_17356);
and U17931 (N_17931,N_17387,N_17037);
nand U17932 (N_17932,N_17086,N_17477);
or U17933 (N_17933,N_17319,N_17430);
and U17934 (N_17934,N_17229,N_17404);
or U17935 (N_17935,N_17008,N_17085);
nand U17936 (N_17936,N_17071,N_17210);
and U17937 (N_17937,N_17384,N_17463);
or U17938 (N_17938,N_17308,N_17236);
and U17939 (N_17939,N_17157,N_17112);
nand U17940 (N_17940,N_17490,N_17160);
or U17941 (N_17941,N_17087,N_17096);
nand U17942 (N_17942,N_17283,N_17314);
xnor U17943 (N_17943,N_17223,N_17260);
and U17944 (N_17944,N_17446,N_17377);
and U17945 (N_17945,N_17351,N_17437);
nand U17946 (N_17946,N_17343,N_17419);
nand U17947 (N_17947,N_17322,N_17494);
or U17948 (N_17948,N_17380,N_17376);
or U17949 (N_17949,N_17320,N_17019);
and U17950 (N_17950,N_17054,N_17429);
nor U17951 (N_17951,N_17364,N_17164);
xor U17952 (N_17952,N_17224,N_17104);
and U17953 (N_17953,N_17245,N_17284);
and U17954 (N_17954,N_17238,N_17087);
nand U17955 (N_17955,N_17421,N_17192);
nor U17956 (N_17956,N_17211,N_17116);
nor U17957 (N_17957,N_17061,N_17223);
and U17958 (N_17958,N_17235,N_17014);
and U17959 (N_17959,N_17463,N_17380);
nand U17960 (N_17960,N_17375,N_17074);
nor U17961 (N_17961,N_17041,N_17284);
nor U17962 (N_17962,N_17283,N_17131);
nand U17963 (N_17963,N_17014,N_17451);
nor U17964 (N_17964,N_17027,N_17271);
nor U17965 (N_17965,N_17002,N_17095);
or U17966 (N_17966,N_17450,N_17018);
nor U17967 (N_17967,N_17330,N_17241);
nor U17968 (N_17968,N_17256,N_17164);
or U17969 (N_17969,N_17112,N_17027);
or U17970 (N_17970,N_17381,N_17112);
or U17971 (N_17971,N_17153,N_17284);
nor U17972 (N_17972,N_17341,N_17157);
nor U17973 (N_17973,N_17219,N_17456);
xnor U17974 (N_17974,N_17474,N_17424);
or U17975 (N_17975,N_17461,N_17303);
nand U17976 (N_17976,N_17294,N_17325);
and U17977 (N_17977,N_17268,N_17404);
xor U17978 (N_17978,N_17302,N_17209);
nand U17979 (N_17979,N_17213,N_17133);
nand U17980 (N_17980,N_17455,N_17489);
nand U17981 (N_17981,N_17085,N_17310);
and U17982 (N_17982,N_17394,N_17396);
or U17983 (N_17983,N_17099,N_17376);
and U17984 (N_17984,N_17316,N_17490);
nor U17985 (N_17985,N_17030,N_17135);
xor U17986 (N_17986,N_17398,N_17390);
nand U17987 (N_17987,N_17125,N_17078);
and U17988 (N_17988,N_17355,N_17060);
nor U17989 (N_17989,N_17401,N_17119);
nor U17990 (N_17990,N_17402,N_17325);
and U17991 (N_17991,N_17186,N_17325);
nor U17992 (N_17992,N_17119,N_17402);
or U17993 (N_17993,N_17111,N_17246);
and U17994 (N_17994,N_17009,N_17307);
or U17995 (N_17995,N_17006,N_17340);
or U17996 (N_17996,N_17115,N_17338);
xor U17997 (N_17997,N_17075,N_17010);
nor U17998 (N_17998,N_17113,N_17020);
or U17999 (N_17999,N_17177,N_17382);
nor U18000 (N_18000,N_17630,N_17542);
and U18001 (N_18001,N_17561,N_17699);
and U18002 (N_18002,N_17940,N_17763);
and U18003 (N_18003,N_17778,N_17689);
or U18004 (N_18004,N_17524,N_17633);
nand U18005 (N_18005,N_17797,N_17785);
nor U18006 (N_18006,N_17678,N_17752);
and U18007 (N_18007,N_17596,N_17794);
nand U18008 (N_18008,N_17599,N_17767);
nand U18009 (N_18009,N_17625,N_17818);
nor U18010 (N_18010,N_17620,N_17855);
xor U18011 (N_18011,N_17878,N_17803);
nand U18012 (N_18012,N_17607,N_17842);
and U18013 (N_18013,N_17914,N_17694);
and U18014 (N_18014,N_17541,N_17970);
and U18015 (N_18015,N_17745,N_17864);
nand U18016 (N_18016,N_17800,N_17936);
nand U18017 (N_18017,N_17582,N_17823);
or U18018 (N_18018,N_17576,N_17951);
and U18019 (N_18019,N_17747,N_17784);
and U18020 (N_18020,N_17887,N_17693);
nor U18021 (N_18021,N_17727,N_17890);
and U18022 (N_18022,N_17971,N_17941);
or U18023 (N_18023,N_17590,N_17665);
and U18024 (N_18024,N_17816,N_17865);
or U18025 (N_18025,N_17628,N_17698);
or U18026 (N_18026,N_17577,N_17844);
and U18027 (N_18027,N_17733,N_17682);
nand U18028 (N_18028,N_17930,N_17832);
and U18029 (N_18029,N_17775,N_17597);
nor U18030 (N_18030,N_17875,N_17609);
nor U18031 (N_18031,N_17676,N_17945);
or U18032 (N_18032,N_17760,N_17756);
nor U18033 (N_18033,N_17519,N_17925);
xor U18034 (N_18034,N_17514,N_17673);
nand U18035 (N_18035,N_17933,N_17562);
or U18036 (N_18036,N_17725,N_17983);
or U18037 (N_18037,N_17808,N_17737);
nor U18038 (N_18038,N_17907,N_17539);
nor U18039 (N_18039,N_17993,N_17717);
or U18040 (N_18040,N_17639,N_17703);
nor U18041 (N_18041,N_17932,N_17578);
nand U18042 (N_18042,N_17535,N_17776);
nand U18043 (N_18043,N_17764,N_17623);
and U18044 (N_18044,N_17931,N_17642);
nand U18045 (N_18045,N_17575,N_17943);
nor U18046 (N_18046,N_17584,N_17885);
nand U18047 (N_18047,N_17537,N_17598);
nand U18048 (N_18048,N_17669,N_17972);
or U18049 (N_18049,N_17851,N_17627);
nand U18050 (N_18050,N_17616,N_17985);
nand U18051 (N_18051,N_17761,N_17849);
nand U18052 (N_18052,N_17608,N_17568);
and U18053 (N_18053,N_17977,N_17560);
and U18054 (N_18054,N_17949,N_17805);
or U18055 (N_18055,N_17565,N_17548);
and U18056 (N_18056,N_17831,N_17581);
nor U18057 (N_18057,N_17606,N_17999);
and U18058 (N_18058,N_17790,N_17588);
nor U18059 (N_18059,N_17814,N_17801);
nand U18060 (N_18060,N_17768,N_17615);
nor U18061 (N_18061,N_17750,N_17718);
or U18062 (N_18062,N_17518,N_17600);
nand U18063 (N_18063,N_17532,N_17675);
nand U18064 (N_18064,N_17547,N_17545);
nand U18065 (N_18065,N_17886,N_17526);
nand U18066 (N_18066,N_17692,N_17506);
xor U18067 (N_18067,N_17583,N_17722);
nand U18068 (N_18068,N_17815,N_17829);
nor U18069 (N_18069,N_17724,N_17799);
or U18070 (N_18070,N_17869,N_17589);
nand U18071 (N_18071,N_17706,N_17618);
or U18072 (N_18072,N_17570,N_17557);
and U18073 (N_18073,N_17653,N_17896);
nand U18074 (N_18074,N_17729,N_17742);
nand U18075 (N_18075,N_17942,N_17774);
nand U18076 (N_18076,N_17543,N_17874);
nand U18077 (N_18077,N_17923,N_17915);
and U18078 (N_18078,N_17883,N_17839);
nor U18079 (N_18079,N_17683,N_17748);
nor U18080 (N_18080,N_17664,N_17810);
and U18081 (N_18081,N_17796,N_17788);
or U18082 (N_18082,N_17853,N_17515);
nand U18083 (N_18083,N_17751,N_17573);
or U18084 (N_18084,N_17963,N_17846);
nor U18085 (N_18085,N_17837,N_17968);
or U18086 (N_18086,N_17757,N_17713);
nor U18087 (N_18087,N_17732,N_17904);
or U18088 (N_18088,N_17770,N_17605);
or U18089 (N_18089,N_17859,N_17591);
nor U18090 (N_18090,N_17916,N_17826);
and U18091 (N_18091,N_17868,N_17522);
nor U18092 (N_18092,N_17671,N_17922);
and U18093 (N_18093,N_17986,N_17998);
xor U18094 (N_18094,N_17900,N_17964);
xnor U18095 (N_18095,N_17817,N_17586);
nor U18096 (N_18096,N_17786,N_17631);
xnor U18097 (N_18097,N_17622,N_17563);
and U18098 (N_18098,N_17705,N_17828);
nand U18099 (N_18099,N_17680,N_17512);
and U18100 (N_18100,N_17708,N_17804);
nor U18101 (N_18101,N_17989,N_17918);
and U18102 (N_18102,N_17947,N_17656);
nor U18103 (N_18103,N_17688,N_17629);
nor U18104 (N_18104,N_17843,N_17735);
nor U18105 (N_18105,N_17852,N_17956);
nand U18106 (N_18106,N_17861,N_17954);
nor U18107 (N_18107,N_17516,N_17707);
nand U18108 (N_18108,N_17594,N_17822);
or U18109 (N_18109,N_17592,N_17530);
or U18110 (N_18110,N_17677,N_17967);
nor U18111 (N_18111,N_17648,N_17566);
nor U18112 (N_18112,N_17952,N_17635);
xor U18113 (N_18113,N_17659,N_17593);
and U18114 (N_18114,N_17509,N_17882);
nand U18115 (N_18115,N_17789,N_17906);
nand U18116 (N_18116,N_17657,N_17525);
nand U18117 (N_18117,N_17613,N_17579);
or U18118 (N_18118,N_17624,N_17755);
nand U18119 (N_18119,N_17603,N_17979);
and U18120 (N_18120,N_17834,N_17838);
or U18121 (N_18121,N_17667,N_17500);
nor U18122 (N_18122,N_17702,N_17980);
and U18123 (N_18123,N_17715,N_17809);
or U18124 (N_18124,N_17517,N_17641);
nor U18125 (N_18125,N_17958,N_17610);
nor U18126 (N_18126,N_17513,N_17637);
nor U18127 (N_18127,N_17503,N_17546);
nor U18128 (N_18128,N_17674,N_17905);
nor U18129 (N_18129,N_17990,N_17807);
nor U18130 (N_18130,N_17777,N_17644);
nor U18131 (N_18131,N_17529,N_17549);
and U18132 (N_18132,N_17580,N_17569);
xnor U18133 (N_18133,N_17813,N_17731);
nand U18134 (N_18134,N_17962,N_17966);
nand U18135 (N_18135,N_17912,N_17505);
and U18136 (N_18136,N_17772,N_17780);
nor U18137 (N_18137,N_17711,N_17556);
and U18138 (N_18138,N_17877,N_17827);
xnor U18139 (N_18139,N_17661,N_17550);
xnor U18140 (N_18140,N_17898,N_17686);
or U18141 (N_18141,N_17889,N_17798);
and U18142 (N_18142,N_17502,N_17646);
nand U18143 (N_18143,N_17658,N_17771);
and U18144 (N_18144,N_17802,N_17723);
nor U18145 (N_18145,N_17670,N_17924);
nor U18146 (N_18146,N_17783,N_17953);
or U18147 (N_18147,N_17830,N_17531);
and U18148 (N_18148,N_17917,N_17508);
and U18149 (N_18149,N_17626,N_17555);
nor U18150 (N_18150,N_17870,N_17929);
nor U18151 (N_18151,N_17871,N_17833);
nor U18152 (N_18152,N_17921,N_17879);
nor U18153 (N_18153,N_17709,N_17679);
nor U18154 (N_18154,N_17617,N_17651);
nor U18155 (N_18155,N_17988,N_17880);
nand U18156 (N_18156,N_17973,N_17965);
nor U18157 (N_18157,N_17587,N_17551);
and U18158 (N_18158,N_17544,N_17632);
xnor U18159 (N_18159,N_17919,N_17901);
nor U18160 (N_18160,N_17719,N_17939);
nor U18161 (N_18161,N_17510,N_17720);
or U18162 (N_18162,N_17994,N_17523);
or U18163 (N_18163,N_17884,N_17946);
xor U18164 (N_18164,N_17765,N_17976);
and U18165 (N_18165,N_17612,N_17812);
or U18166 (N_18166,N_17974,N_17820);
and U18167 (N_18167,N_17893,N_17781);
and U18168 (N_18168,N_17619,N_17978);
or U18169 (N_18169,N_17860,N_17937);
and U18170 (N_18170,N_17660,N_17895);
nor U18171 (N_18171,N_17913,N_17858);
nand U18172 (N_18172,N_17975,N_17716);
and U18173 (N_18173,N_17684,N_17521);
xor U18174 (N_18174,N_17749,N_17981);
or U18175 (N_18175,N_17636,N_17754);
xor U18176 (N_18176,N_17595,N_17773);
nand U18177 (N_18177,N_17740,N_17911);
and U18178 (N_18178,N_17643,N_17554);
and U18179 (N_18179,N_17553,N_17738);
and U18180 (N_18180,N_17856,N_17696);
xor U18181 (N_18181,N_17638,N_17564);
or U18182 (N_18182,N_17504,N_17695);
and U18183 (N_18183,N_17928,N_17903);
and U18184 (N_18184,N_17996,N_17690);
or U18185 (N_18185,N_17841,N_17938);
or U18186 (N_18186,N_17654,N_17961);
and U18187 (N_18187,N_17668,N_17959);
nor U18188 (N_18188,N_17567,N_17663);
or U18189 (N_18189,N_17845,N_17850);
nand U18190 (N_18190,N_17655,N_17908);
and U18191 (N_18191,N_17872,N_17854);
xor U18192 (N_18192,N_17571,N_17552);
or U18193 (N_18193,N_17769,N_17712);
nor U18194 (N_18194,N_17857,N_17528);
or U18195 (N_18195,N_17662,N_17714);
nor U18196 (N_18196,N_17894,N_17739);
nand U18197 (N_18197,N_17782,N_17645);
or U18198 (N_18198,N_17863,N_17982);
nor U18199 (N_18199,N_17558,N_17795);
and U18200 (N_18200,N_17540,N_17811);
and U18201 (N_18201,N_17585,N_17734);
and U18202 (N_18202,N_17710,N_17793);
nor U18203 (N_18203,N_17867,N_17909);
and U18204 (N_18204,N_17559,N_17899);
nand U18205 (N_18205,N_17960,N_17806);
or U18206 (N_18206,N_17650,N_17927);
nor U18207 (N_18207,N_17501,N_17700);
nand U18208 (N_18208,N_17791,N_17787);
xnor U18209 (N_18209,N_17614,N_17825);
nand U18210 (N_18210,N_17892,N_17934);
nor U18211 (N_18211,N_17697,N_17640);
and U18212 (N_18212,N_17995,N_17873);
nor U18213 (N_18213,N_17991,N_17847);
nand U18214 (N_18214,N_17721,N_17984);
nand U18215 (N_18215,N_17753,N_17681);
xor U18216 (N_18216,N_17891,N_17848);
and U18217 (N_18217,N_17520,N_17741);
and U18218 (N_18218,N_17944,N_17881);
and U18219 (N_18219,N_17920,N_17910);
and U18220 (N_18220,N_17746,N_17821);
xnor U18221 (N_18221,N_17792,N_17672);
nand U18222 (N_18222,N_17536,N_17969);
nand U18223 (N_18223,N_17728,N_17779);
and U18224 (N_18224,N_17876,N_17572);
or U18225 (N_18225,N_17666,N_17730);
nand U18226 (N_18226,N_17534,N_17601);
nor U18227 (N_18227,N_17704,N_17840);
nand U18228 (N_18228,N_17935,N_17743);
or U18229 (N_18229,N_17611,N_17897);
nand U18230 (N_18230,N_17527,N_17926);
nor U18231 (N_18231,N_17602,N_17726);
nand U18232 (N_18232,N_17574,N_17762);
or U18233 (N_18233,N_17948,N_17507);
or U18234 (N_18234,N_17836,N_17758);
nand U18235 (N_18235,N_17634,N_17766);
or U18236 (N_18236,N_17862,N_17997);
xnor U18237 (N_18237,N_17888,N_17736);
nor U18238 (N_18238,N_17649,N_17511);
and U18239 (N_18239,N_17957,N_17691);
and U18240 (N_18240,N_17621,N_17955);
and U18241 (N_18241,N_17866,N_17987);
and U18242 (N_18242,N_17744,N_17835);
and U18243 (N_18243,N_17538,N_17819);
nor U18244 (N_18244,N_17902,N_17604);
nand U18245 (N_18245,N_17701,N_17992);
nor U18246 (N_18246,N_17687,N_17950);
and U18247 (N_18247,N_17824,N_17647);
or U18248 (N_18248,N_17685,N_17533);
and U18249 (N_18249,N_17759,N_17652);
nor U18250 (N_18250,N_17793,N_17628);
nand U18251 (N_18251,N_17747,N_17922);
and U18252 (N_18252,N_17975,N_17869);
or U18253 (N_18253,N_17732,N_17508);
nand U18254 (N_18254,N_17659,N_17961);
and U18255 (N_18255,N_17690,N_17788);
and U18256 (N_18256,N_17542,N_17607);
nand U18257 (N_18257,N_17967,N_17669);
and U18258 (N_18258,N_17944,N_17985);
nand U18259 (N_18259,N_17505,N_17713);
or U18260 (N_18260,N_17511,N_17971);
xor U18261 (N_18261,N_17853,N_17898);
nor U18262 (N_18262,N_17900,N_17963);
and U18263 (N_18263,N_17513,N_17886);
nand U18264 (N_18264,N_17664,N_17891);
xor U18265 (N_18265,N_17633,N_17826);
xnor U18266 (N_18266,N_17752,N_17549);
nor U18267 (N_18267,N_17720,N_17520);
and U18268 (N_18268,N_17559,N_17700);
xnor U18269 (N_18269,N_17583,N_17716);
or U18270 (N_18270,N_17883,N_17935);
or U18271 (N_18271,N_17693,N_17698);
and U18272 (N_18272,N_17787,N_17814);
and U18273 (N_18273,N_17893,N_17714);
xor U18274 (N_18274,N_17946,N_17575);
or U18275 (N_18275,N_17687,N_17609);
or U18276 (N_18276,N_17581,N_17709);
nand U18277 (N_18277,N_17842,N_17577);
nor U18278 (N_18278,N_17704,N_17502);
or U18279 (N_18279,N_17824,N_17611);
or U18280 (N_18280,N_17521,N_17755);
nand U18281 (N_18281,N_17778,N_17923);
nand U18282 (N_18282,N_17634,N_17548);
nor U18283 (N_18283,N_17896,N_17992);
or U18284 (N_18284,N_17527,N_17910);
xor U18285 (N_18285,N_17911,N_17890);
or U18286 (N_18286,N_17818,N_17702);
nand U18287 (N_18287,N_17933,N_17691);
nor U18288 (N_18288,N_17972,N_17938);
nand U18289 (N_18289,N_17636,N_17817);
or U18290 (N_18290,N_17503,N_17787);
nor U18291 (N_18291,N_17851,N_17558);
nor U18292 (N_18292,N_17595,N_17788);
and U18293 (N_18293,N_17707,N_17665);
or U18294 (N_18294,N_17928,N_17846);
or U18295 (N_18295,N_17992,N_17724);
xnor U18296 (N_18296,N_17646,N_17863);
or U18297 (N_18297,N_17999,N_17725);
nand U18298 (N_18298,N_17983,N_17793);
nor U18299 (N_18299,N_17911,N_17616);
or U18300 (N_18300,N_17630,N_17736);
nand U18301 (N_18301,N_17531,N_17813);
nand U18302 (N_18302,N_17701,N_17880);
and U18303 (N_18303,N_17719,N_17829);
or U18304 (N_18304,N_17667,N_17542);
nor U18305 (N_18305,N_17992,N_17689);
nand U18306 (N_18306,N_17971,N_17842);
and U18307 (N_18307,N_17507,N_17598);
xor U18308 (N_18308,N_17553,N_17822);
xor U18309 (N_18309,N_17973,N_17528);
nor U18310 (N_18310,N_17845,N_17970);
xnor U18311 (N_18311,N_17873,N_17802);
nor U18312 (N_18312,N_17955,N_17599);
or U18313 (N_18313,N_17567,N_17926);
and U18314 (N_18314,N_17627,N_17903);
nand U18315 (N_18315,N_17961,N_17882);
and U18316 (N_18316,N_17964,N_17750);
nor U18317 (N_18317,N_17541,N_17941);
nand U18318 (N_18318,N_17796,N_17508);
nor U18319 (N_18319,N_17747,N_17862);
xnor U18320 (N_18320,N_17530,N_17695);
and U18321 (N_18321,N_17723,N_17847);
or U18322 (N_18322,N_17740,N_17585);
nor U18323 (N_18323,N_17792,N_17970);
nand U18324 (N_18324,N_17538,N_17756);
or U18325 (N_18325,N_17868,N_17834);
and U18326 (N_18326,N_17599,N_17604);
or U18327 (N_18327,N_17829,N_17565);
or U18328 (N_18328,N_17809,N_17893);
or U18329 (N_18329,N_17708,N_17905);
nand U18330 (N_18330,N_17720,N_17633);
nand U18331 (N_18331,N_17820,N_17796);
nand U18332 (N_18332,N_17817,N_17938);
or U18333 (N_18333,N_17525,N_17970);
nor U18334 (N_18334,N_17510,N_17594);
nand U18335 (N_18335,N_17585,N_17536);
nand U18336 (N_18336,N_17545,N_17937);
or U18337 (N_18337,N_17964,N_17619);
xnor U18338 (N_18338,N_17709,N_17593);
nand U18339 (N_18339,N_17885,N_17803);
and U18340 (N_18340,N_17826,N_17927);
nor U18341 (N_18341,N_17923,N_17699);
nand U18342 (N_18342,N_17809,N_17596);
or U18343 (N_18343,N_17777,N_17920);
and U18344 (N_18344,N_17683,N_17583);
and U18345 (N_18345,N_17608,N_17918);
nand U18346 (N_18346,N_17815,N_17575);
and U18347 (N_18347,N_17853,N_17691);
nor U18348 (N_18348,N_17929,N_17799);
or U18349 (N_18349,N_17733,N_17508);
nand U18350 (N_18350,N_17664,N_17857);
or U18351 (N_18351,N_17638,N_17584);
or U18352 (N_18352,N_17924,N_17940);
and U18353 (N_18353,N_17981,N_17689);
or U18354 (N_18354,N_17619,N_17900);
nor U18355 (N_18355,N_17976,N_17811);
nand U18356 (N_18356,N_17877,N_17647);
nor U18357 (N_18357,N_17914,N_17611);
nand U18358 (N_18358,N_17983,N_17689);
xnor U18359 (N_18359,N_17777,N_17782);
nor U18360 (N_18360,N_17555,N_17918);
and U18361 (N_18361,N_17759,N_17550);
or U18362 (N_18362,N_17766,N_17833);
or U18363 (N_18363,N_17755,N_17805);
nand U18364 (N_18364,N_17543,N_17871);
nor U18365 (N_18365,N_17794,N_17688);
or U18366 (N_18366,N_17600,N_17869);
nor U18367 (N_18367,N_17853,N_17791);
xor U18368 (N_18368,N_17751,N_17716);
nor U18369 (N_18369,N_17616,N_17855);
and U18370 (N_18370,N_17829,N_17546);
nor U18371 (N_18371,N_17946,N_17637);
and U18372 (N_18372,N_17626,N_17639);
and U18373 (N_18373,N_17702,N_17733);
and U18374 (N_18374,N_17843,N_17700);
nand U18375 (N_18375,N_17648,N_17751);
nor U18376 (N_18376,N_17596,N_17820);
nor U18377 (N_18377,N_17717,N_17934);
and U18378 (N_18378,N_17797,N_17727);
nand U18379 (N_18379,N_17849,N_17659);
or U18380 (N_18380,N_17859,N_17501);
or U18381 (N_18381,N_17867,N_17780);
xnor U18382 (N_18382,N_17813,N_17893);
and U18383 (N_18383,N_17950,N_17808);
xnor U18384 (N_18384,N_17745,N_17615);
and U18385 (N_18385,N_17769,N_17654);
nand U18386 (N_18386,N_17913,N_17973);
nor U18387 (N_18387,N_17626,N_17719);
nand U18388 (N_18388,N_17843,N_17904);
nand U18389 (N_18389,N_17548,N_17733);
or U18390 (N_18390,N_17521,N_17938);
and U18391 (N_18391,N_17883,N_17876);
nand U18392 (N_18392,N_17986,N_17784);
or U18393 (N_18393,N_17649,N_17578);
xnor U18394 (N_18394,N_17592,N_17767);
or U18395 (N_18395,N_17939,N_17614);
nand U18396 (N_18396,N_17837,N_17936);
or U18397 (N_18397,N_17598,N_17781);
nand U18398 (N_18398,N_17843,N_17849);
or U18399 (N_18399,N_17533,N_17963);
xor U18400 (N_18400,N_17688,N_17603);
or U18401 (N_18401,N_17896,N_17541);
xnor U18402 (N_18402,N_17591,N_17945);
and U18403 (N_18403,N_17513,N_17917);
or U18404 (N_18404,N_17907,N_17889);
or U18405 (N_18405,N_17660,N_17529);
and U18406 (N_18406,N_17831,N_17878);
nand U18407 (N_18407,N_17937,N_17951);
nor U18408 (N_18408,N_17570,N_17686);
and U18409 (N_18409,N_17607,N_17545);
xor U18410 (N_18410,N_17834,N_17581);
nor U18411 (N_18411,N_17836,N_17680);
or U18412 (N_18412,N_17663,N_17589);
and U18413 (N_18413,N_17923,N_17947);
nand U18414 (N_18414,N_17640,N_17648);
nand U18415 (N_18415,N_17833,N_17981);
nand U18416 (N_18416,N_17813,N_17839);
nor U18417 (N_18417,N_17699,N_17681);
nand U18418 (N_18418,N_17620,N_17899);
and U18419 (N_18419,N_17507,N_17983);
and U18420 (N_18420,N_17814,N_17527);
xor U18421 (N_18421,N_17850,N_17873);
nand U18422 (N_18422,N_17782,N_17662);
nand U18423 (N_18423,N_17763,N_17643);
or U18424 (N_18424,N_17656,N_17887);
xor U18425 (N_18425,N_17818,N_17909);
and U18426 (N_18426,N_17811,N_17745);
nand U18427 (N_18427,N_17978,N_17543);
nor U18428 (N_18428,N_17649,N_17526);
nor U18429 (N_18429,N_17886,N_17728);
and U18430 (N_18430,N_17554,N_17886);
nand U18431 (N_18431,N_17556,N_17622);
nor U18432 (N_18432,N_17809,N_17606);
nand U18433 (N_18433,N_17877,N_17995);
nand U18434 (N_18434,N_17746,N_17726);
nand U18435 (N_18435,N_17899,N_17636);
nand U18436 (N_18436,N_17785,N_17579);
nor U18437 (N_18437,N_17500,N_17781);
nor U18438 (N_18438,N_17901,N_17557);
and U18439 (N_18439,N_17787,N_17911);
and U18440 (N_18440,N_17579,N_17765);
or U18441 (N_18441,N_17613,N_17669);
or U18442 (N_18442,N_17669,N_17727);
and U18443 (N_18443,N_17695,N_17501);
nor U18444 (N_18444,N_17722,N_17619);
nand U18445 (N_18445,N_17983,N_17589);
nor U18446 (N_18446,N_17817,N_17882);
and U18447 (N_18447,N_17666,N_17959);
and U18448 (N_18448,N_17725,N_17515);
or U18449 (N_18449,N_17545,N_17714);
and U18450 (N_18450,N_17870,N_17835);
or U18451 (N_18451,N_17548,N_17667);
or U18452 (N_18452,N_17617,N_17834);
nand U18453 (N_18453,N_17922,N_17899);
nor U18454 (N_18454,N_17885,N_17594);
nand U18455 (N_18455,N_17692,N_17597);
or U18456 (N_18456,N_17787,N_17632);
or U18457 (N_18457,N_17751,N_17891);
or U18458 (N_18458,N_17718,N_17833);
or U18459 (N_18459,N_17914,N_17836);
and U18460 (N_18460,N_17542,N_17881);
nor U18461 (N_18461,N_17966,N_17647);
and U18462 (N_18462,N_17999,N_17843);
and U18463 (N_18463,N_17758,N_17773);
nor U18464 (N_18464,N_17795,N_17690);
or U18465 (N_18465,N_17868,N_17738);
nand U18466 (N_18466,N_17526,N_17756);
nand U18467 (N_18467,N_17572,N_17828);
and U18468 (N_18468,N_17865,N_17946);
or U18469 (N_18469,N_17851,N_17677);
nand U18470 (N_18470,N_17588,N_17674);
nand U18471 (N_18471,N_17562,N_17925);
nand U18472 (N_18472,N_17762,N_17668);
nor U18473 (N_18473,N_17640,N_17907);
or U18474 (N_18474,N_17563,N_17725);
xor U18475 (N_18475,N_17684,N_17528);
and U18476 (N_18476,N_17783,N_17609);
nand U18477 (N_18477,N_17520,N_17748);
xor U18478 (N_18478,N_17903,N_17733);
or U18479 (N_18479,N_17895,N_17746);
or U18480 (N_18480,N_17901,N_17807);
nand U18481 (N_18481,N_17505,N_17783);
nand U18482 (N_18482,N_17688,N_17616);
and U18483 (N_18483,N_17826,N_17751);
nor U18484 (N_18484,N_17994,N_17661);
or U18485 (N_18485,N_17834,N_17976);
nor U18486 (N_18486,N_17756,N_17706);
and U18487 (N_18487,N_17896,N_17551);
and U18488 (N_18488,N_17617,N_17559);
nand U18489 (N_18489,N_17504,N_17696);
xor U18490 (N_18490,N_17552,N_17630);
or U18491 (N_18491,N_17783,N_17596);
and U18492 (N_18492,N_17651,N_17614);
nor U18493 (N_18493,N_17902,N_17802);
and U18494 (N_18494,N_17543,N_17892);
xor U18495 (N_18495,N_17863,N_17503);
and U18496 (N_18496,N_17686,N_17843);
nor U18497 (N_18497,N_17780,N_17686);
nand U18498 (N_18498,N_17888,N_17861);
nand U18499 (N_18499,N_17656,N_17532);
or U18500 (N_18500,N_18106,N_18280);
or U18501 (N_18501,N_18051,N_18085);
xnor U18502 (N_18502,N_18036,N_18407);
and U18503 (N_18503,N_18068,N_18107);
nor U18504 (N_18504,N_18015,N_18398);
or U18505 (N_18505,N_18228,N_18286);
or U18506 (N_18506,N_18098,N_18420);
nor U18507 (N_18507,N_18208,N_18447);
and U18508 (N_18508,N_18457,N_18462);
or U18509 (N_18509,N_18124,N_18460);
nor U18510 (N_18510,N_18092,N_18181);
or U18511 (N_18511,N_18197,N_18472);
nor U18512 (N_18512,N_18191,N_18234);
nand U18513 (N_18513,N_18105,N_18287);
xor U18514 (N_18514,N_18161,N_18395);
and U18515 (N_18515,N_18031,N_18469);
or U18516 (N_18516,N_18296,N_18301);
nand U18517 (N_18517,N_18086,N_18331);
xor U18518 (N_18518,N_18353,N_18461);
and U18519 (N_18519,N_18174,N_18293);
and U18520 (N_18520,N_18361,N_18401);
and U18521 (N_18521,N_18499,N_18064);
nand U18522 (N_18522,N_18422,N_18254);
or U18523 (N_18523,N_18049,N_18219);
nand U18524 (N_18524,N_18414,N_18243);
nor U18525 (N_18525,N_18396,N_18229);
nand U18526 (N_18526,N_18081,N_18003);
and U18527 (N_18527,N_18483,N_18385);
nor U18528 (N_18528,N_18135,N_18404);
or U18529 (N_18529,N_18316,N_18405);
nand U18530 (N_18530,N_18364,N_18334);
nand U18531 (N_18531,N_18156,N_18346);
nand U18532 (N_18532,N_18160,N_18299);
and U18533 (N_18533,N_18194,N_18445);
nand U18534 (N_18534,N_18452,N_18166);
or U18535 (N_18535,N_18162,N_18115);
and U18536 (N_18536,N_18290,N_18476);
nand U18537 (N_18537,N_18063,N_18355);
nand U18538 (N_18538,N_18159,N_18378);
or U18539 (N_18539,N_18410,N_18260);
and U18540 (N_18540,N_18300,N_18180);
nand U18541 (N_18541,N_18455,N_18087);
xor U18542 (N_18542,N_18070,N_18377);
nand U18543 (N_18543,N_18247,N_18204);
nand U18544 (N_18544,N_18200,N_18103);
nand U18545 (N_18545,N_18285,N_18205);
or U18546 (N_18546,N_18266,N_18419);
nor U18547 (N_18547,N_18215,N_18177);
nor U18548 (N_18548,N_18305,N_18348);
or U18549 (N_18549,N_18237,N_18345);
or U18550 (N_18550,N_18139,N_18391);
nor U18551 (N_18551,N_18210,N_18190);
nor U18552 (N_18552,N_18065,N_18328);
and U18553 (N_18553,N_18487,N_18265);
nand U18554 (N_18554,N_18335,N_18492);
nor U18555 (N_18555,N_18477,N_18203);
or U18556 (N_18556,N_18123,N_18044);
or U18557 (N_18557,N_18148,N_18446);
nor U18558 (N_18558,N_18009,N_18226);
nand U18559 (N_18559,N_18479,N_18415);
nand U18560 (N_18560,N_18173,N_18431);
and U18561 (N_18561,N_18357,N_18143);
and U18562 (N_18562,N_18365,N_18111);
and U18563 (N_18563,N_18451,N_18034);
and U18564 (N_18564,N_18302,N_18272);
nor U18565 (N_18565,N_18221,N_18320);
nand U18566 (N_18566,N_18062,N_18186);
nand U18567 (N_18567,N_18425,N_18045);
nand U18568 (N_18568,N_18350,N_18141);
or U18569 (N_18569,N_18110,N_18012);
and U18570 (N_18570,N_18038,N_18011);
xor U18571 (N_18571,N_18198,N_18091);
and U18572 (N_18572,N_18449,N_18052);
and U18573 (N_18573,N_18144,N_18120);
xnor U18574 (N_18574,N_18187,N_18137);
nor U18575 (N_18575,N_18040,N_18430);
or U18576 (N_18576,N_18375,N_18104);
or U18577 (N_18577,N_18374,N_18056);
nand U18578 (N_18578,N_18027,N_18261);
nand U18579 (N_18579,N_18471,N_18060);
nor U18580 (N_18580,N_18257,N_18488);
or U18581 (N_18581,N_18278,N_18019);
and U18582 (N_18582,N_18321,N_18403);
nor U18583 (N_18583,N_18498,N_18312);
or U18584 (N_18584,N_18050,N_18354);
nor U18585 (N_18585,N_18369,N_18292);
nand U18586 (N_18586,N_18069,N_18362);
nor U18587 (N_18587,N_18310,N_18214);
or U18588 (N_18588,N_18084,N_18408);
and U18589 (N_18589,N_18494,N_18146);
nand U18590 (N_18590,N_18154,N_18035);
and U18591 (N_18591,N_18225,N_18182);
and U18592 (N_18592,N_18356,N_18307);
nand U18593 (N_18593,N_18444,N_18039);
nand U18594 (N_18594,N_18133,N_18251);
or U18595 (N_18595,N_18493,N_18380);
or U18596 (N_18596,N_18399,N_18317);
nand U18597 (N_18597,N_18170,N_18347);
nand U18598 (N_18598,N_18400,N_18128);
and U18599 (N_18599,N_18097,N_18206);
nor U18600 (N_18600,N_18417,N_18413);
or U18601 (N_18601,N_18435,N_18211);
and U18602 (N_18602,N_18196,N_18473);
or U18603 (N_18603,N_18264,N_18037);
nand U18604 (N_18604,N_18061,N_18021);
or U18605 (N_18605,N_18439,N_18179);
and U18606 (N_18606,N_18239,N_18308);
xor U18607 (N_18607,N_18478,N_18256);
and U18608 (N_18608,N_18132,N_18392);
and U18609 (N_18609,N_18474,N_18114);
and U18610 (N_18610,N_18495,N_18298);
nand U18611 (N_18611,N_18245,N_18279);
and U18612 (N_18612,N_18025,N_18231);
nor U18613 (N_18613,N_18394,N_18423);
nand U18614 (N_18614,N_18093,N_18406);
or U18615 (N_18615,N_18121,N_18340);
xnor U18616 (N_18616,N_18450,N_18193);
nand U18617 (N_18617,N_18250,N_18327);
or U18618 (N_18618,N_18217,N_18288);
xnor U18619 (N_18619,N_18002,N_18426);
nand U18620 (N_18620,N_18443,N_18442);
or U18621 (N_18621,N_18429,N_18017);
nor U18622 (N_18622,N_18384,N_18131);
xnor U18623 (N_18623,N_18157,N_18284);
and U18624 (N_18624,N_18283,N_18195);
or U18625 (N_18625,N_18155,N_18496);
nor U18626 (N_18626,N_18042,N_18441);
or U18627 (N_18627,N_18253,N_18306);
and U18628 (N_18628,N_18233,N_18319);
or U18629 (N_18629,N_18058,N_18158);
nor U18630 (N_18630,N_18094,N_18222);
or U18631 (N_18631,N_18325,N_18269);
or U18632 (N_18632,N_18171,N_18212);
or U18633 (N_18633,N_18289,N_18220);
nor U18634 (N_18634,N_18014,N_18199);
nand U18635 (N_18635,N_18277,N_18013);
nand U18636 (N_18636,N_18329,N_18188);
and U18637 (N_18637,N_18249,N_18454);
xnor U18638 (N_18638,N_18134,N_18163);
and U18639 (N_18639,N_18373,N_18282);
and U18640 (N_18640,N_18150,N_18466);
or U18641 (N_18641,N_18291,N_18475);
and U18642 (N_18642,N_18480,N_18080);
or U18643 (N_18643,N_18418,N_18008);
xor U18644 (N_18644,N_18227,N_18218);
or U18645 (N_18645,N_18048,N_18057);
nor U18646 (N_18646,N_18138,N_18032);
nand U18647 (N_18647,N_18294,N_18341);
nand U18648 (N_18648,N_18102,N_18448);
nand U18649 (N_18649,N_18453,N_18382);
and U18650 (N_18650,N_18349,N_18026);
or U18651 (N_18651,N_18303,N_18076);
nor U18652 (N_18652,N_18022,N_18368);
xor U18653 (N_18653,N_18485,N_18126);
nor U18654 (N_18654,N_18020,N_18344);
nor U18655 (N_18655,N_18088,N_18213);
nand U18656 (N_18656,N_18267,N_18109);
xor U18657 (N_18657,N_18436,N_18053);
or U18658 (N_18658,N_18041,N_18202);
nand U18659 (N_18659,N_18309,N_18016);
or U18660 (N_18660,N_18140,N_18073);
or U18661 (N_18661,N_18127,N_18216);
nor U18662 (N_18662,N_18333,N_18262);
nor U18663 (N_18663,N_18130,N_18484);
nand U18664 (N_18664,N_18388,N_18372);
or U18665 (N_18665,N_18332,N_18255);
nand U18666 (N_18666,N_18491,N_18336);
nand U18667 (N_18667,N_18297,N_18274);
and U18668 (N_18668,N_18175,N_18075);
nor U18669 (N_18669,N_18029,N_18339);
or U18670 (N_18670,N_18077,N_18238);
nor U18671 (N_18671,N_18270,N_18389);
nand U18672 (N_18672,N_18323,N_18047);
nor U18673 (N_18673,N_18152,N_18273);
nor U18674 (N_18674,N_18071,N_18101);
and U18675 (N_18675,N_18242,N_18232);
nand U18676 (N_18676,N_18263,N_18033);
nor U18677 (N_18677,N_18074,N_18004);
or U18678 (N_18678,N_18402,N_18235);
and U18679 (N_18679,N_18351,N_18185);
nand U18680 (N_18680,N_18326,N_18178);
and U18681 (N_18681,N_18024,N_18007);
or U18682 (N_18682,N_18481,N_18464);
or U18683 (N_18683,N_18470,N_18059);
and U18684 (N_18684,N_18304,N_18352);
nor U18685 (N_18685,N_18151,N_18324);
nand U18686 (N_18686,N_18314,N_18363);
nand U18687 (N_18687,N_18437,N_18376);
nand U18688 (N_18688,N_18412,N_18315);
nor U18689 (N_18689,N_18142,N_18268);
and U18690 (N_18690,N_18099,N_18055);
and U18691 (N_18691,N_18164,N_18456);
or U18692 (N_18692,N_18271,N_18259);
nand U18693 (N_18693,N_18189,N_18209);
nand U18694 (N_18694,N_18275,N_18467);
or U18695 (N_18695,N_18082,N_18046);
nand U18696 (N_18696,N_18201,N_18252);
and U18697 (N_18697,N_18183,N_18379);
or U18698 (N_18698,N_18096,N_18005);
nand U18699 (N_18699,N_18486,N_18463);
nor U18700 (N_18700,N_18424,N_18311);
or U18701 (N_18701,N_18427,N_18145);
and U18702 (N_18702,N_18112,N_18122);
nor U18703 (N_18703,N_18397,N_18458);
nand U18704 (N_18704,N_18066,N_18108);
and U18705 (N_18705,N_18416,N_18165);
nor U18706 (N_18706,N_18482,N_18381);
and U18707 (N_18707,N_18386,N_18433);
and U18708 (N_18708,N_18116,N_18095);
or U18709 (N_18709,N_18390,N_18018);
nor U18710 (N_18710,N_18067,N_18072);
nor U18711 (N_18711,N_18147,N_18125);
and U18712 (N_18712,N_18167,N_18030);
nand U18713 (N_18713,N_18010,N_18338);
nand U18714 (N_18714,N_18434,N_18089);
nor U18715 (N_18715,N_18119,N_18118);
xnor U18716 (N_18716,N_18428,N_18000);
nor U18717 (N_18717,N_18313,N_18244);
or U18718 (N_18718,N_18169,N_18176);
nand U18719 (N_18719,N_18241,N_18117);
nand U18720 (N_18720,N_18172,N_18136);
nand U18721 (N_18721,N_18230,N_18236);
nor U18722 (N_18722,N_18421,N_18100);
xnor U18723 (N_18723,N_18330,N_18366);
and U18724 (N_18724,N_18258,N_18459);
nand U18725 (N_18725,N_18440,N_18192);
nor U18726 (N_18726,N_18465,N_18246);
nor U18727 (N_18727,N_18168,N_18043);
and U18728 (N_18728,N_18432,N_18248);
and U18729 (N_18729,N_18409,N_18090);
nand U18730 (N_18730,N_18276,N_18295);
or U18731 (N_18731,N_18497,N_18113);
and U18732 (N_18732,N_18054,N_18149);
xor U18733 (N_18733,N_18393,N_18411);
nor U18734 (N_18734,N_18490,N_18322);
or U18735 (N_18735,N_18028,N_18359);
or U18736 (N_18736,N_18023,N_18468);
nor U18737 (N_18737,N_18343,N_18078);
nand U18738 (N_18738,N_18489,N_18001);
nand U18739 (N_18739,N_18207,N_18438);
and U18740 (N_18740,N_18383,N_18224);
nand U18741 (N_18741,N_18367,N_18153);
xor U18742 (N_18742,N_18184,N_18371);
and U18743 (N_18743,N_18342,N_18079);
and U18744 (N_18744,N_18370,N_18387);
and U18745 (N_18745,N_18083,N_18337);
or U18746 (N_18746,N_18281,N_18360);
nor U18747 (N_18747,N_18129,N_18318);
or U18748 (N_18748,N_18223,N_18358);
nand U18749 (N_18749,N_18240,N_18006);
nand U18750 (N_18750,N_18067,N_18036);
and U18751 (N_18751,N_18186,N_18159);
or U18752 (N_18752,N_18387,N_18384);
or U18753 (N_18753,N_18077,N_18134);
and U18754 (N_18754,N_18214,N_18057);
or U18755 (N_18755,N_18019,N_18104);
nor U18756 (N_18756,N_18144,N_18414);
nand U18757 (N_18757,N_18135,N_18182);
xnor U18758 (N_18758,N_18060,N_18384);
or U18759 (N_18759,N_18239,N_18095);
nor U18760 (N_18760,N_18399,N_18196);
and U18761 (N_18761,N_18208,N_18055);
or U18762 (N_18762,N_18312,N_18054);
or U18763 (N_18763,N_18080,N_18142);
nor U18764 (N_18764,N_18047,N_18260);
nand U18765 (N_18765,N_18039,N_18414);
nand U18766 (N_18766,N_18431,N_18231);
nor U18767 (N_18767,N_18301,N_18271);
nor U18768 (N_18768,N_18006,N_18202);
xor U18769 (N_18769,N_18066,N_18480);
and U18770 (N_18770,N_18339,N_18286);
or U18771 (N_18771,N_18223,N_18436);
or U18772 (N_18772,N_18394,N_18184);
nand U18773 (N_18773,N_18445,N_18203);
and U18774 (N_18774,N_18277,N_18164);
nor U18775 (N_18775,N_18186,N_18245);
xor U18776 (N_18776,N_18263,N_18382);
nor U18777 (N_18777,N_18360,N_18135);
or U18778 (N_18778,N_18443,N_18358);
nand U18779 (N_18779,N_18472,N_18076);
nor U18780 (N_18780,N_18275,N_18335);
and U18781 (N_18781,N_18237,N_18399);
nor U18782 (N_18782,N_18263,N_18408);
and U18783 (N_18783,N_18099,N_18211);
xor U18784 (N_18784,N_18048,N_18308);
nor U18785 (N_18785,N_18222,N_18161);
or U18786 (N_18786,N_18154,N_18256);
nand U18787 (N_18787,N_18281,N_18384);
xnor U18788 (N_18788,N_18036,N_18192);
nand U18789 (N_18789,N_18419,N_18353);
and U18790 (N_18790,N_18312,N_18153);
or U18791 (N_18791,N_18412,N_18018);
nor U18792 (N_18792,N_18377,N_18367);
nand U18793 (N_18793,N_18354,N_18233);
and U18794 (N_18794,N_18250,N_18047);
or U18795 (N_18795,N_18407,N_18362);
nor U18796 (N_18796,N_18183,N_18279);
and U18797 (N_18797,N_18100,N_18289);
or U18798 (N_18798,N_18184,N_18119);
xor U18799 (N_18799,N_18460,N_18045);
nand U18800 (N_18800,N_18356,N_18447);
nand U18801 (N_18801,N_18432,N_18404);
nor U18802 (N_18802,N_18093,N_18458);
xnor U18803 (N_18803,N_18444,N_18317);
xor U18804 (N_18804,N_18053,N_18358);
nor U18805 (N_18805,N_18272,N_18016);
or U18806 (N_18806,N_18410,N_18025);
nor U18807 (N_18807,N_18135,N_18049);
and U18808 (N_18808,N_18029,N_18365);
nand U18809 (N_18809,N_18219,N_18121);
or U18810 (N_18810,N_18219,N_18157);
and U18811 (N_18811,N_18326,N_18320);
nand U18812 (N_18812,N_18123,N_18105);
xor U18813 (N_18813,N_18432,N_18475);
nand U18814 (N_18814,N_18392,N_18390);
nand U18815 (N_18815,N_18469,N_18202);
and U18816 (N_18816,N_18012,N_18170);
nand U18817 (N_18817,N_18264,N_18306);
or U18818 (N_18818,N_18112,N_18015);
nor U18819 (N_18819,N_18334,N_18215);
or U18820 (N_18820,N_18176,N_18287);
or U18821 (N_18821,N_18232,N_18135);
nor U18822 (N_18822,N_18161,N_18116);
and U18823 (N_18823,N_18301,N_18447);
or U18824 (N_18824,N_18381,N_18120);
and U18825 (N_18825,N_18094,N_18400);
and U18826 (N_18826,N_18175,N_18115);
xnor U18827 (N_18827,N_18219,N_18224);
xnor U18828 (N_18828,N_18353,N_18393);
nand U18829 (N_18829,N_18389,N_18469);
or U18830 (N_18830,N_18346,N_18123);
and U18831 (N_18831,N_18269,N_18069);
or U18832 (N_18832,N_18224,N_18391);
or U18833 (N_18833,N_18066,N_18331);
and U18834 (N_18834,N_18449,N_18092);
nor U18835 (N_18835,N_18239,N_18154);
nand U18836 (N_18836,N_18022,N_18066);
and U18837 (N_18837,N_18296,N_18192);
or U18838 (N_18838,N_18125,N_18259);
nand U18839 (N_18839,N_18048,N_18389);
and U18840 (N_18840,N_18476,N_18280);
and U18841 (N_18841,N_18005,N_18028);
and U18842 (N_18842,N_18091,N_18497);
and U18843 (N_18843,N_18333,N_18249);
or U18844 (N_18844,N_18338,N_18167);
nor U18845 (N_18845,N_18363,N_18077);
nand U18846 (N_18846,N_18427,N_18332);
or U18847 (N_18847,N_18223,N_18435);
nor U18848 (N_18848,N_18022,N_18462);
and U18849 (N_18849,N_18348,N_18163);
nand U18850 (N_18850,N_18159,N_18102);
and U18851 (N_18851,N_18156,N_18182);
nand U18852 (N_18852,N_18371,N_18003);
nor U18853 (N_18853,N_18304,N_18466);
and U18854 (N_18854,N_18339,N_18096);
nand U18855 (N_18855,N_18059,N_18066);
or U18856 (N_18856,N_18233,N_18121);
and U18857 (N_18857,N_18497,N_18174);
or U18858 (N_18858,N_18143,N_18195);
and U18859 (N_18859,N_18106,N_18165);
xnor U18860 (N_18860,N_18192,N_18188);
nor U18861 (N_18861,N_18369,N_18160);
nor U18862 (N_18862,N_18299,N_18338);
xnor U18863 (N_18863,N_18374,N_18188);
or U18864 (N_18864,N_18435,N_18279);
xnor U18865 (N_18865,N_18150,N_18065);
or U18866 (N_18866,N_18097,N_18431);
or U18867 (N_18867,N_18201,N_18473);
nor U18868 (N_18868,N_18207,N_18226);
nand U18869 (N_18869,N_18322,N_18070);
nand U18870 (N_18870,N_18273,N_18463);
and U18871 (N_18871,N_18153,N_18026);
and U18872 (N_18872,N_18168,N_18217);
xor U18873 (N_18873,N_18111,N_18133);
and U18874 (N_18874,N_18241,N_18255);
nor U18875 (N_18875,N_18406,N_18361);
nor U18876 (N_18876,N_18265,N_18439);
or U18877 (N_18877,N_18476,N_18150);
or U18878 (N_18878,N_18142,N_18459);
nor U18879 (N_18879,N_18304,N_18170);
and U18880 (N_18880,N_18317,N_18154);
nor U18881 (N_18881,N_18098,N_18286);
or U18882 (N_18882,N_18274,N_18082);
xnor U18883 (N_18883,N_18073,N_18112);
and U18884 (N_18884,N_18413,N_18374);
nand U18885 (N_18885,N_18462,N_18363);
or U18886 (N_18886,N_18348,N_18177);
and U18887 (N_18887,N_18141,N_18070);
and U18888 (N_18888,N_18454,N_18439);
or U18889 (N_18889,N_18485,N_18323);
xor U18890 (N_18890,N_18130,N_18023);
nand U18891 (N_18891,N_18164,N_18022);
or U18892 (N_18892,N_18100,N_18397);
and U18893 (N_18893,N_18483,N_18274);
nand U18894 (N_18894,N_18354,N_18049);
xnor U18895 (N_18895,N_18212,N_18024);
nor U18896 (N_18896,N_18039,N_18435);
xor U18897 (N_18897,N_18358,N_18252);
nand U18898 (N_18898,N_18025,N_18238);
or U18899 (N_18899,N_18135,N_18274);
xnor U18900 (N_18900,N_18224,N_18435);
and U18901 (N_18901,N_18145,N_18017);
and U18902 (N_18902,N_18197,N_18376);
xnor U18903 (N_18903,N_18272,N_18248);
nor U18904 (N_18904,N_18230,N_18294);
and U18905 (N_18905,N_18414,N_18140);
or U18906 (N_18906,N_18265,N_18212);
or U18907 (N_18907,N_18347,N_18371);
nor U18908 (N_18908,N_18173,N_18352);
nand U18909 (N_18909,N_18127,N_18211);
nand U18910 (N_18910,N_18454,N_18181);
and U18911 (N_18911,N_18131,N_18071);
or U18912 (N_18912,N_18168,N_18017);
or U18913 (N_18913,N_18394,N_18387);
xnor U18914 (N_18914,N_18435,N_18475);
xnor U18915 (N_18915,N_18018,N_18436);
nor U18916 (N_18916,N_18115,N_18101);
and U18917 (N_18917,N_18394,N_18266);
and U18918 (N_18918,N_18444,N_18398);
and U18919 (N_18919,N_18170,N_18333);
or U18920 (N_18920,N_18221,N_18402);
nand U18921 (N_18921,N_18485,N_18208);
or U18922 (N_18922,N_18417,N_18045);
xor U18923 (N_18923,N_18072,N_18222);
nand U18924 (N_18924,N_18498,N_18399);
nor U18925 (N_18925,N_18160,N_18046);
or U18926 (N_18926,N_18402,N_18296);
or U18927 (N_18927,N_18487,N_18010);
nor U18928 (N_18928,N_18428,N_18037);
xor U18929 (N_18929,N_18258,N_18322);
and U18930 (N_18930,N_18268,N_18184);
nand U18931 (N_18931,N_18400,N_18146);
nor U18932 (N_18932,N_18063,N_18142);
and U18933 (N_18933,N_18370,N_18410);
or U18934 (N_18934,N_18234,N_18140);
or U18935 (N_18935,N_18348,N_18046);
nand U18936 (N_18936,N_18383,N_18283);
nor U18937 (N_18937,N_18019,N_18023);
or U18938 (N_18938,N_18134,N_18432);
nor U18939 (N_18939,N_18275,N_18167);
xnor U18940 (N_18940,N_18136,N_18198);
xnor U18941 (N_18941,N_18400,N_18255);
or U18942 (N_18942,N_18437,N_18432);
nand U18943 (N_18943,N_18249,N_18097);
nor U18944 (N_18944,N_18167,N_18195);
xor U18945 (N_18945,N_18298,N_18238);
or U18946 (N_18946,N_18155,N_18268);
nor U18947 (N_18947,N_18242,N_18336);
nand U18948 (N_18948,N_18448,N_18385);
nand U18949 (N_18949,N_18086,N_18278);
nand U18950 (N_18950,N_18100,N_18162);
or U18951 (N_18951,N_18204,N_18009);
nand U18952 (N_18952,N_18011,N_18353);
nor U18953 (N_18953,N_18123,N_18371);
nand U18954 (N_18954,N_18394,N_18370);
and U18955 (N_18955,N_18326,N_18317);
and U18956 (N_18956,N_18468,N_18079);
and U18957 (N_18957,N_18100,N_18325);
or U18958 (N_18958,N_18204,N_18074);
nor U18959 (N_18959,N_18042,N_18068);
nand U18960 (N_18960,N_18256,N_18443);
and U18961 (N_18961,N_18035,N_18174);
nand U18962 (N_18962,N_18121,N_18085);
xor U18963 (N_18963,N_18485,N_18476);
nor U18964 (N_18964,N_18226,N_18332);
nor U18965 (N_18965,N_18461,N_18233);
xnor U18966 (N_18966,N_18233,N_18215);
nor U18967 (N_18967,N_18321,N_18174);
or U18968 (N_18968,N_18371,N_18429);
nor U18969 (N_18969,N_18226,N_18123);
and U18970 (N_18970,N_18195,N_18374);
nand U18971 (N_18971,N_18317,N_18278);
or U18972 (N_18972,N_18182,N_18425);
and U18973 (N_18973,N_18059,N_18036);
nor U18974 (N_18974,N_18195,N_18420);
xor U18975 (N_18975,N_18103,N_18007);
or U18976 (N_18976,N_18117,N_18212);
nor U18977 (N_18977,N_18383,N_18041);
xor U18978 (N_18978,N_18022,N_18483);
nand U18979 (N_18979,N_18458,N_18384);
xor U18980 (N_18980,N_18327,N_18004);
nor U18981 (N_18981,N_18155,N_18087);
or U18982 (N_18982,N_18331,N_18403);
or U18983 (N_18983,N_18286,N_18488);
or U18984 (N_18984,N_18218,N_18315);
nor U18985 (N_18985,N_18136,N_18385);
and U18986 (N_18986,N_18033,N_18429);
or U18987 (N_18987,N_18345,N_18078);
and U18988 (N_18988,N_18046,N_18404);
and U18989 (N_18989,N_18359,N_18230);
xnor U18990 (N_18990,N_18070,N_18307);
xor U18991 (N_18991,N_18008,N_18484);
xnor U18992 (N_18992,N_18084,N_18175);
and U18993 (N_18993,N_18174,N_18273);
nand U18994 (N_18994,N_18408,N_18129);
or U18995 (N_18995,N_18237,N_18356);
or U18996 (N_18996,N_18413,N_18483);
and U18997 (N_18997,N_18244,N_18038);
or U18998 (N_18998,N_18085,N_18397);
or U18999 (N_18999,N_18338,N_18348);
nor U19000 (N_19000,N_18810,N_18736);
and U19001 (N_19001,N_18958,N_18693);
and U19002 (N_19002,N_18643,N_18556);
xor U19003 (N_19003,N_18915,N_18602);
xnor U19004 (N_19004,N_18960,N_18663);
nand U19005 (N_19005,N_18593,N_18666);
nor U19006 (N_19006,N_18940,N_18947);
nand U19007 (N_19007,N_18750,N_18879);
nand U19008 (N_19008,N_18838,N_18636);
and U19009 (N_19009,N_18873,N_18922);
and U19010 (N_19010,N_18896,N_18665);
nand U19011 (N_19011,N_18789,N_18704);
nor U19012 (N_19012,N_18951,N_18820);
or U19013 (N_19013,N_18728,N_18936);
nor U19014 (N_19014,N_18723,N_18536);
nand U19015 (N_19015,N_18824,N_18858);
nor U19016 (N_19016,N_18897,N_18982);
and U19017 (N_19017,N_18970,N_18521);
or U19018 (N_19018,N_18702,N_18613);
and U19019 (N_19019,N_18829,N_18932);
or U19020 (N_19020,N_18833,N_18575);
nor U19021 (N_19021,N_18560,N_18972);
xnor U19022 (N_19022,N_18884,N_18800);
or U19023 (N_19023,N_18684,N_18524);
nor U19024 (N_19024,N_18755,N_18866);
or U19025 (N_19025,N_18757,N_18679);
nand U19026 (N_19026,N_18577,N_18853);
xor U19027 (N_19027,N_18671,N_18880);
nor U19028 (N_19028,N_18886,N_18738);
nor U19029 (N_19029,N_18737,N_18538);
nand U19030 (N_19030,N_18984,N_18851);
and U19031 (N_19031,N_18875,N_18517);
xnor U19032 (N_19032,N_18823,N_18615);
nand U19033 (N_19033,N_18759,N_18802);
and U19034 (N_19034,N_18742,N_18659);
and U19035 (N_19035,N_18513,N_18504);
nor U19036 (N_19036,N_18770,N_18911);
and U19037 (N_19037,N_18998,N_18986);
nand U19038 (N_19038,N_18701,N_18834);
and U19039 (N_19039,N_18542,N_18821);
nor U19040 (N_19040,N_18928,N_18836);
and U19041 (N_19041,N_18927,N_18943);
xor U19042 (N_19042,N_18610,N_18990);
and U19043 (N_19043,N_18786,N_18959);
and U19044 (N_19044,N_18758,N_18596);
nor U19045 (N_19045,N_18657,N_18890);
nor U19046 (N_19046,N_18744,N_18988);
nor U19047 (N_19047,N_18599,N_18623);
and U19048 (N_19048,N_18780,N_18777);
or U19049 (N_19049,N_18839,N_18871);
nand U19050 (N_19050,N_18712,N_18653);
and U19051 (N_19051,N_18867,N_18969);
nand U19052 (N_19052,N_18992,N_18640);
nor U19053 (N_19053,N_18557,N_18796);
nor U19054 (N_19054,N_18814,N_18539);
xor U19055 (N_19055,N_18963,N_18715);
or U19056 (N_19056,N_18798,N_18501);
or U19057 (N_19057,N_18555,N_18919);
nor U19058 (N_19058,N_18692,N_18957);
and U19059 (N_19059,N_18850,N_18816);
nor U19060 (N_19060,N_18717,N_18606);
nor U19061 (N_19061,N_18601,N_18722);
or U19062 (N_19062,N_18845,N_18545);
nand U19063 (N_19063,N_18648,N_18803);
or U19064 (N_19064,N_18893,N_18888);
nand U19065 (N_19065,N_18627,N_18804);
xor U19066 (N_19066,N_18697,N_18551);
nand U19067 (N_19067,N_18881,N_18587);
and U19068 (N_19068,N_18872,N_18929);
nor U19069 (N_19069,N_18509,N_18918);
xnor U19070 (N_19070,N_18864,N_18968);
xor U19071 (N_19071,N_18526,N_18774);
or U19072 (N_19072,N_18832,N_18731);
or U19073 (N_19073,N_18638,N_18892);
and U19074 (N_19074,N_18726,N_18903);
nand U19075 (N_19075,N_18690,N_18865);
and U19076 (N_19076,N_18905,N_18748);
xnor U19077 (N_19077,N_18732,N_18908);
nand U19078 (N_19078,N_18724,N_18632);
or U19079 (N_19079,N_18568,N_18978);
and U19080 (N_19080,N_18764,N_18512);
nor U19081 (N_19081,N_18916,N_18554);
and U19082 (N_19082,N_18569,N_18700);
nand U19083 (N_19083,N_18926,N_18869);
and U19084 (N_19084,N_18544,N_18614);
nor U19085 (N_19085,N_18719,N_18725);
or U19086 (N_19086,N_18582,N_18914);
or U19087 (N_19087,N_18518,N_18909);
nor U19088 (N_19088,N_18565,N_18868);
nor U19089 (N_19089,N_18625,N_18583);
nand U19090 (N_19090,N_18797,N_18733);
nand U19091 (N_19091,N_18809,N_18920);
and U19092 (N_19092,N_18787,N_18841);
nand U19093 (N_19093,N_18706,N_18654);
and U19094 (N_19094,N_18688,N_18508);
nor U19095 (N_19095,N_18637,N_18877);
and U19096 (N_19096,N_18756,N_18953);
xor U19097 (N_19097,N_18598,N_18678);
and U19098 (N_19098,N_18674,N_18727);
or U19099 (N_19099,N_18751,N_18891);
or U19100 (N_19100,N_18549,N_18535);
or U19101 (N_19101,N_18580,N_18664);
nand U19102 (N_19102,N_18946,N_18793);
or U19103 (N_19103,N_18779,N_18511);
nand U19104 (N_19104,N_18973,N_18955);
and U19105 (N_19105,N_18937,N_18686);
xor U19106 (N_19106,N_18807,N_18989);
or U19107 (N_19107,N_18516,N_18948);
and U19108 (N_19108,N_18740,N_18574);
or U19109 (N_19109,N_18910,N_18933);
nand U19110 (N_19110,N_18673,N_18954);
nor U19111 (N_19111,N_18677,N_18621);
nand U19112 (N_19112,N_18694,N_18618);
nand U19113 (N_19113,N_18894,N_18695);
nand U19114 (N_19114,N_18620,N_18527);
and U19115 (N_19115,N_18778,N_18540);
or U19116 (N_19116,N_18730,N_18856);
nand U19117 (N_19117,N_18572,N_18707);
xor U19118 (N_19118,N_18876,N_18644);
or U19119 (N_19119,N_18548,N_18710);
nand U19120 (N_19120,N_18862,N_18771);
or U19121 (N_19121,N_18626,N_18848);
nand U19122 (N_19122,N_18528,N_18533);
nor U19123 (N_19123,N_18541,N_18588);
and U19124 (N_19124,N_18805,N_18981);
nand U19125 (N_19125,N_18604,N_18600);
nor U19126 (N_19126,N_18961,N_18772);
nand U19127 (N_19127,N_18590,N_18925);
nor U19128 (N_19128,N_18849,N_18641);
and U19129 (N_19129,N_18578,N_18831);
or U19130 (N_19130,N_18660,N_18938);
nor U19131 (N_19131,N_18612,N_18964);
nor U19132 (N_19132,N_18912,N_18752);
nand U19133 (N_19133,N_18622,N_18515);
nand U19134 (N_19134,N_18519,N_18965);
or U19135 (N_19135,N_18505,N_18785);
xor U19136 (N_19136,N_18899,N_18506);
nand U19137 (N_19137,N_18983,N_18675);
nor U19138 (N_19138,N_18815,N_18633);
or U19139 (N_19139,N_18776,N_18768);
and U19140 (N_19140,N_18503,N_18882);
nand U19141 (N_19141,N_18931,N_18979);
and U19142 (N_19142,N_18507,N_18564);
nand U19143 (N_19143,N_18628,N_18962);
nand U19144 (N_19144,N_18558,N_18617);
nor U19145 (N_19145,N_18543,N_18788);
xor U19146 (N_19146,N_18883,N_18826);
nand U19147 (N_19147,N_18840,N_18502);
nand U19148 (N_19148,N_18563,N_18591);
nor U19149 (N_19149,N_18642,N_18993);
or U19150 (N_19150,N_18949,N_18714);
xor U19151 (N_19151,N_18523,N_18561);
nand U19152 (N_19152,N_18645,N_18586);
nand U19153 (N_19153,N_18682,N_18913);
and U19154 (N_19154,N_18611,N_18837);
xor U19155 (N_19155,N_18629,N_18799);
and U19156 (N_19156,N_18552,N_18830);
and U19157 (N_19157,N_18656,N_18670);
and U19158 (N_19158,N_18795,N_18874);
and U19159 (N_19159,N_18531,N_18945);
nor U19160 (N_19160,N_18843,N_18822);
nand U19161 (N_19161,N_18980,N_18828);
and U19162 (N_19162,N_18597,N_18608);
and U19163 (N_19163,N_18801,N_18818);
xnor U19164 (N_19164,N_18902,N_18765);
xnor U19165 (N_19165,N_18781,N_18975);
and U19166 (N_19166,N_18844,N_18650);
or U19167 (N_19167,N_18534,N_18889);
and U19168 (N_19168,N_18579,N_18753);
nor U19169 (N_19169,N_18749,N_18952);
or U19170 (N_19170,N_18746,N_18649);
or U19171 (N_19171,N_18589,N_18835);
nand U19172 (N_19172,N_18861,N_18683);
nor U19173 (N_19173,N_18775,N_18529);
and U19174 (N_19174,N_18584,N_18860);
xnor U19175 (N_19175,N_18716,N_18939);
nand U19176 (N_19176,N_18974,N_18729);
or U19177 (N_19177,N_18901,N_18699);
or U19178 (N_19178,N_18607,N_18635);
and U19179 (N_19179,N_18500,N_18741);
nor U19180 (N_19180,N_18530,N_18991);
or U19181 (N_19181,N_18669,N_18680);
or U19182 (N_19182,N_18720,N_18687);
or U19183 (N_19183,N_18827,N_18647);
xnor U19184 (N_19184,N_18935,N_18944);
or U19185 (N_19185,N_18718,N_18576);
nor U19186 (N_19186,N_18655,N_18760);
or U19187 (N_19187,N_18857,N_18739);
nand U19188 (N_19188,N_18811,N_18782);
or U19189 (N_19189,N_18999,N_18976);
or U19190 (N_19190,N_18514,N_18956);
and U19191 (N_19191,N_18791,N_18870);
nand U19192 (N_19192,N_18941,N_18696);
xor U19193 (N_19193,N_18651,N_18689);
and U19194 (N_19194,N_18977,N_18825);
nor U19195 (N_19195,N_18652,N_18773);
or U19196 (N_19196,N_18658,N_18705);
nand U19197 (N_19197,N_18971,N_18676);
and U19198 (N_19198,N_18573,N_18747);
and U19199 (N_19199,N_18698,N_18546);
nand U19200 (N_19200,N_18924,N_18852);
or U19201 (N_19201,N_18537,N_18808);
or U19202 (N_19202,N_18847,N_18895);
or U19203 (N_19203,N_18609,N_18790);
or U19204 (N_19204,N_18592,N_18603);
nor U19205 (N_19205,N_18906,N_18846);
xor U19206 (N_19206,N_18996,N_18721);
nor U19207 (N_19207,N_18783,N_18594);
and U19208 (N_19208,N_18639,N_18942);
and U19209 (N_19209,N_18930,N_18662);
nand U19210 (N_19210,N_18734,N_18743);
nor U19211 (N_19211,N_18631,N_18685);
and U19212 (N_19212,N_18806,N_18985);
and U19213 (N_19213,N_18709,N_18708);
nor U19214 (N_19214,N_18668,N_18522);
or U19215 (N_19215,N_18761,N_18898);
and U19216 (N_19216,N_18532,N_18547);
xor U19217 (N_19217,N_18624,N_18994);
xnor U19218 (N_19218,N_18819,N_18566);
nor U19219 (N_19219,N_18987,N_18812);
nand U19220 (N_19220,N_18713,N_18763);
xor U19221 (N_19221,N_18967,N_18817);
nor U19222 (N_19222,N_18784,N_18754);
nor U19223 (N_19223,N_18745,N_18691);
nor U19224 (N_19224,N_18966,N_18711);
and U19225 (N_19225,N_18585,N_18735);
nor U19226 (N_19226,N_18842,N_18525);
nand U19227 (N_19227,N_18995,N_18885);
and U19228 (N_19228,N_18510,N_18923);
and U19229 (N_19229,N_18934,N_18646);
nor U19230 (N_19230,N_18766,N_18559);
xnor U19231 (N_19231,N_18917,N_18667);
or U19232 (N_19232,N_18997,N_18854);
nand U19233 (N_19233,N_18855,N_18550);
nand U19234 (N_19234,N_18634,N_18681);
or U19235 (N_19235,N_18570,N_18703);
nor U19236 (N_19236,N_18605,N_18921);
and U19237 (N_19237,N_18630,N_18553);
nand U19238 (N_19238,N_18907,N_18661);
xor U19239 (N_19239,N_18767,N_18762);
or U19240 (N_19240,N_18794,N_18904);
or U19241 (N_19241,N_18567,N_18672);
nor U19242 (N_19242,N_18878,N_18616);
nand U19243 (N_19243,N_18900,N_18520);
and U19244 (N_19244,N_18562,N_18792);
and U19245 (N_19245,N_18619,N_18950);
nor U19246 (N_19246,N_18571,N_18813);
nand U19247 (N_19247,N_18595,N_18581);
nor U19248 (N_19248,N_18863,N_18859);
nand U19249 (N_19249,N_18769,N_18887);
and U19250 (N_19250,N_18746,N_18927);
nor U19251 (N_19251,N_18564,N_18741);
nand U19252 (N_19252,N_18920,N_18932);
nor U19253 (N_19253,N_18889,N_18878);
or U19254 (N_19254,N_18593,N_18580);
or U19255 (N_19255,N_18925,N_18585);
nand U19256 (N_19256,N_18544,N_18840);
or U19257 (N_19257,N_18962,N_18517);
nand U19258 (N_19258,N_18535,N_18854);
xor U19259 (N_19259,N_18524,N_18596);
or U19260 (N_19260,N_18980,N_18954);
nand U19261 (N_19261,N_18721,N_18704);
xor U19262 (N_19262,N_18963,N_18724);
and U19263 (N_19263,N_18967,N_18901);
xor U19264 (N_19264,N_18861,N_18685);
or U19265 (N_19265,N_18899,N_18570);
xnor U19266 (N_19266,N_18596,N_18600);
and U19267 (N_19267,N_18579,N_18622);
and U19268 (N_19268,N_18753,N_18856);
and U19269 (N_19269,N_18828,N_18802);
and U19270 (N_19270,N_18607,N_18976);
or U19271 (N_19271,N_18771,N_18629);
or U19272 (N_19272,N_18774,N_18747);
or U19273 (N_19273,N_18537,N_18953);
nor U19274 (N_19274,N_18714,N_18832);
nor U19275 (N_19275,N_18502,N_18572);
xor U19276 (N_19276,N_18924,N_18627);
xor U19277 (N_19277,N_18553,N_18706);
and U19278 (N_19278,N_18681,N_18705);
or U19279 (N_19279,N_18982,N_18633);
nand U19280 (N_19280,N_18637,N_18662);
nand U19281 (N_19281,N_18748,N_18856);
nand U19282 (N_19282,N_18889,N_18681);
or U19283 (N_19283,N_18760,N_18892);
and U19284 (N_19284,N_18514,N_18966);
or U19285 (N_19285,N_18891,N_18533);
nor U19286 (N_19286,N_18884,N_18943);
and U19287 (N_19287,N_18641,N_18915);
or U19288 (N_19288,N_18711,N_18507);
or U19289 (N_19289,N_18756,N_18619);
nor U19290 (N_19290,N_18758,N_18620);
nand U19291 (N_19291,N_18924,N_18692);
xor U19292 (N_19292,N_18699,N_18847);
nand U19293 (N_19293,N_18909,N_18982);
or U19294 (N_19294,N_18605,N_18580);
and U19295 (N_19295,N_18698,N_18773);
and U19296 (N_19296,N_18621,N_18528);
nand U19297 (N_19297,N_18984,N_18657);
xnor U19298 (N_19298,N_18605,N_18764);
and U19299 (N_19299,N_18511,N_18596);
nor U19300 (N_19300,N_18852,N_18699);
nor U19301 (N_19301,N_18649,N_18905);
or U19302 (N_19302,N_18990,N_18865);
nand U19303 (N_19303,N_18688,N_18727);
xor U19304 (N_19304,N_18846,N_18955);
or U19305 (N_19305,N_18638,N_18535);
and U19306 (N_19306,N_18543,N_18570);
nand U19307 (N_19307,N_18644,N_18955);
or U19308 (N_19308,N_18571,N_18924);
and U19309 (N_19309,N_18911,N_18681);
or U19310 (N_19310,N_18602,N_18895);
xnor U19311 (N_19311,N_18856,N_18614);
and U19312 (N_19312,N_18919,N_18787);
nor U19313 (N_19313,N_18952,N_18719);
nand U19314 (N_19314,N_18875,N_18759);
and U19315 (N_19315,N_18922,N_18764);
or U19316 (N_19316,N_18804,N_18917);
nor U19317 (N_19317,N_18759,N_18747);
nor U19318 (N_19318,N_18640,N_18503);
nor U19319 (N_19319,N_18895,N_18983);
and U19320 (N_19320,N_18747,N_18761);
nand U19321 (N_19321,N_18667,N_18772);
xor U19322 (N_19322,N_18962,N_18777);
and U19323 (N_19323,N_18788,N_18520);
and U19324 (N_19324,N_18957,N_18705);
and U19325 (N_19325,N_18615,N_18641);
nand U19326 (N_19326,N_18608,N_18658);
nand U19327 (N_19327,N_18584,N_18826);
nor U19328 (N_19328,N_18500,N_18929);
xor U19329 (N_19329,N_18781,N_18624);
nand U19330 (N_19330,N_18675,N_18551);
or U19331 (N_19331,N_18966,N_18524);
or U19332 (N_19332,N_18834,N_18757);
or U19333 (N_19333,N_18559,N_18591);
and U19334 (N_19334,N_18812,N_18925);
nor U19335 (N_19335,N_18913,N_18890);
nor U19336 (N_19336,N_18832,N_18975);
nor U19337 (N_19337,N_18983,N_18653);
nor U19338 (N_19338,N_18880,N_18805);
or U19339 (N_19339,N_18726,N_18555);
and U19340 (N_19340,N_18944,N_18706);
nand U19341 (N_19341,N_18936,N_18882);
and U19342 (N_19342,N_18890,N_18846);
xnor U19343 (N_19343,N_18766,N_18647);
and U19344 (N_19344,N_18589,N_18575);
xnor U19345 (N_19345,N_18730,N_18917);
nor U19346 (N_19346,N_18975,N_18995);
or U19347 (N_19347,N_18557,N_18528);
or U19348 (N_19348,N_18590,N_18563);
and U19349 (N_19349,N_18943,N_18982);
and U19350 (N_19350,N_18897,N_18961);
and U19351 (N_19351,N_18619,N_18647);
nor U19352 (N_19352,N_18815,N_18991);
xnor U19353 (N_19353,N_18694,N_18857);
nor U19354 (N_19354,N_18575,N_18738);
or U19355 (N_19355,N_18848,N_18976);
nor U19356 (N_19356,N_18873,N_18538);
nor U19357 (N_19357,N_18550,N_18587);
or U19358 (N_19358,N_18703,N_18721);
xnor U19359 (N_19359,N_18758,N_18788);
nor U19360 (N_19360,N_18771,N_18609);
and U19361 (N_19361,N_18533,N_18554);
or U19362 (N_19362,N_18642,N_18887);
nand U19363 (N_19363,N_18537,N_18757);
nor U19364 (N_19364,N_18905,N_18792);
and U19365 (N_19365,N_18924,N_18847);
nor U19366 (N_19366,N_18942,N_18610);
or U19367 (N_19367,N_18662,N_18847);
nand U19368 (N_19368,N_18575,N_18939);
nor U19369 (N_19369,N_18901,N_18782);
nand U19370 (N_19370,N_18993,N_18980);
nor U19371 (N_19371,N_18813,N_18812);
nand U19372 (N_19372,N_18783,N_18889);
and U19373 (N_19373,N_18781,N_18520);
nor U19374 (N_19374,N_18622,N_18706);
xnor U19375 (N_19375,N_18668,N_18955);
and U19376 (N_19376,N_18877,N_18728);
nand U19377 (N_19377,N_18889,N_18774);
or U19378 (N_19378,N_18611,N_18989);
or U19379 (N_19379,N_18709,N_18596);
nand U19380 (N_19380,N_18731,N_18732);
and U19381 (N_19381,N_18720,N_18797);
or U19382 (N_19382,N_18543,N_18822);
nor U19383 (N_19383,N_18723,N_18521);
and U19384 (N_19384,N_18740,N_18897);
nor U19385 (N_19385,N_18734,N_18695);
nand U19386 (N_19386,N_18972,N_18839);
and U19387 (N_19387,N_18703,N_18893);
nand U19388 (N_19388,N_18980,N_18658);
or U19389 (N_19389,N_18522,N_18693);
and U19390 (N_19390,N_18935,N_18614);
and U19391 (N_19391,N_18526,N_18797);
or U19392 (N_19392,N_18545,N_18503);
nor U19393 (N_19393,N_18895,N_18902);
or U19394 (N_19394,N_18544,N_18611);
or U19395 (N_19395,N_18635,N_18746);
xnor U19396 (N_19396,N_18599,N_18521);
or U19397 (N_19397,N_18948,N_18833);
nor U19398 (N_19398,N_18514,N_18786);
xor U19399 (N_19399,N_18533,N_18928);
and U19400 (N_19400,N_18970,N_18809);
or U19401 (N_19401,N_18627,N_18873);
and U19402 (N_19402,N_18725,N_18643);
nand U19403 (N_19403,N_18626,N_18806);
xnor U19404 (N_19404,N_18869,N_18634);
nand U19405 (N_19405,N_18785,N_18759);
or U19406 (N_19406,N_18772,N_18639);
and U19407 (N_19407,N_18822,N_18718);
nor U19408 (N_19408,N_18763,N_18907);
or U19409 (N_19409,N_18779,N_18682);
or U19410 (N_19410,N_18582,N_18609);
and U19411 (N_19411,N_18542,N_18520);
nor U19412 (N_19412,N_18839,N_18634);
and U19413 (N_19413,N_18923,N_18707);
nor U19414 (N_19414,N_18839,N_18516);
nand U19415 (N_19415,N_18511,N_18595);
nor U19416 (N_19416,N_18974,N_18634);
or U19417 (N_19417,N_18684,N_18575);
and U19418 (N_19418,N_18883,N_18976);
or U19419 (N_19419,N_18952,N_18938);
xnor U19420 (N_19420,N_18961,N_18564);
and U19421 (N_19421,N_18787,N_18648);
xnor U19422 (N_19422,N_18756,N_18890);
nand U19423 (N_19423,N_18586,N_18982);
or U19424 (N_19424,N_18548,N_18927);
and U19425 (N_19425,N_18855,N_18566);
nor U19426 (N_19426,N_18588,N_18564);
nand U19427 (N_19427,N_18588,N_18609);
nand U19428 (N_19428,N_18660,N_18606);
and U19429 (N_19429,N_18960,N_18502);
or U19430 (N_19430,N_18913,N_18997);
nand U19431 (N_19431,N_18694,N_18651);
nand U19432 (N_19432,N_18886,N_18953);
and U19433 (N_19433,N_18728,N_18544);
or U19434 (N_19434,N_18504,N_18992);
nor U19435 (N_19435,N_18897,N_18802);
xnor U19436 (N_19436,N_18773,N_18736);
or U19437 (N_19437,N_18633,N_18967);
nand U19438 (N_19438,N_18949,N_18725);
nand U19439 (N_19439,N_18518,N_18656);
and U19440 (N_19440,N_18900,N_18501);
nor U19441 (N_19441,N_18509,N_18760);
nand U19442 (N_19442,N_18694,N_18751);
or U19443 (N_19443,N_18504,N_18622);
and U19444 (N_19444,N_18823,N_18756);
and U19445 (N_19445,N_18645,N_18807);
or U19446 (N_19446,N_18724,N_18797);
or U19447 (N_19447,N_18879,N_18780);
and U19448 (N_19448,N_18963,N_18955);
and U19449 (N_19449,N_18726,N_18922);
or U19450 (N_19450,N_18672,N_18859);
nor U19451 (N_19451,N_18629,N_18606);
nand U19452 (N_19452,N_18520,N_18898);
xnor U19453 (N_19453,N_18603,N_18604);
or U19454 (N_19454,N_18806,N_18992);
nand U19455 (N_19455,N_18684,N_18696);
nand U19456 (N_19456,N_18524,N_18508);
nor U19457 (N_19457,N_18633,N_18763);
nand U19458 (N_19458,N_18891,N_18738);
nor U19459 (N_19459,N_18536,N_18721);
and U19460 (N_19460,N_18598,N_18854);
and U19461 (N_19461,N_18809,N_18969);
and U19462 (N_19462,N_18636,N_18723);
and U19463 (N_19463,N_18513,N_18588);
nor U19464 (N_19464,N_18513,N_18531);
or U19465 (N_19465,N_18811,N_18715);
and U19466 (N_19466,N_18691,N_18694);
or U19467 (N_19467,N_18842,N_18953);
nand U19468 (N_19468,N_18602,N_18623);
and U19469 (N_19469,N_18759,N_18673);
nor U19470 (N_19470,N_18609,N_18531);
and U19471 (N_19471,N_18866,N_18579);
nand U19472 (N_19472,N_18526,N_18916);
and U19473 (N_19473,N_18852,N_18715);
nand U19474 (N_19474,N_18508,N_18589);
and U19475 (N_19475,N_18825,N_18702);
nor U19476 (N_19476,N_18882,N_18528);
and U19477 (N_19477,N_18734,N_18732);
and U19478 (N_19478,N_18994,N_18576);
and U19479 (N_19479,N_18986,N_18537);
and U19480 (N_19480,N_18506,N_18836);
and U19481 (N_19481,N_18568,N_18543);
nand U19482 (N_19482,N_18734,N_18973);
or U19483 (N_19483,N_18956,N_18645);
nor U19484 (N_19484,N_18871,N_18915);
nand U19485 (N_19485,N_18624,N_18782);
nor U19486 (N_19486,N_18775,N_18796);
and U19487 (N_19487,N_18636,N_18600);
nor U19488 (N_19488,N_18677,N_18704);
xnor U19489 (N_19489,N_18985,N_18568);
nor U19490 (N_19490,N_18907,N_18630);
xor U19491 (N_19491,N_18565,N_18559);
nand U19492 (N_19492,N_18608,N_18734);
and U19493 (N_19493,N_18836,N_18996);
and U19494 (N_19494,N_18682,N_18725);
nor U19495 (N_19495,N_18854,N_18519);
nand U19496 (N_19496,N_18966,N_18511);
and U19497 (N_19497,N_18777,N_18844);
nand U19498 (N_19498,N_18642,N_18696);
nand U19499 (N_19499,N_18936,N_18561);
nor U19500 (N_19500,N_19264,N_19275);
and U19501 (N_19501,N_19340,N_19008);
or U19502 (N_19502,N_19079,N_19060);
nand U19503 (N_19503,N_19114,N_19042);
nand U19504 (N_19504,N_19150,N_19417);
or U19505 (N_19505,N_19404,N_19333);
nand U19506 (N_19506,N_19483,N_19414);
nand U19507 (N_19507,N_19122,N_19199);
nand U19508 (N_19508,N_19377,N_19294);
nand U19509 (N_19509,N_19397,N_19400);
or U19510 (N_19510,N_19039,N_19229);
xor U19511 (N_19511,N_19019,N_19031);
and U19512 (N_19512,N_19044,N_19286);
nor U19513 (N_19513,N_19211,N_19312);
xnor U19514 (N_19514,N_19452,N_19260);
nor U19515 (N_19515,N_19255,N_19098);
and U19516 (N_19516,N_19296,N_19054);
or U19517 (N_19517,N_19219,N_19324);
or U19518 (N_19518,N_19066,N_19425);
and U19519 (N_19519,N_19259,N_19497);
and U19520 (N_19520,N_19029,N_19491);
or U19521 (N_19521,N_19041,N_19252);
nand U19522 (N_19522,N_19330,N_19113);
and U19523 (N_19523,N_19071,N_19089);
and U19524 (N_19524,N_19266,N_19184);
nand U19525 (N_19525,N_19043,N_19261);
or U19526 (N_19526,N_19145,N_19231);
nand U19527 (N_19527,N_19327,N_19316);
and U19528 (N_19528,N_19137,N_19123);
nor U19529 (N_19529,N_19283,N_19139);
or U19530 (N_19530,N_19362,N_19126);
or U19531 (N_19531,N_19059,N_19157);
or U19532 (N_19532,N_19461,N_19015);
xnor U19533 (N_19533,N_19434,N_19195);
nor U19534 (N_19534,N_19180,N_19418);
nor U19535 (N_19535,N_19445,N_19273);
nor U19536 (N_19536,N_19276,N_19131);
nand U19537 (N_19537,N_19057,N_19058);
nor U19538 (N_19538,N_19037,N_19393);
and U19539 (N_19539,N_19336,N_19119);
nor U19540 (N_19540,N_19419,N_19171);
or U19541 (N_19541,N_19392,N_19238);
xor U19542 (N_19542,N_19099,N_19115);
nor U19543 (N_19543,N_19435,N_19136);
or U19544 (N_19544,N_19111,N_19205);
or U19545 (N_19545,N_19153,N_19374);
nand U19546 (N_19546,N_19475,N_19421);
or U19547 (N_19547,N_19247,N_19314);
xnor U19548 (N_19548,N_19350,N_19226);
xnor U19549 (N_19549,N_19167,N_19258);
or U19550 (N_19550,N_19378,N_19407);
nor U19551 (N_19551,N_19192,N_19103);
nand U19552 (N_19552,N_19141,N_19242);
nor U19553 (N_19553,N_19280,N_19128);
xor U19554 (N_19554,N_19177,N_19228);
nor U19555 (N_19555,N_19225,N_19121);
nor U19556 (N_19556,N_19320,N_19262);
and U19557 (N_19557,N_19387,N_19292);
and U19558 (N_19558,N_19170,N_19040);
nor U19559 (N_19559,N_19299,N_19420);
or U19560 (N_19560,N_19028,N_19000);
nand U19561 (N_19561,N_19210,N_19460);
nor U19562 (N_19562,N_19013,N_19490);
nor U19563 (N_19563,N_19035,N_19376);
and U19564 (N_19564,N_19168,N_19014);
and U19565 (N_19565,N_19117,N_19036);
and U19566 (N_19566,N_19334,N_19457);
nand U19567 (N_19567,N_19124,N_19279);
and U19568 (N_19568,N_19156,N_19337);
nor U19569 (N_19569,N_19001,N_19110);
nand U19570 (N_19570,N_19061,N_19402);
and U19571 (N_19571,N_19482,N_19133);
and U19572 (N_19572,N_19118,N_19464);
and U19573 (N_19573,N_19458,N_19317);
and U19574 (N_19574,N_19391,N_19045);
nor U19575 (N_19575,N_19386,N_19290);
and U19576 (N_19576,N_19331,N_19453);
nand U19577 (N_19577,N_19096,N_19382);
nand U19578 (N_19578,N_19499,N_19351);
and U19579 (N_19579,N_19467,N_19289);
and U19580 (N_19580,N_19183,N_19373);
nand U19581 (N_19581,N_19318,N_19053);
nand U19582 (N_19582,N_19097,N_19143);
and U19583 (N_19583,N_19193,N_19429);
nor U19584 (N_19584,N_19249,N_19448);
nor U19585 (N_19585,N_19257,N_19227);
and U19586 (N_19586,N_19284,N_19415);
nand U19587 (N_19587,N_19194,N_19438);
and U19588 (N_19588,N_19295,N_19368);
or U19589 (N_19589,N_19465,N_19138);
and U19590 (N_19590,N_19010,N_19152);
and U19591 (N_19591,N_19451,N_19088);
nand U19592 (N_19592,N_19367,N_19070);
and U19593 (N_19593,N_19485,N_19388);
and U19594 (N_19594,N_19444,N_19024);
and U19595 (N_19595,N_19178,N_19263);
and U19596 (N_19596,N_19006,N_19078);
nand U19597 (N_19597,N_19161,N_19248);
and U19598 (N_19598,N_19056,N_19081);
nor U19599 (N_19599,N_19215,N_19106);
xor U19600 (N_19600,N_19379,N_19309);
nand U19601 (N_19601,N_19441,N_19271);
nand U19602 (N_19602,N_19343,N_19495);
or U19603 (N_19603,N_19162,N_19033);
nor U19604 (N_19604,N_19307,N_19241);
xor U19605 (N_19605,N_19086,N_19109);
xor U19606 (N_19606,N_19322,N_19147);
or U19607 (N_19607,N_19481,N_19370);
nand U19608 (N_19608,N_19394,N_19371);
or U19609 (N_19609,N_19403,N_19342);
or U19610 (N_19610,N_19220,N_19017);
and U19611 (N_19611,N_19234,N_19354);
nor U19612 (N_19612,N_19470,N_19038);
nand U19613 (N_19613,N_19338,N_19052);
and U19614 (N_19614,N_19236,N_19101);
xor U19615 (N_19615,N_19197,N_19108);
nor U19616 (N_19616,N_19065,N_19357);
xnor U19617 (N_19617,N_19450,N_19004);
nor U19618 (N_19618,N_19233,N_19440);
nand U19619 (N_19619,N_19218,N_19237);
nor U19620 (N_19620,N_19068,N_19353);
nand U19621 (N_19621,N_19206,N_19486);
xnor U19622 (N_19622,N_19426,N_19213);
nand U19623 (N_19623,N_19256,N_19472);
or U19624 (N_19624,N_19149,N_19186);
nand U19625 (N_19625,N_19478,N_19332);
nor U19626 (N_19626,N_19127,N_19468);
xnor U19627 (N_19627,N_19191,N_19423);
nand U19628 (N_19628,N_19254,N_19090);
xor U19629 (N_19629,N_19087,N_19454);
nand U19630 (N_19630,N_19442,N_19094);
or U19631 (N_19631,N_19174,N_19428);
and U19632 (N_19632,N_19265,N_19329);
xor U19633 (N_19633,N_19480,N_19072);
nand U19634 (N_19634,N_19411,N_19185);
or U19635 (N_19635,N_19047,N_19496);
or U19636 (N_19636,N_19319,N_19134);
xnor U19637 (N_19637,N_19020,N_19239);
nand U19638 (N_19638,N_19055,N_19268);
and U19639 (N_19639,N_19462,N_19463);
nor U19640 (N_19640,N_19356,N_19176);
nand U19641 (N_19641,N_19471,N_19422);
nor U19642 (N_19642,N_19477,N_19344);
and U19643 (N_19643,N_19146,N_19204);
nand U19644 (N_19644,N_19196,N_19437);
nor U19645 (N_19645,N_19278,N_19120);
or U19646 (N_19646,N_19365,N_19446);
and U19647 (N_19647,N_19409,N_19433);
nand U19648 (N_19648,N_19214,N_19396);
or U19649 (N_19649,N_19075,N_19315);
or U19650 (N_19650,N_19169,N_19083);
and U19651 (N_19651,N_19251,N_19303);
nor U19652 (N_19652,N_19148,N_19160);
and U19653 (N_19653,N_19172,N_19240);
nand U19654 (N_19654,N_19125,N_19436);
and U19655 (N_19655,N_19355,N_19287);
nor U19656 (N_19656,N_19381,N_19005);
nor U19657 (N_19657,N_19372,N_19476);
nand U19658 (N_19658,N_19474,N_19449);
nor U19659 (N_19659,N_19200,N_19140);
nand U19660 (N_19660,N_19144,N_19455);
xnor U19661 (N_19661,N_19363,N_19401);
and U19662 (N_19662,N_19107,N_19298);
or U19663 (N_19663,N_19395,N_19027);
nor U19664 (N_19664,N_19085,N_19484);
nor U19665 (N_19665,N_19003,N_19216);
nand U19666 (N_19666,N_19092,N_19305);
nand U19667 (N_19667,N_19253,N_19439);
nand U19668 (N_19668,N_19235,N_19328);
and U19669 (N_19669,N_19269,N_19100);
and U19670 (N_19670,N_19424,N_19369);
or U19671 (N_19671,N_19012,N_19282);
or U19672 (N_19672,N_19026,N_19281);
nand U19673 (N_19673,N_19189,N_19300);
and U19674 (N_19674,N_19223,N_19416);
nor U19675 (N_19675,N_19095,N_19212);
nand U19676 (N_19676,N_19456,N_19142);
xnor U19677 (N_19677,N_19306,N_19224);
xor U19678 (N_19678,N_19166,N_19188);
or U19679 (N_19679,N_19366,N_19132);
nor U19680 (N_19680,N_19492,N_19018);
nand U19681 (N_19681,N_19375,N_19301);
nor U19682 (N_19682,N_19104,N_19341);
nand U19683 (N_19683,N_19202,N_19201);
or U19684 (N_19684,N_19349,N_19359);
xor U19685 (N_19685,N_19181,N_19165);
nor U19686 (N_19686,N_19347,N_19022);
or U19687 (N_19687,N_19348,N_19431);
nor U19688 (N_19688,N_19390,N_19410);
xnor U19689 (N_19689,N_19105,N_19048);
or U19690 (N_19690,N_19297,N_19339);
or U19691 (N_19691,N_19073,N_19002);
or U19692 (N_19692,N_19313,N_19067);
or U19693 (N_19693,N_19064,N_19291);
nor U19694 (N_19694,N_19062,N_19032);
or U19695 (N_19695,N_19361,N_19326);
or U19696 (N_19696,N_19209,N_19245);
xor U19697 (N_19697,N_19198,N_19345);
nand U19698 (N_19698,N_19335,N_19288);
nand U19699 (N_19699,N_19389,N_19405);
nand U19700 (N_19700,N_19116,N_19173);
or U19701 (N_19701,N_19063,N_19473);
and U19702 (N_19702,N_19159,N_19091);
and U19703 (N_19703,N_19250,N_19267);
nand U19704 (N_19704,N_19221,N_19102);
xor U19705 (N_19705,N_19222,N_19077);
and U19706 (N_19706,N_19398,N_19302);
xnor U19707 (N_19707,N_19208,N_19084);
nand U19708 (N_19708,N_19182,N_19025);
or U19709 (N_19709,N_19074,N_19154);
or U19710 (N_19710,N_19246,N_19230);
or U19711 (N_19711,N_19459,N_19479);
nand U19712 (N_19712,N_19380,N_19155);
or U19713 (N_19713,N_19408,N_19488);
and U19714 (N_19714,N_19443,N_19270);
nor U19715 (N_19715,N_19030,N_19011);
or U19716 (N_19716,N_19399,N_19207);
nand U19717 (N_19717,N_19430,N_19346);
nand U19718 (N_19718,N_19413,N_19244);
xor U19719 (N_19719,N_19323,N_19384);
nor U19720 (N_19720,N_19325,N_19023);
nand U19721 (N_19721,N_19076,N_19164);
nand U19722 (N_19722,N_19272,N_19308);
xnor U19723 (N_19723,N_19469,N_19217);
nand U19724 (N_19724,N_19051,N_19179);
nor U19725 (N_19725,N_19360,N_19129);
and U19726 (N_19726,N_19321,N_19158);
nor U19727 (N_19727,N_19447,N_19494);
xnor U19728 (N_19728,N_19310,N_19069);
nand U19729 (N_19729,N_19358,N_19082);
nand U19730 (N_19730,N_19112,N_19489);
nor U19731 (N_19731,N_19304,N_19163);
or U19732 (N_19732,N_19187,N_19093);
nor U19733 (N_19733,N_19427,N_19151);
nand U19734 (N_19734,N_19487,N_19175);
or U19735 (N_19735,N_19130,N_19232);
nand U19736 (N_19736,N_19412,N_19034);
nand U19737 (N_19737,N_19466,N_19352);
or U19738 (N_19738,N_19406,N_19009);
and U19739 (N_19739,N_19243,N_19046);
nand U19740 (N_19740,N_19080,N_19190);
or U19741 (N_19741,N_19049,N_19274);
xor U19742 (N_19742,N_19432,N_19021);
nor U19743 (N_19743,N_19383,N_19016);
and U19744 (N_19744,N_19385,N_19498);
and U19745 (N_19745,N_19493,N_19007);
and U19746 (N_19746,N_19203,N_19364);
nand U19747 (N_19747,N_19293,N_19135);
nand U19748 (N_19748,N_19050,N_19277);
nand U19749 (N_19749,N_19311,N_19285);
and U19750 (N_19750,N_19076,N_19080);
or U19751 (N_19751,N_19130,N_19047);
nor U19752 (N_19752,N_19430,N_19011);
nand U19753 (N_19753,N_19295,N_19314);
or U19754 (N_19754,N_19417,N_19403);
or U19755 (N_19755,N_19254,N_19499);
nand U19756 (N_19756,N_19013,N_19223);
or U19757 (N_19757,N_19439,N_19207);
nand U19758 (N_19758,N_19062,N_19474);
nand U19759 (N_19759,N_19489,N_19121);
or U19760 (N_19760,N_19155,N_19445);
and U19761 (N_19761,N_19278,N_19185);
or U19762 (N_19762,N_19329,N_19495);
xnor U19763 (N_19763,N_19482,N_19164);
or U19764 (N_19764,N_19306,N_19042);
and U19765 (N_19765,N_19285,N_19135);
nand U19766 (N_19766,N_19266,N_19340);
nor U19767 (N_19767,N_19229,N_19036);
xnor U19768 (N_19768,N_19110,N_19383);
and U19769 (N_19769,N_19371,N_19338);
or U19770 (N_19770,N_19468,N_19484);
xnor U19771 (N_19771,N_19200,N_19466);
nand U19772 (N_19772,N_19183,N_19165);
nand U19773 (N_19773,N_19395,N_19009);
nor U19774 (N_19774,N_19321,N_19092);
nor U19775 (N_19775,N_19388,N_19314);
nor U19776 (N_19776,N_19485,N_19087);
xor U19777 (N_19777,N_19089,N_19318);
and U19778 (N_19778,N_19135,N_19171);
nor U19779 (N_19779,N_19325,N_19089);
nor U19780 (N_19780,N_19317,N_19234);
nand U19781 (N_19781,N_19356,N_19226);
nor U19782 (N_19782,N_19278,N_19495);
nand U19783 (N_19783,N_19073,N_19364);
or U19784 (N_19784,N_19048,N_19009);
nor U19785 (N_19785,N_19338,N_19068);
xor U19786 (N_19786,N_19189,N_19358);
nand U19787 (N_19787,N_19179,N_19483);
and U19788 (N_19788,N_19079,N_19109);
nor U19789 (N_19789,N_19325,N_19141);
xnor U19790 (N_19790,N_19021,N_19425);
nand U19791 (N_19791,N_19078,N_19401);
nand U19792 (N_19792,N_19474,N_19168);
nand U19793 (N_19793,N_19359,N_19423);
nor U19794 (N_19794,N_19093,N_19009);
or U19795 (N_19795,N_19215,N_19234);
or U19796 (N_19796,N_19293,N_19423);
nor U19797 (N_19797,N_19406,N_19036);
nand U19798 (N_19798,N_19299,N_19339);
or U19799 (N_19799,N_19322,N_19333);
nor U19800 (N_19800,N_19073,N_19072);
nor U19801 (N_19801,N_19460,N_19101);
and U19802 (N_19802,N_19448,N_19494);
or U19803 (N_19803,N_19020,N_19206);
xnor U19804 (N_19804,N_19350,N_19188);
or U19805 (N_19805,N_19304,N_19331);
or U19806 (N_19806,N_19232,N_19368);
nand U19807 (N_19807,N_19335,N_19006);
and U19808 (N_19808,N_19109,N_19369);
or U19809 (N_19809,N_19149,N_19388);
nand U19810 (N_19810,N_19029,N_19338);
nor U19811 (N_19811,N_19192,N_19116);
nand U19812 (N_19812,N_19279,N_19194);
xor U19813 (N_19813,N_19478,N_19433);
and U19814 (N_19814,N_19391,N_19256);
or U19815 (N_19815,N_19333,N_19337);
or U19816 (N_19816,N_19491,N_19452);
or U19817 (N_19817,N_19345,N_19426);
nor U19818 (N_19818,N_19275,N_19017);
or U19819 (N_19819,N_19399,N_19079);
nand U19820 (N_19820,N_19323,N_19133);
nand U19821 (N_19821,N_19295,N_19390);
and U19822 (N_19822,N_19283,N_19432);
nand U19823 (N_19823,N_19125,N_19465);
nor U19824 (N_19824,N_19233,N_19483);
nor U19825 (N_19825,N_19161,N_19140);
and U19826 (N_19826,N_19441,N_19433);
nor U19827 (N_19827,N_19374,N_19498);
nand U19828 (N_19828,N_19227,N_19418);
nand U19829 (N_19829,N_19150,N_19399);
or U19830 (N_19830,N_19027,N_19077);
or U19831 (N_19831,N_19469,N_19162);
or U19832 (N_19832,N_19202,N_19081);
nand U19833 (N_19833,N_19250,N_19386);
and U19834 (N_19834,N_19437,N_19378);
or U19835 (N_19835,N_19263,N_19088);
and U19836 (N_19836,N_19270,N_19438);
nor U19837 (N_19837,N_19404,N_19090);
and U19838 (N_19838,N_19106,N_19123);
nor U19839 (N_19839,N_19164,N_19156);
nor U19840 (N_19840,N_19291,N_19480);
or U19841 (N_19841,N_19476,N_19365);
nand U19842 (N_19842,N_19284,N_19333);
or U19843 (N_19843,N_19109,N_19223);
xnor U19844 (N_19844,N_19233,N_19408);
or U19845 (N_19845,N_19231,N_19328);
nor U19846 (N_19846,N_19065,N_19451);
or U19847 (N_19847,N_19108,N_19037);
and U19848 (N_19848,N_19011,N_19418);
xor U19849 (N_19849,N_19412,N_19429);
nor U19850 (N_19850,N_19278,N_19178);
xnor U19851 (N_19851,N_19061,N_19054);
nand U19852 (N_19852,N_19231,N_19394);
and U19853 (N_19853,N_19285,N_19283);
nor U19854 (N_19854,N_19237,N_19224);
or U19855 (N_19855,N_19241,N_19446);
nor U19856 (N_19856,N_19302,N_19381);
or U19857 (N_19857,N_19292,N_19009);
nand U19858 (N_19858,N_19184,N_19403);
or U19859 (N_19859,N_19214,N_19025);
and U19860 (N_19860,N_19367,N_19072);
nand U19861 (N_19861,N_19146,N_19344);
or U19862 (N_19862,N_19369,N_19254);
nor U19863 (N_19863,N_19254,N_19456);
nand U19864 (N_19864,N_19307,N_19402);
xnor U19865 (N_19865,N_19298,N_19216);
or U19866 (N_19866,N_19383,N_19438);
or U19867 (N_19867,N_19294,N_19391);
nand U19868 (N_19868,N_19151,N_19085);
nand U19869 (N_19869,N_19155,N_19356);
nor U19870 (N_19870,N_19256,N_19323);
or U19871 (N_19871,N_19378,N_19122);
nand U19872 (N_19872,N_19332,N_19042);
nor U19873 (N_19873,N_19021,N_19433);
or U19874 (N_19874,N_19103,N_19115);
nor U19875 (N_19875,N_19336,N_19021);
and U19876 (N_19876,N_19052,N_19465);
or U19877 (N_19877,N_19142,N_19013);
and U19878 (N_19878,N_19188,N_19098);
nor U19879 (N_19879,N_19114,N_19096);
nand U19880 (N_19880,N_19060,N_19131);
and U19881 (N_19881,N_19183,N_19045);
nor U19882 (N_19882,N_19406,N_19267);
xor U19883 (N_19883,N_19057,N_19259);
and U19884 (N_19884,N_19092,N_19430);
nand U19885 (N_19885,N_19088,N_19184);
or U19886 (N_19886,N_19342,N_19448);
or U19887 (N_19887,N_19303,N_19033);
nand U19888 (N_19888,N_19336,N_19266);
nand U19889 (N_19889,N_19077,N_19112);
nand U19890 (N_19890,N_19386,N_19006);
nor U19891 (N_19891,N_19232,N_19106);
nor U19892 (N_19892,N_19416,N_19498);
nor U19893 (N_19893,N_19151,N_19377);
or U19894 (N_19894,N_19203,N_19368);
and U19895 (N_19895,N_19113,N_19345);
nand U19896 (N_19896,N_19388,N_19165);
xor U19897 (N_19897,N_19022,N_19240);
and U19898 (N_19898,N_19398,N_19150);
and U19899 (N_19899,N_19369,N_19216);
and U19900 (N_19900,N_19209,N_19013);
and U19901 (N_19901,N_19103,N_19216);
nor U19902 (N_19902,N_19174,N_19259);
or U19903 (N_19903,N_19204,N_19301);
nand U19904 (N_19904,N_19174,N_19054);
nand U19905 (N_19905,N_19345,N_19125);
or U19906 (N_19906,N_19366,N_19393);
nor U19907 (N_19907,N_19289,N_19072);
nor U19908 (N_19908,N_19411,N_19068);
nand U19909 (N_19909,N_19376,N_19436);
nor U19910 (N_19910,N_19307,N_19076);
nor U19911 (N_19911,N_19099,N_19202);
or U19912 (N_19912,N_19358,N_19207);
or U19913 (N_19913,N_19131,N_19377);
xnor U19914 (N_19914,N_19203,N_19161);
or U19915 (N_19915,N_19058,N_19031);
nand U19916 (N_19916,N_19475,N_19169);
nor U19917 (N_19917,N_19279,N_19049);
xnor U19918 (N_19918,N_19434,N_19482);
nand U19919 (N_19919,N_19249,N_19127);
nand U19920 (N_19920,N_19398,N_19499);
or U19921 (N_19921,N_19312,N_19446);
nand U19922 (N_19922,N_19486,N_19183);
or U19923 (N_19923,N_19314,N_19044);
nor U19924 (N_19924,N_19279,N_19438);
nand U19925 (N_19925,N_19195,N_19201);
nor U19926 (N_19926,N_19085,N_19444);
xnor U19927 (N_19927,N_19131,N_19263);
and U19928 (N_19928,N_19270,N_19440);
or U19929 (N_19929,N_19438,N_19060);
nand U19930 (N_19930,N_19425,N_19312);
nand U19931 (N_19931,N_19202,N_19166);
xnor U19932 (N_19932,N_19203,N_19125);
nand U19933 (N_19933,N_19497,N_19430);
nor U19934 (N_19934,N_19080,N_19349);
nor U19935 (N_19935,N_19052,N_19355);
nand U19936 (N_19936,N_19069,N_19308);
or U19937 (N_19937,N_19450,N_19375);
and U19938 (N_19938,N_19329,N_19307);
xnor U19939 (N_19939,N_19038,N_19432);
xor U19940 (N_19940,N_19116,N_19304);
or U19941 (N_19941,N_19118,N_19041);
nand U19942 (N_19942,N_19157,N_19054);
and U19943 (N_19943,N_19028,N_19321);
and U19944 (N_19944,N_19000,N_19362);
and U19945 (N_19945,N_19407,N_19135);
nor U19946 (N_19946,N_19204,N_19098);
nor U19947 (N_19947,N_19347,N_19064);
and U19948 (N_19948,N_19421,N_19205);
nand U19949 (N_19949,N_19187,N_19499);
or U19950 (N_19950,N_19177,N_19466);
nor U19951 (N_19951,N_19362,N_19089);
xor U19952 (N_19952,N_19164,N_19438);
or U19953 (N_19953,N_19338,N_19195);
nor U19954 (N_19954,N_19470,N_19120);
or U19955 (N_19955,N_19136,N_19172);
nand U19956 (N_19956,N_19215,N_19243);
nor U19957 (N_19957,N_19311,N_19448);
xnor U19958 (N_19958,N_19062,N_19475);
xnor U19959 (N_19959,N_19085,N_19194);
or U19960 (N_19960,N_19445,N_19201);
or U19961 (N_19961,N_19356,N_19151);
xnor U19962 (N_19962,N_19233,N_19246);
nor U19963 (N_19963,N_19019,N_19025);
nor U19964 (N_19964,N_19067,N_19415);
and U19965 (N_19965,N_19448,N_19015);
or U19966 (N_19966,N_19117,N_19302);
nand U19967 (N_19967,N_19030,N_19480);
nor U19968 (N_19968,N_19083,N_19016);
and U19969 (N_19969,N_19026,N_19468);
nand U19970 (N_19970,N_19019,N_19018);
nand U19971 (N_19971,N_19165,N_19288);
xnor U19972 (N_19972,N_19125,N_19268);
and U19973 (N_19973,N_19252,N_19437);
nand U19974 (N_19974,N_19457,N_19291);
or U19975 (N_19975,N_19380,N_19415);
and U19976 (N_19976,N_19128,N_19181);
nor U19977 (N_19977,N_19382,N_19392);
nand U19978 (N_19978,N_19191,N_19160);
nand U19979 (N_19979,N_19288,N_19444);
nor U19980 (N_19980,N_19225,N_19254);
or U19981 (N_19981,N_19036,N_19297);
or U19982 (N_19982,N_19032,N_19043);
nand U19983 (N_19983,N_19129,N_19044);
or U19984 (N_19984,N_19481,N_19444);
or U19985 (N_19985,N_19474,N_19310);
nand U19986 (N_19986,N_19420,N_19111);
and U19987 (N_19987,N_19486,N_19428);
or U19988 (N_19988,N_19016,N_19463);
or U19989 (N_19989,N_19336,N_19247);
nand U19990 (N_19990,N_19431,N_19022);
nor U19991 (N_19991,N_19141,N_19385);
and U19992 (N_19992,N_19281,N_19030);
and U19993 (N_19993,N_19243,N_19384);
nor U19994 (N_19994,N_19175,N_19191);
and U19995 (N_19995,N_19325,N_19027);
xor U19996 (N_19996,N_19179,N_19117);
nand U19997 (N_19997,N_19113,N_19439);
or U19998 (N_19998,N_19365,N_19374);
or U19999 (N_19999,N_19412,N_19104);
nand U20000 (N_20000,N_19541,N_19860);
nor U20001 (N_20001,N_19795,N_19813);
xnor U20002 (N_20002,N_19861,N_19705);
nand U20003 (N_20003,N_19605,N_19547);
nor U20004 (N_20004,N_19846,N_19582);
or U20005 (N_20005,N_19730,N_19986);
nor U20006 (N_20006,N_19727,N_19634);
and U20007 (N_20007,N_19517,N_19820);
nor U20008 (N_20008,N_19892,N_19809);
nand U20009 (N_20009,N_19803,N_19557);
xnor U20010 (N_20010,N_19504,N_19949);
nand U20011 (N_20011,N_19982,N_19937);
nor U20012 (N_20012,N_19510,N_19755);
nand U20013 (N_20013,N_19881,N_19550);
and U20014 (N_20014,N_19689,N_19816);
nand U20015 (N_20015,N_19643,N_19930);
and U20016 (N_20016,N_19704,N_19542);
or U20017 (N_20017,N_19945,N_19874);
or U20018 (N_20018,N_19898,N_19878);
or U20019 (N_20019,N_19528,N_19680);
and U20020 (N_20020,N_19978,N_19926);
and U20021 (N_20021,N_19902,N_19909);
or U20022 (N_20022,N_19932,N_19800);
nor U20023 (N_20023,N_19645,N_19920);
nor U20024 (N_20024,N_19774,N_19931);
and U20025 (N_20025,N_19770,N_19654);
nor U20026 (N_20026,N_19596,N_19951);
nor U20027 (N_20027,N_19533,N_19628);
nor U20028 (N_20028,N_19658,N_19501);
xnor U20029 (N_20029,N_19888,N_19530);
and U20030 (N_20030,N_19839,N_19642);
and U20031 (N_20031,N_19551,N_19996);
and U20032 (N_20032,N_19841,N_19783);
or U20033 (N_20033,N_19655,N_19619);
xnor U20034 (N_20034,N_19999,N_19757);
nor U20035 (N_20035,N_19553,N_19821);
nand U20036 (N_20036,N_19767,N_19769);
xor U20037 (N_20037,N_19500,N_19648);
and U20038 (N_20038,N_19649,N_19956);
or U20039 (N_20039,N_19880,N_19873);
xor U20040 (N_20040,N_19641,N_19670);
nand U20041 (N_20041,N_19725,N_19682);
nand U20042 (N_20042,N_19879,N_19513);
nand U20043 (N_20043,N_19815,N_19918);
xor U20044 (N_20044,N_19904,N_19693);
xnor U20045 (N_20045,N_19636,N_19721);
nand U20046 (N_20046,N_19690,N_19685);
nand U20047 (N_20047,N_19984,N_19611);
nand U20048 (N_20048,N_19968,N_19589);
and U20049 (N_20049,N_19538,N_19561);
and U20050 (N_20050,N_19570,N_19775);
nor U20051 (N_20051,N_19614,N_19586);
or U20052 (N_20052,N_19985,N_19762);
and U20053 (N_20053,N_19992,N_19671);
nor U20054 (N_20054,N_19600,N_19876);
nor U20055 (N_20055,N_19965,N_19509);
or U20056 (N_20056,N_19975,N_19919);
nor U20057 (N_20057,N_19793,N_19905);
or U20058 (N_20058,N_19679,N_19805);
or U20059 (N_20059,N_19971,N_19806);
nand U20060 (N_20060,N_19523,N_19691);
or U20061 (N_20061,N_19778,N_19872);
nand U20062 (N_20062,N_19753,N_19777);
and U20063 (N_20063,N_19781,N_19980);
and U20064 (N_20064,N_19663,N_19540);
or U20065 (N_20065,N_19864,N_19866);
or U20066 (N_20066,N_19592,N_19745);
and U20067 (N_20067,N_19626,N_19632);
nor U20068 (N_20068,N_19773,N_19812);
nor U20069 (N_20069,N_19667,N_19531);
and U20070 (N_20070,N_19681,N_19676);
nand U20071 (N_20071,N_19807,N_19970);
nand U20072 (N_20072,N_19894,N_19752);
nand U20073 (N_20073,N_19695,N_19917);
xnor U20074 (N_20074,N_19532,N_19733);
nand U20075 (N_20075,N_19644,N_19673);
or U20076 (N_20076,N_19928,N_19903);
nor U20077 (N_20077,N_19855,N_19686);
nand U20078 (N_20078,N_19683,N_19871);
nor U20079 (N_20079,N_19884,N_19943);
nand U20080 (N_20080,N_19665,N_19997);
nor U20081 (N_20081,N_19936,N_19732);
or U20082 (N_20082,N_19606,N_19857);
xnor U20083 (N_20083,N_19656,N_19722);
nor U20084 (N_20084,N_19955,N_19837);
nand U20085 (N_20085,N_19507,N_19870);
nand U20086 (N_20086,N_19948,N_19647);
nand U20087 (N_20087,N_19572,N_19818);
and U20088 (N_20088,N_19962,N_19520);
or U20089 (N_20089,N_19651,N_19906);
nand U20090 (N_20090,N_19838,N_19819);
or U20091 (N_20091,N_19941,N_19741);
nand U20092 (N_20092,N_19579,N_19785);
nand U20093 (N_20093,N_19843,N_19895);
or U20094 (N_20094,N_19696,N_19766);
or U20095 (N_20095,N_19938,N_19811);
and U20096 (N_20096,N_19739,N_19633);
nand U20097 (N_20097,N_19604,N_19743);
and U20098 (N_20098,N_19516,N_19758);
or U20099 (N_20099,N_19735,N_19684);
or U20100 (N_20100,N_19840,N_19719);
nand U20101 (N_20101,N_19525,N_19503);
or U20102 (N_20102,N_19953,N_19768);
and U20103 (N_20103,N_19529,N_19581);
and U20104 (N_20104,N_19590,N_19567);
and U20105 (N_20105,N_19574,N_19521);
nand U20106 (N_20106,N_19519,N_19585);
nand U20107 (N_20107,N_19786,N_19502);
or U20108 (N_20108,N_19573,N_19833);
nand U20109 (N_20109,N_19865,N_19858);
nand U20110 (N_20110,N_19921,N_19674);
and U20111 (N_20111,N_19568,N_19896);
nand U20112 (N_20112,N_19908,N_19973);
and U20113 (N_20113,N_19830,N_19694);
and U20114 (N_20114,N_19514,N_19713);
xor U20115 (N_20115,N_19802,N_19964);
nand U20116 (N_20116,N_19615,N_19701);
nor U20117 (N_20117,N_19867,N_19669);
xnor U20118 (N_20118,N_19933,N_19979);
or U20119 (N_20119,N_19637,N_19848);
nand U20120 (N_20120,N_19515,N_19749);
nor U20121 (N_20121,N_19737,N_19765);
nor U20122 (N_20122,N_19844,N_19534);
nand U20123 (N_20123,N_19672,N_19863);
xnor U20124 (N_20124,N_19664,N_19899);
nor U20125 (N_20125,N_19627,N_19527);
nand U20126 (N_20126,N_19804,N_19912);
xnor U20127 (N_20127,N_19823,N_19708);
or U20128 (N_20128,N_19554,N_19960);
xor U20129 (N_20129,N_19677,N_19620);
nand U20130 (N_20130,N_19607,N_19524);
and U20131 (N_20131,N_19635,N_19729);
nand U20132 (N_20132,N_19958,N_19886);
or U20133 (N_20133,N_19856,N_19624);
xnor U20134 (N_20134,N_19961,N_19666);
and U20135 (N_20135,N_19559,N_19522);
or U20136 (N_20136,N_19911,N_19703);
nand U20137 (N_20137,N_19709,N_19613);
and U20138 (N_20138,N_19817,N_19789);
nor U20139 (N_20139,N_19990,N_19814);
nand U20140 (N_20140,N_19575,N_19782);
and U20141 (N_20141,N_19639,N_19983);
nand U20142 (N_20142,N_19697,N_19560);
and U20143 (N_20143,N_19969,N_19720);
and U20144 (N_20144,N_19652,N_19834);
and U20145 (N_20145,N_19712,N_19772);
nor U20146 (N_20146,N_19678,N_19610);
xor U20147 (N_20147,N_19646,N_19734);
and U20148 (N_20148,N_19631,N_19890);
or U20149 (N_20149,N_19850,N_19508);
nand U20150 (N_20150,N_19593,N_19959);
nand U20151 (N_20151,N_19927,N_19854);
or U20152 (N_20152,N_19609,N_19847);
nor U20153 (N_20153,N_19638,N_19788);
or U20154 (N_20154,N_19728,N_19954);
nand U20155 (N_20155,N_19603,N_19535);
and U20156 (N_20156,N_19750,N_19602);
and U20157 (N_20157,N_19849,N_19944);
or U20158 (N_20158,N_19711,N_19588);
and U20159 (N_20159,N_19562,N_19915);
nor U20160 (N_20160,N_19976,N_19594);
nand U20161 (N_20161,N_19763,N_19836);
and U20162 (N_20162,N_19660,N_19564);
nor U20163 (N_20163,N_19640,N_19947);
nand U20164 (N_20164,N_19612,N_19731);
and U20165 (N_20165,N_19952,N_19842);
and U20166 (N_20166,N_19591,N_19548);
xor U20167 (N_20167,N_19736,N_19875);
or U20168 (N_20168,N_19630,N_19717);
or U20169 (N_20169,N_19563,N_19577);
nor U20170 (N_20170,N_19887,N_19511);
nor U20171 (N_20171,N_19650,N_19893);
and U20172 (N_20172,N_19852,N_19518);
nand U20173 (N_20173,N_19580,N_19756);
and U20174 (N_20174,N_19549,N_19707);
xor U20175 (N_20175,N_19558,N_19761);
and U20176 (N_20176,N_19827,N_19826);
or U20177 (N_20177,N_19718,N_19784);
xnor U20178 (N_20178,N_19608,N_19617);
or U20179 (N_20179,N_19897,N_19539);
or U20180 (N_20180,N_19710,N_19618);
or U20181 (N_20181,N_19877,N_19966);
xnor U20182 (N_20182,N_19883,N_19692);
nor U20183 (N_20183,N_19747,N_19862);
and U20184 (N_20184,N_19859,N_19601);
or U20185 (N_20185,N_19543,N_19832);
or U20186 (N_20186,N_19885,N_19702);
or U20187 (N_20187,N_19578,N_19565);
nand U20188 (N_20188,N_19923,N_19963);
nand U20189 (N_20189,N_19796,N_19714);
xnor U20190 (N_20190,N_19584,N_19993);
xor U20191 (N_20191,N_19913,N_19662);
nand U20192 (N_20192,N_19653,N_19587);
and U20193 (N_20193,N_19835,N_19506);
or U20194 (N_20194,N_19910,N_19576);
or U20195 (N_20195,N_19657,N_19698);
nor U20196 (N_20196,N_19598,N_19723);
xnor U20197 (N_20197,N_19790,N_19629);
nand U20198 (N_20198,N_19566,N_19889);
nor U20199 (N_20199,N_19668,N_19597);
or U20200 (N_20200,N_19799,N_19661);
nor U20201 (N_20201,N_19925,N_19780);
or U20202 (N_20202,N_19829,N_19792);
nor U20203 (N_20203,N_19791,N_19569);
or U20204 (N_20204,N_19748,N_19798);
or U20205 (N_20205,N_19744,N_19740);
nand U20206 (N_20206,N_19544,N_19760);
or U20207 (N_20207,N_19505,N_19746);
nor U20208 (N_20208,N_19801,N_19981);
xor U20209 (N_20209,N_19616,N_19512);
and U20210 (N_20210,N_19779,N_19688);
nand U20211 (N_20211,N_19942,N_19810);
xor U20212 (N_20212,N_19764,N_19939);
or U20213 (N_20213,N_19808,N_19715);
and U20214 (N_20214,N_19845,N_19991);
xnor U20215 (N_20215,N_19716,N_19950);
nor U20216 (N_20216,N_19940,N_19555);
nand U20217 (N_20217,N_19891,N_19995);
and U20218 (N_20218,N_19935,N_19797);
nand U20219 (N_20219,N_19552,N_19687);
nand U20220 (N_20220,N_19831,N_19571);
and U20221 (N_20221,N_19901,N_19623);
nor U20222 (N_20222,N_19595,N_19726);
or U20223 (N_20223,N_19851,N_19699);
or U20224 (N_20224,N_19526,N_19972);
nand U20225 (N_20225,N_19868,N_19700);
nor U20226 (N_20226,N_19869,N_19853);
or U20227 (N_20227,N_19922,N_19622);
nor U20228 (N_20228,N_19934,N_19583);
or U20229 (N_20229,N_19882,N_19974);
nand U20230 (N_20230,N_19546,N_19536);
and U20231 (N_20231,N_19825,N_19599);
or U20232 (N_20232,N_19659,N_19924);
nand U20233 (N_20233,N_19989,N_19537);
nor U20234 (N_20234,N_19771,N_19545);
nor U20235 (N_20235,N_19957,N_19625);
nor U20236 (N_20236,N_19759,N_19742);
or U20237 (N_20237,N_19907,N_19724);
and U20238 (N_20238,N_19776,N_19994);
and U20239 (N_20239,N_19914,N_19822);
and U20240 (N_20240,N_19988,N_19998);
or U20241 (N_20241,N_19900,N_19977);
and U20242 (N_20242,N_19621,N_19787);
nand U20243 (N_20243,N_19675,N_19946);
nor U20244 (N_20244,N_19828,N_19929);
nor U20245 (N_20245,N_19967,N_19751);
xnor U20246 (N_20246,N_19706,N_19754);
nand U20247 (N_20247,N_19824,N_19556);
and U20248 (N_20248,N_19738,N_19987);
or U20249 (N_20249,N_19916,N_19794);
and U20250 (N_20250,N_19803,N_19857);
and U20251 (N_20251,N_19693,N_19875);
and U20252 (N_20252,N_19850,N_19935);
and U20253 (N_20253,N_19771,N_19847);
and U20254 (N_20254,N_19822,N_19871);
or U20255 (N_20255,N_19966,N_19585);
and U20256 (N_20256,N_19659,N_19675);
or U20257 (N_20257,N_19881,N_19825);
nor U20258 (N_20258,N_19918,N_19643);
xor U20259 (N_20259,N_19842,N_19686);
nand U20260 (N_20260,N_19568,N_19577);
or U20261 (N_20261,N_19703,N_19907);
nand U20262 (N_20262,N_19652,N_19705);
nand U20263 (N_20263,N_19945,N_19776);
and U20264 (N_20264,N_19973,N_19809);
nor U20265 (N_20265,N_19745,N_19772);
and U20266 (N_20266,N_19890,N_19550);
nand U20267 (N_20267,N_19851,N_19789);
nor U20268 (N_20268,N_19638,N_19885);
xor U20269 (N_20269,N_19783,N_19663);
nand U20270 (N_20270,N_19650,N_19856);
nor U20271 (N_20271,N_19518,N_19751);
xor U20272 (N_20272,N_19584,N_19960);
xnor U20273 (N_20273,N_19787,N_19888);
xnor U20274 (N_20274,N_19747,N_19611);
or U20275 (N_20275,N_19660,N_19771);
nor U20276 (N_20276,N_19702,N_19962);
and U20277 (N_20277,N_19938,N_19511);
nor U20278 (N_20278,N_19645,N_19672);
and U20279 (N_20279,N_19655,N_19579);
or U20280 (N_20280,N_19724,N_19586);
nand U20281 (N_20281,N_19767,N_19532);
nand U20282 (N_20282,N_19910,N_19625);
and U20283 (N_20283,N_19510,N_19716);
and U20284 (N_20284,N_19875,N_19822);
xor U20285 (N_20285,N_19890,N_19841);
nand U20286 (N_20286,N_19561,N_19849);
or U20287 (N_20287,N_19617,N_19753);
and U20288 (N_20288,N_19793,N_19546);
and U20289 (N_20289,N_19668,N_19944);
nor U20290 (N_20290,N_19752,N_19889);
nand U20291 (N_20291,N_19592,N_19807);
and U20292 (N_20292,N_19868,N_19846);
and U20293 (N_20293,N_19519,N_19818);
nor U20294 (N_20294,N_19566,N_19558);
and U20295 (N_20295,N_19807,N_19801);
nor U20296 (N_20296,N_19590,N_19584);
nand U20297 (N_20297,N_19863,N_19942);
and U20298 (N_20298,N_19792,N_19982);
nand U20299 (N_20299,N_19656,N_19783);
nor U20300 (N_20300,N_19505,N_19534);
and U20301 (N_20301,N_19594,N_19502);
nand U20302 (N_20302,N_19848,N_19519);
or U20303 (N_20303,N_19882,N_19649);
xnor U20304 (N_20304,N_19737,N_19662);
nor U20305 (N_20305,N_19888,N_19731);
and U20306 (N_20306,N_19861,N_19841);
nor U20307 (N_20307,N_19941,N_19954);
xor U20308 (N_20308,N_19932,N_19885);
or U20309 (N_20309,N_19571,N_19865);
nand U20310 (N_20310,N_19632,N_19672);
nand U20311 (N_20311,N_19995,N_19710);
or U20312 (N_20312,N_19516,N_19564);
and U20313 (N_20313,N_19659,N_19949);
or U20314 (N_20314,N_19578,N_19624);
nand U20315 (N_20315,N_19742,N_19660);
nand U20316 (N_20316,N_19717,N_19560);
and U20317 (N_20317,N_19510,N_19968);
xor U20318 (N_20318,N_19776,N_19562);
nand U20319 (N_20319,N_19762,N_19784);
nor U20320 (N_20320,N_19712,N_19931);
and U20321 (N_20321,N_19796,N_19938);
and U20322 (N_20322,N_19639,N_19737);
xor U20323 (N_20323,N_19841,N_19522);
nor U20324 (N_20324,N_19725,N_19953);
xor U20325 (N_20325,N_19594,N_19806);
and U20326 (N_20326,N_19781,N_19987);
nor U20327 (N_20327,N_19868,N_19663);
nor U20328 (N_20328,N_19761,N_19519);
nor U20329 (N_20329,N_19796,N_19807);
and U20330 (N_20330,N_19695,N_19884);
or U20331 (N_20331,N_19501,N_19768);
nor U20332 (N_20332,N_19589,N_19747);
nand U20333 (N_20333,N_19530,N_19736);
nor U20334 (N_20334,N_19899,N_19715);
and U20335 (N_20335,N_19600,N_19750);
or U20336 (N_20336,N_19784,N_19853);
or U20337 (N_20337,N_19642,N_19547);
xnor U20338 (N_20338,N_19570,N_19894);
or U20339 (N_20339,N_19911,N_19796);
nand U20340 (N_20340,N_19717,N_19840);
or U20341 (N_20341,N_19991,N_19834);
or U20342 (N_20342,N_19586,N_19927);
xnor U20343 (N_20343,N_19960,N_19764);
and U20344 (N_20344,N_19863,N_19918);
and U20345 (N_20345,N_19741,N_19681);
nand U20346 (N_20346,N_19556,N_19813);
nor U20347 (N_20347,N_19683,N_19534);
xnor U20348 (N_20348,N_19523,N_19684);
or U20349 (N_20349,N_19879,N_19736);
xor U20350 (N_20350,N_19915,N_19535);
xnor U20351 (N_20351,N_19744,N_19749);
nand U20352 (N_20352,N_19682,N_19862);
or U20353 (N_20353,N_19959,N_19798);
nand U20354 (N_20354,N_19689,N_19663);
and U20355 (N_20355,N_19789,N_19864);
nand U20356 (N_20356,N_19580,N_19660);
nor U20357 (N_20357,N_19997,N_19773);
nor U20358 (N_20358,N_19807,N_19749);
xnor U20359 (N_20359,N_19934,N_19839);
or U20360 (N_20360,N_19973,N_19982);
nand U20361 (N_20361,N_19878,N_19670);
nor U20362 (N_20362,N_19634,N_19808);
or U20363 (N_20363,N_19551,N_19674);
nor U20364 (N_20364,N_19790,N_19988);
nor U20365 (N_20365,N_19709,N_19652);
and U20366 (N_20366,N_19580,N_19748);
nand U20367 (N_20367,N_19889,N_19939);
or U20368 (N_20368,N_19544,N_19585);
nor U20369 (N_20369,N_19727,N_19834);
or U20370 (N_20370,N_19652,N_19789);
nor U20371 (N_20371,N_19601,N_19627);
and U20372 (N_20372,N_19589,N_19710);
and U20373 (N_20373,N_19879,N_19812);
nor U20374 (N_20374,N_19917,N_19830);
xor U20375 (N_20375,N_19514,N_19899);
or U20376 (N_20376,N_19955,N_19833);
nand U20377 (N_20377,N_19511,N_19990);
or U20378 (N_20378,N_19795,N_19728);
nand U20379 (N_20379,N_19582,N_19599);
and U20380 (N_20380,N_19554,N_19680);
or U20381 (N_20381,N_19944,N_19755);
nand U20382 (N_20382,N_19563,N_19901);
and U20383 (N_20383,N_19588,N_19556);
or U20384 (N_20384,N_19738,N_19905);
nor U20385 (N_20385,N_19577,N_19808);
nand U20386 (N_20386,N_19738,N_19863);
and U20387 (N_20387,N_19612,N_19515);
and U20388 (N_20388,N_19643,N_19965);
and U20389 (N_20389,N_19514,N_19682);
and U20390 (N_20390,N_19521,N_19611);
nand U20391 (N_20391,N_19800,N_19564);
and U20392 (N_20392,N_19720,N_19556);
nand U20393 (N_20393,N_19654,N_19583);
or U20394 (N_20394,N_19704,N_19521);
nor U20395 (N_20395,N_19777,N_19615);
nor U20396 (N_20396,N_19751,N_19663);
or U20397 (N_20397,N_19935,N_19625);
nor U20398 (N_20398,N_19519,N_19922);
and U20399 (N_20399,N_19516,N_19999);
or U20400 (N_20400,N_19613,N_19985);
nand U20401 (N_20401,N_19692,N_19852);
nor U20402 (N_20402,N_19504,N_19814);
nor U20403 (N_20403,N_19636,N_19520);
nor U20404 (N_20404,N_19548,N_19976);
and U20405 (N_20405,N_19596,N_19677);
and U20406 (N_20406,N_19558,N_19915);
or U20407 (N_20407,N_19691,N_19978);
and U20408 (N_20408,N_19580,N_19516);
nor U20409 (N_20409,N_19640,N_19733);
nand U20410 (N_20410,N_19903,N_19752);
or U20411 (N_20411,N_19896,N_19718);
or U20412 (N_20412,N_19898,N_19821);
and U20413 (N_20413,N_19882,N_19635);
and U20414 (N_20414,N_19971,N_19922);
or U20415 (N_20415,N_19958,N_19789);
and U20416 (N_20416,N_19844,N_19705);
xnor U20417 (N_20417,N_19724,N_19606);
or U20418 (N_20418,N_19970,N_19589);
xor U20419 (N_20419,N_19578,N_19949);
and U20420 (N_20420,N_19732,N_19871);
xor U20421 (N_20421,N_19519,N_19752);
or U20422 (N_20422,N_19897,N_19706);
or U20423 (N_20423,N_19792,N_19517);
nor U20424 (N_20424,N_19586,N_19928);
and U20425 (N_20425,N_19706,N_19774);
or U20426 (N_20426,N_19888,N_19653);
nor U20427 (N_20427,N_19677,N_19790);
nand U20428 (N_20428,N_19591,N_19851);
nor U20429 (N_20429,N_19750,N_19624);
and U20430 (N_20430,N_19540,N_19850);
or U20431 (N_20431,N_19980,N_19787);
nand U20432 (N_20432,N_19662,N_19505);
or U20433 (N_20433,N_19851,N_19988);
nand U20434 (N_20434,N_19990,N_19580);
nand U20435 (N_20435,N_19541,N_19574);
and U20436 (N_20436,N_19953,N_19502);
nand U20437 (N_20437,N_19979,N_19573);
xor U20438 (N_20438,N_19770,N_19937);
and U20439 (N_20439,N_19851,N_19519);
and U20440 (N_20440,N_19763,N_19745);
nand U20441 (N_20441,N_19962,N_19740);
or U20442 (N_20442,N_19979,N_19810);
nor U20443 (N_20443,N_19799,N_19687);
and U20444 (N_20444,N_19785,N_19885);
and U20445 (N_20445,N_19935,N_19825);
nand U20446 (N_20446,N_19880,N_19538);
nand U20447 (N_20447,N_19780,N_19929);
nor U20448 (N_20448,N_19880,N_19559);
nand U20449 (N_20449,N_19547,N_19533);
nand U20450 (N_20450,N_19993,N_19561);
and U20451 (N_20451,N_19557,N_19833);
nand U20452 (N_20452,N_19501,N_19697);
nand U20453 (N_20453,N_19786,N_19997);
or U20454 (N_20454,N_19690,N_19597);
or U20455 (N_20455,N_19935,N_19963);
and U20456 (N_20456,N_19652,N_19901);
nor U20457 (N_20457,N_19984,N_19950);
xor U20458 (N_20458,N_19872,N_19511);
and U20459 (N_20459,N_19986,N_19746);
and U20460 (N_20460,N_19591,N_19688);
xnor U20461 (N_20461,N_19639,N_19945);
and U20462 (N_20462,N_19910,N_19558);
nor U20463 (N_20463,N_19795,N_19842);
and U20464 (N_20464,N_19606,N_19608);
xor U20465 (N_20465,N_19718,N_19950);
nor U20466 (N_20466,N_19929,N_19937);
or U20467 (N_20467,N_19805,N_19826);
xnor U20468 (N_20468,N_19767,N_19574);
or U20469 (N_20469,N_19572,N_19903);
and U20470 (N_20470,N_19721,N_19577);
nor U20471 (N_20471,N_19568,N_19720);
or U20472 (N_20472,N_19929,N_19913);
nand U20473 (N_20473,N_19915,N_19669);
nand U20474 (N_20474,N_19991,N_19988);
nand U20475 (N_20475,N_19600,N_19911);
or U20476 (N_20476,N_19786,N_19891);
nand U20477 (N_20477,N_19590,N_19808);
nor U20478 (N_20478,N_19893,N_19736);
or U20479 (N_20479,N_19675,N_19844);
or U20480 (N_20480,N_19657,N_19628);
and U20481 (N_20481,N_19776,N_19538);
and U20482 (N_20482,N_19608,N_19554);
and U20483 (N_20483,N_19653,N_19793);
and U20484 (N_20484,N_19764,N_19988);
xor U20485 (N_20485,N_19638,N_19846);
or U20486 (N_20486,N_19516,N_19638);
nor U20487 (N_20487,N_19890,N_19792);
xnor U20488 (N_20488,N_19728,N_19781);
or U20489 (N_20489,N_19893,N_19634);
nor U20490 (N_20490,N_19832,N_19519);
or U20491 (N_20491,N_19536,N_19740);
nor U20492 (N_20492,N_19938,N_19675);
or U20493 (N_20493,N_19782,N_19684);
and U20494 (N_20494,N_19568,N_19644);
nor U20495 (N_20495,N_19884,N_19641);
nor U20496 (N_20496,N_19990,N_19933);
nand U20497 (N_20497,N_19525,N_19674);
and U20498 (N_20498,N_19835,N_19577);
and U20499 (N_20499,N_19508,N_19605);
and U20500 (N_20500,N_20428,N_20069);
nor U20501 (N_20501,N_20418,N_20484);
nand U20502 (N_20502,N_20376,N_20413);
and U20503 (N_20503,N_20127,N_20393);
xor U20504 (N_20504,N_20173,N_20474);
or U20505 (N_20505,N_20449,N_20200);
nand U20506 (N_20506,N_20171,N_20036);
and U20507 (N_20507,N_20190,N_20311);
or U20508 (N_20508,N_20280,N_20232);
nand U20509 (N_20509,N_20142,N_20361);
nand U20510 (N_20510,N_20080,N_20191);
and U20511 (N_20511,N_20192,N_20250);
xor U20512 (N_20512,N_20004,N_20068);
nor U20513 (N_20513,N_20446,N_20128);
nor U20514 (N_20514,N_20107,N_20156);
nor U20515 (N_20515,N_20424,N_20022);
nor U20516 (N_20516,N_20199,N_20015);
or U20517 (N_20517,N_20287,N_20329);
xnor U20518 (N_20518,N_20347,N_20243);
or U20519 (N_20519,N_20365,N_20468);
nand U20520 (N_20520,N_20388,N_20444);
nand U20521 (N_20521,N_20319,N_20000);
or U20522 (N_20522,N_20220,N_20315);
or U20523 (N_20523,N_20033,N_20497);
xor U20524 (N_20524,N_20088,N_20348);
nor U20525 (N_20525,N_20317,N_20202);
nand U20526 (N_20526,N_20102,N_20229);
nor U20527 (N_20527,N_20327,N_20059);
nor U20528 (N_20528,N_20414,N_20115);
nand U20529 (N_20529,N_20155,N_20164);
and U20530 (N_20530,N_20270,N_20344);
or U20531 (N_20531,N_20209,N_20025);
nor U20532 (N_20532,N_20321,N_20300);
xnor U20533 (N_20533,N_20216,N_20111);
xnor U20534 (N_20534,N_20046,N_20044);
xnor U20535 (N_20535,N_20104,N_20244);
xor U20536 (N_20536,N_20053,N_20378);
xnor U20537 (N_20537,N_20212,N_20379);
xor U20538 (N_20538,N_20441,N_20362);
nor U20539 (N_20539,N_20149,N_20399);
or U20540 (N_20540,N_20482,N_20346);
and U20541 (N_20541,N_20373,N_20066);
nand U20542 (N_20542,N_20029,N_20358);
xnor U20543 (N_20543,N_20041,N_20175);
nand U20544 (N_20544,N_20451,N_20279);
and U20545 (N_20545,N_20230,N_20206);
nand U20546 (N_20546,N_20406,N_20481);
nand U20547 (N_20547,N_20296,N_20304);
xnor U20548 (N_20548,N_20057,N_20081);
or U20549 (N_20549,N_20110,N_20272);
xor U20550 (N_20550,N_20407,N_20288);
xor U20551 (N_20551,N_20219,N_20040);
nor U20552 (N_20552,N_20387,N_20178);
nor U20553 (N_20553,N_20062,N_20457);
xor U20554 (N_20554,N_20345,N_20383);
and U20555 (N_20555,N_20491,N_20495);
nor U20556 (N_20556,N_20089,N_20119);
nand U20557 (N_20557,N_20332,N_20403);
nand U20558 (N_20558,N_20204,N_20284);
and U20559 (N_20559,N_20218,N_20483);
nand U20560 (N_20560,N_20231,N_20008);
nand U20561 (N_20561,N_20355,N_20283);
or U20562 (N_20562,N_20374,N_20034);
or U20563 (N_20563,N_20225,N_20159);
or U20564 (N_20564,N_20236,N_20063);
nand U20565 (N_20565,N_20124,N_20245);
and U20566 (N_20566,N_20078,N_20120);
and U20567 (N_20567,N_20443,N_20012);
and U20568 (N_20568,N_20181,N_20179);
nand U20569 (N_20569,N_20459,N_20145);
and U20570 (N_20570,N_20343,N_20445);
and U20571 (N_20571,N_20377,N_20135);
or U20572 (N_20572,N_20334,N_20342);
and U20573 (N_20573,N_20290,N_20152);
nand U20574 (N_20574,N_20055,N_20177);
nor U20575 (N_20575,N_20341,N_20167);
nor U20576 (N_20576,N_20038,N_20065);
and U20577 (N_20577,N_20282,N_20086);
and U20578 (N_20578,N_20480,N_20305);
nand U20579 (N_20579,N_20401,N_20289);
nor U20580 (N_20580,N_20411,N_20281);
or U20581 (N_20581,N_20356,N_20415);
nand U20582 (N_20582,N_20074,N_20479);
or U20583 (N_20583,N_20137,N_20467);
nor U20584 (N_20584,N_20370,N_20096);
nor U20585 (N_20585,N_20163,N_20189);
nor U20586 (N_20586,N_20248,N_20368);
nor U20587 (N_20587,N_20075,N_20409);
nand U20588 (N_20588,N_20326,N_20151);
and U20589 (N_20589,N_20252,N_20242);
nor U20590 (N_20590,N_20490,N_20486);
nor U20591 (N_20591,N_20260,N_20228);
or U20592 (N_20592,N_20306,N_20113);
and U20593 (N_20593,N_20032,N_20150);
or U20594 (N_20594,N_20463,N_20211);
or U20595 (N_20595,N_20275,N_20003);
nor U20596 (N_20596,N_20299,N_20043);
or U20597 (N_20597,N_20349,N_20052);
or U20598 (N_20598,N_20324,N_20234);
nand U20599 (N_20599,N_20313,N_20099);
nand U20600 (N_20600,N_20256,N_20352);
nor U20601 (N_20601,N_20011,N_20391);
nand U20602 (N_20602,N_20237,N_20440);
nand U20603 (N_20603,N_20070,N_20169);
nor U20604 (N_20604,N_20475,N_20316);
nor U20605 (N_20605,N_20117,N_20223);
and U20606 (N_20606,N_20339,N_20442);
nand U20607 (N_20607,N_20277,N_20461);
and U20608 (N_20608,N_20372,N_20337);
or U20609 (N_20609,N_20360,N_20121);
nor U20610 (N_20610,N_20194,N_20101);
and U20611 (N_20611,N_20002,N_20071);
or U20612 (N_20612,N_20083,N_20477);
xor U20613 (N_20613,N_20438,N_20076);
nand U20614 (N_20614,N_20450,N_20494);
nand U20615 (N_20615,N_20359,N_20241);
and U20616 (N_20616,N_20161,N_20126);
xnor U20617 (N_20617,N_20251,N_20437);
and U20618 (N_20618,N_20257,N_20464);
xnor U20619 (N_20619,N_20073,N_20478);
xnor U20620 (N_20620,N_20402,N_20026);
nand U20621 (N_20621,N_20143,N_20364);
or U20622 (N_20622,N_20196,N_20049);
or U20623 (N_20623,N_20447,N_20350);
nor U20624 (N_20624,N_20172,N_20154);
and U20625 (N_20625,N_20489,N_20278);
nor U20626 (N_20626,N_20238,N_20139);
nand U20627 (N_20627,N_20087,N_20453);
and U20628 (N_20628,N_20462,N_20427);
xnor U20629 (N_20629,N_20213,N_20006);
or U20630 (N_20630,N_20499,N_20405);
or U20631 (N_20631,N_20235,N_20056);
and U20632 (N_20632,N_20146,N_20476);
or U20633 (N_20633,N_20058,N_20331);
or U20634 (N_20634,N_20203,N_20129);
nand U20635 (N_20635,N_20157,N_20488);
and U20636 (N_20636,N_20123,N_20197);
and U20637 (N_20637,N_20125,N_20103);
nor U20638 (N_20638,N_20013,N_20431);
xnor U20639 (N_20639,N_20395,N_20408);
nor U20640 (N_20640,N_20091,N_20430);
nand U20641 (N_20641,N_20318,N_20295);
nor U20642 (N_20642,N_20353,N_20381);
nor U20643 (N_20643,N_20335,N_20136);
nor U20644 (N_20644,N_20094,N_20466);
nand U20645 (N_20645,N_20274,N_20118);
nand U20646 (N_20646,N_20470,N_20493);
nand U20647 (N_20647,N_20116,N_20310);
or U20648 (N_20648,N_20487,N_20222);
nor U20649 (N_20649,N_20404,N_20498);
nor U20650 (N_20650,N_20144,N_20357);
nand U20651 (N_20651,N_20389,N_20269);
xor U20652 (N_20652,N_20018,N_20434);
nand U20653 (N_20653,N_20254,N_20323);
nor U20654 (N_20654,N_20185,N_20108);
nor U20655 (N_20655,N_20294,N_20007);
nand U20656 (N_20656,N_20338,N_20291);
nor U20657 (N_20657,N_20182,N_20233);
or U20658 (N_20658,N_20336,N_20208);
and U20659 (N_20659,N_20239,N_20024);
nor U20660 (N_20660,N_20227,N_20133);
or U20661 (N_20661,N_20258,N_20263);
nand U20662 (N_20662,N_20425,N_20385);
nor U20663 (N_20663,N_20226,N_20363);
or U20664 (N_20664,N_20456,N_20485);
and U20665 (N_20665,N_20293,N_20448);
or U20666 (N_20666,N_20308,N_20077);
and U20667 (N_20667,N_20384,N_20469);
nand U20668 (N_20668,N_20421,N_20247);
or U20669 (N_20669,N_20097,N_20367);
nand U20670 (N_20670,N_20390,N_20035);
nor U20671 (N_20671,N_20435,N_20009);
or U20672 (N_20672,N_20106,N_20286);
nor U20673 (N_20673,N_20410,N_20165);
nand U20674 (N_20674,N_20186,N_20166);
nand U20675 (N_20675,N_20187,N_20392);
nor U20676 (N_20676,N_20039,N_20354);
and U20677 (N_20677,N_20174,N_20031);
or U20678 (N_20678,N_20100,N_20303);
or U20679 (N_20679,N_20264,N_20412);
xor U20680 (N_20680,N_20021,N_20224);
or U20681 (N_20681,N_20047,N_20153);
xnor U20682 (N_20682,N_20105,N_20134);
nor U20683 (N_20683,N_20176,N_20325);
nand U20684 (N_20684,N_20168,N_20394);
nand U20685 (N_20685,N_20017,N_20312);
and U20686 (N_20686,N_20201,N_20267);
or U20687 (N_20687,N_20268,N_20060);
nor U20688 (N_20688,N_20465,N_20210);
nand U20689 (N_20689,N_20050,N_20183);
and U20690 (N_20690,N_20330,N_20417);
or U20691 (N_20691,N_20439,N_20375);
and U20692 (N_20692,N_20188,N_20042);
nor U20693 (N_20693,N_20432,N_20386);
nand U20694 (N_20694,N_20028,N_20147);
and U20695 (N_20695,N_20221,N_20051);
nand U20696 (N_20696,N_20048,N_20214);
nor U20697 (N_20697,N_20265,N_20285);
or U20698 (N_20698,N_20473,N_20093);
or U20699 (N_20699,N_20320,N_20001);
or U20700 (N_20700,N_20422,N_20369);
xnor U20701 (N_20701,N_20130,N_20416);
or U20702 (N_20702,N_20140,N_20030);
and U20703 (N_20703,N_20458,N_20122);
xnor U20704 (N_20704,N_20433,N_20061);
nor U20705 (N_20705,N_20072,N_20396);
and U20706 (N_20706,N_20454,N_20255);
or U20707 (N_20707,N_20382,N_20020);
nor U20708 (N_20708,N_20198,N_20085);
nor U20709 (N_20709,N_20114,N_20095);
nand U20710 (N_20710,N_20132,N_20092);
nor U20711 (N_20711,N_20351,N_20160);
or U20712 (N_20712,N_20309,N_20240);
or U20713 (N_20713,N_20082,N_20207);
nor U20714 (N_20714,N_20302,N_20141);
or U20715 (N_20715,N_20067,N_20027);
nand U20716 (N_20716,N_20215,N_20333);
or U20717 (N_20717,N_20398,N_20301);
xor U20718 (N_20718,N_20064,N_20148);
nor U20719 (N_20719,N_20246,N_20259);
xor U20720 (N_20720,N_20340,N_20322);
nor U20721 (N_20721,N_20426,N_20005);
nand U20722 (N_20722,N_20423,N_20184);
and U20723 (N_20723,N_20471,N_20271);
nor U20724 (N_20724,N_20162,N_20037);
nor U20725 (N_20725,N_20366,N_20014);
or U20726 (N_20726,N_20380,N_20455);
nand U20727 (N_20727,N_20109,N_20266);
nand U20728 (N_20728,N_20079,N_20016);
nor U20729 (N_20729,N_20193,N_20131);
nand U20730 (N_20730,N_20496,N_20276);
nand U20731 (N_20731,N_20371,N_20420);
and U20732 (N_20732,N_20297,N_20217);
and U20733 (N_20733,N_20253,N_20195);
nand U20734 (N_20734,N_20472,N_20419);
nor U20735 (N_20735,N_20262,N_20010);
xor U20736 (N_20736,N_20180,N_20273);
or U20737 (N_20737,N_20170,N_20328);
and U20738 (N_20738,N_20261,N_20054);
nand U20739 (N_20739,N_20158,N_20460);
nor U20740 (N_20740,N_20023,N_20307);
xnor U20741 (N_20741,N_20292,N_20452);
nor U20742 (N_20742,N_20045,N_20429);
nand U20743 (N_20743,N_20098,N_20138);
or U20744 (N_20744,N_20112,N_20397);
and U20745 (N_20745,N_20205,N_20492);
nor U20746 (N_20746,N_20084,N_20019);
nor U20747 (N_20747,N_20436,N_20298);
nand U20748 (N_20748,N_20249,N_20314);
or U20749 (N_20749,N_20090,N_20400);
and U20750 (N_20750,N_20380,N_20199);
and U20751 (N_20751,N_20289,N_20383);
nor U20752 (N_20752,N_20031,N_20200);
nand U20753 (N_20753,N_20021,N_20451);
or U20754 (N_20754,N_20443,N_20106);
xnor U20755 (N_20755,N_20400,N_20158);
nor U20756 (N_20756,N_20351,N_20476);
or U20757 (N_20757,N_20363,N_20046);
xor U20758 (N_20758,N_20385,N_20345);
or U20759 (N_20759,N_20243,N_20264);
xnor U20760 (N_20760,N_20171,N_20471);
or U20761 (N_20761,N_20006,N_20394);
nand U20762 (N_20762,N_20495,N_20254);
and U20763 (N_20763,N_20342,N_20029);
or U20764 (N_20764,N_20061,N_20263);
and U20765 (N_20765,N_20021,N_20435);
or U20766 (N_20766,N_20200,N_20157);
and U20767 (N_20767,N_20432,N_20466);
or U20768 (N_20768,N_20282,N_20446);
or U20769 (N_20769,N_20314,N_20118);
xnor U20770 (N_20770,N_20219,N_20353);
or U20771 (N_20771,N_20415,N_20037);
nand U20772 (N_20772,N_20240,N_20445);
and U20773 (N_20773,N_20473,N_20213);
and U20774 (N_20774,N_20179,N_20169);
nor U20775 (N_20775,N_20046,N_20162);
or U20776 (N_20776,N_20336,N_20454);
or U20777 (N_20777,N_20144,N_20269);
or U20778 (N_20778,N_20189,N_20096);
nor U20779 (N_20779,N_20115,N_20040);
nand U20780 (N_20780,N_20206,N_20470);
and U20781 (N_20781,N_20158,N_20363);
or U20782 (N_20782,N_20370,N_20453);
nand U20783 (N_20783,N_20455,N_20247);
nand U20784 (N_20784,N_20443,N_20000);
nor U20785 (N_20785,N_20358,N_20164);
xnor U20786 (N_20786,N_20292,N_20042);
xnor U20787 (N_20787,N_20204,N_20122);
xnor U20788 (N_20788,N_20431,N_20363);
nand U20789 (N_20789,N_20047,N_20460);
nand U20790 (N_20790,N_20450,N_20376);
nor U20791 (N_20791,N_20276,N_20123);
or U20792 (N_20792,N_20476,N_20280);
and U20793 (N_20793,N_20215,N_20337);
nor U20794 (N_20794,N_20044,N_20479);
xnor U20795 (N_20795,N_20220,N_20205);
nand U20796 (N_20796,N_20049,N_20019);
and U20797 (N_20797,N_20108,N_20284);
or U20798 (N_20798,N_20181,N_20285);
nand U20799 (N_20799,N_20452,N_20088);
nand U20800 (N_20800,N_20394,N_20319);
xor U20801 (N_20801,N_20186,N_20376);
or U20802 (N_20802,N_20470,N_20145);
or U20803 (N_20803,N_20464,N_20417);
nand U20804 (N_20804,N_20280,N_20099);
and U20805 (N_20805,N_20324,N_20487);
nor U20806 (N_20806,N_20142,N_20228);
and U20807 (N_20807,N_20168,N_20274);
and U20808 (N_20808,N_20475,N_20026);
and U20809 (N_20809,N_20303,N_20048);
nor U20810 (N_20810,N_20097,N_20217);
or U20811 (N_20811,N_20087,N_20163);
and U20812 (N_20812,N_20166,N_20366);
nand U20813 (N_20813,N_20250,N_20215);
nor U20814 (N_20814,N_20462,N_20449);
nor U20815 (N_20815,N_20289,N_20328);
or U20816 (N_20816,N_20372,N_20251);
or U20817 (N_20817,N_20298,N_20462);
or U20818 (N_20818,N_20207,N_20210);
and U20819 (N_20819,N_20008,N_20160);
nand U20820 (N_20820,N_20416,N_20021);
nand U20821 (N_20821,N_20499,N_20221);
nand U20822 (N_20822,N_20202,N_20284);
and U20823 (N_20823,N_20473,N_20376);
xnor U20824 (N_20824,N_20362,N_20395);
and U20825 (N_20825,N_20386,N_20036);
and U20826 (N_20826,N_20410,N_20043);
nand U20827 (N_20827,N_20257,N_20301);
or U20828 (N_20828,N_20219,N_20420);
or U20829 (N_20829,N_20116,N_20032);
or U20830 (N_20830,N_20379,N_20106);
or U20831 (N_20831,N_20170,N_20157);
or U20832 (N_20832,N_20060,N_20334);
or U20833 (N_20833,N_20314,N_20289);
and U20834 (N_20834,N_20387,N_20184);
xor U20835 (N_20835,N_20251,N_20309);
and U20836 (N_20836,N_20251,N_20375);
nand U20837 (N_20837,N_20405,N_20009);
nor U20838 (N_20838,N_20292,N_20038);
and U20839 (N_20839,N_20173,N_20080);
nor U20840 (N_20840,N_20001,N_20069);
xnor U20841 (N_20841,N_20484,N_20072);
xor U20842 (N_20842,N_20372,N_20098);
nand U20843 (N_20843,N_20450,N_20196);
nor U20844 (N_20844,N_20135,N_20020);
or U20845 (N_20845,N_20315,N_20181);
and U20846 (N_20846,N_20292,N_20291);
nor U20847 (N_20847,N_20377,N_20454);
and U20848 (N_20848,N_20246,N_20127);
nand U20849 (N_20849,N_20117,N_20172);
xor U20850 (N_20850,N_20241,N_20440);
and U20851 (N_20851,N_20044,N_20164);
nand U20852 (N_20852,N_20004,N_20019);
or U20853 (N_20853,N_20228,N_20378);
nor U20854 (N_20854,N_20188,N_20438);
nand U20855 (N_20855,N_20003,N_20010);
nand U20856 (N_20856,N_20213,N_20036);
nand U20857 (N_20857,N_20487,N_20216);
xor U20858 (N_20858,N_20170,N_20228);
and U20859 (N_20859,N_20281,N_20485);
nand U20860 (N_20860,N_20400,N_20419);
nor U20861 (N_20861,N_20309,N_20426);
nand U20862 (N_20862,N_20330,N_20123);
nor U20863 (N_20863,N_20187,N_20390);
and U20864 (N_20864,N_20027,N_20437);
nand U20865 (N_20865,N_20067,N_20473);
or U20866 (N_20866,N_20445,N_20114);
and U20867 (N_20867,N_20271,N_20156);
nor U20868 (N_20868,N_20208,N_20100);
and U20869 (N_20869,N_20368,N_20037);
nand U20870 (N_20870,N_20471,N_20129);
and U20871 (N_20871,N_20463,N_20023);
and U20872 (N_20872,N_20099,N_20408);
and U20873 (N_20873,N_20239,N_20020);
nand U20874 (N_20874,N_20461,N_20149);
or U20875 (N_20875,N_20139,N_20297);
xnor U20876 (N_20876,N_20496,N_20010);
xnor U20877 (N_20877,N_20438,N_20295);
nand U20878 (N_20878,N_20306,N_20336);
and U20879 (N_20879,N_20088,N_20193);
xnor U20880 (N_20880,N_20386,N_20159);
and U20881 (N_20881,N_20398,N_20431);
and U20882 (N_20882,N_20228,N_20432);
or U20883 (N_20883,N_20265,N_20089);
or U20884 (N_20884,N_20412,N_20055);
nand U20885 (N_20885,N_20338,N_20250);
nor U20886 (N_20886,N_20311,N_20392);
nand U20887 (N_20887,N_20168,N_20496);
or U20888 (N_20888,N_20364,N_20000);
and U20889 (N_20889,N_20089,N_20470);
nand U20890 (N_20890,N_20190,N_20109);
nor U20891 (N_20891,N_20496,N_20242);
nor U20892 (N_20892,N_20379,N_20322);
and U20893 (N_20893,N_20189,N_20059);
xor U20894 (N_20894,N_20092,N_20072);
and U20895 (N_20895,N_20260,N_20361);
and U20896 (N_20896,N_20302,N_20289);
xor U20897 (N_20897,N_20298,N_20067);
or U20898 (N_20898,N_20446,N_20457);
and U20899 (N_20899,N_20101,N_20442);
xnor U20900 (N_20900,N_20449,N_20081);
nand U20901 (N_20901,N_20088,N_20278);
nand U20902 (N_20902,N_20100,N_20489);
and U20903 (N_20903,N_20097,N_20401);
xor U20904 (N_20904,N_20169,N_20333);
or U20905 (N_20905,N_20493,N_20080);
nor U20906 (N_20906,N_20174,N_20125);
nor U20907 (N_20907,N_20192,N_20263);
or U20908 (N_20908,N_20325,N_20380);
nor U20909 (N_20909,N_20488,N_20209);
or U20910 (N_20910,N_20162,N_20369);
and U20911 (N_20911,N_20225,N_20215);
nand U20912 (N_20912,N_20031,N_20215);
xor U20913 (N_20913,N_20419,N_20438);
and U20914 (N_20914,N_20088,N_20221);
nor U20915 (N_20915,N_20048,N_20039);
or U20916 (N_20916,N_20224,N_20421);
nand U20917 (N_20917,N_20158,N_20125);
or U20918 (N_20918,N_20265,N_20185);
or U20919 (N_20919,N_20284,N_20188);
or U20920 (N_20920,N_20179,N_20459);
and U20921 (N_20921,N_20035,N_20467);
nand U20922 (N_20922,N_20375,N_20358);
or U20923 (N_20923,N_20486,N_20104);
nand U20924 (N_20924,N_20157,N_20299);
xnor U20925 (N_20925,N_20325,N_20191);
or U20926 (N_20926,N_20385,N_20200);
and U20927 (N_20927,N_20124,N_20465);
nor U20928 (N_20928,N_20332,N_20115);
nand U20929 (N_20929,N_20108,N_20449);
nand U20930 (N_20930,N_20171,N_20152);
xor U20931 (N_20931,N_20149,N_20360);
and U20932 (N_20932,N_20373,N_20393);
and U20933 (N_20933,N_20101,N_20360);
and U20934 (N_20934,N_20271,N_20097);
nor U20935 (N_20935,N_20192,N_20308);
or U20936 (N_20936,N_20162,N_20273);
nand U20937 (N_20937,N_20054,N_20424);
and U20938 (N_20938,N_20257,N_20243);
xnor U20939 (N_20939,N_20409,N_20296);
nand U20940 (N_20940,N_20358,N_20269);
nand U20941 (N_20941,N_20337,N_20112);
or U20942 (N_20942,N_20387,N_20279);
or U20943 (N_20943,N_20193,N_20475);
nor U20944 (N_20944,N_20461,N_20105);
nor U20945 (N_20945,N_20300,N_20465);
or U20946 (N_20946,N_20055,N_20146);
nor U20947 (N_20947,N_20165,N_20324);
nand U20948 (N_20948,N_20286,N_20479);
and U20949 (N_20949,N_20312,N_20142);
xor U20950 (N_20950,N_20241,N_20064);
xor U20951 (N_20951,N_20070,N_20182);
nor U20952 (N_20952,N_20317,N_20384);
or U20953 (N_20953,N_20233,N_20378);
and U20954 (N_20954,N_20467,N_20358);
xor U20955 (N_20955,N_20482,N_20383);
and U20956 (N_20956,N_20247,N_20456);
nor U20957 (N_20957,N_20034,N_20444);
and U20958 (N_20958,N_20415,N_20314);
or U20959 (N_20959,N_20498,N_20109);
or U20960 (N_20960,N_20498,N_20452);
xor U20961 (N_20961,N_20021,N_20385);
nor U20962 (N_20962,N_20328,N_20390);
and U20963 (N_20963,N_20292,N_20108);
and U20964 (N_20964,N_20086,N_20062);
xnor U20965 (N_20965,N_20169,N_20085);
or U20966 (N_20966,N_20245,N_20469);
and U20967 (N_20967,N_20047,N_20099);
or U20968 (N_20968,N_20094,N_20044);
nand U20969 (N_20969,N_20031,N_20196);
xor U20970 (N_20970,N_20393,N_20033);
and U20971 (N_20971,N_20298,N_20005);
nand U20972 (N_20972,N_20424,N_20130);
and U20973 (N_20973,N_20232,N_20265);
nand U20974 (N_20974,N_20141,N_20089);
or U20975 (N_20975,N_20262,N_20216);
nor U20976 (N_20976,N_20149,N_20346);
nor U20977 (N_20977,N_20490,N_20492);
or U20978 (N_20978,N_20030,N_20159);
or U20979 (N_20979,N_20187,N_20453);
and U20980 (N_20980,N_20076,N_20486);
nor U20981 (N_20981,N_20476,N_20392);
nor U20982 (N_20982,N_20216,N_20255);
xnor U20983 (N_20983,N_20343,N_20136);
xor U20984 (N_20984,N_20402,N_20002);
nor U20985 (N_20985,N_20139,N_20398);
or U20986 (N_20986,N_20031,N_20177);
nand U20987 (N_20987,N_20417,N_20118);
and U20988 (N_20988,N_20409,N_20381);
nor U20989 (N_20989,N_20078,N_20382);
nand U20990 (N_20990,N_20422,N_20207);
nand U20991 (N_20991,N_20253,N_20100);
nor U20992 (N_20992,N_20021,N_20069);
or U20993 (N_20993,N_20459,N_20398);
or U20994 (N_20994,N_20394,N_20380);
nor U20995 (N_20995,N_20425,N_20218);
or U20996 (N_20996,N_20024,N_20281);
or U20997 (N_20997,N_20381,N_20302);
and U20998 (N_20998,N_20094,N_20013);
nor U20999 (N_20999,N_20310,N_20396);
nor U21000 (N_21000,N_20761,N_20844);
and U21001 (N_21001,N_20720,N_20803);
and U21002 (N_21002,N_20617,N_20830);
or U21003 (N_21003,N_20620,N_20807);
nor U21004 (N_21004,N_20582,N_20922);
and U21005 (N_21005,N_20762,N_20929);
and U21006 (N_21006,N_20948,N_20590);
nor U21007 (N_21007,N_20504,N_20687);
nand U21008 (N_21008,N_20974,N_20505);
or U21009 (N_21009,N_20667,N_20961);
or U21010 (N_21010,N_20842,N_20580);
and U21011 (N_21011,N_20649,N_20541);
nand U21012 (N_21012,N_20622,N_20771);
nand U21013 (N_21013,N_20852,N_20659);
nand U21014 (N_21014,N_20584,N_20663);
or U21015 (N_21015,N_20797,N_20875);
or U21016 (N_21016,N_20958,N_20769);
xnor U21017 (N_21017,N_20655,N_20650);
nor U21018 (N_21018,N_20833,N_20967);
nor U21019 (N_21019,N_20630,N_20774);
or U21020 (N_21020,N_20568,N_20999);
nor U21021 (N_21021,N_20828,N_20837);
and U21022 (N_21022,N_20968,N_20749);
nor U21023 (N_21023,N_20506,N_20735);
and U21024 (N_21024,N_20954,N_20933);
nand U21025 (N_21025,N_20819,N_20514);
xnor U21026 (N_21026,N_20795,N_20942);
or U21027 (N_21027,N_20754,N_20614);
and U21028 (N_21028,N_20581,N_20500);
and U21029 (N_21029,N_20938,N_20935);
nor U21030 (N_21030,N_20585,N_20544);
xnor U21031 (N_21031,N_20755,N_20882);
nor U21032 (N_21032,N_20678,N_20546);
nand U21033 (N_21033,N_20950,N_20986);
nand U21034 (N_21034,N_20936,N_20587);
and U21035 (N_21035,N_20731,N_20664);
nand U21036 (N_21036,N_20710,N_20751);
nand U21037 (N_21037,N_20524,N_20870);
nand U21038 (N_21038,N_20530,N_20701);
or U21039 (N_21039,N_20560,N_20536);
and U21040 (N_21040,N_20717,N_20684);
nand U21041 (N_21041,N_20539,N_20892);
and U21042 (N_21042,N_20962,N_20734);
xnor U21043 (N_21043,N_20733,N_20704);
xor U21044 (N_21044,N_20848,N_20785);
and U21045 (N_21045,N_20865,N_20522);
or U21046 (N_21046,N_20854,N_20953);
nor U21047 (N_21047,N_20592,N_20910);
nor U21048 (N_21048,N_20977,N_20941);
nor U21049 (N_21049,N_20610,N_20995);
and U21050 (N_21050,N_20537,N_20752);
nor U21051 (N_21051,N_20960,N_20681);
nor U21052 (N_21052,N_20728,N_20851);
nand U21053 (N_21053,N_20683,N_20697);
xor U21054 (N_21054,N_20674,N_20594);
nor U21055 (N_21055,N_20793,N_20786);
xnor U21056 (N_21056,N_20745,N_20725);
or U21057 (N_21057,N_20703,N_20934);
xnor U21058 (N_21058,N_20662,N_20850);
nor U21059 (N_21059,N_20689,N_20586);
nor U21060 (N_21060,N_20548,N_20742);
or U21061 (N_21061,N_20577,N_20509);
nor U21062 (N_21062,N_20966,N_20576);
nand U21063 (N_21063,N_20740,N_20949);
and U21064 (N_21064,N_20783,N_20897);
nand U21065 (N_21065,N_20644,N_20519);
nor U21066 (N_21066,N_20790,N_20713);
or U21067 (N_21067,N_20503,N_20721);
nand U21068 (N_21068,N_20893,N_20711);
nor U21069 (N_21069,N_20794,N_20920);
xnor U21070 (N_21070,N_20691,N_20832);
and U21071 (N_21071,N_20944,N_20562);
nor U21072 (N_21072,N_20824,N_20518);
and U21073 (N_21073,N_20887,N_20979);
and U21074 (N_21074,N_20903,N_20839);
xnor U21075 (N_21075,N_20998,N_20545);
xor U21076 (N_21076,N_20955,N_20779);
or U21077 (N_21077,N_20975,N_20706);
or U21078 (N_21078,N_20940,N_20712);
and U21079 (N_21079,N_20613,N_20528);
and U21080 (N_21080,N_20923,N_20772);
nor U21081 (N_21081,N_20906,N_20916);
nand U21082 (N_21082,N_20588,N_20931);
xnor U21083 (N_21083,N_20616,N_20700);
xnor U21084 (N_21084,N_20798,N_20909);
nand U21085 (N_21085,N_20991,N_20969);
and U21086 (N_21086,N_20727,N_20557);
nor U21087 (N_21087,N_20692,N_20778);
and U21088 (N_21088,N_20997,N_20859);
nand U21089 (N_21089,N_20781,N_20987);
nand U21090 (N_21090,N_20653,N_20829);
nor U21091 (N_21091,N_20627,N_20766);
nand U21092 (N_21092,N_20512,N_20973);
xor U21093 (N_21093,N_20787,N_20891);
or U21094 (N_21094,N_20855,N_20729);
nor U21095 (N_21095,N_20708,N_20812);
and U21096 (N_21096,N_20623,N_20993);
nand U21097 (N_21097,N_20589,N_20699);
or U21098 (N_21098,N_20531,N_20996);
or U21099 (N_21099,N_20715,N_20648);
nor U21100 (N_21100,N_20563,N_20640);
xnor U21101 (N_21101,N_20682,N_20804);
nand U21102 (N_21102,N_20972,N_20543);
or U21103 (N_21103,N_20513,N_20867);
and U21104 (N_21104,N_20707,N_20860);
or U21105 (N_21105,N_20881,N_20567);
nor U21106 (N_21106,N_20921,N_20809);
and U21107 (N_21107,N_20709,N_20880);
or U21108 (N_21108,N_20652,N_20789);
and U21109 (N_21109,N_20719,N_20843);
and U21110 (N_21110,N_20671,N_20877);
xnor U21111 (N_21111,N_20963,N_20680);
or U21112 (N_21112,N_20527,N_20750);
nand U21113 (N_21113,N_20773,N_20970);
or U21114 (N_21114,N_20716,N_20657);
and U21115 (N_21115,N_20964,N_20615);
nand U21116 (N_21116,N_20561,N_20796);
nor U21117 (N_21117,N_20775,N_20814);
nand U21118 (N_21118,N_20869,N_20912);
nor U21119 (N_21119,N_20510,N_20874);
and U21120 (N_21120,N_20813,N_20628);
and U21121 (N_21121,N_20672,N_20917);
nand U21122 (N_21122,N_20904,N_20746);
and U21123 (N_21123,N_20939,N_20930);
or U21124 (N_21124,N_20547,N_20722);
nor U21125 (N_21125,N_20937,N_20511);
or U21126 (N_21126,N_20611,N_20638);
nor U21127 (N_21127,N_20951,N_20591);
or U21128 (N_21128,N_20827,N_20694);
or U21129 (N_21129,N_20702,N_20911);
or U21130 (N_21130,N_20925,N_20756);
and U21131 (N_21131,N_20846,N_20575);
and U21132 (N_21132,N_20501,N_20744);
nor U21133 (N_21133,N_20943,N_20619);
or U21134 (N_21134,N_20924,N_20792);
nor U21135 (N_21135,N_20947,N_20758);
nand U21136 (N_21136,N_20805,N_20669);
nor U21137 (N_21137,N_20840,N_20820);
and U21138 (N_21138,N_20743,N_20621);
or U21139 (N_21139,N_20905,N_20811);
nand U21140 (N_21140,N_20926,N_20660);
or U21141 (N_21141,N_20757,N_20551);
nand U21142 (N_21142,N_20515,N_20836);
nand U21143 (N_21143,N_20686,N_20978);
nand U21144 (N_21144,N_20676,N_20873);
xor U21145 (N_21145,N_20888,N_20945);
or U21146 (N_21146,N_20864,N_20606);
xor U21147 (N_21147,N_20673,N_20521);
and U21148 (N_21148,N_20826,N_20693);
and U21149 (N_21149,N_20777,N_20520);
nor U21150 (N_21150,N_20635,N_20834);
nand U21151 (N_21151,N_20845,N_20738);
nor U21152 (N_21152,N_20508,N_20685);
nand U21153 (N_21153,N_20760,N_20858);
nor U21154 (N_21154,N_20884,N_20724);
nor U21155 (N_21155,N_20886,N_20876);
and U21156 (N_21156,N_20806,N_20553);
nand U21157 (N_21157,N_20989,N_20688);
or U21158 (N_21158,N_20889,N_20776);
nand U21159 (N_21159,N_20992,N_20643);
or U21160 (N_21160,N_20841,N_20646);
and U21161 (N_21161,N_20571,N_20965);
nand U21162 (N_21162,N_20639,N_20932);
nand U21163 (N_21163,N_20570,N_20516);
nor U21164 (N_21164,N_20782,N_20915);
nor U21165 (N_21165,N_20853,N_20647);
nand U21166 (N_21166,N_20668,N_20636);
xor U21167 (N_21167,N_20983,N_20868);
nand U21168 (N_21168,N_20698,N_20849);
or U21169 (N_21169,N_20651,N_20759);
or U21170 (N_21170,N_20677,N_20661);
and U21171 (N_21171,N_20894,N_20583);
nand U21172 (N_21172,N_20885,N_20573);
nand U21173 (N_21173,N_20872,N_20831);
or U21174 (N_21174,N_20624,N_20637);
nand U21175 (N_21175,N_20654,N_20791);
or U21176 (N_21176,N_20533,N_20718);
or U21177 (N_21177,N_20626,N_20695);
xnor U21178 (N_21178,N_20629,N_20632);
or U21179 (N_21179,N_20984,N_20602);
or U21180 (N_21180,N_20665,N_20780);
or U21181 (N_21181,N_20612,N_20770);
nand U21182 (N_21182,N_20784,N_20538);
or U21183 (N_21183,N_20641,N_20634);
nand U21184 (N_21184,N_20818,N_20607);
xnor U21185 (N_21185,N_20788,N_20866);
and U21186 (N_21186,N_20666,N_20633);
and U21187 (N_21187,N_20604,N_20631);
and U21188 (N_21188,N_20994,N_20861);
nand U21189 (N_21189,N_20747,N_20670);
nand U21190 (N_21190,N_20625,N_20908);
nand U21191 (N_21191,N_20705,N_20605);
nor U21192 (N_21192,N_20618,N_20579);
or U21193 (N_21193,N_20928,N_20597);
nor U21194 (N_21194,N_20569,N_20822);
nand U21195 (N_21195,N_20816,N_20726);
nand U21196 (N_21196,N_20835,N_20558);
nand U21197 (N_21197,N_20971,N_20601);
or U21198 (N_21198,N_20550,N_20981);
and U21199 (N_21199,N_20507,N_20566);
nor U21200 (N_21200,N_20914,N_20554);
and U21201 (N_21201,N_20863,N_20800);
or U21202 (N_21202,N_20609,N_20927);
nor U21203 (N_21203,N_20907,N_20603);
nand U21204 (N_21204,N_20764,N_20748);
and U21205 (N_21205,N_20957,N_20901);
and U21206 (N_21206,N_20919,N_20825);
nand U21207 (N_21207,N_20879,N_20898);
and U21208 (N_21208,N_20810,N_20767);
nor U21209 (N_21209,N_20952,N_20608);
nor U21210 (N_21210,N_20801,N_20817);
nand U21211 (N_21211,N_20542,N_20896);
or U21212 (N_21212,N_20535,N_20847);
or U21213 (N_21213,N_20990,N_20976);
nand U21214 (N_21214,N_20815,N_20730);
nor U21215 (N_21215,N_20883,N_20862);
nor U21216 (N_21216,N_20526,N_20723);
nor U21217 (N_21217,N_20549,N_20690);
nor U21218 (N_21218,N_20599,N_20565);
xnor U21219 (N_21219,N_20808,N_20529);
and U21220 (N_21220,N_20918,N_20890);
nor U21221 (N_21221,N_20857,N_20517);
or U21222 (N_21222,N_20902,N_20564);
and U21223 (N_21223,N_20895,N_20900);
nor U21224 (N_21224,N_20736,N_20753);
or U21225 (N_21225,N_20823,N_20679);
or U21226 (N_21226,N_20574,N_20534);
nor U21227 (N_21227,N_20595,N_20593);
nor U21228 (N_21228,N_20982,N_20598);
nand U21229 (N_21229,N_20821,N_20765);
nand U21230 (N_21230,N_20656,N_20642);
nand U21231 (N_21231,N_20600,N_20956);
nand U21232 (N_21232,N_20899,N_20871);
and U21233 (N_21233,N_20556,N_20658);
nor U21234 (N_21234,N_20959,N_20572);
nor U21235 (N_21235,N_20596,N_20525);
nand U21236 (N_21236,N_20985,N_20555);
and U21237 (N_21237,N_20768,N_20502);
or U21238 (N_21238,N_20523,N_20946);
nor U21239 (N_21239,N_20737,N_20799);
nor U21240 (N_21240,N_20540,N_20675);
nor U21241 (N_21241,N_20980,N_20732);
nand U21242 (N_21242,N_20532,N_20552);
or U21243 (N_21243,N_20645,N_20856);
or U21244 (N_21244,N_20741,N_20913);
or U21245 (N_21245,N_20696,N_20988);
or U21246 (N_21246,N_20578,N_20763);
xnor U21247 (N_21247,N_20739,N_20559);
xor U21248 (N_21248,N_20838,N_20878);
nand U21249 (N_21249,N_20714,N_20802);
nand U21250 (N_21250,N_20887,N_20617);
or U21251 (N_21251,N_20798,N_20790);
nand U21252 (N_21252,N_20942,N_20962);
nor U21253 (N_21253,N_20505,N_20812);
and U21254 (N_21254,N_20619,N_20569);
and U21255 (N_21255,N_20994,N_20794);
or U21256 (N_21256,N_20683,N_20719);
nand U21257 (N_21257,N_20825,N_20849);
and U21258 (N_21258,N_20937,N_20996);
nor U21259 (N_21259,N_20682,N_20508);
nand U21260 (N_21260,N_20993,N_20973);
nor U21261 (N_21261,N_20913,N_20782);
and U21262 (N_21262,N_20885,N_20662);
nand U21263 (N_21263,N_20816,N_20999);
nand U21264 (N_21264,N_20748,N_20763);
nor U21265 (N_21265,N_20786,N_20911);
nor U21266 (N_21266,N_20879,N_20767);
xor U21267 (N_21267,N_20659,N_20879);
nand U21268 (N_21268,N_20606,N_20974);
nor U21269 (N_21269,N_20714,N_20521);
nor U21270 (N_21270,N_20615,N_20748);
or U21271 (N_21271,N_20761,N_20882);
nand U21272 (N_21272,N_20595,N_20749);
xnor U21273 (N_21273,N_20514,N_20938);
nand U21274 (N_21274,N_20683,N_20864);
or U21275 (N_21275,N_20500,N_20984);
nand U21276 (N_21276,N_20968,N_20896);
nand U21277 (N_21277,N_20825,N_20685);
or U21278 (N_21278,N_20627,N_20530);
nor U21279 (N_21279,N_20913,N_20509);
and U21280 (N_21280,N_20972,N_20870);
and U21281 (N_21281,N_20728,N_20793);
or U21282 (N_21282,N_20843,N_20508);
nor U21283 (N_21283,N_20552,N_20688);
and U21284 (N_21284,N_20570,N_20672);
and U21285 (N_21285,N_20729,N_20520);
xor U21286 (N_21286,N_20986,N_20717);
nor U21287 (N_21287,N_20990,N_20912);
nor U21288 (N_21288,N_20764,N_20956);
nor U21289 (N_21289,N_20717,N_20749);
or U21290 (N_21290,N_20895,N_20933);
or U21291 (N_21291,N_20993,N_20773);
or U21292 (N_21292,N_20804,N_20640);
nand U21293 (N_21293,N_20983,N_20988);
nand U21294 (N_21294,N_20619,N_20653);
nand U21295 (N_21295,N_20860,N_20782);
and U21296 (N_21296,N_20908,N_20964);
nor U21297 (N_21297,N_20512,N_20644);
nor U21298 (N_21298,N_20900,N_20632);
nand U21299 (N_21299,N_20623,N_20859);
nand U21300 (N_21300,N_20778,N_20909);
nor U21301 (N_21301,N_20656,N_20756);
and U21302 (N_21302,N_20917,N_20573);
xnor U21303 (N_21303,N_20928,N_20678);
nor U21304 (N_21304,N_20711,N_20780);
or U21305 (N_21305,N_20958,N_20914);
nor U21306 (N_21306,N_20505,N_20810);
nor U21307 (N_21307,N_20853,N_20631);
and U21308 (N_21308,N_20526,N_20985);
nor U21309 (N_21309,N_20916,N_20604);
nor U21310 (N_21310,N_20823,N_20785);
xnor U21311 (N_21311,N_20759,N_20726);
or U21312 (N_21312,N_20760,N_20553);
and U21313 (N_21313,N_20733,N_20596);
xor U21314 (N_21314,N_20592,N_20702);
nor U21315 (N_21315,N_20735,N_20838);
and U21316 (N_21316,N_20728,N_20532);
and U21317 (N_21317,N_20655,N_20591);
nor U21318 (N_21318,N_20820,N_20798);
nand U21319 (N_21319,N_20782,N_20720);
xor U21320 (N_21320,N_20504,N_20662);
or U21321 (N_21321,N_20985,N_20578);
and U21322 (N_21322,N_20866,N_20632);
and U21323 (N_21323,N_20666,N_20592);
nor U21324 (N_21324,N_20846,N_20941);
and U21325 (N_21325,N_20784,N_20548);
nand U21326 (N_21326,N_20955,N_20870);
xor U21327 (N_21327,N_20626,N_20557);
nand U21328 (N_21328,N_20516,N_20536);
and U21329 (N_21329,N_20751,N_20952);
nand U21330 (N_21330,N_20702,N_20602);
xor U21331 (N_21331,N_20714,N_20824);
nor U21332 (N_21332,N_20968,N_20626);
nor U21333 (N_21333,N_20707,N_20603);
or U21334 (N_21334,N_20961,N_20670);
nand U21335 (N_21335,N_20806,N_20551);
nand U21336 (N_21336,N_20942,N_20705);
nand U21337 (N_21337,N_20557,N_20670);
or U21338 (N_21338,N_20854,N_20712);
or U21339 (N_21339,N_20583,N_20791);
nor U21340 (N_21340,N_20841,N_20831);
xor U21341 (N_21341,N_20756,N_20873);
or U21342 (N_21342,N_20917,N_20894);
xnor U21343 (N_21343,N_20696,N_20614);
and U21344 (N_21344,N_20910,N_20724);
or U21345 (N_21345,N_20944,N_20981);
nor U21346 (N_21346,N_20504,N_20578);
or U21347 (N_21347,N_20808,N_20681);
nor U21348 (N_21348,N_20800,N_20798);
or U21349 (N_21349,N_20658,N_20543);
nand U21350 (N_21350,N_20730,N_20708);
and U21351 (N_21351,N_20794,N_20779);
or U21352 (N_21352,N_20924,N_20615);
nor U21353 (N_21353,N_20917,N_20999);
nand U21354 (N_21354,N_20930,N_20665);
or U21355 (N_21355,N_20597,N_20744);
nor U21356 (N_21356,N_20917,N_20933);
xor U21357 (N_21357,N_20663,N_20902);
and U21358 (N_21358,N_20819,N_20659);
nand U21359 (N_21359,N_20992,N_20838);
or U21360 (N_21360,N_20616,N_20864);
and U21361 (N_21361,N_20579,N_20954);
or U21362 (N_21362,N_20552,N_20556);
nand U21363 (N_21363,N_20781,N_20673);
and U21364 (N_21364,N_20799,N_20765);
nand U21365 (N_21365,N_20907,N_20861);
and U21366 (N_21366,N_20580,N_20846);
nand U21367 (N_21367,N_20726,N_20879);
nand U21368 (N_21368,N_20789,N_20739);
nand U21369 (N_21369,N_20955,N_20760);
xnor U21370 (N_21370,N_20589,N_20796);
nand U21371 (N_21371,N_20659,N_20932);
nor U21372 (N_21372,N_20816,N_20889);
nor U21373 (N_21373,N_20837,N_20876);
nor U21374 (N_21374,N_20963,N_20668);
or U21375 (N_21375,N_20608,N_20912);
nand U21376 (N_21376,N_20833,N_20540);
nand U21377 (N_21377,N_20894,N_20990);
or U21378 (N_21378,N_20580,N_20781);
nand U21379 (N_21379,N_20965,N_20708);
or U21380 (N_21380,N_20552,N_20993);
nor U21381 (N_21381,N_20999,N_20579);
nor U21382 (N_21382,N_20850,N_20737);
xnor U21383 (N_21383,N_20850,N_20992);
nand U21384 (N_21384,N_20628,N_20576);
nor U21385 (N_21385,N_20694,N_20670);
nor U21386 (N_21386,N_20819,N_20584);
nor U21387 (N_21387,N_20874,N_20742);
nand U21388 (N_21388,N_20622,N_20692);
nand U21389 (N_21389,N_20546,N_20819);
and U21390 (N_21390,N_20923,N_20600);
nand U21391 (N_21391,N_20776,N_20848);
and U21392 (N_21392,N_20878,N_20844);
xor U21393 (N_21393,N_20915,N_20955);
nor U21394 (N_21394,N_20793,N_20947);
or U21395 (N_21395,N_20922,N_20729);
nand U21396 (N_21396,N_20633,N_20763);
xor U21397 (N_21397,N_20865,N_20530);
or U21398 (N_21398,N_20633,N_20954);
nand U21399 (N_21399,N_20828,N_20631);
or U21400 (N_21400,N_20533,N_20772);
or U21401 (N_21401,N_20796,N_20635);
or U21402 (N_21402,N_20635,N_20922);
nand U21403 (N_21403,N_20897,N_20792);
xnor U21404 (N_21404,N_20537,N_20878);
nand U21405 (N_21405,N_20977,N_20976);
and U21406 (N_21406,N_20542,N_20532);
xnor U21407 (N_21407,N_20931,N_20987);
nand U21408 (N_21408,N_20874,N_20664);
xor U21409 (N_21409,N_20744,N_20734);
and U21410 (N_21410,N_20802,N_20977);
or U21411 (N_21411,N_20687,N_20529);
nand U21412 (N_21412,N_20892,N_20961);
and U21413 (N_21413,N_20974,N_20735);
and U21414 (N_21414,N_20559,N_20526);
nand U21415 (N_21415,N_20801,N_20672);
nand U21416 (N_21416,N_20551,N_20848);
and U21417 (N_21417,N_20689,N_20940);
and U21418 (N_21418,N_20593,N_20669);
nand U21419 (N_21419,N_20971,N_20872);
and U21420 (N_21420,N_20976,N_20614);
or U21421 (N_21421,N_20649,N_20521);
nor U21422 (N_21422,N_20978,N_20934);
nand U21423 (N_21423,N_20874,N_20659);
and U21424 (N_21424,N_20717,N_20921);
xnor U21425 (N_21425,N_20970,N_20629);
or U21426 (N_21426,N_20751,N_20829);
or U21427 (N_21427,N_20621,N_20519);
or U21428 (N_21428,N_20820,N_20787);
and U21429 (N_21429,N_20537,N_20918);
nand U21430 (N_21430,N_20737,N_20709);
nand U21431 (N_21431,N_20715,N_20759);
and U21432 (N_21432,N_20788,N_20740);
xor U21433 (N_21433,N_20552,N_20561);
or U21434 (N_21434,N_20525,N_20945);
or U21435 (N_21435,N_20984,N_20554);
nand U21436 (N_21436,N_20647,N_20522);
xor U21437 (N_21437,N_20696,N_20532);
nor U21438 (N_21438,N_20712,N_20687);
nand U21439 (N_21439,N_20801,N_20614);
and U21440 (N_21440,N_20791,N_20632);
nor U21441 (N_21441,N_20795,N_20869);
or U21442 (N_21442,N_20701,N_20801);
nor U21443 (N_21443,N_20504,N_20756);
nand U21444 (N_21444,N_20900,N_20953);
nor U21445 (N_21445,N_20500,N_20640);
nor U21446 (N_21446,N_20940,N_20906);
nand U21447 (N_21447,N_20974,N_20915);
nor U21448 (N_21448,N_20969,N_20604);
or U21449 (N_21449,N_20837,N_20951);
nor U21450 (N_21450,N_20762,N_20526);
nor U21451 (N_21451,N_20781,N_20636);
and U21452 (N_21452,N_20853,N_20719);
nor U21453 (N_21453,N_20513,N_20612);
nor U21454 (N_21454,N_20633,N_20595);
or U21455 (N_21455,N_20534,N_20739);
nand U21456 (N_21456,N_20851,N_20754);
xnor U21457 (N_21457,N_20729,N_20782);
xnor U21458 (N_21458,N_20706,N_20749);
or U21459 (N_21459,N_20928,N_20852);
nand U21460 (N_21460,N_20712,N_20522);
nand U21461 (N_21461,N_20893,N_20667);
nor U21462 (N_21462,N_20517,N_20589);
or U21463 (N_21463,N_20729,N_20710);
nor U21464 (N_21464,N_20734,N_20719);
or U21465 (N_21465,N_20807,N_20522);
xnor U21466 (N_21466,N_20998,N_20570);
nand U21467 (N_21467,N_20696,N_20585);
nor U21468 (N_21468,N_20536,N_20559);
xor U21469 (N_21469,N_20536,N_20738);
or U21470 (N_21470,N_20755,N_20610);
nand U21471 (N_21471,N_20953,N_20694);
and U21472 (N_21472,N_20925,N_20916);
and U21473 (N_21473,N_20613,N_20563);
or U21474 (N_21474,N_20732,N_20510);
or U21475 (N_21475,N_20823,N_20800);
nor U21476 (N_21476,N_20926,N_20580);
or U21477 (N_21477,N_20915,N_20625);
nand U21478 (N_21478,N_20584,N_20944);
nand U21479 (N_21479,N_20569,N_20710);
or U21480 (N_21480,N_20612,N_20574);
and U21481 (N_21481,N_20875,N_20760);
or U21482 (N_21482,N_20811,N_20980);
and U21483 (N_21483,N_20815,N_20622);
nand U21484 (N_21484,N_20526,N_20844);
or U21485 (N_21485,N_20917,N_20911);
or U21486 (N_21486,N_20943,N_20911);
xor U21487 (N_21487,N_20615,N_20635);
xnor U21488 (N_21488,N_20832,N_20889);
nor U21489 (N_21489,N_20741,N_20684);
nand U21490 (N_21490,N_20951,N_20533);
or U21491 (N_21491,N_20971,N_20765);
or U21492 (N_21492,N_20958,N_20940);
xor U21493 (N_21493,N_20798,N_20519);
and U21494 (N_21494,N_20558,N_20616);
xnor U21495 (N_21495,N_20955,N_20843);
nand U21496 (N_21496,N_20616,N_20634);
or U21497 (N_21497,N_20530,N_20885);
or U21498 (N_21498,N_20948,N_20936);
and U21499 (N_21499,N_20559,N_20723);
xnor U21500 (N_21500,N_21263,N_21250);
nor U21501 (N_21501,N_21113,N_21122);
nor U21502 (N_21502,N_21292,N_21481);
xor U21503 (N_21503,N_21178,N_21309);
xor U21504 (N_21504,N_21044,N_21325);
nand U21505 (N_21505,N_21395,N_21487);
or U21506 (N_21506,N_21156,N_21240);
and U21507 (N_21507,N_21143,N_21125);
nand U21508 (N_21508,N_21329,N_21304);
nand U21509 (N_21509,N_21248,N_21008);
nand U21510 (N_21510,N_21389,N_21251);
nand U21511 (N_21511,N_21343,N_21406);
nand U21512 (N_21512,N_21147,N_21047);
nor U21513 (N_21513,N_21215,N_21187);
and U21514 (N_21514,N_21166,N_21085);
nor U21515 (N_21515,N_21444,N_21064);
nand U21516 (N_21516,N_21277,N_21203);
nand U21517 (N_21517,N_21446,N_21477);
nand U21518 (N_21518,N_21238,N_21267);
nand U21519 (N_21519,N_21480,N_21126);
or U21520 (N_21520,N_21317,N_21114);
and U21521 (N_21521,N_21077,N_21124);
nand U21522 (N_21522,N_21453,N_21073);
and U21523 (N_21523,N_21378,N_21375);
nand U21524 (N_21524,N_21297,N_21040);
and U21525 (N_21525,N_21377,N_21014);
nand U21526 (N_21526,N_21318,N_21167);
xnor U21527 (N_21527,N_21239,N_21342);
nor U21528 (N_21528,N_21399,N_21458);
nand U21529 (N_21529,N_21495,N_21025);
nor U21530 (N_21530,N_21404,N_21182);
nand U21531 (N_21531,N_21148,N_21271);
nor U21532 (N_21532,N_21473,N_21053);
or U21533 (N_21533,N_21435,N_21293);
and U21534 (N_21534,N_21123,N_21265);
nand U21535 (N_21535,N_21408,N_21130);
and U21536 (N_21536,N_21099,N_21189);
nor U21537 (N_21537,N_21041,N_21157);
nand U21538 (N_21538,N_21264,N_21321);
and U21539 (N_21539,N_21291,N_21242);
nand U21540 (N_21540,N_21045,N_21288);
and U21541 (N_21541,N_21367,N_21266);
nand U21542 (N_21542,N_21048,N_21362);
nand U21543 (N_21543,N_21348,N_21440);
nor U21544 (N_21544,N_21411,N_21005);
or U21545 (N_21545,N_21015,N_21051);
nand U21546 (N_21546,N_21307,N_21419);
nor U21547 (N_21547,N_21352,N_21088);
xor U21548 (N_21548,N_21455,N_21349);
nor U21549 (N_21549,N_21163,N_21384);
nor U21550 (N_21550,N_21360,N_21192);
or U21551 (N_21551,N_21154,N_21368);
or U21552 (N_21552,N_21018,N_21094);
xnor U21553 (N_21553,N_21082,N_21387);
and U21554 (N_21554,N_21306,N_21494);
nor U21555 (N_21555,N_21075,N_21165);
xor U21556 (N_21556,N_21485,N_21465);
or U21557 (N_21557,N_21020,N_21424);
nand U21558 (N_21558,N_21057,N_21247);
or U21559 (N_21559,N_21228,N_21017);
and U21560 (N_21560,N_21497,N_21115);
nand U21561 (N_21561,N_21185,N_21137);
and U21562 (N_21562,N_21102,N_21139);
or U21563 (N_21563,N_21338,N_21209);
nor U21564 (N_21564,N_21393,N_21245);
nor U21565 (N_21565,N_21086,N_21398);
xnor U21566 (N_21566,N_21168,N_21207);
or U21567 (N_21567,N_21253,N_21069);
nor U21568 (N_21568,N_21451,N_21422);
nor U21569 (N_21569,N_21090,N_21350);
nand U21570 (N_21570,N_21030,N_21391);
or U21571 (N_21571,N_21300,N_21272);
or U21572 (N_21572,N_21080,N_21294);
or U21573 (N_21573,N_21110,N_21109);
nor U21574 (N_21574,N_21002,N_21042);
and U21575 (N_21575,N_21149,N_21146);
and U21576 (N_21576,N_21258,N_21347);
or U21577 (N_21577,N_21260,N_21356);
and U21578 (N_21578,N_21442,N_21478);
and U21579 (N_21579,N_21161,N_21438);
and U21580 (N_21580,N_21326,N_21198);
nor U21581 (N_21581,N_21417,N_21131);
nor U21582 (N_21582,N_21308,N_21474);
and U21583 (N_21583,N_21006,N_21046);
and U21584 (N_21584,N_21078,N_21032);
and U21585 (N_21585,N_21132,N_21327);
and U21586 (N_21586,N_21281,N_21276);
nand U21587 (N_21587,N_21211,N_21496);
xor U21588 (N_21588,N_21268,N_21400);
or U21589 (N_21589,N_21336,N_21394);
nand U21590 (N_21590,N_21358,N_21074);
nand U21591 (N_21591,N_21434,N_21108);
and U21592 (N_21592,N_21106,N_21230);
nor U21593 (N_21593,N_21289,N_21369);
or U21594 (N_21594,N_21103,N_21013);
nor U21595 (N_21595,N_21364,N_21096);
nor U21596 (N_21596,N_21246,N_21426);
xor U21597 (N_21597,N_21062,N_21221);
nor U21598 (N_21598,N_21205,N_21463);
nor U21599 (N_21599,N_21470,N_21035);
and U21600 (N_21600,N_21299,N_21144);
nand U21601 (N_21601,N_21060,N_21379);
nand U21602 (N_21602,N_21070,N_21202);
nand U21603 (N_21603,N_21218,N_21031);
nand U21604 (N_21604,N_21216,N_21019);
nand U21605 (N_21605,N_21244,N_21186);
nand U21606 (N_21606,N_21081,N_21098);
and U21607 (N_21607,N_21101,N_21493);
and U21608 (N_21608,N_21104,N_21208);
nand U21609 (N_21609,N_21488,N_21012);
nand U21610 (N_21610,N_21427,N_21397);
nand U21611 (N_21611,N_21100,N_21199);
nor U21612 (N_21612,N_21409,N_21471);
and U21613 (N_21613,N_21127,N_21024);
and U21614 (N_21614,N_21227,N_21357);
nand U21615 (N_21615,N_21311,N_21283);
nand U21616 (N_21616,N_21105,N_21155);
nor U21617 (N_21617,N_21193,N_21055);
nor U21618 (N_21618,N_21340,N_21022);
nand U21619 (N_21619,N_21302,N_21036);
nor U21620 (N_21620,N_21092,N_21310);
and U21621 (N_21621,N_21217,N_21180);
nor U21622 (N_21622,N_21436,N_21231);
nand U21623 (N_21623,N_21007,N_21043);
and U21624 (N_21624,N_21175,N_21286);
and U21625 (N_21625,N_21396,N_21441);
or U21626 (N_21626,N_21232,N_21275);
nand U21627 (N_21627,N_21344,N_21412);
and U21628 (N_21628,N_21009,N_21003);
nor U21629 (N_21629,N_21392,N_21313);
nor U21630 (N_21630,N_21191,N_21261);
nor U21631 (N_21631,N_21469,N_21213);
nand U21632 (N_21632,N_21120,N_21382);
nand U21633 (N_21633,N_21170,N_21116);
and U21634 (N_21634,N_21454,N_21499);
and U21635 (N_21635,N_21095,N_21079);
nand U21636 (N_21636,N_21459,N_21256);
nand U21637 (N_21637,N_21407,N_21461);
nor U21638 (N_21638,N_21235,N_21129);
and U21639 (N_21639,N_21162,N_21111);
nor U21640 (N_21640,N_21179,N_21087);
nor U21641 (N_21641,N_21121,N_21016);
or U21642 (N_21642,N_21049,N_21363);
xnor U21643 (N_21643,N_21449,N_21462);
nand U21644 (N_21644,N_21257,N_21486);
and U21645 (N_21645,N_21373,N_21330);
nand U21646 (N_21646,N_21158,N_21401);
nand U21647 (N_21647,N_21204,N_21445);
or U21648 (N_21648,N_21195,N_21320);
or U21649 (N_21649,N_21135,N_21091);
nor U21650 (N_21650,N_21214,N_21021);
or U21651 (N_21651,N_21405,N_21038);
and U21652 (N_21652,N_21403,N_21374);
or U21653 (N_21653,N_21278,N_21134);
or U21654 (N_21654,N_21443,N_21262);
or U21655 (N_21655,N_21476,N_21439);
and U21656 (N_21656,N_21071,N_21421);
nor U21657 (N_21657,N_21492,N_21252);
and U21658 (N_21658,N_21067,N_21249);
and U21659 (N_21659,N_21093,N_21468);
or U21660 (N_21660,N_21464,N_21222);
xnor U21661 (N_21661,N_21010,N_21328);
and U21662 (N_21662,N_21353,N_21151);
nand U21663 (N_21663,N_21491,N_21118);
nand U21664 (N_21664,N_21065,N_21433);
nor U21665 (N_21665,N_21447,N_21270);
or U21666 (N_21666,N_21279,N_21365);
and U21667 (N_21667,N_21410,N_21174);
nand U21668 (N_21668,N_21037,N_21141);
and U21669 (N_21669,N_21072,N_21346);
and U21670 (N_21670,N_21431,N_21282);
nor U21671 (N_21671,N_21437,N_21223);
nand U21672 (N_21672,N_21425,N_21243);
xnor U21673 (N_21673,N_21273,N_21066);
or U21674 (N_21674,N_21152,N_21226);
or U21675 (N_21675,N_21254,N_21402);
xnor U21676 (N_21676,N_21084,N_21176);
nand U21677 (N_21677,N_21483,N_21172);
nand U21678 (N_21678,N_21333,N_21386);
and U21679 (N_21679,N_21298,N_21322);
nor U21680 (N_21680,N_21448,N_21415);
or U21681 (N_21681,N_21039,N_21224);
nand U21682 (N_21682,N_21316,N_21190);
and U21683 (N_21683,N_21490,N_21196);
and U21684 (N_21684,N_21169,N_21475);
or U21685 (N_21685,N_21107,N_21484);
or U21686 (N_21686,N_21324,N_21285);
or U21687 (N_21687,N_21376,N_21136);
nand U21688 (N_21688,N_21140,N_21117);
xor U21689 (N_21689,N_21089,N_21390);
nor U21690 (N_21690,N_21388,N_21219);
nand U21691 (N_21691,N_21206,N_21068);
nand U21692 (N_21692,N_21112,N_21430);
nand U21693 (N_21693,N_21413,N_21429);
nand U21694 (N_21694,N_21160,N_21332);
or U21695 (N_21695,N_21335,N_21351);
nor U21696 (N_21696,N_21201,N_21050);
nand U21697 (N_21697,N_21380,N_21418);
or U21698 (N_21698,N_21366,N_21138);
nand U21699 (N_21699,N_21128,N_21381);
nor U21700 (N_21700,N_21414,N_21269);
nor U21701 (N_21701,N_21200,N_21133);
nand U21702 (N_21702,N_21029,N_21159);
and U21703 (N_21703,N_21457,N_21056);
nor U21704 (N_21704,N_21063,N_21312);
nand U21705 (N_21705,N_21303,N_21150);
xor U21706 (N_21706,N_21076,N_21234);
or U21707 (N_21707,N_21355,N_21371);
and U21708 (N_21708,N_21472,N_21339);
and U21709 (N_21709,N_21450,N_21173);
or U21710 (N_21710,N_21280,N_21027);
nand U21711 (N_21711,N_21331,N_21059);
or U21712 (N_21712,N_21423,N_21482);
nand U21713 (N_21713,N_21004,N_21337);
nand U21714 (N_21714,N_21181,N_21498);
nor U21715 (N_21715,N_21194,N_21210);
and U21716 (N_21716,N_21034,N_21428);
xnor U21717 (N_21717,N_21001,N_21334);
nand U21718 (N_21718,N_21290,N_21023);
or U21719 (N_21719,N_21197,N_21177);
xor U21720 (N_21720,N_21188,N_21052);
and U21721 (N_21721,N_21054,N_21153);
nor U21722 (N_21722,N_21164,N_21058);
or U21723 (N_21723,N_21323,N_21183);
and U21724 (N_21724,N_21212,N_21370);
or U21725 (N_21725,N_21314,N_21284);
xor U21726 (N_21726,N_21341,N_21460);
and U21727 (N_21727,N_21489,N_21225);
or U21728 (N_21728,N_21241,N_21142);
and U21729 (N_21729,N_21383,N_21000);
and U21730 (N_21730,N_21033,N_21259);
xnor U21731 (N_21731,N_21295,N_21296);
or U21732 (N_21732,N_21011,N_21119);
and U21733 (N_21733,N_21301,N_21274);
xnor U21734 (N_21734,N_21184,N_21385);
nor U21735 (N_21735,N_21229,N_21452);
or U21736 (N_21736,N_21026,N_21097);
nand U21737 (N_21737,N_21420,N_21255);
and U21738 (N_21738,N_21466,N_21359);
nor U21739 (N_21739,N_21028,N_21145);
nor U21740 (N_21740,N_21432,N_21372);
and U21741 (N_21741,N_21345,N_21361);
nand U21742 (N_21742,N_21237,N_21354);
nand U21743 (N_21743,N_21305,N_21479);
or U21744 (N_21744,N_21083,N_21416);
nor U21745 (N_21745,N_21467,N_21061);
nor U21746 (N_21746,N_21220,N_21319);
nand U21747 (N_21747,N_21171,N_21236);
nor U21748 (N_21748,N_21315,N_21287);
or U21749 (N_21749,N_21233,N_21456);
xor U21750 (N_21750,N_21324,N_21473);
nand U21751 (N_21751,N_21177,N_21169);
and U21752 (N_21752,N_21061,N_21457);
or U21753 (N_21753,N_21328,N_21418);
nor U21754 (N_21754,N_21202,N_21177);
nand U21755 (N_21755,N_21377,N_21418);
and U21756 (N_21756,N_21455,N_21209);
xnor U21757 (N_21757,N_21426,N_21023);
and U21758 (N_21758,N_21272,N_21464);
and U21759 (N_21759,N_21094,N_21482);
nand U21760 (N_21760,N_21184,N_21146);
or U21761 (N_21761,N_21334,N_21234);
nand U21762 (N_21762,N_21051,N_21467);
nand U21763 (N_21763,N_21281,N_21487);
and U21764 (N_21764,N_21154,N_21356);
nor U21765 (N_21765,N_21279,N_21354);
nor U21766 (N_21766,N_21087,N_21382);
nor U21767 (N_21767,N_21072,N_21284);
nor U21768 (N_21768,N_21037,N_21409);
nor U21769 (N_21769,N_21439,N_21154);
nor U21770 (N_21770,N_21113,N_21480);
xnor U21771 (N_21771,N_21393,N_21195);
nand U21772 (N_21772,N_21338,N_21422);
nand U21773 (N_21773,N_21353,N_21080);
or U21774 (N_21774,N_21151,N_21167);
xor U21775 (N_21775,N_21091,N_21179);
nand U21776 (N_21776,N_21032,N_21295);
or U21777 (N_21777,N_21487,N_21131);
and U21778 (N_21778,N_21422,N_21261);
or U21779 (N_21779,N_21477,N_21346);
nor U21780 (N_21780,N_21017,N_21434);
and U21781 (N_21781,N_21120,N_21008);
or U21782 (N_21782,N_21206,N_21211);
nor U21783 (N_21783,N_21325,N_21341);
or U21784 (N_21784,N_21038,N_21369);
and U21785 (N_21785,N_21088,N_21496);
and U21786 (N_21786,N_21432,N_21069);
or U21787 (N_21787,N_21274,N_21106);
nor U21788 (N_21788,N_21403,N_21429);
or U21789 (N_21789,N_21044,N_21131);
nor U21790 (N_21790,N_21105,N_21067);
nor U21791 (N_21791,N_21174,N_21168);
nand U21792 (N_21792,N_21457,N_21143);
nor U21793 (N_21793,N_21072,N_21482);
and U21794 (N_21794,N_21158,N_21208);
nand U21795 (N_21795,N_21397,N_21164);
nor U21796 (N_21796,N_21186,N_21219);
nor U21797 (N_21797,N_21241,N_21353);
or U21798 (N_21798,N_21172,N_21197);
nand U21799 (N_21799,N_21021,N_21185);
nand U21800 (N_21800,N_21284,N_21439);
and U21801 (N_21801,N_21475,N_21119);
and U21802 (N_21802,N_21038,N_21260);
nand U21803 (N_21803,N_21380,N_21370);
nor U21804 (N_21804,N_21246,N_21082);
and U21805 (N_21805,N_21155,N_21138);
nor U21806 (N_21806,N_21261,N_21381);
nand U21807 (N_21807,N_21155,N_21363);
and U21808 (N_21808,N_21324,N_21240);
nand U21809 (N_21809,N_21204,N_21307);
or U21810 (N_21810,N_21287,N_21497);
nand U21811 (N_21811,N_21037,N_21484);
xnor U21812 (N_21812,N_21095,N_21182);
nor U21813 (N_21813,N_21280,N_21326);
nand U21814 (N_21814,N_21136,N_21462);
nor U21815 (N_21815,N_21246,N_21337);
nand U21816 (N_21816,N_21371,N_21006);
or U21817 (N_21817,N_21418,N_21296);
and U21818 (N_21818,N_21299,N_21337);
xor U21819 (N_21819,N_21163,N_21267);
or U21820 (N_21820,N_21402,N_21385);
nand U21821 (N_21821,N_21248,N_21007);
and U21822 (N_21822,N_21461,N_21369);
nor U21823 (N_21823,N_21421,N_21324);
nand U21824 (N_21824,N_21135,N_21462);
and U21825 (N_21825,N_21246,N_21326);
nor U21826 (N_21826,N_21496,N_21485);
nand U21827 (N_21827,N_21327,N_21492);
nor U21828 (N_21828,N_21063,N_21437);
nor U21829 (N_21829,N_21421,N_21349);
nand U21830 (N_21830,N_21238,N_21486);
nor U21831 (N_21831,N_21384,N_21363);
nand U21832 (N_21832,N_21312,N_21425);
nor U21833 (N_21833,N_21174,N_21380);
or U21834 (N_21834,N_21178,N_21016);
xnor U21835 (N_21835,N_21131,N_21242);
or U21836 (N_21836,N_21374,N_21195);
nor U21837 (N_21837,N_21320,N_21480);
nor U21838 (N_21838,N_21171,N_21338);
or U21839 (N_21839,N_21444,N_21161);
and U21840 (N_21840,N_21363,N_21464);
nand U21841 (N_21841,N_21085,N_21053);
or U21842 (N_21842,N_21334,N_21395);
nand U21843 (N_21843,N_21119,N_21429);
xnor U21844 (N_21844,N_21482,N_21092);
nand U21845 (N_21845,N_21397,N_21263);
and U21846 (N_21846,N_21092,N_21198);
and U21847 (N_21847,N_21072,N_21146);
nor U21848 (N_21848,N_21058,N_21169);
or U21849 (N_21849,N_21302,N_21431);
nor U21850 (N_21850,N_21076,N_21380);
nor U21851 (N_21851,N_21401,N_21459);
or U21852 (N_21852,N_21304,N_21218);
and U21853 (N_21853,N_21455,N_21035);
nor U21854 (N_21854,N_21373,N_21103);
xnor U21855 (N_21855,N_21171,N_21480);
nand U21856 (N_21856,N_21209,N_21491);
nor U21857 (N_21857,N_21407,N_21078);
nand U21858 (N_21858,N_21484,N_21212);
or U21859 (N_21859,N_21170,N_21028);
nand U21860 (N_21860,N_21220,N_21363);
and U21861 (N_21861,N_21200,N_21096);
or U21862 (N_21862,N_21455,N_21322);
and U21863 (N_21863,N_21286,N_21329);
and U21864 (N_21864,N_21484,N_21077);
nor U21865 (N_21865,N_21456,N_21464);
or U21866 (N_21866,N_21354,N_21231);
nand U21867 (N_21867,N_21392,N_21023);
nor U21868 (N_21868,N_21137,N_21224);
or U21869 (N_21869,N_21131,N_21217);
nor U21870 (N_21870,N_21373,N_21358);
nand U21871 (N_21871,N_21352,N_21085);
nor U21872 (N_21872,N_21056,N_21296);
or U21873 (N_21873,N_21348,N_21338);
nand U21874 (N_21874,N_21419,N_21148);
nor U21875 (N_21875,N_21037,N_21272);
nor U21876 (N_21876,N_21178,N_21105);
or U21877 (N_21877,N_21084,N_21215);
and U21878 (N_21878,N_21142,N_21453);
nor U21879 (N_21879,N_21278,N_21464);
nand U21880 (N_21880,N_21205,N_21020);
nor U21881 (N_21881,N_21227,N_21119);
nand U21882 (N_21882,N_21132,N_21073);
or U21883 (N_21883,N_21246,N_21186);
nor U21884 (N_21884,N_21409,N_21048);
and U21885 (N_21885,N_21320,N_21355);
or U21886 (N_21886,N_21397,N_21015);
nand U21887 (N_21887,N_21229,N_21031);
or U21888 (N_21888,N_21287,N_21327);
and U21889 (N_21889,N_21482,N_21166);
nand U21890 (N_21890,N_21252,N_21034);
nand U21891 (N_21891,N_21446,N_21144);
or U21892 (N_21892,N_21186,N_21281);
nand U21893 (N_21893,N_21488,N_21483);
and U21894 (N_21894,N_21491,N_21389);
nand U21895 (N_21895,N_21367,N_21122);
or U21896 (N_21896,N_21414,N_21018);
or U21897 (N_21897,N_21435,N_21321);
nor U21898 (N_21898,N_21477,N_21315);
nor U21899 (N_21899,N_21193,N_21373);
xor U21900 (N_21900,N_21433,N_21360);
and U21901 (N_21901,N_21262,N_21163);
and U21902 (N_21902,N_21074,N_21081);
or U21903 (N_21903,N_21292,N_21416);
and U21904 (N_21904,N_21018,N_21475);
nor U21905 (N_21905,N_21145,N_21054);
nor U21906 (N_21906,N_21437,N_21002);
xor U21907 (N_21907,N_21382,N_21397);
nor U21908 (N_21908,N_21248,N_21283);
nor U21909 (N_21909,N_21090,N_21056);
xnor U21910 (N_21910,N_21029,N_21409);
xnor U21911 (N_21911,N_21067,N_21330);
nand U21912 (N_21912,N_21055,N_21003);
nand U21913 (N_21913,N_21095,N_21175);
xnor U21914 (N_21914,N_21450,N_21428);
xnor U21915 (N_21915,N_21292,N_21246);
xnor U21916 (N_21916,N_21252,N_21344);
nand U21917 (N_21917,N_21422,N_21065);
nor U21918 (N_21918,N_21454,N_21036);
or U21919 (N_21919,N_21308,N_21101);
nand U21920 (N_21920,N_21277,N_21290);
nor U21921 (N_21921,N_21201,N_21326);
and U21922 (N_21922,N_21113,N_21153);
and U21923 (N_21923,N_21406,N_21045);
and U21924 (N_21924,N_21346,N_21464);
and U21925 (N_21925,N_21087,N_21163);
and U21926 (N_21926,N_21257,N_21040);
nand U21927 (N_21927,N_21295,N_21329);
or U21928 (N_21928,N_21291,N_21127);
nand U21929 (N_21929,N_21431,N_21311);
or U21930 (N_21930,N_21218,N_21130);
or U21931 (N_21931,N_21002,N_21250);
nor U21932 (N_21932,N_21313,N_21037);
nor U21933 (N_21933,N_21472,N_21312);
and U21934 (N_21934,N_21375,N_21187);
nor U21935 (N_21935,N_21297,N_21047);
or U21936 (N_21936,N_21417,N_21139);
nand U21937 (N_21937,N_21042,N_21004);
or U21938 (N_21938,N_21322,N_21230);
and U21939 (N_21939,N_21448,N_21006);
nand U21940 (N_21940,N_21283,N_21315);
nor U21941 (N_21941,N_21196,N_21480);
nor U21942 (N_21942,N_21212,N_21271);
and U21943 (N_21943,N_21152,N_21336);
or U21944 (N_21944,N_21459,N_21420);
nor U21945 (N_21945,N_21482,N_21104);
and U21946 (N_21946,N_21303,N_21050);
nand U21947 (N_21947,N_21176,N_21409);
nand U21948 (N_21948,N_21399,N_21038);
nor U21949 (N_21949,N_21256,N_21003);
and U21950 (N_21950,N_21465,N_21473);
nor U21951 (N_21951,N_21335,N_21412);
or U21952 (N_21952,N_21374,N_21222);
xnor U21953 (N_21953,N_21385,N_21440);
xor U21954 (N_21954,N_21471,N_21332);
nor U21955 (N_21955,N_21041,N_21413);
xnor U21956 (N_21956,N_21310,N_21130);
nor U21957 (N_21957,N_21002,N_21407);
nand U21958 (N_21958,N_21396,N_21103);
and U21959 (N_21959,N_21294,N_21406);
or U21960 (N_21960,N_21154,N_21403);
or U21961 (N_21961,N_21201,N_21162);
xnor U21962 (N_21962,N_21154,N_21011);
nand U21963 (N_21963,N_21388,N_21326);
nand U21964 (N_21964,N_21010,N_21254);
or U21965 (N_21965,N_21338,N_21233);
or U21966 (N_21966,N_21258,N_21075);
or U21967 (N_21967,N_21160,N_21495);
nor U21968 (N_21968,N_21435,N_21339);
or U21969 (N_21969,N_21291,N_21151);
nor U21970 (N_21970,N_21238,N_21343);
nand U21971 (N_21971,N_21214,N_21257);
nor U21972 (N_21972,N_21395,N_21316);
nand U21973 (N_21973,N_21240,N_21235);
and U21974 (N_21974,N_21288,N_21236);
or U21975 (N_21975,N_21356,N_21006);
or U21976 (N_21976,N_21260,N_21430);
nor U21977 (N_21977,N_21008,N_21259);
nor U21978 (N_21978,N_21343,N_21308);
and U21979 (N_21979,N_21292,N_21042);
and U21980 (N_21980,N_21172,N_21241);
nand U21981 (N_21981,N_21201,N_21217);
nand U21982 (N_21982,N_21049,N_21118);
nand U21983 (N_21983,N_21337,N_21134);
or U21984 (N_21984,N_21251,N_21104);
and U21985 (N_21985,N_21063,N_21414);
and U21986 (N_21986,N_21259,N_21032);
nand U21987 (N_21987,N_21398,N_21208);
nand U21988 (N_21988,N_21418,N_21079);
nand U21989 (N_21989,N_21018,N_21150);
nand U21990 (N_21990,N_21493,N_21433);
and U21991 (N_21991,N_21344,N_21242);
xnor U21992 (N_21992,N_21235,N_21321);
nand U21993 (N_21993,N_21411,N_21428);
and U21994 (N_21994,N_21057,N_21375);
and U21995 (N_21995,N_21354,N_21350);
nor U21996 (N_21996,N_21055,N_21104);
nor U21997 (N_21997,N_21043,N_21291);
and U21998 (N_21998,N_21456,N_21371);
nand U21999 (N_21999,N_21322,N_21392);
nand U22000 (N_22000,N_21855,N_21553);
nor U22001 (N_22001,N_21997,N_21751);
and U22002 (N_22002,N_21584,N_21575);
or U22003 (N_22003,N_21673,N_21873);
or U22004 (N_22004,N_21629,N_21608);
and U22005 (N_22005,N_21984,N_21941);
and U22006 (N_22006,N_21870,N_21927);
and U22007 (N_22007,N_21709,N_21819);
or U22008 (N_22008,N_21630,N_21983);
xor U22009 (N_22009,N_21979,N_21681);
and U22010 (N_22010,N_21521,N_21913);
nor U22011 (N_22011,N_21660,N_21885);
or U22012 (N_22012,N_21602,N_21882);
nand U22013 (N_22013,N_21864,N_21563);
nor U22014 (N_22014,N_21957,N_21613);
or U22015 (N_22015,N_21947,N_21515);
nor U22016 (N_22016,N_21924,N_21916);
or U22017 (N_22017,N_21793,N_21974);
nor U22018 (N_22018,N_21918,N_21606);
and U22019 (N_22019,N_21771,N_21768);
nor U22020 (N_22020,N_21999,N_21926);
and U22021 (N_22021,N_21671,N_21654);
or U22022 (N_22022,N_21952,N_21726);
nor U22023 (N_22023,N_21626,N_21933);
xnor U22024 (N_22024,N_21954,N_21544);
or U22025 (N_22025,N_21994,N_21605);
or U22026 (N_22026,N_21734,N_21991);
and U22027 (N_22027,N_21646,N_21794);
and U22028 (N_22028,N_21600,N_21756);
nand U22029 (N_22029,N_21808,N_21677);
nor U22030 (N_22030,N_21839,N_21937);
xor U22031 (N_22031,N_21776,N_21877);
or U22032 (N_22032,N_21825,N_21818);
nand U22033 (N_22033,N_21534,N_21538);
nand U22034 (N_22034,N_21852,N_21610);
xor U22035 (N_22035,N_21783,N_21902);
nor U22036 (N_22036,N_21977,N_21850);
nand U22037 (N_22037,N_21583,N_21814);
or U22038 (N_22038,N_21594,N_21901);
or U22039 (N_22039,N_21505,N_21732);
nand U22040 (N_22040,N_21787,N_21883);
or U22041 (N_22041,N_21747,N_21944);
nand U22042 (N_22042,N_21722,N_21878);
nand U22043 (N_22043,N_21841,N_21692);
nand U22044 (N_22044,N_21807,N_21507);
and U22045 (N_22045,N_21762,N_21548);
or U22046 (N_22046,N_21533,N_21661);
or U22047 (N_22047,N_21909,N_21614);
nand U22048 (N_22048,N_21628,N_21921);
nand U22049 (N_22049,N_21840,N_21767);
nand U22050 (N_22050,N_21580,N_21942);
or U22051 (N_22051,N_21753,N_21844);
nor U22052 (N_22052,N_21915,N_21863);
xor U22053 (N_22053,N_21728,N_21639);
nand U22054 (N_22054,N_21955,N_21737);
nor U22055 (N_22055,N_21890,N_21694);
and U22056 (N_22056,N_21817,N_21667);
or U22057 (N_22057,N_21791,N_21826);
nor U22058 (N_22058,N_21510,N_21607);
nor U22059 (N_22059,N_21898,N_21688);
nor U22060 (N_22060,N_21648,N_21752);
nand U22061 (N_22061,N_21953,N_21874);
xnor U22062 (N_22062,N_21867,N_21821);
nor U22063 (N_22063,N_21532,N_21590);
nor U22064 (N_22064,N_21919,N_21653);
nor U22065 (N_22065,N_21846,N_21573);
xor U22066 (N_22066,N_21558,N_21788);
or U22067 (N_22067,N_21812,N_21778);
nand U22068 (N_22068,N_21589,N_21781);
nor U22069 (N_22069,N_21823,N_21931);
or U22070 (N_22070,N_21950,N_21830);
nor U22071 (N_22071,N_21854,N_21765);
and U22072 (N_22072,N_21509,N_21685);
nand U22073 (N_22073,N_21718,N_21743);
and U22074 (N_22074,N_21739,N_21985);
nand U22075 (N_22075,N_21888,N_21966);
and U22076 (N_22076,N_21861,N_21615);
and U22077 (N_22077,N_21832,N_21755);
nor U22078 (N_22078,N_21849,N_21655);
xnor U22079 (N_22079,N_21559,N_21552);
or U22080 (N_22080,N_21662,N_21535);
and U22081 (N_22081,N_21705,N_21881);
nor U22082 (N_22082,N_21784,N_21690);
xor U22083 (N_22083,N_21570,N_21960);
and U22084 (N_22084,N_21813,N_21623);
nor U22085 (N_22085,N_21893,N_21581);
or U22086 (N_22086,N_21631,N_21750);
nor U22087 (N_22087,N_21820,N_21634);
or U22088 (N_22088,N_21550,N_21892);
or U22089 (N_22089,N_21706,N_21522);
nor U22090 (N_22090,N_21514,N_21635);
nand U22091 (N_22091,N_21990,N_21665);
nand U22092 (N_22092,N_21982,N_21545);
nand U22093 (N_22093,N_21922,N_21633);
xnor U22094 (N_22094,N_21556,N_21551);
or U22095 (N_22095,N_21757,N_21658);
or U22096 (N_22096,N_21780,N_21712);
xor U22097 (N_22097,N_21934,N_21619);
nand U22098 (N_22098,N_21569,N_21847);
and U22099 (N_22099,N_21714,N_21592);
and U22100 (N_22100,N_21541,N_21764);
or U22101 (N_22101,N_21586,N_21572);
and U22102 (N_22102,N_21704,N_21799);
or U22103 (N_22103,N_21988,N_21987);
nor U22104 (N_22104,N_21622,N_21809);
or U22105 (N_22105,N_21891,N_21956);
or U22106 (N_22106,N_21880,N_21696);
and U22107 (N_22107,N_21785,N_21993);
nand U22108 (N_22108,N_21822,N_21645);
nand U22109 (N_22109,N_21806,N_21659);
nand U22110 (N_22110,N_21872,N_21742);
or U22111 (N_22111,N_21708,N_21568);
or U22112 (N_22112,N_21989,N_21961);
and U22113 (N_22113,N_21504,N_21511);
or U22114 (N_22114,N_21731,N_21998);
nor U22115 (N_22115,N_21502,N_21930);
xnor U22116 (N_22116,N_21679,N_21682);
or U22117 (N_22117,N_21560,N_21876);
xnor U22118 (N_22118,N_21506,N_21981);
nand U22119 (N_22119,N_21740,N_21946);
and U22120 (N_22120,N_21640,N_21903);
or U22121 (N_22121,N_21700,N_21908);
or U22122 (N_22122,N_21896,N_21958);
or U22123 (N_22123,N_21674,N_21678);
nor U22124 (N_22124,N_21699,N_21729);
or U22125 (N_22125,N_21805,N_21547);
or U22126 (N_22126,N_21798,N_21695);
xor U22127 (N_22127,N_21929,N_21702);
or U22128 (N_22128,N_21576,N_21627);
nand U22129 (N_22129,N_21815,N_21748);
and U22130 (N_22130,N_21656,N_21663);
or U22131 (N_22131,N_21795,N_21831);
and U22132 (N_22132,N_21760,N_21759);
or U22133 (N_22133,N_21668,N_21527);
and U22134 (N_22134,N_21860,N_21777);
and U22135 (N_22135,N_21680,N_21536);
or U22136 (N_22136,N_21526,N_21666);
xnor U22137 (N_22137,N_21632,N_21717);
xnor U22138 (N_22138,N_21604,N_21828);
nor U22139 (N_22139,N_21936,N_21683);
nand U22140 (N_22140,N_21508,N_21554);
and U22141 (N_22141,N_21995,N_21932);
nand U22142 (N_22142,N_21889,N_21766);
nand U22143 (N_22143,N_21657,N_21843);
nor U22144 (N_22144,N_21624,N_21968);
and U22145 (N_22145,N_21561,N_21897);
and U22146 (N_22146,N_21736,N_21923);
nand U22147 (N_22147,N_21693,N_21625);
nor U22148 (N_22148,N_21928,N_21720);
nor U22149 (N_22149,N_21910,N_21528);
and U22150 (N_22150,N_21962,N_21925);
nand U22151 (N_22151,N_21804,N_21567);
nand U22152 (N_22152,N_21676,N_21963);
and U22153 (N_22153,N_21911,N_21557);
or U22154 (N_22154,N_21986,N_21859);
and U22155 (N_22155,N_21851,N_21786);
and U22156 (N_22156,N_21517,N_21647);
and U22157 (N_22157,N_21912,N_21618);
and U22158 (N_22158,N_21578,N_21858);
and U22159 (N_22159,N_21672,N_21862);
nor U22160 (N_22160,N_21789,N_21675);
or U22161 (N_22161,N_21698,N_21866);
nor U22162 (N_22162,N_21827,N_21723);
xor U22163 (N_22163,N_21976,N_21503);
nor U22164 (N_22164,N_21621,N_21810);
nor U22165 (N_22165,N_21713,N_21745);
nand U22166 (N_22166,N_21543,N_21500);
nand U22167 (N_22167,N_21530,N_21727);
nand U22168 (N_22168,N_21501,N_21643);
xnor U22169 (N_22169,N_21642,N_21865);
nor U22170 (N_22170,N_21733,N_21687);
and U22171 (N_22171,N_21721,N_21894);
and U22172 (N_22172,N_21920,N_21711);
nor U22173 (N_22173,N_21939,N_21996);
nor U22174 (N_22174,N_21595,N_21638);
nor U22175 (N_22175,N_21649,N_21582);
or U22176 (N_22176,N_21591,N_21574);
and U22177 (N_22177,N_21636,N_21965);
nand U22178 (N_22178,N_21973,N_21773);
nor U22179 (N_22179,N_21587,N_21803);
nor U22180 (N_22180,N_21971,N_21644);
xnor U22181 (N_22181,N_21875,N_21524);
nand U22182 (N_22182,N_21564,N_21758);
xor U22183 (N_22183,N_21829,N_21585);
nand U22184 (N_22184,N_21900,N_21964);
xor U22185 (N_22185,N_21761,N_21887);
xnor U22186 (N_22186,N_21703,N_21691);
and U22187 (N_22187,N_21970,N_21801);
nand U22188 (N_22188,N_21738,N_21907);
nand U22189 (N_22189,N_21641,N_21725);
nor U22190 (N_22190,N_21774,N_21571);
and U22191 (N_22191,N_21686,N_21652);
or U22192 (N_22192,N_21797,N_21565);
and U22193 (N_22193,N_21518,N_21537);
nand U22194 (N_22194,N_21669,N_21519);
or U22195 (N_22195,N_21938,N_21904);
nor U22196 (N_22196,N_21617,N_21601);
and U22197 (N_22197,N_21972,N_21857);
and U22198 (N_22198,N_21992,N_21612);
or U22199 (N_22199,N_21520,N_21539);
nand U22200 (N_22200,N_21792,N_21802);
nor U22201 (N_22201,N_21744,N_21837);
xor U22202 (N_22202,N_21790,N_21651);
or U22203 (N_22203,N_21512,N_21833);
and U22204 (N_22204,N_21868,N_21746);
or U22205 (N_22205,N_21741,N_21869);
xor U22206 (N_22206,N_21945,N_21555);
nand U22207 (N_22207,N_21967,N_21513);
or U22208 (N_22208,N_21597,N_21879);
nand U22209 (N_22209,N_21684,N_21664);
xor U22210 (N_22210,N_21531,N_21853);
xnor U22211 (N_22211,N_21609,N_21782);
nand U22212 (N_22212,N_21730,N_21980);
xor U22213 (N_22213,N_21525,N_21588);
and U22214 (N_22214,N_21701,N_21735);
and U22215 (N_22215,N_21914,N_21775);
nor U22216 (N_22216,N_21542,N_21710);
and U22217 (N_22217,N_21611,N_21770);
nor U22218 (N_22218,N_21779,N_21834);
nand U22219 (N_22219,N_21838,N_21516);
xnor U22220 (N_22220,N_21824,N_21689);
or U22221 (N_22221,N_21577,N_21523);
or U22222 (N_22222,N_21562,N_21905);
or U22223 (N_22223,N_21724,N_21836);
and U22224 (N_22224,N_21899,N_21951);
nor U22225 (N_22225,N_21754,N_21707);
or U22226 (N_22226,N_21884,N_21715);
nand U22227 (N_22227,N_21603,N_21845);
or U22228 (N_22228,N_21637,N_21975);
or U22229 (N_22229,N_21856,N_21895);
nor U22230 (N_22230,N_21796,N_21697);
xor U22231 (N_22231,N_21763,N_21616);
or U22232 (N_22232,N_21540,N_21620);
and U22233 (N_22233,N_21579,N_21811);
and U22234 (N_22234,N_21749,N_21549);
and U22235 (N_22235,N_21842,N_21940);
xor U22236 (N_22236,N_21835,N_21978);
nand U22237 (N_22237,N_21906,N_21599);
nand U22238 (N_22238,N_21670,N_21917);
nor U22239 (N_22239,N_21772,N_21719);
nand U22240 (N_22240,N_21598,N_21769);
or U22241 (N_22241,N_21948,N_21650);
nor U22242 (N_22242,N_21529,N_21871);
nor U22243 (N_22243,N_21716,N_21848);
nand U22244 (N_22244,N_21943,N_21816);
nor U22245 (N_22245,N_21800,N_21596);
and U22246 (N_22246,N_21593,N_21935);
nor U22247 (N_22247,N_21886,N_21566);
or U22248 (N_22248,N_21949,N_21546);
nor U22249 (N_22249,N_21969,N_21959);
and U22250 (N_22250,N_21551,N_21684);
nand U22251 (N_22251,N_21824,N_21734);
or U22252 (N_22252,N_21597,N_21963);
nor U22253 (N_22253,N_21751,N_21978);
nor U22254 (N_22254,N_21726,N_21612);
and U22255 (N_22255,N_21627,N_21522);
or U22256 (N_22256,N_21970,N_21674);
xnor U22257 (N_22257,N_21791,N_21836);
or U22258 (N_22258,N_21760,N_21946);
and U22259 (N_22259,N_21536,N_21721);
nand U22260 (N_22260,N_21865,N_21777);
nand U22261 (N_22261,N_21563,N_21767);
xnor U22262 (N_22262,N_21623,N_21626);
nor U22263 (N_22263,N_21943,N_21529);
or U22264 (N_22264,N_21504,N_21966);
nand U22265 (N_22265,N_21855,N_21951);
or U22266 (N_22266,N_21566,N_21565);
and U22267 (N_22267,N_21563,N_21744);
nor U22268 (N_22268,N_21852,N_21753);
and U22269 (N_22269,N_21877,N_21742);
nor U22270 (N_22270,N_21693,N_21972);
and U22271 (N_22271,N_21505,N_21985);
nor U22272 (N_22272,N_21940,N_21878);
and U22273 (N_22273,N_21847,N_21653);
or U22274 (N_22274,N_21993,N_21852);
nand U22275 (N_22275,N_21806,N_21500);
and U22276 (N_22276,N_21921,N_21690);
nand U22277 (N_22277,N_21710,N_21963);
and U22278 (N_22278,N_21502,N_21571);
or U22279 (N_22279,N_21839,N_21851);
and U22280 (N_22280,N_21682,N_21786);
nor U22281 (N_22281,N_21700,N_21559);
nor U22282 (N_22282,N_21655,N_21702);
and U22283 (N_22283,N_21874,N_21618);
or U22284 (N_22284,N_21902,N_21813);
xor U22285 (N_22285,N_21748,N_21614);
and U22286 (N_22286,N_21660,N_21762);
nor U22287 (N_22287,N_21924,N_21652);
and U22288 (N_22288,N_21641,N_21727);
and U22289 (N_22289,N_21635,N_21679);
or U22290 (N_22290,N_21808,N_21901);
and U22291 (N_22291,N_21877,N_21763);
nand U22292 (N_22292,N_21974,N_21644);
and U22293 (N_22293,N_21821,N_21942);
and U22294 (N_22294,N_21611,N_21886);
xnor U22295 (N_22295,N_21858,N_21613);
nand U22296 (N_22296,N_21528,N_21960);
nor U22297 (N_22297,N_21850,N_21795);
or U22298 (N_22298,N_21932,N_21698);
or U22299 (N_22299,N_21595,N_21831);
nor U22300 (N_22300,N_21990,N_21843);
xnor U22301 (N_22301,N_21944,N_21580);
and U22302 (N_22302,N_21702,N_21774);
and U22303 (N_22303,N_21789,N_21738);
xnor U22304 (N_22304,N_21650,N_21983);
xor U22305 (N_22305,N_21626,N_21617);
and U22306 (N_22306,N_21955,N_21639);
or U22307 (N_22307,N_21728,N_21548);
or U22308 (N_22308,N_21521,N_21522);
and U22309 (N_22309,N_21752,N_21850);
nor U22310 (N_22310,N_21559,N_21697);
nor U22311 (N_22311,N_21651,N_21823);
nand U22312 (N_22312,N_21770,N_21636);
nand U22313 (N_22313,N_21561,N_21682);
or U22314 (N_22314,N_21755,N_21890);
xnor U22315 (N_22315,N_21811,N_21958);
or U22316 (N_22316,N_21707,N_21830);
xnor U22317 (N_22317,N_21709,N_21859);
nand U22318 (N_22318,N_21947,N_21654);
or U22319 (N_22319,N_21605,N_21501);
or U22320 (N_22320,N_21728,N_21717);
nand U22321 (N_22321,N_21958,N_21898);
and U22322 (N_22322,N_21961,N_21982);
and U22323 (N_22323,N_21894,N_21673);
and U22324 (N_22324,N_21852,N_21589);
and U22325 (N_22325,N_21946,N_21680);
and U22326 (N_22326,N_21510,N_21995);
or U22327 (N_22327,N_21921,N_21834);
nand U22328 (N_22328,N_21573,N_21802);
nor U22329 (N_22329,N_21579,N_21713);
nand U22330 (N_22330,N_21747,N_21846);
nand U22331 (N_22331,N_21795,N_21887);
or U22332 (N_22332,N_21567,N_21982);
xnor U22333 (N_22333,N_21766,N_21646);
nor U22334 (N_22334,N_21549,N_21810);
nor U22335 (N_22335,N_21990,N_21574);
and U22336 (N_22336,N_21592,N_21753);
nand U22337 (N_22337,N_21832,N_21704);
nand U22338 (N_22338,N_21782,N_21928);
or U22339 (N_22339,N_21669,N_21752);
nand U22340 (N_22340,N_21791,N_21545);
and U22341 (N_22341,N_21937,N_21586);
nor U22342 (N_22342,N_21993,N_21703);
xnor U22343 (N_22343,N_21597,N_21510);
and U22344 (N_22344,N_21718,N_21966);
and U22345 (N_22345,N_21630,N_21633);
or U22346 (N_22346,N_21974,N_21828);
nor U22347 (N_22347,N_21583,N_21786);
nand U22348 (N_22348,N_21689,N_21830);
nor U22349 (N_22349,N_21775,N_21506);
or U22350 (N_22350,N_21682,N_21507);
nand U22351 (N_22351,N_21954,N_21702);
or U22352 (N_22352,N_21860,N_21755);
nor U22353 (N_22353,N_21686,N_21908);
and U22354 (N_22354,N_21790,N_21942);
and U22355 (N_22355,N_21816,N_21849);
nand U22356 (N_22356,N_21673,N_21591);
and U22357 (N_22357,N_21876,N_21534);
and U22358 (N_22358,N_21638,N_21949);
nor U22359 (N_22359,N_21821,N_21973);
and U22360 (N_22360,N_21770,N_21599);
xor U22361 (N_22361,N_21792,N_21844);
nor U22362 (N_22362,N_21555,N_21978);
nand U22363 (N_22363,N_21668,N_21770);
and U22364 (N_22364,N_21956,N_21772);
nor U22365 (N_22365,N_21909,N_21623);
and U22366 (N_22366,N_21620,N_21568);
and U22367 (N_22367,N_21516,N_21801);
or U22368 (N_22368,N_21943,N_21915);
nand U22369 (N_22369,N_21860,N_21667);
and U22370 (N_22370,N_21589,N_21680);
and U22371 (N_22371,N_21993,N_21680);
and U22372 (N_22372,N_21538,N_21596);
and U22373 (N_22373,N_21677,N_21772);
and U22374 (N_22374,N_21754,N_21833);
and U22375 (N_22375,N_21649,N_21981);
nor U22376 (N_22376,N_21967,N_21929);
or U22377 (N_22377,N_21969,N_21514);
nor U22378 (N_22378,N_21814,N_21823);
and U22379 (N_22379,N_21605,N_21930);
nand U22380 (N_22380,N_21724,N_21936);
and U22381 (N_22381,N_21825,N_21835);
nand U22382 (N_22382,N_21961,N_21924);
nand U22383 (N_22383,N_21999,N_21868);
nor U22384 (N_22384,N_21510,N_21898);
nand U22385 (N_22385,N_21980,N_21572);
or U22386 (N_22386,N_21570,N_21543);
and U22387 (N_22387,N_21724,N_21912);
nor U22388 (N_22388,N_21686,N_21552);
and U22389 (N_22389,N_21547,N_21531);
xor U22390 (N_22390,N_21881,N_21563);
nand U22391 (N_22391,N_21733,N_21643);
or U22392 (N_22392,N_21626,N_21912);
xor U22393 (N_22393,N_21677,N_21618);
nor U22394 (N_22394,N_21673,N_21581);
nand U22395 (N_22395,N_21827,N_21610);
or U22396 (N_22396,N_21817,N_21801);
nor U22397 (N_22397,N_21517,N_21650);
or U22398 (N_22398,N_21584,N_21887);
nor U22399 (N_22399,N_21742,N_21572);
nor U22400 (N_22400,N_21530,N_21615);
or U22401 (N_22401,N_21803,N_21644);
nor U22402 (N_22402,N_21840,N_21638);
nand U22403 (N_22403,N_21531,N_21778);
nand U22404 (N_22404,N_21830,N_21750);
nand U22405 (N_22405,N_21713,N_21832);
or U22406 (N_22406,N_21680,N_21944);
nand U22407 (N_22407,N_21550,N_21655);
xnor U22408 (N_22408,N_21584,N_21826);
and U22409 (N_22409,N_21645,N_21508);
and U22410 (N_22410,N_21861,N_21658);
nor U22411 (N_22411,N_21547,N_21791);
nand U22412 (N_22412,N_21576,N_21818);
or U22413 (N_22413,N_21857,N_21716);
or U22414 (N_22414,N_21785,N_21559);
and U22415 (N_22415,N_21847,N_21992);
and U22416 (N_22416,N_21742,N_21957);
or U22417 (N_22417,N_21692,N_21892);
nand U22418 (N_22418,N_21862,N_21721);
nor U22419 (N_22419,N_21855,N_21505);
and U22420 (N_22420,N_21652,N_21562);
and U22421 (N_22421,N_21933,N_21932);
nor U22422 (N_22422,N_21853,N_21521);
xor U22423 (N_22423,N_21925,N_21887);
and U22424 (N_22424,N_21659,N_21503);
nor U22425 (N_22425,N_21638,N_21819);
nand U22426 (N_22426,N_21991,N_21557);
xor U22427 (N_22427,N_21673,N_21787);
nor U22428 (N_22428,N_21849,N_21888);
and U22429 (N_22429,N_21598,N_21987);
nand U22430 (N_22430,N_21903,N_21951);
and U22431 (N_22431,N_21921,N_21721);
and U22432 (N_22432,N_21533,N_21698);
and U22433 (N_22433,N_21886,N_21920);
or U22434 (N_22434,N_21776,N_21621);
nor U22435 (N_22435,N_21561,N_21805);
and U22436 (N_22436,N_21840,N_21668);
and U22437 (N_22437,N_21907,N_21668);
and U22438 (N_22438,N_21594,N_21821);
or U22439 (N_22439,N_21743,N_21670);
nand U22440 (N_22440,N_21531,N_21834);
nand U22441 (N_22441,N_21995,N_21593);
nand U22442 (N_22442,N_21598,N_21919);
or U22443 (N_22443,N_21561,N_21649);
and U22444 (N_22444,N_21549,N_21723);
nand U22445 (N_22445,N_21682,N_21739);
and U22446 (N_22446,N_21680,N_21596);
nand U22447 (N_22447,N_21805,N_21824);
xnor U22448 (N_22448,N_21579,N_21969);
xnor U22449 (N_22449,N_21745,N_21575);
and U22450 (N_22450,N_21779,N_21698);
or U22451 (N_22451,N_21670,N_21947);
and U22452 (N_22452,N_21884,N_21686);
and U22453 (N_22453,N_21753,N_21617);
or U22454 (N_22454,N_21565,N_21834);
or U22455 (N_22455,N_21829,N_21563);
nor U22456 (N_22456,N_21957,N_21981);
nand U22457 (N_22457,N_21937,N_21818);
nand U22458 (N_22458,N_21962,N_21541);
nand U22459 (N_22459,N_21883,N_21860);
and U22460 (N_22460,N_21633,N_21860);
nand U22461 (N_22461,N_21531,N_21631);
and U22462 (N_22462,N_21547,N_21835);
or U22463 (N_22463,N_21598,N_21848);
nor U22464 (N_22464,N_21982,N_21591);
nand U22465 (N_22465,N_21883,N_21875);
nand U22466 (N_22466,N_21702,N_21967);
or U22467 (N_22467,N_21656,N_21884);
nor U22468 (N_22468,N_21765,N_21700);
or U22469 (N_22469,N_21657,N_21873);
nor U22470 (N_22470,N_21591,N_21917);
xnor U22471 (N_22471,N_21915,N_21544);
nor U22472 (N_22472,N_21888,N_21727);
and U22473 (N_22473,N_21709,N_21951);
xnor U22474 (N_22474,N_21589,N_21844);
or U22475 (N_22475,N_21527,N_21960);
nand U22476 (N_22476,N_21782,N_21965);
or U22477 (N_22477,N_21792,N_21672);
or U22478 (N_22478,N_21996,N_21612);
nor U22479 (N_22479,N_21623,N_21675);
and U22480 (N_22480,N_21788,N_21804);
nor U22481 (N_22481,N_21998,N_21893);
nand U22482 (N_22482,N_21889,N_21633);
and U22483 (N_22483,N_21755,N_21783);
nor U22484 (N_22484,N_21937,N_21678);
and U22485 (N_22485,N_21624,N_21505);
nand U22486 (N_22486,N_21846,N_21844);
nor U22487 (N_22487,N_21956,N_21763);
nor U22488 (N_22488,N_21920,N_21945);
nand U22489 (N_22489,N_21605,N_21957);
xnor U22490 (N_22490,N_21568,N_21505);
nor U22491 (N_22491,N_21605,N_21512);
nand U22492 (N_22492,N_21807,N_21968);
or U22493 (N_22493,N_21984,N_21996);
xnor U22494 (N_22494,N_21636,N_21875);
and U22495 (N_22495,N_21715,N_21523);
or U22496 (N_22496,N_21783,N_21532);
nand U22497 (N_22497,N_21617,N_21744);
nand U22498 (N_22498,N_21909,N_21771);
and U22499 (N_22499,N_21770,N_21949);
nor U22500 (N_22500,N_22134,N_22390);
nor U22501 (N_22501,N_22219,N_22458);
nand U22502 (N_22502,N_22466,N_22262);
nor U22503 (N_22503,N_22359,N_22397);
or U22504 (N_22504,N_22131,N_22374);
nor U22505 (N_22505,N_22427,N_22209);
or U22506 (N_22506,N_22423,N_22136);
nand U22507 (N_22507,N_22204,N_22017);
nand U22508 (N_22508,N_22127,N_22454);
nand U22509 (N_22509,N_22403,N_22072);
and U22510 (N_22510,N_22206,N_22269);
nor U22511 (N_22511,N_22101,N_22405);
nand U22512 (N_22512,N_22177,N_22163);
and U22513 (N_22513,N_22160,N_22468);
nor U22514 (N_22514,N_22291,N_22042);
and U22515 (N_22515,N_22023,N_22078);
or U22516 (N_22516,N_22325,N_22333);
or U22517 (N_22517,N_22254,N_22259);
or U22518 (N_22518,N_22272,N_22214);
and U22519 (N_22519,N_22106,N_22271);
and U22520 (N_22520,N_22222,N_22370);
xor U22521 (N_22521,N_22159,N_22296);
nand U22522 (N_22522,N_22074,N_22183);
xor U22523 (N_22523,N_22290,N_22084);
nor U22524 (N_22524,N_22158,N_22292);
nand U22525 (N_22525,N_22103,N_22249);
and U22526 (N_22526,N_22276,N_22348);
nor U22527 (N_22527,N_22426,N_22257);
or U22528 (N_22528,N_22231,N_22172);
and U22529 (N_22529,N_22012,N_22373);
nor U22530 (N_22530,N_22137,N_22425);
and U22531 (N_22531,N_22030,N_22489);
or U22532 (N_22532,N_22494,N_22335);
and U22533 (N_22533,N_22297,N_22171);
or U22534 (N_22534,N_22300,N_22413);
or U22535 (N_22535,N_22008,N_22429);
nand U22536 (N_22536,N_22176,N_22245);
and U22537 (N_22537,N_22059,N_22303);
nand U22538 (N_22538,N_22490,N_22221);
xor U22539 (N_22539,N_22394,N_22393);
nand U22540 (N_22540,N_22298,N_22071);
nor U22541 (N_22541,N_22323,N_22332);
or U22542 (N_22542,N_22380,N_22420);
nor U22543 (N_22543,N_22057,N_22308);
or U22544 (N_22544,N_22069,N_22355);
nor U22545 (N_22545,N_22382,N_22418);
xor U22546 (N_22546,N_22428,N_22058);
or U22547 (N_22547,N_22174,N_22217);
nor U22548 (N_22548,N_22266,N_22117);
and U22549 (N_22549,N_22138,N_22463);
nor U22550 (N_22550,N_22493,N_22089);
and U22551 (N_22551,N_22470,N_22419);
nand U22552 (N_22552,N_22144,N_22318);
and U22553 (N_22553,N_22284,N_22295);
xnor U22554 (N_22554,N_22476,N_22436);
nand U22555 (N_22555,N_22422,N_22327);
xor U22556 (N_22556,N_22343,N_22304);
nor U22557 (N_22557,N_22396,N_22368);
nor U22558 (N_22558,N_22313,N_22047);
and U22559 (N_22559,N_22180,N_22184);
and U22560 (N_22560,N_22309,N_22379);
nand U22561 (N_22561,N_22312,N_22481);
nand U22562 (N_22562,N_22234,N_22268);
and U22563 (N_22563,N_22478,N_22113);
and U22564 (N_22564,N_22242,N_22414);
or U22565 (N_22565,N_22079,N_22337);
nor U22566 (N_22566,N_22377,N_22369);
or U22567 (N_22567,N_22031,N_22310);
and U22568 (N_22568,N_22239,N_22086);
and U22569 (N_22569,N_22181,N_22263);
and U22570 (N_22570,N_22256,N_22255);
xor U22571 (N_22571,N_22019,N_22415);
and U22572 (N_22572,N_22020,N_22210);
or U22573 (N_22573,N_22479,N_22356);
nand U22574 (N_22574,N_22366,N_22139);
nand U22575 (N_22575,N_22378,N_22015);
nand U22576 (N_22576,N_22022,N_22041);
or U22577 (N_22577,N_22224,N_22472);
nor U22578 (N_22578,N_22093,N_22046);
xnor U22579 (N_22579,N_22035,N_22142);
or U22580 (N_22580,N_22462,N_22109);
nor U22581 (N_22581,N_22143,N_22112);
or U22582 (N_22582,N_22275,N_22218);
xor U22583 (N_22583,N_22252,N_22100);
or U22584 (N_22584,N_22153,N_22044);
or U22585 (N_22585,N_22484,N_22339);
nor U22586 (N_22586,N_22431,N_22213);
xnor U22587 (N_22587,N_22365,N_22237);
or U22588 (N_22588,N_22443,N_22293);
or U22589 (N_22589,N_22013,N_22082);
and U22590 (N_22590,N_22164,N_22126);
or U22591 (N_22591,N_22205,N_22111);
xor U22592 (N_22592,N_22361,N_22483);
or U22593 (N_22593,N_22283,N_22280);
xnor U22594 (N_22594,N_22445,N_22498);
or U22595 (N_22595,N_22357,N_22354);
or U22596 (N_22596,N_22442,N_22179);
or U22597 (N_22597,N_22444,N_22320);
or U22598 (N_22598,N_22457,N_22401);
and U22599 (N_22599,N_22386,N_22149);
and U22600 (N_22600,N_22238,N_22133);
and U22601 (N_22601,N_22167,N_22244);
nand U22602 (N_22602,N_22384,N_22471);
nand U22603 (N_22603,N_22288,N_22199);
nand U22604 (N_22604,N_22099,N_22034);
and U22605 (N_22605,N_22371,N_22192);
xnor U22606 (N_22606,N_22324,N_22408);
nor U22607 (N_22607,N_22329,N_22250);
or U22608 (N_22608,N_22311,N_22102);
or U22609 (N_22609,N_22236,N_22220);
nand U22610 (N_22610,N_22438,N_22014);
nor U22611 (N_22611,N_22480,N_22452);
nand U22612 (N_22612,N_22281,N_22389);
nand U22613 (N_22613,N_22246,N_22273);
or U22614 (N_22614,N_22228,N_22416);
nor U22615 (N_22615,N_22215,N_22145);
nor U22616 (N_22616,N_22486,N_22289);
nor U22617 (N_22617,N_22331,N_22054);
or U22618 (N_22618,N_22216,N_22460);
and U22619 (N_22619,N_22437,N_22116);
or U22620 (N_22620,N_22433,N_22066);
and U22621 (N_22621,N_22340,N_22182);
xnor U22622 (N_22622,N_22441,N_22195);
xnor U22623 (N_22623,N_22383,N_22169);
nor U22624 (N_22624,N_22287,N_22132);
xnor U22625 (N_22625,N_22187,N_22026);
or U22626 (N_22626,N_22207,N_22347);
nand U22627 (N_22627,N_22388,N_22000);
and U22628 (N_22628,N_22118,N_22417);
nand U22629 (N_22629,N_22248,N_22051);
nand U22630 (N_22630,N_22274,N_22060);
and U22631 (N_22631,N_22029,N_22162);
nand U22632 (N_22632,N_22186,N_22338);
or U22633 (N_22633,N_22038,N_22391);
nand U22634 (N_22634,N_22077,N_22449);
and U22635 (N_22635,N_22439,N_22260);
xor U22636 (N_22636,N_22277,N_22170);
or U22637 (N_22637,N_22049,N_22253);
or U22638 (N_22638,N_22201,N_22240);
nor U22639 (N_22639,N_22451,N_22372);
or U22640 (N_22640,N_22406,N_22353);
or U22641 (N_22641,N_22130,N_22261);
nand U22642 (N_22642,N_22385,N_22191);
nor U22643 (N_22643,N_22342,N_22197);
nor U22644 (N_22644,N_22226,N_22070);
nand U22645 (N_22645,N_22010,N_22025);
or U22646 (N_22646,N_22203,N_22007);
nor U22647 (N_22647,N_22473,N_22032);
or U22648 (N_22648,N_22152,N_22251);
and U22649 (N_22649,N_22302,N_22392);
nand U22650 (N_22650,N_22140,N_22122);
nor U22651 (N_22651,N_22161,N_22211);
nor U22652 (N_22652,N_22430,N_22367);
nor U22653 (N_22653,N_22005,N_22487);
or U22654 (N_22654,N_22033,N_22028);
nor U22655 (N_22655,N_22105,N_22461);
or U22656 (N_22656,N_22196,N_22083);
nor U22657 (N_22657,N_22267,N_22350);
and U22658 (N_22658,N_22168,N_22052);
or U22659 (N_22659,N_22063,N_22027);
or U22660 (N_22660,N_22120,N_22062);
xnor U22661 (N_22661,N_22344,N_22003);
nor U22662 (N_22662,N_22227,N_22056);
and U22663 (N_22663,N_22230,N_22349);
nand U22664 (N_22664,N_22440,N_22004);
and U22665 (N_22665,N_22307,N_22055);
nor U22666 (N_22666,N_22381,N_22096);
xnor U22667 (N_22667,N_22037,N_22185);
and U22668 (N_22668,N_22067,N_22435);
nand U22669 (N_22669,N_22154,N_22114);
and U22670 (N_22670,N_22175,N_22402);
and U22671 (N_22671,N_22061,N_22050);
or U22672 (N_22672,N_22097,N_22173);
and U22673 (N_22673,N_22125,N_22068);
or U22674 (N_22674,N_22194,N_22006);
or U22675 (N_22675,N_22024,N_22235);
and U22676 (N_22676,N_22212,N_22200);
nand U22677 (N_22677,N_22075,N_22317);
nor U22678 (N_22678,N_22225,N_22364);
nor U22679 (N_22679,N_22482,N_22363);
nand U22680 (N_22680,N_22135,N_22156);
nand U22681 (N_22681,N_22410,N_22404);
or U22682 (N_22682,N_22314,N_22198);
or U22683 (N_22683,N_22285,N_22157);
nand U22684 (N_22684,N_22001,N_22474);
nand U22685 (N_22685,N_22351,N_22155);
or U22686 (N_22686,N_22475,N_22421);
or U22687 (N_22687,N_22081,N_22306);
nor U22688 (N_22688,N_22301,N_22232);
nand U22689 (N_22689,N_22341,N_22048);
and U22690 (N_22690,N_22328,N_22223);
nand U22691 (N_22691,N_22459,N_22018);
nand U22692 (N_22692,N_22039,N_22115);
and U22693 (N_22693,N_22319,N_22465);
xor U22694 (N_22694,N_22264,N_22279);
xnor U22695 (N_22695,N_22088,N_22352);
or U22696 (N_22696,N_22098,N_22305);
or U22697 (N_22697,N_22124,N_22085);
or U22698 (N_22698,N_22009,N_22040);
nand U22699 (N_22699,N_22188,N_22002);
nand U22700 (N_22700,N_22147,N_22464);
nor U22701 (N_22701,N_22178,N_22467);
or U22702 (N_22702,N_22488,N_22434);
nand U22703 (N_22703,N_22166,N_22053);
or U22704 (N_22704,N_22450,N_22499);
and U22705 (N_22705,N_22315,N_22286);
nor U22706 (N_22706,N_22491,N_22412);
nor U22707 (N_22707,N_22278,N_22073);
nor U22708 (N_22708,N_22036,N_22330);
xnor U22709 (N_22709,N_22095,N_22129);
nor U22710 (N_22710,N_22326,N_22165);
and U22711 (N_22711,N_22080,N_22360);
nor U22712 (N_22712,N_22150,N_22294);
nand U22713 (N_22713,N_22497,N_22011);
and U22714 (N_22714,N_22243,N_22448);
or U22715 (N_22715,N_22043,N_22065);
and U22716 (N_22716,N_22092,N_22456);
or U22717 (N_22717,N_22110,N_22090);
or U22718 (N_22718,N_22411,N_22399);
nand U22719 (N_22719,N_22123,N_22193);
xor U22720 (N_22720,N_22477,N_22492);
or U22721 (N_22721,N_22202,N_22495);
xnor U22722 (N_22722,N_22241,N_22299);
nand U22723 (N_22723,N_22021,N_22146);
or U22724 (N_22724,N_22104,N_22447);
nand U22725 (N_22725,N_22407,N_22375);
nor U22726 (N_22726,N_22282,N_22119);
nor U22727 (N_22727,N_22455,N_22121);
or U22728 (N_22728,N_22258,N_22398);
and U22729 (N_22729,N_22345,N_22376);
or U22730 (N_22730,N_22107,N_22233);
nor U22731 (N_22731,N_22094,N_22141);
xnor U22732 (N_22732,N_22432,N_22322);
and U22733 (N_22733,N_22108,N_22076);
nor U22734 (N_22734,N_22496,N_22453);
and U22735 (N_22735,N_22424,N_22336);
or U22736 (N_22736,N_22016,N_22064);
or U22737 (N_22737,N_22247,N_22148);
nand U22738 (N_22738,N_22189,N_22270);
nor U22739 (N_22739,N_22387,N_22446);
nand U22740 (N_22740,N_22045,N_22358);
nand U22741 (N_22741,N_22229,N_22400);
xor U22742 (N_22742,N_22190,N_22321);
or U22743 (N_22743,N_22334,N_22265);
xor U22744 (N_22744,N_22128,N_22469);
xnor U22745 (N_22745,N_22087,N_22316);
and U22746 (N_22746,N_22346,N_22485);
nand U22747 (N_22747,N_22208,N_22362);
nand U22748 (N_22748,N_22395,N_22409);
or U22749 (N_22749,N_22091,N_22151);
xor U22750 (N_22750,N_22107,N_22187);
and U22751 (N_22751,N_22080,N_22113);
nand U22752 (N_22752,N_22146,N_22362);
nand U22753 (N_22753,N_22401,N_22317);
and U22754 (N_22754,N_22245,N_22310);
xor U22755 (N_22755,N_22349,N_22418);
or U22756 (N_22756,N_22164,N_22173);
nor U22757 (N_22757,N_22217,N_22344);
and U22758 (N_22758,N_22243,N_22401);
and U22759 (N_22759,N_22113,N_22288);
and U22760 (N_22760,N_22291,N_22384);
nand U22761 (N_22761,N_22104,N_22136);
xor U22762 (N_22762,N_22125,N_22024);
or U22763 (N_22763,N_22480,N_22211);
and U22764 (N_22764,N_22399,N_22104);
and U22765 (N_22765,N_22459,N_22174);
nor U22766 (N_22766,N_22000,N_22307);
nor U22767 (N_22767,N_22216,N_22437);
or U22768 (N_22768,N_22441,N_22481);
xor U22769 (N_22769,N_22279,N_22310);
or U22770 (N_22770,N_22473,N_22298);
and U22771 (N_22771,N_22492,N_22411);
or U22772 (N_22772,N_22286,N_22413);
nor U22773 (N_22773,N_22372,N_22343);
nor U22774 (N_22774,N_22398,N_22474);
nand U22775 (N_22775,N_22118,N_22184);
nor U22776 (N_22776,N_22048,N_22181);
or U22777 (N_22777,N_22352,N_22454);
and U22778 (N_22778,N_22463,N_22098);
nor U22779 (N_22779,N_22383,N_22043);
and U22780 (N_22780,N_22217,N_22194);
nor U22781 (N_22781,N_22141,N_22479);
and U22782 (N_22782,N_22403,N_22001);
and U22783 (N_22783,N_22223,N_22213);
or U22784 (N_22784,N_22141,N_22160);
or U22785 (N_22785,N_22418,N_22166);
and U22786 (N_22786,N_22137,N_22146);
and U22787 (N_22787,N_22455,N_22216);
nand U22788 (N_22788,N_22457,N_22179);
nand U22789 (N_22789,N_22464,N_22111);
nand U22790 (N_22790,N_22399,N_22162);
nor U22791 (N_22791,N_22387,N_22206);
or U22792 (N_22792,N_22399,N_22432);
nor U22793 (N_22793,N_22362,N_22443);
and U22794 (N_22794,N_22165,N_22055);
and U22795 (N_22795,N_22274,N_22187);
nor U22796 (N_22796,N_22311,N_22151);
or U22797 (N_22797,N_22013,N_22311);
or U22798 (N_22798,N_22155,N_22052);
and U22799 (N_22799,N_22452,N_22335);
or U22800 (N_22800,N_22353,N_22475);
nand U22801 (N_22801,N_22237,N_22305);
or U22802 (N_22802,N_22285,N_22068);
nor U22803 (N_22803,N_22116,N_22029);
and U22804 (N_22804,N_22109,N_22359);
nor U22805 (N_22805,N_22480,N_22046);
and U22806 (N_22806,N_22273,N_22078);
nor U22807 (N_22807,N_22393,N_22103);
and U22808 (N_22808,N_22473,N_22309);
or U22809 (N_22809,N_22377,N_22456);
nand U22810 (N_22810,N_22364,N_22145);
nand U22811 (N_22811,N_22025,N_22429);
or U22812 (N_22812,N_22068,N_22063);
or U22813 (N_22813,N_22001,N_22443);
nand U22814 (N_22814,N_22410,N_22405);
nor U22815 (N_22815,N_22068,N_22048);
and U22816 (N_22816,N_22037,N_22194);
and U22817 (N_22817,N_22160,N_22349);
or U22818 (N_22818,N_22461,N_22219);
nor U22819 (N_22819,N_22080,N_22079);
nand U22820 (N_22820,N_22302,N_22221);
nor U22821 (N_22821,N_22405,N_22119);
nand U22822 (N_22822,N_22086,N_22206);
or U22823 (N_22823,N_22101,N_22384);
nor U22824 (N_22824,N_22378,N_22201);
nand U22825 (N_22825,N_22400,N_22482);
nor U22826 (N_22826,N_22367,N_22011);
xor U22827 (N_22827,N_22196,N_22221);
and U22828 (N_22828,N_22372,N_22092);
nor U22829 (N_22829,N_22396,N_22467);
xor U22830 (N_22830,N_22024,N_22144);
nand U22831 (N_22831,N_22182,N_22042);
nor U22832 (N_22832,N_22414,N_22210);
nor U22833 (N_22833,N_22407,N_22023);
and U22834 (N_22834,N_22479,N_22377);
and U22835 (N_22835,N_22118,N_22380);
nor U22836 (N_22836,N_22233,N_22002);
nor U22837 (N_22837,N_22077,N_22416);
and U22838 (N_22838,N_22499,N_22289);
nor U22839 (N_22839,N_22420,N_22077);
nand U22840 (N_22840,N_22116,N_22396);
or U22841 (N_22841,N_22238,N_22294);
nand U22842 (N_22842,N_22189,N_22489);
or U22843 (N_22843,N_22349,N_22319);
nand U22844 (N_22844,N_22050,N_22193);
nor U22845 (N_22845,N_22279,N_22165);
and U22846 (N_22846,N_22104,N_22099);
xnor U22847 (N_22847,N_22470,N_22365);
nand U22848 (N_22848,N_22131,N_22020);
nor U22849 (N_22849,N_22460,N_22415);
or U22850 (N_22850,N_22003,N_22112);
or U22851 (N_22851,N_22066,N_22012);
xor U22852 (N_22852,N_22361,N_22087);
nor U22853 (N_22853,N_22382,N_22064);
nand U22854 (N_22854,N_22291,N_22050);
nand U22855 (N_22855,N_22043,N_22119);
and U22856 (N_22856,N_22003,N_22295);
or U22857 (N_22857,N_22070,N_22033);
or U22858 (N_22858,N_22456,N_22003);
or U22859 (N_22859,N_22416,N_22456);
or U22860 (N_22860,N_22089,N_22423);
nand U22861 (N_22861,N_22188,N_22428);
nor U22862 (N_22862,N_22004,N_22299);
nand U22863 (N_22863,N_22081,N_22180);
or U22864 (N_22864,N_22122,N_22048);
and U22865 (N_22865,N_22092,N_22247);
nor U22866 (N_22866,N_22143,N_22428);
nand U22867 (N_22867,N_22176,N_22125);
or U22868 (N_22868,N_22017,N_22351);
nor U22869 (N_22869,N_22490,N_22382);
nor U22870 (N_22870,N_22186,N_22008);
and U22871 (N_22871,N_22219,N_22117);
nor U22872 (N_22872,N_22241,N_22222);
nand U22873 (N_22873,N_22253,N_22112);
and U22874 (N_22874,N_22371,N_22410);
nor U22875 (N_22875,N_22204,N_22135);
or U22876 (N_22876,N_22327,N_22259);
nor U22877 (N_22877,N_22210,N_22343);
and U22878 (N_22878,N_22069,N_22081);
nand U22879 (N_22879,N_22320,N_22336);
nor U22880 (N_22880,N_22270,N_22249);
nor U22881 (N_22881,N_22005,N_22135);
and U22882 (N_22882,N_22260,N_22391);
and U22883 (N_22883,N_22199,N_22146);
and U22884 (N_22884,N_22202,N_22084);
nor U22885 (N_22885,N_22166,N_22105);
nor U22886 (N_22886,N_22130,N_22158);
and U22887 (N_22887,N_22177,N_22055);
and U22888 (N_22888,N_22160,N_22385);
and U22889 (N_22889,N_22171,N_22314);
nand U22890 (N_22890,N_22386,N_22344);
xnor U22891 (N_22891,N_22352,N_22098);
or U22892 (N_22892,N_22275,N_22017);
nand U22893 (N_22893,N_22219,N_22148);
nor U22894 (N_22894,N_22005,N_22467);
nand U22895 (N_22895,N_22410,N_22107);
nor U22896 (N_22896,N_22032,N_22200);
and U22897 (N_22897,N_22071,N_22063);
nand U22898 (N_22898,N_22497,N_22061);
nand U22899 (N_22899,N_22278,N_22147);
nor U22900 (N_22900,N_22307,N_22117);
xor U22901 (N_22901,N_22454,N_22005);
xor U22902 (N_22902,N_22435,N_22003);
nor U22903 (N_22903,N_22049,N_22393);
and U22904 (N_22904,N_22360,N_22414);
and U22905 (N_22905,N_22149,N_22163);
nand U22906 (N_22906,N_22272,N_22259);
or U22907 (N_22907,N_22229,N_22456);
or U22908 (N_22908,N_22058,N_22279);
and U22909 (N_22909,N_22419,N_22230);
and U22910 (N_22910,N_22409,N_22002);
nand U22911 (N_22911,N_22361,N_22427);
or U22912 (N_22912,N_22411,N_22310);
nor U22913 (N_22913,N_22263,N_22144);
or U22914 (N_22914,N_22268,N_22032);
and U22915 (N_22915,N_22434,N_22463);
and U22916 (N_22916,N_22308,N_22204);
nand U22917 (N_22917,N_22449,N_22155);
and U22918 (N_22918,N_22096,N_22499);
nand U22919 (N_22919,N_22308,N_22177);
or U22920 (N_22920,N_22144,N_22061);
nand U22921 (N_22921,N_22289,N_22209);
or U22922 (N_22922,N_22321,N_22305);
nand U22923 (N_22923,N_22397,N_22300);
and U22924 (N_22924,N_22354,N_22276);
and U22925 (N_22925,N_22053,N_22277);
xor U22926 (N_22926,N_22237,N_22254);
or U22927 (N_22927,N_22300,N_22358);
nand U22928 (N_22928,N_22305,N_22486);
or U22929 (N_22929,N_22115,N_22320);
or U22930 (N_22930,N_22393,N_22194);
nand U22931 (N_22931,N_22170,N_22303);
nor U22932 (N_22932,N_22361,N_22479);
xnor U22933 (N_22933,N_22362,N_22497);
or U22934 (N_22934,N_22154,N_22226);
or U22935 (N_22935,N_22001,N_22320);
nor U22936 (N_22936,N_22420,N_22356);
nand U22937 (N_22937,N_22100,N_22155);
nor U22938 (N_22938,N_22469,N_22358);
nand U22939 (N_22939,N_22084,N_22064);
xnor U22940 (N_22940,N_22482,N_22254);
nor U22941 (N_22941,N_22170,N_22013);
and U22942 (N_22942,N_22242,N_22081);
xor U22943 (N_22943,N_22113,N_22120);
nor U22944 (N_22944,N_22063,N_22057);
or U22945 (N_22945,N_22293,N_22115);
or U22946 (N_22946,N_22367,N_22195);
or U22947 (N_22947,N_22006,N_22069);
and U22948 (N_22948,N_22276,N_22141);
and U22949 (N_22949,N_22153,N_22372);
or U22950 (N_22950,N_22131,N_22047);
or U22951 (N_22951,N_22104,N_22076);
nand U22952 (N_22952,N_22444,N_22293);
and U22953 (N_22953,N_22415,N_22477);
nor U22954 (N_22954,N_22477,N_22039);
xnor U22955 (N_22955,N_22182,N_22462);
and U22956 (N_22956,N_22070,N_22162);
xnor U22957 (N_22957,N_22304,N_22259);
or U22958 (N_22958,N_22370,N_22149);
or U22959 (N_22959,N_22395,N_22138);
or U22960 (N_22960,N_22348,N_22469);
nand U22961 (N_22961,N_22297,N_22078);
or U22962 (N_22962,N_22461,N_22157);
nor U22963 (N_22963,N_22336,N_22420);
xor U22964 (N_22964,N_22284,N_22241);
nand U22965 (N_22965,N_22015,N_22433);
and U22966 (N_22966,N_22381,N_22368);
nor U22967 (N_22967,N_22262,N_22240);
or U22968 (N_22968,N_22333,N_22389);
nand U22969 (N_22969,N_22271,N_22204);
or U22970 (N_22970,N_22152,N_22338);
nor U22971 (N_22971,N_22088,N_22296);
or U22972 (N_22972,N_22293,N_22176);
nand U22973 (N_22973,N_22363,N_22049);
nor U22974 (N_22974,N_22424,N_22083);
or U22975 (N_22975,N_22313,N_22066);
or U22976 (N_22976,N_22169,N_22232);
xnor U22977 (N_22977,N_22390,N_22337);
nor U22978 (N_22978,N_22383,N_22152);
nor U22979 (N_22979,N_22439,N_22321);
and U22980 (N_22980,N_22271,N_22491);
or U22981 (N_22981,N_22472,N_22104);
and U22982 (N_22982,N_22374,N_22073);
or U22983 (N_22983,N_22344,N_22457);
or U22984 (N_22984,N_22399,N_22397);
xor U22985 (N_22985,N_22255,N_22384);
nand U22986 (N_22986,N_22126,N_22000);
or U22987 (N_22987,N_22116,N_22123);
or U22988 (N_22988,N_22341,N_22206);
nand U22989 (N_22989,N_22111,N_22354);
and U22990 (N_22990,N_22142,N_22360);
and U22991 (N_22991,N_22170,N_22171);
nor U22992 (N_22992,N_22349,N_22212);
or U22993 (N_22993,N_22176,N_22441);
nand U22994 (N_22994,N_22029,N_22167);
nor U22995 (N_22995,N_22121,N_22354);
nor U22996 (N_22996,N_22072,N_22357);
or U22997 (N_22997,N_22296,N_22056);
nor U22998 (N_22998,N_22156,N_22493);
nor U22999 (N_22999,N_22052,N_22278);
nor U23000 (N_23000,N_22830,N_22944);
or U23001 (N_23001,N_22972,N_22615);
nand U23002 (N_23002,N_22882,N_22949);
nand U23003 (N_23003,N_22870,N_22618);
and U23004 (N_23004,N_22666,N_22504);
xnor U23005 (N_23005,N_22675,N_22969);
or U23006 (N_23006,N_22913,N_22769);
xnor U23007 (N_23007,N_22650,N_22814);
or U23008 (N_23008,N_22823,N_22794);
xnor U23009 (N_23009,N_22608,N_22693);
or U23010 (N_23010,N_22674,N_22942);
nand U23011 (N_23011,N_22593,N_22788);
or U23012 (N_23012,N_22585,N_22662);
nor U23013 (N_23013,N_22835,N_22992);
or U23014 (N_23014,N_22810,N_22710);
and U23015 (N_23015,N_22565,N_22600);
nor U23016 (N_23016,N_22854,N_22657);
and U23017 (N_23017,N_22754,N_22701);
or U23018 (N_23018,N_22957,N_22645);
xor U23019 (N_23019,N_22812,N_22587);
nand U23020 (N_23020,N_22519,N_22917);
nor U23021 (N_23021,N_22563,N_22603);
nand U23022 (N_23022,N_22885,N_22793);
or U23023 (N_23023,N_22592,N_22890);
nor U23024 (N_23024,N_22895,N_22622);
and U23025 (N_23025,N_22583,N_22781);
or U23026 (N_23026,N_22926,N_22838);
nor U23027 (N_23027,N_22633,N_22771);
nor U23028 (N_23028,N_22652,N_22968);
and U23029 (N_23029,N_22514,N_22667);
nor U23030 (N_23030,N_22651,N_22685);
or U23031 (N_23031,N_22979,N_22982);
xnor U23032 (N_23032,N_22877,N_22828);
or U23033 (N_23033,N_22959,N_22620);
xor U23034 (N_23034,N_22889,N_22530);
or U23035 (N_23035,N_22998,N_22680);
and U23036 (N_23036,N_22630,N_22930);
nor U23037 (N_23037,N_22862,N_22910);
nand U23038 (N_23038,N_22602,N_22574);
nor U23039 (N_23039,N_22786,N_22797);
xnor U23040 (N_23040,N_22661,N_22768);
and U23041 (N_23041,N_22948,N_22819);
or U23042 (N_23042,N_22632,N_22643);
and U23043 (N_23043,N_22967,N_22860);
nand U23044 (N_23044,N_22804,N_22744);
nand U23045 (N_23045,N_22761,N_22550);
and U23046 (N_23046,N_22941,N_22834);
or U23047 (N_23047,N_22976,N_22737);
nand U23048 (N_23048,N_22871,N_22720);
nand U23049 (N_23049,N_22881,N_22730);
or U23050 (N_23050,N_22699,N_22509);
nand U23051 (N_23051,N_22755,N_22919);
and U23052 (N_23052,N_22783,N_22855);
and U23053 (N_23053,N_22590,N_22866);
nor U23054 (N_23054,N_22561,N_22690);
or U23055 (N_23055,N_22527,N_22821);
nand U23056 (N_23056,N_22596,N_22525);
or U23057 (N_23057,N_22907,N_22987);
or U23058 (N_23058,N_22807,N_22933);
nand U23059 (N_23059,N_22845,N_22824);
xor U23060 (N_23060,N_22663,N_22532);
nand U23061 (N_23061,N_22626,N_22859);
or U23062 (N_23062,N_22902,N_22562);
nand U23063 (N_23063,N_22880,N_22642);
nand U23064 (N_23064,N_22865,N_22879);
nand U23065 (N_23065,N_22545,N_22557);
and U23066 (N_23066,N_22923,N_22659);
nand U23067 (N_23067,N_22612,N_22997);
nor U23068 (N_23068,N_22503,N_22813);
nand U23069 (N_23069,N_22507,N_22637);
or U23070 (N_23070,N_22799,N_22578);
or U23071 (N_23071,N_22617,N_22999);
nand U23072 (N_23072,N_22715,N_22805);
nand U23073 (N_23073,N_22544,N_22964);
and U23074 (N_23074,N_22966,N_22742);
nor U23075 (N_23075,N_22961,N_22739);
nor U23076 (N_23076,N_22521,N_22539);
nor U23077 (N_23077,N_22552,N_22897);
and U23078 (N_23078,N_22773,N_22806);
nor U23079 (N_23079,N_22767,N_22611);
xor U23080 (N_23080,N_22653,N_22770);
and U23081 (N_23081,N_22639,N_22660);
nor U23082 (N_23082,N_22713,N_22875);
or U23083 (N_23083,N_22702,N_22887);
and U23084 (N_23084,N_22908,N_22581);
or U23085 (N_23085,N_22597,N_22975);
nand U23086 (N_23086,N_22546,N_22533);
nor U23087 (N_23087,N_22502,N_22529);
nor U23088 (N_23088,N_22747,N_22709);
nand U23089 (N_23089,N_22683,N_22576);
and U23090 (N_23090,N_22517,N_22748);
or U23091 (N_23091,N_22842,N_22990);
xnor U23092 (N_23092,N_22672,N_22665);
and U23093 (N_23093,N_22832,N_22912);
nand U23094 (N_23094,N_22506,N_22993);
or U23095 (N_23095,N_22569,N_22974);
nor U23096 (N_23096,N_22869,N_22759);
or U23097 (N_23097,N_22695,N_22896);
and U23098 (N_23098,N_22678,N_22989);
nand U23099 (N_23099,N_22648,N_22756);
nand U23100 (N_23100,N_22853,N_22836);
or U23101 (N_23101,N_22820,N_22635);
and U23102 (N_23102,N_22803,N_22753);
and U23103 (N_23103,N_22850,N_22582);
nor U23104 (N_23104,N_22595,N_22684);
xor U23105 (N_23105,N_22681,N_22757);
xnor U23106 (N_23106,N_22852,N_22556);
nand U23107 (N_23107,N_22634,N_22627);
or U23108 (N_23108,N_22591,N_22536);
and U23109 (N_23109,N_22973,N_22548);
and U23110 (N_23110,N_22641,N_22570);
or U23111 (N_23111,N_22722,N_22559);
nor U23112 (N_23112,N_22861,N_22741);
or U23113 (N_23113,N_22796,N_22534);
nand U23114 (N_23114,N_22621,N_22929);
nor U23115 (N_23115,N_22687,N_22868);
or U23116 (N_23116,N_22558,N_22523);
and U23117 (N_23117,N_22873,N_22732);
or U23118 (N_23118,N_22724,N_22981);
nor U23119 (N_23119,N_22963,N_22790);
nand U23120 (N_23120,N_22631,N_22577);
nor U23121 (N_23121,N_22671,N_22656);
nand U23122 (N_23122,N_22554,N_22886);
nand U23123 (N_23123,N_22856,N_22679);
and U23124 (N_23124,N_22745,N_22945);
nand U23125 (N_23125,N_22943,N_22847);
or U23126 (N_23126,N_22782,N_22738);
or U23127 (N_23127,N_22851,N_22646);
nand U23128 (N_23128,N_22613,N_22700);
nor U23129 (N_23129,N_22827,N_22924);
and U23130 (N_23130,N_22760,N_22716);
and U23131 (N_23131,N_22694,N_22515);
nand U23132 (N_23132,N_22909,N_22616);
and U23133 (N_23133,N_22867,N_22547);
and U23134 (N_23134,N_22795,N_22901);
and U23135 (N_23135,N_22735,N_22995);
nand U23136 (N_23136,N_22727,N_22644);
nor U23137 (N_23137,N_22891,N_22607);
or U23138 (N_23138,N_22524,N_22543);
xnor U23139 (N_23139,N_22594,N_22844);
or U23140 (N_23140,N_22884,N_22704);
or U23141 (N_23141,N_22691,N_22991);
nor U23142 (N_23142,N_22752,N_22697);
xor U23143 (N_23143,N_22780,N_22531);
nor U23144 (N_23144,N_22958,N_22726);
nor U23145 (N_23145,N_22934,N_22636);
nor U23146 (N_23146,N_22876,N_22765);
nand U23147 (N_23147,N_22927,N_22588);
or U23148 (N_23148,N_22996,N_22888);
or U23149 (N_23149,N_22816,N_22586);
and U23150 (N_23150,N_22640,N_22937);
nor U23151 (N_23151,N_22516,N_22785);
and U23152 (N_23152,N_22980,N_22655);
nand U23153 (N_23153,N_22899,N_22826);
or U23154 (N_23154,N_22677,N_22668);
xor U23155 (N_23155,N_22654,N_22936);
nor U23156 (N_23156,N_22571,N_22921);
xnor U23157 (N_23157,N_22688,N_22540);
nand U23158 (N_23158,N_22956,N_22609);
nand U23159 (N_23159,N_22864,N_22601);
nand U23160 (N_23160,N_22802,N_22914);
nand U23161 (N_23161,N_22553,N_22686);
xor U23162 (N_23162,N_22736,N_22606);
nand U23163 (N_23163,N_22692,N_22822);
or U23164 (N_23164,N_22985,N_22815);
and U23165 (N_23165,N_22772,N_22918);
or U23166 (N_23166,N_22833,N_22817);
and U23167 (N_23167,N_22508,N_22728);
and U23168 (N_23168,N_22915,N_22589);
xor U23169 (N_23169,N_22751,N_22811);
nor U23170 (N_23170,N_22510,N_22743);
nor U23171 (N_23171,N_22818,N_22900);
and U23172 (N_23172,N_22955,N_22787);
and U23173 (N_23173,N_22746,N_22706);
nor U23174 (N_23174,N_22708,N_22954);
nor U23175 (N_23175,N_22638,N_22872);
or U23176 (N_23176,N_22673,N_22535);
nor U23177 (N_23177,N_22705,N_22874);
or U23178 (N_23178,N_22831,N_22784);
nor U23179 (N_23179,N_22960,N_22808);
xor U23180 (N_23180,N_22729,N_22733);
or U23181 (N_23181,N_22809,N_22689);
or U23182 (N_23182,N_22777,N_22779);
nor U23183 (N_23183,N_22717,N_22848);
nand U23184 (N_23184,N_22658,N_22501);
nand U23185 (N_23185,N_22837,N_22623);
and U23186 (N_23186,N_22555,N_22841);
nand U23187 (N_23187,N_22572,N_22549);
xor U23188 (N_23188,N_22696,N_22714);
nor U23189 (N_23189,N_22763,N_22749);
and U23190 (N_23190,N_22892,N_22986);
nand U23191 (N_23191,N_22711,N_22707);
or U23192 (N_23192,N_22953,N_22800);
nor U23193 (N_23193,N_22664,N_22505);
nand U23194 (N_23194,N_22628,N_22647);
nand U23195 (N_23195,N_22863,N_22946);
nand U23196 (N_23196,N_22858,N_22526);
and U23197 (N_23197,N_22575,N_22721);
nor U23198 (N_23198,N_22584,N_22843);
and U23199 (N_23199,N_22940,N_22764);
or U23200 (N_23200,N_22573,N_22723);
nor U23201 (N_23201,N_22932,N_22938);
xnor U23202 (N_23202,N_22894,N_22719);
nor U23203 (N_23203,N_22537,N_22906);
and U23204 (N_23204,N_22878,N_22977);
and U23205 (N_23205,N_22703,N_22580);
or U23206 (N_23206,N_22984,N_22935);
or U23207 (N_23207,N_22846,N_22625);
nand U23208 (N_23208,N_22669,N_22551);
or U23209 (N_23209,N_22916,N_22792);
and U23210 (N_23210,N_22566,N_22965);
nor U23211 (N_23211,N_22560,N_22712);
and U23212 (N_23212,N_22528,N_22791);
and U23213 (N_23213,N_22978,N_22750);
nand U23214 (N_23214,N_22905,N_22541);
nand U23215 (N_23215,N_22758,N_22994);
and U23216 (N_23216,N_22564,N_22512);
and U23217 (N_23217,N_22513,N_22798);
or U23218 (N_23218,N_22789,N_22538);
nor U23219 (N_23219,N_22950,N_22962);
nor U23220 (N_23220,N_22518,N_22839);
and U23221 (N_23221,N_22928,N_22766);
nor U23222 (N_23222,N_22542,N_22775);
and U23223 (N_23223,N_22579,N_22567);
xor U23224 (N_23224,N_22988,N_22947);
or U23225 (N_23225,N_22500,N_22952);
or U23226 (N_23226,N_22734,N_22670);
nand U23227 (N_23227,N_22825,N_22718);
nor U23228 (N_23228,N_22951,N_22925);
or U23229 (N_23229,N_22931,N_22970);
and U23230 (N_23230,N_22605,N_22522);
and U23231 (N_23231,N_22676,N_22599);
or U23232 (N_23232,N_22598,N_22801);
and U23233 (N_23233,N_22614,N_22903);
nand U23234 (N_23234,N_22511,N_22762);
nor U23235 (N_23235,N_22778,N_22849);
or U23236 (N_23236,N_22911,N_22520);
and U23237 (N_23237,N_22725,N_22857);
or U23238 (N_23238,N_22604,N_22776);
or U23239 (N_23239,N_22920,N_22624);
nor U23240 (N_23240,N_22682,N_22883);
xor U23241 (N_23241,N_22649,N_22922);
nor U23242 (N_23242,N_22983,N_22898);
nand U23243 (N_23243,N_22568,N_22619);
or U23244 (N_23244,N_22971,N_22774);
or U23245 (N_23245,N_22893,N_22904);
nand U23246 (N_23246,N_22731,N_22829);
and U23247 (N_23247,N_22698,N_22629);
or U23248 (N_23248,N_22740,N_22610);
or U23249 (N_23249,N_22840,N_22939);
xnor U23250 (N_23250,N_22945,N_22901);
or U23251 (N_23251,N_22753,N_22899);
nand U23252 (N_23252,N_22565,N_22941);
nand U23253 (N_23253,N_22648,N_22802);
nand U23254 (N_23254,N_22658,N_22516);
or U23255 (N_23255,N_22951,N_22883);
nor U23256 (N_23256,N_22670,N_22601);
or U23257 (N_23257,N_22694,N_22693);
and U23258 (N_23258,N_22820,N_22577);
nand U23259 (N_23259,N_22718,N_22557);
nand U23260 (N_23260,N_22699,N_22566);
or U23261 (N_23261,N_22954,N_22966);
nand U23262 (N_23262,N_22652,N_22965);
and U23263 (N_23263,N_22532,N_22909);
and U23264 (N_23264,N_22726,N_22874);
and U23265 (N_23265,N_22651,N_22843);
xnor U23266 (N_23266,N_22539,N_22983);
or U23267 (N_23267,N_22987,N_22533);
and U23268 (N_23268,N_22630,N_22860);
and U23269 (N_23269,N_22942,N_22816);
or U23270 (N_23270,N_22991,N_22723);
or U23271 (N_23271,N_22546,N_22959);
and U23272 (N_23272,N_22648,N_22538);
and U23273 (N_23273,N_22969,N_22533);
nand U23274 (N_23274,N_22865,N_22759);
nor U23275 (N_23275,N_22600,N_22841);
and U23276 (N_23276,N_22730,N_22719);
nor U23277 (N_23277,N_22927,N_22839);
and U23278 (N_23278,N_22534,N_22949);
nand U23279 (N_23279,N_22799,N_22796);
or U23280 (N_23280,N_22766,N_22569);
nand U23281 (N_23281,N_22749,N_22969);
nor U23282 (N_23282,N_22656,N_22838);
or U23283 (N_23283,N_22551,N_22859);
nor U23284 (N_23284,N_22534,N_22889);
nor U23285 (N_23285,N_22566,N_22743);
nor U23286 (N_23286,N_22572,N_22795);
nor U23287 (N_23287,N_22651,N_22913);
and U23288 (N_23288,N_22902,N_22740);
or U23289 (N_23289,N_22662,N_22911);
or U23290 (N_23290,N_22569,N_22968);
nand U23291 (N_23291,N_22529,N_22672);
or U23292 (N_23292,N_22827,N_22660);
xnor U23293 (N_23293,N_22990,N_22943);
xnor U23294 (N_23294,N_22729,N_22860);
nor U23295 (N_23295,N_22772,N_22781);
nand U23296 (N_23296,N_22524,N_22790);
and U23297 (N_23297,N_22788,N_22806);
xnor U23298 (N_23298,N_22770,N_22649);
and U23299 (N_23299,N_22981,N_22526);
nand U23300 (N_23300,N_22898,N_22673);
nor U23301 (N_23301,N_22553,N_22801);
nand U23302 (N_23302,N_22716,N_22814);
and U23303 (N_23303,N_22592,N_22678);
and U23304 (N_23304,N_22820,N_22547);
and U23305 (N_23305,N_22510,N_22502);
nor U23306 (N_23306,N_22892,N_22862);
or U23307 (N_23307,N_22935,N_22994);
and U23308 (N_23308,N_22555,N_22913);
nand U23309 (N_23309,N_22981,N_22794);
nand U23310 (N_23310,N_22740,N_22934);
and U23311 (N_23311,N_22718,N_22748);
nand U23312 (N_23312,N_22787,N_22730);
nand U23313 (N_23313,N_22755,N_22944);
nand U23314 (N_23314,N_22998,N_22760);
nor U23315 (N_23315,N_22900,N_22527);
or U23316 (N_23316,N_22564,N_22519);
or U23317 (N_23317,N_22724,N_22951);
xnor U23318 (N_23318,N_22945,N_22651);
nand U23319 (N_23319,N_22543,N_22998);
or U23320 (N_23320,N_22704,N_22995);
xor U23321 (N_23321,N_22573,N_22920);
nand U23322 (N_23322,N_22838,N_22650);
or U23323 (N_23323,N_22592,N_22914);
or U23324 (N_23324,N_22800,N_22652);
nor U23325 (N_23325,N_22837,N_22675);
or U23326 (N_23326,N_22649,N_22572);
xnor U23327 (N_23327,N_22590,N_22740);
and U23328 (N_23328,N_22946,N_22818);
or U23329 (N_23329,N_22829,N_22582);
nand U23330 (N_23330,N_22741,N_22945);
nor U23331 (N_23331,N_22718,N_22826);
or U23332 (N_23332,N_22995,N_22703);
nand U23333 (N_23333,N_22692,N_22518);
and U23334 (N_23334,N_22606,N_22697);
nor U23335 (N_23335,N_22861,N_22733);
nor U23336 (N_23336,N_22936,N_22849);
or U23337 (N_23337,N_22997,N_22787);
nor U23338 (N_23338,N_22557,N_22500);
or U23339 (N_23339,N_22915,N_22789);
nor U23340 (N_23340,N_22532,N_22830);
nand U23341 (N_23341,N_22539,N_22956);
nand U23342 (N_23342,N_22778,N_22920);
and U23343 (N_23343,N_22523,N_22560);
or U23344 (N_23344,N_22679,N_22665);
nor U23345 (N_23345,N_22576,N_22592);
or U23346 (N_23346,N_22565,N_22674);
nand U23347 (N_23347,N_22999,N_22780);
nand U23348 (N_23348,N_22922,N_22972);
nand U23349 (N_23349,N_22510,N_22675);
nor U23350 (N_23350,N_22912,N_22933);
and U23351 (N_23351,N_22954,N_22813);
nand U23352 (N_23352,N_22878,N_22979);
and U23353 (N_23353,N_22871,N_22783);
nor U23354 (N_23354,N_22907,N_22644);
or U23355 (N_23355,N_22715,N_22683);
or U23356 (N_23356,N_22516,N_22717);
and U23357 (N_23357,N_22809,N_22835);
nand U23358 (N_23358,N_22842,N_22798);
or U23359 (N_23359,N_22861,N_22691);
and U23360 (N_23360,N_22861,N_22878);
or U23361 (N_23361,N_22548,N_22717);
and U23362 (N_23362,N_22850,N_22912);
nand U23363 (N_23363,N_22818,N_22597);
and U23364 (N_23364,N_22814,N_22997);
nor U23365 (N_23365,N_22878,N_22881);
nor U23366 (N_23366,N_22511,N_22971);
nand U23367 (N_23367,N_22603,N_22818);
nand U23368 (N_23368,N_22938,N_22870);
and U23369 (N_23369,N_22613,N_22541);
nor U23370 (N_23370,N_22697,N_22957);
nand U23371 (N_23371,N_22974,N_22815);
xnor U23372 (N_23372,N_22833,N_22903);
nor U23373 (N_23373,N_22918,N_22929);
and U23374 (N_23374,N_22899,N_22940);
xnor U23375 (N_23375,N_22875,N_22991);
nor U23376 (N_23376,N_22963,N_22755);
or U23377 (N_23377,N_22847,N_22675);
nand U23378 (N_23378,N_22572,N_22906);
and U23379 (N_23379,N_22745,N_22539);
nor U23380 (N_23380,N_22789,N_22661);
and U23381 (N_23381,N_22607,N_22987);
xnor U23382 (N_23382,N_22941,N_22966);
nor U23383 (N_23383,N_22868,N_22616);
or U23384 (N_23384,N_22841,N_22709);
or U23385 (N_23385,N_22676,N_22967);
nor U23386 (N_23386,N_22712,N_22979);
and U23387 (N_23387,N_22568,N_22997);
xnor U23388 (N_23388,N_22529,N_22991);
nor U23389 (N_23389,N_22739,N_22513);
or U23390 (N_23390,N_22719,N_22542);
nor U23391 (N_23391,N_22778,N_22758);
nand U23392 (N_23392,N_22602,N_22646);
xnor U23393 (N_23393,N_22679,N_22966);
or U23394 (N_23394,N_22939,N_22847);
nand U23395 (N_23395,N_22975,N_22963);
and U23396 (N_23396,N_22973,N_22840);
or U23397 (N_23397,N_22693,N_22573);
and U23398 (N_23398,N_22910,N_22693);
or U23399 (N_23399,N_22932,N_22841);
and U23400 (N_23400,N_22667,N_22673);
or U23401 (N_23401,N_22864,N_22648);
nand U23402 (N_23402,N_22673,N_22850);
xor U23403 (N_23403,N_22723,N_22629);
and U23404 (N_23404,N_22851,N_22578);
nand U23405 (N_23405,N_22818,N_22691);
and U23406 (N_23406,N_22849,N_22581);
or U23407 (N_23407,N_22859,N_22964);
or U23408 (N_23408,N_22846,N_22811);
and U23409 (N_23409,N_22969,N_22912);
and U23410 (N_23410,N_22582,N_22572);
nand U23411 (N_23411,N_22873,N_22680);
and U23412 (N_23412,N_22942,N_22989);
nand U23413 (N_23413,N_22930,N_22956);
or U23414 (N_23414,N_22695,N_22693);
or U23415 (N_23415,N_22511,N_22752);
nand U23416 (N_23416,N_22591,N_22593);
or U23417 (N_23417,N_22871,N_22917);
xor U23418 (N_23418,N_22719,N_22993);
or U23419 (N_23419,N_22523,N_22590);
or U23420 (N_23420,N_22642,N_22997);
nor U23421 (N_23421,N_22889,N_22857);
or U23422 (N_23422,N_22930,N_22544);
or U23423 (N_23423,N_22831,N_22600);
and U23424 (N_23424,N_22639,N_22848);
and U23425 (N_23425,N_22917,N_22815);
nand U23426 (N_23426,N_22586,N_22883);
and U23427 (N_23427,N_22504,N_22849);
nor U23428 (N_23428,N_22583,N_22967);
nand U23429 (N_23429,N_22698,N_22631);
xnor U23430 (N_23430,N_22875,N_22719);
and U23431 (N_23431,N_22580,N_22603);
nand U23432 (N_23432,N_22566,N_22955);
nor U23433 (N_23433,N_22923,N_22866);
or U23434 (N_23434,N_22619,N_22878);
and U23435 (N_23435,N_22799,N_22808);
nand U23436 (N_23436,N_22823,N_22747);
or U23437 (N_23437,N_22659,N_22865);
nor U23438 (N_23438,N_22800,N_22656);
nand U23439 (N_23439,N_22858,N_22504);
nor U23440 (N_23440,N_22910,N_22730);
and U23441 (N_23441,N_22730,N_22836);
and U23442 (N_23442,N_22528,N_22862);
nand U23443 (N_23443,N_22874,N_22928);
and U23444 (N_23444,N_22638,N_22613);
nand U23445 (N_23445,N_22878,N_22800);
xor U23446 (N_23446,N_22882,N_22697);
or U23447 (N_23447,N_22514,N_22962);
nor U23448 (N_23448,N_22580,N_22838);
nand U23449 (N_23449,N_22626,N_22511);
nor U23450 (N_23450,N_22964,N_22806);
and U23451 (N_23451,N_22501,N_22893);
or U23452 (N_23452,N_22608,N_22937);
or U23453 (N_23453,N_22945,N_22916);
nand U23454 (N_23454,N_22566,N_22501);
nor U23455 (N_23455,N_22752,N_22611);
nor U23456 (N_23456,N_22625,N_22920);
nand U23457 (N_23457,N_22534,N_22813);
or U23458 (N_23458,N_22529,N_22807);
xnor U23459 (N_23459,N_22548,N_22774);
nor U23460 (N_23460,N_22923,N_22532);
xnor U23461 (N_23461,N_22727,N_22559);
and U23462 (N_23462,N_22513,N_22668);
nor U23463 (N_23463,N_22560,N_22658);
or U23464 (N_23464,N_22529,N_22694);
or U23465 (N_23465,N_22804,N_22943);
nor U23466 (N_23466,N_22720,N_22805);
and U23467 (N_23467,N_22712,N_22728);
and U23468 (N_23468,N_22845,N_22832);
nor U23469 (N_23469,N_22568,N_22618);
and U23470 (N_23470,N_22735,N_22520);
or U23471 (N_23471,N_22632,N_22541);
and U23472 (N_23472,N_22545,N_22869);
nand U23473 (N_23473,N_22590,N_22827);
xor U23474 (N_23474,N_22861,N_22975);
or U23475 (N_23475,N_22642,N_22627);
and U23476 (N_23476,N_22615,N_22914);
nor U23477 (N_23477,N_22549,N_22938);
nand U23478 (N_23478,N_22748,N_22849);
nand U23479 (N_23479,N_22975,N_22961);
and U23480 (N_23480,N_22611,N_22801);
nor U23481 (N_23481,N_22606,N_22649);
nor U23482 (N_23482,N_22682,N_22894);
nor U23483 (N_23483,N_22633,N_22559);
or U23484 (N_23484,N_22768,N_22913);
nand U23485 (N_23485,N_22598,N_22704);
nand U23486 (N_23486,N_22638,N_22888);
or U23487 (N_23487,N_22858,N_22817);
and U23488 (N_23488,N_22731,N_22535);
or U23489 (N_23489,N_22947,N_22933);
and U23490 (N_23490,N_22852,N_22893);
nand U23491 (N_23491,N_22768,N_22675);
or U23492 (N_23492,N_22727,N_22696);
or U23493 (N_23493,N_22606,N_22810);
or U23494 (N_23494,N_22898,N_22900);
nand U23495 (N_23495,N_22579,N_22533);
nand U23496 (N_23496,N_22778,N_22648);
or U23497 (N_23497,N_22750,N_22634);
nor U23498 (N_23498,N_22600,N_22842);
and U23499 (N_23499,N_22920,N_22563);
or U23500 (N_23500,N_23345,N_23140);
and U23501 (N_23501,N_23082,N_23486);
or U23502 (N_23502,N_23045,N_23438);
xor U23503 (N_23503,N_23297,N_23404);
nand U23504 (N_23504,N_23236,N_23325);
xor U23505 (N_23505,N_23303,N_23180);
nor U23506 (N_23506,N_23068,N_23284);
xor U23507 (N_23507,N_23204,N_23454);
or U23508 (N_23508,N_23427,N_23280);
nand U23509 (N_23509,N_23027,N_23176);
nor U23510 (N_23510,N_23447,N_23205);
nand U23511 (N_23511,N_23375,N_23075);
and U23512 (N_23512,N_23042,N_23200);
and U23513 (N_23513,N_23097,N_23124);
and U23514 (N_23514,N_23465,N_23321);
nand U23515 (N_23515,N_23142,N_23386);
nand U23516 (N_23516,N_23395,N_23247);
nor U23517 (N_23517,N_23195,N_23231);
nand U23518 (N_23518,N_23130,N_23253);
nor U23519 (N_23519,N_23213,N_23431);
xnor U23520 (N_23520,N_23352,N_23248);
nor U23521 (N_23521,N_23324,N_23105);
nor U23522 (N_23522,N_23242,N_23376);
and U23523 (N_23523,N_23363,N_23432);
nand U23524 (N_23524,N_23466,N_23311);
nor U23525 (N_23525,N_23008,N_23058);
nor U23526 (N_23526,N_23216,N_23127);
and U23527 (N_23527,N_23353,N_23011);
nand U23528 (N_23528,N_23148,N_23425);
and U23529 (N_23529,N_23040,N_23138);
nor U23530 (N_23530,N_23418,N_23389);
xnor U23531 (N_23531,N_23146,N_23391);
and U23532 (N_23532,N_23181,N_23147);
or U23533 (N_23533,N_23250,N_23167);
and U23534 (N_23534,N_23026,N_23372);
or U23535 (N_23535,N_23339,N_23110);
nand U23536 (N_23536,N_23090,N_23334);
and U23537 (N_23537,N_23212,N_23174);
or U23538 (N_23538,N_23330,N_23197);
xnor U23539 (N_23539,N_23349,N_23051);
and U23540 (N_23540,N_23478,N_23215);
nand U23541 (N_23541,N_23202,N_23073);
nor U23542 (N_23542,N_23217,N_23368);
and U23543 (N_23543,N_23166,N_23235);
or U23544 (N_23544,N_23393,N_23317);
nor U23545 (N_23545,N_23054,N_23310);
or U23546 (N_23546,N_23239,N_23126);
nand U23547 (N_23547,N_23025,N_23357);
or U23548 (N_23548,N_23149,N_23030);
or U23549 (N_23549,N_23228,N_23063);
xnor U23550 (N_23550,N_23112,N_23044);
or U23551 (N_23551,N_23493,N_23116);
or U23552 (N_23552,N_23219,N_23473);
nand U23553 (N_23553,N_23207,N_23012);
nand U23554 (N_23554,N_23154,N_23115);
or U23555 (N_23555,N_23382,N_23492);
or U23556 (N_23556,N_23244,N_23078);
and U23557 (N_23557,N_23067,N_23323);
nor U23558 (N_23558,N_23491,N_23394);
or U23559 (N_23559,N_23169,N_23144);
nor U23560 (N_23560,N_23000,N_23245);
nor U23561 (N_23561,N_23287,N_23364);
and U23562 (N_23562,N_23413,N_23064);
or U23563 (N_23563,N_23428,N_23240);
nor U23564 (N_23564,N_23306,N_23016);
xnor U23565 (N_23565,N_23269,N_23474);
and U23566 (N_23566,N_23390,N_23275);
nand U23567 (N_23567,N_23225,N_23077);
or U23568 (N_23568,N_23259,N_23336);
or U23569 (N_23569,N_23398,N_23256);
xor U23570 (N_23570,N_23238,N_23283);
nand U23571 (N_23571,N_23496,N_23276);
or U23572 (N_23572,N_23094,N_23308);
nand U23573 (N_23573,N_23302,N_23305);
nand U23574 (N_23574,N_23237,N_23013);
or U23575 (N_23575,N_23423,N_23314);
or U23576 (N_23576,N_23251,N_23331);
xor U23577 (N_23577,N_23446,N_23087);
or U23578 (N_23578,N_23233,N_23103);
nor U23579 (N_23579,N_23318,N_23189);
nand U23580 (N_23580,N_23348,N_23161);
xnor U23581 (N_23581,N_23397,N_23488);
or U23582 (N_23582,N_23299,N_23050);
nor U23583 (N_23583,N_23028,N_23241);
and U23584 (N_23584,N_23053,N_23261);
nor U23585 (N_23585,N_23358,N_23270);
nor U23586 (N_23586,N_23227,N_23162);
or U23587 (N_23587,N_23484,N_23074);
nand U23588 (N_23588,N_23069,N_23182);
nand U23589 (N_23589,N_23257,N_23096);
or U23590 (N_23590,N_23439,N_23156);
or U23591 (N_23591,N_23265,N_23246);
nand U23592 (N_23592,N_23288,N_23313);
nor U23593 (N_23593,N_23414,N_23099);
nand U23594 (N_23594,N_23061,N_23095);
nor U23595 (N_23595,N_23354,N_23185);
and U23596 (N_23596,N_23290,N_23059);
or U23597 (N_23597,N_23224,N_23274);
or U23598 (N_23598,N_23433,N_23281);
nor U23599 (N_23599,N_23415,N_23451);
xnor U23600 (N_23600,N_23469,N_23495);
nor U23601 (N_23601,N_23457,N_23379);
xnor U23602 (N_23602,N_23029,N_23483);
or U23603 (N_23603,N_23186,N_23043);
and U23604 (N_23604,N_23378,N_23192);
nor U23605 (N_23605,N_23340,N_23292);
or U23606 (N_23606,N_23383,N_23183);
and U23607 (N_23607,N_23020,N_23429);
nor U23608 (N_23608,N_23137,N_23410);
nor U23609 (N_23609,N_23472,N_23201);
and U23610 (N_23610,N_23412,N_23009);
nor U23611 (N_23611,N_23065,N_23057);
or U23612 (N_23612,N_23362,N_23396);
or U23613 (N_23613,N_23298,N_23448);
and U23614 (N_23614,N_23335,N_23277);
nand U23615 (N_23615,N_23464,N_23490);
nand U23616 (N_23616,N_23271,N_23262);
or U23617 (N_23617,N_23449,N_23480);
or U23618 (N_23618,N_23080,N_23346);
nor U23619 (N_23619,N_23135,N_23199);
nor U23620 (N_23620,N_23089,N_23350);
or U23621 (N_23621,N_23360,N_23121);
nand U23622 (N_23622,N_23377,N_23252);
nand U23623 (N_23623,N_23499,N_23341);
nor U23624 (N_23624,N_23031,N_23255);
xnor U23625 (N_23625,N_23343,N_23155);
or U23626 (N_23626,N_23408,N_23017);
nand U23627 (N_23627,N_23208,N_23304);
or U23628 (N_23628,N_23037,N_23387);
or U23629 (N_23629,N_23014,N_23307);
xnor U23630 (N_23630,N_23436,N_23264);
or U23631 (N_23631,N_23039,N_23487);
and U23632 (N_23632,N_23459,N_23111);
nand U23633 (N_23633,N_23294,N_23400);
or U23634 (N_23634,N_23134,N_23117);
and U23635 (N_23635,N_23165,N_23093);
xor U23636 (N_23636,N_23402,N_23467);
nand U23637 (N_23637,N_23361,N_23158);
nand U23638 (N_23638,N_23079,N_23461);
or U23639 (N_23639,N_23273,N_23211);
and U23640 (N_23640,N_23254,N_23196);
and U23641 (N_23641,N_23356,N_23295);
and U23642 (N_23642,N_23108,N_23392);
nand U23643 (N_23643,N_23033,N_23032);
or U23644 (N_23644,N_23084,N_23128);
nor U23645 (N_23645,N_23114,N_23430);
xor U23646 (N_23646,N_23190,N_23132);
nor U23647 (N_23647,N_23036,N_23417);
xor U23648 (N_23648,N_23316,N_23046);
and U23649 (N_23649,N_23333,N_23312);
and U23650 (N_23650,N_23076,N_23326);
nand U23651 (N_23651,N_23191,N_23049);
and U23652 (N_23652,N_23102,N_23218);
and U23653 (N_23653,N_23088,N_23047);
or U23654 (N_23654,N_23293,N_23230);
nor U23655 (N_23655,N_23381,N_23437);
nor U23656 (N_23656,N_23133,N_23003);
xnor U23657 (N_23657,N_23267,N_23206);
nand U23658 (N_23658,N_23403,N_23416);
and U23659 (N_23659,N_23214,N_23220);
or U23660 (N_23660,N_23405,N_23258);
or U23661 (N_23661,N_23101,N_23193);
and U23662 (N_23662,N_23409,N_23388);
nor U23663 (N_23663,N_23477,N_23272);
or U23664 (N_23664,N_23151,N_23419);
and U23665 (N_23665,N_23401,N_23260);
nor U23666 (N_23666,N_23022,N_23291);
xor U23667 (N_23667,N_23475,N_23249);
nand U23668 (N_23668,N_23263,N_23476);
nand U23669 (N_23669,N_23052,N_23406);
nor U23670 (N_23670,N_23168,N_23048);
or U23671 (N_23671,N_23010,N_23315);
nand U23672 (N_23672,N_23226,N_23329);
nor U23673 (N_23673,N_23374,N_23482);
nor U23674 (N_23674,N_23434,N_23422);
and U23675 (N_23675,N_23091,N_23184);
nor U23676 (N_23676,N_23344,N_23479);
or U23677 (N_23677,N_23136,N_23083);
xnor U23678 (N_23678,N_23494,N_23285);
and U23679 (N_23679,N_23489,N_23453);
and U23680 (N_23680,N_23018,N_23178);
nor U23681 (N_23681,N_23337,N_23034);
xnor U23682 (N_23682,N_23369,N_23107);
or U23683 (N_23683,N_23462,N_23384);
and U23684 (N_23684,N_23232,N_23229);
or U23685 (N_23685,N_23266,N_23380);
nor U23686 (N_23686,N_23152,N_23468);
nand U23687 (N_23687,N_23443,N_23338);
nor U23688 (N_23688,N_23385,N_23159);
nand U23689 (N_23689,N_23024,N_23035);
nand U23690 (N_23690,N_23481,N_23268);
and U23691 (N_23691,N_23188,N_23163);
or U23692 (N_23692,N_23455,N_23460);
or U23693 (N_23693,N_23056,N_23109);
nor U23694 (N_23694,N_23426,N_23435);
and U23695 (N_23695,N_23203,N_23210);
nand U23696 (N_23696,N_23309,N_23004);
nand U23697 (N_23697,N_23119,N_23153);
or U23698 (N_23698,N_23365,N_23407);
nor U23699 (N_23699,N_23062,N_23015);
nor U23700 (N_23700,N_23145,N_23021);
and U23701 (N_23701,N_23296,N_23150);
or U23702 (N_23702,N_23002,N_23289);
or U23703 (N_23703,N_23320,N_23005);
or U23704 (N_23704,N_23143,N_23243);
nand U23705 (N_23705,N_23023,N_23399);
or U23706 (N_23706,N_23006,N_23209);
or U23707 (N_23707,N_23328,N_23171);
or U23708 (N_23708,N_23129,N_23113);
nand U23709 (N_23709,N_23411,N_23450);
nand U23710 (N_23710,N_23282,N_23498);
and U23711 (N_23711,N_23444,N_23139);
or U23712 (N_23712,N_23098,N_23198);
or U23713 (N_23713,N_23187,N_23071);
and U23714 (N_23714,N_23007,N_23179);
xor U23715 (N_23715,N_23001,N_23223);
and U23716 (N_23716,N_23445,N_23458);
nand U23717 (N_23717,N_23327,N_23452);
nor U23718 (N_23718,N_23038,N_23279);
nand U23719 (N_23719,N_23359,N_23070);
and U23720 (N_23720,N_23222,N_23485);
and U23721 (N_23721,N_23278,N_23351);
nor U23722 (N_23722,N_23471,N_23300);
and U23723 (N_23723,N_23173,N_23104);
and U23724 (N_23724,N_23131,N_23157);
or U23725 (N_23725,N_23440,N_23081);
nand U23726 (N_23726,N_23055,N_23319);
nor U23727 (N_23727,N_23322,N_23194);
nor U23728 (N_23728,N_23092,N_23177);
nand U23729 (N_23729,N_23123,N_23085);
nor U23730 (N_23730,N_23370,N_23332);
nor U23731 (N_23731,N_23066,N_23421);
nand U23732 (N_23732,N_23342,N_23367);
xor U23733 (N_23733,N_23234,N_23086);
and U23734 (N_23734,N_23355,N_23072);
nor U23735 (N_23735,N_23366,N_23221);
or U23736 (N_23736,N_23060,N_23286);
and U23737 (N_23737,N_23301,N_23463);
nand U23738 (N_23738,N_23456,N_23122);
nor U23739 (N_23739,N_23041,N_23442);
nand U23740 (N_23740,N_23470,N_23175);
nand U23741 (N_23741,N_23118,N_23373);
and U23742 (N_23742,N_23441,N_23371);
nor U23743 (N_23743,N_23120,N_23100);
nor U23744 (N_23744,N_23497,N_23164);
nor U23745 (N_23745,N_23125,N_23172);
nand U23746 (N_23746,N_23424,N_23170);
nor U23747 (N_23747,N_23160,N_23420);
nand U23748 (N_23748,N_23141,N_23106);
nand U23749 (N_23749,N_23019,N_23347);
nor U23750 (N_23750,N_23168,N_23469);
xor U23751 (N_23751,N_23103,N_23195);
nor U23752 (N_23752,N_23114,N_23248);
and U23753 (N_23753,N_23103,N_23172);
or U23754 (N_23754,N_23471,N_23228);
nand U23755 (N_23755,N_23175,N_23282);
and U23756 (N_23756,N_23079,N_23382);
nor U23757 (N_23757,N_23057,N_23015);
nand U23758 (N_23758,N_23403,N_23026);
or U23759 (N_23759,N_23310,N_23274);
nor U23760 (N_23760,N_23317,N_23316);
xor U23761 (N_23761,N_23152,N_23284);
nand U23762 (N_23762,N_23145,N_23471);
or U23763 (N_23763,N_23128,N_23098);
xnor U23764 (N_23764,N_23238,N_23285);
or U23765 (N_23765,N_23073,N_23437);
and U23766 (N_23766,N_23499,N_23290);
nand U23767 (N_23767,N_23064,N_23127);
xor U23768 (N_23768,N_23294,N_23415);
nand U23769 (N_23769,N_23205,N_23089);
nand U23770 (N_23770,N_23466,N_23008);
and U23771 (N_23771,N_23096,N_23225);
and U23772 (N_23772,N_23223,N_23013);
nand U23773 (N_23773,N_23486,N_23421);
or U23774 (N_23774,N_23377,N_23135);
nor U23775 (N_23775,N_23148,N_23121);
nor U23776 (N_23776,N_23118,N_23032);
or U23777 (N_23777,N_23150,N_23289);
and U23778 (N_23778,N_23281,N_23247);
xnor U23779 (N_23779,N_23063,N_23350);
and U23780 (N_23780,N_23142,N_23411);
nor U23781 (N_23781,N_23347,N_23472);
nor U23782 (N_23782,N_23293,N_23324);
nand U23783 (N_23783,N_23119,N_23138);
and U23784 (N_23784,N_23469,N_23170);
and U23785 (N_23785,N_23341,N_23287);
or U23786 (N_23786,N_23172,N_23332);
nand U23787 (N_23787,N_23093,N_23429);
or U23788 (N_23788,N_23187,N_23017);
or U23789 (N_23789,N_23154,N_23392);
nand U23790 (N_23790,N_23293,N_23023);
nand U23791 (N_23791,N_23193,N_23329);
nor U23792 (N_23792,N_23176,N_23280);
nand U23793 (N_23793,N_23307,N_23183);
and U23794 (N_23794,N_23280,N_23033);
and U23795 (N_23795,N_23031,N_23017);
nor U23796 (N_23796,N_23211,N_23411);
and U23797 (N_23797,N_23363,N_23469);
xnor U23798 (N_23798,N_23391,N_23145);
or U23799 (N_23799,N_23040,N_23214);
nor U23800 (N_23800,N_23028,N_23102);
nor U23801 (N_23801,N_23467,N_23415);
or U23802 (N_23802,N_23364,N_23124);
nand U23803 (N_23803,N_23370,N_23167);
and U23804 (N_23804,N_23011,N_23208);
and U23805 (N_23805,N_23106,N_23012);
and U23806 (N_23806,N_23256,N_23060);
or U23807 (N_23807,N_23138,N_23221);
nand U23808 (N_23808,N_23095,N_23357);
and U23809 (N_23809,N_23226,N_23183);
nand U23810 (N_23810,N_23123,N_23048);
nand U23811 (N_23811,N_23275,N_23322);
nor U23812 (N_23812,N_23239,N_23161);
or U23813 (N_23813,N_23053,N_23112);
nand U23814 (N_23814,N_23326,N_23456);
and U23815 (N_23815,N_23386,N_23084);
nor U23816 (N_23816,N_23295,N_23037);
or U23817 (N_23817,N_23471,N_23097);
nand U23818 (N_23818,N_23296,N_23042);
nand U23819 (N_23819,N_23336,N_23342);
nor U23820 (N_23820,N_23431,N_23404);
nor U23821 (N_23821,N_23485,N_23168);
and U23822 (N_23822,N_23007,N_23313);
nand U23823 (N_23823,N_23089,N_23375);
and U23824 (N_23824,N_23276,N_23383);
nand U23825 (N_23825,N_23406,N_23412);
or U23826 (N_23826,N_23091,N_23149);
nand U23827 (N_23827,N_23437,N_23472);
xnor U23828 (N_23828,N_23132,N_23467);
and U23829 (N_23829,N_23312,N_23299);
and U23830 (N_23830,N_23193,N_23166);
and U23831 (N_23831,N_23125,N_23261);
or U23832 (N_23832,N_23475,N_23162);
or U23833 (N_23833,N_23369,N_23255);
nor U23834 (N_23834,N_23173,N_23279);
nor U23835 (N_23835,N_23076,N_23112);
nand U23836 (N_23836,N_23374,N_23023);
or U23837 (N_23837,N_23429,N_23098);
nor U23838 (N_23838,N_23094,N_23164);
or U23839 (N_23839,N_23322,N_23226);
and U23840 (N_23840,N_23214,N_23458);
or U23841 (N_23841,N_23160,N_23347);
and U23842 (N_23842,N_23432,N_23310);
xor U23843 (N_23843,N_23105,N_23392);
and U23844 (N_23844,N_23023,N_23178);
and U23845 (N_23845,N_23078,N_23290);
or U23846 (N_23846,N_23260,N_23413);
and U23847 (N_23847,N_23219,N_23000);
and U23848 (N_23848,N_23420,N_23493);
nand U23849 (N_23849,N_23118,N_23405);
xor U23850 (N_23850,N_23030,N_23246);
nor U23851 (N_23851,N_23189,N_23479);
and U23852 (N_23852,N_23304,N_23453);
nor U23853 (N_23853,N_23110,N_23072);
nor U23854 (N_23854,N_23419,N_23200);
xnor U23855 (N_23855,N_23102,N_23410);
xnor U23856 (N_23856,N_23445,N_23009);
and U23857 (N_23857,N_23393,N_23032);
or U23858 (N_23858,N_23486,N_23442);
nand U23859 (N_23859,N_23267,N_23040);
nand U23860 (N_23860,N_23288,N_23437);
or U23861 (N_23861,N_23012,N_23031);
and U23862 (N_23862,N_23319,N_23422);
or U23863 (N_23863,N_23359,N_23080);
xor U23864 (N_23864,N_23205,N_23046);
or U23865 (N_23865,N_23430,N_23283);
and U23866 (N_23866,N_23354,N_23118);
nor U23867 (N_23867,N_23232,N_23090);
or U23868 (N_23868,N_23015,N_23300);
and U23869 (N_23869,N_23182,N_23269);
nor U23870 (N_23870,N_23166,N_23427);
and U23871 (N_23871,N_23311,N_23204);
nor U23872 (N_23872,N_23157,N_23348);
or U23873 (N_23873,N_23258,N_23423);
and U23874 (N_23874,N_23427,N_23336);
nand U23875 (N_23875,N_23492,N_23079);
nor U23876 (N_23876,N_23007,N_23207);
and U23877 (N_23877,N_23171,N_23059);
nand U23878 (N_23878,N_23468,N_23317);
and U23879 (N_23879,N_23096,N_23460);
and U23880 (N_23880,N_23347,N_23310);
nand U23881 (N_23881,N_23128,N_23100);
and U23882 (N_23882,N_23349,N_23302);
nor U23883 (N_23883,N_23428,N_23140);
nor U23884 (N_23884,N_23470,N_23437);
or U23885 (N_23885,N_23482,N_23158);
and U23886 (N_23886,N_23158,N_23484);
and U23887 (N_23887,N_23402,N_23408);
nor U23888 (N_23888,N_23398,N_23384);
or U23889 (N_23889,N_23045,N_23469);
nand U23890 (N_23890,N_23080,N_23174);
and U23891 (N_23891,N_23319,N_23152);
nand U23892 (N_23892,N_23490,N_23326);
xnor U23893 (N_23893,N_23457,N_23040);
nand U23894 (N_23894,N_23433,N_23083);
nand U23895 (N_23895,N_23070,N_23214);
and U23896 (N_23896,N_23001,N_23033);
nor U23897 (N_23897,N_23137,N_23361);
or U23898 (N_23898,N_23201,N_23492);
nand U23899 (N_23899,N_23075,N_23082);
nor U23900 (N_23900,N_23067,N_23489);
or U23901 (N_23901,N_23137,N_23411);
nand U23902 (N_23902,N_23457,N_23193);
and U23903 (N_23903,N_23172,N_23418);
and U23904 (N_23904,N_23419,N_23495);
nor U23905 (N_23905,N_23003,N_23083);
nor U23906 (N_23906,N_23206,N_23153);
and U23907 (N_23907,N_23310,N_23004);
nor U23908 (N_23908,N_23060,N_23020);
nor U23909 (N_23909,N_23475,N_23141);
and U23910 (N_23910,N_23471,N_23490);
nand U23911 (N_23911,N_23041,N_23316);
nor U23912 (N_23912,N_23313,N_23166);
and U23913 (N_23913,N_23051,N_23115);
nand U23914 (N_23914,N_23151,N_23126);
and U23915 (N_23915,N_23007,N_23401);
nand U23916 (N_23916,N_23442,N_23372);
and U23917 (N_23917,N_23354,N_23206);
and U23918 (N_23918,N_23027,N_23013);
nand U23919 (N_23919,N_23412,N_23364);
nand U23920 (N_23920,N_23387,N_23144);
nand U23921 (N_23921,N_23013,N_23335);
or U23922 (N_23922,N_23399,N_23009);
and U23923 (N_23923,N_23366,N_23171);
nor U23924 (N_23924,N_23285,N_23022);
xor U23925 (N_23925,N_23384,N_23161);
nor U23926 (N_23926,N_23479,N_23227);
nor U23927 (N_23927,N_23097,N_23005);
or U23928 (N_23928,N_23422,N_23295);
or U23929 (N_23929,N_23265,N_23084);
nand U23930 (N_23930,N_23276,N_23045);
xnor U23931 (N_23931,N_23268,N_23023);
and U23932 (N_23932,N_23156,N_23272);
xnor U23933 (N_23933,N_23311,N_23301);
nor U23934 (N_23934,N_23042,N_23022);
and U23935 (N_23935,N_23284,N_23353);
nor U23936 (N_23936,N_23271,N_23142);
nand U23937 (N_23937,N_23278,N_23408);
or U23938 (N_23938,N_23486,N_23122);
nor U23939 (N_23939,N_23013,N_23024);
nor U23940 (N_23940,N_23309,N_23316);
nor U23941 (N_23941,N_23115,N_23422);
and U23942 (N_23942,N_23042,N_23492);
or U23943 (N_23943,N_23042,N_23226);
nor U23944 (N_23944,N_23089,N_23177);
or U23945 (N_23945,N_23192,N_23024);
and U23946 (N_23946,N_23263,N_23393);
nand U23947 (N_23947,N_23084,N_23326);
xnor U23948 (N_23948,N_23282,N_23004);
nand U23949 (N_23949,N_23402,N_23101);
nor U23950 (N_23950,N_23323,N_23305);
nand U23951 (N_23951,N_23319,N_23328);
or U23952 (N_23952,N_23172,N_23443);
nor U23953 (N_23953,N_23060,N_23276);
and U23954 (N_23954,N_23048,N_23081);
or U23955 (N_23955,N_23455,N_23225);
and U23956 (N_23956,N_23325,N_23312);
nor U23957 (N_23957,N_23043,N_23445);
and U23958 (N_23958,N_23103,N_23252);
and U23959 (N_23959,N_23412,N_23478);
or U23960 (N_23960,N_23488,N_23233);
nor U23961 (N_23961,N_23221,N_23444);
or U23962 (N_23962,N_23378,N_23220);
or U23963 (N_23963,N_23383,N_23019);
nand U23964 (N_23964,N_23361,N_23073);
xnor U23965 (N_23965,N_23141,N_23363);
nor U23966 (N_23966,N_23229,N_23017);
and U23967 (N_23967,N_23423,N_23122);
nand U23968 (N_23968,N_23024,N_23366);
and U23969 (N_23969,N_23422,N_23106);
xnor U23970 (N_23970,N_23369,N_23392);
and U23971 (N_23971,N_23317,N_23224);
nand U23972 (N_23972,N_23286,N_23048);
and U23973 (N_23973,N_23330,N_23419);
nand U23974 (N_23974,N_23137,N_23408);
and U23975 (N_23975,N_23229,N_23355);
nor U23976 (N_23976,N_23190,N_23278);
nor U23977 (N_23977,N_23030,N_23193);
nor U23978 (N_23978,N_23057,N_23077);
or U23979 (N_23979,N_23437,N_23184);
nor U23980 (N_23980,N_23358,N_23106);
or U23981 (N_23981,N_23091,N_23146);
nand U23982 (N_23982,N_23041,N_23163);
or U23983 (N_23983,N_23237,N_23344);
and U23984 (N_23984,N_23046,N_23009);
nor U23985 (N_23985,N_23258,N_23477);
nand U23986 (N_23986,N_23215,N_23031);
nand U23987 (N_23987,N_23440,N_23001);
and U23988 (N_23988,N_23358,N_23108);
and U23989 (N_23989,N_23107,N_23362);
nand U23990 (N_23990,N_23306,N_23315);
or U23991 (N_23991,N_23132,N_23286);
or U23992 (N_23992,N_23092,N_23368);
or U23993 (N_23993,N_23164,N_23387);
and U23994 (N_23994,N_23461,N_23123);
nor U23995 (N_23995,N_23210,N_23167);
nand U23996 (N_23996,N_23461,N_23478);
nor U23997 (N_23997,N_23119,N_23117);
and U23998 (N_23998,N_23407,N_23074);
nor U23999 (N_23999,N_23095,N_23261);
nand U24000 (N_24000,N_23640,N_23833);
xor U24001 (N_24001,N_23526,N_23918);
or U24002 (N_24002,N_23873,N_23782);
or U24003 (N_24003,N_23678,N_23767);
nor U24004 (N_24004,N_23956,N_23856);
nand U24005 (N_24005,N_23596,N_23671);
and U24006 (N_24006,N_23629,N_23616);
xor U24007 (N_24007,N_23706,N_23927);
nand U24008 (N_24008,N_23772,N_23999);
or U24009 (N_24009,N_23605,N_23836);
nor U24010 (N_24010,N_23679,N_23689);
and U24011 (N_24011,N_23727,N_23960);
or U24012 (N_24012,N_23949,N_23828);
nor U24013 (N_24013,N_23892,N_23571);
nand U24014 (N_24014,N_23751,N_23842);
or U24015 (N_24015,N_23698,N_23807);
or U24016 (N_24016,N_23834,N_23631);
nand U24017 (N_24017,N_23994,N_23861);
nand U24018 (N_24018,N_23951,N_23974);
and U24019 (N_24019,N_23703,N_23986);
and U24020 (N_24020,N_23800,N_23742);
and U24021 (N_24021,N_23862,N_23749);
nor U24022 (N_24022,N_23915,N_23535);
nor U24023 (N_24023,N_23839,N_23564);
xnor U24024 (N_24024,N_23922,N_23612);
nand U24025 (N_24025,N_23736,N_23619);
nand U24026 (N_24026,N_23843,N_23920);
or U24027 (N_24027,N_23525,N_23634);
nand U24028 (N_24028,N_23938,N_23684);
nand U24029 (N_24029,N_23558,N_23937);
or U24030 (N_24030,N_23648,N_23697);
nand U24031 (N_24031,N_23685,N_23926);
nor U24032 (N_24032,N_23987,N_23904);
nor U24033 (N_24033,N_23868,N_23804);
or U24034 (N_24034,N_23789,N_23917);
xnor U24035 (N_24035,N_23771,N_23660);
nor U24036 (N_24036,N_23667,N_23940);
xnor U24037 (N_24037,N_23528,N_23523);
nor U24038 (N_24038,N_23835,N_23916);
nand U24039 (N_24039,N_23729,N_23863);
nand U24040 (N_24040,N_23810,N_23880);
nand U24041 (N_24041,N_23580,N_23971);
nand U24042 (N_24042,N_23795,N_23981);
nand U24043 (N_24043,N_23841,N_23583);
nand U24044 (N_24044,N_23955,N_23931);
xnor U24045 (N_24045,N_23888,N_23819);
xnor U24046 (N_24046,N_23598,N_23794);
nor U24047 (N_24047,N_23978,N_23552);
or U24048 (N_24048,N_23850,N_23539);
or U24049 (N_24049,N_23876,N_23705);
and U24050 (N_24050,N_23533,N_23693);
nor U24051 (N_24051,N_23519,N_23641);
and U24052 (N_24052,N_23695,N_23658);
nor U24053 (N_24053,N_23781,N_23853);
and U24054 (N_24054,N_23731,N_23811);
or U24055 (N_24055,N_23952,N_23740);
or U24056 (N_24056,N_23633,N_23998);
nor U24057 (N_24057,N_23885,N_23769);
or U24058 (N_24058,N_23874,N_23816);
nor U24059 (N_24059,N_23770,N_23687);
and U24060 (N_24060,N_23893,N_23723);
nor U24061 (N_24061,N_23867,N_23899);
or U24062 (N_24062,N_23883,N_23902);
xor U24063 (N_24063,N_23611,N_23531);
nand U24064 (N_24064,N_23529,N_23959);
or U24065 (N_24065,N_23608,N_23775);
and U24066 (N_24066,N_23919,N_23557);
and U24067 (N_24067,N_23666,N_23713);
nand U24068 (N_24068,N_23607,N_23855);
or U24069 (N_24069,N_23824,N_23502);
nor U24070 (N_24070,N_23562,N_23910);
nand U24071 (N_24071,N_23550,N_23877);
xor U24072 (N_24072,N_23617,N_23501);
nor U24073 (N_24073,N_23936,N_23774);
or U24074 (N_24074,N_23979,N_23948);
or U24075 (N_24075,N_23933,N_23518);
and U24076 (N_24076,N_23548,N_23878);
and U24077 (N_24077,N_23964,N_23623);
xnor U24078 (N_24078,N_23761,N_23638);
and U24079 (N_24079,N_23668,N_23812);
or U24080 (N_24080,N_23965,N_23515);
and U24081 (N_24081,N_23887,N_23722);
or U24082 (N_24082,N_23696,N_23675);
xnor U24083 (N_24083,N_23721,N_23585);
nor U24084 (N_24084,N_23594,N_23815);
nand U24085 (N_24085,N_23872,N_23945);
or U24086 (N_24086,N_23909,N_23813);
xnor U24087 (N_24087,N_23718,N_23553);
and U24088 (N_24088,N_23724,N_23935);
and U24089 (N_24089,N_23676,N_23524);
or U24090 (N_24090,N_23540,N_23882);
nand U24091 (N_24091,N_23559,N_23942);
and U24092 (N_24092,N_23622,N_23983);
or U24093 (N_24093,N_23982,N_23912);
xor U24094 (N_24094,N_23680,N_23980);
nand U24095 (N_24095,N_23790,N_23976);
xor U24096 (N_24096,N_23568,N_23763);
and U24097 (N_24097,N_23954,N_23627);
nand U24098 (N_24098,N_23517,N_23711);
or U24099 (N_24099,N_23766,N_23669);
and U24100 (N_24100,N_23716,N_23646);
xnor U24101 (N_24101,N_23500,N_23972);
or U24102 (N_24102,N_23838,N_23637);
nand U24103 (N_24103,N_23614,N_23615);
nand U24104 (N_24104,N_23726,N_23510);
or U24105 (N_24105,N_23758,N_23532);
nor U24106 (N_24106,N_23601,N_23606);
xnor U24107 (N_24107,N_23664,N_23773);
xnor U24108 (N_24108,N_23822,N_23977);
nor U24109 (N_24109,N_23737,N_23691);
nor U24110 (N_24110,N_23900,N_23506);
xnor U24111 (N_24111,N_23780,N_23563);
nor U24112 (N_24112,N_23603,N_23542);
and U24113 (N_24113,N_23894,N_23673);
or U24114 (N_24114,N_23991,N_23860);
nor U24115 (N_24115,N_23953,N_23655);
or U24116 (N_24116,N_23886,N_23985);
xnor U24117 (N_24117,N_23599,N_23831);
nor U24118 (N_24118,N_23840,N_23674);
and U24119 (N_24119,N_23702,N_23895);
nand U24120 (N_24120,N_23651,N_23516);
nand U24121 (N_24121,N_23587,N_23777);
nand U24122 (N_24122,N_23744,N_23747);
or U24123 (N_24123,N_23597,N_23647);
nor U24124 (N_24124,N_23509,N_23717);
or U24125 (N_24125,N_23848,N_23875);
nor U24126 (N_24126,N_23572,N_23534);
nand U24127 (N_24127,N_23653,N_23707);
nand U24128 (N_24128,N_23681,N_23898);
and U24129 (N_24129,N_23569,N_23712);
or U24130 (N_24130,N_23743,N_23889);
nand U24131 (N_24131,N_23901,N_23549);
or U24132 (N_24132,N_23768,N_23586);
nor U24133 (N_24133,N_23869,N_23941);
and U24134 (N_24134,N_23521,N_23923);
or U24135 (N_24135,N_23595,N_23613);
or U24136 (N_24136,N_23752,N_23970);
nand U24137 (N_24137,N_23968,N_23925);
and U24138 (N_24138,N_23719,N_23665);
nor U24139 (N_24139,N_23830,N_23755);
xnor U24140 (N_24140,N_23939,N_23969);
and U24141 (N_24141,N_23859,N_23930);
or U24142 (N_24142,N_23576,N_23556);
xnor U24143 (N_24143,N_23609,N_23881);
and U24144 (N_24144,N_23546,N_23757);
nor U24145 (N_24145,N_23643,N_23928);
nand U24146 (N_24146,N_23753,N_23791);
nor U24147 (N_24147,N_23715,N_23710);
and U24148 (N_24148,N_23932,N_23659);
and U24149 (N_24149,N_23682,N_23701);
and U24150 (N_24150,N_23688,N_23801);
xor U24151 (N_24151,N_23505,N_23625);
or U24152 (N_24152,N_23750,N_23797);
nand U24153 (N_24153,N_23806,N_23662);
or U24154 (N_24154,N_23765,N_23575);
or U24155 (N_24155,N_23577,N_23778);
nand U24156 (N_24156,N_23589,N_23604);
nor U24157 (N_24157,N_23591,N_23890);
and U24158 (N_24158,N_23908,N_23884);
or U24159 (N_24159,N_23683,N_23512);
nor U24160 (N_24160,N_23686,N_23748);
nor U24161 (N_24161,N_23764,N_23990);
nand U24162 (N_24162,N_23639,N_23924);
nand U24163 (N_24163,N_23690,N_23630);
or U24164 (N_24164,N_23547,N_23738);
and U24165 (N_24165,N_23808,N_23988);
nand U24166 (N_24166,N_23896,N_23913);
nand U24167 (N_24167,N_23796,N_23992);
and U24168 (N_24168,N_23879,N_23624);
nor U24169 (N_24169,N_23997,N_23600);
nand U24170 (N_24170,N_23785,N_23714);
and U24171 (N_24171,N_23802,N_23582);
and U24172 (N_24172,N_23929,N_23820);
or U24173 (N_24173,N_23857,N_23579);
or U24174 (N_24174,N_23903,N_23642);
nor U24175 (N_24175,N_23565,N_23602);
nor U24176 (N_24176,N_23561,N_23864);
or U24177 (N_24177,N_23527,N_23530);
or U24178 (N_24178,N_23851,N_23825);
and U24179 (N_24179,N_23672,N_23537);
and U24180 (N_24180,N_23905,N_23656);
or U24181 (N_24181,N_23832,N_23829);
and U24182 (N_24182,N_23593,N_23805);
nor U24183 (N_24183,N_23844,N_23522);
or U24184 (N_24184,N_23975,N_23581);
and U24185 (N_24185,N_23628,N_23996);
nand U24186 (N_24186,N_23950,N_23733);
nor U24187 (N_24187,N_23745,N_23958);
xor U24188 (N_24188,N_23734,N_23995);
nand U24189 (N_24189,N_23567,N_23650);
or U24190 (N_24190,N_23788,N_23708);
and U24191 (N_24191,N_23943,N_23993);
xnor U24192 (N_24192,N_23618,N_23661);
nor U24193 (N_24193,N_23514,N_23845);
nor U24194 (N_24194,N_23984,N_23827);
and U24195 (N_24195,N_23837,N_23854);
and U24196 (N_24196,N_23520,N_23730);
xor U24197 (N_24197,N_23654,N_23538);
xor U24198 (N_24198,N_23866,N_23632);
nor U24199 (N_24199,N_23946,N_23746);
and U24200 (N_24200,N_23592,N_23652);
nor U24201 (N_24201,N_23677,N_23725);
nand U24202 (N_24202,N_23897,N_23784);
or U24203 (N_24203,N_23545,N_23760);
and U24204 (N_24204,N_23620,N_23793);
nor U24205 (N_24205,N_23741,N_23511);
xor U24206 (N_24206,N_23555,N_23657);
nand U24207 (N_24207,N_23636,N_23759);
nor U24208 (N_24208,N_23792,N_23944);
and U24209 (N_24209,N_23756,N_23649);
nor U24210 (N_24210,N_23911,N_23762);
xor U24211 (N_24211,N_23626,N_23720);
or U24212 (N_24212,N_23566,N_23709);
nand U24213 (N_24213,N_23541,N_23814);
nor U24214 (N_24214,N_23560,N_23551);
nor U24215 (N_24215,N_23739,N_23963);
or U24216 (N_24216,N_23826,N_23786);
or U24217 (N_24217,N_23906,N_23776);
nand U24218 (N_24218,N_23554,N_23973);
nand U24219 (N_24219,N_23821,N_23846);
nor U24220 (N_24220,N_23799,N_23513);
nor U24221 (N_24221,N_23847,N_23735);
nor U24222 (N_24222,N_23645,N_23663);
and U24223 (N_24223,N_23865,N_23728);
and U24224 (N_24224,N_23635,N_23732);
nor U24225 (N_24225,N_23670,N_23590);
and U24226 (N_24226,N_23803,N_23699);
nand U24227 (N_24227,N_23610,N_23694);
nor U24228 (N_24228,N_23503,N_23967);
or U24229 (N_24229,N_23621,N_23809);
nor U24230 (N_24230,N_23798,N_23544);
nand U24231 (N_24231,N_23921,N_23754);
or U24232 (N_24232,N_23961,N_23914);
nand U24233 (N_24233,N_23966,N_23858);
xnor U24234 (N_24234,N_23504,N_23787);
nor U24235 (N_24235,N_23578,N_23871);
nand U24236 (N_24236,N_23573,N_23818);
or U24237 (N_24237,N_23536,N_23644);
nand U24238 (N_24238,N_23907,N_23704);
xnor U24239 (N_24239,N_23957,N_23783);
and U24240 (N_24240,N_23700,N_23989);
nor U24241 (N_24241,N_23947,N_23870);
nand U24242 (N_24242,N_23588,N_23849);
nand U24243 (N_24243,N_23823,N_23692);
and U24244 (N_24244,N_23779,N_23934);
and U24245 (N_24245,N_23570,N_23962);
xnor U24246 (N_24246,N_23817,N_23574);
nor U24247 (N_24247,N_23852,N_23584);
and U24248 (N_24248,N_23891,N_23508);
and U24249 (N_24249,N_23507,N_23543);
xnor U24250 (N_24250,N_23847,N_23751);
nand U24251 (N_24251,N_23501,N_23746);
or U24252 (N_24252,N_23891,N_23636);
or U24253 (N_24253,N_23591,N_23741);
and U24254 (N_24254,N_23810,N_23573);
and U24255 (N_24255,N_23761,N_23985);
nand U24256 (N_24256,N_23582,N_23764);
or U24257 (N_24257,N_23633,N_23717);
nor U24258 (N_24258,N_23579,N_23622);
xor U24259 (N_24259,N_23853,N_23754);
nand U24260 (N_24260,N_23827,N_23753);
and U24261 (N_24261,N_23750,N_23882);
nand U24262 (N_24262,N_23772,N_23649);
and U24263 (N_24263,N_23590,N_23709);
and U24264 (N_24264,N_23917,N_23594);
and U24265 (N_24265,N_23662,N_23582);
nor U24266 (N_24266,N_23523,N_23505);
nand U24267 (N_24267,N_23677,N_23848);
nor U24268 (N_24268,N_23598,N_23947);
xor U24269 (N_24269,N_23946,N_23832);
and U24270 (N_24270,N_23914,N_23778);
and U24271 (N_24271,N_23619,N_23596);
or U24272 (N_24272,N_23537,N_23638);
and U24273 (N_24273,N_23631,N_23696);
or U24274 (N_24274,N_23735,N_23553);
or U24275 (N_24275,N_23828,N_23547);
nor U24276 (N_24276,N_23553,N_23665);
and U24277 (N_24277,N_23811,N_23522);
nor U24278 (N_24278,N_23677,N_23762);
and U24279 (N_24279,N_23826,N_23888);
nand U24280 (N_24280,N_23952,N_23717);
nor U24281 (N_24281,N_23990,N_23943);
or U24282 (N_24282,N_23964,N_23817);
nand U24283 (N_24283,N_23790,N_23675);
or U24284 (N_24284,N_23599,N_23823);
nor U24285 (N_24285,N_23574,N_23617);
or U24286 (N_24286,N_23629,N_23610);
or U24287 (N_24287,N_23641,N_23918);
nor U24288 (N_24288,N_23977,N_23859);
and U24289 (N_24289,N_23579,N_23873);
and U24290 (N_24290,N_23709,N_23520);
xnor U24291 (N_24291,N_23570,N_23501);
and U24292 (N_24292,N_23844,N_23533);
or U24293 (N_24293,N_23582,N_23605);
or U24294 (N_24294,N_23584,N_23747);
xor U24295 (N_24295,N_23707,N_23848);
nand U24296 (N_24296,N_23741,N_23602);
or U24297 (N_24297,N_23906,N_23677);
and U24298 (N_24298,N_23905,N_23504);
and U24299 (N_24299,N_23637,N_23842);
and U24300 (N_24300,N_23599,N_23929);
nor U24301 (N_24301,N_23749,N_23713);
and U24302 (N_24302,N_23945,N_23990);
and U24303 (N_24303,N_23850,N_23928);
and U24304 (N_24304,N_23600,N_23816);
or U24305 (N_24305,N_23652,N_23517);
and U24306 (N_24306,N_23699,N_23833);
nor U24307 (N_24307,N_23556,N_23790);
nor U24308 (N_24308,N_23688,N_23993);
or U24309 (N_24309,N_23917,N_23815);
nor U24310 (N_24310,N_23669,N_23557);
nor U24311 (N_24311,N_23547,N_23514);
or U24312 (N_24312,N_23924,N_23606);
and U24313 (N_24313,N_23551,N_23500);
or U24314 (N_24314,N_23850,N_23561);
or U24315 (N_24315,N_23800,N_23842);
xor U24316 (N_24316,N_23834,N_23676);
nor U24317 (N_24317,N_23866,N_23914);
and U24318 (N_24318,N_23536,N_23615);
and U24319 (N_24319,N_23969,N_23759);
nand U24320 (N_24320,N_23755,N_23858);
nor U24321 (N_24321,N_23665,N_23859);
nand U24322 (N_24322,N_23578,N_23577);
xnor U24323 (N_24323,N_23709,N_23753);
and U24324 (N_24324,N_23544,N_23846);
nand U24325 (N_24325,N_23646,N_23853);
nor U24326 (N_24326,N_23768,N_23991);
or U24327 (N_24327,N_23635,N_23579);
nand U24328 (N_24328,N_23538,N_23979);
and U24329 (N_24329,N_23607,N_23902);
and U24330 (N_24330,N_23603,N_23765);
or U24331 (N_24331,N_23656,N_23636);
nand U24332 (N_24332,N_23722,N_23909);
nor U24333 (N_24333,N_23839,N_23629);
or U24334 (N_24334,N_23989,N_23813);
and U24335 (N_24335,N_23575,N_23527);
nor U24336 (N_24336,N_23732,N_23550);
nor U24337 (N_24337,N_23585,N_23790);
and U24338 (N_24338,N_23522,N_23995);
nand U24339 (N_24339,N_23661,N_23956);
nor U24340 (N_24340,N_23766,N_23714);
and U24341 (N_24341,N_23523,N_23718);
nand U24342 (N_24342,N_23841,N_23752);
nand U24343 (N_24343,N_23907,N_23695);
and U24344 (N_24344,N_23792,N_23698);
and U24345 (N_24345,N_23714,N_23986);
nor U24346 (N_24346,N_23944,N_23671);
and U24347 (N_24347,N_23801,N_23696);
nand U24348 (N_24348,N_23674,N_23569);
nor U24349 (N_24349,N_23964,N_23987);
xnor U24350 (N_24350,N_23701,N_23886);
or U24351 (N_24351,N_23760,N_23985);
and U24352 (N_24352,N_23884,N_23504);
or U24353 (N_24353,N_23535,N_23657);
nand U24354 (N_24354,N_23692,N_23776);
nand U24355 (N_24355,N_23573,N_23932);
nor U24356 (N_24356,N_23522,N_23874);
nand U24357 (N_24357,N_23784,N_23959);
or U24358 (N_24358,N_23973,N_23810);
xor U24359 (N_24359,N_23508,N_23900);
or U24360 (N_24360,N_23952,N_23869);
or U24361 (N_24361,N_23680,N_23890);
or U24362 (N_24362,N_23543,N_23788);
and U24363 (N_24363,N_23727,N_23772);
nor U24364 (N_24364,N_23527,N_23914);
or U24365 (N_24365,N_23735,N_23793);
nor U24366 (N_24366,N_23945,N_23726);
or U24367 (N_24367,N_23841,N_23667);
nand U24368 (N_24368,N_23932,N_23778);
nor U24369 (N_24369,N_23902,N_23858);
nand U24370 (N_24370,N_23551,N_23537);
and U24371 (N_24371,N_23720,N_23675);
or U24372 (N_24372,N_23520,N_23560);
nand U24373 (N_24373,N_23980,N_23602);
nand U24374 (N_24374,N_23967,N_23686);
nor U24375 (N_24375,N_23956,N_23535);
nor U24376 (N_24376,N_23937,N_23707);
xnor U24377 (N_24377,N_23888,N_23929);
xor U24378 (N_24378,N_23740,N_23638);
nor U24379 (N_24379,N_23740,N_23670);
nor U24380 (N_24380,N_23548,N_23982);
nand U24381 (N_24381,N_23709,N_23930);
nand U24382 (N_24382,N_23952,N_23838);
xnor U24383 (N_24383,N_23749,N_23945);
nor U24384 (N_24384,N_23642,N_23820);
and U24385 (N_24385,N_23650,N_23600);
nand U24386 (N_24386,N_23691,N_23733);
nor U24387 (N_24387,N_23522,N_23595);
or U24388 (N_24388,N_23948,N_23907);
nand U24389 (N_24389,N_23980,N_23571);
nor U24390 (N_24390,N_23691,N_23647);
nor U24391 (N_24391,N_23950,N_23620);
nor U24392 (N_24392,N_23608,N_23671);
and U24393 (N_24393,N_23795,N_23688);
nand U24394 (N_24394,N_23914,N_23963);
xnor U24395 (N_24395,N_23758,N_23613);
nor U24396 (N_24396,N_23519,N_23601);
and U24397 (N_24397,N_23743,N_23765);
nor U24398 (N_24398,N_23691,N_23545);
nor U24399 (N_24399,N_23619,N_23920);
or U24400 (N_24400,N_23779,N_23589);
xnor U24401 (N_24401,N_23517,N_23835);
and U24402 (N_24402,N_23504,N_23972);
and U24403 (N_24403,N_23862,N_23681);
and U24404 (N_24404,N_23613,N_23641);
and U24405 (N_24405,N_23836,N_23882);
nor U24406 (N_24406,N_23989,N_23616);
xor U24407 (N_24407,N_23538,N_23915);
xnor U24408 (N_24408,N_23983,N_23930);
and U24409 (N_24409,N_23893,N_23967);
nor U24410 (N_24410,N_23763,N_23727);
xnor U24411 (N_24411,N_23644,N_23718);
and U24412 (N_24412,N_23602,N_23657);
nor U24413 (N_24413,N_23580,N_23726);
nor U24414 (N_24414,N_23768,N_23777);
or U24415 (N_24415,N_23610,N_23602);
nor U24416 (N_24416,N_23611,N_23605);
or U24417 (N_24417,N_23528,N_23519);
or U24418 (N_24418,N_23738,N_23894);
xor U24419 (N_24419,N_23621,N_23864);
nand U24420 (N_24420,N_23916,N_23537);
and U24421 (N_24421,N_23798,N_23818);
nand U24422 (N_24422,N_23952,N_23804);
nand U24423 (N_24423,N_23749,N_23711);
nor U24424 (N_24424,N_23670,N_23846);
or U24425 (N_24425,N_23587,N_23936);
and U24426 (N_24426,N_23577,N_23830);
xor U24427 (N_24427,N_23801,N_23693);
xor U24428 (N_24428,N_23516,N_23856);
and U24429 (N_24429,N_23623,N_23549);
nor U24430 (N_24430,N_23639,N_23955);
nand U24431 (N_24431,N_23705,N_23787);
nor U24432 (N_24432,N_23569,N_23959);
nand U24433 (N_24433,N_23934,N_23693);
and U24434 (N_24434,N_23502,N_23748);
or U24435 (N_24435,N_23584,N_23585);
nor U24436 (N_24436,N_23734,N_23659);
and U24437 (N_24437,N_23503,N_23957);
nor U24438 (N_24438,N_23743,N_23822);
nand U24439 (N_24439,N_23887,N_23894);
nand U24440 (N_24440,N_23507,N_23529);
or U24441 (N_24441,N_23614,N_23520);
nor U24442 (N_24442,N_23933,N_23965);
xnor U24443 (N_24443,N_23866,N_23509);
or U24444 (N_24444,N_23524,N_23521);
and U24445 (N_24445,N_23918,N_23645);
and U24446 (N_24446,N_23778,N_23943);
or U24447 (N_24447,N_23542,N_23697);
or U24448 (N_24448,N_23983,N_23995);
nand U24449 (N_24449,N_23685,N_23905);
nor U24450 (N_24450,N_23859,N_23905);
nand U24451 (N_24451,N_23947,N_23720);
or U24452 (N_24452,N_23695,N_23752);
or U24453 (N_24453,N_23745,N_23761);
and U24454 (N_24454,N_23718,N_23501);
or U24455 (N_24455,N_23672,N_23951);
xor U24456 (N_24456,N_23502,N_23580);
nor U24457 (N_24457,N_23907,N_23993);
nor U24458 (N_24458,N_23640,N_23826);
or U24459 (N_24459,N_23877,N_23918);
nor U24460 (N_24460,N_23605,N_23505);
and U24461 (N_24461,N_23603,N_23631);
nor U24462 (N_24462,N_23521,N_23904);
or U24463 (N_24463,N_23732,N_23657);
or U24464 (N_24464,N_23875,N_23557);
and U24465 (N_24465,N_23957,N_23769);
nor U24466 (N_24466,N_23562,N_23824);
nor U24467 (N_24467,N_23921,N_23672);
and U24468 (N_24468,N_23845,N_23874);
or U24469 (N_24469,N_23939,N_23506);
or U24470 (N_24470,N_23537,N_23955);
and U24471 (N_24471,N_23864,N_23650);
nor U24472 (N_24472,N_23927,N_23909);
or U24473 (N_24473,N_23957,N_23587);
xor U24474 (N_24474,N_23517,N_23618);
nor U24475 (N_24475,N_23784,N_23797);
or U24476 (N_24476,N_23891,N_23957);
xnor U24477 (N_24477,N_23969,N_23681);
nor U24478 (N_24478,N_23634,N_23556);
nor U24479 (N_24479,N_23520,N_23821);
or U24480 (N_24480,N_23959,N_23957);
and U24481 (N_24481,N_23652,N_23803);
or U24482 (N_24482,N_23663,N_23923);
nor U24483 (N_24483,N_23550,N_23928);
nand U24484 (N_24484,N_23986,N_23737);
or U24485 (N_24485,N_23787,N_23664);
xor U24486 (N_24486,N_23727,N_23581);
or U24487 (N_24487,N_23531,N_23668);
nor U24488 (N_24488,N_23776,N_23529);
nand U24489 (N_24489,N_23751,N_23819);
and U24490 (N_24490,N_23882,N_23613);
nand U24491 (N_24491,N_23934,N_23708);
nor U24492 (N_24492,N_23555,N_23878);
nand U24493 (N_24493,N_23653,N_23760);
nand U24494 (N_24494,N_23542,N_23579);
or U24495 (N_24495,N_23627,N_23824);
nor U24496 (N_24496,N_23844,N_23708);
nor U24497 (N_24497,N_23721,N_23993);
and U24498 (N_24498,N_23767,N_23552);
xnor U24499 (N_24499,N_23900,N_23753);
or U24500 (N_24500,N_24381,N_24080);
or U24501 (N_24501,N_24469,N_24045);
nor U24502 (N_24502,N_24444,N_24081);
nand U24503 (N_24503,N_24284,N_24335);
nor U24504 (N_24504,N_24061,N_24231);
and U24505 (N_24505,N_24328,N_24446);
or U24506 (N_24506,N_24115,N_24135);
nand U24507 (N_24507,N_24130,N_24226);
nor U24508 (N_24508,N_24321,N_24464);
nand U24509 (N_24509,N_24288,N_24405);
nor U24510 (N_24510,N_24058,N_24119);
nor U24511 (N_24511,N_24285,N_24268);
xor U24512 (N_24512,N_24267,N_24259);
nand U24513 (N_24513,N_24489,N_24018);
nor U24514 (N_24514,N_24315,N_24352);
and U24515 (N_24515,N_24056,N_24105);
nand U24516 (N_24516,N_24294,N_24498);
or U24517 (N_24517,N_24037,N_24090);
nor U24518 (N_24518,N_24176,N_24133);
nor U24519 (N_24519,N_24095,N_24302);
or U24520 (N_24520,N_24363,N_24232);
or U24521 (N_24521,N_24024,N_24006);
or U24522 (N_24522,N_24383,N_24374);
and U24523 (N_24523,N_24162,N_24209);
nand U24524 (N_24524,N_24438,N_24454);
and U24525 (N_24525,N_24425,N_24424);
xnor U24526 (N_24526,N_24083,N_24218);
and U24527 (N_24527,N_24034,N_24307);
and U24528 (N_24528,N_24141,N_24341);
and U24529 (N_24529,N_24370,N_24409);
and U24530 (N_24530,N_24017,N_24166);
or U24531 (N_24531,N_24369,N_24487);
nand U24532 (N_24532,N_24255,N_24089);
or U24533 (N_24533,N_24210,N_24099);
nand U24534 (N_24534,N_24091,N_24170);
nor U24535 (N_24535,N_24174,N_24493);
nor U24536 (N_24536,N_24477,N_24295);
nor U24537 (N_24537,N_24350,N_24411);
nor U24538 (N_24538,N_24296,N_24180);
nand U24539 (N_24539,N_24479,N_24450);
and U24540 (N_24540,N_24338,N_24276);
and U24541 (N_24541,N_24159,N_24376);
nor U24542 (N_24542,N_24153,N_24320);
and U24543 (N_24543,N_24154,N_24336);
nand U24544 (N_24544,N_24447,N_24217);
nor U24545 (N_24545,N_24216,N_24113);
or U24546 (N_24546,N_24474,N_24007);
nand U24547 (N_24547,N_24012,N_24325);
nor U24548 (N_24548,N_24029,N_24401);
or U24549 (N_24549,N_24165,N_24392);
and U24550 (N_24550,N_24497,N_24048);
or U24551 (N_24551,N_24275,N_24264);
nor U24552 (N_24552,N_24142,N_24459);
nor U24553 (N_24553,N_24312,N_24291);
nor U24554 (N_24554,N_24238,N_24262);
and U24555 (N_24555,N_24421,N_24011);
or U24556 (N_24556,N_24175,N_24345);
nor U24557 (N_24557,N_24414,N_24234);
nand U24558 (N_24558,N_24127,N_24195);
nor U24559 (N_24559,N_24125,N_24388);
xnor U24560 (N_24560,N_24049,N_24208);
nor U24561 (N_24561,N_24440,N_24377);
and U24562 (N_24562,N_24179,N_24040);
or U24563 (N_24563,N_24239,N_24423);
nand U24564 (N_24564,N_24389,N_24213);
or U24565 (N_24565,N_24198,N_24279);
nor U24566 (N_24566,N_24185,N_24396);
nor U24567 (N_24567,N_24160,N_24094);
nor U24568 (N_24568,N_24346,N_24106);
xor U24569 (N_24569,N_24437,N_24043);
or U24570 (N_24570,N_24257,N_24261);
nor U24571 (N_24571,N_24164,N_24281);
nand U24572 (N_24572,N_24413,N_24362);
and U24573 (N_24573,N_24270,N_24023);
nand U24574 (N_24574,N_24458,N_24373);
nor U24575 (N_24575,N_24220,N_24455);
nor U24576 (N_24576,N_24399,N_24204);
and U24577 (N_24577,N_24055,N_24301);
nand U24578 (N_24578,N_24044,N_24087);
xor U24579 (N_24579,N_24138,N_24177);
or U24580 (N_24580,N_24072,N_24104);
nor U24581 (N_24581,N_24112,N_24330);
nand U24582 (N_24582,N_24453,N_24151);
or U24583 (N_24583,N_24380,N_24282);
nand U24584 (N_24584,N_24486,N_24491);
or U24585 (N_24585,N_24070,N_24355);
or U24586 (N_24586,N_24173,N_24327);
or U24587 (N_24587,N_24286,N_24078);
and U24588 (N_24588,N_24416,N_24054);
or U24589 (N_24589,N_24111,N_24365);
xor U24590 (N_24590,N_24121,N_24131);
nor U24591 (N_24591,N_24030,N_24499);
and U24592 (N_24592,N_24168,N_24186);
or U24593 (N_24593,N_24269,N_24475);
or U24594 (N_24594,N_24129,N_24434);
xnor U24595 (N_24595,N_24071,N_24062);
or U24596 (N_24596,N_24225,N_24371);
nand U24597 (N_24597,N_24260,N_24236);
or U24598 (N_24598,N_24467,N_24169);
or U24599 (N_24599,N_24445,N_24337);
nor U24600 (N_24600,N_24379,N_24488);
nor U24601 (N_24601,N_24188,N_24344);
nor U24602 (N_24602,N_24123,N_24274);
xnor U24603 (N_24603,N_24435,N_24323);
or U24604 (N_24604,N_24100,N_24098);
nor U24605 (N_24605,N_24155,N_24067);
and U24606 (N_24606,N_24429,N_24351);
xor U24607 (N_24607,N_24481,N_24184);
nor U24608 (N_24608,N_24490,N_24485);
or U24609 (N_24609,N_24200,N_24266);
and U24610 (N_24610,N_24248,N_24258);
and U24611 (N_24611,N_24400,N_24036);
xor U24612 (N_24612,N_24244,N_24026);
nand U24613 (N_24613,N_24163,N_24457);
or U24614 (N_24614,N_24065,N_24375);
xnor U24615 (N_24615,N_24367,N_24110);
or U24616 (N_24616,N_24410,N_24317);
nand U24617 (N_24617,N_24229,N_24240);
nand U24618 (N_24618,N_24033,N_24386);
nor U24619 (N_24619,N_24496,N_24342);
nor U24620 (N_24620,N_24347,N_24366);
nor U24621 (N_24621,N_24003,N_24283);
nor U24622 (N_24622,N_24382,N_24339);
or U24623 (N_24623,N_24158,N_24107);
nor U24624 (N_24624,N_24309,N_24197);
and U24625 (N_24625,N_24057,N_24390);
and U24626 (N_24626,N_24357,N_24332);
nand U24627 (N_24627,N_24117,N_24356);
or U24628 (N_24628,N_24292,N_24418);
nand U24629 (N_24629,N_24066,N_24265);
and U24630 (N_24630,N_24349,N_24230);
and U24631 (N_24631,N_24436,N_24465);
or U24632 (N_24632,N_24172,N_24093);
or U24633 (N_24633,N_24466,N_24406);
and U24634 (N_24634,N_24076,N_24428);
xnor U24635 (N_24635,N_24441,N_24224);
nand U24636 (N_24636,N_24451,N_24157);
or U24637 (N_24637,N_24181,N_24103);
and U24638 (N_24638,N_24422,N_24308);
nor U24639 (N_24639,N_24387,N_24042);
nor U24640 (N_24640,N_24092,N_24136);
xor U24641 (N_24641,N_24074,N_24476);
and U24642 (N_24642,N_24047,N_24187);
or U24643 (N_24643,N_24319,N_24201);
or U24644 (N_24644,N_24427,N_24391);
nor U24645 (N_24645,N_24063,N_24073);
xor U24646 (N_24646,N_24102,N_24364);
nand U24647 (N_24647,N_24235,N_24009);
and U24648 (N_24648,N_24306,N_24182);
or U24649 (N_24649,N_24452,N_24008);
or U24650 (N_24650,N_24334,N_24463);
and U24651 (N_24651,N_24252,N_24359);
xor U24652 (N_24652,N_24132,N_24233);
or U24653 (N_24653,N_24120,N_24395);
nor U24654 (N_24654,N_24482,N_24417);
xnor U24655 (N_24655,N_24430,N_24211);
nor U24656 (N_24656,N_24118,N_24075);
and U24657 (N_24657,N_24096,N_24191);
nor U24658 (N_24658,N_24189,N_24031);
nand U24659 (N_24659,N_24140,N_24397);
and U24660 (N_24660,N_24254,N_24223);
and U24661 (N_24661,N_24245,N_24039);
nand U24662 (N_24662,N_24004,N_24331);
nor U24663 (N_24663,N_24271,N_24456);
nor U24664 (N_24664,N_24122,N_24041);
nor U24665 (N_24665,N_24368,N_24426);
xnor U24666 (N_24666,N_24412,N_24206);
nand U24667 (N_24667,N_24484,N_24263);
nand U24668 (N_24668,N_24084,N_24237);
nor U24669 (N_24669,N_24082,N_24214);
and U24670 (N_24670,N_24014,N_24303);
nor U24671 (N_24671,N_24431,N_24404);
or U24672 (N_24672,N_24468,N_24203);
nand U24673 (N_24673,N_24473,N_24300);
or U24674 (N_24674,N_24207,N_24495);
nand U24675 (N_24675,N_24097,N_24432);
or U24676 (N_24676,N_24290,N_24318);
nor U24677 (N_24677,N_24035,N_24150);
and U24678 (N_24678,N_24013,N_24215);
and U24679 (N_24679,N_24384,N_24183);
nor U24680 (N_24680,N_24228,N_24433);
nand U24681 (N_24681,N_24360,N_24101);
nor U24682 (N_24682,N_24147,N_24287);
nor U24683 (N_24683,N_24146,N_24193);
nor U24684 (N_24684,N_24448,N_24253);
nand U24685 (N_24685,N_24116,N_24134);
nand U24686 (N_24686,N_24394,N_24354);
or U24687 (N_24687,N_24333,N_24402);
and U24688 (N_24688,N_24152,N_24086);
or U24689 (N_24689,N_24016,N_24143);
nor U24690 (N_24690,N_24298,N_24273);
nor U24691 (N_24691,N_24088,N_24322);
nor U24692 (N_24692,N_24114,N_24190);
and U24693 (N_24693,N_24472,N_24311);
or U24694 (N_24694,N_24398,N_24324);
xor U24695 (N_24695,N_24247,N_24439);
nor U24696 (N_24696,N_24053,N_24407);
nor U24697 (N_24697,N_24002,N_24109);
nor U24698 (N_24698,N_24478,N_24242);
and U24699 (N_24699,N_24156,N_24348);
nand U24700 (N_24700,N_24205,N_24408);
nor U24701 (N_24701,N_24251,N_24196);
xnor U24702 (N_24702,N_24415,N_24494);
nor U24703 (N_24703,N_24167,N_24278);
nor U24704 (N_24704,N_24137,N_24372);
nor U24705 (N_24705,N_24246,N_24001);
nand U24706 (N_24706,N_24419,N_24028);
nor U24707 (N_24707,N_24480,N_24199);
nand U24708 (N_24708,N_24343,N_24243);
nand U24709 (N_24709,N_24241,N_24005);
or U24710 (N_24710,N_24161,N_24293);
or U24711 (N_24711,N_24124,N_24492);
nor U24712 (N_24712,N_24052,N_24015);
xnor U24713 (N_24713,N_24222,N_24149);
nor U24714 (N_24714,N_24250,N_24171);
and U24715 (N_24715,N_24144,N_24219);
or U24716 (N_24716,N_24000,N_24314);
nand U24717 (N_24717,N_24126,N_24462);
nand U24718 (N_24718,N_24064,N_24289);
nand U24719 (N_24719,N_24378,N_24272);
xor U24720 (N_24720,N_24050,N_24192);
nand U24721 (N_24721,N_24256,N_24461);
or U24722 (N_24722,N_24358,N_24305);
nor U24723 (N_24723,N_24460,N_24060);
or U24724 (N_24724,N_24032,N_24340);
or U24725 (N_24725,N_24145,N_24128);
nand U24726 (N_24726,N_24326,N_24077);
and U24727 (N_24727,N_24025,N_24046);
nand U24728 (N_24728,N_24449,N_24310);
nor U24729 (N_24729,N_24483,N_24443);
xnor U24730 (N_24730,N_24393,N_24022);
nand U24731 (N_24731,N_24202,N_24212);
or U24732 (N_24732,N_24470,N_24353);
nand U24733 (N_24733,N_24148,N_24403);
nand U24734 (N_24734,N_24316,N_24297);
nor U24735 (N_24735,N_24304,N_24299);
nor U24736 (N_24736,N_24019,N_24420);
xnor U24737 (N_24737,N_24021,N_24068);
and U24738 (N_24738,N_24059,N_24079);
or U24739 (N_24739,N_24280,N_24010);
and U24740 (N_24740,N_24249,N_24221);
nand U24741 (N_24741,N_24442,N_24085);
or U24742 (N_24742,N_24051,N_24227);
nor U24743 (N_24743,N_24178,N_24329);
nor U24744 (N_24744,N_24027,N_24194);
and U24745 (N_24745,N_24139,N_24385);
xor U24746 (N_24746,N_24108,N_24038);
nand U24747 (N_24747,N_24277,N_24020);
nor U24748 (N_24748,N_24069,N_24361);
nand U24749 (N_24749,N_24313,N_24471);
nor U24750 (N_24750,N_24045,N_24451);
nand U24751 (N_24751,N_24070,N_24204);
and U24752 (N_24752,N_24482,N_24285);
nor U24753 (N_24753,N_24416,N_24324);
nor U24754 (N_24754,N_24026,N_24381);
nor U24755 (N_24755,N_24344,N_24064);
nor U24756 (N_24756,N_24398,N_24029);
and U24757 (N_24757,N_24326,N_24274);
xor U24758 (N_24758,N_24228,N_24247);
nor U24759 (N_24759,N_24417,N_24469);
and U24760 (N_24760,N_24458,N_24221);
nand U24761 (N_24761,N_24106,N_24403);
or U24762 (N_24762,N_24399,N_24035);
nor U24763 (N_24763,N_24439,N_24399);
and U24764 (N_24764,N_24040,N_24288);
nor U24765 (N_24765,N_24105,N_24170);
nor U24766 (N_24766,N_24335,N_24184);
or U24767 (N_24767,N_24216,N_24318);
nand U24768 (N_24768,N_24378,N_24096);
or U24769 (N_24769,N_24074,N_24168);
xnor U24770 (N_24770,N_24083,N_24023);
xor U24771 (N_24771,N_24363,N_24475);
nor U24772 (N_24772,N_24386,N_24209);
nand U24773 (N_24773,N_24126,N_24015);
or U24774 (N_24774,N_24475,N_24045);
nand U24775 (N_24775,N_24340,N_24073);
xor U24776 (N_24776,N_24344,N_24391);
nand U24777 (N_24777,N_24108,N_24426);
nor U24778 (N_24778,N_24448,N_24321);
and U24779 (N_24779,N_24362,N_24404);
nand U24780 (N_24780,N_24483,N_24376);
xor U24781 (N_24781,N_24048,N_24207);
or U24782 (N_24782,N_24142,N_24225);
nand U24783 (N_24783,N_24247,N_24152);
nor U24784 (N_24784,N_24397,N_24007);
nor U24785 (N_24785,N_24244,N_24061);
nand U24786 (N_24786,N_24250,N_24325);
nand U24787 (N_24787,N_24462,N_24465);
and U24788 (N_24788,N_24357,N_24245);
nor U24789 (N_24789,N_24050,N_24055);
nor U24790 (N_24790,N_24140,N_24077);
and U24791 (N_24791,N_24194,N_24477);
xnor U24792 (N_24792,N_24262,N_24404);
or U24793 (N_24793,N_24312,N_24118);
and U24794 (N_24794,N_24428,N_24151);
or U24795 (N_24795,N_24093,N_24480);
nand U24796 (N_24796,N_24453,N_24271);
nor U24797 (N_24797,N_24250,N_24085);
nand U24798 (N_24798,N_24351,N_24223);
and U24799 (N_24799,N_24126,N_24410);
or U24800 (N_24800,N_24385,N_24392);
nor U24801 (N_24801,N_24180,N_24239);
and U24802 (N_24802,N_24395,N_24102);
xor U24803 (N_24803,N_24387,N_24279);
nor U24804 (N_24804,N_24087,N_24386);
and U24805 (N_24805,N_24397,N_24180);
xnor U24806 (N_24806,N_24228,N_24067);
nand U24807 (N_24807,N_24195,N_24048);
nor U24808 (N_24808,N_24472,N_24353);
nand U24809 (N_24809,N_24079,N_24364);
or U24810 (N_24810,N_24356,N_24002);
and U24811 (N_24811,N_24085,N_24434);
nor U24812 (N_24812,N_24171,N_24261);
or U24813 (N_24813,N_24394,N_24237);
and U24814 (N_24814,N_24096,N_24006);
xnor U24815 (N_24815,N_24188,N_24429);
nand U24816 (N_24816,N_24007,N_24322);
and U24817 (N_24817,N_24454,N_24343);
and U24818 (N_24818,N_24410,N_24435);
and U24819 (N_24819,N_24361,N_24124);
and U24820 (N_24820,N_24085,N_24121);
or U24821 (N_24821,N_24363,N_24308);
nor U24822 (N_24822,N_24211,N_24478);
nor U24823 (N_24823,N_24080,N_24372);
xnor U24824 (N_24824,N_24047,N_24226);
and U24825 (N_24825,N_24430,N_24003);
nand U24826 (N_24826,N_24065,N_24453);
nor U24827 (N_24827,N_24032,N_24182);
or U24828 (N_24828,N_24141,N_24379);
nor U24829 (N_24829,N_24465,N_24127);
or U24830 (N_24830,N_24189,N_24455);
nor U24831 (N_24831,N_24361,N_24173);
or U24832 (N_24832,N_24467,N_24063);
nand U24833 (N_24833,N_24014,N_24479);
or U24834 (N_24834,N_24356,N_24422);
xnor U24835 (N_24835,N_24280,N_24192);
xnor U24836 (N_24836,N_24034,N_24485);
nor U24837 (N_24837,N_24403,N_24185);
nor U24838 (N_24838,N_24046,N_24317);
and U24839 (N_24839,N_24261,N_24350);
or U24840 (N_24840,N_24179,N_24083);
nand U24841 (N_24841,N_24089,N_24029);
nor U24842 (N_24842,N_24413,N_24005);
nor U24843 (N_24843,N_24430,N_24239);
nand U24844 (N_24844,N_24263,N_24363);
and U24845 (N_24845,N_24209,N_24034);
or U24846 (N_24846,N_24455,N_24004);
or U24847 (N_24847,N_24272,N_24386);
nand U24848 (N_24848,N_24457,N_24312);
and U24849 (N_24849,N_24070,N_24146);
and U24850 (N_24850,N_24435,N_24347);
nor U24851 (N_24851,N_24038,N_24411);
xor U24852 (N_24852,N_24378,N_24334);
or U24853 (N_24853,N_24008,N_24039);
or U24854 (N_24854,N_24290,N_24486);
and U24855 (N_24855,N_24269,N_24289);
and U24856 (N_24856,N_24011,N_24457);
and U24857 (N_24857,N_24454,N_24370);
or U24858 (N_24858,N_24459,N_24288);
xor U24859 (N_24859,N_24287,N_24184);
xor U24860 (N_24860,N_24251,N_24076);
nor U24861 (N_24861,N_24422,N_24083);
and U24862 (N_24862,N_24397,N_24107);
xor U24863 (N_24863,N_24384,N_24086);
nor U24864 (N_24864,N_24133,N_24424);
and U24865 (N_24865,N_24236,N_24112);
or U24866 (N_24866,N_24362,N_24364);
and U24867 (N_24867,N_24161,N_24199);
or U24868 (N_24868,N_24170,N_24041);
nand U24869 (N_24869,N_24362,N_24456);
nor U24870 (N_24870,N_24139,N_24475);
nor U24871 (N_24871,N_24177,N_24017);
nor U24872 (N_24872,N_24230,N_24397);
nand U24873 (N_24873,N_24014,N_24224);
or U24874 (N_24874,N_24481,N_24400);
or U24875 (N_24875,N_24355,N_24015);
nand U24876 (N_24876,N_24219,N_24099);
xnor U24877 (N_24877,N_24435,N_24188);
nand U24878 (N_24878,N_24319,N_24408);
xnor U24879 (N_24879,N_24197,N_24234);
xor U24880 (N_24880,N_24331,N_24246);
nor U24881 (N_24881,N_24016,N_24267);
or U24882 (N_24882,N_24243,N_24072);
nand U24883 (N_24883,N_24431,N_24213);
nor U24884 (N_24884,N_24026,N_24208);
and U24885 (N_24885,N_24177,N_24057);
xor U24886 (N_24886,N_24369,N_24429);
or U24887 (N_24887,N_24437,N_24158);
nor U24888 (N_24888,N_24475,N_24020);
or U24889 (N_24889,N_24143,N_24418);
and U24890 (N_24890,N_24315,N_24031);
or U24891 (N_24891,N_24468,N_24362);
or U24892 (N_24892,N_24340,N_24240);
nand U24893 (N_24893,N_24371,N_24272);
nor U24894 (N_24894,N_24244,N_24210);
or U24895 (N_24895,N_24156,N_24055);
and U24896 (N_24896,N_24405,N_24471);
or U24897 (N_24897,N_24240,N_24385);
or U24898 (N_24898,N_24491,N_24337);
nand U24899 (N_24899,N_24230,N_24495);
nor U24900 (N_24900,N_24066,N_24409);
or U24901 (N_24901,N_24039,N_24268);
nor U24902 (N_24902,N_24389,N_24378);
nor U24903 (N_24903,N_24370,N_24290);
and U24904 (N_24904,N_24288,N_24094);
and U24905 (N_24905,N_24211,N_24246);
xnor U24906 (N_24906,N_24342,N_24114);
and U24907 (N_24907,N_24002,N_24499);
nand U24908 (N_24908,N_24213,N_24198);
nand U24909 (N_24909,N_24365,N_24226);
nand U24910 (N_24910,N_24191,N_24407);
nor U24911 (N_24911,N_24123,N_24340);
nor U24912 (N_24912,N_24306,N_24191);
or U24913 (N_24913,N_24098,N_24423);
and U24914 (N_24914,N_24011,N_24101);
nand U24915 (N_24915,N_24258,N_24151);
and U24916 (N_24916,N_24182,N_24435);
nor U24917 (N_24917,N_24353,N_24373);
or U24918 (N_24918,N_24325,N_24025);
or U24919 (N_24919,N_24457,N_24099);
or U24920 (N_24920,N_24364,N_24031);
xnor U24921 (N_24921,N_24045,N_24035);
nand U24922 (N_24922,N_24158,N_24228);
and U24923 (N_24923,N_24324,N_24291);
nand U24924 (N_24924,N_24450,N_24387);
nor U24925 (N_24925,N_24224,N_24385);
or U24926 (N_24926,N_24087,N_24312);
and U24927 (N_24927,N_24396,N_24086);
nand U24928 (N_24928,N_24423,N_24034);
or U24929 (N_24929,N_24442,N_24357);
nor U24930 (N_24930,N_24017,N_24082);
or U24931 (N_24931,N_24135,N_24068);
and U24932 (N_24932,N_24294,N_24367);
nand U24933 (N_24933,N_24352,N_24367);
nor U24934 (N_24934,N_24218,N_24182);
and U24935 (N_24935,N_24230,N_24011);
xnor U24936 (N_24936,N_24358,N_24141);
xnor U24937 (N_24937,N_24431,N_24333);
nor U24938 (N_24938,N_24307,N_24393);
nor U24939 (N_24939,N_24402,N_24091);
and U24940 (N_24940,N_24191,N_24421);
nand U24941 (N_24941,N_24309,N_24333);
or U24942 (N_24942,N_24211,N_24429);
nor U24943 (N_24943,N_24198,N_24284);
and U24944 (N_24944,N_24031,N_24218);
xnor U24945 (N_24945,N_24150,N_24189);
and U24946 (N_24946,N_24017,N_24072);
xor U24947 (N_24947,N_24115,N_24383);
nand U24948 (N_24948,N_24032,N_24362);
and U24949 (N_24949,N_24210,N_24067);
nand U24950 (N_24950,N_24419,N_24436);
nand U24951 (N_24951,N_24177,N_24124);
nor U24952 (N_24952,N_24167,N_24105);
or U24953 (N_24953,N_24117,N_24136);
nand U24954 (N_24954,N_24498,N_24300);
or U24955 (N_24955,N_24496,N_24331);
and U24956 (N_24956,N_24305,N_24024);
nor U24957 (N_24957,N_24350,N_24386);
or U24958 (N_24958,N_24458,N_24032);
and U24959 (N_24959,N_24479,N_24017);
and U24960 (N_24960,N_24457,N_24356);
nand U24961 (N_24961,N_24034,N_24208);
nor U24962 (N_24962,N_24407,N_24319);
nand U24963 (N_24963,N_24256,N_24339);
and U24964 (N_24964,N_24087,N_24029);
nor U24965 (N_24965,N_24397,N_24458);
nand U24966 (N_24966,N_24039,N_24311);
or U24967 (N_24967,N_24190,N_24074);
nor U24968 (N_24968,N_24477,N_24248);
or U24969 (N_24969,N_24415,N_24272);
or U24970 (N_24970,N_24477,N_24311);
nor U24971 (N_24971,N_24476,N_24171);
or U24972 (N_24972,N_24359,N_24488);
nand U24973 (N_24973,N_24408,N_24148);
nor U24974 (N_24974,N_24368,N_24227);
and U24975 (N_24975,N_24287,N_24078);
nor U24976 (N_24976,N_24391,N_24279);
and U24977 (N_24977,N_24103,N_24344);
and U24978 (N_24978,N_24263,N_24108);
nand U24979 (N_24979,N_24101,N_24032);
nor U24980 (N_24980,N_24431,N_24106);
or U24981 (N_24981,N_24285,N_24190);
and U24982 (N_24982,N_24023,N_24222);
or U24983 (N_24983,N_24011,N_24156);
and U24984 (N_24984,N_24241,N_24425);
nand U24985 (N_24985,N_24386,N_24133);
nand U24986 (N_24986,N_24365,N_24363);
nand U24987 (N_24987,N_24237,N_24330);
or U24988 (N_24988,N_24079,N_24264);
or U24989 (N_24989,N_24497,N_24137);
or U24990 (N_24990,N_24394,N_24154);
nand U24991 (N_24991,N_24083,N_24333);
nor U24992 (N_24992,N_24044,N_24456);
nand U24993 (N_24993,N_24234,N_24431);
nor U24994 (N_24994,N_24337,N_24031);
nor U24995 (N_24995,N_24032,N_24365);
and U24996 (N_24996,N_24487,N_24298);
xor U24997 (N_24997,N_24087,N_24272);
or U24998 (N_24998,N_24035,N_24023);
nor U24999 (N_24999,N_24144,N_24075);
nor UO_0 (O_0,N_24834,N_24997);
and UO_1 (O_1,N_24500,N_24794);
or UO_2 (O_2,N_24601,N_24906);
nand UO_3 (O_3,N_24687,N_24513);
nand UO_4 (O_4,N_24713,N_24824);
nand UO_5 (O_5,N_24909,N_24791);
xor UO_6 (O_6,N_24890,N_24869);
or UO_7 (O_7,N_24952,N_24857);
nor UO_8 (O_8,N_24755,N_24522);
nand UO_9 (O_9,N_24995,N_24837);
and UO_10 (O_10,N_24682,N_24940);
and UO_11 (O_11,N_24569,N_24514);
or UO_12 (O_12,N_24836,N_24889);
nand UO_13 (O_13,N_24547,N_24655);
or UO_14 (O_14,N_24550,N_24955);
or UO_15 (O_15,N_24705,N_24849);
or UO_16 (O_16,N_24663,N_24701);
nand UO_17 (O_17,N_24598,N_24638);
nor UO_18 (O_18,N_24776,N_24935);
or UO_19 (O_19,N_24628,N_24826);
or UO_20 (O_20,N_24786,N_24504);
or UO_21 (O_21,N_24694,N_24662);
xor UO_22 (O_22,N_24936,N_24803);
and UO_23 (O_23,N_24648,N_24905);
xor UO_24 (O_24,N_24654,N_24901);
nor UO_25 (O_25,N_24767,N_24549);
nor UO_26 (O_26,N_24829,N_24691);
and UO_27 (O_27,N_24542,N_24925);
and UO_28 (O_28,N_24949,N_24641);
nand UO_29 (O_29,N_24808,N_24611);
and UO_30 (O_30,N_24528,N_24702);
nand UO_31 (O_31,N_24804,N_24552);
or UO_32 (O_32,N_24576,N_24593);
nand UO_33 (O_33,N_24548,N_24765);
nand UO_34 (O_34,N_24976,N_24966);
nor UO_35 (O_35,N_24977,N_24895);
and UO_36 (O_36,N_24914,N_24572);
and UO_37 (O_37,N_24879,N_24560);
and UO_38 (O_38,N_24639,N_24902);
and UO_39 (O_39,N_24630,N_24562);
and UO_40 (O_40,N_24679,N_24689);
nor UO_41 (O_41,N_24831,N_24554);
xnor UO_42 (O_42,N_24850,N_24810);
and UO_43 (O_43,N_24659,N_24861);
nand UO_44 (O_44,N_24880,N_24922);
and UO_45 (O_45,N_24932,N_24590);
or UO_46 (O_46,N_24874,N_24555);
nand UO_47 (O_47,N_24722,N_24627);
or UO_48 (O_48,N_24969,N_24657);
nand UO_49 (O_49,N_24870,N_24941);
or UO_50 (O_50,N_24759,N_24757);
and UO_51 (O_51,N_24983,N_24600);
nand UO_52 (O_52,N_24573,N_24944);
nor UO_53 (O_53,N_24723,N_24884);
nor UO_54 (O_54,N_24825,N_24948);
or UO_55 (O_55,N_24915,N_24678);
and UO_56 (O_56,N_24896,N_24758);
nor UO_57 (O_57,N_24762,N_24798);
or UO_58 (O_58,N_24970,N_24529);
and UO_59 (O_59,N_24649,N_24636);
or UO_60 (O_60,N_24832,N_24957);
or UO_61 (O_61,N_24737,N_24992);
or UO_62 (O_62,N_24809,N_24581);
nor UO_63 (O_63,N_24621,N_24530);
nand UO_64 (O_64,N_24629,N_24833);
and UO_65 (O_65,N_24586,N_24877);
nand UO_66 (O_66,N_24766,N_24646);
or UO_67 (O_67,N_24887,N_24864);
nor UO_68 (O_68,N_24811,N_24644);
nand UO_69 (O_69,N_24930,N_24579);
nand UO_70 (O_70,N_24945,N_24728);
and UO_71 (O_71,N_24635,N_24990);
or UO_72 (O_72,N_24647,N_24715);
or UO_73 (O_73,N_24704,N_24669);
nand UO_74 (O_74,N_24599,N_24744);
and UO_75 (O_75,N_24816,N_24607);
nor UO_76 (O_76,N_24721,N_24815);
nand UO_77 (O_77,N_24946,N_24615);
or UO_78 (O_78,N_24753,N_24821);
and UO_79 (O_79,N_24622,N_24531);
and UO_80 (O_80,N_24508,N_24929);
or UO_81 (O_81,N_24517,N_24671);
nand UO_82 (O_82,N_24760,N_24817);
nand UO_83 (O_83,N_24942,N_24726);
nor UO_84 (O_84,N_24911,N_24703);
nor UO_85 (O_85,N_24975,N_24852);
xor UO_86 (O_86,N_24602,N_24670);
or UO_87 (O_87,N_24751,N_24637);
or UO_88 (O_88,N_24674,N_24873);
and UO_89 (O_89,N_24754,N_24891);
and UO_90 (O_90,N_24656,N_24954);
nor UO_91 (O_91,N_24892,N_24551);
or UO_92 (O_92,N_24968,N_24592);
nor UO_93 (O_93,N_24652,N_24510);
nor UO_94 (O_94,N_24899,N_24782);
or UO_95 (O_95,N_24783,N_24988);
nor UO_96 (O_96,N_24841,N_24994);
nor UO_97 (O_97,N_24677,N_24720);
xor UO_98 (O_98,N_24750,N_24675);
and UO_99 (O_99,N_24960,N_24958);
and UO_100 (O_100,N_24535,N_24516);
or UO_101 (O_101,N_24708,N_24749);
and UO_102 (O_102,N_24545,N_24734);
xor UO_103 (O_103,N_24511,N_24814);
nand UO_104 (O_104,N_24790,N_24537);
or UO_105 (O_105,N_24640,N_24792);
or UO_106 (O_106,N_24540,N_24764);
nor UO_107 (O_107,N_24616,N_24743);
nor UO_108 (O_108,N_24653,N_24688);
nor UO_109 (O_109,N_24680,N_24871);
or UO_110 (O_110,N_24741,N_24978);
or UO_111 (O_111,N_24863,N_24919);
or UO_112 (O_112,N_24700,N_24806);
and UO_113 (O_113,N_24835,N_24574);
and UO_114 (O_114,N_24979,N_24541);
xor UO_115 (O_115,N_24718,N_24985);
or UO_116 (O_116,N_24575,N_24706);
nor UO_117 (O_117,N_24756,N_24842);
xor UO_118 (O_118,N_24605,N_24921);
or UO_119 (O_119,N_24591,N_24822);
or UO_120 (O_120,N_24546,N_24855);
nor UO_121 (O_121,N_24931,N_24724);
nor UO_122 (O_122,N_24926,N_24732);
and UO_123 (O_123,N_24882,N_24774);
and UO_124 (O_124,N_24924,N_24736);
nor UO_125 (O_125,N_24533,N_24578);
nand UO_126 (O_126,N_24904,N_24559);
nor UO_127 (O_127,N_24557,N_24643);
or UO_128 (O_128,N_24987,N_24568);
xnor UO_129 (O_129,N_24916,N_24933);
nor UO_130 (O_130,N_24866,N_24563);
and UO_131 (O_131,N_24735,N_24784);
nor UO_132 (O_132,N_24710,N_24623);
nand UO_133 (O_133,N_24739,N_24897);
nand UO_134 (O_134,N_24927,N_24827);
or UO_135 (O_135,N_24881,N_24594);
and UO_136 (O_136,N_24779,N_24502);
nand UO_137 (O_137,N_24507,N_24519);
nand UO_138 (O_138,N_24520,N_24672);
nand UO_139 (O_139,N_24707,N_24878);
nand UO_140 (O_140,N_24799,N_24597);
nor UO_141 (O_141,N_24862,N_24717);
nand UO_142 (O_142,N_24585,N_24730);
or UO_143 (O_143,N_24947,N_24544);
nor UO_144 (O_144,N_24634,N_24570);
nor UO_145 (O_145,N_24830,N_24626);
xnor UO_146 (O_146,N_24609,N_24613);
nor UO_147 (O_147,N_24795,N_24773);
nor UO_148 (O_148,N_24769,N_24604);
and UO_149 (O_149,N_24738,N_24772);
nor UO_150 (O_150,N_24571,N_24534);
xnor UO_151 (O_151,N_24650,N_24631);
nor UO_152 (O_152,N_24617,N_24780);
nor UO_153 (O_153,N_24854,N_24807);
nor UO_154 (O_154,N_24812,N_24625);
nor UO_155 (O_155,N_24633,N_24698);
or UO_156 (O_156,N_24939,N_24989);
or UO_157 (O_157,N_24785,N_24577);
xnor UO_158 (O_158,N_24819,N_24860);
or UO_159 (O_159,N_24912,N_24962);
nand UO_160 (O_160,N_24917,N_24991);
and UO_161 (O_161,N_24883,N_24610);
or UO_162 (O_162,N_24888,N_24789);
nand UO_163 (O_163,N_24972,N_24908);
and UO_164 (O_164,N_24768,N_24984);
nor UO_165 (O_165,N_24553,N_24763);
xnor UO_166 (O_166,N_24839,N_24538);
or UO_167 (O_167,N_24587,N_24527);
and UO_168 (O_168,N_24771,N_24660);
nand UO_169 (O_169,N_24745,N_24651);
or UO_170 (O_170,N_24847,N_24971);
nor UO_171 (O_171,N_24567,N_24853);
nor UO_172 (O_172,N_24521,N_24982);
nor UO_173 (O_173,N_24748,N_24711);
nor UO_174 (O_174,N_24907,N_24943);
nor UO_175 (O_175,N_24561,N_24885);
nand UO_176 (O_176,N_24580,N_24661);
nand UO_177 (O_177,N_24894,N_24886);
nand UO_178 (O_178,N_24856,N_24525);
and UO_179 (O_179,N_24843,N_24618);
or UO_180 (O_180,N_24781,N_24953);
nand UO_181 (O_181,N_24918,N_24658);
and UO_182 (O_182,N_24934,N_24589);
xnor UO_183 (O_183,N_24965,N_24693);
and UO_184 (O_184,N_24539,N_24667);
nor UO_185 (O_185,N_24999,N_24777);
or UO_186 (O_186,N_24859,N_24595);
nand UO_187 (O_187,N_24800,N_24963);
nand UO_188 (O_188,N_24910,N_24747);
and UO_189 (O_189,N_24828,N_24683);
nand UO_190 (O_190,N_24614,N_24797);
nor UO_191 (O_191,N_24526,N_24981);
nor UO_192 (O_192,N_24608,N_24716);
and UO_193 (O_193,N_24690,N_24823);
or UO_194 (O_194,N_24588,N_24596);
xor UO_195 (O_195,N_24729,N_24501);
nand UO_196 (O_196,N_24556,N_24685);
or UO_197 (O_197,N_24875,N_24505);
nand UO_198 (O_198,N_24903,N_24928);
or UO_199 (O_199,N_24956,N_24668);
nand UO_200 (O_200,N_24973,N_24787);
xnor UO_201 (O_201,N_24950,N_24900);
and UO_202 (O_202,N_24536,N_24619);
xnor UO_203 (O_203,N_24712,N_24523);
or UO_204 (O_204,N_24733,N_24583);
or UO_205 (O_205,N_24692,N_24788);
or UO_206 (O_206,N_24512,N_24565);
and UO_207 (O_207,N_24503,N_24673);
or UO_208 (O_208,N_24778,N_24612);
or UO_209 (O_209,N_24967,N_24898);
nand UO_210 (O_210,N_24506,N_24714);
nor UO_211 (O_211,N_24980,N_24996);
nor UO_212 (O_212,N_24813,N_24603);
nand UO_213 (O_213,N_24558,N_24665);
nor UO_214 (O_214,N_24820,N_24846);
nand UO_215 (O_215,N_24775,N_24838);
nand UO_216 (O_216,N_24686,N_24796);
or UO_217 (O_217,N_24872,N_24699);
and UO_218 (O_218,N_24740,N_24725);
nand UO_219 (O_219,N_24893,N_24937);
xor UO_220 (O_220,N_24564,N_24584);
xor UO_221 (O_221,N_24606,N_24509);
or UO_222 (O_222,N_24746,N_24876);
nand UO_223 (O_223,N_24642,N_24818);
nor UO_224 (O_224,N_24696,N_24620);
nand UO_225 (O_225,N_24845,N_24697);
nand UO_226 (O_226,N_24974,N_24913);
or UO_227 (O_227,N_24731,N_24695);
and UO_228 (O_228,N_24951,N_24865);
and UO_229 (O_229,N_24998,N_24684);
or UO_230 (O_230,N_24752,N_24761);
xor UO_231 (O_231,N_24848,N_24645);
xor UO_232 (O_232,N_24805,N_24664);
and UO_233 (O_233,N_24719,N_24770);
or UO_234 (O_234,N_24840,N_24518);
or UO_235 (O_235,N_24543,N_24867);
and UO_236 (O_236,N_24666,N_24676);
nor UO_237 (O_237,N_24993,N_24923);
nand UO_238 (O_238,N_24844,N_24582);
nor UO_239 (O_239,N_24868,N_24851);
nor UO_240 (O_240,N_24727,N_24961);
nor UO_241 (O_241,N_24524,N_24801);
nor UO_242 (O_242,N_24632,N_24566);
or UO_243 (O_243,N_24986,N_24858);
nand UO_244 (O_244,N_24938,N_24532);
xor UO_245 (O_245,N_24624,N_24515);
and UO_246 (O_246,N_24920,N_24681);
or UO_247 (O_247,N_24964,N_24793);
and UO_248 (O_248,N_24742,N_24959);
and UO_249 (O_249,N_24709,N_24802);
or UO_250 (O_250,N_24701,N_24807);
or UO_251 (O_251,N_24662,N_24937);
nor UO_252 (O_252,N_24700,N_24780);
and UO_253 (O_253,N_24564,N_24929);
xor UO_254 (O_254,N_24672,N_24689);
nor UO_255 (O_255,N_24742,N_24773);
and UO_256 (O_256,N_24905,N_24951);
and UO_257 (O_257,N_24871,N_24597);
nand UO_258 (O_258,N_24859,N_24733);
and UO_259 (O_259,N_24962,N_24838);
nor UO_260 (O_260,N_24901,N_24653);
xnor UO_261 (O_261,N_24695,N_24912);
nor UO_262 (O_262,N_24566,N_24694);
nor UO_263 (O_263,N_24869,N_24615);
nand UO_264 (O_264,N_24926,N_24935);
nand UO_265 (O_265,N_24622,N_24795);
or UO_266 (O_266,N_24928,N_24979);
nand UO_267 (O_267,N_24698,N_24780);
or UO_268 (O_268,N_24630,N_24931);
and UO_269 (O_269,N_24688,N_24998);
or UO_270 (O_270,N_24623,N_24573);
or UO_271 (O_271,N_24604,N_24594);
or UO_272 (O_272,N_24576,N_24861);
or UO_273 (O_273,N_24782,N_24850);
nand UO_274 (O_274,N_24725,N_24788);
or UO_275 (O_275,N_24764,N_24990);
nor UO_276 (O_276,N_24622,N_24657);
and UO_277 (O_277,N_24753,N_24701);
nand UO_278 (O_278,N_24845,N_24519);
nand UO_279 (O_279,N_24749,N_24965);
and UO_280 (O_280,N_24603,N_24936);
and UO_281 (O_281,N_24584,N_24691);
nand UO_282 (O_282,N_24945,N_24997);
nor UO_283 (O_283,N_24696,N_24949);
nand UO_284 (O_284,N_24679,N_24572);
or UO_285 (O_285,N_24727,N_24681);
and UO_286 (O_286,N_24863,N_24628);
and UO_287 (O_287,N_24938,N_24616);
nand UO_288 (O_288,N_24754,N_24892);
and UO_289 (O_289,N_24944,N_24543);
nand UO_290 (O_290,N_24928,N_24759);
and UO_291 (O_291,N_24939,N_24766);
nand UO_292 (O_292,N_24923,N_24628);
nand UO_293 (O_293,N_24926,N_24860);
nand UO_294 (O_294,N_24562,N_24732);
and UO_295 (O_295,N_24948,N_24979);
and UO_296 (O_296,N_24537,N_24735);
nand UO_297 (O_297,N_24797,N_24764);
or UO_298 (O_298,N_24774,N_24809);
and UO_299 (O_299,N_24645,N_24719);
and UO_300 (O_300,N_24694,N_24749);
nand UO_301 (O_301,N_24647,N_24609);
and UO_302 (O_302,N_24995,N_24513);
and UO_303 (O_303,N_24733,N_24605);
nand UO_304 (O_304,N_24781,N_24918);
xnor UO_305 (O_305,N_24760,N_24996);
nand UO_306 (O_306,N_24644,N_24684);
nor UO_307 (O_307,N_24958,N_24653);
nand UO_308 (O_308,N_24733,N_24666);
nand UO_309 (O_309,N_24821,N_24993);
or UO_310 (O_310,N_24530,N_24615);
or UO_311 (O_311,N_24786,N_24513);
and UO_312 (O_312,N_24821,N_24792);
nand UO_313 (O_313,N_24827,N_24831);
and UO_314 (O_314,N_24739,N_24953);
and UO_315 (O_315,N_24776,N_24819);
nand UO_316 (O_316,N_24676,N_24617);
nor UO_317 (O_317,N_24975,N_24640);
nor UO_318 (O_318,N_24820,N_24882);
or UO_319 (O_319,N_24686,N_24565);
nand UO_320 (O_320,N_24804,N_24680);
nor UO_321 (O_321,N_24855,N_24582);
nor UO_322 (O_322,N_24784,N_24592);
and UO_323 (O_323,N_24683,N_24564);
nor UO_324 (O_324,N_24993,N_24599);
nor UO_325 (O_325,N_24661,N_24785);
or UO_326 (O_326,N_24513,N_24699);
nor UO_327 (O_327,N_24980,N_24593);
nor UO_328 (O_328,N_24850,N_24973);
xnor UO_329 (O_329,N_24826,N_24974);
nand UO_330 (O_330,N_24559,N_24617);
nand UO_331 (O_331,N_24815,N_24798);
and UO_332 (O_332,N_24733,N_24777);
nor UO_333 (O_333,N_24858,N_24742);
nor UO_334 (O_334,N_24664,N_24852);
nor UO_335 (O_335,N_24884,N_24670);
xor UO_336 (O_336,N_24680,N_24913);
nand UO_337 (O_337,N_24826,N_24967);
nor UO_338 (O_338,N_24892,N_24697);
or UO_339 (O_339,N_24976,N_24859);
nor UO_340 (O_340,N_24527,N_24606);
and UO_341 (O_341,N_24683,N_24697);
xor UO_342 (O_342,N_24860,N_24687);
nor UO_343 (O_343,N_24638,N_24628);
nor UO_344 (O_344,N_24919,N_24803);
xor UO_345 (O_345,N_24637,N_24657);
or UO_346 (O_346,N_24896,N_24765);
or UO_347 (O_347,N_24833,N_24670);
nor UO_348 (O_348,N_24814,N_24807);
nand UO_349 (O_349,N_24577,N_24701);
nand UO_350 (O_350,N_24503,N_24665);
and UO_351 (O_351,N_24961,N_24937);
nor UO_352 (O_352,N_24730,N_24827);
and UO_353 (O_353,N_24770,N_24961);
or UO_354 (O_354,N_24723,N_24832);
nor UO_355 (O_355,N_24961,N_24537);
nand UO_356 (O_356,N_24775,N_24674);
nand UO_357 (O_357,N_24725,N_24915);
or UO_358 (O_358,N_24759,N_24643);
and UO_359 (O_359,N_24744,N_24877);
or UO_360 (O_360,N_24609,N_24662);
nor UO_361 (O_361,N_24771,N_24580);
nand UO_362 (O_362,N_24852,N_24816);
and UO_363 (O_363,N_24721,N_24601);
or UO_364 (O_364,N_24538,N_24584);
xor UO_365 (O_365,N_24806,N_24542);
and UO_366 (O_366,N_24600,N_24598);
nor UO_367 (O_367,N_24929,N_24969);
nor UO_368 (O_368,N_24871,N_24639);
and UO_369 (O_369,N_24699,N_24763);
or UO_370 (O_370,N_24898,N_24686);
nand UO_371 (O_371,N_24607,N_24941);
and UO_372 (O_372,N_24649,N_24943);
nor UO_373 (O_373,N_24747,N_24653);
and UO_374 (O_374,N_24696,N_24648);
and UO_375 (O_375,N_24936,N_24911);
nand UO_376 (O_376,N_24901,N_24863);
nand UO_377 (O_377,N_24686,N_24559);
nand UO_378 (O_378,N_24885,N_24944);
nor UO_379 (O_379,N_24931,N_24912);
and UO_380 (O_380,N_24794,N_24600);
and UO_381 (O_381,N_24656,N_24700);
nand UO_382 (O_382,N_24654,N_24664);
or UO_383 (O_383,N_24608,N_24817);
and UO_384 (O_384,N_24807,N_24994);
or UO_385 (O_385,N_24652,N_24557);
nand UO_386 (O_386,N_24725,N_24666);
nand UO_387 (O_387,N_24891,N_24744);
and UO_388 (O_388,N_24767,N_24633);
nand UO_389 (O_389,N_24904,N_24981);
or UO_390 (O_390,N_24785,N_24769);
nand UO_391 (O_391,N_24679,N_24501);
nor UO_392 (O_392,N_24611,N_24766);
and UO_393 (O_393,N_24966,N_24757);
or UO_394 (O_394,N_24799,N_24636);
and UO_395 (O_395,N_24625,N_24594);
nor UO_396 (O_396,N_24898,N_24513);
nand UO_397 (O_397,N_24556,N_24541);
nand UO_398 (O_398,N_24890,N_24949);
nand UO_399 (O_399,N_24848,N_24798);
nor UO_400 (O_400,N_24984,N_24932);
or UO_401 (O_401,N_24589,N_24512);
xnor UO_402 (O_402,N_24542,N_24724);
nor UO_403 (O_403,N_24703,N_24574);
xnor UO_404 (O_404,N_24940,N_24662);
nor UO_405 (O_405,N_24898,N_24519);
and UO_406 (O_406,N_24702,N_24543);
nand UO_407 (O_407,N_24912,N_24635);
nor UO_408 (O_408,N_24895,N_24814);
or UO_409 (O_409,N_24618,N_24804);
and UO_410 (O_410,N_24814,N_24696);
nand UO_411 (O_411,N_24625,N_24897);
and UO_412 (O_412,N_24735,N_24906);
or UO_413 (O_413,N_24586,N_24553);
or UO_414 (O_414,N_24540,N_24553);
nor UO_415 (O_415,N_24694,N_24970);
and UO_416 (O_416,N_24879,N_24979);
and UO_417 (O_417,N_24900,N_24838);
and UO_418 (O_418,N_24623,N_24794);
or UO_419 (O_419,N_24532,N_24992);
nand UO_420 (O_420,N_24846,N_24763);
nor UO_421 (O_421,N_24526,N_24614);
or UO_422 (O_422,N_24910,N_24780);
and UO_423 (O_423,N_24602,N_24587);
nor UO_424 (O_424,N_24951,N_24744);
nand UO_425 (O_425,N_24567,N_24683);
and UO_426 (O_426,N_24970,N_24547);
nor UO_427 (O_427,N_24712,N_24765);
nand UO_428 (O_428,N_24535,N_24514);
nor UO_429 (O_429,N_24794,N_24720);
or UO_430 (O_430,N_24782,N_24702);
nor UO_431 (O_431,N_24841,N_24586);
or UO_432 (O_432,N_24514,N_24877);
nor UO_433 (O_433,N_24599,N_24600);
nor UO_434 (O_434,N_24940,N_24844);
or UO_435 (O_435,N_24593,N_24933);
nand UO_436 (O_436,N_24999,N_24673);
and UO_437 (O_437,N_24922,N_24707);
and UO_438 (O_438,N_24776,N_24829);
nand UO_439 (O_439,N_24598,N_24780);
and UO_440 (O_440,N_24587,N_24839);
or UO_441 (O_441,N_24749,N_24839);
nor UO_442 (O_442,N_24787,N_24722);
xnor UO_443 (O_443,N_24839,N_24942);
nand UO_444 (O_444,N_24812,N_24527);
and UO_445 (O_445,N_24950,N_24934);
nand UO_446 (O_446,N_24849,N_24542);
and UO_447 (O_447,N_24864,N_24762);
and UO_448 (O_448,N_24569,N_24649);
nand UO_449 (O_449,N_24933,N_24603);
xnor UO_450 (O_450,N_24608,N_24724);
or UO_451 (O_451,N_24817,N_24804);
and UO_452 (O_452,N_24526,N_24560);
nand UO_453 (O_453,N_24535,N_24965);
nand UO_454 (O_454,N_24993,N_24854);
or UO_455 (O_455,N_24638,N_24707);
nor UO_456 (O_456,N_24528,N_24692);
nand UO_457 (O_457,N_24820,N_24737);
nand UO_458 (O_458,N_24824,N_24628);
nand UO_459 (O_459,N_24605,N_24591);
or UO_460 (O_460,N_24925,N_24866);
and UO_461 (O_461,N_24760,N_24823);
nor UO_462 (O_462,N_24580,N_24780);
and UO_463 (O_463,N_24986,N_24812);
nand UO_464 (O_464,N_24991,N_24901);
nor UO_465 (O_465,N_24679,N_24599);
or UO_466 (O_466,N_24988,N_24885);
nand UO_467 (O_467,N_24782,N_24657);
nand UO_468 (O_468,N_24741,N_24881);
nor UO_469 (O_469,N_24840,N_24732);
and UO_470 (O_470,N_24807,N_24828);
and UO_471 (O_471,N_24702,N_24779);
nand UO_472 (O_472,N_24943,N_24792);
nor UO_473 (O_473,N_24593,N_24541);
nor UO_474 (O_474,N_24935,N_24941);
and UO_475 (O_475,N_24546,N_24701);
and UO_476 (O_476,N_24770,N_24850);
and UO_477 (O_477,N_24755,N_24952);
xnor UO_478 (O_478,N_24892,N_24663);
nor UO_479 (O_479,N_24876,N_24921);
xnor UO_480 (O_480,N_24917,N_24979);
or UO_481 (O_481,N_24758,N_24951);
and UO_482 (O_482,N_24614,N_24915);
nand UO_483 (O_483,N_24825,N_24739);
nor UO_484 (O_484,N_24846,N_24787);
nand UO_485 (O_485,N_24509,N_24800);
nand UO_486 (O_486,N_24632,N_24720);
xor UO_487 (O_487,N_24809,N_24718);
nor UO_488 (O_488,N_24628,N_24579);
nor UO_489 (O_489,N_24507,N_24737);
xnor UO_490 (O_490,N_24869,N_24734);
or UO_491 (O_491,N_24558,N_24786);
and UO_492 (O_492,N_24729,N_24594);
or UO_493 (O_493,N_24939,N_24502);
nand UO_494 (O_494,N_24840,N_24791);
nand UO_495 (O_495,N_24920,N_24648);
xor UO_496 (O_496,N_24529,N_24537);
nor UO_497 (O_497,N_24902,N_24849);
and UO_498 (O_498,N_24544,N_24821);
nor UO_499 (O_499,N_24856,N_24673);
or UO_500 (O_500,N_24548,N_24907);
and UO_501 (O_501,N_24895,N_24992);
nor UO_502 (O_502,N_24724,N_24795);
nand UO_503 (O_503,N_24951,N_24759);
xor UO_504 (O_504,N_24981,N_24976);
nor UO_505 (O_505,N_24619,N_24625);
and UO_506 (O_506,N_24554,N_24742);
xor UO_507 (O_507,N_24897,N_24920);
and UO_508 (O_508,N_24513,N_24855);
or UO_509 (O_509,N_24534,N_24643);
nor UO_510 (O_510,N_24885,N_24560);
xor UO_511 (O_511,N_24794,N_24855);
and UO_512 (O_512,N_24638,N_24528);
nor UO_513 (O_513,N_24717,N_24913);
and UO_514 (O_514,N_24726,N_24972);
nand UO_515 (O_515,N_24937,N_24987);
and UO_516 (O_516,N_24907,N_24928);
or UO_517 (O_517,N_24953,N_24885);
and UO_518 (O_518,N_24823,N_24800);
or UO_519 (O_519,N_24990,N_24915);
nor UO_520 (O_520,N_24758,N_24902);
and UO_521 (O_521,N_24573,N_24896);
nor UO_522 (O_522,N_24869,N_24580);
nand UO_523 (O_523,N_24540,N_24645);
and UO_524 (O_524,N_24737,N_24673);
nand UO_525 (O_525,N_24850,N_24931);
nor UO_526 (O_526,N_24903,N_24987);
nor UO_527 (O_527,N_24611,N_24872);
xor UO_528 (O_528,N_24862,N_24752);
nand UO_529 (O_529,N_24619,N_24527);
nand UO_530 (O_530,N_24732,N_24968);
or UO_531 (O_531,N_24949,N_24967);
nand UO_532 (O_532,N_24716,N_24584);
xor UO_533 (O_533,N_24768,N_24692);
xnor UO_534 (O_534,N_24873,N_24630);
nor UO_535 (O_535,N_24635,N_24839);
nand UO_536 (O_536,N_24687,N_24615);
or UO_537 (O_537,N_24544,N_24944);
or UO_538 (O_538,N_24911,N_24886);
nor UO_539 (O_539,N_24861,N_24840);
or UO_540 (O_540,N_24506,N_24827);
or UO_541 (O_541,N_24560,N_24605);
or UO_542 (O_542,N_24624,N_24824);
xnor UO_543 (O_543,N_24950,N_24990);
and UO_544 (O_544,N_24932,N_24729);
or UO_545 (O_545,N_24744,N_24701);
nor UO_546 (O_546,N_24793,N_24610);
and UO_547 (O_547,N_24918,N_24951);
nor UO_548 (O_548,N_24903,N_24846);
and UO_549 (O_549,N_24701,N_24769);
nand UO_550 (O_550,N_24649,N_24537);
or UO_551 (O_551,N_24902,N_24782);
nor UO_552 (O_552,N_24811,N_24630);
or UO_553 (O_553,N_24588,N_24934);
nand UO_554 (O_554,N_24965,N_24515);
and UO_555 (O_555,N_24818,N_24553);
nor UO_556 (O_556,N_24747,N_24958);
or UO_557 (O_557,N_24628,N_24856);
or UO_558 (O_558,N_24633,N_24923);
and UO_559 (O_559,N_24641,N_24880);
nor UO_560 (O_560,N_24672,N_24700);
or UO_561 (O_561,N_24657,N_24525);
nand UO_562 (O_562,N_24750,N_24606);
or UO_563 (O_563,N_24791,N_24511);
nor UO_564 (O_564,N_24644,N_24655);
nor UO_565 (O_565,N_24926,N_24701);
nor UO_566 (O_566,N_24830,N_24968);
nand UO_567 (O_567,N_24716,N_24544);
or UO_568 (O_568,N_24692,N_24942);
or UO_569 (O_569,N_24801,N_24500);
nor UO_570 (O_570,N_24740,N_24610);
nor UO_571 (O_571,N_24529,N_24766);
and UO_572 (O_572,N_24905,N_24742);
xor UO_573 (O_573,N_24551,N_24759);
nor UO_574 (O_574,N_24651,N_24831);
or UO_575 (O_575,N_24975,N_24559);
and UO_576 (O_576,N_24694,N_24998);
nand UO_577 (O_577,N_24751,N_24857);
nand UO_578 (O_578,N_24823,N_24912);
nor UO_579 (O_579,N_24956,N_24513);
or UO_580 (O_580,N_24581,N_24984);
and UO_581 (O_581,N_24616,N_24521);
and UO_582 (O_582,N_24696,N_24673);
or UO_583 (O_583,N_24886,N_24777);
nand UO_584 (O_584,N_24805,N_24548);
or UO_585 (O_585,N_24522,N_24549);
and UO_586 (O_586,N_24913,N_24666);
nor UO_587 (O_587,N_24828,N_24934);
or UO_588 (O_588,N_24508,N_24987);
or UO_589 (O_589,N_24995,N_24611);
nor UO_590 (O_590,N_24861,N_24782);
or UO_591 (O_591,N_24847,N_24637);
nand UO_592 (O_592,N_24928,N_24590);
and UO_593 (O_593,N_24971,N_24717);
and UO_594 (O_594,N_24572,N_24641);
xnor UO_595 (O_595,N_24803,N_24504);
nand UO_596 (O_596,N_24966,N_24803);
or UO_597 (O_597,N_24869,N_24814);
or UO_598 (O_598,N_24613,N_24966);
xor UO_599 (O_599,N_24928,N_24910);
or UO_600 (O_600,N_24652,N_24817);
and UO_601 (O_601,N_24918,N_24521);
and UO_602 (O_602,N_24895,N_24784);
nor UO_603 (O_603,N_24955,N_24575);
nor UO_604 (O_604,N_24726,N_24791);
and UO_605 (O_605,N_24697,N_24689);
or UO_606 (O_606,N_24592,N_24512);
nor UO_607 (O_607,N_24568,N_24939);
or UO_608 (O_608,N_24953,N_24890);
nor UO_609 (O_609,N_24761,N_24711);
xor UO_610 (O_610,N_24798,N_24819);
nor UO_611 (O_611,N_24601,N_24878);
and UO_612 (O_612,N_24697,N_24827);
or UO_613 (O_613,N_24639,N_24681);
and UO_614 (O_614,N_24559,N_24758);
nand UO_615 (O_615,N_24600,N_24547);
xnor UO_616 (O_616,N_24776,N_24753);
nor UO_617 (O_617,N_24790,N_24958);
or UO_618 (O_618,N_24571,N_24859);
or UO_619 (O_619,N_24833,N_24745);
or UO_620 (O_620,N_24861,N_24860);
and UO_621 (O_621,N_24635,N_24544);
xnor UO_622 (O_622,N_24560,N_24570);
or UO_623 (O_623,N_24640,N_24702);
nand UO_624 (O_624,N_24853,N_24513);
nand UO_625 (O_625,N_24903,N_24731);
nor UO_626 (O_626,N_24745,N_24695);
nand UO_627 (O_627,N_24671,N_24862);
nand UO_628 (O_628,N_24808,N_24779);
nand UO_629 (O_629,N_24826,N_24689);
nand UO_630 (O_630,N_24677,N_24853);
xor UO_631 (O_631,N_24866,N_24519);
xnor UO_632 (O_632,N_24993,N_24546);
nand UO_633 (O_633,N_24561,N_24767);
or UO_634 (O_634,N_24562,N_24723);
nor UO_635 (O_635,N_24972,N_24936);
xnor UO_636 (O_636,N_24610,N_24972);
nand UO_637 (O_637,N_24966,N_24638);
or UO_638 (O_638,N_24625,N_24968);
nand UO_639 (O_639,N_24983,N_24740);
and UO_640 (O_640,N_24974,N_24766);
or UO_641 (O_641,N_24881,N_24570);
and UO_642 (O_642,N_24883,N_24863);
nor UO_643 (O_643,N_24875,N_24637);
nand UO_644 (O_644,N_24829,N_24958);
nand UO_645 (O_645,N_24682,N_24667);
nand UO_646 (O_646,N_24785,N_24560);
and UO_647 (O_647,N_24862,N_24587);
nor UO_648 (O_648,N_24701,N_24533);
nor UO_649 (O_649,N_24765,N_24511);
nand UO_650 (O_650,N_24726,N_24933);
and UO_651 (O_651,N_24681,N_24761);
nand UO_652 (O_652,N_24529,N_24503);
nor UO_653 (O_653,N_24634,N_24970);
xnor UO_654 (O_654,N_24667,N_24646);
nor UO_655 (O_655,N_24721,N_24725);
nand UO_656 (O_656,N_24949,N_24936);
nand UO_657 (O_657,N_24785,N_24685);
and UO_658 (O_658,N_24534,N_24893);
nand UO_659 (O_659,N_24957,N_24629);
and UO_660 (O_660,N_24638,N_24998);
nand UO_661 (O_661,N_24870,N_24830);
nor UO_662 (O_662,N_24683,N_24775);
xnor UO_663 (O_663,N_24827,N_24696);
and UO_664 (O_664,N_24543,N_24993);
and UO_665 (O_665,N_24967,N_24882);
xnor UO_666 (O_666,N_24993,N_24745);
nand UO_667 (O_667,N_24815,N_24552);
or UO_668 (O_668,N_24984,N_24861);
xnor UO_669 (O_669,N_24764,N_24607);
nor UO_670 (O_670,N_24951,N_24515);
nand UO_671 (O_671,N_24747,N_24681);
xnor UO_672 (O_672,N_24725,N_24805);
or UO_673 (O_673,N_24940,N_24952);
xor UO_674 (O_674,N_24870,N_24811);
xnor UO_675 (O_675,N_24847,N_24607);
and UO_676 (O_676,N_24875,N_24641);
and UO_677 (O_677,N_24885,N_24875);
and UO_678 (O_678,N_24603,N_24706);
nand UO_679 (O_679,N_24992,N_24997);
and UO_680 (O_680,N_24634,N_24560);
nor UO_681 (O_681,N_24519,N_24668);
and UO_682 (O_682,N_24876,N_24631);
nand UO_683 (O_683,N_24669,N_24762);
and UO_684 (O_684,N_24553,N_24904);
nand UO_685 (O_685,N_24507,N_24585);
nor UO_686 (O_686,N_24776,N_24970);
nand UO_687 (O_687,N_24947,N_24903);
nor UO_688 (O_688,N_24527,N_24624);
and UO_689 (O_689,N_24966,N_24837);
and UO_690 (O_690,N_24898,N_24926);
and UO_691 (O_691,N_24810,N_24927);
and UO_692 (O_692,N_24549,N_24995);
nor UO_693 (O_693,N_24765,N_24958);
xor UO_694 (O_694,N_24510,N_24997);
nand UO_695 (O_695,N_24633,N_24931);
and UO_696 (O_696,N_24863,N_24659);
nand UO_697 (O_697,N_24900,N_24958);
xnor UO_698 (O_698,N_24923,N_24925);
xnor UO_699 (O_699,N_24663,N_24673);
nor UO_700 (O_700,N_24530,N_24905);
nand UO_701 (O_701,N_24508,N_24669);
and UO_702 (O_702,N_24706,N_24669);
and UO_703 (O_703,N_24518,N_24865);
or UO_704 (O_704,N_24993,N_24642);
and UO_705 (O_705,N_24998,N_24766);
or UO_706 (O_706,N_24711,N_24760);
nand UO_707 (O_707,N_24838,N_24500);
nor UO_708 (O_708,N_24714,N_24502);
nand UO_709 (O_709,N_24957,N_24586);
and UO_710 (O_710,N_24591,N_24823);
or UO_711 (O_711,N_24850,N_24832);
nand UO_712 (O_712,N_24564,N_24961);
or UO_713 (O_713,N_24669,N_24866);
or UO_714 (O_714,N_24901,N_24792);
and UO_715 (O_715,N_24506,N_24867);
nor UO_716 (O_716,N_24661,N_24677);
or UO_717 (O_717,N_24612,N_24875);
nand UO_718 (O_718,N_24859,N_24796);
nand UO_719 (O_719,N_24628,N_24567);
xor UO_720 (O_720,N_24520,N_24556);
and UO_721 (O_721,N_24753,N_24682);
nor UO_722 (O_722,N_24601,N_24907);
and UO_723 (O_723,N_24519,N_24851);
nor UO_724 (O_724,N_24963,N_24787);
nor UO_725 (O_725,N_24634,N_24685);
or UO_726 (O_726,N_24860,N_24546);
and UO_727 (O_727,N_24733,N_24952);
and UO_728 (O_728,N_24784,N_24708);
xor UO_729 (O_729,N_24563,N_24646);
nor UO_730 (O_730,N_24942,N_24712);
and UO_731 (O_731,N_24819,N_24744);
and UO_732 (O_732,N_24921,N_24532);
and UO_733 (O_733,N_24721,N_24811);
nand UO_734 (O_734,N_24548,N_24605);
xnor UO_735 (O_735,N_24750,N_24637);
nand UO_736 (O_736,N_24692,N_24624);
nor UO_737 (O_737,N_24803,N_24558);
nand UO_738 (O_738,N_24692,N_24536);
or UO_739 (O_739,N_24886,N_24933);
or UO_740 (O_740,N_24641,N_24538);
nor UO_741 (O_741,N_24711,N_24745);
and UO_742 (O_742,N_24845,N_24694);
or UO_743 (O_743,N_24676,N_24863);
nand UO_744 (O_744,N_24773,N_24805);
nor UO_745 (O_745,N_24856,N_24912);
and UO_746 (O_746,N_24983,N_24835);
or UO_747 (O_747,N_24789,N_24963);
nor UO_748 (O_748,N_24577,N_24819);
and UO_749 (O_749,N_24518,N_24702);
nor UO_750 (O_750,N_24917,N_24799);
nand UO_751 (O_751,N_24778,N_24705);
and UO_752 (O_752,N_24602,N_24801);
nand UO_753 (O_753,N_24541,N_24822);
or UO_754 (O_754,N_24692,N_24965);
or UO_755 (O_755,N_24979,N_24779);
and UO_756 (O_756,N_24538,N_24924);
nand UO_757 (O_757,N_24878,N_24824);
nor UO_758 (O_758,N_24627,N_24535);
or UO_759 (O_759,N_24848,N_24824);
nor UO_760 (O_760,N_24797,N_24914);
nor UO_761 (O_761,N_24623,N_24920);
xor UO_762 (O_762,N_24725,N_24832);
and UO_763 (O_763,N_24613,N_24766);
and UO_764 (O_764,N_24844,N_24793);
nor UO_765 (O_765,N_24799,N_24679);
nor UO_766 (O_766,N_24639,N_24597);
nor UO_767 (O_767,N_24534,N_24913);
nor UO_768 (O_768,N_24996,N_24999);
nor UO_769 (O_769,N_24754,N_24859);
xor UO_770 (O_770,N_24986,N_24674);
or UO_771 (O_771,N_24794,N_24899);
or UO_772 (O_772,N_24773,N_24710);
xor UO_773 (O_773,N_24755,N_24913);
nor UO_774 (O_774,N_24645,N_24658);
nor UO_775 (O_775,N_24971,N_24864);
and UO_776 (O_776,N_24855,N_24747);
or UO_777 (O_777,N_24519,N_24830);
nand UO_778 (O_778,N_24568,N_24924);
nand UO_779 (O_779,N_24548,N_24899);
xnor UO_780 (O_780,N_24762,N_24883);
nand UO_781 (O_781,N_24711,N_24591);
nand UO_782 (O_782,N_24664,N_24709);
nand UO_783 (O_783,N_24562,N_24660);
or UO_784 (O_784,N_24876,N_24560);
or UO_785 (O_785,N_24728,N_24845);
xor UO_786 (O_786,N_24941,N_24611);
or UO_787 (O_787,N_24786,N_24915);
or UO_788 (O_788,N_24660,N_24556);
or UO_789 (O_789,N_24661,N_24790);
nor UO_790 (O_790,N_24789,N_24818);
nand UO_791 (O_791,N_24600,N_24538);
nand UO_792 (O_792,N_24731,N_24995);
nand UO_793 (O_793,N_24540,N_24560);
or UO_794 (O_794,N_24895,N_24725);
and UO_795 (O_795,N_24554,N_24663);
nor UO_796 (O_796,N_24648,N_24661);
and UO_797 (O_797,N_24851,N_24515);
nor UO_798 (O_798,N_24904,N_24854);
nand UO_799 (O_799,N_24636,N_24574);
nand UO_800 (O_800,N_24604,N_24833);
nor UO_801 (O_801,N_24778,N_24724);
nor UO_802 (O_802,N_24649,N_24955);
and UO_803 (O_803,N_24975,N_24774);
nand UO_804 (O_804,N_24566,N_24727);
and UO_805 (O_805,N_24643,N_24781);
xor UO_806 (O_806,N_24545,N_24643);
xor UO_807 (O_807,N_24670,N_24858);
or UO_808 (O_808,N_24621,N_24882);
or UO_809 (O_809,N_24930,N_24551);
nor UO_810 (O_810,N_24785,N_24888);
nor UO_811 (O_811,N_24738,N_24851);
xnor UO_812 (O_812,N_24977,N_24631);
or UO_813 (O_813,N_24792,N_24986);
nor UO_814 (O_814,N_24627,N_24767);
nor UO_815 (O_815,N_24935,N_24637);
xnor UO_816 (O_816,N_24666,N_24737);
or UO_817 (O_817,N_24549,N_24551);
nor UO_818 (O_818,N_24765,N_24971);
nor UO_819 (O_819,N_24639,N_24889);
or UO_820 (O_820,N_24592,N_24989);
nand UO_821 (O_821,N_24606,N_24975);
nor UO_822 (O_822,N_24846,N_24774);
or UO_823 (O_823,N_24565,N_24698);
and UO_824 (O_824,N_24872,N_24850);
nand UO_825 (O_825,N_24592,N_24686);
nand UO_826 (O_826,N_24938,N_24622);
and UO_827 (O_827,N_24631,N_24686);
nor UO_828 (O_828,N_24632,N_24623);
nand UO_829 (O_829,N_24617,N_24701);
xor UO_830 (O_830,N_24626,N_24637);
or UO_831 (O_831,N_24614,N_24932);
and UO_832 (O_832,N_24840,N_24719);
or UO_833 (O_833,N_24591,N_24933);
or UO_834 (O_834,N_24556,N_24537);
and UO_835 (O_835,N_24852,N_24511);
xor UO_836 (O_836,N_24771,N_24954);
xor UO_837 (O_837,N_24679,N_24911);
nand UO_838 (O_838,N_24977,N_24928);
and UO_839 (O_839,N_24957,N_24537);
and UO_840 (O_840,N_24559,N_24546);
or UO_841 (O_841,N_24657,N_24592);
and UO_842 (O_842,N_24652,N_24538);
xor UO_843 (O_843,N_24774,N_24828);
or UO_844 (O_844,N_24918,N_24587);
nand UO_845 (O_845,N_24861,N_24508);
nand UO_846 (O_846,N_24967,N_24867);
or UO_847 (O_847,N_24568,N_24941);
nand UO_848 (O_848,N_24691,N_24524);
nor UO_849 (O_849,N_24686,N_24930);
nor UO_850 (O_850,N_24638,N_24580);
and UO_851 (O_851,N_24654,N_24779);
nor UO_852 (O_852,N_24524,N_24573);
and UO_853 (O_853,N_24594,N_24524);
nor UO_854 (O_854,N_24869,N_24889);
and UO_855 (O_855,N_24562,N_24816);
nand UO_856 (O_856,N_24908,N_24538);
and UO_857 (O_857,N_24595,N_24708);
nand UO_858 (O_858,N_24625,N_24617);
nor UO_859 (O_859,N_24698,N_24713);
nand UO_860 (O_860,N_24538,N_24980);
xnor UO_861 (O_861,N_24707,N_24784);
nand UO_862 (O_862,N_24654,N_24562);
xnor UO_863 (O_863,N_24556,N_24911);
nand UO_864 (O_864,N_24783,N_24701);
or UO_865 (O_865,N_24555,N_24707);
and UO_866 (O_866,N_24944,N_24697);
nand UO_867 (O_867,N_24661,N_24820);
nor UO_868 (O_868,N_24944,N_24702);
or UO_869 (O_869,N_24859,N_24626);
nor UO_870 (O_870,N_24699,N_24758);
xnor UO_871 (O_871,N_24819,N_24598);
and UO_872 (O_872,N_24900,N_24885);
or UO_873 (O_873,N_24864,N_24679);
nand UO_874 (O_874,N_24763,N_24726);
xor UO_875 (O_875,N_24821,N_24681);
nor UO_876 (O_876,N_24910,N_24759);
nor UO_877 (O_877,N_24600,N_24756);
or UO_878 (O_878,N_24790,N_24768);
nand UO_879 (O_879,N_24789,N_24565);
or UO_880 (O_880,N_24632,N_24962);
or UO_881 (O_881,N_24964,N_24674);
nor UO_882 (O_882,N_24833,N_24824);
nor UO_883 (O_883,N_24591,N_24714);
nor UO_884 (O_884,N_24812,N_24702);
xnor UO_885 (O_885,N_24861,N_24774);
nand UO_886 (O_886,N_24823,N_24901);
nand UO_887 (O_887,N_24839,N_24606);
nand UO_888 (O_888,N_24827,N_24569);
nand UO_889 (O_889,N_24867,N_24913);
or UO_890 (O_890,N_24612,N_24726);
or UO_891 (O_891,N_24533,N_24500);
and UO_892 (O_892,N_24609,N_24776);
and UO_893 (O_893,N_24508,N_24983);
and UO_894 (O_894,N_24548,N_24837);
nand UO_895 (O_895,N_24658,N_24844);
or UO_896 (O_896,N_24584,N_24505);
and UO_897 (O_897,N_24531,N_24597);
nand UO_898 (O_898,N_24799,N_24863);
nor UO_899 (O_899,N_24722,N_24839);
nand UO_900 (O_900,N_24744,N_24688);
or UO_901 (O_901,N_24945,N_24692);
nand UO_902 (O_902,N_24650,N_24855);
nand UO_903 (O_903,N_24671,N_24554);
nor UO_904 (O_904,N_24610,N_24642);
or UO_905 (O_905,N_24757,N_24518);
nand UO_906 (O_906,N_24768,N_24737);
nor UO_907 (O_907,N_24762,N_24973);
or UO_908 (O_908,N_24659,N_24590);
xnor UO_909 (O_909,N_24862,N_24856);
and UO_910 (O_910,N_24827,N_24989);
or UO_911 (O_911,N_24505,N_24630);
nand UO_912 (O_912,N_24808,N_24552);
nand UO_913 (O_913,N_24604,N_24690);
or UO_914 (O_914,N_24629,N_24911);
nand UO_915 (O_915,N_24632,N_24629);
xnor UO_916 (O_916,N_24878,N_24503);
xor UO_917 (O_917,N_24524,N_24673);
nand UO_918 (O_918,N_24973,N_24507);
and UO_919 (O_919,N_24848,N_24532);
nor UO_920 (O_920,N_24867,N_24920);
nand UO_921 (O_921,N_24955,N_24941);
and UO_922 (O_922,N_24711,N_24865);
and UO_923 (O_923,N_24725,N_24677);
xnor UO_924 (O_924,N_24953,N_24678);
nand UO_925 (O_925,N_24970,N_24514);
nor UO_926 (O_926,N_24590,N_24717);
or UO_927 (O_927,N_24912,N_24982);
xor UO_928 (O_928,N_24748,N_24666);
or UO_929 (O_929,N_24601,N_24542);
or UO_930 (O_930,N_24543,N_24507);
and UO_931 (O_931,N_24779,N_24764);
and UO_932 (O_932,N_24640,N_24847);
nor UO_933 (O_933,N_24781,N_24636);
or UO_934 (O_934,N_24663,N_24693);
or UO_935 (O_935,N_24827,N_24984);
or UO_936 (O_936,N_24981,N_24578);
nand UO_937 (O_937,N_24568,N_24821);
xnor UO_938 (O_938,N_24969,N_24961);
nand UO_939 (O_939,N_24997,N_24845);
and UO_940 (O_940,N_24968,N_24863);
or UO_941 (O_941,N_24563,N_24855);
or UO_942 (O_942,N_24600,N_24899);
or UO_943 (O_943,N_24626,N_24773);
or UO_944 (O_944,N_24725,N_24739);
or UO_945 (O_945,N_24697,N_24524);
nor UO_946 (O_946,N_24766,N_24858);
nor UO_947 (O_947,N_24637,N_24834);
nor UO_948 (O_948,N_24686,N_24705);
nor UO_949 (O_949,N_24775,N_24501);
or UO_950 (O_950,N_24800,N_24807);
nand UO_951 (O_951,N_24880,N_24645);
and UO_952 (O_952,N_24506,N_24870);
nor UO_953 (O_953,N_24814,N_24767);
nand UO_954 (O_954,N_24987,N_24604);
or UO_955 (O_955,N_24847,N_24796);
nor UO_956 (O_956,N_24862,N_24875);
and UO_957 (O_957,N_24631,N_24867);
and UO_958 (O_958,N_24524,N_24601);
and UO_959 (O_959,N_24659,N_24514);
or UO_960 (O_960,N_24503,N_24977);
or UO_961 (O_961,N_24504,N_24870);
nand UO_962 (O_962,N_24757,N_24997);
xor UO_963 (O_963,N_24525,N_24506);
nor UO_964 (O_964,N_24716,N_24656);
or UO_965 (O_965,N_24562,N_24638);
or UO_966 (O_966,N_24611,N_24545);
and UO_967 (O_967,N_24875,N_24547);
nor UO_968 (O_968,N_24552,N_24852);
or UO_969 (O_969,N_24950,N_24971);
and UO_970 (O_970,N_24673,N_24566);
nand UO_971 (O_971,N_24971,N_24676);
and UO_972 (O_972,N_24764,N_24730);
and UO_973 (O_973,N_24531,N_24718);
and UO_974 (O_974,N_24906,N_24661);
nand UO_975 (O_975,N_24528,N_24958);
xor UO_976 (O_976,N_24824,N_24800);
nand UO_977 (O_977,N_24815,N_24888);
nand UO_978 (O_978,N_24577,N_24861);
or UO_979 (O_979,N_24812,N_24943);
and UO_980 (O_980,N_24710,N_24842);
nand UO_981 (O_981,N_24829,N_24737);
nand UO_982 (O_982,N_24683,N_24715);
or UO_983 (O_983,N_24988,N_24714);
or UO_984 (O_984,N_24687,N_24528);
nor UO_985 (O_985,N_24798,N_24622);
nor UO_986 (O_986,N_24591,N_24872);
nand UO_987 (O_987,N_24536,N_24661);
or UO_988 (O_988,N_24734,N_24838);
nand UO_989 (O_989,N_24811,N_24587);
xnor UO_990 (O_990,N_24644,N_24503);
or UO_991 (O_991,N_24874,N_24969);
or UO_992 (O_992,N_24623,N_24806);
nor UO_993 (O_993,N_24699,N_24609);
and UO_994 (O_994,N_24809,N_24504);
and UO_995 (O_995,N_24570,N_24962);
and UO_996 (O_996,N_24728,N_24559);
nor UO_997 (O_997,N_24835,N_24694);
nor UO_998 (O_998,N_24565,N_24728);
and UO_999 (O_999,N_24738,N_24740);
nand UO_1000 (O_1000,N_24654,N_24840);
nor UO_1001 (O_1001,N_24671,N_24822);
nand UO_1002 (O_1002,N_24539,N_24636);
nand UO_1003 (O_1003,N_24522,N_24688);
nand UO_1004 (O_1004,N_24850,N_24602);
nand UO_1005 (O_1005,N_24801,N_24628);
and UO_1006 (O_1006,N_24663,N_24743);
nand UO_1007 (O_1007,N_24620,N_24799);
and UO_1008 (O_1008,N_24983,N_24554);
or UO_1009 (O_1009,N_24600,N_24874);
or UO_1010 (O_1010,N_24642,N_24686);
or UO_1011 (O_1011,N_24538,N_24579);
and UO_1012 (O_1012,N_24588,N_24612);
nor UO_1013 (O_1013,N_24998,N_24574);
nand UO_1014 (O_1014,N_24729,N_24819);
nand UO_1015 (O_1015,N_24704,N_24573);
nor UO_1016 (O_1016,N_24999,N_24664);
and UO_1017 (O_1017,N_24969,N_24686);
and UO_1018 (O_1018,N_24845,N_24573);
xor UO_1019 (O_1019,N_24522,N_24738);
or UO_1020 (O_1020,N_24967,N_24600);
or UO_1021 (O_1021,N_24564,N_24681);
nor UO_1022 (O_1022,N_24555,N_24751);
nand UO_1023 (O_1023,N_24543,N_24717);
nor UO_1024 (O_1024,N_24510,N_24502);
and UO_1025 (O_1025,N_24651,N_24660);
nand UO_1026 (O_1026,N_24726,N_24698);
and UO_1027 (O_1027,N_24717,N_24703);
or UO_1028 (O_1028,N_24874,N_24996);
or UO_1029 (O_1029,N_24639,N_24789);
nor UO_1030 (O_1030,N_24781,N_24782);
nor UO_1031 (O_1031,N_24862,N_24954);
nor UO_1032 (O_1032,N_24756,N_24718);
nand UO_1033 (O_1033,N_24709,N_24793);
and UO_1034 (O_1034,N_24746,N_24948);
or UO_1035 (O_1035,N_24744,N_24771);
nor UO_1036 (O_1036,N_24707,N_24685);
or UO_1037 (O_1037,N_24807,N_24529);
or UO_1038 (O_1038,N_24942,N_24503);
or UO_1039 (O_1039,N_24500,N_24704);
and UO_1040 (O_1040,N_24616,N_24777);
nand UO_1041 (O_1041,N_24939,N_24952);
or UO_1042 (O_1042,N_24676,N_24808);
and UO_1043 (O_1043,N_24633,N_24658);
xor UO_1044 (O_1044,N_24642,N_24921);
nand UO_1045 (O_1045,N_24732,N_24734);
nor UO_1046 (O_1046,N_24935,N_24806);
and UO_1047 (O_1047,N_24704,N_24582);
nand UO_1048 (O_1048,N_24982,N_24839);
or UO_1049 (O_1049,N_24922,N_24502);
and UO_1050 (O_1050,N_24645,N_24982);
nor UO_1051 (O_1051,N_24923,N_24781);
or UO_1052 (O_1052,N_24631,N_24727);
nand UO_1053 (O_1053,N_24544,N_24698);
or UO_1054 (O_1054,N_24888,N_24757);
or UO_1055 (O_1055,N_24886,N_24870);
xnor UO_1056 (O_1056,N_24706,N_24617);
or UO_1057 (O_1057,N_24771,N_24553);
nand UO_1058 (O_1058,N_24764,N_24747);
and UO_1059 (O_1059,N_24704,N_24753);
nor UO_1060 (O_1060,N_24524,N_24631);
nor UO_1061 (O_1061,N_24709,N_24810);
nor UO_1062 (O_1062,N_24580,N_24710);
nand UO_1063 (O_1063,N_24523,N_24911);
and UO_1064 (O_1064,N_24931,N_24844);
xor UO_1065 (O_1065,N_24962,N_24628);
nand UO_1066 (O_1066,N_24994,N_24945);
or UO_1067 (O_1067,N_24989,N_24812);
or UO_1068 (O_1068,N_24829,N_24984);
nand UO_1069 (O_1069,N_24920,N_24555);
nand UO_1070 (O_1070,N_24938,N_24880);
nand UO_1071 (O_1071,N_24859,N_24851);
nand UO_1072 (O_1072,N_24891,N_24861);
and UO_1073 (O_1073,N_24968,N_24906);
nor UO_1074 (O_1074,N_24681,N_24884);
or UO_1075 (O_1075,N_24836,N_24541);
nand UO_1076 (O_1076,N_24905,N_24524);
and UO_1077 (O_1077,N_24729,N_24695);
and UO_1078 (O_1078,N_24990,N_24942);
nand UO_1079 (O_1079,N_24630,N_24882);
and UO_1080 (O_1080,N_24782,N_24950);
nor UO_1081 (O_1081,N_24960,N_24568);
nand UO_1082 (O_1082,N_24880,N_24944);
nand UO_1083 (O_1083,N_24953,N_24945);
and UO_1084 (O_1084,N_24874,N_24628);
or UO_1085 (O_1085,N_24541,N_24626);
nor UO_1086 (O_1086,N_24727,N_24685);
nor UO_1087 (O_1087,N_24733,N_24793);
xor UO_1088 (O_1088,N_24553,N_24827);
nor UO_1089 (O_1089,N_24886,N_24696);
or UO_1090 (O_1090,N_24824,N_24566);
or UO_1091 (O_1091,N_24871,N_24688);
nand UO_1092 (O_1092,N_24665,N_24544);
nor UO_1093 (O_1093,N_24681,N_24998);
nand UO_1094 (O_1094,N_24551,N_24861);
nand UO_1095 (O_1095,N_24665,N_24911);
nor UO_1096 (O_1096,N_24769,N_24771);
or UO_1097 (O_1097,N_24817,N_24996);
or UO_1098 (O_1098,N_24904,N_24591);
xor UO_1099 (O_1099,N_24891,N_24863);
nand UO_1100 (O_1100,N_24715,N_24894);
nand UO_1101 (O_1101,N_24932,N_24906);
xnor UO_1102 (O_1102,N_24608,N_24599);
and UO_1103 (O_1103,N_24815,N_24788);
xnor UO_1104 (O_1104,N_24994,N_24794);
nand UO_1105 (O_1105,N_24742,N_24878);
nor UO_1106 (O_1106,N_24625,N_24900);
nand UO_1107 (O_1107,N_24728,N_24593);
and UO_1108 (O_1108,N_24940,N_24517);
or UO_1109 (O_1109,N_24695,N_24557);
or UO_1110 (O_1110,N_24652,N_24627);
nand UO_1111 (O_1111,N_24854,N_24984);
nand UO_1112 (O_1112,N_24546,N_24730);
and UO_1113 (O_1113,N_24632,N_24673);
or UO_1114 (O_1114,N_24674,N_24647);
and UO_1115 (O_1115,N_24958,N_24581);
or UO_1116 (O_1116,N_24559,N_24814);
nand UO_1117 (O_1117,N_24683,N_24639);
and UO_1118 (O_1118,N_24637,N_24708);
xnor UO_1119 (O_1119,N_24569,N_24611);
nor UO_1120 (O_1120,N_24730,N_24547);
nand UO_1121 (O_1121,N_24794,N_24840);
nor UO_1122 (O_1122,N_24629,N_24751);
and UO_1123 (O_1123,N_24801,N_24926);
and UO_1124 (O_1124,N_24785,N_24857);
nand UO_1125 (O_1125,N_24854,N_24996);
nor UO_1126 (O_1126,N_24643,N_24997);
xnor UO_1127 (O_1127,N_24840,N_24600);
nand UO_1128 (O_1128,N_24873,N_24869);
or UO_1129 (O_1129,N_24733,N_24837);
nand UO_1130 (O_1130,N_24984,N_24607);
xor UO_1131 (O_1131,N_24786,N_24580);
and UO_1132 (O_1132,N_24867,N_24737);
or UO_1133 (O_1133,N_24526,N_24671);
and UO_1134 (O_1134,N_24760,N_24983);
and UO_1135 (O_1135,N_24513,N_24553);
nand UO_1136 (O_1136,N_24504,N_24666);
and UO_1137 (O_1137,N_24775,N_24502);
nor UO_1138 (O_1138,N_24543,N_24830);
nor UO_1139 (O_1139,N_24927,N_24892);
and UO_1140 (O_1140,N_24998,N_24819);
and UO_1141 (O_1141,N_24862,N_24926);
nor UO_1142 (O_1142,N_24574,N_24802);
and UO_1143 (O_1143,N_24970,N_24801);
nor UO_1144 (O_1144,N_24735,N_24971);
nor UO_1145 (O_1145,N_24766,N_24970);
nor UO_1146 (O_1146,N_24502,N_24844);
nand UO_1147 (O_1147,N_24551,N_24651);
nand UO_1148 (O_1148,N_24855,N_24958);
nor UO_1149 (O_1149,N_24799,N_24908);
nand UO_1150 (O_1150,N_24800,N_24726);
nor UO_1151 (O_1151,N_24724,N_24930);
nor UO_1152 (O_1152,N_24956,N_24973);
or UO_1153 (O_1153,N_24526,N_24761);
or UO_1154 (O_1154,N_24505,N_24857);
nand UO_1155 (O_1155,N_24859,N_24879);
nor UO_1156 (O_1156,N_24672,N_24941);
and UO_1157 (O_1157,N_24630,N_24839);
and UO_1158 (O_1158,N_24562,N_24729);
or UO_1159 (O_1159,N_24722,N_24664);
xor UO_1160 (O_1160,N_24871,N_24543);
nand UO_1161 (O_1161,N_24752,N_24538);
nand UO_1162 (O_1162,N_24592,N_24543);
or UO_1163 (O_1163,N_24742,N_24611);
nand UO_1164 (O_1164,N_24574,N_24787);
and UO_1165 (O_1165,N_24515,N_24732);
nand UO_1166 (O_1166,N_24798,N_24634);
and UO_1167 (O_1167,N_24902,N_24871);
nand UO_1168 (O_1168,N_24952,N_24856);
and UO_1169 (O_1169,N_24788,N_24752);
nor UO_1170 (O_1170,N_24549,N_24716);
nor UO_1171 (O_1171,N_24650,N_24997);
nand UO_1172 (O_1172,N_24738,N_24920);
nor UO_1173 (O_1173,N_24933,N_24653);
and UO_1174 (O_1174,N_24996,N_24794);
and UO_1175 (O_1175,N_24796,N_24536);
or UO_1176 (O_1176,N_24904,N_24562);
nor UO_1177 (O_1177,N_24715,N_24646);
nand UO_1178 (O_1178,N_24981,N_24678);
xor UO_1179 (O_1179,N_24827,N_24671);
nand UO_1180 (O_1180,N_24519,N_24977);
nand UO_1181 (O_1181,N_24576,N_24539);
and UO_1182 (O_1182,N_24814,N_24992);
nor UO_1183 (O_1183,N_24528,N_24874);
or UO_1184 (O_1184,N_24822,N_24627);
nor UO_1185 (O_1185,N_24769,N_24702);
nor UO_1186 (O_1186,N_24816,N_24637);
nor UO_1187 (O_1187,N_24886,N_24944);
nor UO_1188 (O_1188,N_24941,N_24580);
or UO_1189 (O_1189,N_24868,N_24717);
nand UO_1190 (O_1190,N_24619,N_24849);
nand UO_1191 (O_1191,N_24879,N_24926);
and UO_1192 (O_1192,N_24795,N_24826);
or UO_1193 (O_1193,N_24768,N_24739);
xor UO_1194 (O_1194,N_24977,N_24560);
and UO_1195 (O_1195,N_24831,N_24566);
nor UO_1196 (O_1196,N_24780,N_24825);
and UO_1197 (O_1197,N_24653,N_24514);
nor UO_1198 (O_1198,N_24556,N_24800);
and UO_1199 (O_1199,N_24519,N_24872);
xnor UO_1200 (O_1200,N_24623,N_24880);
and UO_1201 (O_1201,N_24816,N_24983);
or UO_1202 (O_1202,N_24742,N_24827);
nor UO_1203 (O_1203,N_24545,N_24534);
nand UO_1204 (O_1204,N_24967,N_24937);
nor UO_1205 (O_1205,N_24593,N_24753);
and UO_1206 (O_1206,N_24878,N_24992);
nand UO_1207 (O_1207,N_24513,N_24788);
and UO_1208 (O_1208,N_24543,N_24893);
nor UO_1209 (O_1209,N_24627,N_24556);
and UO_1210 (O_1210,N_24602,N_24644);
or UO_1211 (O_1211,N_24563,N_24790);
or UO_1212 (O_1212,N_24517,N_24507);
and UO_1213 (O_1213,N_24569,N_24843);
or UO_1214 (O_1214,N_24643,N_24705);
nand UO_1215 (O_1215,N_24898,N_24584);
and UO_1216 (O_1216,N_24600,N_24979);
nor UO_1217 (O_1217,N_24958,N_24778);
or UO_1218 (O_1218,N_24687,N_24910);
and UO_1219 (O_1219,N_24583,N_24695);
or UO_1220 (O_1220,N_24944,N_24523);
nor UO_1221 (O_1221,N_24862,N_24594);
nor UO_1222 (O_1222,N_24576,N_24596);
or UO_1223 (O_1223,N_24852,N_24749);
nand UO_1224 (O_1224,N_24664,N_24827);
nor UO_1225 (O_1225,N_24641,N_24796);
or UO_1226 (O_1226,N_24989,N_24868);
or UO_1227 (O_1227,N_24854,N_24564);
and UO_1228 (O_1228,N_24855,N_24955);
or UO_1229 (O_1229,N_24759,N_24930);
and UO_1230 (O_1230,N_24979,N_24635);
nand UO_1231 (O_1231,N_24662,N_24746);
nand UO_1232 (O_1232,N_24639,N_24636);
or UO_1233 (O_1233,N_24837,N_24849);
xnor UO_1234 (O_1234,N_24858,N_24652);
and UO_1235 (O_1235,N_24600,N_24906);
or UO_1236 (O_1236,N_24917,N_24724);
nor UO_1237 (O_1237,N_24974,N_24780);
xnor UO_1238 (O_1238,N_24714,N_24643);
and UO_1239 (O_1239,N_24665,N_24595);
nand UO_1240 (O_1240,N_24983,N_24576);
and UO_1241 (O_1241,N_24916,N_24672);
or UO_1242 (O_1242,N_24806,N_24685);
or UO_1243 (O_1243,N_24539,N_24730);
and UO_1244 (O_1244,N_24781,N_24572);
and UO_1245 (O_1245,N_24980,N_24680);
nand UO_1246 (O_1246,N_24968,N_24866);
nand UO_1247 (O_1247,N_24801,N_24735);
and UO_1248 (O_1248,N_24842,N_24991);
nand UO_1249 (O_1249,N_24751,N_24745);
nand UO_1250 (O_1250,N_24657,N_24870);
and UO_1251 (O_1251,N_24809,N_24707);
nor UO_1252 (O_1252,N_24515,N_24767);
and UO_1253 (O_1253,N_24613,N_24610);
and UO_1254 (O_1254,N_24663,N_24803);
or UO_1255 (O_1255,N_24855,N_24678);
nand UO_1256 (O_1256,N_24799,N_24981);
nand UO_1257 (O_1257,N_24676,N_24540);
nor UO_1258 (O_1258,N_24828,N_24723);
nand UO_1259 (O_1259,N_24668,N_24528);
nand UO_1260 (O_1260,N_24684,N_24505);
or UO_1261 (O_1261,N_24687,N_24980);
nor UO_1262 (O_1262,N_24821,N_24965);
nor UO_1263 (O_1263,N_24733,N_24590);
and UO_1264 (O_1264,N_24569,N_24576);
and UO_1265 (O_1265,N_24675,N_24545);
and UO_1266 (O_1266,N_24712,N_24503);
and UO_1267 (O_1267,N_24723,N_24502);
and UO_1268 (O_1268,N_24521,N_24940);
nand UO_1269 (O_1269,N_24993,N_24680);
and UO_1270 (O_1270,N_24879,N_24740);
or UO_1271 (O_1271,N_24902,N_24936);
nand UO_1272 (O_1272,N_24519,N_24983);
xor UO_1273 (O_1273,N_24588,N_24611);
nor UO_1274 (O_1274,N_24720,N_24675);
and UO_1275 (O_1275,N_24999,N_24530);
xnor UO_1276 (O_1276,N_24630,N_24655);
nor UO_1277 (O_1277,N_24846,N_24838);
and UO_1278 (O_1278,N_24551,N_24665);
and UO_1279 (O_1279,N_24587,N_24772);
nor UO_1280 (O_1280,N_24839,N_24658);
or UO_1281 (O_1281,N_24569,N_24944);
nand UO_1282 (O_1282,N_24822,N_24989);
nand UO_1283 (O_1283,N_24734,N_24627);
xnor UO_1284 (O_1284,N_24855,N_24973);
and UO_1285 (O_1285,N_24748,N_24991);
or UO_1286 (O_1286,N_24939,N_24697);
or UO_1287 (O_1287,N_24502,N_24720);
nor UO_1288 (O_1288,N_24826,N_24635);
nand UO_1289 (O_1289,N_24512,N_24842);
nand UO_1290 (O_1290,N_24593,N_24598);
and UO_1291 (O_1291,N_24871,N_24816);
nor UO_1292 (O_1292,N_24738,N_24698);
and UO_1293 (O_1293,N_24733,N_24726);
or UO_1294 (O_1294,N_24545,N_24645);
nor UO_1295 (O_1295,N_24638,N_24582);
and UO_1296 (O_1296,N_24583,N_24588);
and UO_1297 (O_1297,N_24920,N_24501);
or UO_1298 (O_1298,N_24643,N_24899);
nand UO_1299 (O_1299,N_24788,N_24596);
and UO_1300 (O_1300,N_24957,N_24643);
nor UO_1301 (O_1301,N_24571,N_24615);
nand UO_1302 (O_1302,N_24718,N_24887);
or UO_1303 (O_1303,N_24539,N_24661);
nand UO_1304 (O_1304,N_24963,N_24627);
and UO_1305 (O_1305,N_24634,N_24877);
nand UO_1306 (O_1306,N_24771,N_24688);
and UO_1307 (O_1307,N_24874,N_24617);
nand UO_1308 (O_1308,N_24856,N_24902);
or UO_1309 (O_1309,N_24606,N_24514);
nor UO_1310 (O_1310,N_24601,N_24606);
nor UO_1311 (O_1311,N_24910,N_24750);
nor UO_1312 (O_1312,N_24895,N_24790);
nand UO_1313 (O_1313,N_24939,N_24890);
and UO_1314 (O_1314,N_24602,N_24978);
nand UO_1315 (O_1315,N_24961,N_24705);
nor UO_1316 (O_1316,N_24604,N_24549);
nand UO_1317 (O_1317,N_24531,N_24621);
nand UO_1318 (O_1318,N_24612,N_24712);
or UO_1319 (O_1319,N_24760,N_24771);
nand UO_1320 (O_1320,N_24724,N_24927);
or UO_1321 (O_1321,N_24653,N_24655);
nand UO_1322 (O_1322,N_24873,N_24543);
nand UO_1323 (O_1323,N_24584,N_24891);
and UO_1324 (O_1324,N_24756,N_24743);
nand UO_1325 (O_1325,N_24666,N_24849);
and UO_1326 (O_1326,N_24651,N_24549);
or UO_1327 (O_1327,N_24971,N_24594);
nor UO_1328 (O_1328,N_24854,N_24517);
nor UO_1329 (O_1329,N_24935,N_24728);
or UO_1330 (O_1330,N_24943,N_24708);
nand UO_1331 (O_1331,N_24695,N_24837);
and UO_1332 (O_1332,N_24700,N_24758);
and UO_1333 (O_1333,N_24764,N_24979);
and UO_1334 (O_1334,N_24839,N_24753);
and UO_1335 (O_1335,N_24836,N_24687);
nor UO_1336 (O_1336,N_24599,N_24947);
nand UO_1337 (O_1337,N_24887,N_24857);
and UO_1338 (O_1338,N_24608,N_24853);
or UO_1339 (O_1339,N_24634,N_24873);
or UO_1340 (O_1340,N_24858,N_24566);
xor UO_1341 (O_1341,N_24800,N_24675);
nand UO_1342 (O_1342,N_24860,N_24911);
and UO_1343 (O_1343,N_24759,N_24705);
or UO_1344 (O_1344,N_24809,N_24805);
or UO_1345 (O_1345,N_24987,N_24852);
and UO_1346 (O_1346,N_24516,N_24907);
or UO_1347 (O_1347,N_24801,N_24903);
xnor UO_1348 (O_1348,N_24638,N_24664);
or UO_1349 (O_1349,N_24609,N_24735);
xnor UO_1350 (O_1350,N_24887,N_24589);
nor UO_1351 (O_1351,N_24795,N_24546);
or UO_1352 (O_1352,N_24518,N_24788);
or UO_1353 (O_1353,N_24680,N_24867);
nand UO_1354 (O_1354,N_24545,N_24718);
and UO_1355 (O_1355,N_24903,N_24838);
or UO_1356 (O_1356,N_24734,N_24910);
and UO_1357 (O_1357,N_24922,N_24834);
xor UO_1358 (O_1358,N_24844,N_24659);
nor UO_1359 (O_1359,N_24967,N_24871);
and UO_1360 (O_1360,N_24915,N_24864);
and UO_1361 (O_1361,N_24525,N_24904);
and UO_1362 (O_1362,N_24821,N_24833);
xnor UO_1363 (O_1363,N_24918,N_24860);
nand UO_1364 (O_1364,N_24724,N_24900);
nor UO_1365 (O_1365,N_24562,N_24754);
nand UO_1366 (O_1366,N_24858,N_24697);
nor UO_1367 (O_1367,N_24560,N_24733);
or UO_1368 (O_1368,N_24704,N_24799);
and UO_1369 (O_1369,N_24590,N_24519);
xor UO_1370 (O_1370,N_24560,N_24558);
nand UO_1371 (O_1371,N_24717,N_24763);
nor UO_1372 (O_1372,N_24642,N_24627);
nand UO_1373 (O_1373,N_24804,N_24611);
and UO_1374 (O_1374,N_24956,N_24790);
nand UO_1375 (O_1375,N_24788,N_24609);
or UO_1376 (O_1376,N_24706,N_24841);
or UO_1377 (O_1377,N_24837,N_24814);
nor UO_1378 (O_1378,N_24928,N_24769);
or UO_1379 (O_1379,N_24574,N_24701);
nor UO_1380 (O_1380,N_24507,N_24780);
nor UO_1381 (O_1381,N_24700,N_24511);
xnor UO_1382 (O_1382,N_24684,N_24706);
nand UO_1383 (O_1383,N_24887,N_24874);
nor UO_1384 (O_1384,N_24713,N_24569);
nor UO_1385 (O_1385,N_24823,N_24798);
or UO_1386 (O_1386,N_24693,N_24513);
nand UO_1387 (O_1387,N_24617,N_24714);
xnor UO_1388 (O_1388,N_24900,N_24989);
nand UO_1389 (O_1389,N_24769,N_24633);
and UO_1390 (O_1390,N_24762,N_24743);
and UO_1391 (O_1391,N_24538,N_24689);
nor UO_1392 (O_1392,N_24635,N_24797);
nand UO_1393 (O_1393,N_24562,N_24580);
or UO_1394 (O_1394,N_24605,N_24734);
and UO_1395 (O_1395,N_24524,N_24911);
nand UO_1396 (O_1396,N_24687,N_24709);
nor UO_1397 (O_1397,N_24788,N_24696);
or UO_1398 (O_1398,N_24768,N_24716);
nor UO_1399 (O_1399,N_24996,N_24738);
and UO_1400 (O_1400,N_24610,N_24820);
and UO_1401 (O_1401,N_24610,N_24578);
and UO_1402 (O_1402,N_24721,N_24607);
xor UO_1403 (O_1403,N_24820,N_24924);
nor UO_1404 (O_1404,N_24922,N_24630);
xnor UO_1405 (O_1405,N_24609,N_24864);
nand UO_1406 (O_1406,N_24936,N_24572);
nor UO_1407 (O_1407,N_24973,N_24763);
or UO_1408 (O_1408,N_24747,N_24526);
or UO_1409 (O_1409,N_24838,N_24764);
nor UO_1410 (O_1410,N_24871,N_24607);
and UO_1411 (O_1411,N_24837,N_24694);
nor UO_1412 (O_1412,N_24933,N_24753);
nand UO_1413 (O_1413,N_24816,N_24591);
or UO_1414 (O_1414,N_24956,N_24511);
or UO_1415 (O_1415,N_24975,N_24581);
nand UO_1416 (O_1416,N_24860,N_24523);
and UO_1417 (O_1417,N_24827,N_24599);
or UO_1418 (O_1418,N_24827,N_24524);
nand UO_1419 (O_1419,N_24505,N_24646);
nor UO_1420 (O_1420,N_24517,N_24936);
or UO_1421 (O_1421,N_24648,N_24603);
and UO_1422 (O_1422,N_24818,N_24990);
xnor UO_1423 (O_1423,N_24884,N_24928);
nor UO_1424 (O_1424,N_24969,N_24826);
or UO_1425 (O_1425,N_24622,N_24617);
or UO_1426 (O_1426,N_24913,N_24643);
xor UO_1427 (O_1427,N_24811,N_24594);
and UO_1428 (O_1428,N_24893,N_24989);
and UO_1429 (O_1429,N_24659,N_24894);
nand UO_1430 (O_1430,N_24778,N_24956);
nand UO_1431 (O_1431,N_24901,N_24947);
nor UO_1432 (O_1432,N_24592,N_24950);
or UO_1433 (O_1433,N_24793,N_24672);
or UO_1434 (O_1434,N_24883,N_24751);
and UO_1435 (O_1435,N_24890,N_24707);
nor UO_1436 (O_1436,N_24934,N_24928);
and UO_1437 (O_1437,N_24522,N_24767);
and UO_1438 (O_1438,N_24536,N_24560);
and UO_1439 (O_1439,N_24921,N_24513);
or UO_1440 (O_1440,N_24920,N_24603);
nor UO_1441 (O_1441,N_24561,N_24902);
nor UO_1442 (O_1442,N_24564,N_24954);
and UO_1443 (O_1443,N_24683,N_24984);
or UO_1444 (O_1444,N_24934,N_24697);
and UO_1445 (O_1445,N_24909,N_24599);
nor UO_1446 (O_1446,N_24718,N_24648);
or UO_1447 (O_1447,N_24701,N_24521);
or UO_1448 (O_1448,N_24998,N_24782);
nand UO_1449 (O_1449,N_24748,N_24526);
and UO_1450 (O_1450,N_24729,N_24593);
nand UO_1451 (O_1451,N_24764,N_24880);
or UO_1452 (O_1452,N_24654,N_24540);
nor UO_1453 (O_1453,N_24983,N_24676);
and UO_1454 (O_1454,N_24901,N_24705);
or UO_1455 (O_1455,N_24566,N_24926);
nor UO_1456 (O_1456,N_24658,N_24728);
or UO_1457 (O_1457,N_24865,N_24827);
nor UO_1458 (O_1458,N_24819,N_24612);
nand UO_1459 (O_1459,N_24514,N_24518);
xnor UO_1460 (O_1460,N_24843,N_24960);
nor UO_1461 (O_1461,N_24556,N_24922);
and UO_1462 (O_1462,N_24652,N_24925);
nor UO_1463 (O_1463,N_24888,N_24578);
and UO_1464 (O_1464,N_24504,N_24619);
nor UO_1465 (O_1465,N_24976,N_24805);
nor UO_1466 (O_1466,N_24795,N_24991);
xor UO_1467 (O_1467,N_24656,N_24594);
or UO_1468 (O_1468,N_24968,N_24611);
or UO_1469 (O_1469,N_24861,N_24832);
nand UO_1470 (O_1470,N_24858,N_24556);
or UO_1471 (O_1471,N_24539,N_24944);
nor UO_1472 (O_1472,N_24554,N_24939);
nand UO_1473 (O_1473,N_24981,N_24681);
nand UO_1474 (O_1474,N_24941,N_24981);
xnor UO_1475 (O_1475,N_24901,N_24940);
nand UO_1476 (O_1476,N_24834,N_24852);
or UO_1477 (O_1477,N_24681,N_24746);
nand UO_1478 (O_1478,N_24594,N_24738);
and UO_1479 (O_1479,N_24567,N_24842);
and UO_1480 (O_1480,N_24509,N_24909);
or UO_1481 (O_1481,N_24674,N_24567);
or UO_1482 (O_1482,N_24600,N_24762);
nand UO_1483 (O_1483,N_24999,N_24759);
or UO_1484 (O_1484,N_24624,N_24830);
nor UO_1485 (O_1485,N_24804,N_24980);
nand UO_1486 (O_1486,N_24846,N_24983);
or UO_1487 (O_1487,N_24698,N_24801);
and UO_1488 (O_1488,N_24914,N_24682);
nand UO_1489 (O_1489,N_24537,N_24916);
xnor UO_1490 (O_1490,N_24599,N_24795);
or UO_1491 (O_1491,N_24729,N_24766);
or UO_1492 (O_1492,N_24581,N_24594);
nor UO_1493 (O_1493,N_24841,N_24823);
nor UO_1494 (O_1494,N_24741,N_24757);
nand UO_1495 (O_1495,N_24610,N_24812);
nor UO_1496 (O_1496,N_24779,N_24902);
xor UO_1497 (O_1497,N_24822,N_24751);
or UO_1498 (O_1498,N_24798,N_24940);
nand UO_1499 (O_1499,N_24592,N_24877);
nor UO_1500 (O_1500,N_24986,N_24901);
nand UO_1501 (O_1501,N_24612,N_24621);
or UO_1502 (O_1502,N_24908,N_24534);
and UO_1503 (O_1503,N_24612,N_24965);
nor UO_1504 (O_1504,N_24621,N_24666);
nand UO_1505 (O_1505,N_24922,N_24842);
or UO_1506 (O_1506,N_24622,N_24506);
and UO_1507 (O_1507,N_24614,N_24975);
nand UO_1508 (O_1508,N_24908,N_24932);
nor UO_1509 (O_1509,N_24595,N_24782);
and UO_1510 (O_1510,N_24766,N_24602);
and UO_1511 (O_1511,N_24701,N_24736);
and UO_1512 (O_1512,N_24658,N_24503);
or UO_1513 (O_1513,N_24710,N_24782);
nor UO_1514 (O_1514,N_24746,N_24963);
and UO_1515 (O_1515,N_24711,N_24727);
nor UO_1516 (O_1516,N_24508,N_24862);
xor UO_1517 (O_1517,N_24561,N_24522);
nand UO_1518 (O_1518,N_24925,N_24714);
nor UO_1519 (O_1519,N_24689,N_24595);
xor UO_1520 (O_1520,N_24505,N_24730);
nand UO_1521 (O_1521,N_24545,N_24529);
nand UO_1522 (O_1522,N_24575,N_24679);
nand UO_1523 (O_1523,N_24764,N_24983);
and UO_1524 (O_1524,N_24931,N_24744);
and UO_1525 (O_1525,N_24532,N_24520);
xor UO_1526 (O_1526,N_24699,N_24957);
nor UO_1527 (O_1527,N_24587,N_24617);
nand UO_1528 (O_1528,N_24690,N_24938);
and UO_1529 (O_1529,N_24984,N_24702);
xnor UO_1530 (O_1530,N_24830,N_24812);
nand UO_1531 (O_1531,N_24744,N_24738);
xnor UO_1532 (O_1532,N_24869,N_24576);
nor UO_1533 (O_1533,N_24845,N_24605);
xnor UO_1534 (O_1534,N_24827,N_24676);
xor UO_1535 (O_1535,N_24530,N_24980);
nor UO_1536 (O_1536,N_24674,N_24683);
nand UO_1537 (O_1537,N_24664,N_24816);
or UO_1538 (O_1538,N_24918,N_24811);
nor UO_1539 (O_1539,N_24843,N_24754);
nand UO_1540 (O_1540,N_24679,N_24890);
and UO_1541 (O_1541,N_24743,N_24677);
and UO_1542 (O_1542,N_24573,N_24890);
and UO_1543 (O_1543,N_24851,N_24703);
nor UO_1544 (O_1544,N_24684,N_24753);
nand UO_1545 (O_1545,N_24811,N_24984);
xor UO_1546 (O_1546,N_24671,N_24909);
xor UO_1547 (O_1547,N_24561,N_24999);
nor UO_1548 (O_1548,N_24698,N_24849);
nor UO_1549 (O_1549,N_24659,N_24573);
nand UO_1550 (O_1550,N_24616,N_24508);
nor UO_1551 (O_1551,N_24501,N_24642);
and UO_1552 (O_1552,N_24525,N_24958);
nor UO_1553 (O_1553,N_24949,N_24526);
and UO_1554 (O_1554,N_24539,N_24927);
and UO_1555 (O_1555,N_24509,N_24523);
and UO_1556 (O_1556,N_24864,N_24789);
and UO_1557 (O_1557,N_24704,N_24936);
nor UO_1558 (O_1558,N_24960,N_24513);
nand UO_1559 (O_1559,N_24944,N_24777);
nand UO_1560 (O_1560,N_24958,N_24832);
nor UO_1561 (O_1561,N_24921,N_24799);
or UO_1562 (O_1562,N_24922,N_24876);
nor UO_1563 (O_1563,N_24704,N_24986);
nor UO_1564 (O_1564,N_24998,N_24634);
xnor UO_1565 (O_1565,N_24911,N_24896);
nor UO_1566 (O_1566,N_24546,N_24631);
nand UO_1567 (O_1567,N_24820,N_24537);
or UO_1568 (O_1568,N_24720,N_24912);
nor UO_1569 (O_1569,N_24919,N_24535);
nor UO_1570 (O_1570,N_24501,N_24667);
or UO_1571 (O_1571,N_24970,N_24817);
nand UO_1572 (O_1572,N_24768,N_24525);
nand UO_1573 (O_1573,N_24670,N_24776);
and UO_1574 (O_1574,N_24872,N_24853);
and UO_1575 (O_1575,N_24574,N_24822);
or UO_1576 (O_1576,N_24797,N_24962);
or UO_1577 (O_1577,N_24919,N_24773);
or UO_1578 (O_1578,N_24537,N_24539);
nor UO_1579 (O_1579,N_24674,N_24976);
nand UO_1580 (O_1580,N_24601,N_24972);
or UO_1581 (O_1581,N_24736,N_24765);
nand UO_1582 (O_1582,N_24522,N_24824);
or UO_1583 (O_1583,N_24708,N_24989);
nor UO_1584 (O_1584,N_24812,N_24751);
and UO_1585 (O_1585,N_24779,N_24885);
nor UO_1586 (O_1586,N_24830,N_24571);
or UO_1587 (O_1587,N_24667,N_24560);
xnor UO_1588 (O_1588,N_24650,N_24967);
nor UO_1589 (O_1589,N_24947,N_24887);
or UO_1590 (O_1590,N_24930,N_24860);
nor UO_1591 (O_1591,N_24963,N_24669);
xnor UO_1592 (O_1592,N_24785,N_24925);
and UO_1593 (O_1593,N_24580,N_24700);
nor UO_1594 (O_1594,N_24557,N_24830);
and UO_1595 (O_1595,N_24716,N_24556);
or UO_1596 (O_1596,N_24960,N_24899);
nor UO_1597 (O_1597,N_24705,N_24942);
nand UO_1598 (O_1598,N_24661,N_24740);
or UO_1599 (O_1599,N_24865,N_24713);
nor UO_1600 (O_1600,N_24916,N_24527);
and UO_1601 (O_1601,N_24670,N_24945);
nor UO_1602 (O_1602,N_24532,N_24514);
and UO_1603 (O_1603,N_24944,N_24503);
nand UO_1604 (O_1604,N_24538,N_24738);
nor UO_1605 (O_1605,N_24595,N_24721);
nor UO_1606 (O_1606,N_24996,N_24972);
or UO_1607 (O_1607,N_24708,N_24741);
or UO_1608 (O_1608,N_24510,N_24726);
nand UO_1609 (O_1609,N_24962,N_24639);
and UO_1610 (O_1610,N_24794,N_24713);
nand UO_1611 (O_1611,N_24842,N_24548);
or UO_1612 (O_1612,N_24824,N_24720);
nor UO_1613 (O_1613,N_24612,N_24859);
nand UO_1614 (O_1614,N_24965,N_24753);
or UO_1615 (O_1615,N_24702,N_24833);
xor UO_1616 (O_1616,N_24619,N_24533);
or UO_1617 (O_1617,N_24856,N_24555);
xnor UO_1618 (O_1618,N_24876,N_24963);
and UO_1619 (O_1619,N_24971,N_24805);
and UO_1620 (O_1620,N_24844,N_24770);
and UO_1621 (O_1621,N_24975,N_24895);
nand UO_1622 (O_1622,N_24661,N_24897);
nor UO_1623 (O_1623,N_24574,N_24780);
or UO_1624 (O_1624,N_24754,N_24761);
nor UO_1625 (O_1625,N_24952,N_24760);
or UO_1626 (O_1626,N_24807,N_24770);
nand UO_1627 (O_1627,N_24635,N_24873);
xor UO_1628 (O_1628,N_24696,N_24878);
xnor UO_1629 (O_1629,N_24874,N_24883);
nand UO_1630 (O_1630,N_24686,N_24594);
nand UO_1631 (O_1631,N_24955,N_24970);
and UO_1632 (O_1632,N_24728,N_24980);
or UO_1633 (O_1633,N_24844,N_24604);
or UO_1634 (O_1634,N_24759,N_24567);
and UO_1635 (O_1635,N_24629,N_24571);
nor UO_1636 (O_1636,N_24557,N_24712);
or UO_1637 (O_1637,N_24537,N_24789);
or UO_1638 (O_1638,N_24811,N_24849);
nor UO_1639 (O_1639,N_24881,N_24909);
and UO_1640 (O_1640,N_24732,N_24871);
or UO_1641 (O_1641,N_24676,N_24715);
and UO_1642 (O_1642,N_24714,N_24833);
xnor UO_1643 (O_1643,N_24672,N_24837);
or UO_1644 (O_1644,N_24627,N_24745);
nand UO_1645 (O_1645,N_24564,N_24814);
xnor UO_1646 (O_1646,N_24677,N_24797);
and UO_1647 (O_1647,N_24997,N_24641);
nor UO_1648 (O_1648,N_24805,N_24965);
or UO_1649 (O_1649,N_24553,N_24772);
nand UO_1650 (O_1650,N_24591,N_24636);
and UO_1651 (O_1651,N_24628,N_24778);
nor UO_1652 (O_1652,N_24996,N_24902);
xnor UO_1653 (O_1653,N_24603,N_24726);
nand UO_1654 (O_1654,N_24537,N_24669);
nand UO_1655 (O_1655,N_24737,N_24931);
xor UO_1656 (O_1656,N_24748,N_24613);
nand UO_1657 (O_1657,N_24765,N_24881);
nand UO_1658 (O_1658,N_24989,N_24650);
nand UO_1659 (O_1659,N_24630,N_24991);
nand UO_1660 (O_1660,N_24550,N_24990);
or UO_1661 (O_1661,N_24596,N_24841);
nor UO_1662 (O_1662,N_24955,N_24657);
xor UO_1663 (O_1663,N_24504,N_24762);
nor UO_1664 (O_1664,N_24773,N_24937);
xnor UO_1665 (O_1665,N_24801,N_24871);
nand UO_1666 (O_1666,N_24958,N_24621);
and UO_1667 (O_1667,N_24644,N_24626);
or UO_1668 (O_1668,N_24962,N_24551);
nor UO_1669 (O_1669,N_24896,N_24514);
nand UO_1670 (O_1670,N_24595,N_24693);
nand UO_1671 (O_1671,N_24853,N_24620);
nor UO_1672 (O_1672,N_24722,N_24846);
nor UO_1673 (O_1673,N_24683,N_24500);
nor UO_1674 (O_1674,N_24530,N_24933);
and UO_1675 (O_1675,N_24922,N_24809);
and UO_1676 (O_1676,N_24904,N_24636);
xnor UO_1677 (O_1677,N_24639,N_24591);
or UO_1678 (O_1678,N_24738,N_24830);
nor UO_1679 (O_1679,N_24854,N_24867);
and UO_1680 (O_1680,N_24740,N_24666);
nor UO_1681 (O_1681,N_24811,N_24905);
nor UO_1682 (O_1682,N_24827,N_24957);
xor UO_1683 (O_1683,N_24584,N_24590);
and UO_1684 (O_1684,N_24565,N_24556);
or UO_1685 (O_1685,N_24513,N_24913);
and UO_1686 (O_1686,N_24785,N_24863);
nor UO_1687 (O_1687,N_24582,N_24593);
or UO_1688 (O_1688,N_24534,N_24576);
or UO_1689 (O_1689,N_24897,N_24910);
and UO_1690 (O_1690,N_24510,N_24500);
nor UO_1691 (O_1691,N_24844,N_24569);
or UO_1692 (O_1692,N_24938,N_24680);
and UO_1693 (O_1693,N_24575,N_24510);
nand UO_1694 (O_1694,N_24601,N_24540);
and UO_1695 (O_1695,N_24527,N_24795);
or UO_1696 (O_1696,N_24975,N_24843);
nand UO_1697 (O_1697,N_24831,N_24529);
nor UO_1698 (O_1698,N_24970,N_24685);
or UO_1699 (O_1699,N_24884,N_24937);
or UO_1700 (O_1700,N_24566,N_24719);
and UO_1701 (O_1701,N_24889,N_24768);
or UO_1702 (O_1702,N_24651,N_24768);
or UO_1703 (O_1703,N_24857,N_24662);
and UO_1704 (O_1704,N_24977,N_24716);
or UO_1705 (O_1705,N_24746,N_24682);
nand UO_1706 (O_1706,N_24880,N_24630);
or UO_1707 (O_1707,N_24674,N_24924);
xnor UO_1708 (O_1708,N_24647,N_24617);
and UO_1709 (O_1709,N_24843,N_24528);
xor UO_1710 (O_1710,N_24787,N_24691);
and UO_1711 (O_1711,N_24550,N_24800);
xor UO_1712 (O_1712,N_24730,N_24914);
xnor UO_1713 (O_1713,N_24725,N_24647);
nor UO_1714 (O_1714,N_24654,N_24512);
xnor UO_1715 (O_1715,N_24520,N_24853);
or UO_1716 (O_1716,N_24606,N_24928);
nand UO_1717 (O_1717,N_24970,N_24643);
nand UO_1718 (O_1718,N_24870,N_24996);
and UO_1719 (O_1719,N_24881,N_24651);
or UO_1720 (O_1720,N_24690,N_24619);
and UO_1721 (O_1721,N_24575,N_24843);
xnor UO_1722 (O_1722,N_24633,N_24909);
or UO_1723 (O_1723,N_24576,N_24963);
and UO_1724 (O_1724,N_24599,N_24830);
or UO_1725 (O_1725,N_24949,N_24981);
nand UO_1726 (O_1726,N_24673,N_24644);
or UO_1727 (O_1727,N_24545,N_24860);
xor UO_1728 (O_1728,N_24527,N_24736);
nand UO_1729 (O_1729,N_24827,N_24996);
xor UO_1730 (O_1730,N_24935,N_24615);
xor UO_1731 (O_1731,N_24670,N_24785);
and UO_1732 (O_1732,N_24620,N_24773);
and UO_1733 (O_1733,N_24642,N_24887);
nor UO_1734 (O_1734,N_24643,N_24771);
and UO_1735 (O_1735,N_24738,N_24548);
nand UO_1736 (O_1736,N_24840,N_24875);
nor UO_1737 (O_1737,N_24593,N_24898);
nand UO_1738 (O_1738,N_24989,N_24535);
nand UO_1739 (O_1739,N_24717,N_24713);
nand UO_1740 (O_1740,N_24906,N_24908);
xnor UO_1741 (O_1741,N_24914,N_24712);
nor UO_1742 (O_1742,N_24579,N_24747);
and UO_1743 (O_1743,N_24775,N_24828);
nor UO_1744 (O_1744,N_24620,N_24896);
or UO_1745 (O_1745,N_24711,N_24968);
or UO_1746 (O_1746,N_24750,N_24927);
xnor UO_1747 (O_1747,N_24942,N_24543);
or UO_1748 (O_1748,N_24725,N_24532);
or UO_1749 (O_1749,N_24690,N_24552);
nor UO_1750 (O_1750,N_24900,N_24921);
nand UO_1751 (O_1751,N_24783,N_24992);
nand UO_1752 (O_1752,N_24855,N_24795);
nand UO_1753 (O_1753,N_24867,N_24804);
or UO_1754 (O_1754,N_24998,N_24988);
nand UO_1755 (O_1755,N_24796,N_24680);
nor UO_1756 (O_1756,N_24874,N_24602);
or UO_1757 (O_1757,N_24849,N_24595);
xnor UO_1758 (O_1758,N_24838,N_24767);
nand UO_1759 (O_1759,N_24817,N_24840);
or UO_1760 (O_1760,N_24855,N_24938);
nand UO_1761 (O_1761,N_24529,N_24942);
xnor UO_1762 (O_1762,N_24881,N_24864);
or UO_1763 (O_1763,N_24997,N_24680);
or UO_1764 (O_1764,N_24778,N_24983);
xor UO_1765 (O_1765,N_24880,N_24569);
and UO_1766 (O_1766,N_24840,N_24742);
nor UO_1767 (O_1767,N_24527,N_24761);
and UO_1768 (O_1768,N_24740,N_24712);
nand UO_1769 (O_1769,N_24614,N_24754);
or UO_1770 (O_1770,N_24760,N_24586);
and UO_1771 (O_1771,N_24810,N_24602);
nor UO_1772 (O_1772,N_24536,N_24941);
nand UO_1773 (O_1773,N_24663,N_24882);
or UO_1774 (O_1774,N_24619,N_24747);
nor UO_1775 (O_1775,N_24990,N_24505);
or UO_1776 (O_1776,N_24949,N_24666);
nand UO_1777 (O_1777,N_24942,N_24786);
and UO_1778 (O_1778,N_24824,N_24541);
and UO_1779 (O_1779,N_24706,N_24588);
or UO_1780 (O_1780,N_24949,N_24898);
and UO_1781 (O_1781,N_24707,N_24941);
nand UO_1782 (O_1782,N_24734,N_24982);
nor UO_1783 (O_1783,N_24771,N_24560);
and UO_1784 (O_1784,N_24985,N_24570);
nand UO_1785 (O_1785,N_24999,N_24514);
nor UO_1786 (O_1786,N_24589,N_24642);
and UO_1787 (O_1787,N_24794,N_24929);
xnor UO_1788 (O_1788,N_24803,N_24615);
nor UO_1789 (O_1789,N_24781,N_24831);
and UO_1790 (O_1790,N_24870,N_24640);
or UO_1791 (O_1791,N_24686,N_24513);
nor UO_1792 (O_1792,N_24995,N_24578);
nand UO_1793 (O_1793,N_24744,N_24850);
nand UO_1794 (O_1794,N_24912,N_24540);
xor UO_1795 (O_1795,N_24820,N_24502);
nor UO_1796 (O_1796,N_24923,N_24800);
and UO_1797 (O_1797,N_24673,N_24548);
nor UO_1798 (O_1798,N_24674,N_24575);
nor UO_1799 (O_1799,N_24849,N_24681);
nor UO_1800 (O_1800,N_24733,N_24904);
and UO_1801 (O_1801,N_24990,N_24622);
nor UO_1802 (O_1802,N_24724,N_24539);
or UO_1803 (O_1803,N_24579,N_24850);
and UO_1804 (O_1804,N_24905,N_24932);
and UO_1805 (O_1805,N_24597,N_24584);
nor UO_1806 (O_1806,N_24841,N_24555);
nand UO_1807 (O_1807,N_24586,N_24917);
or UO_1808 (O_1808,N_24764,N_24519);
nor UO_1809 (O_1809,N_24643,N_24818);
nor UO_1810 (O_1810,N_24744,N_24767);
xnor UO_1811 (O_1811,N_24734,N_24864);
nand UO_1812 (O_1812,N_24564,N_24723);
or UO_1813 (O_1813,N_24966,N_24635);
xor UO_1814 (O_1814,N_24655,N_24698);
nand UO_1815 (O_1815,N_24729,N_24767);
nand UO_1816 (O_1816,N_24562,N_24519);
and UO_1817 (O_1817,N_24976,N_24931);
and UO_1818 (O_1818,N_24769,N_24692);
nor UO_1819 (O_1819,N_24729,N_24613);
nor UO_1820 (O_1820,N_24674,N_24862);
nor UO_1821 (O_1821,N_24856,N_24675);
nor UO_1822 (O_1822,N_24958,N_24865);
nor UO_1823 (O_1823,N_24817,N_24626);
or UO_1824 (O_1824,N_24547,N_24772);
nor UO_1825 (O_1825,N_24870,N_24585);
nand UO_1826 (O_1826,N_24805,N_24635);
xor UO_1827 (O_1827,N_24560,N_24757);
and UO_1828 (O_1828,N_24556,N_24975);
or UO_1829 (O_1829,N_24523,N_24867);
and UO_1830 (O_1830,N_24993,N_24610);
nand UO_1831 (O_1831,N_24856,N_24648);
nand UO_1832 (O_1832,N_24921,N_24886);
and UO_1833 (O_1833,N_24506,N_24572);
nor UO_1834 (O_1834,N_24679,N_24792);
or UO_1835 (O_1835,N_24687,N_24685);
and UO_1836 (O_1836,N_24979,N_24881);
and UO_1837 (O_1837,N_24809,N_24622);
nand UO_1838 (O_1838,N_24520,N_24885);
nand UO_1839 (O_1839,N_24753,N_24500);
nand UO_1840 (O_1840,N_24701,N_24858);
nor UO_1841 (O_1841,N_24733,N_24626);
xor UO_1842 (O_1842,N_24738,N_24563);
nand UO_1843 (O_1843,N_24574,N_24519);
or UO_1844 (O_1844,N_24900,N_24877);
nor UO_1845 (O_1845,N_24556,N_24903);
nand UO_1846 (O_1846,N_24854,N_24663);
nor UO_1847 (O_1847,N_24966,N_24848);
or UO_1848 (O_1848,N_24567,N_24829);
or UO_1849 (O_1849,N_24689,N_24728);
nor UO_1850 (O_1850,N_24561,N_24572);
and UO_1851 (O_1851,N_24853,N_24785);
and UO_1852 (O_1852,N_24835,N_24760);
or UO_1853 (O_1853,N_24630,N_24724);
nand UO_1854 (O_1854,N_24995,N_24563);
nor UO_1855 (O_1855,N_24635,N_24773);
xnor UO_1856 (O_1856,N_24877,N_24503);
nand UO_1857 (O_1857,N_24551,N_24883);
nor UO_1858 (O_1858,N_24695,N_24522);
xnor UO_1859 (O_1859,N_24986,N_24957);
and UO_1860 (O_1860,N_24543,N_24553);
nand UO_1861 (O_1861,N_24812,N_24886);
and UO_1862 (O_1862,N_24947,N_24799);
or UO_1863 (O_1863,N_24787,N_24944);
nand UO_1864 (O_1864,N_24543,N_24546);
and UO_1865 (O_1865,N_24721,N_24572);
nand UO_1866 (O_1866,N_24872,N_24995);
nor UO_1867 (O_1867,N_24607,N_24532);
nand UO_1868 (O_1868,N_24586,N_24909);
nand UO_1869 (O_1869,N_24584,N_24925);
and UO_1870 (O_1870,N_24801,N_24722);
nand UO_1871 (O_1871,N_24603,N_24908);
nor UO_1872 (O_1872,N_24615,N_24992);
or UO_1873 (O_1873,N_24685,N_24635);
and UO_1874 (O_1874,N_24697,N_24891);
and UO_1875 (O_1875,N_24560,N_24632);
and UO_1876 (O_1876,N_24521,N_24564);
nor UO_1877 (O_1877,N_24563,N_24523);
nor UO_1878 (O_1878,N_24914,N_24903);
and UO_1879 (O_1879,N_24653,N_24609);
and UO_1880 (O_1880,N_24573,N_24595);
xor UO_1881 (O_1881,N_24610,N_24913);
or UO_1882 (O_1882,N_24601,N_24769);
nand UO_1883 (O_1883,N_24955,N_24523);
nor UO_1884 (O_1884,N_24978,N_24877);
and UO_1885 (O_1885,N_24642,N_24927);
and UO_1886 (O_1886,N_24923,N_24605);
nand UO_1887 (O_1887,N_24676,N_24518);
and UO_1888 (O_1888,N_24926,N_24539);
nor UO_1889 (O_1889,N_24709,N_24525);
nand UO_1890 (O_1890,N_24835,N_24836);
and UO_1891 (O_1891,N_24948,N_24526);
nor UO_1892 (O_1892,N_24695,N_24828);
and UO_1893 (O_1893,N_24617,N_24836);
nor UO_1894 (O_1894,N_24985,N_24827);
xnor UO_1895 (O_1895,N_24816,N_24557);
and UO_1896 (O_1896,N_24748,N_24906);
xor UO_1897 (O_1897,N_24614,N_24664);
and UO_1898 (O_1898,N_24766,N_24691);
or UO_1899 (O_1899,N_24636,N_24583);
nand UO_1900 (O_1900,N_24688,N_24521);
or UO_1901 (O_1901,N_24810,N_24731);
or UO_1902 (O_1902,N_24782,N_24705);
and UO_1903 (O_1903,N_24589,N_24791);
and UO_1904 (O_1904,N_24542,N_24567);
nor UO_1905 (O_1905,N_24612,N_24639);
or UO_1906 (O_1906,N_24935,N_24873);
nand UO_1907 (O_1907,N_24686,N_24626);
nand UO_1908 (O_1908,N_24881,N_24553);
or UO_1909 (O_1909,N_24795,N_24883);
nor UO_1910 (O_1910,N_24532,N_24836);
or UO_1911 (O_1911,N_24569,N_24988);
nor UO_1912 (O_1912,N_24539,N_24974);
nor UO_1913 (O_1913,N_24972,N_24575);
or UO_1914 (O_1914,N_24721,N_24503);
nand UO_1915 (O_1915,N_24877,N_24599);
or UO_1916 (O_1916,N_24874,N_24943);
or UO_1917 (O_1917,N_24633,N_24878);
nor UO_1918 (O_1918,N_24597,N_24717);
nor UO_1919 (O_1919,N_24972,N_24889);
and UO_1920 (O_1920,N_24634,N_24602);
xnor UO_1921 (O_1921,N_24527,N_24780);
nor UO_1922 (O_1922,N_24846,N_24523);
and UO_1923 (O_1923,N_24726,N_24604);
nand UO_1924 (O_1924,N_24779,N_24839);
nand UO_1925 (O_1925,N_24899,N_24722);
nor UO_1926 (O_1926,N_24771,N_24850);
nor UO_1927 (O_1927,N_24664,N_24514);
or UO_1928 (O_1928,N_24651,N_24982);
nor UO_1929 (O_1929,N_24967,N_24628);
nand UO_1930 (O_1930,N_24727,N_24774);
nand UO_1931 (O_1931,N_24719,N_24854);
or UO_1932 (O_1932,N_24819,N_24920);
nor UO_1933 (O_1933,N_24806,N_24641);
xor UO_1934 (O_1934,N_24859,N_24882);
and UO_1935 (O_1935,N_24888,N_24614);
nand UO_1936 (O_1936,N_24903,N_24508);
nor UO_1937 (O_1937,N_24985,N_24934);
and UO_1938 (O_1938,N_24804,N_24942);
nand UO_1939 (O_1939,N_24762,N_24905);
xnor UO_1940 (O_1940,N_24905,N_24538);
nor UO_1941 (O_1941,N_24982,N_24522);
nand UO_1942 (O_1942,N_24577,N_24664);
xor UO_1943 (O_1943,N_24992,N_24866);
nor UO_1944 (O_1944,N_24902,N_24614);
nand UO_1945 (O_1945,N_24625,N_24942);
nor UO_1946 (O_1946,N_24986,N_24740);
nand UO_1947 (O_1947,N_24591,N_24979);
and UO_1948 (O_1948,N_24791,N_24993);
or UO_1949 (O_1949,N_24739,N_24806);
or UO_1950 (O_1950,N_24851,N_24992);
and UO_1951 (O_1951,N_24549,N_24843);
xor UO_1952 (O_1952,N_24767,N_24788);
xnor UO_1953 (O_1953,N_24892,N_24694);
and UO_1954 (O_1954,N_24781,N_24921);
nor UO_1955 (O_1955,N_24717,N_24851);
xnor UO_1956 (O_1956,N_24867,N_24693);
nand UO_1957 (O_1957,N_24531,N_24871);
and UO_1958 (O_1958,N_24506,N_24632);
or UO_1959 (O_1959,N_24834,N_24904);
or UO_1960 (O_1960,N_24594,N_24644);
and UO_1961 (O_1961,N_24969,N_24592);
and UO_1962 (O_1962,N_24633,N_24520);
nor UO_1963 (O_1963,N_24715,N_24876);
and UO_1964 (O_1964,N_24572,N_24933);
nand UO_1965 (O_1965,N_24510,N_24967);
nand UO_1966 (O_1966,N_24866,N_24620);
or UO_1967 (O_1967,N_24706,N_24741);
xnor UO_1968 (O_1968,N_24762,N_24681);
and UO_1969 (O_1969,N_24797,N_24973);
or UO_1970 (O_1970,N_24750,N_24548);
nand UO_1971 (O_1971,N_24701,N_24758);
nand UO_1972 (O_1972,N_24778,N_24858);
and UO_1973 (O_1973,N_24702,N_24868);
and UO_1974 (O_1974,N_24691,N_24786);
and UO_1975 (O_1975,N_24942,N_24755);
nand UO_1976 (O_1976,N_24510,N_24854);
nand UO_1977 (O_1977,N_24758,N_24645);
or UO_1978 (O_1978,N_24711,N_24700);
or UO_1979 (O_1979,N_24674,N_24928);
xnor UO_1980 (O_1980,N_24540,N_24867);
and UO_1981 (O_1981,N_24801,N_24743);
nor UO_1982 (O_1982,N_24604,N_24624);
and UO_1983 (O_1983,N_24595,N_24745);
nor UO_1984 (O_1984,N_24500,N_24810);
nor UO_1985 (O_1985,N_24984,N_24913);
nand UO_1986 (O_1986,N_24518,N_24667);
and UO_1987 (O_1987,N_24848,N_24545);
and UO_1988 (O_1988,N_24666,N_24986);
or UO_1989 (O_1989,N_24825,N_24541);
xnor UO_1990 (O_1990,N_24769,N_24884);
nor UO_1991 (O_1991,N_24673,N_24683);
nand UO_1992 (O_1992,N_24834,N_24963);
nor UO_1993 (O_1993,N_24718,N_24696);
or UO_1994 (O_1994,N_24741,N_24971);
and UO_1995 (O_1995,N_24721,N_24760);
and UO_1996 (O_1996,N_24519,N_24779);
xnor UO_1997 (O_1997,N_24627,N_24986);
nand UO_1998 (O_1998,N_24993,N_24842);
nor UO_1999 (O_1999,N_24617,N_24528);
nor UO_2000 (O_2000,N_24875,N_24503);
xor UO_2001 (O_2001,N_24615,N_24618);
nor UO_2002 (O_2002,N_24845,N_24700);
xnor UO_2003 (O_2003,N_24893,N_24982);
nor UO_2004 (O_2004,N_24663,N_24811);
and UO_2005 (O_2005,N_24737,N_24994);
or UO_2006 (O_2006,N_24860,N_24528);
or UO_2007 (O_2007,N_24553,N_24932);
nand UO_2008 (O_2008,N_24983,N_24733);
or UO_2009 (O_2009,N_24520,N_24770);
nand UO_2010 (O_2010,N_24950,N_24845);
nand UO_2011 (O_2011,N_24671,N_24995);
nor UO_2012 (O_2012,N_24847,N_24941);
nand UO_2013 (O_2013,N_24568,N_24885);
and UO_2014 (O_2014,N_24635,N_24738);
and UO_2015 (O_2015,N_24784,N_24941);
or UO_2016 (O_2016,N_24693,N_24668);
and UO_2017 (O_2017,N_24807,N_24868);
or UO_2018 (O_2018,N_24586,N_24727);
nor UO_2019 (O_2019,N_24642,N_24834);
nor UO_2020 (O_2020,N_24541,N_24701);
nor UO_2021 (O_2021,N_24900,N_24846);
xor UO_2022 (O_2022,N_24529,N_24738);
nor UO_2023 (O_2023,N_24631,N_24562);
nor UO_2024 (O_2024,N_24514,N_24882);
xor UO_2025 (O_2025,N_24626,N_24972);
or UO_2026 (O_2026,N_24594,N_24786);
and UO_2027 (O_2027,N_24779,N_24679);
nor UO_2028 (O_2028,N_24842,N_24907);
and UO_2029 (O_2029,N_24757,N_24664);
nand UO_2030 (O_2030,N_24586,N_24594);
and UO_2031 (O_2031,N_24587,N_24993);
or UO_2032 (O_2032,N_24759,N_24921);
nand UO_2033 (O_2033,N_24569,N_24970);
xnor UO_2034 (O_2034,N_24877,N_24647);
or UO_2035 (O_2035,N_24659,N_24609);
xnor UO_2036 (O_2036,N_24771,N_24908);
nand UO_2037 (O_2037,N_24506,N_24757);
nand UO_2038 (O_2038,N_24928,N_24540);
xnor UO_2039 (O_2039,N_24936,N_24912);
nand UO_2040 (O_2040,N_24912,N_24661);
or UO_2041 (O_2041,N_24775,N_24830);
nand UO_2042 (O_2042,N_24617,N_24899);
nand UO_2043 (O_2043,N_24601,N_24889);
and UO_2044 (O_2044,N_24525,N_24943);
and UO_2045 (O_2045,N_24610,N_24678);
and UO_2046 (O_2046,N_24559,N_24804);
or UO_2047 (O_2047,N_24580,N_24898);
nor UO_2048 (O_2048,N_24730,N_24884);
nor UO_2049 (O_2049,N_24551,N_24702);
nor UO_2050 (O_2050,N_24524,N_24815);
nand UO_2051 (O_2051,N_24532,N_24509);
xor UO_2052 (O_2052,N_24765,N_24665);
nand UO_2053 (O_2053,N_24866,N_24951);
and UO_2054 (O_2054,N_24870,N_24696);
or UO_2055 (O_2055,N_24624,N_24777);
nor UO_2056 (O_2056,N_24842,N_24537);
xor UO_2057 (O_2057,N_24549,N_24558);
and UO_2058 (O_2058,N_24809,N_24706);
nor UO_2059 (O_2059,N_24754,N_24717);
nand UO_2060 (O_2060,N_24893,N_24653);
xor UO_2061 (O_2061,N_24621,N_24633);
nand UO_2062 (O_2062,N_24980,N_24917);
or UO_2063 (O_2063,N_24999,N_24995);
nor UO_2064 (O_2064,N_24892,N_24752);
nand UO_2065 (O_2065,N_24650,N_24932);
nand UO_2066 (O_2066,N_24857,N_24830);
nor UO_2067 (O_2067,N_24572,N_24819);
xnor UO_2068 (O_2068,N_24595,N_24597);
xnor UO_2069 (O_2069,N_24998,N_24803);
nor UO_2070 (O_2070,N_24721,N_24586);
and UO_2071 (O_2071,N_24510,N_24673);
nand UO_2072 (O_2072,N_24888,N_24799);
nor UO_2073 (O_2073,N_24912,N_24885);
xor UO_2074 (O_2074,N_24816,N_24873);
and UO_2075 (O_2075,N_24678,N_24729);
xor UO_2076 (O_2076,N_24971,N_24786);
and UO_2077 (O_2077,N_24618,N_24812);
or UO_2078 (O_2078,N_24673,N_24942);
xnor UO_2079 (O_2079,N_24619,N_24719);
and UO_2080 (O_2080,N_24614,N_24786);
nand UO_2081 (O_2081,N_24619,N_24975);
xor UO_2082 (O_2082,N_24683,N_24588);
nor UO_2083 (O_2083,N_24516,N_24810);
or UO_2084 (O_2084,N_24703,N_24775);
or UO_2085 (O_2085,N_24954,N_24815);
or UO_2086 (O_2086,N_24618,N_24577);
nand UO_2087 (O_2087,N_24860,N_24637);
or UO_2088 (O_2088,N_24803,N_24975);
or UO_2089 (O_2089,N_24668,N_24530);
nor UO_2090 (O_2090,N_24916,N_24950);
nor UO_2091 (O_2091,N_24849,N_24624);
xor UO_2092 (O_2092,N_24884,N_24900);
nor UO_2093 (O_2093,N_24508,N_24683);
and UO_2094 (O_2094,N_24730,N_24667);
or UO_2095 (O_2095,N_24966,N_24679);
nor UO_2096 (O_2096,N_24824,N_24801);
xnor UO_2097 (O_2097,N_24736,N_24648);
nand UO_2098 (O_2098,N_24505,N_24501);
and UO_2099 (O_2099,N_24926,N_24903);
nor UO_2100 (O_2100,N_24953,N_24625);
nor UO_2101 (O_2101,N_24996,N_24989);
and UO_2102 (O_2102,N_24985,N_24997);
nor UO_2103 (O_2103,N_24914,N_24698);
or UO_2104 (O_2104,N_24509,N_24994);
nor UO_2105 (O_2105,N_24595,N_24999);
nand UO_2106 (O_2106,N_24727,N_24617);
and UO_2107 (O_2107,N_24672,N_24545);
nand UO_2108 (O_2108,N_24615,N_24619);
or UO_2109 (O_2109,N_24656,N_24659);
and UO_2110 (O_2110,N_24534,N_24536);
or UO_2111 (O_2111,N_24818,N_24952);
and UO_2112 (O_2112,N_24757,N_24647);
nand UO_2113 (O_2113,N_24902,N_24635);
nand UO_2114 (O_2114,N_24927,N_24983);
nor UO_2115 (O_2115,N_24560,N_24941);
nor UO_2116 (O_2116,N_24845,N_24898);
and UO_2117 (O_2117,N_24706,N_24626);
nor UO_2118 (O_2118,N_24995,N_24698);
nand UO_2119 (O_2119,N_24908,N_24934);
nor UO_2120 (O_2120,N_24897,N_24798);
nand UO_2121 (O_2121,N_24642,N_24792);
nor UO_2122 (O_2122,N_24739,N_24554);
or UO_2123 (O_2123,N_24869,N_24813);
xnor UO_2124 (O_2124,N_24905,N_24690);
nor UO_2125 (O_2125,N_24832,N_24764);
or UO_2126 (O_2126,N_24977,N_24752);
nor UO_2127 (O_2127,N_24996,N_24663);
or UO_2128 (O_2128,N_24565,N_24835);
and UO_2129 (O_2129,N_24804,N_24908);
and UO_2130 (O_2130,N_24846,N_24995);
nor UO_2131 (O_2131,N_24786,N_24767);
and UO_2132 (O_2132,N_24863,N_24990);
and UO_2133 (O_2133,N_24949,N_24971);
nor UO_2134 (O_2134,N_24981,N_24884);
xnor UO_2135 (O_2135,N_24822,N_24631);
or UO_2136 (O_2136,N_24945,N_24625);
xor UO_2137 (O_2137,N_24523,N_24924);
xor UO_2138 (O_2138,N_24828,N_24707);
nor UO_2139 (O_2139,N_24645,N_24863);
nor UO_2140 (O_2140,N_24967,N_24758);
and UO_2141 (O_2141,N_24706,N_24562);
and UO_2142 (O_2142,N_24993,N_24657);
nor UO_2143 (O_2143,N_24624,N_24828);
and UO_2144 (O_2144,N_24904,N_24728);
xnor UO_2145 (O_2145,N_24922,N_24642);
xor UO_2146 (O_2146,N_24661,N_24866);
nand UO_2147 (O_2147,N_24973,N_24520);
nor UO_2148 (O_2148,N_24582,N_24597);
nor UO_2149 (O_2149,N_24595,N_24525);
nor UO_2150 (O_2150,N_24568,N_24519);
and UO_2151 (O_2151,N_24989,N_24986);
nor UO_2152 (O_2152,N_24644,N_24516);
or UO_2153 (O_2153,N_24565,N_24807);
xor UO_2154 (O_2154,N_24719,N_24613);
and UO_2155 (O_2155,N_24587,N_24511);
nand UO_2156 (O_2156,N_24606,N_24572);
xor UO_2157 (O_2157,N_24863,N_24605);
and UO_2158 (O_2158,N_24827,N_24612);
or UO_2159 (O_2159,N_24637,N_24944);
or UO_2160 (O_2160,N_24621,N_24965);
or UO_2161 (O_2161,N_24564,N_24638);
or UO_2162 (O_2162,N_24974,N_24577);
or UO_2163 (O_2163,N_24842,N_24825);
nand UO_2164 (O_2164,N_24661,N_24928);
nor UO_2165 (O_2165,N_24938,N_24659);
or UO_2166 (O_2166,N_24504,N_24563);
or UO_2167 (O_2167,N_24986,N_24528);
nand UO_2168 (O_2168,N_24694,N_24972);
or UO_2169 (O_2169,N_24762,N_24631);
nand UO_2170 (O_2170,N_24915,N_24781);
nand UO_2171 (O_2171,N_24600,N_24761);
or UO_2172 (O_2172,N_24655,N_24953);
and UO_2173 (O_2173,N_24628,N_24618);
xor UO_2174 (O_2174,N_24641,N_24569);
xnor UO_2175 (O_2175,N_24871,N_24907);
or UO_2176 (O_2176,N_24585,N_24933);
nor UO_2177 (O_2177,N_24866,N_24835);
xnor UO_2178 (O_2178,N_24557,N_24873);
nand UO_2179 (O_2179,N_24754,N_24715);
or UO_2180 (O_2180,N_24675,N_24613);
nor UO_2181 (O_2181,N_24932,N_24967);
xnor UO_2182 (O_2182,N_24605,N_24780);
and UO_2183 (O_2183,N_24867,N_24952);
nand UO_2184 (O_2184,N_24790,N_24804);
nor UO_2185 (O_2185,N_24563,N_24695);
or UO_2186 (O_2186,N_24716,N_24766);
or UO_2187 (O_2187,N_24855,N_24548);
and UO_2188 (O_2188,N_24610,N_24724);
or UO_2189 (O_2189,N_24564,N_24710);
and UO_2190 (O_2190,N_24690,N_24851);
nor UO_2191 (O_2191,N_24951,N_24577);
nand UO_2192 (O_2192,N_24519,N_24819);
or UO_2193 (O_2193,N_24702,N_24621);
or UO_2194 (O_2194,N_24784,N_24663);
and UO_2195 (O_2195,N_24669,N_24586);
or UO_2196 (O_2196,N_24700,N_24554);
or UO_2197 (O_2197,N_24624,N_24609);
nand UO_2198 (O_2198,N_24925,N_24789);
nor UO_2199 (O_2199,N_24893,N_24860);
nand UO_2200 (O_2200,N_24775,N_24500);
nor UO_2201 (O_2201,N_24936,N_24905);
or UO_2202 (O_2202,N_24705,N_24934);
and UO_2203 (O_2203,N_24742,N_24791);
nand UO_2204 (O_2204,N_24853,N_24565);
nand UO_2205 (O_2205,N_24679,N_24520);
and UO_2206 (O_2206,N_24947,N_24911);
or UO_2207 (O_2207,N_24502,N_24997);
nor UO_2208 (O_2208,N_24880,N_24668);
nand UO_2209 (O_2209,N_24771,N_24697);
nand UO_2210 (O_2210,N_24867,N_24590);
or UO_2211 (O_2211,N_24565,N_24619);
nor UO_2212 (O_2212,N_24798,N_24943);
nor UO_2213 (O_2213,N_24644,N_24984);
and UO_2214 (O_2214,N_24535,N_24726);
or UO_2215 (O_2215,N_24846,N_24661);
nand UO_2216 (O_2216,N_24679,N_24764);
nor UO_2217 (O_2217,N_24731,N_24821);
xnor UO_2218 (O_2218,N_24753,N_24840);
nor UO_2219 (O_2219,N_24646,N_24724);
nand UO_2220 (O_2220,N_24765,N_24532);
or UO_2221 (O_2221,N_24930,N_24939);
xor UO_2222 (O_2222,N_24646,N_24824);
xor UO_2223 (O_2223,N_24535,N_24876);
nor UO_2224 (O_2224,N_24823,N_24503);
nor UO_2225 (O_2225,N_24891,N_24718);
xnor UO_2226 (O_2226,N_24502,N_24517);
and UO_2227 (O_2227,N_24928,N_24627);
nand UO_2228 (O_2228,N_24751,N_24635);
or UO_2229 (O_2229,N_24835,N_24587);
and UO_2230 (O_2230,N_24934,N_24880);
xor UO_2231 (O_2231,N_24579,N_24783);
nor UO_2232 (O_2232,N_24565,N_24811);
and UO_2233 (O_2233,N_24667,N_24602);
xnor UO_2234 (O_2234,N_24976,N_24771);
nand UO_2235 (O_2235,N_24855,N_24716);
nand UO_2236 (O_2236,N_24960,N_24900);
or UO_2237 (O_2237,N_24552,N_24656);
and UO_2238 (O_2238,N_24522,N_24728);
nor UO_2239 (O_2239,N_24672,N_24910);
nand UO_2240 (O_2240,N_24510,N_24786);
nor UO_2241 (O_2241,N_24545,N_24582);
or UO_2242 (O_2242,N_24669,N_24945);
xnor UO_2243 (O_2243,N_24925,N_24898);
or UO_2244 (O_2244,N_24731,N_24915);
nor UO_2245 (O_2245,N_24881,N_24785);
and UO_2246 (O_2246,N_24671,N_24722);
and UO_2247 (O_2247,N_24504,N_24627);
nor UO_2248 (O_2248,N_24827,N_24737);
or UO_2249 (O_2249,N_24599,N_24866);
nor UO_2250 (O_2250,N_24678,N_24563);
xor UO_2251 (O_2251,N_24684,N_24798);
or UO_2252 (O_2252,N_24523,N_24613);
or UO_2253 (O_2253,N_24582,N_24876);
or UO_2254 (O_2254,N_24994,N_24984);
and UO_2255 (O_2255,N_24579,N_24934);
nor UO_2256 (O_2256,N_24718,N_24631);
or UO_2257 (O_2257,N_24557,N_24675);
or UO_2258 (O_2258,N_24807,N_24962);
nor UO_2259 (O_2259,N_24692,N_24634);
nand UO_2260 (O_2260,N_24992,N_24847);
nor UO_2261 (O_2261,N_24570,N_24544);
nor UO_2262 (O_2262,N_24717,N_24926);
nand UO_2263 (O_2263,N_24628,N_24719);
xnor UO_2264 (O_2264,N_24755,N_24801);
or UO_2265 (O_2265,N_24989,N_24818);
or UO_2266 (O_2266,N_24711,N_24859);
or UO_2267 (O_2267,N_24604,N_24601);
or UO_2268 (O_2268,N_24551,N_24885);
and UO_2269 (O_2269,N_24702,N_24925);
or UO_2270 (O_2270,N_24732,N_24909);
and UO_2271 (O_2271,N_24986,N_24752);
nor UO_2272 (O_2272,N_24929,N_24948);
and UO_2273 (O_2273,N_24599,N_24596);
and UO_2274 (O_2274,N_24749,N_24666);
or UO_2275 (O_2275,N_24813,N_24817);
nor UO_2276 (O_2276,N_24676,N_24839);
nor UO_2277 (O_2277,N_24816,N_24978);
or UO_2278 (O_2278,N_24941,N_24690);
or UO_2279 (O_2279,N_24910,N_24699);
xnor UO_2280 (O_2280,N_24583,N_24595);
nor UO_2281 (O_2281,N_24501,N_24793);
nand UO_2282 (O_2282,N_24962,N_24523);
nand UO_2283 (O_2283,N_24625,N_24745);
or UO_2284 (O_2284,N_24513,N_24587);
and UO_2285 (O_2285,N_24659,N_24686);
or UO_2286 (O_2286,N_24960,N_24989);
or UO_2287 (O_2287,N_24820,N_24812);
and UO_2288 (O_2288,N_24922,N_24890);
or UO_2289 (O_2289,N_24976,N_24883);
xnor UO_2290 (O_2290,N_24885,N_24871);
xor UO_2291 (O_2291,N_24639,N_24855);
or UO_2292 (O_2292,N_24902,N_24610);
nand UO_2293 (O_2293,N_24945,N_24570);
or UO_2294 (O_2294,N_24957,N_24589);
or UO_2295 (O_2295,N_24962,N_24711);
nor UO_2296 (O_2296,N_24867,N_24890);
nand UO_2297 (O_2297,N_24926,N_24892);
nor UO_2298 (O_2298,N_24609,N_24821);
nor UO_2299 (O_2299,N_24891,N_24876);
and UO_2300 (O_2300,N_24922,N_24592);
or UO_2301 (O_2301,N_24580,N_24748);
nor UO_2302 (O_2302,N_24577,N_24530);
nand UO_2303 (O_2303,N_24590,N_24727);
or UO_2304 (O_2304,N_24797,N_24572);
or UO_2305 (O_2305,N_24513,N_24617);
and UO_2306 (O_2306,N_24556,N_24852);
and UO_2307 (O_2307,N_24829,N_24815);
xnor UO_2308 (O_2308,N_24963,N_24674);
and UO_2309 (O_2309,N_24863,N_24588);
and UO_2310 (O_2310,N_24888,N_24928);
nor UO_2311 (O_2311,N_24622,N_24762);
nand UO_2312 (O_2312,N_24814,N_24729);
nor UO_2313 (O_2313,N_24669,N_24566);
nor UO_2314 (O_2314,N_24689,N_24833);
or UO_2315 (O_2315,N_24737,N_24586);
and UO_2316 (O_2316,N_24581,N_24714);
nor UO_2317 (O_2317,N_24561,N_24513);
nor UO_2318 (O_2318,N_24726,N_24950);
nand UO_2319 (O_2319,N_24583,N_24531);
or UO_2320 (O_2320,N_24640,N_24588);
or UO_2321 (O_2321,N_24638,N_24575);
nor UO_2322 (O_2322,N_24838,N_24891);
or UO_2323 (O_2323,N_24516,N_24911);
or UO_2324 (O_2324,N_24809,N_24560);
xor UO_2325 (O_2325,N_24769,N_24664);
nand UO_2326 (O_2326,N_24718,N_24693);
nor UO_2327 (O_2327,N_24609,N_24945);
and UO_2328 (O_2328,N_24763,N_24557);
nand UO_2329 (O_2329,N_24529,N_24621);
nand UO_2330 (O_2330,N_24969,N_24923);
nor UO_2331 (O_2331,N_24772,N_24763);
and UO_2332 (O_2332,N_24794,N_24765);
nor UO_2333 (O_2333,N_24652,N_24500);
nor UO_2334 (O_2334,N_24894,N_24806);
nor UO_2335 (O_2335,N_24597,N_24960);
nor UO_2336 (O_2336,N_24515,N_24673);
nor UO_2337 (O_2337,N_24580,N_24993);
or UO_2338 (O_2338,N_24578,N_24605);
and UO_2339 (O_2339,N_24680,N_24906);
or UO_2340 (O_2340,N_24835,N_24876);
nand UO_2341 (O_2341,N_24953,N_24588);
and UO_2342 (O_2342,N_24802,N_24910);
or UO_2343 (O_2343,N_24875,N_24947);
or UO_2344 (O_2344,N_24755,N_24774);
nor UO_2345 (O_2345,N_24516,N_24512);
nand UO_2346 (O_2346,N_24808,N_24574);
nor UO_2347 (O_2347,N_24988,N_24587);
nor UO_2348 (O_2348,N_24611,N_24951);
or UO_2349 (O_2349,N_24629,N_24860);
nor UO_2350 (O_2350,N_24716,N_24706);
or UO_2351 (O_2351,N_24979,N_24570);
nor UO_2352 (O_2352,N_24933,N_24841);
nand UO_2353 (O_2353,N_24929,N_24790);
and UO_2354 (O_2354,N_24601,N_24976);
xnor UO_2355 (O_2355,N_24879,N_24866);
nor UO_2356 (O_2356,N_24941,N_24959);
nor UO_2357 (O_2357,N_24917,N_24657);
nand UO_2358 (O_2358,N_24601,N_24794);
xnor UO_2359 (O_2359,N_24575,N_24600);
and UO_2360 (O_2360,N_24743,N_24566);
nand UO_2361 (O_2361,N_24540,N_24931);
nor UO_2362 (O_2362,N_24624,N_24745);
nand UO_2363 (O_2363,N_24534,N_24574);
and UO_2364 (O_2364,N_24802,N_24642);
and UO_2365 (O_2365,N_24722,N_24809);
nor UO_2366 (O_2366,N_24596,N_24810);
nand UO_2367 (O_2367,N_24557,N_24898);
nor UO_2368 (O_2368,N_24658,N_24801);
and UO_2369 (O_2369,N_24970,N_24760);
xnor UO_2370 (O_2370,N_24925,N_24543);
or UO_2371 (O_2371,N_24690,N_24856);
and UO_2372 (O_2372,N_24937,N_24691);
nand UO_2373 (O_2373,N_24527,N_24679);
or UO_2374 (O_2374,N_24539,N_24520);
nor UO_2375 (O_2375,N_24924,N_24754);
nor UO_2376 (O_2376,N_24793,N_24912);
or UO_2377 (O_2377,N_24744,N_24884);
nand UO_2378 (O_2378,N_24612,N_24635);
or UO_2379 (O_2379,N_24921,N_24613);
or UO_2380 (O_2380,N_24700,N_24827);
and UO_2381 (O_2381,N_24544,N_24704);
or UO_2382 (O_2382,N_24872,N_24655);
and UO_2383 (O_2383,N_24933,N_24714);
and UO_2384 (O_2384,N_24889,N_24659);
nand UO_2385 (O_2385,N_24703,N_24513);
and UO_2386 (O_2386,N_24946,N_24584);
nand UO_2387 (O_2387,N_24881,N_24557);
and UO_2388 (O_2388,N_24951,N_24982);
or UO_2389 (O_2389,N_24558,N_24691);
and UO_2390 (O_2390,N_24906,N_24905);
or UO_2391 (O_2391,N_24889,N_24835);
or UO_2392 (O_2392,N_24626,N_24942);
nor UO_2393 (O_2393,N_24645,N_24878);
and UO_2394 (O_2394,N_24621,N_24573);
or UO_2395 (O_2395,N_24772,N_24770);
xor UO_2396 (O_2396,N_24571,N_24812);
nor UO_2397 (O_2397,N_24685,N_24794);
nor UO_2398 (O_2398,N_24928,N_24731);
or UO_2399 (O_2399,N_24909,N_24916);
nand UO_2400 (O_2400,N_24971,N_24922);
nand UO_2401 (O_2401,N_24889,N_24748);
xnor UO_2402 (O_2402,N_24962,N_24803);
and UO_2403 (O_2403,N_24854,N_24884);
or UO_2404 (O_2404,N_24735,N_24524);
and UO_2405 (O_2405,N_24801,N_24968);
and UO_2406 (O_2406,N_24586,N_24968);
and UO_2407 (O_2407,N_24736,N_24620);
or UO_2408 (O_2408,N_24888,N_24690);
nor UO_2409 (O_2409,N_24815,N_24887);
xor UO_2410 (O_2410,N_24511,N_24606);
and UO_2411 (O_2411,N_24814,N_24879);
nor UO_2412 (O_2412,N_24607,N_24555);
nor UO_2413 (O_2413,N_24782,N_24868);
and UO_2414 (O_2414,N_24821,N_24967);
and UO_2415 (O_2415,N_24553,N_24524);
or UO_2416 (O_2416,N_24681,N_24682);
or UO_2417 (O_2417,N_24644,N_24641);
nand UO_2418 (O_2418,N_24644,N_24585);
and UO_2419 (O_2419,N_24598,N_24691);
or UO_2420 (O_2420,N_24946,N_24820);
xor UO_2421 (O_2421,N_24804,N_24654);
xor UO_2422 (O_2422,N_24847,N_24935);
or UO_2423 (O_2423,N_24688,N_24642);
or UO_2424 (O_2424,N_24589,N_24987);
xor UO_2425 (O_2425,N_24568,N_24550);
or UO_2426 (O_2426,N_24602,N_24748);
nor UO_2427 (O_2427,N_24975,N_24857);
nor UO_2428 (O_2428,N_24691,N_24680);
and UO_2429 (O_2429,N_24929,N_24710);
nand UO_2430 (O_2430,N_24678,N_24898);
and UO_2431 (O_2431,N_24646,N_24560);
or UO_2432 (O_2432,N_24815,N_24589);
nand UO_2433 (O_2433,N_24690,N_24743);
nor UO_2434 (O_2434,N_24575,N_24809);
and UO_2435 (O_2435,N_24879,N_24747);
or UO_2436 (O_2436,N_24885,N_24578);
or UO_2437 (O_2437,N_24585,N_24744);
and UO_2438 (O_2438,N_24578,N_24671);
nand UO_2439 (O_2439,N_24645,N_24779);
nand UO_2440 (O_2440,N_24694,N_24659);
nand UO_2441 (O_2441,N_24623,N_24517);
xnor UO_2442 (O_2442,N_24719,N_24853);
or UO_2443 (O_2443,N_24726,N_24811);
and UO_2444 (O_2444,N_24510,N_24745);
nand UO_2445 (O_2445,N_24794,N_24861);
nand UO_2446 (O_2446,N_24718,N_24937);
nor UO_2447 (O_2447,N_24525,N_24611);
or UO_2448 (O_2448,N_24875,N_24886);
and UO_2449 (O_2449,N_24968,N_24756);
nand UO_2450 (O_2450,N_24659,N_24838);
or UO_2451 (O_2451,N_24979,N_24817);
and UO_2452 (O_2452,N_24709,N_24824);
nand UO_2453 (O_2453,N_24835,N_24758);
nand UO_2454 (O_2454,N_24680,N_24909);
nor UO_2455 (O_2455,N_24823,N_24775);
nor UO_2456 (O_2456,N_24600,N_24882);
nor UO_2457 (O_2457,N_24683,N_24996);
nand UO_2458 (O_2458,N_24772,N_24790);
xnor UO_2459 (O_2459,N_24859,N_24574);
or UO_2460 (O_2460,N_24758,N_24666);
nor UO_2461 (O_2461,N_24989,N_24662);
and UO_2462 (O_2462,N_24519,N_24878);
and UO_2463 (O_2463,N_24586,N_24634);
and UO_2464 (O_2464,N_24818,N_24612);
nand UO_2465 (O_2465,N_24859,N_24759);
xnor UO_2466 (O_2466,N_24895,N_24857);
xor UO_2467 (O_2467,N_24735,N_24856);
and UO_2468 (O_2468,N_24818,N_24979);
or UO_2469 (O_2469,N_24589,N_24652);
nand UO_2470 (O_2470,N_24768,N_24873);
or UO_2471 (O_2471,N_24595,N_24741);
nand UO_2472 (O_2472,N_24961,N_24639);
nor UO_2473 (O_2473,N_24514,N_24758);
nor UO_2474 (O_2474,N_24957,N_24557);
nand UO_2475 (O_2475,N_24961,N_24559);
nand UO_2476 (O_2476,N_24956,N_24788);
nand UO_2477 (O_2477,N_24962,N_24994);
nand UO_2478 (O_2478,N_24661,N_24628);
nor UO_2479 (O_2479,N_24901,N_24935);
nand UO_2480 (O_2480,N_24773,N_24962);
or UO_2481 (O_2481,N_24598,N_24729);
nand UO_2482 (O_2482,N_24507,N_24982);
or UO_2483 (O_2483,N_24646,N_24738);
nor UO_2484 (O_2484,N_24577,N_24682);
or UO_2485 (O_2485,N_24589,N_24574);
nor UO_2486 (O_2486,N_24897,N_24645);
and UO_2487 (O_2487,N_24918,N_24667);
and UO_2488 (O_2488,N_24611,N_24631);
or UO_2489 (O_2489,N_24539,N_24640);
nand UO_2490 (O_2490,N_24540,N_24969);
nor UO_2491 (O_2491,N_24872,N_24520);
nor UO_2492 (O_2492,N_24821,N_24807);
and UO_2493 (O_2493,N_24713,N_24544);
nand UO_2494 (O_2494,N_24657,N_24543);
or UO_2495 (O_2495,N_24890,N_24842);
xnor UO_2496 (O_2496,N_24534,N_24765);
nand UO_2497 (O_2497,N_24819,N_24682);
or UO_2498 (O_2498,N_24968,N_24841);
or UO_2499 (O_2499,N_24621,N_24779);
nor UO_2500 (O_2500,N_24581,N_24944);
nand UO_2501 (O_2501,N_24664,N_24906);
nor UO_2502 (O_2502,N_24540,N_24631);
xnor UO_2503 (O_2503,N_24840,N_24574);
or UO_2504 (O_2504,N_24563,N_24585);
and UO_2505 (O_2505,N_24686,N_24873);
xor UO_2506 (O_2506,N_24756,N_24515);
and UO_2507 (O_2507,N_24869,N_24554);
or UO_2508 (O_2508,N_24616,N_24746);
xor UO_2509 (O_2509,N_24630,N_24646);
nor UO_2510 (O_2510,N_24529,N_24899);
or UO_2511 (O_2511,N_24877,N_24817);
and UO_2512 (O_2512,N_24743,N_24632);
and UO_2513 (O_2513,N_24786,N_24728);
or UO_2514 (O_2514,N_24995,N_24891);
nand UO_2515 (O_2515,N_24981,N_24935);
or UO_2516 (O_2516,N_24788,N_24992);
and UO_2517 (O_2517,N_24630,N_24828);
or UO_2518 (O_2518,N_24604,N_24628);
nor UO_2519 (O_2519,N_24976,N_24929);
nor UO_2520 (O_2520,N_24535,N_24613);
nand UO_2521 (O_2521,N_24832,N_24508);
and UO_2522 (O_2522,N_24551,N_24925);
or UO_2523 (O_2523,N_24652,N_24861);
xor UO_2524 (O_2524,N_24811,N_24649);
and UO_2525 (O_2525,N_24925,N_24505);
xor UO_2526 (O_2526,N_24889,N_24921);
and UO_2527 (O_2527,N_24618,N_24851);
and UO_2528 (O_2528,N_24802,N_24588);
xor UO_2529 (O_2529,N_24591,N_24958);
and UO_2530 (O_2530,N_24540,N_24597);
nor UO_2531 (O_2531,N_24939,N_24520);
nor UO_2532 (O_2532,N_24987,N_24793);
nor UO_2533 (O_2533,N_24644,N_24966);
and UO_2534 (O_2534,N_24957,N_24574);
or UO_2535 (O_2535,N_24549,N_24935);
nand UO_2536 (O_2536,N_24850,N_24862);
nor UO_2537 (O_2537,N_24922,N_24930);
or UO_2538 (O_2538,N_24760,N_24624);
nand UO_2539 (O_2539,N_24687,N_24542);
nor UO_2540 (O_2540,N_24983,N_24505);
nand UO_2541 (O_2541,N_24510,N_24853);
nor UO_2542 (O_2542,N_24746,N_24747);
and UO_2543 (O_2543,N_24895,N_24518);
nor UO_2544 (O_2544,N_24896,N_24890);
and UO_2545 (O_2545,N_24750,N_24575);
nand UO_2546 (O_2546,N_24508,N_24940);
nand UO_2547 (O_2547,N_24963,N_24584);
or UO_2548 (O_2548,N_24759,N_24748);
or UO_2549 (O_2549,N_24857,N_24571);
xor UO_2550 (O_2550,N_24789,N_24595);
nor UO_2551 (O_2551,N_24916,N_24828);
nand UO_2552 (O_2552,N_24746,N_24671);
and UO_2553 (O_2553,N_24582,N_24955);
and UO_2554 (O_2554,N_24682,N_24958);
or UO_2555 (O_2555,N_24637,N_24772);
and UO_2556 (O_2556,N_24533,N_24514);
nor UO_2557 (O_2557,N_24994,N_24691);
nand UO_2558 (O_2558,N_24982,N_24967);
nand UO_2559 (O_2559,N_24980,N_24907);
or UO_2560 (O_2560,N_24727,N_24854);
nor UO_2561 (O_2561,N_24703,N_24529);
xor UO_2562 (O_2562,N_24802,N_24872);
nand UO_2563 (O_2563,N_24539,N_24795);
nor UO_2564 (O_2564,N_24831,N_24568);
nand UO_2565 (O_2565,N_24805,N_24767);
nand UO_2566 (O_2566,N_24840,N_24851);
and UO_2567 (O_2567,N_24598,N_24874);
or UO_2568 (O_2568,N_24872,N_24719);
or UO_2569 (O_2569,N_24930,N_24706);
nor UO_2570 (O_2570,N_24708,N_24939);
nor UO_2571 (O_2571,N_24795,N_24747);
or UO_2572 (O_2572,N_24712,N_24728);
and UO_2573 (O_2573,N_24622,N_24994);
xnor UO_2574 (O_2574,N_24769,N_24693);
and UO_2575 (O_2575,N_24763,N_24740);
and UO_2576 (O_2576,N_24794,N_24558);
and UO_2577 (O_2577,N_24961,N_24786);
xnor UO_2578 (O_2578,N_24984,N_24599);
and UO_2579 (O_2579,N_24598,N_24997);
and UO_2580 (O_2580,N_24560,N_24773);
nand UO_2581 (O_2581,N_24919,N_24622);
and UO_2582 (O_2582,N_24783,N_24673);
nor UO_2583 (O_2583,N_24531,N_24869);
or UO_2584 (O_2584,N_24509,N_24607);
nor UO_2585 (O_2585,N_24586,N_24609);
nand UO_2586 (O_2586,N_24814,N_24770);
nor UO_2587 (O_2587,N_24721,N_24990);
nor UO_2588 (O_2588,N_24950,N_24967);
nor UO_2589 (O_2589,N_24969,N_24965);
or UO_2590 (O_2590,N_24511,N_24500);
nor UO_2591 (O_2591,N_24732,N_24932);
nor UO_2592 (O_2592,N_24521,N_24631);
nor UO_2593 (O_2593,N_24981,N_24644);
and UO_2594 (O_2594,N_24849,N_24683);
nand UO_2595 (O_2595,N_24954,N_24700);
and UO_2596 (O_2596,N_24685,N_24810);
nand UO_2597 (O_2597,N_24648,N_24777);
and UO_2598 (O_2598,N_24507,N_24665);
nor UO_2599 (O_2599,N_24600,N_24692);
nand UO_2600 (O_2600,N_24779,N_24810);
and UO_2601 (O_2601,N_24731,N_24627);
nor UO_2602 (O_2602,N_24571,N_24794);
nor UO_2603 (O_2603,N_24847,N_24903);
nor UO_2604 (O_2604,N_24780,N_24516);
or UO_2605 (O_2605,N_24603,N_24973);
and UO_2606 (O_2606,N_24808,N_24798);
nand UO_2607 (O_2607,N_24943,N_24589);
nand UO_2608 (O_2608,N_24961,N_24765);
and UO_2609 (O_2609,N_24977,N_24598);
nor UO_2610 (O_2610,N_24889,N_24586);
nand UO_2611 (O_2611,N_24843,N_24906);
nand UO_2612 (O_2612,N_24793,N_24972);
nor UO_2613 (O_2613,N_24901,N_24687);
nand UO_2614 (O_2614,N_24999,N_24965);
nand UO_2615 (O_2615,N_24571,N_24870);
and UO_2616 (O_2616,N_24658,N_24779);
or UO_2617 (O_2617,N_24637,N_24697);
or UO_2618 (O_2618,N_24675,N_24758);
nor UO_2619 (O_2619,N_24955,N_24681);
nor UO_2620 (O_2620,N_24587,N_24844);
and UO_2621 (O_2621,N_24642,N_24612);
nor UO_2622 (O_2622,N_24905,N_24745);
nor UO_2623 (O_2623,N_24967,N_24918);
or UO_2624 (O_2624,N_24742,N_24980);
and UO_2625 (O_2625,N_24521,N_24562);
and UO_2626 (O_2626,N_24697,N_24645);
and UO_2627 (O_2627,N_24743,N_24963);
nand UO_2628 (O_2628,N_24722,N_24805);
and UO_2629 (O_2629,N_24797,N_24541);
nor UO_2630 (O_2630,N_24650,N_24931);
nand UO_2631 (O_2631,N_24955,N_24608);
nand UO_2632 (O_2632,N_24551,N_24879);
nor UO_2633 (O_2633,N_24941,N_24500);
nor UO_2634 (O_2634,N_24692,N_24909);
and UO_2635 (O_2635,N_24707,N_24606);
nand UO_2636 (O_2636,N_24525,N_24554);
nor UO_2637 (O_2637,N_24957,N_24836);
nand UO_2638 (O_2638,N_24989,N_24711);
nor UO_2639 (O_2639,N_24724,N_24899);
nand UO_2640 (O_2640,N_24692,N_24857);
and UO_2641 (O_2641,N_24737,N_24932);
or UO_2642 (O_2642,N_24571,N_24819);
and UO_2643 (O_2643,N_24551,N_24731);
nor UO_2644 (O_2644,N_24825,N_24935);
and UO_2645 (O_2645,N_24604,N_24961);
nand UO_2646 (O_2646,N_24944,N_24769);
and UO_2647 (O_2647,N_24731,N_24623);
and UO_2648 (O_2648,N_24854,N_24722);
and UO_2649 (O_2649,N_24854,N_24583);
or UO_2650 (O_2650,N_24787,N_24892);
nor UO_2651 (O_2651,N_24873,N_24504);
and UO_2652 (O_2652,N_24834,N_24940);
nand UO_2653 (O_2653,N_24924,N_24659);
xnor UO_2654 (O_2654,N_24854,N_24753);
nor UO_2655 (O_2655,N_24509,N_24521);
and UO_2656 (O_2656,N_24672,N_24805);
or UO_2657 (O_2657,N_24638,N_24737);
nor UO_2658 (O_2658,N_24649,N_24628);
nand UO_2659 (O_2659,N_24743,N_24643);
xnor UO_2660 (O_2660,N_24622,N_24525);
nor UO_2661 (O_2661,N_24664,N_24891);
or UO_2662 (O_2662,N_24883,N_24807);
nor UO_2663 (O_2663,N_24532,N_24541);
or UO_2664 (O_2664,N_24567,N_24649);
nor UO_2665 (O_2665,N_24609,N_24580);
nand UO_2666 (O_2666,N_24878,N_24740);
nand UO_2667 (O_2667,N_24515,N_24657);
nand UO_2668 (O_2668,N_24749,N_24533);
nand UO_2669 (O_2669,N_24692,N_24822);
or UO_2670 (O_2670,N_24623,N_24779);
or UO_2671 (O_2671,N_24788,N_24999);
or UO_2672 (O_2672,N_24955,N_24978);
nor UO_2673 (O_2673,N_24951,N_24556);
xor UO_2674 (O_2674,N_24874,N_24974);
nand UO_2675 (O_2675,N_24962,N_24567);
and UO_2676 (O_2676,N_24749,N_24586);
nand UO_2677 (O_2677,N_24906,N_24603);
nand UO_2678 (O_2678,N_24802,N_24530);
nand UO_2679 (O_2679,N_24873,N_24749);
or UO_2680 (O_2680,N_24678,N_24936);
nor UO_2681 (O_2681,N_24668,N_24864);
and UO_2682 (O_2682,N_24943,N_24666);
or UO_2683 (O_2683,N_24685,N_24793);
xnor UO_2684 (O_2684,N_24981,N_24914);
or UO_2685 (O_2685,N_24670,N_24627);
xor UO_2686 (O_2686,N_24900,N_24656);
nand UO_2687 (O_2687,N_24940,N_24999);
and UO_2688 (O_2688,N_24711,N_24766);
nand UO_2689 (O_2689,N_24731,N_24728);
nand UO_2690 (O_2690,N_24781,N_24731);
and UO_2691 (O_2691,N_24607,N_24712);
nor UO_2692 (O_2692,N_24599,N_24749);
and UO_2693 (O_2693,N_24814,N_24517);
nand UO_2694 (O_2694,N_24572,N_24924);
nor UO_2695 (O_2695,N_24686,N_24557);
xnor UO_2696 (O_2696,N_24878,N_24840);
and UO_2697 (O_2697,N_24927,N_24972);
and UO_2698 (O_2698,N_24938,N_24572);
and UO_2699 (O_2699,N_24794,N_24721);
nor UO_2700 (O_2700,N_24908,N_24513);
nand UO_2701 (O_2701,N_24926,N_24725);
nand UO_2702 (O_2702,N_24609,N_24901);
and UO_2703 (O_2703,N_24584,N_24830);
nand UO_2704 (O_2704,N_24522,N_24761);
nor UO_2705 (O_2705,N_24915,N_24821);
nor UO_2706 (O_2706,N_24564,N_24758);
nor UO_2707 (O_2707,N_24928,N_24523);
or UO_2708 (O_2708,N_24545,N_24966);
or UO_2709 (O_2709,N_24532,N_24692);
xnor UO_2710 (O_2710,N_24594,N_24910);
and UO_2711 (O_2711,N_24798,N_24888);
or UO_2712 (O_2712,N_24860,N_24536);
xor UO_2713 (O_2713,N_24587,N_24864);
and UO_2714 (O_2714,N_24725,N_24816);
and UO_2715 (O_2715,N_24659,N_24581);
or UO_2716 (O_2716,N_24974,N_24937);
nor UO_2717 (O_2717,N_24566,N_24822);
nor UO_2718 (O_2718,N_24543,N_24969);
and UO_2719 (O_2719,N_24940,N_24690);
nor UO_2720 (O_2720,N_24899,N_24888);
xnor UO_2721 (O_2721,N_24568,N_24551);
nand UO_2722 (O_2722,N_24629,N_24535);
nor UO_2723 (O_2723,N_24637,N_24515);
or UO_2724 (O_2724,N_24960,N_24686);
xnor UO_2725 (O_2725,N_24809,N_24800);
and UO_2726 (O_2726,N_24880,N_24858);
nor UO_2727 (O_2727,N_24860,N_24504);
nor UO_2728 (O_2728,N_24905,N_24526);
or UO_2729 (O_2729,N_24956,N_24771);
nor UO_2730 (O_2730,N_24703,N_24802);
or UO_2731 (O_2731,N_24970,N_24588);
or UO_2732 (O_2732,N_24648,N_24765);
and UO_2733 (O_2733,N_24614,N_24735);
and UO_2734 (O_2734,N_24921,N_24535);
and UO_2735 (O_2735,N_24522,N_24922);
nor UO_2736 (O_2736,N_24911,N_24714);
nand UO_2737 (O_2737,N_24560,N_24970);
nand UO_2738 (O_2738,N_24676,N_24941);
or UO_2739 (O_2739,N_24597,N_24666);
or UO_2740 (O_2740,N_24672,N_24607);
xnor UO_2741 (O_2741,N_24703,N_24569);
or UO_2742 (O_2742,N_24734,N_24559);
nor UO_2743 (O_2743,N_24946,N_24763);
nor UO_2744 (O_2744,N_24692,N_24948);
nand UO_2745 (O_2745,N_24590,N_24917);
nor UO_2746 (O_2746,N_24916,N_24832);
nand UO_2747 (O_2747,N_24929,N_24585);
or UO_2748 (O_2748,N_24640,N_24711);
nor UO_2749 (O_2749,N_24648,N_24694);
and UO_2750 (O_2750,N_24694,N_24895);
or UO_2751 (O_2751,N_24929,N_24756);
nor UO_2752 (O_2752,N_24655,N_24802);
nor UO_2753 (O_2753,N_24911,N_24711);
nand UO_2754 (O_2754,N_24926,N_24626);
nor UO_2755 (O_2755,N_24781,N_24926);
nand UO_2756 (O_2756,N_24664,N_24716);
nand UO_2757 (O_2757,N_24980,N_24592);
nand UO_2758 (O_2758,N_24574,N_24873);
nor UO_2759 (O_2759,N_24745,N_24844);
nor UO_2760 (O_2760,N_24905,N_24874);
nand UO_2761 (O_2761,N_24838,N_24635);
nor UO_2762 (O_2762,N_24923,N_24688);
and UO_2763 (O_2763,N_24904,N_24958);
or UO_2764 (O_2764,N_24807,N_24875);
or UO_2765 (O_2765,N_24582,N_24500);
nor UO_2766 (O_2766,N_24541,N_24547);
or UO_2767 (O_2767,N_24758,N_24729);
xnor UO_2768 (O_2768,N_24708,N_24679);
xnor UO_2769 (O_2769,N_24603,N_24650);
or UO_2770 (O_2770,N_24819,N_24995);
or UO_2771 (O_2771,N_24848,N_24872);
or UO_2772 (O_2772,N_24811,N_24677);
and UO_2773 (O_2773,N_24861,N_24592);
nor UO_2774 (O_2774,N_24554,N_24641);
nor UO_2775 (O_2775,N_24909,N_24606);
nand UO_2776 (O_2776,N_24845,N_24578);
and UO_2777 (O_2777,N_24966,N_24624);
nor UO_2778 (O_2778,N_24693,N_24521);
and UO_2779 (O_2779,N_24967,N_24702);
and UO_2780 (O_2780,N_24757,N_24684);
nand UO_2781 (O_2781,N_24688,N_24518);
or UO_2782 (O_2782,N_24968,N_24910);
or UO_2783 (O_2783,N_24980,N_24672);
nand UO_2784 (O_2784,N_24798,N_24699);
or UO_2785 (O_2785,N_24863,N_24705);
and UO_2786 (O_2786,N_24597,N_24746);
nor UO_2787 (O_2787,N_24885,N_24794);
or UO_2788 (O_2788,N_24841,N_24838);
and UO_2789 (O_2789,N_24932,N_24546);
or UO_2790 (O_2790,N_24718,N_24571);
or UO_2791 (O_2791,N_24769,N_24966);
and UO_2792 (O_2792,N_24795,N_24988);
nand UO_2793 (O_2793,N_24731,N_24658);
xor UO_2794 (O_2794,N_24532,N_24543);
nor UO_2795 (O_2795,N_24627,N_24762);
xnor UO_2796 (O_2796,N_24828,N_24734);
nor UO_2797 (O_2797,N_24911,N_24632);
or UO_2798 (O_2798,N_24770,N_24533);
and UO_2799 (O_2799,N_24772,N_24908);
or UO_2800 (O_2800,N_24870,N_24619);
and UO_2801 (O_2801,N_24670,N_24744);
or UO_2802 (O_2802,N_24501,N_24595);
xor UO_2803 (O_2803,N_24703,N_24931);
nand UO_2804 (O_2804,N_24825,N_24863);
or UO_2805 (O_2805,N_24703,N_24571);
nor UO_2806 (O_2806,N_24781,N_24817);
xnor UO_2807 (O_2807,N_24568,N_24975);
and UO_2808 (O_2808,N_24592,N_24819);
and UO_2809 (O_2809,N_24601,N_24798);
nand UO_2810 (O_2810,N_24727,N_24940);
xnor UO_2811 (O_2811,N_24527,N_24799);
or UO_2812 (O_2812,N_24654,N_24663);
nand UO_2813 (O_2813,N_24933,N_24794);
and UO_2814 (O_2814,N_24521,N_24861);
and UO_2815 (O_2815,N_24522,N_24968);
nor UO_2816 (O_2816,N_24749,N_24915);
or UO_2817 (O_2817,N_24915,N_24737);
nor UO_2818 (O_2818,N_24970,N_24601);
xnor UO_2819 (O_2819,N_24865,N_24973);
nand UO_2820 (O_2820,N_24827,N_24613);
or UO_2821 (O_2821,N_24827,N_24739);
nor UO_2822 (O_2822,N_24574,N_24564);
and UO_2823 (O_2823,N_24636,N_24651);
nand UO_2824 (O_2824,N_24558,N_24857);
and UO_2825 (O_2825,N_24740,N_24694);
and UO_2826 (O_2826,N_24751,N_24990);
nor UO_2827 (O_2827,N_24845,N_24816);
xnor UO_2828 (O_2828,N_24944,N_24767);
xnor UO_2829 (O_2829,N_24707,N_24771);
and UO_2830 (O_2830,N_24771,N_24884);
and UO_2831 (O_2831,N_24837,N_24724);
or UO_2832 (O_2832,N_24653,N_24560);
or UO_2833 (O_2833,N_24984,N_24617);
nand UO_2834 (O_2834,N_24509,N_24889);
nand UO_2835 (O_2835,N_24923,N_24976);
nor UO_2836 (O_2836,N_24712,N_24969);
nand UO_2837 (O_2837,N_24537,N_24900);
and UO_2838 (O_2838,N_24973,N_24871);
or UO_2839 (O_2839,N_24814,N_24932);
nor UO_2840 (O_2840,N_24836,N_24761);
nor UO_2841 (O_2841,N_24753,N_24794);
and UO_2842 (O_2842,N_24927,N_24526);
and UO_2843 (O_2843,N_24931,N_24778);
or UO_2844 (O_2844,N_24873,N_24622);
and UO_2845 (O_2845,N_24874,N_24991);
nor UO_2846 (O_2846,N_24909,N_24931);
and UO_2847 (O_2847,N_24657,N_24908);
or UO_2848 (O_2848,N_24903,N_24816);
nand UO_2849 (O_2849,N_24780,N_24954);
or UO_2850 (O_2850,N_24952,N_24513);
or UO_2851 (O_2851,N_24960,N_24973);
or UO_2852 (O_2852,N_24603,N_24934);
and UO_2853 (O_2853,N_24642,N_24828);
nand UO_2854 (O_2854,N_24545,N_24521);
nand UO_2855 (O_2855,N_24570,N_24913);
nand UO_2856 (O_2856,N_24561,N_24740);
or UO_2857 (O_2857,N_24862,N_24580);
or UO_2858 (O_2858,N_24678,N_24721);
and UO_2859 (O_2859,N_24787,N_24665);
nor UO_2860 (O_2860,N_24719,N_24644);
and UO_2861 (O_2861,N_24753,N_24716);
nand UO_2862 (O_2862,N_24585,N_24891);
or UO_2863 (O_2863,N_24538,N_24763);
nand UO_2864 (O_2864,N_24639,N_24514);
or UO_2865 (O_2865,N_24658,N_24874);
or UO_2866 (O_2866,N_24775,N_24897);
nand UO_2867 (O_2867,N_24677,N_24549);
nand UO_2868 (O_2868,N_24865,N_24963);
or UO_2869 (O_2869,N_24887,N_24556);
nand UO_2870 (O_2870,N_24887,N_24696);
or UO_2871 (O_2871,N_24531,N_24732);
nand UO_2872 (O_2872,N_24678,N_24889);
or UO_2873 (O_2873,N_24882,N_24618);
or UO_2874 (O_2874,N_24728,N_24647);
nor UO_2875 (O_2875,N_24650,N_24503);
or UO_2876 (O_2876,N_24859,N_24775);
and UO_2877 (O_2877,N_24942,N_24774);
xor UO_2878 (O_2878,N_24723,N_24574);
or UO_2879 (O_2879,N_24696,N_24531);
and UO_2880 (O_2880,N_24777,N_24991);
nand UO_2881 (O_2881,N_24898,N_24983);
and UO_2882 (O_2882,N_24683,N_24974);
nand UO_2883 (O_2883,N_24978,N_24771);
nand UO_2884 (O_2884,N_24902,N_24586);
nand UO_2885 (O_2885,N_24679,N_24780);
or UO_2886 (O_2886,N_24615,N_24941);
nand UO_2887 (O_2887,N_24665,N_24772);
nand UO_2888 (O_2888,N_24900,N_24987);
xnor UO_2889 (O_2889,N_24524,N_24896);
xor UO_2890 (O_2890,N_24852,N_24684);
nor UO_2891 (O_2891,N_24765,N_24539);
and UO_2892 (O_2892,N_24961,N_24999);
nor UO_2893 (O_2893,N_24986,N_24932);
nor UO_2894 (O_2894,N_24789,N_24772);
nor UO_2895 (O_2895,N_24774,N_24543);
or UO_2896 (O_2896,N_24506,N_24508);
and UO_2897 (O_2897,N_24672,N_24564);
and UO_2898 (O_2898,N_24729,N_24618);
or UO_2899 (O_2899,N_24961,N_24752);
and UO_2900 (O_2900,N_24806,N_24586);
nand UO_2901 (O_2901,N_24723,N_24615);
nand UO_2902 (O_2902,N_24852,N_24673);
and UO_2903 (O_2903,N_24820,N_24630);
and UO_2904 (O_2904,N_24511,N_24505);
or UO_2905 (O_2905,N_24814,N_24976);
or UO_2906 (O_2906,N_24624,N_24601);
and UO_2907 (O_2907,N_24503,N_24780);
and UO_2908 (O_2908,N_24818,N_24561);
and UO_2909 (O_2909,N_24513,N_24681);
nand UO_2910 (O_2910,N_24607,N_24502);
or UO_2911 (O_2911,N_24680,N_24727);
nor UO_2912 (O_2912,N_24777,N_24663);
and UO_2913 (O_2913,N_24919,N_24688);
nand UO_2914 (O_2914,N_24940,N_24823);
nand UO_2915 (O_2915,N_24644,N_24995);
nand UO_2916 (O_2916,N_24596,N_24907);
xnor UO_2917 (O_2917,N_24788,N_24914);
and UO_2918 (O_2918,N_24772,N_24771);
or UO_2919 (O_2919,N_24958,N_24802);
or UO_2920 (O_2920,N_24908,N_24562);
and UO_2921 (O_2921,N_24981,N_24888);
nor UO_2922 (O_2922,N_24561,N_24953);
and UO_2923 (O_2923,N_24552,N_24908);
nor UO_2924 (O_2924,N_24640,N_24609);
or UO_2925 (O_2925,N_24988,N_24748);
nor UO_2926 (O_2926,N_24540,N_24926);
nand UO_2927 (O_2927,N_24504,N_24868);
nor UO_2928 (O_2928,N_24794,N_24510);
or UO_2929 (O_2929,N_24867,N_24731);
xor UO_2930 (O_2930,N_24653,N_24857);
nand UO_2931 (O_2931,N_24938,N_24918);
or UO_2932 (O_2932,N_24926,N_24710);
or UO_2933 (O_2933,N_24936,N_24537);
and UO_2934 (O_2934,N_24840,N_24524);
nand UO_2935 (O_2935,N_24655,N_24859);
or UO_2936 (O_2936,N_24647,N_24713);
nand UO_2937 (O_2937,N_24887,N_24602);
nor UO_2938 (O_2938,N_24775,N_24592);
nor UO_2939 (O_2939,N_24831,N_24997);
xnor UO_2940 (O_2940,N_24529,N_24706);
and UO_2941 (O_2941,N_24714,N_24580);
xnor UO_2942 (O_2942,N_24964,N_24619);
nand UO_2943 (O_2943,N_24977,N_24510);
or UO_2944 (O_2944,N_24768,N_24829);
or UO_2945 (O_2945,N_24667,N_24529);
or UO_2946 (O_2946,N_24736,N_24895);
xor UO_2947 (O_2947,N_24515,N_24760);
and UO_2948 (O_2948,N_24793,N_24924);
xnor UO_2949 (O_2949,N_24972,N_24876);
and UO_2950 (O_2950,N_24538,N_24564);
nor UO_2951 (O_2951,N_24547,N_24731);
and UO_2952 (O_2952,N_24579,N_24878);
and UO_2953 (O_2953,N_24825,N_24711);
and UO_2954 (O_2954,N_24689,N_24507);
nor UO_2955 (O_2955,N_24909,N_24676);
and UO_2956 (O_2956,N_24788,N_24792);
or UO_2957 (O_2957,N_24989,N_24712);
nor UO_2958 (O_2958,N_24769,N_24993);
and UO_2959 (O_2959,N_24717,N_24771);
and UO_2960 (O_2960,N_24666,N_24661);
or UO_2961 (O_2961,N_24847,N_24660);
or UO_2962 (O_2962,N_24700,N_24970);
xor UO_2963 (O_2963,N_24595,N_24984);
and UO_2964 (O_2964,N_24847,N_24925);
and UO_2965 (O_2965,N_24764,N_24521);
xnor UO_2966 (O_2966,N_24971,N_24884);
nor UO_2967 (O_2967,N_24544,N_24692);
nand UO_2968 (O_2968,N_24968,N_24807);
and UO_2969 (O_2969,N_24700,N_24993);
nand UO_2970 (O_2970,N_24975,N_24899);
or UO_2971 (O_2971,N_24646,N_24683);
or UO_2972 (O_2972,N_24866,N_24960);
and UO_2973 (O_2973,N_24527,N_24514);
nand UO_2974 (O_2974,N_24791,N_24874);
and UO_2975 (O_2975,N_24760,N_24944);
or UO_2976 (O_2976,N_24676,N_24536);
or UO_2977 (O_2977,N_24778,N_24888);
or UO_2978 (O_2978,N_24585,N_24782);
xnor UO_2979 (O_2979,N_24841,N_24542);
and UO_2980 (O_2980,N_24636,N_24999);
or UO_2981 (O_2981,N_24601,N_24692);
and UO_2982 (O_2982,N_24727,N_24924);
nand UO_2983 (O_2983,N_24781,N_24587);
and UO_2984 (O_2984,N_24696,N_24742);
or UO_2985 (O_2985,N_24854,N_24607);
nand UO_2986 (O_2986,N_24697,N_24530);
xnor UO_2987 (O_2987,N_24785,N_24733);
and UO_2988 (O_2988,N_24732,N_24903);
and UO_2989 (O_2989,N_24794,N_24968);
xor UO_2990 (O_2990,N_24577,N_24875);
xor UO_2991 (O_2991,N_24595,N_24683);
nor UO_2992 (O_2992,N_24775,N_24572);
or UO_2993 (O_2993,N_24992,N_24672);
xor UO_2994 (O_2994,N_24858,N_24694);
nand UO_2995 (O_2995,N_24681,N_24560);
and UO_2996 (O_2996,N_24683,N_24858);
and UO_2997 (O_2997,N_24517,N_24972);
or UO_2998 (O_2998,N_24916,N_24805);
nand UO_2999 (O_2999,N_24507,N_24814);
endmodule