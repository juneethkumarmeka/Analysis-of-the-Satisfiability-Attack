module basic_750_5000_1000_2_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2501,N_2502,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2543,N_2544,N_2546,N_2547,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2566,N_2567,N_2568,N_2569,N_2571,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2584,N_2586,N_2588,N_2589,N_2590,N_2591,N_2592,N_2594,N_2595,N_2596,N_2597,N_2598,N_2600,N_2601,N_2602,N_2603,N_2604,N_2607,N_2608,N_2609,N_2611,N_2613,N_2614,N_2616,N_2617,N_2619,N_2620,N_2621,N_2623,N_2624,N_2625,N_2626,N_2629,N_2630,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2645,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2664,N_2665,N_2666,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2693,N_2694,N_2696,N_2698,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2714,N_2716,N_2718,N_2719,N_2720,N_2722,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2759,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2771,N_2772,N_2773,N_2774,N_2776,N_2777,N_2779,N_2780,N_2781,N_2783,N_2785,N_2787,N_2788,N_2789,N_2793,N_2794,N_2796,N_2798,N_2799,N_2800,N_2804,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2829,N_2830,N_2833,N_2834,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2845,N_2846,N_2847,N_2848,N_2851,N_2852,N_2853,N_2855,N_2856,N_2857,N_2859,N_2862,N_2863,N_2865,N_2866,N_2867,N_2870,N_2872,N_2873,N_2874,N_2875,N_2876,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2887,N_2888,N_2890,N_2891,N_2892,N_2894,N_2895,N_2896,N_2897,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2909,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2941,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2954,N_2955,N_2956,N_2957,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2978,N_2979,N_2980,N_2981,N_2982,N_2984,N_2985,N_2986,N_2988,N_2989,N_2990,N_2991,N_2993,N_2994,N_2995,N_2997,N_2998,N_2999,N_3001,N_3002,N_3003,N_3004,N_3006,N_3007,N_3008,N_3009,N_3010,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3019,N_3020,N_3021,N_3023,N_3024,N_3026,N_3027,N_3028,N_3029,N_3030,N_3032,N_3034,N_3035,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3044,N_3046,N_3047,N_3048,N_3049,N_3050,N_3052,N_3053,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3073,N_3074,N_3075,N_3077,N_3078,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3087,N_3088,N_3089,N_3090,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3101,N_3102,N_3104,N_3106,N_3107,N_3108,N_3110,N_3112,N_3113,N_3115,N_3116,N_3117,N_3119,N_3120,N_3121,N_3122,N_3123,N_3125,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3136,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3145,N_3146,N_3148,N_3150,N_3152,N_3153,N_3156,N_3158,N_3159,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3178,N_3179,N_3180,N_3182,N_3186,N_3188,N_3189,N_3190,N_3193,N_3194,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3235,N_3237,N_3238,N_3239,N_3240,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3252,N_3254,N_3255,N_3257,N_3258,N_3260,N_3261,N_3262,N_3263,N_3264,N_3267,N_3269,N_3270,N_3271,N_3272,N_3273,N_3276,N_3278,N_3280,N_3281,N_3282,N_3283,N_3285,N_3286,N_3287,N_3289,N_3291,N_3292,N_3294,N_3295,N_3298,N_3299,N_3300,N_3302,N_3303,N_3305,N_3306,N_3307,N_3308,N_3310,N_3311,N_3314,N_3318,N_3321,N_3322,N_3323,N_3324,N_3325,N_3327,N_3328,N_3329,N_3330,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3342,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3366,N_3368,N_3369,N_3370,N_3372,N_3373,N_3375,N_3376,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3390,N_3391,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3431,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3447,N_3448,N_3450,N_3451,N_3452,N_3453,N_3454,N_3457,N_3458,N_3459,N_3462,N_3463,N_3465,N_3468,N_3469,N_3472,N_3473,N_3474,N_3476,N_3477,N_3478,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3499,N_3500,N_3501,N_3502,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3511,N_3512,N_3514,N_3515,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3530,N_3532,N_3534,N_3536,N_3537,N_3538,N_3539,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3548,N_3549,N_3550,N_3551,N_3552,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3580,N_3582,N_3583,N_3584,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3601,N_3602,N_3604,N_3605,N_3607,N_3608,N_3609,N_3610,N_3611,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3627,N_3628,N_3629,N_3630,N_3631,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3643,N_3644,N_3646,N_3647,N_3648,N_3652,N_3653,N_3654,N_3655,N_3656,N_3658,N_3659,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3706,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3717,N_3718,N_3720,N_3721,N_3722,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3732,N_3734,N_3735,N_3736,N_3737,N_3740,N_3741,N_3742,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3758,N_3759,N_3764,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3776,N_3777,N_3779,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3798,N_3799,N_3800,N_3801,N_3802,N_3804,N_3805,N_3806,N_3808,N_3809,N_3810,N_3811,N_3813,N_3814,N_3816,N_3817,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3846,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3867,N_3868,N_3869,N_3871,N_3872,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3896,N_3897,N_3898,N_3899,N_3901,N_3902,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3914,N_3916,N_3917,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3946,N_3947,N_3948,N_3950,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3963,N_3964,N_3966,N_3967,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3982,N_3983,N_3984,N_3985,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4010,N_4011,N_4012,N_4013,N_4014,N_4017,N_4018,N_4019,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4038,N_4039,N_4040,N_4041,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4058,N_4059,N_4060,N_4061,N_4063,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4074,N_4075,N_4076,N_4077,N_4079,N_4080,N_4082,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4101,N_4103,N_4105,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4115,N_4117,N_4118,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4131,N_4132,N_4133,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4175,N_4176,N_4177,N_4178,N_4179,N_4181,N_4182,N_4183,N_4184,N_4185,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4202,N_4203,N_4204,N_4205,N_4207,N_4208,N_4210,N_4211,N_4212,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4249,N_4250,N_4254,N_4255,N_4257,N_4259,N_4261,N_4262,N_4264,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4300,N_4301,N_4302,N_4303,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4322,N_4323,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4341,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4352,N_4355,N_4356,N_4357,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4376,N_4377,N_4378,N_4379,N_4380,N_4382,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4403,N_4404,N_4407,N_4408,N_4410,N_4411,N_4412,N_4413,N_4415,N_4416,N_4417,N_4418,N_4420,N_4421,N_4422,N_4423,N_4426,N_4427,N_4428,N_4430,N_4431,N_4432,N_4433,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4442,N_4444,N_4445,N_4447,N_4448,N_4449,N_4451,N_4452,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4484,N_4485,N_4487,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4498,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4515,N_4516,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4525,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4535,N_4536,N_4537,N_4538,N_4539,N_4541,N_4542,N_4543,N_4544,N_4546,N_4547,N_4548,N_4549,N_4551,N_4552,N_4553,N_4554,N_4556,N_4557,N_4558,N_4560,N_4562,N_4563,N_4564,N_4568,N_4569,N_4570,N_4571,N_4573,N_4574,N_4575,N_4577,N_4578,N_4581,N_4582,N_4583,N_4584,N_4586,N_4587,N_4588,N_4589,N_4590,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4662,N_4663,N_4664,N_4665,N_4666,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4681,N_4682,N_4683,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4703,N_4704,N_4705,N_4706,N_4707,N_4709,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4730,N_4732,N_4733,N_4734,N_4738,N_4739,N_4741,N_4742,N_4745,N_4746,N_4747,N_4748,N_4750,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4769,N_4770,N_4771,N_4778,N_4780,N_4782,N_4783,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4821,N_4822,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4843,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4859,N_4860,N_4861,N_4862,N_4863,N_4865,N_4866,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4880,N_4881,N_4884,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4909,N_4911,N_4912,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4923,N_4925,N_4926,N_4928,N_4929,N_4930,N_4931,N_4932,N_4934,N_4935,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4959,N_4962,N_4963,N_4965,N_4968,N_4969,N_4971,N_4972,N_4975,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4998,N_4999;
or U0 (N_0,In_189,In_207);
nor U1 (N_1,In_404,In_616);
and U2 (N_2,In_469,In_584);
nand U3 (N_3,In_468,In_261);
nand U4 (N_4,In_515,In_139);
or U5 (N_5,In_561,In_722);
nor U6 (N_6,In_219,In_321);
nand U7 (N_7,In_683,In_618);
or U8 (N_8,In_62,In_319);
nand U9 (N_9,In_113,In_576);
or U10 (N_10,In_500,In_425);
nor U11 (N_11,In_605,In_262);
or U12 (N_12,In_33,In_441);
or U13 (N_13,In_669,In_549);
nand U14 (N_14,In_108,In_484);
nand U15 (N_15,In_744,In_288);
or U16 (N_16,In_512,In_123);
nor U17 (N_17,In_396,In_309);
xnor U18 (N_18,In_638,In_213);
xnor U19 (N_19,In_229,In_349);
nor U20 (N_20,In_294,In_32);
and U21 (N_21,In_25,In_373);
nand U22 (N_22,In_491,In_677);
or U23 (N_23,In_643,In_43);
and U24 (N_24,In_22,In_58);
nand U25 (N_25,In_240,In_444);
nand U26 (N_26,In_271,In_347);
nor U27 (N_27,In_475,In_285);
and U28 (N_28,In_436,In_276);
nor U29 (N_29,In_335,In_486);
and U30 (N_30,In_641,In_171);
nand U31 (N_31,In_450,In_16);
nand U32 (N_32,In_52,In_231);
xnor U33 (N_33,In_367,In_144);
xor U34 (N_34,In_185,In_375);
and U35 (N_35,In_466,In_84);
or U36 (N_36,In_42,In_79);
and U37 (N_37,In_740,In_145);
xnor U38 (N_38,In_173,In_600);
or U39 (N_39,In_354,In_37);
xnor U40 (N_40,In_274,In_483);
xnor U41 (N_41,In_521,In_199);
xor U42 (N_42,In_719,In_27);
or U43 (N_43,In_275,In_615);
nor U44 (N_44,In_608,In_380);
or U45 (N_45,In_745,In_57);
xnor U46 (N_46,In_7,In_534);
xnor U47 (N_47,In_585,In_53);
nor U48 (N_48,In_518,In_730);
nor U49 (N_49,In_104,In_502);
nor U50 (N_50,In_44,In_426);
nand U51 (N_51,In_266,In_673);
nand U52 (N_52,In_405,In_545);
nand U53 (N_53,In_47,In_642);
or U54 (N_54,In_381,In_140);
or U55 (N_55,In_41,In_617);
or U56 (N_56,In_298,In_465);
and U57 (N_57,In_190,In_333);
nand U58 (N_58,In_738,In_519);
or U59 (N_59,In_313,In_726);
or U60 (N_60,In_118,In_350);
nand U61 (N_61,In_149,In_485);
nand U62 (N_62,In_657,In_334);
or U63 (N_63,In_133,In_581);
nand U64 (N_64,In_676,In_270);
xnor U65 (N_65,In_143,In_248);
nor U66 (N_66,In_157,In_451);
nand U67 (N_67,In_329,In_131);
and U68 (N_68,In_324,In_65);
or U69 (N_69,In_12,In_201);
nand U70 (N_70,In_242,In_328);
nand U71 (N_71,In_222,In_645);
nor U72 (N_72,In_660,In_6);
and U73 (N_73,In_714,In_307);
and U74 (N_74,In_682,In_269);
nor U75 (N_75,In_297,In_135);
or U76 (N_76,In_147,In_579);
nand U77 (N_77,In_202,In_359);
and U78 (N_78,In_5,In_568);
and U79 (N_79,In_177,In_564);
nor U80 (N_80,In_402,In_110);
xor U81 (N_81,In_287,In_83);
nor U82 (N_82,In_556,In_458);
or U83 (N_83,In_137,In_453);
and U84 (N_84,In_394,In_280);
xnor U85 (N_85,In_296,In_454);
or U86 (N_86,In_416,In_40);
and U87 (N_87,In_629,In_665);
nor U88 (N_88,In_300,In_371);
xnor U89 (N_89,In_24,In_172);
and U90 (N_90,In_169,In_387);
and U91 (N_91,In_66,In_746);
or U92 (N_92,In_161,In_70);
nor U93 (N_93,In_245,In_395);
or U94 (N_94,In_96,In_675);
and U95 (N_95,In_604,In_538);
nor U96 (N_96,In_279,In_476);
and U97 (N_97,In_655,In_178);
nand U98 (N_98,In_644,In_221);
and U99 (N_99,In_13,In_86);
or U100 (N_100,In_734,In_567);
and U101 (N_101,In_667,In_390);
nor U102 (N_102,In_663,In_166);
xor U103 (N_103,In_739,In_244);
and U104 (N_104,In_136,In_412);
xnor U105 (N_105,In_102,In_666);
and U106 (N_106,In_174,In_376);
xor U107 (N_107,In_107,In_409);
and U108 (N_108,In_293,In_610);
and U109 (N_109,In_434,In_372);
nor U110 (N_110,In_204,In_23);
or U111 (N_111,In_303,In_210);
and U112 (N_112,In_640,In_747);
nand U113 (N_113,In_81,In_685);
nor U114 (N_114,In_536,In_315);
and U115 (N_115,In_115,In_68);
nor U116 (N_116,In_693,In_277);
nor U117 (N_117,In_619,In_708);
nor U118 (N_118,In_181,In_11);
xor U119 (N_119,In_662,In_494);
and U120 (N_120,In_195,In_314);
and U121 (N_121,In_537,In_284);
and U122 (N_122,In_748,In_712);
or U123 (N_123,In_64,In_217);
nor U124 (N_124,In_624,In_716);
nand U125 (N_125,In_393,In_457);
nor U126 (N_126,In_478,In_256);
nor U127 (N_127,In_595,In_493);
and U128 (N_128,In_415,In_48);
nand U129 (N_129,In_659,In_449);
nor U130 (N_130,In_208,In_607);
xnor U131 (N_131,In_92,In_695);
nor U132 (N_132,In_656,In_463);
or U133 (N_133,In_341,In_689);
xnor U134 (N_134,In_743,In_156);
and U135 (N_135,In_382,In_723);
and U136 (N_136,In_499,In_742);
or U137 (N_137,In_191,In_80);
nand U138 (N_138,In_700,In_732);
or U139 (N_139,In_226,In_291);
or U140 (N_140,In_82,In_87);
xor U141 (N_141,In_525,In_715);
and U142 (N_142,In_541,In_370);
xor U143 (N_143,In_330,In_649);
nand U144 (N_144,In_348,In_238);
nor U145 (N_145,In_430,In_482);
and U146 (N_146,In_322,In_472);
nand U147 (N_147,In_109,In_305);
or U148 (N_148,In_433,In_130);
or U149 (N_149,In_255,In_527);
and U150 (N_150,In_148,In_99);
or U151 (N_151,In_127,In_516);
nand U152 (N_152,In_524,In_292);
nor U153 (N_153,In_146,In_510);
nand U154 (N_154,In_481,In_193);
xor U155 (N_155,In_681,In_150);
nand U156 (N_156,In_180,In_498);
nor U157 (N_157,In_327,In_421);
or U158 (N_158,In_264,In_282);
xnor U159 (N_159,In_551,In_1);
nand U160 (N_160,In_223,In_623);
nand U161 (N_161,In_165,In_211);
nor U162 (N_162,In_614,In_508);
or U163 (N_163,In_507,In_386);
xor U164 (N_164,In_557,In_250);
nor U165 (N_165,In_105,In_384);
or U166 (N_166,In_206,In_365);
nor U167 (N_167,In_635,In_205);
nand U168 (N_168,In_186,In_357);
nor U169 (N_169,In_124,In_340);
nor U170 (N_170,In_119,In_184);
nand U171 (N_171,In_111,In_273);
or U172 (N_172,In_2,In_630);
nand U173 (N_173,In_35,In_306);
or U174 (N_174,In_580,In_397);
and U175 (N_175,In_492,In_560);
or U176 (N_176,In_533,In_575);
xnor U177 (N_177,In_325,In_95);
or U178 (N_178,In_749,In_338);
or U179 (N_179,In_632,In_114);
nor U180 (N_180,In_227,In_710);
nor U181 (N_181,In_578,In_661);
or U182 (N_182,In_346,In_69);
nand U183 (N_183,In_310,In_258);
nand U184 (N_184,In_489,In_603);
xor U185 (N_185,In_21,In_59);
and U186 (N_186,In_299,In_162);
nand U187 (N_187,In_429,In_592);
or U188 (N_188,In_265,In_601);
and U189 (N_189,In_364,In_406);
and U190 (N_190,In_511,In_668);
and U191 (N_191,In_593,In_652);
or U192 (N_192,In_729,In_741);
xor U193 (N_193,In_4,In_236);
nand U194 (N_194,In_420,In_63);
or U195 (N_195,In_437,In_132);
nor U196 (N_196,In_56,In_461);
nor U197 (N_197,In_563,In_535);
nor U198 (N_198,In_352,In_696);
nand U199 (N_199,In_553,In_0);
nor U200 (N_200,In_308,In_260);
nand U201 (N_201,In_368,In_398);
and U202 (N_202,In_142,In_170);
or U203 (N_203,In_112,In_344);
xnor U204 (N_204,In_399,In_621);
and U205 (N_205,In_237,In_724);
and U206 (N_206,In_411,In_474);
xor U207 (N_207,In_197,In_163);
nor U208 (N_208,In_257,In_312);
and U209 (N_209,In_428,In_230);
and U210 (N_210,In_501,In_464);
and U211 (N_211,In_116,In_548);
or U212 (N_212,In_323,In_117);
nor U213 (N_213,In_459,In_471);
and U214 (N_214,In_736,In_639);
xor U215 (N_215,In_234,In_636);
xnor U216 (N_216,In_268,In_383);
or U217 (N_217,In_259,In_9);
nor U218 (N_218,In_54,In_414);
nor U219 (N_219,In_517,In_559);
and U220 (N_220,In_456,In_215);
nor U221 (N_221,In_241,In_717);
nand U222 (N_222,In_71,In_462);
nand U223 (N_223,In_495,In_628);
nor U224 (N_224,In_570,In_634);
nor U225 (N_225,In_243,In_597);
or U226 (N_226,In_77,In_562);
and U227 (N_227,In_671,In_153);
nand U228 (N_228,In_467,In_20);
and U229 (N_229,In_74,In_709);
nand U230 (N_230,In_224,In_196);
nor U231 (N_231,In_684,In_573);
or U232 (N_232,In_733,In_546);
or U233 (N_233,In_304,In_154);
or U234 (N_234,In_218,In_417);
nor U235 (N_235,In_680,In_439);
and U236 (N_236,In_403,In_203);
nand U237 (N_237,In_3,In_91);
nand U238 (N_238,In_289,In_342);
and U239 (N_239,In_530,In_674);
xor U240 (N_240,In_89,In_232);
or U241 (N_241,In_361,In_168);
nor U242 (N_242,In_28,In_703);
and U243 (N_243,In_49,In_612);
nor U244 (N_244,In_427,In_721);
nor U245 (N_245,In_249,In_209);
and U246 (N_246,In_141,In_34);
xor U247 (N_247,In_735,In_252);
nand U248 (N_248,In_187,In_392);
nand U249 (N_249,In_8,In_690);
nand U250 (N_250,In_737,In_355);
nand U251 (N_251,In_97,In_692);
xnor U252 (N_252,In_488,In_725);
and U253 (N_253,In_122,In_72);
xnor U254 (N_254,In_331,In_336);
nand U255 (N_255,In_295,In_611);
nor U256 (N_256,In_718,In_424);
xor U257 (N_257,In_251,In_633);
or U258 (N_258,In_46,In_694);
and U259 (N_259,In_631,In_151);
and U260 (N_260,In_45,In_36);
or U261 (N_261,In_159,In_360);
nor U262 (N_262,In_594,In_326);
xor U263 (N_263,In_18,In_620);
or U264 (N_264,In_128,In_701);
xor U265 (N_265,In_212,In_496);
nand U266 (N_266,In_94,In_351);
nor U267 (N_267,In_10,In_532);
and U268 (N_268,In_30,In_129);
and U269 (N_269,In_39,In_650);
and U270 (N_270,In_67,In_528);
or U271 (N_271,In_423,In_379);
nor U272 (N_272,In_599,In_198);
nand U273 (N_273,In_278,In_699);
nor U274 (N_274,In_418,In_26);
nand U275 (N_275,In_552,In_106);
xor U276 (N_276,In_353,In_391);
and U277 (N_277,In_51,In_550);
and U278 (N_278,In_233,In_435);
nand U279 (N_279,In_267,In_60);
and U280 (N_280,In_369,In_448);
or U281 (N_281,In_554,In_73);
nor U282 (N_282,In_686,In_526);
nand U283 (N_283,In_598,In_90);
nand U284 (N_284,In_509,In_571);
and U285 (N_285,In_555,In_558);
nand U286 (N_286,In_179,In_687);
and U287 (N_287,In_506,In_192);
or U288 (N_288,In_75,In_514);
nand U289 (N_289,In_574,In_317);
or U290 (N_290,In_214,In_320);
nand U291 (N_291,In_419,In_164);
or U292 (N_292,In_378,In_125);
nor U293 (N_293,In_477,In_272);
or U294 (N_294,In_126,In_235);
nor U295 (N_295,In_290,In_410);
or U296 (N_296,In_706,In_490);
or U297 (N_297,In_422,In_672);
nand U298 (N_298,In_401,In_679);
xnor U299 (N_299,In_316,In_627);
nor U300 (N_300,In_586,In_100);
and U301 (N_301,In_505,In_589);
nand U302 (N_302,In_566,In_432);
nand U303 (N_303,In_446,In_588);
nor U304 (N_304,In_286,In_670);
or U305 (N_305,In_93,In_407);
and U306 (N_306,In_363,In_720);
nand U307 (N_307,In_622,In_625);
xor U308 (N_308,In_253,In_543);
nor U309 (N_309,In_440,In_470);
or U310 (N_310,In_374,In_200);
nor U311 (N_311,In_487,In_152);
nand U312 (N_312,In_311,In_626);
or U313 (N_313,In_473,In_572);
or U314 (N_314,In_155,In_158);
nand U315 (N_315,In_697,In_332);
or U316 (N_316,In_513,In_76);
or U317 (N_317,In_455,In_61);
xnor U318 (N_318,In_731,In_577);
or U319 (N_319,In_228,In_539);
xor U320 (N_320,In_691,In_590);
nand U321 (N_321,In_160,In_175);
and U322 (N_322,In_318,In_400);
nand U323 (N_323,In_19,In_120);
nand U324 (N_324,In_569,In_583);
and U325 (N_325,In_283,In_188);
xor U326 (N_326,In_176,In_358);
nand U327 (N_327,In_591,In_678);
nand U328 (N_328,In_713,In_648);
nor U329 (N_329,In_688,In_31);
or U330 (N_330,In_587,In_452);
and U331 (N_331,In_98,In_345);
and U332 (N_332,In_651,In_431);
nor U333 (N_333,In_653,In_366);
nand U334 (N_334,In_522,In_389);
and U335 (N_335,In_388,In_443);
xnor U336 (N_336,In_704,In_246);
or U337 (N_337,In_225,In_220);
nand U338 (N_338,In_602,In_194);
or U339 (N_339,In_377,In_503);
nor U340 (N_340,In_606,In_263);
xor U341 (N_341,In_413,In_609);
nand U342 (N_342,In_658,In_216);
nand U343 (N_343,In_582,In_103);
nor U344 (N_344,In_88,In_356);
nand U345 (N_345,In_447,In_167);
nand U346 (N_346,In_239,In_408);
nand U347 (N_347,In_460,In_183);
and U348 (N_348,In_520,In_121);
nand U349 (N_349,In_637,In_301);
and U350 (N_350,In_385,In_711);
xor U351 (N_351,In_337,In_14);
nor U352 (N_352,In_547,In_702);
or U353 (N_353,In_302,In_497);
nor U354 (N_354,In_38,In_698);
xnor U355 (N_355,In_55,In_646);
nor U356 (N_356,In_728,In_479);
or U357 (N_357,In_540,In_445);
nor U358 (N_358,In_15,In_17);
nor U359 (N_359,In_654,In_664);
or U360 (N_360,In_247,In_705);
nor U361 (N_361,In_438,In_138);
nand U362 (N_362,In_254,In_281);
nor U363 (N_363,In_362,In_544);
nand U364 (N_364,In_531,In_29);
nor U365 (N_365,In_78,In_523);
or U366 (N_366,In_50,In_182);
and U367 (N_367,In_442,In_85);
or U368 (N_368,In_504,In_134);
nand U369 (N_369,In_613,In_343);
or U370 (N_370,In_727,In_565);
nand U371 (N_371,In_707,In_101);
nor U372 (N_372,In_529,In_596);
nor U373 (N_373,In_647,In_480);
nor U374 (N_374,In_339,In_542);
and U375 (N_375,In_80,In_723);
nand U376 (N_376,In_205,In_585);
or U377 (N_377,In_217,In_315);
nand U378 (N_378,In_735,In_116);
nand U379 (N_379,In_588,In_743);
nor U380 (N_380,In_256,In_68);
and U381 (N_381,In_16,In_672);
nand U382 (N_382,In_654,In_647);
or U383 (N_383,In_740,In_616);
nor U384 (N_384,In_233,In_627);
or U385 (N_385,In_678,In_544);
nand U386 (N_386,In_494,In_695);
and U387 (N_387,In_448,In_169);
or U388 (N_388,In_524,In_480);
xnor U389 (N_389,In_318,In_202);
nor U390 (N_390,In_440,In_507);
nor U391 (N_391,In_247,In_206);
or U392 (N_392,In_444,In_107);
or U393 (N_393,In_105,In_579);
nor U394 (N_394,In_513,In_118);
nand U395 (N_395,In_628,In_600);
or U396 (N_396,In_590,In_95);
and U397 (N_397,In_378,In_387);
xnor U398 (N_398,In_621,In_432);
nand U399 (N_399,In_575,In_105);
nor U400 (N_400,In_172,In_282);
and U401 (N_401,In_78,In_143);
and U402 (N_402,In_264,In_16);
xnor U403 (N_403,In_253,In_715);
or U404 (N_404,In_228,In_555);
and U405 (N_405,In_509,In_399);
nor U406 (N_406,In_444,In_635);
or U407 (N_407,In_584,In_306);
or U408 (N_408,In_502,In_418);
or U409 (N_409,In_359,In_351);
nand U410 (N_410,In_194,In_221);
xnor U411 (N_411,In_119,In_24);
and U412 (N_412,In_102,In_186);
nor U413 (N_413,In_229,In_65);
nor U414 (N_414,In_374,In_160);
xor U415 (N_415,In_413,In_256);
and U416 (N_416,In_161,In_50);
nor U417 (N_417,In_746,In_378);
nand U418 (N_418,In_226,In_79);
and U419 (N_419,In_533,In_680);
and U420 (N_420,In_595,In_248);
nor U421 (N_421,In_271,In_69);
and U422 (N_422,In_714,In_388);
nor U423 (N_423,In_318,In_558);
nand U424 (N_424,In_260,In_706);
nor U425 (N_425,In_480,In_304);
or U426 (N_426,In_301,In_529);
nor U427 (N_427,In_562,In_32);
or U428 (N_428,In_722,In_636);
and U429 (N_429,In_75,In_73);
and U430 (N_430,In_166,In_412);
or U431 (N_431,In_65,In_115);
and U432 (N_432,In_595,In_126);
or U433 (N_433,In_63,In_517);
or U434 (N_434,In_574,In_474);
nand U435 (N_435,In_132,In_293);
and U436 (N_436,In_410,In_748);
or U437 (N_437,In_674,In_245);
nor U438 (N_438,In_91,In_514);
or U439 (N_439,In_182,In_384);
and U440 (N_440,In_298,In_49);
nand U441 (N_441,In_323,In_245);
or U442 (N_442,In_571,In_9);
or U443 (N_443,In_409,In_417);
or U444 (N_444,In_604,In_133);
or U445 (N_445,In_418,In_244);
or U446 (N_446,In_675,In_442);
nand U447 (N_447,In_14,In_710);
nand U448 (N_448,In_669,In_602);
and U449 (N_449,In_21,In_346);
or U450 (N_450,In_6,In_335);
nand U451 (N_451,In_597,In_45);
and U452 (N_452,In_80,In_23);
or U453 (N_453,In_348,In_241);
or U454 (N_454,In_346,In_569);
or U455 (N_455,In_68,In_241);
and U456 (N_456,In_672,In_615);
or U457 (N_457,In_371,In_123);
nand U458 (N_458,In_557,In_538);
nand U459 (N_459,In_206,In_39);
nand U460 (N_460,In_664,In_363);
nor U461 (N_461,In_577,In_186);
and U462 (N_462,In_267,In_381);
and U463 (N_463,In_120,In_616);
and U464 (N_464,In_529,In_425);
nor U465 (N_465,In_141,In_700);
and U466 (N_466,In_687,In_700);
and U467 (N_467,In_578,In_616);
and U468 (N_468,In_341,In_498);
or U469 (N_469,In_510,In_675);
and U470 (N_470,In_104,In_647);
and U471 (N_471,In_741,In_124);
and U472 (N_472,In_640,In_100);
nand U473 (N_473,In_621,In_420);
nand U474 (N_474,In_719,In_154);
xor U475 (N_475,In_234,In_684);
or U476 (N_476,In_594,In_661);
xnor U477 (N_477,In_531,In_711);
nand U478 (N_478,In_591,In_612);
and U479 (N_479,In_683,In_169);
nor U480 (N_480,In_590,In_196);
nand U481 (N_481,In_313,In_590);
and U482 (N_482,In_498,In_29);
and U483 (N_483,In_198,In_596);
and U484 (N_484,In_565,In_306);
nor U485 (N_485,In_281,In_524);
nand U486 (N_486,In_193,In_59);
or U487 (N_487,In_111,In_240);
xnor U488 (N_488,In_234,In_567);
nor U489 (N_489,In_606,In_472);
xnor U490 (N_490,In_688,In_59);
or U491 (N_491,In_582,In_113);
and U492 (N_492,In_362,In_243);
xor U493 (N_493,In_487,In_25);
nand U494 (N_494,In_579,In_205);
or U495 (N_495,In_240,In_351);
nand U496 (N_496,In_686,In_593);
xor U497 (N_497,In_435,In_349);
or U498 (N_498,In_324,In_529);
nand U499 (N_499,In_23,In_410);
xnor U500 (N_500,In_686,In_612);
nor U501 (N_501,In_648,In_440);
nor U502 (N_502,In_430,In_553);
xnor U503 (N_503,In_646,In_59);
xnor U504 (N_504,In_23,In_424);
nor U505 (N_505,In_553,In_297);
nor U506 (N_506,In_591,In_72);
xor U507 (N_507,In_607,In_537);
xor U508 (N_508,In_490,In_261);
nor U509 (N_509,In_340,In_200);
xnor U510 (N_510,In_253,In_460);
or U511 (N_511,In_207,In_727);
nor U512 (N_512,In_535,In_282);
or U513 (N_513,In_554,In_206);
and U514 (N_514,In_570,In_255);
or U515 (N_515,In_291,In_181);
nand U516 (N_516,In_612,In_589);
nor U517 (N_517,In_383,In_590);
nor U518 (N_518,In_297,In_698);
or U519 (N_519,In_311,In_112);
and U520 (N_520,In_315,In_328);
or U521 (N_521,In_556,In_282);
and U522 (N_522,In_594,In_180);
nand U523 (N_523,In_555,In_346);
nand U524 (N_524,In_611,In_686);
xor U525 (N_525,In_535,In_65);
xor U526 (N_526,In_43,In_79);
and U527 (N_527,In_698,In_702);
or U528 (N_528,In_236,In_737);
or U529 (N_529,In_544,In_589);
nor U530 (N_530,In_293,In_383);
and U531 (N_531,In_606,In_391);
or U532 (N_532,In_205,In_514);
nand U533 (N_533,In_263,In_79);
xor U534 (N_534,In_186,In_645);
and U535 (N_535,In_605,In_395);
and U536 (N_536,In_102,In_644);
nand U537 (N_537,In_169,In_287);
nand U538 (N_538,In_195,In_163);
nor U539 (N_539,In_202,In_209);
nor U540 (N_540,In_477,In_341);
nor U541 (N_541,In_487,In_522);
nor U542 (N_542,In_1,In_603);
or U543 (N_543,In_304,In_342);
nand U544 (N_544,In_526,In_354);
nor U545 (N_545,In_153,In_466);
or U546 (N_546,In_302,In_540);
or U547 (N_547,In_12,In_596);
nor U548 (N_548,In_121,In_629);
and U549 (N_549,In_391,In_514);
and U550 (N_550,In_617,In_404);
nand U551 (N_551,In_511,In_223);
nor U552 (N_552,In_8,In_748);
or U553 (N_553,In_495,In_366);
nor U554 (N_554,In_261,In_677);
or U555 (N_555,In_643,In_503);
xnor U556 (N_556,In_378,In_266);
nand U557 (N_557,In_22,In_286);
or U558 (N_558,In_736,In_70);
and U559 (N_559,In_178,In_689);
nor U560 (N_560,In_730,In_585);
xnor U561 (N_561,In_128,In_495);
and U562 (N_562,In_338,In_721);
or U563 (N_563,In_216,In_619);
nor U564 (N_564,In_611,In_522);
nand U565 (N_565,In_159,In_195);
nor U566 (N_566,In_680,In_391);
or U567 (N_567,In_301,In_11);
and U568 (N_568,In_579,In_488);
xnor U569 (N_569,In_159,In_336);
nor U570 (N_570,In_203,In_545);
nor U571 (N_571,In_460,In_404);
and U572 (N_572,In_217,In_49);
or U573 (N_573,In_548,In_738);
or U574 (N_574,In_569,In_348);
and U575 (N_575,In_213,In_611);
and U576 (N_576,In_4,In_627);
nand U577 (N_577,In_518,In_3);
nand U578 (N_578,In_13,In_321);
nand U579 (N_579,In_686,In_292);
and U580 (N_580,In_507,In_697);
xnor U581 (N_581,In_734,In_389);
and U582 (N_582,In_452,In_504);
and U583 (N_583,In_37,In_562);
or U584 (N_584,In_290,In_65);
and U585 (N_585,In_478,In_468);
nand U586 (N_586,In_140,In_577);
nand U587 (N_587,In_34,In_306);
or U588 (N_588,In_740,In_336);
xnor U589 (N_589,In_326,In_354);
and U590 (N_590,In_64,In_74);
xnor U591 (N_591,In_567,In_520);
or U592 (N_592,In_130,In_412);
xnor U593 (N_593,In_611,In_389);
nor U594 (N_594,In_248,In_572);
nand U595 (N_595,In_206,In_255);
nand U596 (N_596,In_588,In_323);
and U597 (N_597,In_690,In_726);
and U598 (N_598,In_564,In_299);
nor U599 (N_599,In_348,In_304);
or U600 (N_600,In_492,In_694);
and U601 (N_601,In_147,In_243);
or U602 (N_602,In_149,In_326);
or U603 (N_603,In_188,In_24);
nor U604 (N_604,In_535,In_226);
nand U605 (N_605,In_214,In_197);
or U606 (N_606,In_219,In_494);
nand U607 (N_607,In_366,In_625);
and U608 (N_608,In_317,In_204);
and U609 (N_609,In_200,In_134);
nand U610 (N_610,In_191,In_89);
nand U611 (N_611,In_412,In_479);
and U612 (N_612,In_129,In_540);
nand U613 (N_613,In_337,In_673);
nand U614 (N_614,In_591,In_297);
nand U615 (N_615,In_574,In_571);
nand U616 (N_616,In_521,In_117);
and U617 (N_617,In_207,In_525);
nand U618 (N_618,In_16,In_149);
nor U619 (N_619,In_134,In_144);
and U620 (N_620,In_119,In_172);
nor U621 (N_621,In_357,In_628);
or U622 (N_622,In_432,In_638);
xor U623 (N_623,In_650,In_176);
nor U624 (N_624,In_721,In_158);
and U625 (N_625,In_490,In_362);
and U626 (N_626,In_552,In_226);
xnor U627 (N_627,In_184,In_125);
and U628 (N_628,In_0,In_147);
and U629 (N_629,In_315,In_465);
or U630 (N_630,In_502,In_507);
nor U631 (N_631,In_667,In_183);
and U632 (N_632,In_39,In_230);
or U633 (N_633,In_19,In_589);
nand U634 (N_634,In_345,In_393);
nand U635 (N_635,In_360,In_710);
nand U636 (N_636,In_685,In_607);
xor U637 (N_637,In_292,In_489);
nand U638 (N_638,In_642,In_279);
nand U639 (N_639,In_576,In_505);
nor U640 (N_640,In_267,In_697);
xnor U641 (N_641,In_521,In_469);
or U642 (N_642,In_311,In_531);
and U643 (N_643,In_158,In_466);
or U644 (N_644,In_82,In_505);
nor U645 (N_645,In_219,In_27);
nor U646 (N_646,In_714,In_639);
nand U647 (N_647,In_456,In_327);
nand U648 (N_648,In_628,In_577);
or U649 (N_649,In_489,In_458);
nand U650 (N_650,In_701,In_193);
nor U651 (N_651,In_299,In_710);
nand U652 (N_652,In_580,In_706);
nor U653 (N_653,In_133,In_565);
nor U654 (N_654,In_440,In_289);
nor U655 (N_655,In_254,In_393);
nand U656 (N_656,In_728,In_558);
or U657 (N_657,In_137,In_22);
or U658 (N_658,In_210,In_325);
nand U659 (N_659,In_553,In_335);
nand U660 (N_660,In_343,In_191);
nor U661 (N_661,In_94,In_380);
or U662 (N_662,In_285,In_382);
nor U663 (N_663,In_45,In_423);
or U664 (N_664,In_715,In_84);
nor U665 (N_665,In_544,In_721);
or U666 (N_666,In_78,In_610);
nor U667 (N_667,In_173,In_105);
or U668 (N_668,In_198,In_420);
xnor U669 (N_669,In_371,In_118);
nor U670 (N_670,In_624,In_93);
xor U671 (N_671,In_27,In_148);
xor U672 (N_672,In_222,In_658);
nand U673 (N_673,In_532,In_26);
or U674 (N_674,In_586,In_368);
and U675 (N_675,In_657,In_228);
nor U676 (N_676,In_287,In_649);
or U677 (N_677,In_657,In_427);
nor U678 (N_678,In_418,In_35);
nand U679 (N_679,In_689,In_575);
and U680 (N_680,In_485,In_565);
xnor U681 (N_681,In_302,In_89);
nand U682 (N_682,In_439,In_73);
nor U683 (N_683,In_29,In_38);
and U684 (N_684,In_622,In_344);
nor U685 (N_685,In_372,In_441);
nand U686 (N_686,In_179,In_310);
and U687 (N_687,In_232,In_497);
nand U688 (N_688,In_354,In_703);
nand U689 (N_689,In_154,In_688);
xnor U690 (N_690,In_685,In_229);
nand U691 (N_691,In_524,In_301);
or U692 (N_692,In_579,In_338);
or U693 (N_693,In_676,In_22);
xnor U694 (N_694,In_63,In_362);
nand U695 (N_695,In_97,In_544);
xnor U696 (N_696,In_625,In_162);
or U697 (N_697,In_199,In_194);
nor U698 (N_698,In_637,In_320);
xor U699 (N_699,In_376,In_686);
or U700 (N_700,In_406,In_367);
or U701 (N_701,In_400,In_85);
nand U702 (N_702,In_153,In_379);
and U703 (N_703,In_300,In_174);
nand U704 (N_704,In_92,In_51);
nor U705 (N_705,In_104,In_650);
nand U706 (N_706,In_409,In_126);
or U707 (N_707,In_647,In_227);
nand U708 (N_708,In_348,In_7);
nand U709 (N_709,In_685,In_261);
nand U710 (N_710,In_693,In_587);
and U711 (N_711,In_395,In_477);
nor U712 (N_712,In_582,In_57);
or U713 (N_713,In_156,In_705);
and U714 (N_714,In_72,In_336);
and U715 (N_715,In_50,In_694);
and U716 (N_716,In_8,In_40);
or U717 (N_717,In_487,In_440);
or U718 (N_718,In_16,In_210);
xnor U719 (N_719,In_420,In_53);
nor U720 (N_720,In_552,In_155);
nor U721 (N_721,In_329,In_390);
nor U722 (N_722,In_667,In_454);
nor U723 (N_723,In_381,In_150);
and U724 (N_724,In_489,In_209);
nor U725 (N_725,In_743,In_63);
nand U726 (N_726,In_116,In_450);
or U727 (N_727,In_395,In_727);
or U728 (N_728,In_654,In_514);
nand U729 (N_729,In_545,In_465);
nand U730 (N_730,In_236,In_640);
nor U731 (N_731,In_161,In_244);
or U732 (N_732,In_293,In_207);
nand U733 (N_733,In_513,In_589);
or U734 (N_734,In_548,In_465);
nand U735 (N_735,In_711,In_656);
and U736 (N_736,In_346,In_609);
or U737 (N_737,In_743,In_549);
and U738 (N_738,In_419,In_687);
xor U739 (N_739,In_339,In_739);
and U740 (N_740,In_492,In_621);
nor U741 (N_741,In_440,In_355);
nor U742 (N_742,In_717,In_667);
nor U743 (N_743,In_368,In_655);
nor U744 (N_744,In_370,In_256);
or U745 (N_745,In_18,In_222);
nand U746 (N_746,In_6,In_710);
nor U747 (N_747,In_45,In_477);
nand U748 (N_748,In_526,In_666);
xor U749 (N_749,In_234,In_173);
nor U750 (N_750,In_492,In_10);
or U751 (N_751,In_651,In_654);
or U752 (N_752,In_71,In_192);
nor U753 (N_753,In_614,In_275);
nand U754 (N_754,In_713,In_172);
xnor U755 (N_755,In_417,In_558);
or U756 (N_756,In_331,In_152);
or U757 (N_757,In_563,In_616);
or U758 (N_758,In_513,In_423);
nand U759 (N_759,In_324,In_443);
or U760 (N_760,In_482,In_527);
and U761 (N_761,In_356,In_623);
nor U762 (N_762,In_418,In_440);
xor U763 (N_763,In_402,In_132);
nand U764 (N_764,In_522,In_434);
or U765 (N_765,In_226,In_585);
nand U766 (N_766,In_126,In_573);
nor U767 (N_767,In_518,In_713);
xor U768 (N_768,In_329,In_629);
and U769 (N_769,In_341,In_674);
nor U770 (N_770,In_360,In_522);
nand U771 (N_771,In_387,In_302);
and U772 (N_772,In_287,In_377);
nor U773 (N_773,In_619,In_350);
xnor U774 (N_774,In_74,In_582);
xor U775 (N_775,In_302,In_269);
xor U776 (N_776,In_449,In_230);
nor U777 (N_777,In_712,In_732);
nand U778 (N_778,In_121,In_391);
xor U779 (N_779,In_653,In_516);
and U780 (N_780,In_657,In_534);
or U781 (N_781,In_255,In_482);
nand U782 (N_782,In_566,In_567);
and U783 (N_783,In_91,In_435);
nor U784 (N_784,In_454,In_201);
nor U785 (N_785,In_13,In_289);
nor U786 (N_786,In_352,In_300);
and U787 (N_787,In_425,In_435);
nor U788 (N_788,In_51,In_192);
nand U789 (N_789,In_662,In_577);
or U790 (N_790,In_664,In_482);
and U791 (N_791,In_505,In_441);
xnor U792 (N_792,In_111,In_505);
or U793 (N_793,In_484,In_725);
or U794 (N_794,In_211,In_400);
nor U795 (N_795,In_36,In_91);
xnor U796 (N_796,In_475,In_576);
or U797 (N_797,In_747,In_420);
xor U798 (N_798,In_416,In_145);
or U799 (N_799,In_740,In_284);
nor U800 (N_800,In_736,In_40);
and U801 (N_801,In_273,In_581);
nand U802 (N_802,In_489,In_113);
or U803 (N_803,In_289,In_456);
nor U804 (N_804,In_713,In_609);
nor U805 (N_805,In_54,In_178);
xor U806 (N_806,In_302,In_23);
and U807 (N_807,In_457,In_556);
and U808 (N_808,In_704,In_316);
or U809 (N_809,In_423,In_174);
nand U810 (N_810,In_137,In_585);
nor U811 (N_811,In_449,In_139);
nand U812 (N_812,In_254,In_627);
nor U813 (N_813,In_340,In_653);
nor U814 (N_814,In_701,In_319);
xnor U815 (N_815,In_721,In_390);
nor U816 (N_816,In_291,In_494);
and U817 (N_817,In_152,In_650);
or U818 (N_818,In_4,In_21);
nor U819 (N_819,In_324,In_430);
nor U820 (N_820,In_349,In_562);
nand U821 (N_821,In_525,In_620);
and U822 (N_822,In_231,In_301);
and U823 (N_823,In_587,In_447);
or U824 (N_824,In_616,In_80);
nor U825 (N_825,In_201,In_145);
nor U826 (N_826,In_16,In_152);
or U827 (N_827,In_303,In_28);
nand U828 (N_828,In_441,In_49);
or U829 (N_829,In_670,In_487);
nand U830 (N_830,In_730,In_313);
nand U831 (N_831,In_536,In_541);
or U832 (N_832,In_723,In_187);
and U833 (N_833,In_731,In_228);
and U834 (N_834,In_614,In_365);
or U835 (N_835,In_146,In_218);
xor U836 (N_836,In_17,In_443);
nand U837 (N_837,In_63,In_243);
nand U838 (N_838,In_472,In_139);
and U839 (N_839,In_24,In_32);
xor U840 (N_840,In_305,In_18);
xor U841 (N_841,In_523,In_711);
nand U842 (N_842,In_199,In_16);
or U843 (N_843,In_421,In_483);
nor U844 (N_844,In_502,In_598);
nand U845 (N_845,In_682,In_307);
nand U846 (N_846,In_315,In_162);
or U847 (N_847,In_144,In_108);
nand U848 (N_848,In_542,In_86);
xnor U849 (N_849,In_332,In_97);
nor U850 (N_850,In_481,In_440);
and U851 (N_851,In_378,In_228);
nand U852 (N_852,In_76,In_325);
or U853 (N_853,In_413,In_318);
nand U854 (N_854,In_360,In_337);
nor U855 (N_855,In_49,In_588);
nand U856 (N_856,In_695,In_129);
nand U857 (N_857,In_201,In_621);
and U858 (N_858,In_224,In_517);
and U859 (N_859,In_444,In_10);
nand U860 (N_860,In_461,In_393);
or U861 (N_861,In_124,In_195);
or U862 (N_862,In_237,In_439);
nor U863 (N_863,In_25,In_113);
nor U864 (N_864,In_146,In_570);
nor U865 (N_865,In_533,In_550);
and U866 (N_866,In_694,In_195);
nand U867 (N_867,In_64,In_363);
or U868 (N_868,In_405,In_710);
nand U869 (N_869,In_619,In_461);
nor U870 (N_870,In_655,In_494);
and U871 (N_871,In_489,In_284);
xnor U872 (N_872,In_348,In_592);
nor U873 (N_873,In_231,In_74);
nor U874 (N_874,In_715,In_536);
and U875 (N_875,In_675,In_290);
or U876 (N_876,In_272,In_144);
nor U877 (N_877,In_570,In_42);
nand U878 (N_878,In_681,In_734);
nand U879 (N_879,In_17,In_402);
and U880 (N_880,In_383,In_182);
and U881 (N_881,In_594,In_221);
and U882 (N_882,In_734,In_316);
nor U883 (N_883,In_227,In_368);
or U884 (N_884,In_664,In_76);
nand U885 (N_885,In_227,In_64);
or U886 (N_886,In_431,In_406);
or U887 (N_887,In_114,In_540);
xor U888 (N_888,In_251,In_3);
or U889 (N_889,In_221,In_274);
nor U890 (N_890,In_441,In_706);
or U891 (N_891,In_8,In_611);
or U892 (N_892,In_730,In_447);
xor U893 (N_893,In_237,In_584);
nor U894 (N_894,In_740,In_330);
or U895 (N_895,In_398,In_643);
and U896 (N_896,In_223,In_429);
or U897 (N_897,In_513,In_109);
xor U898 (N_898,In_553,In_462);
nor U899 (N_899,In_737,In_177);
nor U900 (N_900,In_428,In_635);
xor U901 (N_901,In_286,In_735);
or U902 (N_902,In_393,In_228);
nor U903 (N_903,In_122,In_391);
nor U904 (N_904,In_291,In_719);
and U905 (N_905,In_192,In_186);
nor U906 (N_906,In_653,In_379);
xor U907 (N_907,In_665,In_734);
nor U908 (N_908,In_165,In_696);
and U909 (N_909,In_30,In_208);
nor U910 (N_910,In_134,In_549);
nand U911 (N_911,In_555,In_443);
xor U912 (N_912,In_326,In_603);
or U913 (N_913,In_540,In_537);
nand U914 (N_914,In_143,In_228);
or U915 (N_915,In_161,In_313);
nand U916 (N_916,In_1,In_218);
nor U917 (N_917,In_699,In_234);
nand U918 (N_918,In_65,In_192);
nor U919 (N_919,In_675,In_375);
and U920 (N_920,In_283,In_209);
and U921 (N_921,In_650,In_100);
nand U922 (N_922,In_319,In_181);
or U923 (N_923,In_433,In_711);
and U924 (N_924,In_323,In_30);
nor U925 (N_925,In_175,In_600);
or U926 (N_926,In_515,In_57);
nand U927 (N_927,In_362,In_749);
and U928 (N_928,In_206,In_585);
and U929 (N_929,In_336,In_621);
or U930 (N_930,In_89,In_672);
nand U931 (N_931,In_640,In_299);
or U932 (N_932,In_234,In_15);
and U933 (N_933,In_587,In_197);
and U934 (N_934,In_592,In_717);
and U935 (N_935,In_349,In_548);
nand U936 (N_936,In_327,In_432);
or U937 (N_937,In_665,In_46);
nand U938 (N_938,In_145,In_163);
and U939 (N_939,In_75,In_3);
nand U940 (N_940,In_708,In_203);
or U941 (N_941,In_80,In_223);
nand U942 (N_942,In_706,In_475);
nor U943 (N_943,In_357,In_263);
nor U944 (N_944,In_43,In_33);
or U945 (N_945,In_480,In_517);
and U946 (N_946,In_734,In_84);
and U947 (N_947,In_304,In_502);
xor U948 (N_948,In_20,In_173);
and U949 (N_949,In_224,In_413);
nor U950 (N_950,In_288,In_711);
nor U951 (N_951,In_276,In_569);
and U952 (N_952,In_90,In_737);
or U953 (N_953,In_155,In_68);
xnor U954 (N_954,In_251,In_200);
or U955 (N_955,In_249,In_522);
and U956 (N_956,In_443,In_309);
nand U957 (N_957,In_611,In_575);
nand U958 (N_958,In_175,In_162);
nor U959 (N_959,In_609,In_113);
nor U960 (N_960,In_420,In_299);
nor U961 (N_961,In_269,In_225);
nor U962 (N_962,In_277,In_181);
nor U963 (N_963,In_153,In_692);
nand U964 (N_964,In_95,In_532);
nand U965 (N_965,In_496,In_523);
xnor U966 (N_966,In_36,In_669);
and U967 (N_967,In_389,In_448);
xnor U968 (N_968,In_74,In_502);
nor U969 (N_969,In_217,In_348);
nand U970 (N_970,In_218,In_651);
nand U971 (N_971,In_68,In_744);
nor U972 (N_972,In_119,In_441);
nor U973 (N_973,In_450,In_89);
nand U974 (N_974,In_213,In_572);
or U975 (N_975,In_64,In_591);
nand U976 (N_976,In_408,In_327);
and U977 (N_977,In_117,In_295);
nor U978 (N_978,In_195,In_167);
nor U979 (N_979,In_716,In_18);
xnor U980 (N_980,In_484,In_516);
nor U981 (N_981,In_696,In_637);
xor U982 (N_982,In_172,In_377);
and U983 (N_983,In_219,In_507);
and U984 (N_984,In_356,In_497);
and U985 (N_985,In_716,In_119);
nor U986 (N_986,In_681,In_11);
or U987 (N_987,In_532,In_370);
nor U988 (N_988,In_551,In_353);
nand U989 (N_989,In_558,In_265);
or U990 (N_990,In_105,In_83);
or U991 (N_991,In_280,In_46);
nand U992 (N_992,In_569,In_724);
xor U993 (N_993,In_204,In_243);
or U994 (N_994,In_524,In_52);
and U995 (N_995,In_165,In_588);
and U996 (N_996,In_728,In_106);
and U997 (N_997,In_80,In_214);
or U998 (N_998,In_168,In_549);
or U999 (N_999,In_184,In_545);
nand U1000 (N_1000,In_648,In_730);
or U1001 (N_1001,In_574,In_197);
xor U1002 (N_1002,In_243,In_65);
or U1003 (N_1003,In_610,In_265);
or U1004 (N_1004,In_573,In_471);
and U1005 (N_1005,In_55,In_542);
nand U1006 (N_1006,In_397,In_398);
nor U1007 (N_1007,In_217,In_325);
nor U1008 (N_1008,In_181,In_372);
nand U1009 (N_1009,In_381,In_262);
and U1010 (N_1010,In_137,In_632);
nand U1011 (N_1011,In_494,In_217);
nor U1012 (N_1012,In_205,In_554);
or U1013 (N_1013,In_168,In_14);
nand U1014 (N_1014,In_323,In_551);
and U1015 (N_1015,In_551,In_227);
or U1016 (N_1016,In_162,In_96);
and U1017 (N_1017,In_552,In_379);
and U1018 (N_1018,In_426,In_292);
nand U1019 (N_1019,In_235,In_169);
and U1020 (N_1020,In_0,In_7);
nand U1021 (N_1021,In_94,In_602);
or U1022 (N_1022,In_230,In_277);
nand U1023 (N_1023,In_233,In_497);
or U1024 (N_1024,In_691,In_276);
xnor U1025 (N_1025,In_227,In_150);
or U1026 (N_1026,In_250,In_210);
nor U1027 (N_1027,In_252,In_519);
or U1028 (N_1028,In_667,In_590);
xor U1029 (N_1029,In_82,In_617);
or U1030 (N_1030,In_488,In_371);
xor U1031 (N_1031,In_323,In_543);
nor U1032 (N_1032,In_487,In_142);
and U1033 (N_1033,In_150,In_127);
nor U1034 (N_1034,In_207,In_541);
and U1035 (N_1035,In_177,In_406);
and U1036 (N_1036,In_147,In_743);
nand U1037 (N_1037,In_290,In_710);
and U1038 (N_1038,In_33,In_240);
and U1039 (N_1039,In_140,In_330);
or U1040 (N_1040,In_37,In_165);
nor U1041 (N_1041,In_382,In_384);
nor U1042 (N_1042,In_410,In_274);
nor U1043 (N_1043,In_725,In_509);
nand U1044 (N_1044,In_12,In_300);
nor U1045 (N_1045,In_148,In_137);
and U1046 (N_1046,In_488,In_146);
and U1047 (N_1047,In_375,In_171);
nand U1048 (N_1048,In_737,In_123);
and U1049 (N_1049,In_130,In_103);
or U1050 (N_1050,In_33,In_71);
nor U1051 (N_1051,In_557,In_616);
and U1052 (N_1052,In_454,In_589);
or U1053 (N_1053,In_64,In_634);
and U1054 (N_1054,In_78,In_651);
or U1055 (N_1055,In_233,In_727);
and U1056 (N_1056,In_448,In_710);
and U1057 (N_1057,In_408,In_494);
and U1058 (N_1058,In_247,In_238);
nand U1059 (N_1059,In_320,In_617);
nand U1060 (N_1060,In_218,In_77);
and U1061 (N_1061,In_173,In_61);
or U1062 (N_1062,In_16,In_87);
xor U1063 (N_1063,In_544,In_529);
and U1064 (N_1064,In_433,In_617);
and U1065 (N_1065,In_78,In_342);
nand U1066 (N_1066,In_338,In_278);
and U1067 (N_1067,In_568,In_467);
nand U1068 (N_1068,In_373,In_618);
nand U1069 (N_1069,In_604,In_493);
xor U1070 (N_1070,In_404,In_73);
xor U1071 (N_1071,In_164,In_167);
xnor U1072 (N_1072,In_252,In_595);
or U1073 (N_1073,In_625,In_485);
or U1074 (N_1074,In_644,In_243);
and U1075 (N_1075,In_631,In_370);
or U1076 (N_1076,In_561,In_205);
nand U1077 (N_1077,In_198,In_720);
nor U1078 (N_1078,In_323,In_301);
and U1079 (N_1079,In_306,In_415);
nor U1080 (N_1080,In_270,In_152);
nand U1081 (N_1081,In_698,In_525);
nand U1082 (N_1082,In_432,In_143);
nor U1083 (N_1083,In_242,In_582);
or U1084 (N_1084,In_656,In_193);
nand U1085 (N_1085,In_319,In_43);
xnor U1086 (N_1086,In_708,In_497);
nor U1087 (N_1087,In_76,In_523);
nor U1088 (N_1088,In_638,In_226);
nand U1089 (N_1089,In_40,In_36);
nor U1090 (N_1090,In_687,In_574);
xnor U1091 (N_1091,In_521,In_411);
or U1092 (N_1092,In_743,In_196);
and U1093 (N_1093,In_229,In_267);
nand U1094 (N_1094,In_256,In_702);
and U1095 (N_1095,In_265,In_576);
or U1096 (N_1096,In_98,In_106);
or U1097 (N_1097,In_113,In_207);
or U1098 (N_1098,In_16,In_482);
xor U1099 (N_1099,In_412,In_348);
nor U1100 (N_1100,In_392,In_530);
or U1101 (N_1101,In_734,In_338);
nand U1102 (N_1102,In_279,In_614);
nor U1103 (N_1103,In_352,In_385);
nand U1104 (N_1104,In_156,In_486);
and U1105 (N_1105,In_729,In_210);
xnor U1106 (N_1106,In_660,In_375);
and U1107 (N_1107,In_709,In_137);
nor U1108 (N_1108,In_138,In_131);
nand U1109 (N_1109,In_508,In_682);
nor U1110 (N_1110,In_39,In_264);
nand U1111 (N_1111,In_645,In_631);
nand U1112 (N_1112,In_520,In_570);
nand U1113 (N_1113,In_598,In_703);
nand U1114 (N_1114,In_116,In_335);
nor U1115 (N_1115,In_650,In_105);
nand U1116 (N_1116,In_60,In_726);
nand U1117 (N_1117,In_448,In_167);
nor U1118 (N_1118,In_669,In_640);
or U1119 (N_1119,In_64,In_721);
nor U1120 (N_1120,In_38,In_466);
nand U1121 (N_1121,In_52,In_199);
nor U1122 (N_1122,In_102,In_396);
or U1123 (N_1123,In_707,In_149);
nand U1124 (N_1124,In_8,In_601);
nor U1125 (N_1125,In_575,In_437);
nand U1126 (N_1126,In_195,In_261);
or U1127 (N_1127,In_272,In_380);
nor U1128 (N_1128,In_459,In_368);
or U1129 (N_1129,In_427,In_458);
nor U1130 (N_1130,In_273,In_322);
or U1131 (N_1131,In_540,In_642);
or U1132 (N_1132,In_449,In_713);
nand U1133 (N_1133,In_156,In_123);
nor U1134 (N_1134,In_460,In_495);
nor U1135 (N_1135,In_11,In_620);
and U1136 (N_1136,In_207,In_549);
nand U1137 (N_1137,In_103,In_196);
and U1138 (N_1138,In_324,In_242);
and U1139 (N_1139,In_143,In_333);
xnor U1140 (N_1140,In_567,In_596);
nand U1141 (N_1141,In_315,In_653);
or U1142 (N_1142,In_549,In_511);
nor U1143 (N_1143,In_194,In_25);
nand U1144 (N_1144,In_8,In_495);
nand U1145 (N_1145,In_59,In_33);
nor U1146 (N_1146,In_28,In_146);
nor U1147 (N_1147,In_301,In_72);
or U1148 (N_1148,In_140,In_523);
or U1149 (N_1149,In_416,In_400);
nor U1150 (N_1150,In_567,In_662);
nand U1151 (N_1151,In_616,In_570);
nand U1152 (N_1152,In_396,In_478);
nor U1153 (N_1153,In_669,In_618);
and U1154 (N_1154,In_480,In_649);
nand U1155 (N_1155,In_205,In_34);
or U1156 (N_1156,In_582,In_210);
nand U1157 (N_1157,In_474,In_185);
nor U1158 (N_1158,In_0,In_86);
nor U1159 (N_1159,In_736,In_47);
and U1160 (N_1160,In_707,In_160);
nor U1161 (N_1161,In_600,In_107);
and U1162 (N_1162,In_41,In_400);
nor U1163 (N_1163,In_480,In_562);
nor U1164 (N_1164,In_617,In_461);
nand U1165 (N_1165,In_187,In_220);
nor U1166 (N_1166,In_620,In_677);
nand U1167 (N_1167,In_492,In_58);
nor U1168 (N_1168,In_227,In_118);
nand U1169 (N_1169,In_218,In_332);
and U1170 (N_1170,In_586,In_301);
nand U1171 (N_1171,In_125,In_390);
or U1172 (N_1172,In_39,In_24);
or U1173 (N_1173,In_77,In_243);
nand U1174 (N_1174,In_241,In_552);
xor U1175 (N_1175,In_622,In_146);
and U1176 (N_1176,In_364,In_380);
nor U1177 (N_1177,In_265,In_706);
nand U1178 (N_1178,In_246,In_339);
and U1179 (N_1179,In_681,In_564);
nor U1180 (N_1180,In_23,In_413);
or U1181 (N_1181,In_324,In_132);
nand U1182 (N_1182,In_616,In_287);
and U1183 (N_1183,In_343,In_335);
nand U1184 (N_1184,In_739,In_392);
and U1185 (N_1185,In_295,In_42);
nor U1186 (N_1186,In_99,In_24);
nand U1187 (N_1187,In_552,In_232);
nand U1188 (N_1188,In_667,In_662);
or U1189 (N_1189,In_229,In_677);
nand U1190 (N_1190,In_247,In_307);
nand U1191 (N_1191,In_687,In_704);
and U1192 (N_1192,In_320,In_37);
xor U1193 (N_1193,In_555,In_357);
xor U1194 (N_1194,In_622,In_152);
nand U1195 (N_1195,In_132,In_669);
nand U1196 (N_1196,In_255,In_196);
nand U1197 (N_1197,In_585,In_565);
and U1198 (N_1198,In_728,In_422);
nor U1199 (N_1199,In_620,In_425);
nand U1200 (N_1200,In_204,In_218);
nand U1201 (N_1201,In_193,In_655);
and U1202 (N_1202,In_659,In_538);
or U1203 (N_1203,In_106,In_626);
nor U1204 (N_1204,In_540,In_117);
nand U1205 (N_1205,In_233,In_458);
nor U1206 (N_1206,In_698,In_665);
nand U1207 (N_1207,In_57,In_422);
and U1208 (N_1208,In_313,In_659);
or U1209 (N_1209,In_510,In_88);
nand U1210 (N_1210,In_18,In_57);
or U1211 (N_1211,In_223,In_640);
nor U1212 (N_1212,In_32,In_69);
nand U1213 (N_1213,In_324,In_257);
nand U1214 (N_1214,In_304,In_715);
nor U1215 (N_1215,In_552,In_478);
nor U1216 (N_1216,In_328,In_210);
nand U1217 (N_1217,In_705,In_146);
nor U1218 (N_1218,In_100,In_730);
nor U1219 (N_1219,In_202,In_229);
or U1220 (N_1220,In_13,In_652);
nor U1221 (N_1221,In_391,In_362);
and U1222 (N_1222,In_228,In_185);
nor U1223 (N_1223,In_747,In_253);
and U1224 (N_1224,In_729,In_349);
nand U1225 (N_1225,In_201,In_182);
nand U1226 (N_1226,In_521,In_270);
or U1227 (N_1227,In_260,In_145);
nand U1228 (N_1228,In_493,In_669);
nand U1229 (N_1229,In_467,In_102);
nor U1230 (N_1230,In_130,In_181);
nor U1231 (N_1231,In_388,In_415);
nand U1232 (N_1232,In_293,In_306);
nand U1233 (N_1233,In_566,In_686);
or U1234 (N_1234,In_694,In_579);
nand U1235 (N_1235,In_702,In_713);
nor U1236 (N_1236,In_418,In_538);
nand U1237 (N_1237,In_345,In_336);
nor U1238 (N_1238,In_728,In_321);
and U1239 (N_1239,In_303,In_699);
or U1240 (N_1240,In_395,In_416);
nand U1241 (N_1241,In_88,In_95);
nor U1242 (N_1242,In_563,In_362);
and U1243 (N_1243,In_135,In_44);
nor U1244 (N_1244,In_519,In_735);
xnor U1245 (N_1245,In_660,In_272);
and U1246 (N_1246,In_106,In_276);
and U1247 (N_1247,In_654,In_391);
and U1248 (N_1248,In_430,In_740);
or U1249 (N_1249,In_71,In_616);
and U1250 (N_1250,In_264,In_307);
or U1251 (N_1251,In_151,In_58);
and U1252 (N_1252,In_565,In_249);
and U1253 (N_1253,In_277,In_574);
and U1254 (N_1254,In_687,In_369);
nand U1255 (N_1255,In_502,In_624);
nor U1256 (N_1256,In_539,In_83);
and U1257 (N_1257,In_32,In_39);
and U1258 (N_1258,In_718,In_239);
or U1259 (N_1259,In_110,In_554);
nand U1260 (N_1260,In_671,In_623);
xor U1261 (N_1261,In_553,In_123);
xnor U1262 (N_1262,In_367,In_373);
and U1263 (N_1263,In_731,In_290);
xor U1264 (N_1264,In_33,In_248);
nor U1265 (N_1265,In_99,In_101);
nor U1266 (N_1266,In_486,In_596);
or U1267 (N_1267,In_724,In_670);
nor U1268 (N_1268,In_386,In_440);
nand U1269 (N_1269,In_159,In_460);
nor U1270 (N_1270,In_409,In_477);
nand U1271 (N_1271,In_231,In_132);
or U1272 (N_1272,In_267,In_669);
or U1273 (N_1273,In_671,In_496);
nand U1274 (N_1274,In_48,In_480);
or U1275 (N_1275,In_302,In_203);
xnor U1276 (N_1276,In_224,In_23);
nand U1277 (N_1277,In_43,In_386);
or U1278 (N_1278,In_64,In_228);
or U1279 (N_1279,In_508,In_48);
nor U1280 (N_1280,In_118,In_509);
and U1281 (N_1281,In_731,In_88);
nand U1282 (N_1282,In_97,In_555);
nand U1283 (N_1283,In_286,In_256);
nand U1284 (N_1284,In_727,In_701);
nand U1285 (N_1285,In_399,In_11);
nor U1286 (N_1286,In_381,In_270);
nor U1287 (N_1287,In_732,In_704);
nand U1288 (N_1288,In_292,In_42);
nor U1289 (N_1289,In_509,In_200);
or U1290 (N_1290,In_315,In_424);
or U1291 (N_1291,In_608,In_298);
and U1292 (N_1292,In_706,In_37);
or U1293 (N_1293,In_10,In_109);
and U1294 (N_1294,In_612,In_166);
and U1295 (N_1295,In_30,In_288);
nor U1296 (N_1296,In_207,In_488);
or U1297 (N_1297,In_479,In_157);
and U1298 (N_1298,In_247,In_456);
xnor U1299 (N_1299,In_477,In_668);
or U1300 (N_1300,In_357,In_709);
and U1301 (N_1301,In_533,In_127);
and U1302 (N_1302,In_507,In_587);
xnor U1303 (N_1303,In_429,In_197);
nor U1304 (N_1304,In_739,In_64);
or U1305 (N_1305,In_372,In_517);
nand U1306 (N_1306,In_503,In_349);
or U1307 (N_1307,In_316,In_553);
nor U1308 (N_1308,In_155,In_611);
nor U1309 (N_1309,In_26,In_733);
nand U1310 (N_1310,In_432,In_219);
nor U1311 (N_1311,In_156,In_49);
nand U1312 (N_1312,In_441,In_644);
or U1313 (N_1313,In_485,In_290);
nand U1314 (N_1314,In_528,In_411);
and U1315 (N_1315,In_35,In_679);
xor U1316 (N_1316,In_12,In_396);
or U1317 (N_1317,In_277,In_384);
nor U1318 (N_1318,In_442,In_614);
or U1319 (N_1319,In_595,In_606);
nand U1320 (N_1320,In_456,In_484);
xor U1321 (N_1321,In_444,In_233);
nor U1322 (N_1322,In_107,In_519);
nand U1323 (N_1323,In_390,In_534);
and U1324 (N_1324,In_105,In_185);
and U1325 (N_1325,In_276,In_665);
and U1326 (N_1326,In_426,In_412);
nand U1327 (N_1327,In_237,In_320);
nand U1328 (N_1328,In_277,In_109);
nand U1329 (N_1329,In_200,In_228);
or U1330 (N_1330,In_435,In_699);
and U1331 (N_1331,In_250,In_514);
or U1332 (N_1332,In_470,In_133);
xnor U1333 (N_1333,In_743,In_647);
or U1334 (N_1334,In_460,In_524);
nand U1335 (N_1335,In_155,In_421);
nor U1336 (N_1336,In_114,In_607);
nand U1337 (N_1337,In_650,In_704);
nand U1338 (N_1338,In_94,In_445);
or U1339 (N_1339,In_697,In_681);
or U1340 (N_1340,In_98,In_663);
nor U1341 (N_1341,In_613,In_306);
and U1342 (N_1342,In_484,In_34);
xor U1343 (N_1343,In_325,In_390);
nor U1344 (N_1344,In_108,In_160);
or U1345 (N_1345,In_278,In_383);
or U1346 (N_1346,In_529,In_122);
nand U1347 (N_1347,In_709,In_26);
nand U1348 (N_1348,In_215,In_166);
or U1349 (N_1349,In_578,In_543);
and U1350 (N_1350,In_645,In_246);
xnor U1351 (N_1351,In_168,In_315);
or U1352 (N_1352,In_534,In_165);
nand U1353 (N_1353,In_669,In_353);
or U1354 (N_1354,In_284,In_98);
nor U1355 (N_1355,In_36,In_342);
or U1356 (N_1356,In_280,In_721);
or U1357 (N_1357,In_533,In_587);
nand U1358 (N_1358,In_95,In_647);
nor U1359 (N_1359,In_160,In_78);
nor U1360 (N_1360,In_9,In_308);
xor U1361 (N_1361,In_67,In_737);
and U1362 (N_1362,In_657,In_684);
and U1363 (N_1363,In_99,In_592);
nand U1364 (N_1364,In_482,In_678);
nand U1365 (N_1365,In_31,In_652);
or U1366 (N_1366,In_317,In_637);
or U1367 (N_1367,In_391,In_497);
and U1368 (N_1368,In_451,In_596);
xor U1369 (N_1369,In_719,In_616);
nand U1370 (N_1370,In_558,In_421);
nor U1371 (N_1371,In_405,In_348);
or U1372 (N_1372,In_211,In_637);
nand U1373 (N_1373,In_635,In_464);
nand U1374 (N_1374,In_616,In_657);
nor U1375 (N_1375,In_374,In_137);
and U1376 (N_1376,In_313,In_262);
nand U1377 (N_1377,In_571,In_163);
nand U1378 (N_1378,In_203,In_620);
xor U1379 (N_1379,In_436,In_475);
and U1380 (N_1380,In_291,In_731);
and U1381 (N_1381,In_500,In_324);
nand U1382 (N_1382,In_420,In_24);
nor U1383 (N_1383,In_10,In_124);
nand U1384 (N_1384,In_98,In_587);
nor U1385 (N_1385,In_522,In_255);
nor U1386 (N_1386,In_611,In_617);
or U1387 (N_1387,In_560,In_374);
and U1388 (N_1388,In_333,In_52);
and U1389 (N_1389,In_651,In_709);
and U1390 (N_1390,In_453,In_549);
nor U1391 (N_1391,In_320,In_77);
or U1392 (N_1392,In_32,In_43);
xnor U1393 (N_1393,In_137,In_256);
and U1394 (N_1394,In_154,In_67);
or U1395 (N_1395,In_185,In_726);
nor U1396 (N_1396,In_631,In_326);
or U1397 (N_1397,In_65,In_745);
or U1398 (N_1398,In_406,In_451);
or U1399 (N_1399,In_498,In_740);
nor U1400 (N_1400,In_465,In_23);
or U1401 (N_1401,In_370,In_642);
or U1402 (N_1402,In_265,In_247);
nor U1403 (N_1403,In_80,In_571);
or U1404 (N_1404,In_402,In_78);
xor U1405 (N_1405,In_574,In_119);
or U1406 (N_1406,In_710,In_10);
nor U1407 (N_1407,In_529,In_193);
nand U1408 (N_1408,In_602,In_273);
and U1409 (N_1409,In_395,In_37);
and U1410 (N_1410,In_108,In_326);
xnor U1411 (N_1411,In_18,In_191);
nor U1412 (N_1412,In_507,In_469);
and U1413 (N_1413,In_576,In_165);
or U1414 (N_1414,In_540,In_692);
and U1415 (N_1415,In_468,In_370);
and U1416 (N_1416,In_207,In_476);
or U1417 (N_1417,In_155,In_398);
and U1418 (N_1418,In_406,In_636);
nand U1419 (N_1419,In_499,In_165);
nor U1420 (N_1420,In_139,In_426);
xor U1421 (N_1421,In_571,In_103);
nand U1422 (N_1422,In_126,In_255);
nor U1423 (N_1423,In_665,In_457);
or U1424 (N_1424,In_395,In_474);
or U1425 (N_1425,In_229,In_12);
nor U1426 (N_1426,In_665,In_185);
and U1427 (N_1427,In_456,In_746);
or U1428 (N_1428,In_233,In_331);
or U1429 (N_1429,In_728,In_372);
nand U1430 (N_1430,In_161,In_234);
and U1431 (N_1431,In_444,In_505);
xor U1432 (N_1432,In_354,In_541);
nand U1433 (N_1433,In_327,In_263);
nand U1434 (N_1434,In_442,In_547);
nor U1435 (N_1435,In_159,In_373);
nand U1436 (N_1436,In_511,In_116);
or U1437 (N_1437,In_285,In_652);
nor U1438 (N_1438,In_523,In_576);
and U1439 (N_1439,In_456,In_489);
and U1440 (N_1440,In_34,In_661);
and U1441 (N_1441,In_680,In_432);
and U1442 (N_1442,In_461,In_291);
and U1443 (N_1443,In_497,In_225);
nand U1444 (N_1444,In_598,In_521);
or U1445 (N_1445,In_110,In_91);
or U1446 (N_1446,In_656,In_407);
nand U1447 (N_1447,In_312,In_101);
nor U1448 (N_1448,In_95,In_113);
nor U1449 (N_1449,In_388,In_85);
or U1450 (N_1450,In_532,In_250);
and U1451 (N_1451,In_394,In_731);
nor U1452 (N_1452,In_653,In_13);
nand U1453 (N_1453,In_749,In_343);
nor U1454 (N_1454,In_718,In_300);
and U1455 (N_1455,In_372,In_617);
nand U1456 (N_1456,In_17,In_738);
nand U1457 (N_1457,In_486,In_147);
and U1458 (N_1458,In_282,In_391);
or U1459 (N_1459,In_201,In_181);
and U1460 (N_1460,In_14,In_272);
nor U1461 (N_1461,In_207,In_156);
or U1462 (N_1462,In_453,In_300);
or U1463 (N_1463,In_130,In_78);
or U1464 (N_1464,In_279,In_645);
nor U1465 (N_1465,In_385,In_282);
nor U1466 (N_1466,In_740,In_674);
xnor U1467 (N_1467,In_171,In_235);
and U1468 (N_1468,In_740,In_585);
nand U1469 (N_1469,In_507,In_506);
nand U1470 (N_1470,In_151,In_252);
nor U1471 (N_1471,In_155,In_66);
nor U1472 (N_1472,In_359,In_173);
and U1473 (N_1473,In_436,In_637);
and U1474 (N_1474,In_719,In_602);
or U1475 (N_1475,In_1,In_647);
xnor U1476 (N_1476,In_336,In_571);
xor U1477 (N_1477,In_139,In_542);
or U1478 (N_1478,In_12,In_5);
nor U1479 (N_1479,In_29,In_497);
xnor U1480 (N_1480,In_396,In_579);
nor U1481 (N_1481,In_408,In_333);
or U1482 (N_1482,In_594,In_402);
or U1483 (N_1483,In_487,In_164);
or U1484 (N_1484,In_305,In_572);
and U1485 (N_1485,In_585,In_516);
and U1486 (N_1486,In_376,In_741);
or U1487 (N_1487,In_361,In_0);
nand U1488 (N_1488,In_303,In_514);
or U1489 (N_1489,In_82,In_243);
or U1490 (N_1490,In_411,In_67);
or U1491 (N_1491,In_596,In_62);
and U1492 (N_1492,In_747,In_579);
and U1493 (N_1493,In_479,In_270);
or U1494 (N_1494,In_529,In_198);
nand U1495 (N_1495,In_658,In_217);
or U1496 (N_1496,In_67,In_659);
or U1497 (N_1497,In_241,In_453);
and U1498 (N_1498,In_541,In_379);
or U1499 (N_1499,In_137,In_590);
nand U1500 (N_1500,In_73,In_222);
xor U1501 (N_1501,In_629,In_615);
or U1502 (N_1502,In_447,In_644);
nand U1503 (N_1503,In_56,In_468);
and U1504 (N_1504,In_196,In_550);
or U1505 (N_1505,In_453,In_464);
nand U1506 (N_1506,In_72,In_121);
or U1507 (N_1507,In_457,In_693);
nor U1508 (N_1508,In_76,In_366);
nor U1509 (N_1509,In_508,In_706);
or U1510 (N_1510,In_642,In_412);
or U1511 (N_1511,In_447,In_698);
or U1512 (N_1512,In_417,In_556);
nor U1513 (N_1513,In_640,In_467);
or U1514 (N_1514,In_341,In_430);
nand U1515 (N_1515,In_31,In_599);
or U1516 (N_1516,In_176,In_621);
and U1517 (N_1517,In_313,In_745);
nand U1518 (N_1518,In_160,In_588);
nor U1519 (N_1519,In_7,In_189);
and U1520 (N_1520,In_40,In_661);
or U1521 (N_1521,In_697,In_704);
nand U1522 (N_1522,In_220,In_475);
or U1523 (N_1523,In_61,In_222);
and U1524 (N_1524,In_67,In_677);
and U1525 (N_1525,In_635,In_713);
and U1526 (N_1526,In_744,In_33);
nand U1527 (N_1527,In_382,In_443);
and U1528 (N_1528,In_89,In_258);
nor U1529 (N_1529,In_45,In_579);
xnor U1530 (N_1530,In_121,In_574);
nand U1531 (N_1531,In_252,In_382);
nor U1532 (N_1532,In_430,In_308);
and U1533 (N_1533,In_705,In_541);
nor U1534 (N_1534,In_370,In_320);
nand U1535 (N_1535,In_461,In_224);
xnor U1536 (N_1536,In_59,In_317);
or U1537 (N_1537,In_230,In_286);
or U1538 (N_1538,In_358,In_114);
and U1539 (N_1539,In_672,In_64);
nor U1540 (N_1540,In_141,In_613);
and U1541 (N_1541,In_181,In_136);
and U1542 (N_1542,In_85,In_335);
or U1543 (N_1543,In_296,In_145);
nor U1544 (N_1544,In_243,In_164);
nand U1545 (N_1545,In_551,In_700);
nand U1546 (N_1546,In_260,In_98);
nor U1547 (N_1547,In_651,In_439);
nand U1548 (N_1548,In_396,In_256);
nor U1549 (N_1549,In_643,In_268);
nand U1550 (N_1550,In_245,In_624);
nor U1551 (N_1551,In_41,In_91);
xnor U1552 (N_1552,In_137,In_166);
nor U1553 (N_1553,In_419,In_583);
or U1554 (N_1554,In_376,In_223);
xnor U1555 (N_1555,In_37,In_541);
or U1556 (N_1556,In_410,In_168);
or U1557 (N_1557,In_573,In_287);
nor U1558 (N_1558,In_63,In_401);
and U1559 (N_1559,In_453,In_368);
or U1560 (N_1560,In_325,In_420);
and U1561 (N_1561,In_106,In_201);
and U1562 (N_1562,In_401,In_265);
nand U1563 (N_1563,In_711,In_448);
nand U1564 (N_1564,In_547,In_684);
or U1565 (N_1565,In_48,In_378);
or U1566 (N_1566,In_407,In_146);
and U1567 (N_1567,In_723,In_106);
and U1568 (N_1568,In_359,In_566);
and U1569 (N_1569,In_364,In_58);
and U1570 (N_1570,In_17,In_150);
nor U1571 (N_1571,In_740,In_646);
nand U1572 (N_1572,In_509,In_540);
xor U1573 (N_1573,In_304,In_614);
xnor U1574 (N_1574,In_206,In_256);
nor U1575 (N_1575,In_90,In_579);
and U1576 (N_1576,In_181,In_288);
nor U1577 (N_1577,In_312,In_27);
or U1578 (N_1578,In_493,In_290);
and U1579 (N_1579,In_683,In_499);
nor U1580 (N_1580,In_33,In_682);
nand U1581 (N_1581,In_395,In_100);
nor U1582 (N_1582,In_710,In_689);
nand U1583 (N_1583,In_511,In_553);
nor U1584 (N_1584,In_102,In_747);
nand U1585 (N_1585,In_543,In_30);
nor U1586 (N_1586,In_237,In_353);
xor U1587 (N_1587,In_257,In_526);
nor U1588 (N_1588,In_312,In_581);
or U1589 (N_1589,In_431,In_78);
nand U1590 (N_1590,In_365,In_348);
nand U1591 (N_1591,In_268,In_465);
and U1592 (N_1592,In_626,In_212);
or U1593 (N_1593,In_155,In_175);
and U1594 (N_1594,In_109,In_100);
nand U1595 (N_1595,In_276,In_387);
nand U1596 (N_1596,In_550,In_653);
nor U1597 (N_1597,In_425,In_717);
and U1598 (N_1598,In_343,In_164);
or U1599 (N_1599,In_323,In_105);
and U1600 (N_1600,In_366,In_697);
or U1601 (N_1601,In_636,In_517);
nor U1602 (N_1602,In_345,In_24);
nor U1603 (N_1603,In_586,In_138);
and U1604 (N_1604,In_689,In_522);
nand U1605 (N_1605,In_244,In_317);
and U1606 (N_1606,In_22,In_358);
and U1607 (N_1607,In_420,In_376);
nand U1608 (N_1608,In_601,In_568);
and U1609 (N_1609,In_387,In_129);
nor U1610 (N_1610,In_532,In_298);
xnor U1611 (N_1611,In_619,In_300);
and U1612 (N_1612,In_227,In_497);
nor U1613 (N_1613,In_353,In_118);
nor U1614 (N_1614,In_295,In_230);
and U1615 (N_1615,In_545,In_128);
or U1616 (N_1616,In_331,In_179);
and U1617 (N_1617,In_222,In_325);
and U1618 (N_1618,In_448,In_734);
nor U1619 (N_1619,In_206,In_508);
and U1620 (N_1620,In_742,In_184);
nand U1621 (N_1621,In_508,In_0);
nand U1622 (N_1622,In_468,In_30);
nor U1623 (N_1623,In_227,In_674);
xnor U1624 (N_1624,In_375,In_228);
nor U1625 (N_1625,In_649,In_741);
nor U1626 (N_1626,In_697,In_103);
xnor U1627 (N_1627,In_283,In_159);
or U1628 (N_1628,In_419,In_450);
nor U1629 (N_1629,In_119,In_512);
nor U1630 (N_1630,In_288,In_719);
nand U1631 (N_1631,In_452,In_398);
nand U1632 (N_1632,In_411,In_178);
and U1633 (N_1633,In_451,In_77);
or U1634 (N_1634,In_651,In_571);
nand U1635 (N_1635,In_437,In_651);
nand U1636 (N_1636,In_570,In_292);
nor U1637 (N_1637,In_186,In_646);
or U1638 (N_1638,In_477,In_746);
or U1639 (N_1639,In_443,In_194);
nor U1640 (N_1640,In_363,In_138);
xnor U1641 (N_1641,In_307,In_640);
and U1642 (N_1642,In_286,In_60);
nor U1643 (N_1643,In_655,In_211);
and U1644 (N_1644,In_9,In_500);
nand U1645 (N_1645,In_228,In_84);
nand U1646 (N_1646,In_734,In_52);
and U1647 (N_1647,In_559,In_12);
xor U1648 (N_1648,In_131,In_23);
and U1649 (N_1649,In_31,In_55);
and U1650 (N_1650,In_359,In_435);
nand U1651 (N_1651,In_309,In_251);
or U1652 (N_1652,In_362,In_562);
xnor U1653 (N_1653,In_691,In_519);
or U1654 (N_1654,In_206,In_567);
or U1655 (N_1655,In_666,In_392);
or U1656 (N_1656,In_188,In_245);
nor U1657 (N_1657,In_637,In_312);
or U1658 (N_1658,In_387,In_100);
nand U1659 (N_1659,In_121,In_221);
nor U1660 (N_1660,In_613,In_425);
nand U1661 (N_1661,In_496,In_521);
and U1662 (N_1662,In_525,In_722);
xor U1663 (N_1663,In_429,In_348);
nor U1664 (N_1664,In_290,In_147);
or U1665 (N_1665,In_709,In_667);
nor U1666 (N_1666,In_676,In_454);
nand U1667 (N_1667,In_315,In_382);
nor U1668 (N_1668,In_219,In_4);
or U1669 (N_1669,In_178,In_361);
and U1670 (N_1670,In_655,In_136);
or U1671 (N_1671,In_204,In_715);
and U1672 (N_1672,In_627,In_26);
nor U1673 (N_1673,In_238,In_301);
nand U1674 (N_1674,In_326,In_59);
nand U1675 (N_1675,In_138,In_66);
nand U1676 (N_1676,In_395,In_649);
nor U1677 (N_1677,In_485,In_702);
and U1678 (N_1678,In_642,In_167);
xor U1679 (N_1679,In_244,In_456);
nor U1680 (N_1680,In_298,In_61);
or U1681 (N_1681,In_173,In_651);
or U1682 (N_1682,In_51,In_229);
nand U1683 (N_1683,In_306,In_345);
and U1684 (N_1684,In_191,In_75);
nor U1685 (N_1685,In_32,In_621);
or U1686 (N_1686,In_131,In_117);
and U1687 (N_1687,In_387,In_516);
or U1688 (N_1688,In_50,In_345);
nor U1689 (N_1689,In_311,In_64);
xor U1690 (N_1690,In_609,In_643);
nor U1691 (N_1691,In_717,In_399);
nor U1692 (N_1692,In_175,In_553);
or U1693 (N_1693,In_416,In_265);
or U1694 (N_1694,In_256,In_41);
or U1695 (N_1695,In_184,In_461);
and U1696 (N_1696,In_436,In_70);
and U1697 (N_1697,In_252,In_470);
and U1698 (N_1698,In_650,In_26);
xor U1699 (N_1699,In_536,In_320);
nor U1700 (N_1700,In_153,In_410);
nand U1701 (N_1701,In_655,In_686);
and U1702 (N_1702,In_329,In_594);
nand U1703 (N_1703,In_371,In_420);
or U1704 (N_1704,In_532,In_56);
nand U1705 (N_1705,In_589,In_472);
and U1706 (N_1706,In_636,In_616);
and U1707 (N_1707,In_267,In_302);
nor U1708 (N_1708,In_196,In_151);
nor U1709 (N_1709,In_42,In_263);
xor U1710 (N_1710,In_193,In_552);
nor U1711 (N_1711,In_721,In_331);
nor U1712 (N_1712,In_90,In_20);
nor U1713 (N_1713,In_746,In_27);
nand U1714 (N_1714,In_667,In_188);
xnor U1715 (N_1715,In_345,In_171);
nor U1716 (N_1716,In_181,In_41);
or U1717 (N_1717,In_632,In_420);
or U1718 (N_1718,In_632,In_491);
nor U1719 (N_1719,In_426,In_326);
or U1720 (N_1720,In_378,In_531);
or U1721 (N_1721,In_140,In_42);
or U1722 (N_1722,In_717,In_191);
nor U1723 (N_1723,In_280,In_88);
nand U1724 (N_1724,In_134,In_559);
and U1725 (N_1725,In_395,In_587);
xnor U1726 (N_1726,In_4,In_300);
nor U1727 (N_1727,In_578,In_47);
and U1728 (N_1728,In_450,In_206);
and U1729 (N_1729,In_217,In_127);
nor U1730 (N_1730,In_523,In_169);
and U1731 (N_1731,In_276,In_710);
nand U1732 (N_1732,In_339,In_482);
or U1733 (N_1733,In_15,In_571);
nor U1734 (N_1734,In_345,In_225);
and U1735 (N_1735,In_589,In_304);
or U1736 (N_1736,In_324,In_520);
nand U1737 (N_1737,In_221,In_484);
nor U1738 (N_1738,In_157,In_500);
nor U1739 (N_1739,In_700,In_167);
nand U1740 (N_1740,In_716,In_141);
nor U1741 (N_1741,In_120,In_113);
nand U1742 (N_1742,In_182,In_38);
nand U1743 (N_1743,In_645,In_360);
nor U1744 (N_1744,In_454,In_257);
nand U1745 (N_1745,In_713,In_748);
nand U1746 (N_1746,In_420,In_44);
nand U1747 (N_1747,In_743,In_279);
nor U1748 (N_1748,In_501,In_194);
nand U1749 (N_1749,In_621,In_723);
nand U1750 (N_1750,In_203,In_494);
nand U1751 (N_1751,In_431,In_596);
and U1752 (N_1752,In_596,In_575);
nor U1753 (N_1753,In_219,In_131);
and U1754 (N_1754,In_198,In_96);
nor U1755 (N_1755,In_540,In_612);
and U1756 (N_1756,In_527,In_419);
or U1757 (N_1757,In_403,In_271);
nand U1758 (N_1758,In_466,In_232);
and U1759 (N_1759,In_476,In_19);
xor U1760 (N_1760,In_275,In_222);
nand U1761 (N_1761,In_475,In_437);
and U1762 (N_1762,In_137,In_3);
and U1763 (N_1763,In_525,In_199);
nand U1764 (N_1764,In_97,In_670);
and U1765 (N_1765,In_22,In_432);
or U1766 (N_1766,In_512,In_397);
or U1767 (N_1767,In_696,In_301);
or U1768 (N_1768,In_534,In_492);
and U1769 (N_1769,In_107,In_183);
nand U1770 (N_1770,In_523,In_583);
or U1771 (N_1771,In_618,In_120);
or U1772 (N_1772,In_712,In_680);
and U1773 (N_1773,In_210,In_486);
nor U1774 (N_1774,In_486,In_591);
and U1775 (N_1775,In_125,In_521);
nor U1776 (N_1776,In_157,In_510);
and U1777 (N_1777,In_624,In_546);
and U1778 (N_1778,In_465,In_604);
and U1779 (N_1779,In_637,In_263);
nand U1780 (N_1780,In_119,In_223);
and U1781 (N_1781,In_394,In_499);
or U1782 (N_1782,In_482,In_375);
or U1783 (N_1783,In_493,In_498);
or U1784 (N_1784,In_374,In_575);
nor U1785 (N_1785,In_250,In_643);
or U1786 (N_1786,In_75,In_420);
or U1787 (N_1787,In_208,In_480);
nand U1788 (N_1788,In_662,In_433);
and U1789 (N_1789,In_445,In_198);
nand U1790 (N_1790,In_229,In_104);
and U1791 (N_1791,In_585,In_607);
nor U1792 (N_1792,In_24,In_322);
and U1793 (N_1793,In_568,In_741);
nand U1794 (N_1794,In_406,In_509);
and U1795 (N_1795,In_704,In_600);
nand U1796 (N_1796,In_471,In_499);
or U1797 (N_1797,In_300,In_471);
nand U1798 (N_1798,In_676,In_55);
and U1799 (N_1799,In_710,In_292);
nand U1800 (N_1800,In_684,In_346);
or U1801 (N_1801,In_638,In_13);
nor U1802 (N_1802,In_346,In_286);
and U1803 (N_1803,In_142,In_28);
and U1804 (N_1804,In_340,In_81);
nand U1805 (N_1805,In_583,In_490);
and U1806 (N_1806,In_433,In_518);
nand U1807 (N_1807,In_61,In_701);
xnor U1808 (N_1808,In_610,In_385);
or U1809 (N_1809,In_530,In_16);
nor U1810 (N_1810,In_699,In_573);
nand U1811 (N_1811,In_197,In_328);
nor U1812 (N_1812,In_306,In_323);
nor U1813 (N_1813,In_200,In_343);
and U1814 (N_1814,In_126,In_56);
nor U1815 (N_1815,In_373,In_723);
or U1816 (N_1816,In_517,In_604);
and U1817 (N_1817,In_529,In_39);
or U1818 (N_1818,In_18,In_731);
nor U1819 (N_1819,In_13,In_97);
nand U1820 (N_1820,In_695,In_8);
and U1821 (N_1821,In_105,In_356);
nor U1822 (N_1822,In_68,In_290);
nor U1823 (N_1823,In_15,In_371);
nand U1824 (N_1824,In_33,In_711);
and U1825 (N_1825,In_54,In_682);
nand U1826 (N_1826,In_200,In_261);
nor U1827 (N_1827,In_191,In_290);
nor U1828 (N_1828,In_647,In_416);
nand U1829 (N_1829,In_191,In_32);
nand U1830 (N_1830,In_242,In_368);
nand U1831 (N_1831,In_162,In_732);
or U1832 (N_1832,In_741,In_244);
or U1833 (N_1833,In_54,In_199);
nand U1834 (N_1834,In_246,In_262);
nand U1835 (N_1835,In_63,In_561);
nand U1836 (N_1836,In_605,In_483);
and U1837 (N_1837,In_728,In_233);
or U1838 (N_1838,In_638,In_224);
or U1839 (N_1839,In_420,In_22);
or U1840 (N_1840,In_643,In_491);
nand U1841 (N_1841,In_627,In_476);
or U1842 (N_1842,In_675,In_102);
and U1843 (N_1843,In_616,In_707);
and U1844 (N_1844,In_150,In_154);
nor U1845 (N_1845,In_470,In_58);
and U1846 (N_1846,In_480,In_323);
nor U1847 (N_1847,In_263,In_253);
nand U1848 (N_1848,In_530,In_50);
and U1849 (N_1849,In_660,In_128);
xor U1850 (N_1850,In_707,In_60);
nor U1851 (N_1851,In_644,In_587);
nand U1852 (N_1852,In_391,In_215);
nor U1853 (N_1853,In_692,In_7);
nor U1854 (N_1854,In_734,In_504);
nor U1855 (N_1855,In_541,In_517);
nand U1856 (N_1856,In_507,In_29);
nor U1857 (N_1857,In_492,In_592);
nor U1858 (N_1858,In_657,In_506);
and U1859 (N_1859,In_12,In_149);
nor U1860 (N_1860,In_49,In_438);
nand U1861 (N_1861,In_549,In_206);
or U1862 (N_1862,In_701,In_411);
or U1863 (N_1863,In_541,In_71);
nand U1864 (N_1864,In_123,In_427);
nand U1865 (N_1865,In_365,In_407);
xnor U1866 (N_1866,In_402,In_637);
nor U1867 (N_1867,In_306,In_219);
nor U1868 (N_1868,In_353,In_70);
nor U1869 (N_1869,In_238,In_59);
and U1870 (N_1870,In_578,In_571);
nor U1871 (N_1871,In_655,In_389);
nor U1872 (N_1872,In_177,In_418);
and U1873 (N_1873,In_572,In_480);
nor U1874 (N_1874,In_320,In_621);
nor U1875 (N_1875,In_612,In_261);
or U1876 (N_1876,In_173,In_472);
nor U1877 (N_1877,In_46,In_736);
xnor U1878 (N_1878,In_700,In_214);
and U1879 (N_1879,In_273,In_154);
nor U1880 (N_1880,In_74,In_700);
xor U1881 (N_1881,In_295,In_742);
or U1882 (N_1882,In_662,In_76);
or U1883 (N_1883,In_718,In_543);
nand U1884 (N_1884,In_225,In_47);
nand U1885 (N_1885,In_582,In_300);
or U1886 (N_1886,In_42,In_297);
nand U1887 (N_1887,In_645,In_705);
or U1888 (N_1888,In_223,In_309);
nand U1889 (N_1889,In_108,In_146);
or U1890 (N_1890,In_253,In_12);
or U1891 (N_1891,In_351,In_457);
or U1892 (N_1892,In_338,In_249);
xor U1893 (N_1893,In_173,In_586);
nand U1894 (N_1894,In_489,In_420);
nand U1895 (N_1895,In_654,In_524);
nand U1896 (N_1896,In_555,In_179);
nand U1897 (N_1897,In_611,In_120);
and U1898 (N_1898,In_678,In_561);
or U1899 (N_1899,In_88,In_432);
and U1900 (N_1900,In_625,In_533);
nor U1901 (N_1901,In_194,In_14);
nand U1902 (N_1902,In_267,In_147);
nand U1903 (N_1903,In_246,In_76);
nand U1904 (N_1904,In_69,In_314);
nor U1905 (N_1905,In_6,In_269);
and U1906 (N_1906,In_726,In_53);
or U1907 (N_1907,In_147,In_186);
nor U1908 (N_1908,In_324,In_118);
nand U1909 (N_1909,In_400,In_77);
nor U1910 (N_1910,In_516,In_511);
or U1911 (N_1911,In_406,In_280);
nor U1912 (N_1912,In_559,In_339);
nand U1913 (N_1913,In_337,In_606);
or U1914 (N_1914,In_370,In_542);
nor U1915 (N_1915,In_597,In_9);
or U1916 (N_1916,In_431,In_121);
and U1917 (N_1917,In_578,In_492);
nand U1918 (N_1918,In_600,In_305);
nand U1919 (N_1919,In_432,In_491);
nand U1920 (N_1920,In_594,In_378);
nand U1921 (N_1921,In_259,In_183);
or U1922 (N_1922,In_202,In_437);
and U1923 (N_1923,In_448,In_247);
nand U1924 (N_1924,In_726,In_326);
nand U1925 (N_1925,In_734,In_523);
xnor U1926 (N_1926,In_699,In_471);
nand U1927 (N_1927,In_128,In_578);
and U1928 (N_1928,In_594,In_733);
and U1929 (N_1929,In_249,In_265);
xnor U1930 (N_1930,In_54,In_381);
and U1931 (N_1931,In_416,In_399);
nor U1932 (N_1932,In_587,In_186);
and U1933 (N_1933,In_529,In_136);
and U1934 (N_1934,In_413,In_168);
nor U1935 (N_1935,In_329,In_259);
or U1936 (N_1936,In_438,In_111);
nor U1937 (N_1937,In_31,In_137);
or U1938 (N_1938,In_553,In_676);
nand U1939 (N_1939,In_699,In_655);
nand U1940 (N_1940,In_42,In_700);
nand U1941 (N_1941,In_517,In_665);
nor U1942 (N_1942,In_12,In_174);
nand U1943 (N_1943,In_400,In_436);
and U1944 (N_1944,In_176,In_540);
nand U1945 (N_1945,In_359,In_398);
nand U1946 (N_1946,In_734,In_433);
nand U1947 (N_1947,In_593,In_670);
and U1948 (N_1948,In_199,In_623);
nand U1949 (N_1949,In_583,In_367);
nor U1950 (N_1950,In_283,In_48);
nand U1951 (N_1951,In_310,In_256);
nor U1952 (N_1952,In_259,In_161);
and U1953 (N_1953,In_663,In_631);
nor U1954 (N_1954,In_536,In_153);
nor U1955 (N_1955,In_378,In_23);
or U1956 (N_1956,In_482,In_611);
and U1957 (N_1957,In_646,In_40);
xnor U1958 (N_1958,In_182,In_97);
nand U1959 (N_1959,In_741,In_297);
nor U1960 (N_1960,In_99,In_172);
or U1961 (N_1961,In_266,In_135);
and U1962 (N_1962,In_0,In_96);
and U1963 (N_1963,In_587,In_671);
or U1964 (N_1964,In_634,In_290);
or U1965 (N_1965,In_36,In_309);
nor U1966 (N_1966,In_450,In_654);
xor U1967 (N_1967,In_99,In_236);
nor U1968 (N_1968,In_393,In_36);
nor U1969 (N_1969,In_71,In_485);
nand U1970 (N_1970,In_278,In_677);
or U1971 (N_1971,In_487,In_294);
and U1972 (N_1972,In_335,In_380);
xor U1973 (N_1973,In_528,In_498);
nand U1974 (N_1974,In_712,In_414);
nand U1975 (N_1975,In_647,In_380);
xor U1976 (N_1976,In_444,In_689);
and U1977 (N_1977,In_192,In_216);
nor U1978 (N_1978,In_340,In_319);
nand U1979 (N_1979,In_639,In_547);
or U1980 (N_1980,In_56,In_3);
or U1981 (N_1981,In_567,In_723);
nand U1982 (N_1982,In_382,In_11);
nand U1983 (N_1983,In_606,In_361);
or U1984 (N_1984,In_90,In_430);
nand U1985 (N_1985,In_556,In_63);
xor U1986 (N_1986,In_58,In_655);
nand U1987 (N_1987,In_484,In_408);
nor U1988 (N_1988,In_634,In_12);
and U1989 (N_1989,In_525,In_193);
xnor U1990 (N_1990,In_321,In_716);
xnor U1991 (N_1991,In_341,In_547);
or U1992 (N_1992,In_126,In_95);
or U1993 (N_1993,In_29,In_418);
xor U1994 (N_1994,In_340,In_397);
nor U1995 (N_1995,In_425,In_370);
or U1996 (N_1996,In_361,In_569);
nor U1997 (N_1997,In_656,In_127);
nand U1998 (N_1998,In_585,In_660);
and U1999 (N_1999,In_492,In_673);
or U2000 (N_2000,In_359,In_148);
nor U2001 (N_2001,In_732,In_374);
nand U2002 (N_2002,In_516,In_453);
nand U2003 (N_2003,In_621,In_579);
and U2004 (N_2004,In_601,In_664);
and U2005 (N_2005,In_395,In_706);
nor U2006 (N_2006,In_223,In_616);
and U2007 (N_2007,In_603,In_109);
or U2008 (N_2008,In_645,In_486);
or U2009 (N_2009,In_145,In_571);
nor U2010 (N_2010,In_506,In_93);
nand U2011 (N_2011,In_165,In_705);
or U2012 (N_2012,In_64,In_158);
xor U2013 (N_2013,In_210,In_62);
nor U2014 (N_2014,In_399,In_354);
nor U2015 (N_2015,In_584,In_554);
xor U2016 (N_2016,In_59,In_642);
xnor U2017 (N_2017,In_468,In_520);
nor U2018 (N_2018,In_20,In_42);
xor U2019 (N_2019,In_0,In_589);
nor U2020 (N_2020,In_2,In_314);
nor U2021 (N_2021,In_8,In_59);
nand U2022 (N_2022,In_714,In_41);
nand U2023 (N_2023,In_527,In_231);
nor U2024 (N_2024,In_706,In_184);
xnor U2025 (N_2025,In_198,In_226);
nor U2026 (N_2026,In_471,In_655);
nor U2027 (N_2027,In_158,In_56);
xor U2028 (N_2028,In_340,In_286);
nor U2029 (N_2029,In_635,In_692);
nor U2030 (N_2030,In_655,In_729);
nor U2031 (N_2031,In_162,In_334);
and U2032 (N_2032,In_736,In_151);
nand U2033 (N_2033,In_316,In_550);
and U2034 (N_2034,In_167,In_589);
xnor U2035 (N_2035,In_348,In_501);
and U2036 (N_2036,In_405,In_726);
and U2037 (N_2037,In_620,In_636);
nand U2038 (N_2038,In_718,In_665);
xor U2039 (N_2039,In_91,In_634);
nor U2040 (N_2040,In_335,In_601);
and U2041 (N_2041,In_718,In_278);
nand U2042 (N_2042,In_452,In_212);
and U2043 (N_2043,In_338,In_453);
or U2044 (N_2044,In_336,In_202);
or U2045 (N_2045,In_549,In_417);
or U2046 (N_2046,In_703,In_726);
and U2047 (N_2047,In_71,In_552);
or U2048 (N_2048,In_456,In_11);
nor U2049 (N_2049,In_340,In_84);
nand U2050 (N_2050,In_166,In_96);
nand U2051 (N_2051,In_493,In_169);
nand U2052 (N_2052,In_745,In_52);
nor U2053 (N_2053,In_371,In_96);
and U2054 (N_2054,In_478,In_8);
or U2055 (N_2055,In_192,In_33);
nor U2056 (N_2056,In_7,In_300);
or U2057 (N_2057,In_349,In_578);
xnor U2058 (N_2058,In_469,In_363);
nor U2059 (N_2059,In_471,In_290);
xnor U2060 (N_2060,In_464,In_617);
or U2061 (N_2061,In_695,In_462);
and U2062 (N_2062,In_80,In_558);
nand U2063 (N_2063,In_572,In_692);
and U2064 (N_2064,In_452,In_457);
nand U2065 (N_2065,In_742,In_595);
nand U2066 (N_2066,In_235,In_459);
nand U2067 (N_2067,In_116,In_76);
or U2068 (N_2068,In_397,In_264);
nand U2069 (N_2069,In_638,In_148);
and U2070 (N_2070,In_214,In_407);
nor U2071 (N_2071,In_352,In_611);
nand U2072 (N_2072,In_274,In_21);
or U2073 (N_2073,In_654,In_63);
nor U2074 (N_2074,In_713,In_157);
and U2075 (N_2075,In_90,In_63);
and U2076 (N_2076,In_522,In_150);
xor U2077 (N_2077,In_191,In_640);
nor U2078 (N_2078,In_531,In_131);
nor U2079 (N_2079,In_554,In_696);
and U2080 (N_2080,In_232,In_48);
or U2081 (N_2081,In_671,In_162);
and U2082 (N_2082,In_404,In_692);
and U2083 (N_2083,In_39,In_619);
or U2084 (N_2084,In_618,In_641);
nand U2085 (N_2085,In_560,In_320);
or U2086 (N_2086,In_370,In_373);
nor U2087 (N_2087,In_470,In_705);
nor U2088 (N_2088,In_616,In_685);
or U2089 (N_2089,In_154,In_683);
nand U2090 (N_2090,In_481,In_56);
and U2091 (N_2091,In_15,In_727);
nand U2092 (N_2092,In_661,In_257);
xor U2093 (N_2093,In_41,In_747);
or U2094 (N_2094,In_262,In_409);
or U2095 (N_2095,In_4,In_115);
nand U2096 (N_2096,In_512,In_58);
and U2097 (N_2097,In_279,In_656);
and U2098 (N_2098,In_554,In_124);
nand U2099 (N_2099,In_711,In_643);
and U2100 (N_2100,In_423,In_464);
or U2101 (N_2101,In_456,In_402);
nor U2102 (N_2102,In_518,In_448);
or U2103 (N_2103,In_94,In_394);
nand U2104 (N_2104,In_723,In_320);
nand U2105 (N_2105,In_543,In_141);
and U2106 (N_2106,In_278,In_183);
nand U2107 (N_2107,In_389,In_124);
nor U2108 (N_2108,In_274,In_334);
nand U2109 (N_2109,In_650,In_484);
or U2110 (N_2110,In_2,In_387);
or U2111 (N_2111,In_328,In_311);
nand U2112 (N_2112,In_593,In_414);
and U2113 (N_2113,In_170,In_599);
nor U2114 (N_2114,In_484,In_602);
and U2115 (N_2115,In_317,In_543);
and U2116 (N_2116,In_459,In_585);
nor U2117 (N_2117,In_440,In_723);
or U2118 (N_2118,In_171,In_272);
or U2119 (N_2119,In_104,In_596);
nor U2120 (N_2120,In_574,In_168);
or U2121 (N_2121,In_255,In_223);
or U2122 (N_2122,In_341,In_602);
or U2123 (N_2123,In_448,In_377);
nor U2124 (N_2124,In_217,In_551);
nor U2125 (N_2125,In_272,In_647);
or U2126 (N_2126,In_432,In_579);
nor U2127 (N_2127,In_192,In_459);
and U2128 (N_2128,In_150,In_354);
or U2129 (N_2129,In_459,In_438);
or U2130 (N_2130,In_17,In_112);
and U2131 (N_2131,In_724,In_412);
xor U2132 (N_2132,In_471,In_708);
and U2133 (N_2133,In_513,In_579);
xor U2134 (N_2134,In_321,In_76);
nand U2135 (N_2135,In_44,In_546);
or U2136 (N_2136,In_231,In_190);
nor U2137 (N_2137,In_198,In_507);
nand U2138 (N_2138,In_54,In_501);
nand U2139 (N_2139,In_722,In_592);
xnor U2140 (N_2140,In_26,In_112);
xor U2141 (N_2141,In_405,In_127);
and U2142 (N_2142,In_718,In_439);
or U2143 (N_2143,In_141,In_686);
and U2144 (N_2144,In_140,In_557);
or U2145 (N_2145,In_373,In_17);
or U2146 (N_2146,In_582,In_686);
nand U2147 (N_2147,In_256,In_14);
nand U2148 (N_2148,In_398,In_177);
nor U2149 (N_2149,In_465,In_508);
or U2150 (N_2150,In_320,In_227);
xor U2151 (N_2151,In_184,In_611);
and U2152 (N_2152,In_443,In_734);
xnor U2153 (N_2153,In_74,In_710);
and U2154 (N_2154,In_318,In_553);
and U2155 (N_2155,In_330,In_137);
nor U2156 (N_2156,In_270,In_51);
xor U2157 (N_2157,In_375,In_112);
nor U2158 (N_2158,In_514,In_434);
nor U2159 (N_2159,In_382,In_184);
nor U2160 (N_2160,In_716,In_37);
nand U2161 (N_2161,In_122,In_505);
or U2162 (N_2162,In_223,In_242);
and U2163 (N_2163,In_657,In_725);
nand U2164 (N_2164,In_512,In_385);
and U2165 (N_2165,In_160,In_732);
and U2166 (N_2166,In_415,In_594);
nor U2167 (N_2167,In_481,In_40);
nand U2168 (N_2168,In_674,In_158);
nand U2169 (N_2169,In_547,In_570);
and U2170 (N_2170,In_528,In_670);
and U2171 (N_2171,In_193,In_676);
nand U2172 (N_2172,In_589,In_470);
nor U2173 (N_2173,In_312,In_289);
xnor U2174 (N_2174,In_543,In_571);
or U2175 (N_2175,In_461,In_336);
and U2176 (N_2176,In_247,In_220);
nor U2177 (N_2177,In_206,In_749);
and U2178 (N_2178,In_442,In_392);
nand U2179 (N_2179,In_182,In_202);
or U2180 (N_2180,In_705,In_244);
nor U2181 (N_2181,In_198,In_742);
or U2182 (N_2182,In_579,In_724);
or U2183 (N_2183,In_366,In_674);
nor U2184 (N_2184,In_533,In_701);
and U2185 (N_2185,In_724,In_700);
xnor U2186 (N_2186,In_701,In_577);
and U2187 (N_2187,In_345,In_605);
or U2188 (N_2188,In_344,In_437);
or U2189 (N_2189,In_61,In_430);
nor U2190 (N_2190,In_725,In_637);
or U2191 (N_2191,In_351,In_444);
nor U2192 (N_2192,In_140,In_260);
or U2193 (N_2193,In_735,In_74);
nand U2194 (N_2194,In_493,In_92);
and U2195 (N_2195,In_418,In_715);
and U2196 (N_2196,In_436,In_593);
and U2197 (N_2197,In_449,In_543);
xor U2198 (N_2198,In_708,In_232);
nand U2199 (N_2199,In_729,In_711);
or U2200 (N_2200,In_516,In_544);
or U2201 (N_2201,In_699,In_226);
or U2202 (N_2202,In_615,In_226);
or U2203 (N_2203,In_330,In_465);
xor U2204 (N_2204,In_579,In_585);
nor U2205 (N_2205,In_23,In_249);
nor U2206 (N_2206,In_515,In_732);
and U2207 (N_2207,In_227,In_403);
xor U2208 (N_2208,In_140,In_526);
and U2209 (N_2209,In_749,In_26);
or U2210 (N_2210,In_198,In_739);
or U2211 (N_2211,In_721,In_103);
or U2212 (N_2212,In_309,In_696);
or U2213 (N_2213,In_576,In_371);
or U2214 (N_2214,In_375,In_399);
nor U2215 (N_2215,In_626,In_488);
and U2216 (N_2216,In_122,In_681);
and U2217 (N_2217,In_654,In_115);
and U2218 (N_2218,In_431,In_629);
and U2219 (N_2219,In_131,In_382);
or U2220 (N_2220,In_392,In_546);
nor U2221 (N_2221,In_605,In_19);
and U2222 (N_2222,In_415,In_598);
or U2223 (N_2223,In_368,In_659);
and U2224 (N_2224,In_660,In_1);
nand U2225 (N_2225,In_515,In_189);
or U2226 (N_2226,In_11,In_375);
or U2227 (N_2227,In_233,In_445);
or U2228 (N_2228,In_226,In_233);
nand U2229 (N_2229,In_78,In_176);
nand U2230 (N_2230,In_673,In_729);
or U2231 (N_2231,In_423,In_584);
and U2232 (N_2232,In_546,In_309);
or U2233 (N_2233,In_239,In_502);
nand U2234 (N_2234,In_507,In_72);
nor U2235 (N_2235,In_725,In_366);
nor U2236 (N_2236,In_381,In_613);
nor U2237 (N_2237,In_316,In_106);
nor U2238 (N_2238,In_515,In_486);
or U2239 (N_2239,In_554,In_356);
and U2240 (N_2240,In_501,In_260);
or U2241 (N_2241,In_610,In_99);
nor U2242 (N_2242,In_281,In_23);
xnor U2243 (N_2243,In_688,In_749);
or U2244 (N_2244,In_247,In_159);
nand U2245 (N_2245,In_520,In_256);
nand U2246 (N_2246,In_265,In_695);
or U2247 (N_2247,In_389,In_548);
and U2248 (N_2248,In_244,In_410);
and U2249 (N_2249,In_335,In_726);
and U2250 (N_2250,In_362,In_259);
nand U2251 (N_2251,In_10,In_633);
nand U2252 (N_2252,In_195,In_715);
xor U2253 (N_2253,In_206,In_638);
or U2254 (N_2254,In_497,In_6);
nand U2255 (N_2255,In_611,In_170);
and U2256 (N_2256,In_197,In_281);
nor U2257 (N_2257,In_570,In_693);
or U2258 (N_2258,In_25,In_199);
nor U2259 (N_2259,In_76,In_708);
nand U2260 (N_2260,In_1,In_366);
nand U2261 (N_2261,In_157,In_182);
xnor U2262 (N_2262,In_380,In_499);
nor U2263 (N_2263,In_64,In_153);
nor U2264 (N_2264,In_674,In_255);
and U2265 (N_2265,In_665,In_283);
xor U2266 (N_2266,In_686,In_135);
xor U2267 (N_2267,In_498,In_335);
nand U2268 (N_2268,In_277,In_398);
or U2269 (N_2269,In_204,In_401);
xnor U2270 (N_2270,In_176,In_451);
nand U2271 (N_2271,In_191,In_234);
and U2272 (N_2272,In_116,In_710);
xnor U2273 (N_2273,In_216,In_606);
xor U2274 (N_2274,In_542,In_503);
or U2275 (N_2275,In_371,In_356);
nand U2276 (N_2276,In_88,In_660);
xor U2277 (N_2277,In_578,In_351);
nor U2278 (N_2278,In_677,In_512);
xnor U2279 (N_2279,In_167,In_289);
nand U2280 (N_2280,In_692,In_210);
and U2281 (N_2281,In_680,In_94);
and U2282 (N_2282,In_443,In_313);
and U2283 (N_2283,In_207,In_491);
nand U2284 (N_2284,In_166,In_227);
nor U2285 (N_2285,In_649,In_309);
and U2286 (N_2286,In_309,In_606);
nand U2287 (N_2287,In_157,In_324);
xnor U2288 (N_2288,In_521,In_684);
nor U2289 (N_2289,In_576,In_72);
and U2290 (N_2290,In_555,In_286);
nor U2291 (N_2291,In_625,In_571);
nand U2292 (N_2292,In_521,In_134);
nand U2293 (N_2293,In_407,In_563);
or U2294 (N_2294,In_492,In_312);
nor U2295 (N_2295,In_28,In_364);
nor U2296 (N_2296,In_134,In_715);
xnor U2297 (N_2297,In_226,In_483);
nor U2298 (N_2298,In_174,In_424);
xnor U2299 (N_2299,In_618,In_104);
xnor U2300 (N_2300,In_692,In_337);
xor U2301 (N_2301,In_474,In_539);
or U2302 (N_2302,In_545,In_179);
nor U2303 (N_2303,In_177,In_335);
xnor U2304 (N_2304,In_293,In_80);
nand U2305 (N_2305,In_254,In_98);
or U2306 (N_2306,In_529,In_14);
nand U2307 (N_2307,In_393,In_56);
nand U2308 (N_2308,In_114,In_245);
nand U2309 (N_2309,In_378,In_570);
or U2310 (N_2310,In_157,In_27);
or U2311 (N_2311,In_678,In_628);
or U2312 (N_2312,In_558,In_120);
and U2313 (N_2313,In_692,In_726);
and U2314 (N_2314,In_345,In_421);
or U2315 (N_2315,In_596,In_19);
nand U2316 (N_2316,In_359,In_237);
nor U2317 (N_2317,In_188,In_473);
nor U2318 (N_2318,In_357,In_307);
nand U2319 (N_2319,In_322,In_390);
nand U2320 (N_2320,In_565,In_356);
xor U2321 (N_2321,In_724,In_689);
and U2322 (N_2322,In_240,In_682);
nand U2323 (N_2323,In_691,In_139);
nor U2324 (N_2324,In_648,In_487);
nor U2325 (N_2325,In_540,In_14);
and U2326 (N_2326,In_386,In_400);
and U2327 (N_2327,In_430,In_568);
or U2328 (N_2328,In_122,In_601);
and U2329 (N_2329,In_49,In_727);
nand U2330 (N_2330,In_331,In_409);
nand U2331 (N_2331,In_329,In_103);
nand U2332 (N_2332,In_4,In_637);
nand U2333 (N_2333,In_426,In_177);
nor U2334 (N_2334,In_93,In_420);
nand U2335 (N_2335,In_103,In_426);
nand U2336 (N_2336,In_93,In_121);
xnor U2337 (N_2337,In_528,In_261);
nand U2338 (N_2338,In_582,In_147);
nor U2339 (N_2339,In_444,In_328);
xor U2340 (N_2340,In_535,In_476);
or U2341 (N_2341,In_555,In_72);
xor U2342 (N_2342,In_48,In_167);
and U2343 (N_2343,In_560,In_72);
xor U2344 (N_2344,In_181,In_517);
nand U2345 (N_2345,In_660,In_679);
and U2346 (N_2346,In_407,In_687);
and U2347 (N_2347,In_464,In_272);
or U2348 (N_2348,In_15,In_558);
and U2349 (N_2349,In_652,In_173);
and U2350 (N_2350,In_567,In_394);
or U2351 (N_2351,In_230,In_687);
xnor U2352 (N_2352,In_372,In_471);
nor U2353 (N_2353,In_394,In_675);
nor U2354 (N_2354,In_232,In_159);
and U2355 (N_2355,In_189,In_472);
and U2356 (N_2356,In_539,In_747);
nor U2357 (N_2357,In_303,In_39);
xor U2358 (N_2358,In_61,In_500);
nand U2359 (N_2359,In_232,In_421);
nor U2360 (N_2360,In_697,In_10);
and U2361 (N_2361,In_328,In_208);
and U2362 (N_2362,In_683,In_682);
or U2363 (N_2363,In_263,In_378);
nand U2364 (N_2364,In_432,In_285);
nor U2365 (N_2365,In_565,In_552);
or U2366 (N_2366,In_500,In_180);
or U2367 (N_2367,In_128,In_368);
and U2368 (N_2368,In_244,In_590);
or U2369 (N_2369,In_522,In_192);
nand U2370 (N_2370,In_105,In_440);
nand U2371 (N_2371,In_366,In_431);
or U2372 (N_2372,In_34,In_573);
or U2373 (N_2373,In_46,In_146);
or U2374 (N_2374,In_313,In_537);
nand U2375 (N_2375,In_720,In_56);
nor U2376 (N_2376,In_308,In_720);
and U2377 (N_2377,In_608,In_550);
nand U2378 (N_2378,In_215,In_383);
and U2379 (N_2379,In_184,In_561);
xor U2380 (N_2380,In_459,In_487);
nand U2381 (N_2381,In_552,In_288);
nor U2382 (N_2382,In_728,In_629);
and U2383 (N_2383,In_460,In_514);
and U2384 (N_2384,In_700,In_301);
nor U2385 (N_2385,In_539,In_469);
or U2386 (N_2386,In_680,In_513);
nand U2387 (N_2387,In_541,In_551);
or U2388 (N_2388,In_14,In_651);
xnor U2389 (N_2389,In_738,In_30);
or U2390 (N_2390,In_284,In_656);
or U2391 (N_2391,In_428,In_432);
nand U2392 (N_2392,In_444,In_748);
and U2393 (N_2393,In_355,In_256);
nand U2394 (N_2394,In_541,In_341);
nand U2395 (N_2395,In_740,In_142);
or U2396 (N_2396,In_57,In_585);
and U2397 (N_2397,In_199,In_123);
nand U2398 (N_2398,In_431,In_661);
and U2399 (N_2399,In_29,In_221);
nor U2400 (N_2400,In_537,In_619);
nand U2401 (N_2401,In_97,In_454);
or U2402 (N_2402,In_250,In_553);
and U2403 (N_2403,In_560,In_335);
and U2404 (N_2404,In_359,In_502);
nor U2405 (N_2405,In_649,In_432);
nand U2406 (N_2406,In_219,In_735);
or U2407 (N_2407,In_672,In_326);
xnor U2408 (N_2408,In_159,In_11);
nor U2409 (N_2409,In_247,In_441);
or U2410 (N_2410,In_72,In_66);
and U2411 (N_2411,In_655,In_120);
nor U2412 (N_2412,In_472,In_58);
and U2413 (N_2413,In_211,In_710);
nor U2414 (N_2414,In_354,In_298);
or U2415 (N_2415,In_424,In_434);
nor U2416 (N_2416,In_350,In_230);
nor U2417 (N_2417,In_162,In_594);
and U2418 (N_2418,In_424,In_142);
nor U2419 (N_2419,In_724,In_536);
nand U2420 (N_2420,In_117,In_127);
or U2421 (N_2421,In_361,In_589);
nand U2422 (N_2422,In_277,In_311);
nor U2423 (N_2423,In_348,In_224);
and U2424 (N_2424,In_158,In_290);
nand U2425 (N_2425,In_605,In_164);
nor U2426 (N_2426,In_478,In_1);
or U2427 (N_2427,In_298,In_541);
nand U2428 (N_2428,In_64,In_366);
and U2429 (N_2429,In_506,In_88);
or U2430 (N_2430,In_301,In_568);
and U2431 (N_2431,In_265,In_466);
or U2432 (N_2432,In_694,In_327);
xnor U2433 (N_2433,In_663,In_59);
or U2434 (N_2434,In_23,In_316);
xor U2435 (N_2435,In_612,In_649);
nor U2436 (N_2436,In_355,In_59);
nor U2437 (N_2437,In_537,In_272);
nor U2438 (N_2438,In_300,In_175);
nand U2439 (N_2439,In_484,In_707);
and U2440 (N_2440,In_477,In_632);
and U2441 (N_2441,In_110,In_705);
nand U2442 (N_2442,In_427,In_290);
nand U2443 (N_2443,In_153,In_112);
nor U2444 (N_2444,In_586,In_201);
nand U2445 (N_2445,In_437,In_577);
xor U2446 (N_2446,In_575,In_162);
xor U2447 (N_2447,In_523,In_185);
and U2448 (N_2448,In_105,In_615);
and U2449 (N_2449,In_518,In_231);
and U2450 (N_2450,In_156,In_538);
nor U2451 (N_2451,In_596,In_503);
xnor U2452 (N_2452,In_326,In_369);
or U2453 (N_2453,In_224,In_679);
nand U2454 (N_2454,In_123,In_658);
nand U2455 (N_2455,In_350,In_268);
or U2456 (N_2456,In_303,In_268);
nand U2457 (N_2457,In_622,In_685);
nand U2458 (N_2458,In_550,In_667);
or U2459 (N_2459,In_215,In_233);
or U2460 (N_2460,In_743,In_468);
nand U2461 (N_2461,In_211,In_497);
xnor U2462 (N_2462,In_529,In_593);
or U2463 (N_2463,In_712,In_377);
xor U2464 (N_2464,In_376,In_377);
xor U2465 (N_2465,In_426,In_344);
and U2466 (N_2466,In_548,In_186);
and U2467 (N_2467,In_492,In_173);
nand U2468 (N_2468,In_259,In_734);
or U2469 (N_2469,In_62,In_1);
nand U2470 (N_2470,In_543,In_164);
or U2471 (N_2471,In_85,In_30);
nand U2472 (N_2472,In_734,In_158);
and U2473 (N_2473,In_557,In_193);
nand U2474 (N_2474,In_23,In_232);
xnor U2475 (N_2475,In_594,In_40);
nor U2476 (N_2476,In_115,In_271);
nand U2477 (N_2477,In_258,In_316);
and U2478 (N_2478,In_431,In_231);
xor U2479 (N_2479,In_632,In_416);
and U2480 (N_2480,In_244,In_698);
or U2481 (N_2481,In_89,In_552);
and U2482 (N_2482,In_17,In_580);
xor U2483 (N_2483,In_69,In_736);
nand U2484 (N_2484,In_171,In_209);
nand U2485 (N_2485,In_737,In_405);
and U2486 (N_2486,In_356,In_406);
xnor U2487 (N_2487,In_371,In_164);
xnor U2488 (N_2488,In_499,In_491);
and U2489 (N_2489,In_170,In_246);
and U2490 (N_2490,In_112,In_163);
nand U2491 (N_2491,In_421,In_141);
xnor U2492 (N_2492,In_336,In_198);
and U2493 (N_2493,In_298,In_105);
and U2494 (N_2494,In_380,In_459);
and U2495 (N_2495,In_655,In_561);
and U2496 (N_2496,In_497,In_49);
or U2497 (N_2497,In_314,In_177);
nand U2498 (N_2498,In_729,In_459);
nor U2499 (N_2499,In_461,In_653);
nand U2500 (N_2500,N_1799,N_1783);
or U2501 (N_2501,N_97,N_704);
nand U2502 (N_2502,N_1369,N_2037);
nand U2503 (N_2503,N_1360,N_1159);
and U2504 (N_2504,N_668,N_267);
nor U2505 (N_2505,N_424,N_222);
nand U2506 (N_2506,N_268,N_154);
and U2507 (N_2507,N_1509,N_1145);
and U2508 (N_2508,N_730,N_1128);
nand U2509 (N_2509,N_1847,N_2061);
nor U2510 (N_2510,N_944,N_751);
xor U2511 (N_2511,N_1584,N_1703);
xor U2512 (N_2512,N_547,N_408);
nand U2513 (N_2513,N_1324,N_1232);
nand U2514 (N_2514,N_1293,N_1662);
and U2515 (N_2515,N_1184,N_114);
nand U2516 (N_2516,N_2430,N_2383);
and U2517 (N_2517,N_1951,N_647);
nand U2518 (N_2518,N_672,N_61);
nand U2519 (N_2519,N_476,N_1877);
or U2520 (N_2520,N_1316,N_1588);
nand U2521 (N_2521,N_1716,N_1645);
and U2522 (N_2522,N_62,N_1370);
nand U2523 (N_2523,N_2,N_369);
or U2524 (N_2524,N_1601,N_1155);
xor U2525 (N_2525,N_1912,N_592);
and U2526 (N_2526,N_164,N_1607);
or U2527 (N_2527,N_181,N_1380);
nand U2528 (N_2528,N_80,N_823);
nand U2529 (N_2529,N_383,N_2208);
nor U2530 (N_2530,N_1001,N_1220);
nor U2531 (N_2531,N_2457,N_955);
nor U2532 (N_2532,N_2007,N_1253);
nand U2533 (N_2533,N_2235,N_209);
nor U2534 (N_2534,N_1344,N_885);
nor U2535 (N_2535,N_2470,N_2153);
xor U2536 (N_2536,N_1729,N_593);
or U2537 (N_2537,N_1850,N_1261);
xor U2538 (N_2538,N_1759,N_686);
nand U2539 (N_2539,N_1449,N_1243);
nand U2540 (N_2540,N_1735,N_1864);
nand U2541 (N_2541,N_131,N_481);
and U2542 (N_2542,N_2454,N_2310);
nand U2543 (N_2543,N_2452,N_2027);
nand U2544 (N_2544,N_1674,N_652);
xor U2545 (N_2545,N_337,N_859);
or U2546 (N_2546,N_1389,N_937);
nand U2547 (N_2547,N_1162,N_192);
nor U2548 (N_2548,N_2239,N_1970);
xor U2549 (N_2549,N_374,N_1646);
or U2550 (N_2550,N_565,N_1266);
or U2551 (N_2551,N_860,N_2317);
and U2552 (N_2552,N_146,N_230);
or U2553 (N_2553,N_563,N_1887);
and U2554 (N_2554,N_2070,N_1035);
nand U2555 (N_2555,N_67,N_572);
and U2556 (N_2556,N_667,N_2091);
and U2557 (N_2557,N_529,N_1955);
xor U2558 (N_2558,N_48,N_1422);
nand U2559 (N_2559,N_1636,N_1122);
and U2560 (N_2560,N_1577,N_894);
nand U2561 (N_2561,N_1515,N_1121);
nand U2562 (N_2562,N_1846,N_1358);
nand U2563 (N_2563,N_1227,N_1055);
nor U2564 (N_2564,N_1278,N_1530);
nand U2565 (N_2565,N_2339,N_1805);
nor U2566 (N_2566,N_2322,N_2097);
xor U2567 (N_2567,N_1106,N_95);
nor U2568 (N_2568,N_1375,N_1158);
xor U2569 (N_2569,N_486,N_37);
xnor U2570 (N_2570,N_2456,N_604);
and U2571 (N_2571,N_362,N_510);
and U2572 (N_2572,N_1031,N_2067);
xnor U2573 (N_2573,N_1903,N_1342);
nand U2574 (N_2574,N_1057,N_516);
or U2575 (N_2575,N_120,N_2121);
and U2576 (N_2576,N_938,N_579);
nor U2577 (N_2577,N_1394,N_513);
nand U2578 (N_2578,N_1612,N_1032);
and U2579 (N_2579,N_2250,N_1125);
and U2580 (N_2580,N_1284,N_2428);
or U2581 (N_2581,N_2396,N_52);
or U2582 (N_2582,N_2342,N_869);
or U2583 (N_2583,N_653,N_2432);
nand U2584 (N_2584,N_1542,N_465);
nand U2585 (N_2585,N_1295,N_1466);
xor U2586 (N_2586,N_2493,N_1000);
or U2587 (N_2587,N_204,N_2426);
nand U2588 (N_2588,N_1798,N_1407);
xor U2589 (N_2589,N_916,N_1428);
nor U2590 (N_2590,N_241,N_182);
and U2591 (N_2591,N_1061,N_1883);
nor U2592 (N_2592,N_750,N_489);
or U2593 (N_2593,N_2045,N_626);
nor U2594 (N_2594,N_742,N_2006);
nor U2595 (N_2595,N_1708,N_173);
nand U2596 (N_2596,N_2467,N_536);
or U2597 (N_2597,N_1187,N_281);
nor U2598 (N_2598,N_1858,N_1852);
nor U2599 (N_2599,N_307,N_2084);
nand U2600 (N_2600,N_84,N_1787);
nand U2601 (N_2601,N_2032,N_1815);
nor U2602 (N_2602,N_971,N_2170);
nor U2603 (N_2603,N_380,N_545);
nand U2604 (N_2604,N_1445,N_1393);
xnor U2605 (N_2605,N_2159,N_1066);
nand U2606 (N_2606,N_1839,N_1690);
nand U2607 (N_2607,N_445,N_138);
nand U2608 (N_2608,N_976,N_893);
nand U2609 (N_2609,N_189,N_1696);
or U2610 (N_2610,N_846,N_1754);
nor U2611 (N_2611,N_1681,N_770);
or U2612 (N_2612,N_1593,N_2439);
and U2613 (N_2613,N_1873,N_1549);
nor U2614 (N_2614,N_2196,N_733);
or U2615 (N_2615,N_649,N_387);
nor U2616 (N_2616,N_769,N_1913);
and U2617 (N_2617,N_969,N_562);
and U2618 (N_2618,N_1443,N_2053);
nand U2619 (N_2619,N_2217,N_661);
nand U2620 (N_2620,N_806,N_2259);
nand U2621 (N_2621,N_1048,N_79);
nor U2622 (N_2622,N_2017,N_1015);
nand U2623 (N_2623,N_2424,N_124);
and U2624 (N_2624,N_2368,N_240);
and U2625 (N_2625,N_1643,N_835);
nand U2626 (N_2626,N_2323,N_950);
nand U2627 (N_2627,N_2466,N_1596);
and U2628 (N_2628,N_2005,N_1074);
and U2629 (N_2629,N_1201,N_1969);
nor U2630 (N_2630,N_1855,N_345);
nor U2631 (N_2631,N_2230,N_1404);
or U2632 (N_2632,N_538,N_1830);
or U2633 (N_2633,N_928,N_2142);
nand U2634 (N_2634,N_1983,N_883);
nand U2635 (N_2635,N_2035,N_472);
and U2636 (N_2636,N_1533,N_30);
nor U2637 (N_2637,N_258,N_2480);
nand U2638 (N_2638,N_1600,N_283);
and U2639 (N_2639,N_1745,N_225);
nand U2640 (N_2640,N_6,N_190);
and U2641 (N_2641,N_1688,N_435);
nor U2642 (N_2642,N_1939,N_2102);
nand U2643 (N_2643,N_979,N_501);
and U2644 (N_2644,N_1764,N_1575);
nand U2645 (N_2645,N_1651,N_679);
and U2646 (N_2646,N_2023,N_1553);
xnor U2647 (N_2647,N_1896,N_2057);
xnor U2648 (N_2648,N_414,N_841);
nor U2649 (N_2649,N_2338,N_1457);
and U2650 (N_2650,N_537,N_940);
or U2651 (N_2651,N_1478,N_1368);
nor U2652 (N_2652,N_293,N_106);
or U2653 (N_2653,N_1954,N_2205);
nor U2654 (N_2654,N_171,N_1138);
and U2655 (N_2655,N_2346,N_556);
or U2656 (N_2656,N_375,N_2052);
nand U2657 (N_2657,N_543,N_505);
xnor U2658 (N_2658,N_598,N_1685);
or U2659 (N_2659,N_179,N_167);
or U2660 (N_2660,N_567,N_273);
nor U2661 (N_2661,N_546,N_1536);
and U2662 (N_2662,N_1237,N_555);
or U2663 (N_2663,N_1774,N_400);
nor U2664 (N_2664,N_1746,N_1808);
or U2665 (N_2665,N_1981,N_2247);
nor U2666 (N_2666,N_1565,N_1033);
nor U2667 (N_2667,N_735,N_2403);
and U2668 (N_2668,N_824,N_1824);
or U2669 (N_2669,N_450,N_2245);
nand U2670 (N_2670,N_585,N_1838);
xor U2671 (N_2671,N_2445,N_188);
and U2672 (N_2672,N_1788,N_1024);
xnor U2673 (N_2673,N_1297,N_930);
nor U2674 (N_2674,N_334,N_1377);
or U2675 (N_2675,N_474,N_2033);
nand U2676 (N_2676,N_316,N_2331);
nor U2677 (N_2677,N_1107,N_716);
or U2678 (N_2678,N_1854,N_2166);
and U2679 (N_2679,N_868,N_590);
or U2680 (N_2680,N_141,N_1611);
nand U2681 (N_2681,N_2462,N_1521);
nor U2682 (N_2682,N_959,N_1087);
and U2683 (N_2683,N_1019,N_266);
or U2684 (N_2684,N_1137,N_2326);
nor U2685 (N_2685,N_429,N_2270);
nor U2686 (N_2686,N_1231,N_1037);
and U2687 (N_2687,N_386,N_2287);
or U2688 (N_2688,N_927,N_1861);
xnor U2689 (N_2689,N_1627,N_632);
nor U2690 (N_2690,N_2391,N_508);
nand U2691 (N_2691,N_370,N_1283);
or U2692 (N_2692,N_2200,N_2181);
and U2693 (N_2693,N_640,N_1660);
nor U2694 (N_2694,N_625,N_1219);
nand U2695 (N_2695,N_150,N_557);
or U2696 (N_2696,N_1795,N_1492);
and U2697 (N_2697,N_1687,N_1326);
or U2698 (N_2698,N_1712,N_1430);
nor U2699 (N_2699,N_137,N_174);
and U2700 (N_2700,N_2406,N_515);
nand U2701 (N_2701,N_309,N_1144);
or U2702 (N_2702,N_24,N_2193);
and U2703 (N_2703,N_191,N_628);
nand U2704 (N_2704,N_985,N_787);
or U2705 (N_2705,N_44,N_1946);
nor U2706 (N_2706,N_872,N_25);
and U2707 (N_2707,N_558,N_1538);
xnor U2708 (N_2708,N_1263,N_518);
and U2709 (N_2709,N_1308,N_1349);
and U2710 (N_2710,N_2060,N_2114);
nand U2711 (N_2711,N_185,N_2284);
and U2712 (N_2712,N_493,N_402);
xnor U2713 (N_2713,N_2315,N_982);
and U2714 (N_2714,N_1244,N_78);
nor U2715 (N_2715,N_449,N_249);
nand U2716 (N_2716,N_499,N_1561);
and U2717 (N_2717,N_2025,N_368);
nand U2718 (N_2718,N_94,N_1556);
or U2719 (N_2719,N_1817,N_1290);
and U2720 (N_2720,N_1467,N_214);
or U2721 (N_2721,N_288,N_975);
nand U2722 (N_2722,N_977,N_33);
nor U2723 (N_2723,N_1083,N_63);
and U2724 (N_2724,N_411,N_1388);
or U2725 (N_2725,N_1099,N_797);
or U2726 (N_2726,N_327,N_1157);
and U2727 (N_2727,N_1541,N_2260);
or U2728 (N_2728,N_1923,N_330);
or U2729 (N_2729,N_2417,N_352);
and U2730 (N_2730,N_1414,N_2274);
nor U2731 (N_2731,N_2285,N_739);
nand U2732 (N_2732,N_2063,N_1365);
or U2733 (N_2733,N_1669,N_406);
nand U2734 (N_2734,N_1195,N_517);
nor U2735 (N_2735,N_170,N_713);
and U2736 (N_2736,N_1901,N_378);
nor U2737 (N_2737,N_1273,N_788);
nor U2738 (N_2738,N_31,N_1210);
and U2739 (N_2739,N_1989,N_905);
or U2740 (N_2740,N_2293,N_596);
or U2741 (N_2741,N_2248,N_1630);
or U2742 (N_2742,N_365,N_821);
nor U2743 (N_2743,N_1497,N_2115);
nor U2744 (N_2744,N_340,N_1747);
nor U2745 (N_2745,N_2283,N_569);
nand U2746 (N_2746,N_948,N_168);
and U2747 (N_2747,N_506,N_1357);
nor U2748 (N_2748,N_1870,N_287);
and U2749 (N_2749,N_7,N_1329);
nand U2750 (N_2750,N_1768,N_1049);
nand U2751 (N_2751,N_747,N_575);
and U2752 (N_2752,N_40,N_1776);
or U2753 (N_2753,N_1323,N_279);
or U2754 (N_2754,N_2148,N_539);
nand U2755 (N_2755,N_1415,N_2262);
and U2756 (N_2756,N_992,N_728);
nand U2757 (N_2757,N_2316,N_1733);
and U2758 (N_2758,N_798,N_426);
nand U2759 (N_2759,N_1248,N_332);
or U2760 (N_2760,N_1320,N_642);
or U2761 (N_2761,N_2477,N_2253);
nand U2762 (N_2762,N_943,N_1676);
nand U2763 (N_2763,N_754,N_14);
nor U2764 (N_2764,N_158,N_373);
or U2765 (N_2765,N_720,N_570);
nor U2766 (N_2766,N_961,N_2174);
xor U2767 (N_2767,N_2127,N_1914);
and U2768 (N_2768,N_2282,N_2377);
nand U2769 (N_2769,N_1664,N_1834);
and U2770 (N_2770,N_619,N_2358);
or U2771 (N_2771,N_1751,N_740);
and U2772 (N_2772,N_924,N_1406);
and U2773 (N_2773,N_2189,N_2435);
and U2774 (N_2774,N_2381,N_2167);
nand U2775 (N_2775,N_1392,N_1874);
nand U2776 (N_2776,N_932,N_1648);
nand U2777 (N_2777,N_791,N_1447);
xnor U2778 (N_2778,N_2337,N_1390);
and U2779 (N_2779,N_2160,N_528);
xnor U2780 (N_2780,N_1038,N_2072);
nor U2781 (N_2781,N_880,N_662);
nand U2782 (N_2782,N_1331,N_1111);
nor U2783 (N_2783,N_2373,N_1891);
xor U2784 (N_2784,N_576,N_1056);
nor U2785 (N_2785,N_521,N_3);
and U2786 (N_2786,N_1889,N_1285);
nor U2787 (N_2787,N_1828,N_66);
and U2788 (N_2788,N_2042,N_294);
and U2789 (N_2789,N_377,N_2483);
nor U2790 (N_2790,N_487,N_610);
or U2791 (N_2791,N_2175,N_1567);
nand U2792 (N_2792,N_1133,N_301);
or U2793 (N_2793,N_773,N_749);
nor U2794 (N_2794,N_336,N_525);
nor U2795 (N_2795,N_1677,N_1878);
or U2796 (N_2796,N_931,N_669);
and U2797 (N_2797,N_1827,N_882);
or U2798 (N_2798,N_2434,N_2487);
and U2799 (N_2799,N_715,N_1557);
nor U2800 (N_2800,N_1477,N_2416);
nand U2801 (N_2801,N_907,N_1930);
nand U2802 (N_2802,N_989,N_2050);
nor U2803 (N_2803,N_467,N_117);
nand U2804 (N_2804,N_404,N_1080);
nor U2805 (N_2805,N_395,N_1431);
nand U2806 (N_2806,N_1062,N_1282);
nand U2807 (N_2807,N_2471,N_1207);
nor U2808 (N_2808,N_1552,N_2139);
and U2809 (N_2809,N_1013,N_341);
nand U2810 (N_2810,N_857,N_1070);
nor U2811 (N_2811,N_1578,N_1624);
and U2812 (N_2812,N_612,N_1412);
and U2813 (N_2813,N_2078,N_2020);
xor U2814 (N_2814,N_2479,N_83);
nand U2815 (N_2815,N_2440,N_523);
or U2816 (N_2816,N_121,N_1836);
or U2817 (N_2817,N_1490,N_1860);
or U2818 (N_2818,N_211,N_559);
or U2819 (N_2819,N_2036,N_2375);
nor U2820 (N_2820,N_1045,N_1439);
or U2821 (N_2821,N_344,N_2008);
nor U2822 (N_2822,N_420,N_1474);
nor U2823 (N_2823,N_153,N_2179);
nand U2824 (N_2824,N_1863,N_1493);
or U2825 (N_2825,N_437,N_712);
nand U2826 (N_2826,N_2219,N_2028);
nor U2827 (N_2827,N_1671,N_1179);
nand U2828 (N_2828,N_243,N_808);
nor U2829 (N_2829,N_1785,N_1191);
nand U2830 (N_2830,N_1279,N_777);
and U2831 (N_2831,N_1178,N_681);
nand U2832 (N_2832,N_550,N_2103);
nor U2833 (N_2833,N_2224,N_2478);
and U2834 (N_2834,N_68,N_2222);
and U2835 (N_2835,N_727,N_804);
or U2836 (N_2836,N_2438,N_322);
or U2837 (N_2837,N_432,N_278);
or U2838 (N_2838,N_1054,N_1940);
nor U2839 (N_2839,N_1656,N_1103);
nor U2840 (N_2840,N_1338,N_331);
nand U2841 (N_2841,N_1996,N_82);
nor U2842 (N_2842,N_1879,N_691);
and U2843 (N_2843,N_280,N_1088);
nand U2844 (N_2844,N_1719,N_1780);
nand U2845 (N_2845,N_942,N_574);
nor U2846 (N_2846,N_891,N_1161);
nor U2847 (N_2847,N_852,N_1617);
nand U2848 (N_2848,N_469,N_2118);
or U2849 (N_2849,N_603,N_206);
or U2850 (N_2850,N_1315,N_2087);
nand U2851 (N_2851,N_621,N_2231);
and U2852 (N_2852,N_1200,N_744);
nor U2853 (N_2853,N_1194,N_219);
nand U2854 (N_2854,N_1059,N_1090);
xnor U2855 (N_2855,N_1075,N_1108);
and U2856 (N_2856,N_1869,N_65);
and U2857 (N_2857,N_2004,N_589);
nor U2858 (N_2858,N_674,N_2398);
nand U2859 (N_2859,N_1978,N_166);
and U2860 (N_2860,N_2335,N_552);
and U2861 (N_2861,N_195,N_312);
nor U2862 (N_2862,N_2343,N_466);
xor U2863 (N_2863,N_2297,N_542);
or U2864 (N_2864,N_101,N_242);
xor U2865 (N_2865,N_1968,N_1621);
or U2866 (N_2866,N_912,N_1757);
and U2867 (N_2867,N_2108,N_9);
nor U2868 (N_2868,N_1330,N_800);
and U2869 (N_2869,N_1188,N_933);
nand U2870 (N_2870,N_122,N_2360);
nand U2871 (N_2871,N_1794,N_1564);
or U2872 (N_2872,N_2152,N_990);
or U2873 (N_2873,N_425,N_439);
nor U2874 (N_2874,N_1228,N_1260);
or U2875 (N_2875,N_1765,N_151);
nand U2876 (N_2876,N_922,N_1622);
and U2877 (N_2877,N_1101,N_2492);
or U2878 (N_2878,N_1034,N_1772);
nor U2879 (N_2879,N_1420,N_323);
and U2880 (N_2880,N_1508,N_561);
nand U2881 (N_2881,N_946,N_274);
nor U2882 (N_2882,N_381,N_970);
xor U2883 (N_2883,N_987,N_1993);
nand U2884 (N_2884,N_2056,N_165);
and U2885 (N_2885,N_1756,N_615);
nor U2886 (N_2886,N_1892,N_271);
and U2887 (N_2887,N_1673,N_1152);
nand U2888 (N_2888,N_1618,N_2258);
nor U2889 (N_2889,N_1376,N_412);
nand U2890 (N_2890,N_656,N_111);
nor U2891 (N_2891,N_2051,N_996);
nand U2892 (N_2892,N_1257,N_698);
and U2893 (N_2893,N_2289,N_1303);
nand U2894 (N_2894,N_634,N_328);
xor U2895 (N_2895,N_2461,N_390);
nor U2896 (N_2896,N_430,N_1302);
and U2897 (N_2897,N_2228,N_1935);
nor U2898 (N_2898,N_1115,N_2420);
or U2899 (N_2899,N_376,N_1437);
and U2900 (N_2900,N_964,N_2355);
or U2901 (N_2901,N_702,N_1859);
nand U2902 (N_2902,N_1113,N_1829);
or U2903 (N_2903,N_655,N_1766);
nor U2904 (N_2904,N_379,N_361);
xnor U2905 (N_2905,N_1458,N_1398);
nor U2906 (N_2906,N_1845,N_921);
or U2907 (N_2907,N_1566,N_2264);
or U2908 (N_2908,N_866,N_2110);
and U2909 (N_2909,N_2000,N_757);
nand U2910 (N_2910,N_2155,N_2107);
nor U2911 (N_2911,N_701,N_2366);
xor U2912 (N_2912,N_488,N_1400);
nand U2913 (N_2913,N_2472,N_329);
nand U2914 (N_2914,N_867,N_398);
nand U2915 (N_2915,N_201,N_2234);
nor U2916 (N_2916,N_877,N_2216);
or U2917 (N_2917,N_1234,N_317);
nand U2918 (N_2918,N_1176,N_2252);
or U2919 (N_2919,N_588,N_1433);
and U2920 (N_2920,N_318,N_49);
nor U2921 (N_2921,N_2320,N_2085);
nand U2922 (N_2922,N_1555,N_1209);
and U2923 (N_2923,N_1429,N_2117);
and U2924 (N_2924,N_233,N_1701);
and U2925 (N_2925,N_2047,N_1792);
or U2926 (N_2926,N_614,N_1942);
and U2927 (N_2927,N_1820,N_1196);
or U2928 (N_2928,N_147,N_47);
nand U2929 (N_2929,N_1975,N_1314);
nand U2930 (N_2930,N_0,N_1306);
and U2931 (N_2931,N_2229,N_1345);
nand U2932 (N_2932,N_2187,N_436);
nand U2933 (N_2933,N_1175,N_1804);
nand U2934 (N_2934,N_2190,N_229);
nor U2935 (N_2935,N_1706,N_16);
or U2936 (N_2936,N_1097,N_811);
or U2937 (N_2937,N_1217,N_826);
or U2938 (N_2938,N_583,N_913);
nor U2939 (N_2939,N_34,N_237);
nand U2940 (N_2940,N_1713,N_1569);
nand U2941 (N_2941,N_706,N_433);
or U2942 (N_2942,N_908,N_973);
or U2943 (N_2943,N_198,N_926);
and U2944 (N_2944,N_782,N_1652);
and U2945 (N_2945,N_112,N_2133);
and U2946 (N_2946,N_1359,N_651);
and U2947 (N_2947,N_1548,N_1598);
nor U2948 (N_2948,N_1208,N_1026);
nor U2949 (N_2949,N_92,N_496);
and U2950 (N_2950,N_1129,N_721);
xor U2951 (N_2951,N_2495,N_2242);
and U2952 (N_2952,N_1665,N_494);
nand U2953 (N_2953,N_2237,N_2496);
or U2954 (N_2954,N_448,N_396);
nand U2955 (N_2955,N_1205,N_1505);
nor U2956 (N_2956,N_193,N_1897);
or U2957 (N_2957,N_650,N_531);
and U2958 (N_2958,N_2109,N_1763);
or U2959 (N_2959,N_1871,N_2198);
or U2960 (N_2960,N_127,N_1915);
nor U2961 (N_2961,N_1483,N_252);
or U2962 (N_2962,N_74,N_1559);
nand U2963 (N_2963,N_2223,N_1446);
and U2964 (N_2964,N_1654,N_1496);
nand U2965 (N_2965,N_2034,N_1917);
and U2966 (N_2966,N_2201,N_1695);
or U2967 (N_2967,N_915,N_1023);
or U2968 (N_2968,N_2347,N_708);
nand U2969 (N_2969,N_2497,N_890);
and U2970 (N_2970,N_2075,N_1758);
or U2971 (N_2971,N_2312,N_1868);
nor U2972 (N_2972,N_2350,N_1174);
or U2973 (N_2973,N_1378,N_296);
nand U2974 (N_2974,N_723,N_1215);
or U2975 (N_2975,N_1925,N_184);
and U2976 (N_2976,N_719,N_1929);
and U2977 (N_2977,N_1491,N_1614);
and U2978 (N_2978,N_2433,N_1427);
and U2979 (N_2979,N_2494,N_2130);
nor U2980 (N_2980,N_384,N_23);
or U2981 (N_2981,N_1164,N_1203);
nor U2982 (N_2982,N_1341,N_1539);
and U2983 (N_2983,N_1116,N_418);
xor U2984 (N_2984,N_128,N_571);
or U2985 (N_2985,N_69,N_1922);
xor U2986 (N_2986,N_1018,N_532);
xor U2987 (N_2987,N_1050,N_1076);
nor U2988 (N_2988,N_1364,N_1786);
or U2989 (N_2989,N_1988,N_364);
nand U2990 (N_2990,N_664,N_220);
nor U2991 (N_2991,N_1118,N_960);
nand U2992 (N_2992,N_729,N_974);
nor U2993 (N_2993,N_1570,N_1936);
or U2994 (N_2994,N_1047,N_2241);
nor U2995 (N_2995,N_2171,N_1030);
nor U2996 (N_2996,N_81,N_88);
nor U2997 (N_2997,N_1595,N_1843);
nor U2998 (N_2998,N_2275,N_1999);
nand U2999 (N_2999,N_825,N_2268);
nand U3000 (N_3000,N_64,N_736);
nand U3001 (N_3001,N_1945,N_1506);
nor U3002 (N_3002,N_1650,N_1580);
and U3003 (N_3003,N_1518,N_605);
and U3004 (N_3004,N_1503,N_1740);
and U3005 (N_3005,N_1347,N_1004);
or U3006 (N_3006,N_2288,N_236);
nand U3007 (N_3007,N_392,N_2092);
and U3008 (N_3008,N_1616,N_1069);
nor U3009 (N_3009,N_524,N_1348);
and U3010 (N_3010,N_1744,N_382);
or U3011 (N_3011,N_1259,N_1741);
nor U3012 (N_3012,N_876,N_836);
nand U3013 (N_3013,N_774,N_2340);
nor U3014 (N_3014,N_423,N_1327);
and U3015 (N_3015,N_2226,N_1619);
nor U3016 (N_3016,N_246,N_1325);
and U3017 (N_3017,N_1485,N_2038);
or U3018 (N_3018,N_2043,N_453);
or U3019 (N_3019,N_911,N_741);
and U3020 (N_3020,N_1513,N_1060);
or U3021 (N_3021,N_1736,N_1256);
and U3022 (N_3022,N_2380,N_693);
or U3023 (N_3023,N_760,N_2352);
nand U3024 (N_3024,N_2364,N_1318);
nor U3025 (N_3025,N_689,N_1790);
nor U3026 (N_3026,N_856,N_673);
nand U3027 (N_3027,N_658,N_665);
or U3028 (N_3028,N_454,N_289);
xor U3029 (N_3029,N_566,N_587);
and U3030 (N_3030,N_861,N_149);
nand U3031 (N_3031,N_1104,N_2279);
nor U3032 (N_3032,N_2041,N_1216);
and U3033 (N_3033,N_2098,N_1702);
or U3034 (N_3034,N_2123,N_1268);
nor U3035 (N_3035,N_2125,N_1663);
nand U3036 (N_3036,N_1222,N_633);
xor U3037 (N_3037,N_291,N_1867);
and U3038 (N_3038,N_276,N_1192);
nand U3039 (N_3039,N_2124,N_2306);
nor U3040 (N_3040,N_302,N_815);
nand U3041 (N_3041,N_2136,N_831);
xor U3042 (N_3042,N_553,N_677);
or U3043 (N_3043,N_1177,N_22);
nor U3044 (N_3044,N_1486,N_904);
and U3045 (N_3045,N_780,N_577);
and U3046 (N_3046,N_110,N_1748);
xor U3047 (N_3047,N_1098,N_1604);
or U3048 (N_3048,N_308,N_1352);
xnor U3049 (N_3049,N_853,N_1142);
or U3050 (N_3050,N_639,N_1705);
nor U3051 (N_3051,N_1250,N_1534);
nand U3052 (N_3052,N_60,N_1130);
nor U3053 (N_3053,N_2026,N_482);
or U3054 (N_3054,N_155,N_1294);
or U3055 (N_3055,N_1190,N_304);
nor U3056 (N_3056,N_1647,N_1762);
or U3057 (N_3057,N_116,N_1351);
nor U3058 (N_3058,N_2311,N_1507);
or U3059 (N_3059,N_186,N_1481);
and U3060 (N_3060,N_1910,N_459);
or U3061 (N_3061,N_1003,N_253);
or U3062 (N_3062,N_35,N_1720);
nor U3063 (N_3063,N_743,N_275);
nor U3064 (N_3064,N_796,N_1791);
nand U3065 (N_3065,N_2401,N_277);
nand U3066 (N_3066,N_1882,N_2307);
or U3067 (N_3067,N_1626,N_963);
nand U3068 (N_3068,N_135,N_1938);
and U3069 (N_3069,N_507,N_1373);
or U3070 (N_3070,N_1424,N_792);
and U3071 (N_3071,N_696,N_226);
nor U3072 (N_3072,N_879,N_53);
or U3073 (N_3073,N_2202,N_2015);
xor U3074 (N_3074,N_202,N_1147);
or U3075 (N_3075,N_1241,N_1608);
nor U3076 (N_3076,N_1469,N_1381);
nor U3077 (N_3077,N_1997,N_519);
and U3078 (N_3078,N_1806,N_397);
xnor U3079 (N_3079,N_1953,N_1299);
nand U3080 (N_3080,N_2269,N_203);
nor U3081 (N_3081,N_2120,N_1046);
or U3082 (N_3082,N_2176,N_786);
nand U3083 (N_3083,N_1710,N_761);
nand U3084 (N_3084,N_2313,N_2442);
or U3085 (N_3085,N_1737,N_159);
or U3086 (N_3086,N_1707,N_2210);
nand U3087 (N_3087,N_1771,N_1531);
or U3088 (N_3088,N_1949,N_1396);
nand U3089 (N_3089,N_2266,N_520);
nand U3090 (N_3090,N_2386,N_162);
or U3091 (N_3091,N_1840,N_2409);
or U3092 (N_3092,N_629,N_900);
and U3093 (N_3093,N_1831,N_297);
and U3094 (N_3094,N_939,N_1084);
nand U3095 (N_3095,N_2249,N_1148);
nand U3096 (N_3096,N_966,N_91);
nor U3097 (N_3097,N_350,N_1547);
or U3098 (N_3098,N_923,N_478);
nand U3099 (N_3099,N_607,N_1782);
and U3100 (N_3100,N_816,N_1753);
nand U3101 (N_3101,N_1286,N_503);
nand U3102 (N_3102,N_2425,N_901);
xnor U3103 (N_3103,N_779,N_2376);
and U3104 (N_3104,N_410,N_564);
nor U3105 (N_3105,N_1962,N_196);
nor U3106 (N_3106,N_645,N_2156);
or U3107 (N_3107,N_2418,N_1849);
or U3108 (N_3108,N_366,N_458);
xnor U3109 (N_3109,N_2195,N_1025);
and U3110 (N_3110,N_1770,N_2126);
or U3111 (N_3111,N_2390,N_21);
nor U3112 (N_3112,N_1010,N_1875);
and U3113 (N_3113,N_586,N_584);
nand U3114 (N_3114,N_611,N_261);
and U3115 (N_3115,N_259,N_951);
nand U3116 (N_3116,N_697,N_671);
nand U3117 (N_3117,N_2086,N_2162);
nand U3118 (N_3118,N_2140,N_1699);
and U3119 (N_3119,N_886,N_492);
nor U3120 (N_3120,N_2414,N_1073);
nand U3121 (N_3121,N_627,N_1944);
or U3122 (N_3122,N_1775,N_1722);
nor U3123 (N_3123,N_799,N_1535);
nor U3124 (N_3124,N_854,N_1212);
nand U3125 (N_3125,N_1068,N_945);
and U3126 (N_3126,N_1322,N_175);
and U3127 (N_3127,N_290,N_1704);
xnor U3128 (N_3128,N_2227,N_51);
and U3129 (N_3129,N_929,N_1202);
nor U3130 (N_3130,N_1550,N_403);
nand U3131 (N_3131,N_1450,N_142);
and U3132 (N_3132,N_1943,N_2164);
or U3133 (N_3133,N_1463,N_10);
xor U3134 (N_3134,N_631,N_2240);
or U3135 (N_3135,N_421,N_1246);
nor U3136 (N_3136,N_335,N_1473);
or U3137 (N_3137,N_1950,N_75);
nor U3138 (N_3138,N_2173,N_1150);
or U3139 (N_3139,N_512,N_1239);
nor U3140 (N_3140,N_1885,N_984);
and U3141 (N_3141,N_2001,N_1041);
nand U3142 (N_3142,N_1039,N_1029);
nor U3143 (N_3143,N_2066,N_2374);
and U3144 (N_3144,N_1694,N_1750);
nor U3145 (N_3145,N_793,N_1528);
nor U3146 (N_3146,N_2453,N_881);
nand U3147 (N_3147,N_637,N_385);
nand U3148 (N_3148,N_1139,N_2188);
xnor U3149 (N_3149,N_965,N_2415);
nand U3150 (N_3150,N_197,N_775);
xnor U3151 (N_3151,N_54,N_440);
or U3152 (N_3152,N_177,N_1081);
xor U3153 (N_3153,N_2255,N_1908);
or U3154 (N_3154,N_103,N_2336);
xor U3155 (N_3155,N_2341,N_2089);
nand U3156 (N_3156,N_636,N_1972);
and U3157 (N_3157,N_115,N_1634);
nand U3158 (N_3158,N_514,N_707);
or U3159 (N_3159,N_2286,N_2498);
xnor U3160 (N_3160,N_914,N_745);
or U3161 (N_3161,N_338,N_1848);
or U3162 (N_3162,N_212,N_36);
nor U3163 (N_3163,N_1317,N_2135);
nor U3164 (N_3164,N_903,N_443);
and U3165 (N_3165,N_1560,N_737);
and U3166 (N_3166,N_1832,N_2449);
nor U3167 (N_3167,N_2157,N_132);
and U3168 (N_3168,N_1519,N_772);
nor U3169 (N_3169,N_1937,N_1156);
and U3170 (N_3170,N_2044,N_1810);
and U3171 (N_3171,N_2094,N_980);
and U3172 (N_3172,N_2473,N_1511);
or U3173 (N_3173,N_2071,N_1620);
or U3174 (N_3174,N_1123,N_870);
or U3175 (N_3175,N_1451,N_2183);
nor U3176 (N_3176,N_1173,N_130);
and U3177 (N_3177,N_2112,N_2281);
or U3178 (N_3178,N_1906,N_2482);
or U3179 (N_3179,N_1354,N_999);
nand U3180 (N_3180,N_1568,N_1958);
or U3181 (N_3181,N_1992,N_1416);
or U3182 (N_3182,N_1255,N_1168);
and U3183 (N_3183,N_1180,N_157);
or U3184 (N_3184,N_1185,N_648);
nand U3185 (N_3185,N_896,N_1853);
xnor U3186 (N_3186,N_682,N_1361);
and U3187 (N_3187,N_1102,N_676);
or U3188 (N_3188,N_455,N_2019);
or U3189 (N_3189,N_1818,N_1258);
or U3190 (N_3190,N_920,N_1522);
nor U3191 (N_3191,N_865,N_1789);
or U3192 (N_3192,N_1272,N_1153);
nor U3193 (N_3193,N_832,N_1489);
or U3194 (N_3194,N_1426,N_1131);
xnor U3195 (N_3195,N_1374,N_2429);
xnor U3196 (N_3196,N_371,N_50);
or U3197 (N_3197,N_2238,N_2141);
or U3198 (N_3198,N_1402,N_1856);
and U3199 (N_3199,N_1058,N_292);
or U3200 (N_3200,N_1096,N_107);
and U3201 (N_3201,N_2122,N_1040);
and U3202 (N_3202,N_77,N_1558);
nor U3203 (N_3203,N_827,N_2408);
nor U3204 (N_3204,N_1957,N_1213);
or U3205 (N_3205,N_1198,N_1346);
and U3206 (N_3206,N_1623,N_257);
or U3207 (N_3207,N_1931,N_1974);
or U3208 (N_3208,N_1779,N_666);
nand U3209 (N_3209,N_580,N_2254);
nand U3210 (N_3210,N_480,N_962);
nor U3211 (N_3211,N_250,N_1067);
or U3212 (N_3212,N_39,N_299);
and U3213 (N_3213,N_2384,N_2314);
nand U3214 (N_3214,N_1275,N_1410);
nor U3215 (N_3215,N_2161,N_675);
or U3216 (N_3216,N_169,N_1385);
and U3217 (N_3217,N_232,N_2178);
nand U3218 (N_3218,N_1581,N_20);
and U3219 (N_3219,N_2367,N_1761);
xnor U3220 (N_3220,N_1668,N_100);
nor U3221 (N_3221,N_1441,N_1245);
or U3222 (N_3222,N_11,N_2400);
or U3223 (N_3223,N_1635,N_533);
xnor U3224 (N_3224,N_2484,N_695);
nor U3225 (N_3225,N_1807,N_731);
or U3226 (N_3226,N_1543,N_2134);
and U3227 (N_3227,N_573,N_1512);
or U3228 (N_3228,N_484,N_997);
nor U3229 (N_3229,N_2177,N_620);
nand U3230 (N_3230,N_358,N_1918);
or U3231 (N_3231,N_1254,N_1990);
and U3232 (N_3232,N_1709,N_753);
nand U3233 (N_3233,N_1924,N_871);
or U3234 (N_3234,N_972,N_670);
or U3235 (N_3235,N_2387,N_1952);
and U3236 (N_3236,N_711,N_541);
nor U3237 (N_3237,N_2489,N_1366);
nor U3238 (N_3238,N_1905,N_1238);
and U3239 (N_3239,N_251,N_692);
nand U3240 (N_3240,N_357,N_217);
or U3241 (N_3241,N_2191,N_783);
or U3242 (N_3242,N_994,N_2021);
xor U3243 (N_3243,N_2029,N_1265);
nor U3244 (N_3244,N_1526,N_722);
nand U3245 (N_3245,N_1796,N_452);
or U3246 (N_3246,N_123,N_1251);
or U3247 (N_3247,N_89,N_1926);
and U3248 (N_3248,N_427,N_830);
nand U3249 (N_3249,N_2304,N_1963);
nor U3250 (N_3250,N_2321,N_1639);
nand U3251 (N_3251,N_221,N_847);
nand U3252 (N_3252,N_1236,N_245);
or U3253 (N_3253,N_1141,N_784);
and U3254 (N_3254,N_326,N_144);
or U3255 (N_3255,N_1240,N_1339);
nor U3256 (N_3256,N_1452,N_909);
nand U3257 (N_3257,N_1977,N_200);
and U3258 (N_3258,N_2099,N_2054);
and U3259 (N_3259,N_2009,N_1135);
nor U3260 (N_3260,N_820,N_1328);
xor U3261 (N_3261,N_1382,N_1307);
nand U3262 (N_3262,N_247,N_1825);
nand U3263 (N_3263,N_1857,N_597);
or U3264 (N_3264,N_1684,N_145);
nand U3265 (N_3265,N_1340,N_2348);
or U3266 (N_3266,N_1143,N_1979);
nand U3267 (N_3267,N_1335,N_1464);
xor U3268 (N_3268,N_2441,N_227);
and U3269 (N_3269,N_1301,N_235);
or U3270 (N_3270,N_2003,N_2090);
xor U3271 (N_3271,N_1078,N_1998);
nand U3272 (N_3272,N_495,N_978);
nor U3273 (N_3273,N_457,N_981);
or U3274 (N_3274,N_98,N_2058);
or U3275 (N_3275,N_1487,N_1683);
or U3276 (N_3276,N_1632,N_2318);
or U3277 (N_3277,N_1079,N_952);
xnor U3278 (N_3278,N_1609,N_1119);
nor U3279 (N_3279,N_766,N_2443);
nand U3280 (N_3280,N_2407,N_2359);
xor U3281 (N_3281,N_1305,N_1384);
and U3282 (N_3282,N_1689,N_2382);
nand U3283 (N_3283,N_1814,N_897);
and U3284 (N_3284,N_1693,N_1514);
nand U3285 (N_3285,N_269,N_2192);
nor U3286 (N_3286,N_215,N_1933);
nand U3287 (N_3287,N_613,N_1233);
xnor U3288 (N_3288,N_1383,N_2299);
nor U3289 (N_3289,N_2147,N_444);
nand U3290 (N_3290,N_714,N_1304);
or U3291 (N_3291,N_1546,N_1661);
nand U3292 (N_3292,N_1605,N_405);
nand U3293 (N_3293,N_934,N_2199);
nor U3294 (N_3294,N_694,N_2308);
and U3295 (N_3295,N_594,N_349);
and U3296 (N_3296,N_2079,N_2393);
and U3297 (N_3297,N_1615,N_176);
nor U3298 (N_3298,N_1982,N_1523);
and U3299 (N_3299,N_2395,N_1154);
nor U3300 (N_3300,N_809,N_1409);
nor U3301 (N_3301,N_1743,N_2081);
nor U3302 (N_3302,N_1726,N_1909);
nor U3303 (N_3303,N_1865,N_616);
and U3304 (N_3304,N_1372,N_2203);
or U3305 (N_3305,N_1572,N_1961);
xnor U3306 (N_3306,N_355,N_2018);
and U3307 (N_3307,N_1277,N_1641);
or U3308 (N_3308,N_644,N_654);
and U3309 (N_3309,N_623,N_1151);
or U3310 (N_3310,N_1602,N_447);
nor U3311 (N_3311,N_1841,N_1221);
xnor U3312 (N_3312,N_1510,N_1028);
nor U3313 (N_3313,N_1551,N_343);
nand U3314 (N_3314,N_1051,N_342);
and U3315 (N_3315,N_256,N_1453);
and U3316 (N_3316,N_849,N_1071);
or U3317 (N_3317,N_2215,N_2132);
or U3318 (N_3318,N_19,N_2301);
or U3319 (N_3319,N_1252,N_2365);
nor U3320 (N_3320,N_1583,N_1343);
or U3321 (N_3321,N_2180,N_843);
nor U3322 (N_3322,N_560,N_568);
xor U3323 (N_3323,N_129,N_1995);
nand U3324 (N_3324,N_2271,N_428);
nand U3325 (N_3325,N_1900,N_2172);
nand U3326 (N_3326,N_497,N_734);
nand U3327 (N_3327,N_389,N_2333);
or U3328 (N_3328,N_887,N_1517);
or U3329 (N_3329,N_2378,N_2379);
and U3330 (N_3330,N_2291,N_600);
or U3331 (N_3331,N_1494,N_1711);
nand U3332 (N_3332,N_1613,N_1666);
and U3333 (N_3333,N_2068,N_2256);
xor U3334 (N_3334,N_1537,N_1670);
and U3335 (N_3335,N_2276,N_1739);
nor U3336 (N_3336,N_1095,N_785);
xnor U3337 (N_3337,N_199,N_462);
or U3338 (N_3338,N_2392,N_1127);
nand U3339 (N_3339,N_2490,N_2451);
and U3340 (N_3340,N_1866,N_956);
nor U3341 (N_3341,N_464,N_134);
xor U3342 (N_3342,N_477,N_1653);
nand U3343 (N_3343,N_643,N_238);
nand U3344 (N_3344,N_2212,N_1731);
nor U3345 (N_3345,N_732,N_2273);
and U3346 (N_3346,N_687,N_231);
nand U3347 (N_3347,N_314,N_889);
nor U3348 (N_3348,N_602,N_2372);
or U3349 (N_3349,N_2463,N_1092);
nand U3350 (N_3350,N_2149,N_1842);
xnor U3351 (N_3351,N_834,N_1310);
and U3352 (N_3352,N_888,N_2465);
xor U3353 (N_3353,N_534,N_1269);
xor U3354 (N_3354,N_2211,N_86);
and U3355 (N_3355,N_2186,N_2319);
nor U3356 (N_3356,N_409,N_1862);
or U3357 (N_3357,N_810,N_509);
nand U3358 (N_3358,N_554,N_70);
nand U3359 (N_3359,N_875,N_1321);
and U3360 (N_3360,N_446,N_2076);
nor U3361 (N_3361,N_72,N_2327);
nand U3362 (N_3362,N_1760,N_1379);
or U3363 (N_3363,N_1247,N_1082);
and U3364 (N_3364,N_125,N_630);
nor U3365 (N_3365,N_109,N_264);
nor U3366 (N_3366,N_1524,N_1333);
or U3367 (N_3367,N_548,N_286);
xnor U3368 (N_3368,N_1911,N_2437);
or U3369 (N_3369,N_1520,N_1472);
nand U3370 (N_3370,N_461,N_2476);
or U3371 (N_3371,N_684,N_2419);
or U3372 (N_3372,N_460,N_1065);
or U3373 (N_3373,N_1011,N_833);
and U3374 (N_3374,N_2303,N_1994);
nand U3375 (N_3375,N_8,N_38);
nor U3376 (N_3376,N_1440,N_700);
nor U3377 (N_3377,N_2328,N_422);
or U3378 (N_3378,N_1529,N_1163);
nor U3379 (N_3379,N_1484,N_2485);
and U3380 (N_3380,N_2491,N_1124);
xor U3381 (N_3381,N_2362,N_1730);
or U3382 (N_3382,N_391,N_442);
nand U3383 (N_3383,N_394,N_936);
and U3384 (N_3384,N_544,N_2486);
or U3385 (N_3385,N_438,N_2024);
xor U3386 (N_3386,N_2022,N_1967);
nand U3387 (N_3387,N_1525,N_606);
or U3388 (N_3388,N_1904,N_1021);
or U3389 (N_3389,N_85,N_1734);
nor U3390 (N_3390,N_967,N_957);
nand U3391 (N_3391,N_2151,N_183);
or U3392 (N_3392,N_1425,N_899);
nand U3393 (N_3393,N_1362,N_1460);
or U3394 (N_3394,N_339,N_262);
nor U3395 (N_3395,N_618,N_1585);
and U3396 (N_3396,N_1947,N_417);
or U3397 (N_3397,N_1966,N_2468);
nor U3398 (N_3398,N_1886,N_794);
and U3399 (N_3399,N_2232,N_470);
or U3400 (N_3400,N_2280,N_1386);
and U3401 (N_3401,N_1470,N_837);
nor U3402 (N_3402,N_56,N_260);
or U3403 (N_3403,N_2349,N_2411);
and U3404 (N_3404,N_1872,N_1170);
xor U3405 (N_3405,N_2158,N_348);
and U3406 (N_3406,N_244,N_1678);
and U3407 (N_3407,N_1455,N_2168);
nand U3408 (N_3408,N_272,N_2427);
and U3409 (N_3409,N_1941,N_2278);
nand U3410 (N_3410,N_2010,N_2448);
or U3411 (N_3411,N_862,N_2204);
nor U3412 (N_3412,N_2233,N_353);
nand U3413 (N_3413,N_254,N_1226);
nor U3414 (N_3414,N_1271,N_1987);
nor U3415 (N_3415,N_2064,N_1149);
nand U3416 (N_3416,N_139,N_1732);
and U3417 (N_3417,N_2351,N_2065);
nand U3418 (N_3418,N_161,N_1);
nand U3419 (N_3419,N_1971,N_1405);
nand U3420 (N_3420,N_917,N_1438);
nor U3421 (N_3421,N_1387,N_530);
nor U3422 (N_3422,N_1767,N_1920);
nand U3423 (N_3423,N_194,N_315);
nand U3424 (N_3424,N_2184,N_1714);
nor U3425 (N_3425,N_473,N_1752);
and U3426 (N_3426,N_475,N_1633);
nand U3427 (N_3427,N_725,N_143);
nor U3428 (N_3428,N_2455,N_1589);
or U3429 (N_3429,N_1884,N_2246);
or U3430 (N_3430,N_2332,N_763);
xnor U3431 (N_3431,N_1625,N_148);
nand U3432 (N_3432,N_1888,N_1006);
xor U3433 (N_3433,N_954,N_2357);
nor U3434 (N_3434,N_2111,N_850);
or U3435 (N_3435,N_2129,N_795);
nor U3436 (N_3436,N_1197,N_372);
and U3437 (N_3437,N_1742,N_500);
and U3438 (N_3438,N_1397,N_1435);
and U3439 (N_3439,N_346,N_2446);
or U3440 (N_3440,N_748,N_2128);
nor U3441 (N_3441,N_1292,N_320);
and U3442 (N_3442,N_925,N_1242);
or U3443 (N_3443,N_968,N_1803);
xnor U3444 (N_3444,N_947,N_71);
nor U3445 (N_3445,N_2488,N_858);
xnor U3446 (N_3446,N_1355,N_1017);
or U3447 (N_3447,N_840,N_1649);
nand U3448 (N_3448,N_210,N_1582);
or U3449 (N_3449,N_311,N_491);
and U3450 (N_3450,N_2263,N_2296);
or U3451 (N_3451,N_659,N_187);
nand U3452 (N_3452,N_813,N_705);
nor U3453 (N_3453,N_646,N_319);
nand U3454 (N_3454,N_419,N_1027);
and U3455 (N_3455,N_863,N_270);
or U3456 (N_3456,N_1738,N_1005);
and U3457 (N_3457,N_140,N_2404);
and U3458 (N_3458,N_1432,N_1371);
nor U3459 (N_3459,N_1403,N_1563);
nor U3460 (N_3460,N_2458,N_551);
or U3461 (N_3461,N_1391,N_2131);
xnor U3462 (N_3462,N_839,N_1475);
or U3463 (N_3463,N_1270,N_136);
or U3464 (N_3464,N_2046,N_703);
nor U3465 (N_3465,N_752,N_622);
or U3466 (N_3466,N_1899,N_2194);
or U3467 (N_3467,N_1679,N_1395);
nand U3468 (N_3468,N_2143,N_801);
nand U3469 (N_3469,N_1204,N_1105);
nor U3470 (N_3470,N_819,N_814);
nor U3471 (N_3471,N_988,N_822);
nand U3472 (N_3472,N_1399,N_1134);
or U3473 (N_3473,N_2334,N_57);
nor U3474 (N_3474,N_108,N_2305);
nand U3475 (N_3475,N_1659,N_1837);
nand U3476 (N_3476,N_1225,N_2016);
and U3477 (N_3477,N_1959,N_2356);
and U3478 (N_3478,N_1459,N_1146);
nand U3479 (N_3479,N_213,N_126);
and U3480 (N_3480,N_2389,N_1755);
or U3481 (N_3481,N_102,N_1591);
nand U3482 (N_3482,N_1211,N_310);
nor U3483 (N_3483,N_1419,N_2163);
nand U3484 (N_3484,N_46,N_1594);
and U3485 (N_3485,N_1544,N_2302);
and U3486 (N_3486,N_1498,N_2261);
or U3487 (N_3487,N_1717,N_73);
or U3488 (N_3488,N_678,N_1109);
nor U3489 (N_3489,N_1077,N_680);
nand U3490 (N_3490,N_1199,N_2014);
or U3491 (N_3491,N_41,N_1100);
nand U3492 (N_3492,N_2481,N_265);
and U3493 (N_3493,N_1298,N_205);
or U3494 (N_3494,N_2344,N_298);
nand U3495 (N_3495,N_1793,N_771);
xor U3496 (N_3496,N_1044,N_2300);
nor U3497 (N_3497,N_1628,N_1576);
and U3498 (N_3498,N_1022,N_581);
or U3499 (N_3499,N_617,N_527);
nor U3500 (N_3500,N_2225,N_1488);
xor U3501 (N_3501,N_1586,N_953);
or U3502 (N_3502,N_1927,N_958);
and U3503 (N_3503,N_802,N_1984);
or U3504 (N_3504,N_1725,N_1114);
or U3505 (N_3505,N_635,N_2290);
or U3506 (N_3506,N_1193,N_758);
nor U3507 (N_3507,N_1985,N_1692);
or U3508 (N_3508,N_1183,N_471);
nand U3509 (N_3509,N_1686,N_2104);
xor U3510 (N_3510,N_1587,N_1468);
nand U3511 (N_3511,N_1822,N_2423);
xnor U3512 (N_3512,N_838,N_608);
and U3513 (N_3513,N_1631,N_1700);
xnor U3514 (N_3514,N_1172,N_1089);
and U3515 (N_3515,N_1851,N_1960);
nor U3516 (N_3516,N_2447,N_842);
nand U3517 (N_3517,N_776,N_2218);
and U3518 (N_3518,N_1189,N_683);
nor U3519 (N_3519,N_1675,N_2095);
and U3520 (N_3520,N_2105,N_1085);
nor U3521 (N_3521,N_45,N_1337);
nor U3522 (N_3522,N_781,N_1644);
and U3523 (N_3523,N_1826,N_2475);
or U3524 (N_3524,N_1319,N_1291);
and U3525 (N_3525,N_2431,N_2436);
nand U3526 (N_3526,N_1444,N_2012);
nor U3527 (N_3527,N_578,N_463);
or U3528 (N_3528,N_1436,N_2138);
nor U3529 (N_3529,N_709,N_32);
nand U3530 (N_3530,N_1007,N_223);
nand U3531 (N_3531,N_2292,N_324);
nand U3532 (N_3532,N_2257,N_657);
and U3533 (N_3533,N_2002,N_300);
or U3534 (N_3534,N_224,N_1063);
and U3535 (N_3535,N_1721,N_726);
xnor U3536 (N_3536,N_1890,N_1500);
xor U3537 (N_3537,N_1811,N_1223);
nor U3538 (N_3538,N_2221,N_738);
nand U3539 (N_3539,N_2150,N_263);
or U3540 (N_3540,N_27,N_1812);
or U3541 (N_3541,N_1956,N_415);
and U3542 (N_3542,N_2083,N_1727);
nand U3543 (N_3543,N_768,N_535);
and U3544 (N_3544,N_285,N_1160);
xnor U3545 (N_3545,N_874,N_1976);
nand U3546 (N_3546,N_363,N_2106);
nand U3547 (N_3547,N_502,N_2169);
nor U3548 (N_3548,N_43,N_2421);
and U3549 (N_3549,N_993,N_1421);
and U3550 (N_3550,N_1334,N_660);
nor U3551 (N_3551,N_851,N_282);
and U3552 (N_3552,N_699,N_2394);
nor U3553 (N_3553,N_1186,N_2464);
or U3554 (N_3554,N_526,N_1965);
xnor U3555 (N_3555,N_504,N_884);
nand U3556 (N_3556,N_2101,N_2100);
nand U3557 (N_3557,N_803,N_305);
and U3558 (N_3558,N_2422,N_1009);
nand U3559 (N_3559,N_1597,N_983);
nand U3560 (N_3560,N_18,N_1574);
and U3561 (N_3561,N_1784,N_152);
xor U3562 (N_3562,N_1120,N_2385);
and U3563 (N_3563,N_1590,N_4);
or U3564 (N_3564,N_1465,N_248);
xnor U3565 (N_3565,N_2397,N_2154);
and U3566 (N_3566,N_1898,N_2371);
xnor U3567 (N_3567,N_1809,N_1020);
and U3568 (N_3568,N_2353,N_638);
and U3569 (N_3569,N_1476,N_1724);
xnor U3570 (N_3570,N_1723,N_1545);
or U3571 (N_3571,N_1986,N_759);
or U3572 (N_3572,N_1309,N_2345);
and U3573 (N_3573,N_1479,N_118);
nand U3574 (N_3574,N_1554,N_2369);
nor U3575 (N_3575,N_609,N_105);
nand U3576 (N_3576,N_2206,N_1181);
xor U3577 (N_3577,N_2048,N_1264);
xnor U3578 (N_3578,N_2402,N_1042);
nand U3579 (N_3579,N_180,N_755);
nand U3580 (N_3580,N_5,N_234);
nand U3581 (N_3581,N_829,N_228);
nand U3582 (N_3582,N_413,N_2450);
or U3583 (N_3583,N_1350,N_483);
nand U3584 (N_3584,N_1637,N_1262);
nand U3585 (N_3585,N_986,N_718);
or U3586 (N_3586,N_2040,N_17);
or U3587 (N_3587,N_1442,N_1126);
xor U3588 (N_3588,N_2298,N_2388);
nor U3589 (N_3589,N_1821,N_2354);
nor U3590 (N_3590,N_1332,N_1014);
nand U3591 (N_3591,N_549,N_1300);
nand U3592 (N_3592,N_401,N_1276);
nand U3593 (N_3593,N_2082,N_96);
nand U3594 (N_3594,N_1907,N_778);
and U3595 (N_3595,N_724,N_321);
nor U3596 (N_3596,N_1016,N_1504);
nor U3597 (N_3597,N_688,N_1800);
and U3598 (N_3598,N_998,N_2405);
and U3599 (N_3599,N_1274,N_1053);
or U3600 (N_3600,N_367,N_1610);
nor U3601 (N_3601,N_113,N_902);
or U3602 (N_3602,N_239,N_354);
nor U3603 (N_3603,N_1948,N_2295);
nand U3604 (N_3604,N_1182,N_1206);
and U3605 (N_3605,N_765,N_1091);
or U3606 (N_3606,N_399,N_160);
nor U3607 (N_3607,N_690,N_935);
nand U3608 (N_3608,N_1667,N_1894);
and U3609 (N_3609,N_1813,N_434);
nor U3610 (N_3610,N_910,N_1132);
or U3611 (N_3611,N_2209,N_2370);
nand U3612 (N_3612,N_1540,N_87);
or U3613 (N_3613,N_15,N_918);
xnor U3614 (N_3614,N_1691,N_284);
xnor U3615 (N_3615,N_1280,N_1072);
nand U3616 (N_3616,N_1214,N_1002);
nand U3617 (N_3617,N_599,N_2220);
or U3618 (N_3618,N_1136,N_2329);
or U3619 (N_3619,N_1471,N_2062);
and U3620 (N_3620,N_1728,N_828);
and U3621 (N_3621,N_898,N_1401);
nand U3622 (N_3622,N_2165,N_2265);
xnor U3623 (N_3623,N_2459,N_1592);
nor U3624 (N_3624,N_216,N_1224);
nor U3625 (N_3625,N_2277,N_919);
nand U3626 (N_3626,N_178,N_2069);
nor U3627 (N_3627,N_1916,N_451);
and U3628 (N_3628,N_2243,N_1697);
nand U3629 (N_3629,N_1448,N_1311);
or U3630 (N_3630,N_1434,N_1166);
or U3631 (N_3631,N_1773,N_479);
xnor U3632 (N_3632,N_1411,N_2399);
and U3633 (N_3633,N_1461,N_2361);
or U3634 (N_3634,N_817,N_844);
and U3635 (N_3635,N_1110,N_1501);
or U3636 (N_3636,N_873,N_1482);
nand U3637 (N_3637,N_641,N_359);
or U3638 (N_3638,N_1093,N_2413);
nand U3639 (N_3639,N_1844,N_490);
nand U3640 (N_3640,N_388,N_1919);
nand U3641 (N_3641,N_295,N_12);
and U3642 (N_3642,N_2469,N_805);
and U3643 (N_3643,N_1356,N_1629);
and U3644 (N_3644,N_2214,N_1642);
nor U3645 (N_3645,N_1579,N_1336);
nand U3646 (N_3646,N_1012,N_1835);
nand U3647 (N_3647,N_1880,N_1833);
and U3648 (N_3648,N_2030,N_1816);
nor U3649 (N_3649,N_255,N_306);
or U3650 (N_3650,N_1655,N_393);
xnor U3651 (N_3651,N_2324,N_28);
or U3652 (N_3652,N_746,N_1456);
nand U3653 (N_3653,N_1417,N_762);
or U3654 (N_3654,N_347,N_2251);
xor U3655 (N_3655,N_1117,N_591);
and U3656 (N_3656,N_333,N_845);
or U3657 (N_3657,N_1495,N_1777);
or U3658 (N_3658,N_2499,N_2080);
and U3659 (N_3659,N_2244,N_1921);
nand U3660 (N_3660,N_2049,N_2207);
nand U3661 (N_3661,N_1171,N_1480);
nand U3662 (N_3662,N_1532,N_685);
and U3663 (N_3663,N_58,N_2039);
nor U3664 (N_3664,N_1599,N_1749);
nor U3665 (N_3665,N_1052,N_941);
nand U3666 (N_3666,N_1169,N_90);
nand U3667 (N_3667,N_1881,N_163);
and U3668 (N_3668,N_1167,N_119);
and U3669 (N_3669,N_2074,N_1895);
nand U3670 (N_3670,N_485,N_1527);
and U3671 (N_3671,N_895,N_1823);
nor U3672 (N_3672,N_1991,N_991);
xnor U3673 (N_3673,N_2236,N_949);
and U3674 (N_3674,N_1288,N_812);
nor U3675 (N_3675,N_29,N_2460);
nor U3676 (N_3676,N_717,N_2013);
xnor U3677 (N_3677,N_99,N_1876);
or U3678 (N_3678,N_663,N_1296);
or U3679 (N_3679,N_1902,N_2031);
nor U3680 (N_3680,N_1289,N_2412);
nand U3681 (N_3681,N_789,N_878);
and U3682 (N_3682,N_1640,N_1454);
nor U3683 (N_3683,N_2077,N_1964);
and U3684 (N_3684,N_416,N_59);
nor U3685 (N_3685,N_2330,N_1682);
or U3686 (N_3686,N_2073,N_1230);
or U3687 (N_3687,N_1140,N_2096);
nand U3688 (N_3688,N_2363,N_1502);
xor U3689 (N_3689,N_1718,N_2309);
xnor U3690 (N_3690,N_1657,N_93);
nand U3691 (N_3691,N_601,N_2144);
and U3692 (N_3692,N_313,N_208);
or U3693 (N_3693,N_1797,N_13);
nor U3694 (N_3694,N_582,N_441);
nor U3695 (N_3695,N_1112,N_864);
nor U3696 (N_3696,N_1229,N_1235);
nand U3697 (N_3697,N_1094,N_2113);
xnor U3698 (N_3698,N_1980,N_2197);
nand U3699 (N_3699,N_351,N_498);
and U3700 (N_3700,N_906,N_1165);
or U3701 (N_3701,N_1281,N_2474);
and U3702 (N_3702,N_1008,N_1423);
or U3703 (N_3703,N_1573,N_767);
nor U3704 (N_3704,N_1802,N_468);
and U3705 (N_3705,N_1064,N_1680);
or U3706 (N_3706,N_807,N_218);
nand U3707 (N_3707,N_1638,N_55);
xor U3708 (N_3708,N_1418,N_207);
nor U3709 (N_3709,N_1312,N_595);
xor U3710 (N_3710,N_2088,N_995);
and U3711 (N_3711,N_2055,N_1086);
nand U3712 (N_3712,N_2137,N_172);
or U3713 (N_3713,N_1043,N_2185);
and U3714 (N_3714,N_1571,N_1036);
xnor U3715 (N_3715,N_522,N_1287);
or U3716 (N_3716,N_2146,N_42);
nor U3717 (N_3717,N_2410,N_818);
or U3718 (N_3718,N_2011,N_848);
and U3719 (N_3719,N_1562,N_76);
xnor U3720 (N_3720,N_2325,N_2119);
or U3721 (N_3721,N_431,N_540);
nor U3722 (N_3722,N_2213,N_1893);
nor U3723 (N_3723,N_855,N_756);
nor U3724 (N_3724,N_1218,N_325);
xor U3725 (N_3725,N_511,N_1462);
nand U3726 (N_3726,N_1778,N_1769);
xnor U3727 (N_3727,N_1932,N_2294);
nor U3728 (N_3728,N_1819,N_1267);
or U3729 (N_3729,N_710,N_133);
nor U3730 (N_3730,N_2116,N_2444);
nor U3731 (N_3731,N_1606,N_892);
or U3732 (N_3732,N_1658,N_1928);
nand U3733 (N_3733,N_2182,N_1715);
nor U3734 (N_3734,N_303,N_156);
and U3735 (N_3735,N_407,N_1367);
or U3736 (N_3736,N_1934,N_1781);
nand U3737 (N_3737,N_764,N_2267);
or U3738 (N_3738,N_1353,N_2059);
nor U3739 (N_3739,N_1499,N_1698);
nor U3740 (N_3740,N_1413,N_104);
nor U3741 (N_3741,N_1313,N_624);
nand U3742 (N_3742,N_1363,N_1801);
nor U3743 (N_3743,N_356,N_1249);
nand U3744 (N_3744,N_1973,N_1603);
nor U3745 (N_3745,N_2272,N_456);
or U3746 (N_3746,N_2093,N_1516);
nand U3747 (N_3747,N_1672,N_790);
and U3748 (N_3748,N_1408,N_2145);
or U3749 (N_3749,N_360,N_26);
nor U3750 (N_3750,N_2133,N_2056);
or U3751 (N_3751,N_1183,N_2029);
or U3752 (N_3752,N_585,N_360);
and U3753 (N_3753,N_1208,N_683);
nor U3754 (N_3754,N_698,N_509);
and U3755 (N_3755,N_1580,N_158);
xnor U3756 (N_3756,N_1921,N_2494);
or U3757 (N_3757,N_660,N_717);
and U3758 (N_3758,N_232,N_2046);
nand U3759 (N_3759,N_1871,N_2237);
and U3760 (N_3760,N_746,N_1155);
or U3761 (N_3761,N_2204,N_878);
or U3762 (N_3762,N_858,N_2464);
and U3763 (N_3763,N_456,N_972);
and U3764 (N_3764,N_2481,N_430);
nor U3765 (N_3765,N_1545,N_2479);
nand U3766 (N_3766,N_1084,N_854);
and U3767 (N_3767,N_483,N_1736);
or U3768 (N_3768,N_537,N_558);
or U3769 (N_3769,N_1876,N_680);
nor U3770 (N_3770,N_1335,N_897);
or U3771 (N_3771,N_2010,N_1006);
nor U3772 (N_3772,N_2363,N_11);
and U3773 (N_3773,N_385,N_550);
and U3774 (N_3774,N_381,N_418);
nand U3775 (N_3775,N_1801,N_1246);
and U3776 (N_3776,N_1171,N_1505);
or U3777 (N_3777,N_378,N_1267);
or U3778 (N_3778,N_1715,N_629);
and U3779 (N_3779,N_1101,N_1709);
nand U3780 (N_3780,N_2402,N_2134);
nor U3781 (N_3781,N_863,N_1911);
and U3782 (N_3782,N_333,N_2339);
or U3783 (N_3783,N_1888,N_129);
nand U3784 (N_3784,N_1848,N_1454);
nand U3785 (N_3785,N_2466,N_579);
or U3786 (N_3786,N_1632,N_2192);
and U3787 (N_3787,N_763,N_1976);
or U3788 (N_3788,N_298,N_1488);
nor U3789 (N_3789,N_641,N_1628);
or U3790 (N_3790,N_2184,N_1102);
xnor U3791 (N_3791,N_2059,N_729);
or U3792 (N_3792,N_1938,N_2034);
or U3793 (N_3793,N_1979,N_404);
nand U3794 (N_3794,N_37,N_977);
and U3795 (N_3795,N_332,N_2137);
nand U3796 (N_3796,N_2128,N_478);
nand U3797 (N_3797,N_82,N_592);
nand U3798 (N_3798,N_1024,N_2166);
or U3799 (N_3799,N_1239,N_1663);
and U3800 (N_3800,N_1071,N_147);
xor U3801 (N_3801,N_2374,N_1188);
or U3802 (N_3802,N_2269,N_1384);
nor U3803 (N_3803,N_218,N_894);
nor U3804 (N_3804,N_1306,N_217);
nor U3805 (N_3805,N_766,N_2180);
or U3806 (N_3806,N_1396,N_2225);
nor U3807 (N_3807,N_1933,N_2071);
nor U3808 (N_3808,N_2466,N_434);
nand U3809 (N_3809,N_1957,N_1492);
nor U3810 (N_3810,N_316,N_2414);
or U3811 (N_3811,N_78,N_770);
or U3812 (N_3812,N_203,N_1192);
and U3813 (N_3813,N_2399,N_2432);
nand U3814 (N_3814,N_2071,N_1934);
and U3815 (N_3815,N_1822,N_538);
and U3816 (N_3816,N_1334,N_891);
nor U3817 (N_3817,N_624,N_225);
and U3818 (N_3818,N_59,N_1066);
or U3819 (N_3819,N_1290,N_418);
xor U3820 (N_3820,N_64,N_165);
or U3821 (N_3821,N_1263,N_275);
and U3822 (N_3822,N_1703,N_1141);
nand U3823 (N_3823,N_2340,N_813);
xor U3824 (N_3824,N_1036,N_920);
and U3825 (N_3825,N_2172,N_1690);
or U3826 (N_3826,N_853,N_1775);
nand U3827 (N_3827,N_1829,N_1182);
or U3828 (N_3828,N_371,N_2241);
or U3829 (N_3829,N_372,N_1137);
nor U3830 (N_3830,N_2134,N_548);
nand U3831 (N_3831,N_361,N_745);
and U3832 (N_3832,N_1559,N_2421);
xor U3833 (N_3833,N_2294,N_2388);
and U3834 (N_3834,N_93,N_402);
nand U3835 (N_3835,N_478,N_1583);
and U3836 (N_3836,N_271,N_1861);
nor U3837 (N_3837,N_2038,N_649);
or U3838 (N_3838,N_1115,N_2182);
and U3839 (N_3839,N_1218,N_1376);
nor U3840 (N_3840,N_254,N_2447);
nor U3841 (N_3841,N_1357,N_2160);
and U3842 (N_3842,N_1120,N_410);
or U3843 (N_3843,N_342,N_94);
or U3844 (N_3844,N_2333,N_1057);
xnor U3845 (N_3845,N_2462,N_47);
and U3846 (N_3846,N_1513,N_462);
nor U3847 (N_3847,N_504,N_1527);
nand U3848 (N_3848,N_905,N_350);
or U3849 (N_3849,N_1073,N_2153);
nor U3850 (N_3850,N_474,N_109);
and U3851 (N_3851,N_1493,N_409);
or U3852 (N_3852,N_1412,N_2171);
nand U3853 (N_3853,N_1358,N_461);
nor U3854 (N_3854,N_2245,N_1479);
or U3855 (N_3855,N_1136,N_1496);
nand U3856 (N_3856,N_2111,N_1817);
and U3857 (N_3857,N_939,N_2215);
nand U3858 (N_3858,N_855,N_742);
or U3859 (N_3859,N_2349,N_1429);
xnor U3860 (N_3860,N_333,N_1689);
nor U3861 (N_3861,N_1009,N_1131);
nand U3862 (N_3862,N_1907,N_1583);
and U3863 (N_3863,N_2376,N_391);
nor U3864 (N_3864,N_1124,N_1903);
and U3865 (N_3865,N_1515,N_1734);
nor U3866 (N_3866,N_1914,N_1559);
nor U3867 (N_3867,N_1228,N_2260);
nand U3868 (N_3868,N_267,N_649);
nor U3869 (N_3869,N_2410,N_1930);
nor U3870 (N_3870,N_1231,N_452);
or U3871 (N_3871,N_1768,N_964);
nor U3872 (N_3872,N_410,N_860);
nand U3873 (N_3873,N_1613,N_1786);
and U3874 (N_3874,N_1163,N_1442);
nor U3875 (N_3875,N_1349,N_2428);
nand U3876 (N_3876,N_1340,N_2184);
or U3877 (N_3877,N_547,N_2156);
xnor U3878 (N_3878,N_1882,N_79);
nand U3879 (N_3879,N_1668,N_1984);
xnor U3880 (N_3880,N_2380,N_232);
and U3881 (N_3881,N_2400,N_2414);
and U3882 (N_3882,N_2071,N_1036);
or U3883 (N_3883,N_634,N_2339);
or U3884 (N_3884,N_2218,N_693);
or U3885 (N_3885,N_676,N_2190);
and U3886 (N_3886,N_1297,N_395);
xor U3887 (N_3887,N_825,N_1372);
nor U3888 (N_3888,N_711,N_2059);
or U3889 (N_3889,N_503,N_217);
or U3890 (N_3890,N_531,N_1930);
and U3891 (N_3891,N_2203,N_1475);
or U3892 (N_3892,N_1388,N_1269);
or U3893 (N_3893,N_1337,N_1162);
nor U3894 (N_3894,N_317,N_2224);
xor U3895 (N_3895,N_581,N_1788);
xnor U3896 (N_3896,N_2249,N_1394);
and U3897 (N_3897,N_1027,N_99);
nor U3898 (N_3898,N_2096,N_2012);
and U3899 (N_3899,N_2333,N_123);
nor U3900 (N_3900,N_51,N_1332);
or U3901 (N_3901,N_1386,N_1837);
and U3902 (N_3902,N_935,N_1555);
nor U3903 (N_3903,N_2340,N_2448);
nor U3904 (N_3904,N_194,N_514);
nand U3905 (N_3905,N_2190,N_522);
nand U3906 (N_3906,N_960,N_2336);
nand U3907 (N_3907,N_240,N_350);
or U3908 (N_3908,N_1442,N_2374);
or U3909 (N_3909,N_1332,N_2105);
nand U3910 (N_3910,N_844,N_2383);
and U3911 (N_3911,N_377,N_1564);
and U3912 (N_3912,N_1272,N_1748);
nor U3913 (N_3913,N_1761,N_1170);
or U3914 (N_3914,N_2306,N_1866);
nand U3915 (N_3915,N_949,N_1826);
or U3916 (N_3916,N_35,N_2386);
nand U3917 (N_3917,N_2044,N_1392);
and U3918 (N_3918,N_793,N_1385);
nor U3919 (N_3919,N_307,N_980);
nor U3920 (N_3920,N_877,N_1641);
nand U3921 (N_3921,N_231,N_1421);
xor U3922 (N_3922,N_2190,N_2482);
xnor U3923 (N_3923,N_1547,N_1491);
nand U3924 (N_3924,N_572,N_781);
and U3925 (N_3925,N_76,N_1834);
and U3926 (N_3926,N_1323,N_2438);
or U3927 (N_3927,N_2463,N_1472);
nand U3928 (N_3928,N_121,N_1753);
or U3929 (N_3929,N_914,N_1524);
or U3930 (N_3930,N_1264,N_1330);
nand U3931 (N_3931,N_1898,N_350);
nor U3932 (N_3932,N_137,N_205);
nand U3933 (N_3933,N_527,N_881);
nand U3934 (N_3934,N_652,N_618);
and U3935 (N_3935,N_615,N_1039);
or U3936 (N_3936,N_291,N_882);
nor U3937 (N_3937,N_1538,N_1450);
or U3938 (N_3938,N_2122,N_1431);
or U3939 (N_3939,N_943,N_418);
nor U3940 (N_3940,N_1983,N_979);
nand U3941 (N_3941,N_49,N_487);
nor U3942 (N_3942,N_1860,N_1935);
nand U3943 (N_3943,N_2377,N_1080);
or U3944 (N_3944,N_2092,N_1446);
nand U3945 (N_3945,N_148,N_2132);
nor U3946 (N_3946,N_1298,N_2414);
or U3947 (N_3947,N_1619,N_1905);
nor U3948 (N_3948,N_2285,N_164);
nand U3949 (N_3949,N_1103,N_1982);
and U3950 (N_3950,N_593,N_1908);
nor U3951 (N_3951,N_1711,N_1202);
nand U3952 (N_3952,N_255,N_170);
and U3953 (N_3953,N_2184,N_462);
or U3954 (N_3954,N_966,N_1610);
nand U3955 (N_3955,N_144,N_1107);
nor U3956 (N_3956,N_769,N_221);
or U3957 (N_3957,N_788,N_1046);
and U3958 (N_3958,N_1528,N_242);
or U3959 (N_3959,N_432,N_952);
nand U3960 (N_3960,N_57,N_1414);
and U3961 (N_3961,N_174,N_475);
xnor U3962 (N_3962,N_1682,N_2082);
and U3963 (N_3963,N_1701,N_1856);
and U3964 (N_3964,N_2115,N_652);
or U3965 (N_3965,N_1972,N_582);
or U3966 (N_3966,N_1614,N_267);
nor U3967 (N_3967,N_1363,N_84);
nand U3968 (N_3968,N_2113,N_808);
nand U3969 (N_3969,N_2200,N_855);
nand U3970 (N_3970,N_2170,N_1114);
or U3971 (N_3971,N_1751,N_855);
and U3972 (N_3972,N_1968,N_186);
xor U3973 (N_3973,N_2357,N_1025);
or U3974 (N_3974,N_758,N_2424);
and U3975 (N_3975,N_1423,N_996);
nand U3976 (N_3976,N_1894,N_1006);
or U3977 (N_3977,N_2450,N_1690);
or U3978 (N_3978,N_1666,N_224);
or U3979 (N_3979,N_132,N_1715);
and U3980 (N_3980,N_926,N_541);
nor U3981 (N_3981,N_1324,N_780);
xor U3982 (N_3982,N_2140,N_1650);
nor U3983 (N_3983,N_1119,N_1983);
or U3984 (N_3984,N_1274,N_611);
nor U3985 (N_3985,N_1542,N_2289);
and U3986 (N_3986,N_804,N_82);
or U3987 (N_3987,N_2047,N_1265);
nand U3988 (N_3988,N_908,N_2122);
nor U3989 (N_3989,N_812,N_670);
and U3990 (N_3990,N_153,N_2492);
nor U3991 (N_3991,N_1587,N_1351);
or U3992 (N_3992,N_2031,N_1229);
nor U3993 (N_3993,N_1172,N_1278);
nor U3994 (N_3994,N_220,N_1811);
nor U3995 (N_3995,N_2215,N_1269);
and U3996 (N_3996,N_1464,N_613);
and U3997 (N_3997,N_195,N_189);
nor U3998 (N_3998,N_1523,N_182);
or U3999 (N_3999,N_1862,N_2279);
or U4000 (N_4000,N_1880,N_2154);
and U4001 (N_4001,N_445,N_1354);
nor U4002 (N_4002,N_504,N_1100);
nand U4003 (N_4003,N_2475,N_1668);
nand U4004 (N_4004,N_30,N_635);
nand U4005 (N_4005,N_344,N_1321);
or U4006 (N_4006,N_1299,N_1875);
xor U4007 (N_4007,N_2253,N_1507);
or U4008 (N_4008,N_1496,N_1541);
or U4009 (N_4009,N_1115,N_990);
or U4010 (N_4010,N_629,N_2146);
nor U4011 (N_4011,N_2021,N_1350);
nand U4012 (N_4012,N_133,N_1490);
nor U4013 (N_4013,N_1994,N_713);
nand U4014 (N_4014,N_1706,N_656);
nand U4015 (N_4015,N_212,N_583);
nand U4016 (N_4016,N_205,N_484);
or U4017 (N_4017,N_607,N_918);
nand U4018 (N_4018,N_2053,N_868);
and U4019 (N_4019,N_2057,N_1410);
nor U4020 (N_4020,N_868,N_2064);
nor U4021 (N_4021,N_2163,N_373);
or U4022 (N_4022,N_1776,N_1245);
or U4023 (N_4023,N_2384,N_1026);
nand U4024 (N_4024,N_957,N_2021);
nor U4025 (N_4025,N_375,N_721);
or U4026 (N_4026,N_1674,N_2360);
and U4027 (N_4027,N_644,N_937);
nand U4028 (N_4028,N_2333,N_833);
and U4029 (N_4029,N_1486,N_2329);
nor U4030 (N_4030,N_18,N_68);
nor U4031 (N_4031,N_611,N_1298);
and U4032 (N_4032,N_1807,N_411);
and U4033 (N_4033,N_1824,N_1390);
nand U4034 (N_4034,N_868,N_1641);
nand U4035 (N_4035,N_843,N_1131);
or U4036 (N_4036,N_340,N_1676);
nor U4037 (N_4037,N_1584,N_1778);
nand U4038 (N_4038,N_2149,N_1343);
nand U4039 (N_4039,N_958,N_537);
and U4040 (N_4040,N_442,N_1866);
and U4041 (N_4041,N_128,N_601);
or U4042 (N_4042,N_1322,N_2341);
or U4043 (N_4043,N_299,N_460);
xnor U4044 (N_4044,N_2140,N_830);
nor U4045 (N_4045,N_1340,N_1991);
and U4046 (N_4046,N_458,N_1425);
or U4047 (N_4047,N_2097,N_1322);
nor U4048 (N_4048,N_2308,N_1112);
or U4049 (N_4049,N_1675,N_1777);
xor U4050 (N_4050,N_2139,N_371);
nor U4051 (N_4051,N_871,N_1954);
and U4052 (N_4052,N_163,N_148);
or U4053 (N_4053,N_1791,N_938);
or U4054 (N_4054,N_1784,N_1671);
nor U4055 (N_4055,N_757,N_133);
nor U4056 (N_4056,N_1112,N_2052);
xnor U4057 (N_4057,N_973,N_2331);
nand U4058 (N_4058,N_2081,N_2497);
and U4059 (N_4059,N_393,N_1209);
and U4060 (N_4060,N_592,N_2180);
or U4061 (N_4061,N_1289,N_1255);
nand U4062 (N_4062,N_1480,N_598);
or U4063 (N_4063,N_406,N_1792);
and U4064 (N_4064,N_580,N_43);
nand U4065 (N_4065,N_1204,N_944);
xor U4066 (N_4066,N_456,N_887);
and U4067 (N_4067,N_1577,N_2234);
nand U4068 (N_4068,N_1706,N_1998);
or U4069 (N_4069,N_1827,N_2337);
or U4070 (N_4070,N_1989,N_374);
nand U4071 (N_4071,N_596,N_299);
nor U4072 (N_4072,N_87,N_1735);
nor U4073 (N_4073,N_919,N_2470);
xnor U4074 (N_4074,N_2451,N_1243);
and U4075 (N_4075,N_389,N_1084);
or U4076 (N_4076,N_1200,N_24);
and U4077 (N_4077,N_2225,N_2270);
nor U4078 (N_4078,N_1458,N_2097);
or U4079 (N_4079,N_1217,N_1497);
nor U4080 (N_4080,N_932,N_1735);
nand U4081 (N_4081,N_1089,N_1364);
and U4082 (N_4082,N_1988,N_1967);
and U4083 (N_4083,N_85,N_810);
xor U4084 (N_4084,N_979,N_988);
or U4085 (N_4085,N_2033,N_2353);
and U4086 (N_4086,N_266,N_1389);
and U4087 (N_4087,N_2485,N_2209);
and U4088 (N_4088,N_1643,N_1577);
nor U4089 (N_4089,N_42,N_2458);
and U4090 (N_4090,N_987,N_2052);
nand U4091 (N_4091,N_155,N_656);
nand U4092 (N_4092,N_78,N_330);
xor U4093 (N_4093,N_1293,N_846);
nand U4094 (N_4094,N_915,N_2069);
or U4095 (N_4095,N_226,N_1832);
xor U4096 (N_4096,N_1425,N_432);
or U4097 (N_4097,N_1813,N_802);
nor U4098 (N_4098,N_254,N_518);
nor U4099 (N_4099,N_1539,N_1826);
and U4100 (N_4100,N_2284,N_425);
xor U4101 (N_4101,N_188,N_2352);
and U4102 (N_4102,N_1205,N_1988);
and U4103 (N_4103,N_1178,N_1727);
nor U4104 (N_4104,N_724,N_2091);
nor U4105 (N_4105,N_589,N_330);
and U4106 (N_4106,N_628,N_357);
nor U4107 (N_4107,N_92,N_1386);
nor U4108 (N_4108,N_2253,N_1733);
nand U4109 (N_4109,N_798,N_554);
nor U4110 (N_4110,N_314,N_1074);
nor U4111 (N_4111,N_1612,N_669);
nor U4112 (N_4112,N_576,N_2157);
and U4113 (N_4113,N_1933,N_173);
xor U4114 (N_4114,N_1288,N_82);
nor U4115 (N_4115,N_2436,N_1498);
or U4116 (N_4116,N_219,N_2257);
or U4117 (N_4117,N_2158,N_317);
xnor U4118 (N_4118,N_550,N_2114);
nand U4119 (N_4119,N_1107,N_1817);
nor U4120 (N_4120,N_483,N_1715);
and U4121 (N_4121,N_1848,N_1024);
and U4122 (N_4122,N_2315,N_230);
xor U4123 (N_4123,N_967,N_601);
xnor U4124 (N_4124,N_671,N_2418);
nand U4125 (N_4125,N_531,N_424);
or U4126 (N_4126,N_1806,N_2391);
or U4127 (N_4127,N_2493,N_2143);
nor U4128 (N_4128,N_1362,N_65);
and U4129 (N_4129,N_1097,N_574);
nor U4130 (N_4130,N_2054,N_1130);
or U4131 (N_4131,N_688,N_2181);
nor U4132 (N_4132,N_1538,N_1051);
and U4133 (N_4133,N_516,N_1615);
or U4134 (N_4134,N_1094,N_115);
nand U4135 (N_4135,N_795,N_1689);
and U4136 (N_4136,N_1579,N_657);
or U4137 (N_4137,N_515,N_1167);
nand U4138 (N_4138,N_1401,N_1571);
and U4139 (N_4139,N_1051,N_808);
or U4140 (N_4140,N_1736,N_1741);
nor U4141 (N_4141,N_198,N_429);
xnor U4142 (N_4142,N_1863,N_32);
nor U4143 (N_4143,N_138,N_1348);
nand U4144 (N_4144,N_138,N_174);
or U4145 (N_4145,N_1851,N_830);
nand U4146 (N_4146,N_576,N_1843);
nand U4147 (N_4147,N_657,N_961);
and U4148 (N_4148,N_701,N_808);
nor U4149 (N_4149,N_2423,N_1108);
nand U4150 (N_4150,N_2398,N_296);
nor U4151 (N_4151,N_1019,N_686);
nand U4152 (N_4152,N_750,N_112);
nor U4153 (N_4153,N_181,N_865);
nor U4154 (N_4154,N_1696,N_447);
and U4155 (N_4155,N_294,N_1380);
nand U4156 (N_4156,N_2389,N_1625);
and U4157 (N_4157,N_1829,N_622);
nand U4158 (N_4158,N_450,N_206);
nand U4159 (N_4159,N_1647,N_515);
and U4160 (N_4160,N_999,N_1880);
and U4161 (N_4161,N_2140,N_2471);
nor U4162 (N_4162,N_931,N_1611);
xnor U4163 (N_4163,N_477,N_718);
or U4164 (N_4164,N_1935,N_1591);
and U4165 (N_4165,N_1837,N_1087);
xor U4166 (N_4166,N_810,N_1537);
and U4167 (N_4167,N_1097,N_447);
nor U4168 (N_4168,N_2004,N_1502);
nand U4169 (N_4169,N_1568,N_688);
or U4170 (N_4170,N_1636,N_1127);
and U4171 (N_4171,N_1373,N_977);
or U4172 (N_4172,N_1985,N_1080);
and U4173 (N_4173,N_1004,N_1619);
and U4174 (N_4174,N_1333,N_2273);
or U4175 (N_4175,N_2176,N_1333);
nor U4176 (N_4176,N_997,N_1733);
and U4177 (N_4177,N_2005,N_1618);
nor U4178 (N_4178,N_2193,N_1991);
and U4179 (N_4179,N_2483,N_387);
and U4180 (N_4180,N_1920,N_1434);
or U4181 (N_4181,N_1309,N_771);
nand U4182 (N_4182,N_2092,N_1582);
nor U4183 (N_4183,N_1271,N_1766);
and U4184 (N_4184,N_1013,N_2018);
nand U4185 (N_4185,N_2264,N_1512);
or U4186 (N_4186,N_1470,N_814);
nand U4187 (N_4187,N_1036,N_1762);
or U4188 (N_4188,N_765,N_773);
nand U4189 (N_4189,N_1760,N_1578);
nand U4190 (N_4190,N_450,N_75);
and U4191 (N_4191,N_77,N_1061);
nand U4192 (N_4192,N_1318,N_294);
and U4193 (N_4193,N_1391,N_376);
nor U4194 (N_4194,N_49,N_101);
nand U4195 (N_4195,N_1421,N_2429);
and U4196 (N_4196,N_841,N_2161);
or U4197 (N_4197,N_206,N_2463);
xor U4198 (N_4198,N_563,N_1207);
and U4199 (N_4199,N_1563,N_563);
nor U4200 (N_4200,N_1826,N_2488);
nor U4201 (N_4201,N_15,N_2276);
xor U4202 (N_4202,N_576,N_215);
or U4203 (N_4203,N_2382,N_767);
and U4204 (N_4204,N_409,N_843);
xnor U4205 (N_4205,N_389,N_1960);
xor U4206 (N_4206,N_1,N_1962);
nor U4207 (N_4207,N_1173,N_1996);
nor U4208 (N_4208,N_362,N_1682);
or U4209 (N_4209,N_1220,N_1532);
and U4210 (N_4210,N_1115,N_1328);
nor U4211 (N_4211,N_1836,N_2169);
and U4212 (N_4212,N_2320,N_1491);
or U4213 (N_4213,N_1332,N_1974);
and U4214 (N_4214,N_496,N_55);
and U4215 (N_4215,N_346,N_726);
and U4216 (N_4216,N_1040,N_1780);
and U4217 (N_4217,N_294,N_1669);
nand U4218 (N_4218,N_1654,N_678);
xnor U4219 (N_4219,N_1464,N_2460);
or U4220 (N_4220,N_1907,N_294);
nand U4221 (N_4221,N_841,N_1789);
nor U4222 (N_4222,N_758,N_890);
or U4223 (N_4223,N_1220,N_689);
nand U4224 (N_4224,N_1506,N_1155);
or U4225 (N_4225,N_171,N_62);
nor U4226 (N_4226,N_1448,N_1326);
nand U4227 (N_4227,N_2325,N_1147);
and U4228 (N_4228,N_1753,N_1495);
and U4229 (N_4229,N_2205,N_161);
or U4230 (N_4230,N_1392,N_1847);
nor U4231 (N_4231,N_1910,N_51);
and U4232 (N_4232,N_922,N_1058);
nand U4233 (N_4233,N_201,N_2407);
xnor U4234 (N_4234,N_1403,N_2396);
nor U4235 (N_4235,N_390,N_936);
and U4236 (N_4236,N_2114,N_785);
or U4237 (N_4237,N_2464,N_2277);
and U4238 (N_4238,N_515,N_1155);
nor U4239 (N_4239,N_2347,N_112);
or U4240 (N_4240,N_623,N_1463);
nand U4241 (N_4241,N_1446,N_1128);
or U4242 (N_4242,N_2195,N_1473);
nand U4243 (N_4243,N_1772,N_473);
nand U4244 (N_4244,N_98,N_1570);
and U4245 (N_4245,N_873,N_351);
and U4246 (N_4246,N_957,N_1307);
or U4247 (N_4247,N_469,N_1970);
and U4248 (N_4248,N_1036,N_1696);
xor U4249 (N_4249,N_1373,N_1392);
nand U4250 (N_4250,N_2072,N_1170);
and U4251 (N_4251,N_852,N_1965);
and U4252 (N_4252,N_453,N_179);
and U4253 (N_4253,N_686,N_2195);
nor U4254 (N_4254,N_671,N_336);
nand U4255 (N_4255,N_573,N_2465);
nor U4256 (N_4256,N_2064,N_2414);
xor U4257 (N_4257,N_1810,N_1813);
xor U4258 (N_4258,N_1950,N_2438);
and U4259 (N_4259,N_567,N_1335);
xor U4260 (N_4260,N_520,N_420);
nand U4261 (N_4261,N_1741,N_51);
nand U4262 (N_4262,N_1275,N_1903);
nor U4263 (N_4263,N_2074,N_478);
nand U4264 (N_4264,N_1449,N_1939);
xnor U4265 (N_4265,N_376,N_1160);
nand U4266 (N_4266,N_1570,N_565);
nand U4267 (N_4267,N_951,N_1257);
or U4268 (N_4268,N_1384,N_418);
nand U4269 (N_4269,N_2208,N_2046);
nand U4270 (N_4270,N_2458,N_2195);
nor U4271 (N_4271,N_611,N_229);
and U4272 (N_4272,N_71,N_517);
or U4273 (N_4273,N_1128,N_493);
nand U4274 (N_4274,N_1161,N_868);
nand U4275 (N_4275,N_2457,N_1015);
nor U4276 (N_4276,N_2279,N_2261);
and U4277 (N_4277,N_1127,N_1104);
nand U4278 (N_4278,N_1402,N_1632);
or U4279 (N_4279,N_1096,N_2337);
nor U4280 (N_4280,N_241,N_835);
nor U4281 (N_4281,N_971,N_245);
and U4282 (N_4282,N_1539,N_1034);
nor U4283 (N_4283,N_1509,N_552);
nor U4284 (N_4284,N_1180,N_1115);
nor U4285 (N_4285,N_1033,N_116);
or U4286 (N_4286,N_2102,N_449);
or U4287 (N_4287,N_1448,N_1928);
xnor U4288 (N_4288,N_1896,N_1416);
and U4289 (N_4289,N_2187,N_346);
and U4290 (N_4290,N_1634,N_1230);
and U4291 (N_4291,N_1428,N_290);
and U4292 (N_4292,N_1425,N_2121);
or U4293 (N_4293,N_2181,N_1037);
nor U4294 (N_4294,N_2188,N_289);
xor U4295 (N_4295,N_2367,N_576);
nand U4296 (N_4296,N_253,N_1573);
and U4297 (N_4297,N_539,N_410);
nand U4298 (N_4298,N_971,N_766);
nor U4299 (N_4299,N_1110,N_1548);
or U4300 (N_4300,N_623,N_306);
nand U4301 (N_4301,N_1055,N_1585);
nor U4302 (N_4302,N_1367,N_1916);
and U4303 (N_4303,N_256,N_637);
nand U4304 (N_4304,N_2048,N_1881);
and U4305 (N_4305,N_1250,N_19);
nand U4306 (N_4306,N_827,N_1541);
and U4307 (N_4307,N_704,N_335);
or U4308 (N_4308,N_583,N_429);
and U4309 (N_4309,N_1624,N_1947);
nand U4310 (N_4310,N_430,N_840);
and U4311 (N_4311,N_1429,N_1644);
or U4312 (N_4312,N_1853,N_2166);
nand U4313 (N_4313,N_166,N_1522);
nand U4314 (N_4314,N_244,N_245);
and U4315 (N_4315,N_966,N_1570);
or U4316 (N_4316,N_600,N_239);
and U4317 (N_4317,N_2461,N_1129);
nand U4318 (N_4318,N_774,N_2356);
xor U4319 (N_4319,N_2220,N_1715);
or U4320 (N_4320,N_407,N_2362);
nand U4321 (N_4321,N_673,N_2136);
nand U4322 (N_4322,N_1855,N_975);
and U4323 (N_4323,N_2226,N_2340);
nor U4324 (N_4324,N_2236,N_135);
nand U4325 (N_4325,N_1021,N_2447);
and U4326 (N_4326,N_2115,N_367);
nor U4327 (N_4327,N_537,N_989);
nor U4328 (N_4328,N_1998,N_2134);
nand U4329 (N_4329,N_73,N_2015);
and U4330 (N_4330,N_315,N_2407);
nand U4331 (N_4331,N_2184,N_821);
nand U4332 (N_4332,N_1091,N_585);
and U4333 (N_4333,N_1497,N_1381);
and U4334 (N_4334,N_1515,N_2298);
nand U4335 (N_4335,N_1154,N_774);
nand U4336 (N_4336,N_1734,N_2112);
nand U4337 (N_4337,N_915,N_224);
nor U4338 (N_4338,N_594,N_2485);
or U4339 (N_4339,N_159,N_2365);
xnor U4340 (N_4340,N_2200,N_835);
and U4341 (N_4341,N_1107,N_549);
or U4342 (N_4342,N_677,N_614);
or U4343 (N_4343,N_1388,N_1449);
nand U4344 (N_4344,N_489,N_2428);
and U4345 (N_4345,N_1860,N_584);
nand U4346 (N_4346,N_2033,N_1355);
nor U4347 (N_4347,N_109,N_2350);
or U4348 (N_4348,N_274,N_204);
nand U4349 (N_4349,N_155,N_152);
nand U4350 (N_4350,N_185,N_2324);
or U4351 (N_4351,N_2417,N_1651);
xnor U4352 (N_4352,N_847,N_1967);
nand U4353 (N_4353,N_1107,N_1386);
nand U4354 (N_4354,N_1837,N_2245);
and U4355 (N_4355,N_124,N_1914);
nor U4356 (N_4356,N_1585,N_873);
xor U4357 (N_4357,N_1658,N_2287);
nor U4358 (N_4358,N_529,N_338);
or U4359 (N_4359,N_618,N_1594);
or U4360 (N_4360,N_922,N_1882);
or U4361 (N_4361,N_734,N_88);
and U4362 (N_4362,N_731,N_332);
or U4363 (N_4363,N_1801,N_1231);
nand U4364 (N_4364,N_1899,N_1837);
or U4365 (N_4365,N_438,N_35);
and U4366 (N_4366,N_1188,N_2325);
nand U4367 (N_4367,N_1591,N_324);
or U4368 (N_4368,N_1381,N_1298);
and U4369 (N_4369,N_778,N_826);
and U4370 (N_4370,N_1226,N_2483);
nand U4371 (N_4371,N_2365,N_972);
or U4372 (N_4372,N_722,N_1283);
and U4373 (N_4373,N_37,N_368);
and U4374 (N_4374,N_1477,N_905);
or U4375 (N_4375,N_295,N_2215);
nor U4376 (N_4376,N_2077,N_193);
and U4377 (N_4377,N_880,N_723);
and U4378 (N_4378,N_1213,N_743);
and U4379 (N_4379,N_68,N_1522);
and U4380 (N_4380,N_225,N_930);
nand U4381 (N_4381,N_1228,N_1265);
nand U4382 (N_4382,N_22,N_519);
nand U4383 (N_4383,N_2211,N_867);
nor U4384 (N_4384,N_2186,N_697);
or U4385 (N_4385,N_2330,N_874);
nor U4386 (N_4386,N_1841,N_2463);
nand U4387 (N_4387,N_278,N_2012);
nor U4388 (N_4388,N_1119,N_2139);
nor U4389 (N_4389,N_2377,N_1508);
nand U4390 (N_4390,N_192,N_2140);
nor U4391 (N_4391,N_174,N_1232);
or U4392 (N_4392,N_2161,N_2304);
or U4393 (N_4393,N_1728,N_1771);
or U4394 (N_4394,N_2264,N_2378);
and U4395 (N_4395,N_1425,N_501);
nand U4396 (N_4396,N_2214,N_944);
nand U4397 (N_4397,N_2414,N_2489);
or U4398 (N_4398,N_227,N_30);
and U4399 (N_4399,N_1337,N_721);
nor U4400 (N_4400,N_2483,N_231);
xnor U4401 (N_4401,N_166,N_1495);
or U4402 (N_4402,N_1117,N_2093);
nand U4403 (N_4403,N_901,N_288);
nor U4404 (N_4404,N_983,N_2357);
nor U4405 (N_4405,N_52,N_1765);
and U4406 (N_4406,N_2198,N_1937);
xor U4407 (N_4407,N_1732,N_890);
and U4408 (N_4408,N_1888,N_854);
nor U4409 (N_4409,N_979,N_68);
nand U4410 (N_4410,N_729,N_1918);
nand U4411 (N_4411,N_485,N_476);
nand U4412 (N_4412,N_1427,N_1380);
nor U4413 (N_4413,N_1889,N_119);
and U4414 (N_4414,N_1430,N_944);
and U4415 (N_4415,N_873,N_2277);
or U4416 (N_4416,N_2454,N_60);
nor U4417 (N_4417,N_820,N_1035);
or U4418 (N_4418,N_1595,N_1684);
and U4419 (N_4419,N_2333,N_857);
nand U4420 (N_4420,N_2070,N_1654);
and U4421 (N_4421,N_1456,N_2106);
nor U4422 (N_4422,N_603,N_79);
or U4423 (N_4423,N_1605,N_703);
nor U4424 (N_4424,N_152,N_2272);
or U4425 (N_4425,N_1109,N_778);
or U4426 (N_4426,N_1714,N_74);
nor U4427 (N_4427,N_2372,N_205);
nor U4428 (N_4428,N_1843,N_2452);
or U4429 (N_4429,N_459,N_2045);
nand U4430 (N_4430,N_361,N_172);
nor U4431 (N_4431,N_1117,N_392);
nand U4432 (N_4432,N_921,N_502);
or U4433 (N_4433,N_384,N_467);
nor U4434 (N_4434,N_436,N_852);
and U4435 (N_4435,N_432,N_2475);
nand U4436 (N_4436,N_23,N_217);
or U4437 (N_4437,N_227,N_253);
or U4438 (N_4438,N_789,N_1414);
nor U4439 (N_4439,N_356,N_887);
nand U4440 (N_4440,N_844,N_2435);
and U4441 (N_4441,N_1779,N_1195);
nand U4442 (N_4442,N_169,N_1520);
nand U4443 (N_4443,N_576,N_1605);
nand U4444 (N_4444,N_782,N_1590);
and U4445 (N_4445,N_1404,N_1448);
nor U4446 (N_4446,N_2120,N_1284);
and U4447 (N_4447,N_2430,N_2367);
or U4448 (N_4448,N_1065,N_1300);
or U4449 (N_4449,N_1187,N_1378);
and U4450 (N_4450,N_1963,N_1829);
nand U4451 (N_4451,N_676,N_704);
xor U4452 (N_4452,N_2441,N_1240);
nor U4453 (N_4453,N_1700,N_1637);
or U4454 (N_4454,N_1460,N_363);
nor U4455 (N_4455,N_1774,N_2486);
nor U4456 (N_4456,N_1789,N_900);
or U4457 (N_4457,N_67,N_466);
nand U4458 (N_4458,N_664,N_2023);
xnor U4459 (N_4459,N_1101,N_494);
nor U4460 (N_4460,N_476,N_1730);
or U4461 (N_4461,N_2416,N_1938);
and U4462 (N_4462,N_442,N_554);
nor U4463 (N_4463,N_2097,N_336);
and U4464 (N_4464,N_1997,N_862);
nor U4465 (N_4465,N_558,N_821);
nand U4466 (N_4466,N_2394,N_1061);
and U4467 (N_4467,N_1907,N_354);
nor U4468 (N_4468,N_1790,N_1245);
nand U4469 (N_4469,N_803,N_2018);
or U4470 (N_4470,N_336,N_1136);
nor U4471 (N_4471,N_1472,N_2395);
nor U4472 (N_4472,N_1625,N_964);
nand U4473 (N_4473,N_849,N_414);
and U4474 (N_4474,N_666,N_84);
nand U4475 (N_4475,N_626,N_820);
or U4476 (N_4476,N_31,N_928);
xor U4477 (N_4477,N_1664,N_1127);
or U4478 (N_4478,N_1266,N_1085);
or U4479 (N_4479,N_897,N_156);
nand U4480 (N_4480,N_1382,N_745);
xor U4481 (N_4481,N_762,N_275);
and U4482 (N_4482,N_1531,N_617);
nor U4483 (N_4483,N_794,N_514);
xor U4484 (N_4484,N_43,N_1070);
and U4485 (N_4485,N_1002,N_431);
nand U4486 (N_4486,N_1290,N_1276);
or U4487 (N_4487,N_2389,N_2079);
nor U4488 (N_4488,N_935,N_2433);
nor U4489 (N_4489,N_1406,N_721);
and U4490 (N_4490,N_1378,N_58);
or U4491 (N_4491,N_2084,N_96);
nand U4492 (N_4492,N_1184,N_2039);
nor U4493 (N_4493,N_1916,N_1520);
nor U4494 (N_4494,N_1831,N_451);
nand U4495 (N_4495,N_579,N_2478);
nand U4496 (N_4496,N_2211,N_1440);
and U4497 (N_4497,N_1299,N_2208);
xnor U4498 (N_4498,N_389,N_1971);
or U4499 (N_4499,N_1833,N_2016);
nand U4500 (N_4500,N_208,N_978);
nand U4501 (N_4501,N_1213,N_1638);
or U4502 (N_4502,N_569,N_2112);
nand U4503 (N_4503,N_395,N_1040);
or U4504 (N_4504,N_186,N_1476);
or U4505 (N_4505,N_200,N_542);
xnor U4506 (N_4506,N_2116,N_1188);
nand U4507 (N_4507,N_827,N_182);
nand U4508 (N_4508,N_2481,N_1014);
xnor U4509 (N_4509,N_1172,N_802);
or U4510 (N_4510,N_2437,N_95);
nor U4511 (N_4511,N_1631,N_813);
nor U4512 (N_4512,N_408,N_217);
nor U4513 (N_4513,N_437,N_630);
nand U4514 (N_4514,N_937,N_1116);
nand U4515 (N_4515,N_709,N_374);
nor U4516 (N_4516,N_39,N_1130);
and U4517 (N_4517,N_1772,N_264);
and U4518 (N_4518,N_1812,N_1818);
and U4519 (N_4519,N_1492,N_2242);
nor U4520 (N_4520,N_123,N_2132);
and U4521 (N_4521,N_2314,N_377);
and U4522 (N_4522,N_574,N_864);
nand U4523 (N_4523,N_2107,N_218);
or U4524 (N_4524,N_1262,N_279);
nand U4525 (N_4525,N_1807,N_2231);
or U4526 (N_4526,N_1976,N_1445);
or U4527 (N_4527,N_586,N_895);
nand U4528 (N_4528,N_2116,N_2064);
nand U4529 (N_4529,N_1916,N_203);
or U4530 (N_4530,N_1855,N_255);
xnor U4531 (N_4531,N_1895,N_195);
nor U4532 (N_4532,N_1832,N_1607);
and U4533 (N_4533,N_1120,N_384);
nor U4534 (N_4534,N_1513,N_1821);
nand U4535 (N_4535,N_845,N_999);
xnor U4536 (N_4536,N_1768,N_44);
and U4537 (N_4537,N_2406,N_504);
or U4538 (N_4538,N_2060,N_425);
or U4539 (N_4539,N_2181,N_1389);
and U4540 (N_4540,N_640,N_895);
nor U4541 (N_4541,N_1145,N_1338);
xor U4542 (N_4542,N_1588,N_1721);
or U4543 (N_4543,N_1921,N_1145);
nand U4544 (N_4544,N_1239,N_959);
nand U4545 (N_4545,N_554,N_233);
nand U4546 (N_4546,N_349,N_1194);
or U4547 (N_4547,N_1090,N_1635);
xnor U4548 (N_4548,N_1623,N_2326);
and U4549 (N_4549,N_1866,N_1757);
nor U4550 (N_4550,N_2252,N_1840);
nand U4551 (N_4551,N_1626,N_800);
and U4552 (N_4552,N_1855,N_1353);
xor U4553 (N_4553,N_2282,N_1981);
nor U4554 (N_4554,N_1989,N_1827);
or U4555 (N_4555,N_1164,N_98);
nor U4556 (N_4556,N_1025,N_680);
xnor U4557 (N_4557,N_573,N_2257);
nand U4558 (N_4558,N_1245,N_1164);
nor U4559 (N_4559,N_1705,N_207);
nor U4560 (N_4560,N_1665,N_329);
or U4561 (N_4561,N_2246,N_1256);
nor U4562 (N_4562,N_1208,N_811);
and U4563 (N_4563,N_1907,N_951);
xor U4564 (N_4564,N_91,N_1386);
or U4565 (N_4565,N_2274,N_1755);
nand U4566 (N_4566,N_914,N_1919);
nor U4567 (N_4567,N_129,N_1120);
nand U4568 (N_4568,N_1978,N_87);
or U4569 (N_4569,N_234,N_1497);
xnor U4570 (N_4570,N_2211,N_1446);
or U4571 (N_4571,N_1053,N_614);
or U4572 (N_4572,N_1196,N_2132);
nand U4573 (N_4573,N_2076,N_2377);
nand U4574 (N_4574,N_734,N_51);
or U4575 (N_4575,N_948,N_1218);
nor U4576 (N_4576,N_1396,N_1758);
nand U4577 (N_4577,N_707,N_431);
nor U4578 (N_4578,N_537,N_276);
and U4579 (N_4579,N_321,N_960);
and U4580 (N_4580,N_516,N_847);
nor U4581 (N_4581,N_1963,N_32);
nand U4582 (N_4582,N_976,N_532);
or U4583 (N_4583,N_1269,N_1463);
and U4584 (N_4584,N_1317,N_2260);
or U4585 (N_4585,N_258,N_2184);
xnor U4586 (N_4586,N_492,N_2062);
nand U4587 (N_4587,N_1849,N_1298);
and U4588 (N_4588,N_2066,N_2242);
and U4589 (N_4589,N_2350,N_1278);
nand U4590 (N_4590,N_281,N_1003);
nand U4591 (N_4591,N_1686,N_2063);
and U4592 (N_4592,N_1760,N_2008);
and U4593 (N_4593,N_857,N_1523);
nand U4594 (N_4594,N_1461,N_2042);
nand U4595 (N_4595,N_695,N_2201);
xnor U4596 (N_4596,N_2185,N_878);
and U4597 (N_4597,N_2083,N_1146);
nor U4598 (N_4598,N_1293,N_375);
and U4599 (N_4599,N_1061,N_1592);
or U4600 (N_4600,N_2194,N_789);
nor U4601 (N_4601,N_400,N_71);
or U4602 (N_4602,N_276,N_1419);
nor U4603 (N_4603,N_1605,N_456);
and U4604 (N_4604,N_168,N_1026);
or U4605 (N_4605,N_1319,N_241);
nand U4606 (N_4606,N_264,N_2249);
nand U4607 (N_4607,N_1653,N_50);
xor U4608 (N_4608,N_2383,N_1355);
nor U4609 (N_4609,N_783,N_934);
and U4610 (N_4610,N_2090,N_1263);
and U4611 (N_4611,N_2401,N_1963);
and U4612 (N_4612,N_1504,N_319);
nor U4613 (N_4613,N_218,N_129);
nand U4614 (N_4614,N_2455,N_1414);
nor U4615 (N_4615,N_1777,N_442);
or U4616 (N_4616,N_1551,N_392);
and U4617 (N_4617,N_2085,N_1388);
nand U4618 (N_4618,N_2425,N_447);
nand U4619 (N_4619,N_1165,N_2342);
nand U4620 (N_4620,N_2442,N_413);
nand U4621 (N_4621,N_1975,N_855);
and U4622 (N_4622,N_161,N_1187);
nand U4623 (N_4623,N_216,N_551);
or U4624 (N_4624,N_1326,N_796);
nor U4625 (N_4625,N_536,N_1469);
or U4626 (N_4626,N_1748,N_493);
nor U4627 (N_4627,N_652,N_2295);
nor U4628 (N_4628,N_649,N_1452);
nor U4629 (N_4629,N_575,N_1200);
or U4630 (N_4630,N_398,N_8);
nand U4631 (N_4631,N_1990,N_2107);
nor U4632 (N_4632,N_649,N_1940);
or U4633 (N_4633,N_1727,N_739);
or U4634 (N_4634,N_1701,N_1899);
nand U4635 (N_4635,N_1802,N_1199);
and U4636 (N_4636,N_857,N_1403);
nor U4637 (N_4637,N_888,N_856);
nand U4638 (N_4638,N_2243,N_122);
or U4639 (N_4639,N_2331,N_1080);
xor U4640 (N_4640,N_1093,N_59);
or U4641 (N_4641,N_1790,N_89);
or U4642 (N_4642,N_231,N_2144);
nor U4643 (N_4643,N_204,N_1302);
nand U4644 (N_4644,N_2476,N_2156);
and U4645 (N_4645,N_1275,N_2437);
nor U4646 (N_4646,N_2327,N_1822);
nor U4647 (N_4647,N_2217,N_1267);
or U4648 (N_4648,N_2414,N_1485);
or U4649 (N_4649,N_904,N_936);
nor U4650 (N_4650,N_851,N_1009);
or U4651 (N_4651,N_1099,N_1892);
or U4652 (N_4652,N_1551,N_1772);
and U4653 (N_4653,N_116,N_979);
or U4654 (N_4654,N_2246,N_758);
and U4655 (N_4655,N_1619,N_539);
and U4656 (N_4656,N_1434,N_1316);
and U4657 (N_4657,N_1190,N_461);
nand U4658 (N_4658,N_1520,N_1323);
and U4659 (N_4659,N_79,N_1554);
or U4660 (N_4660,N_1787,N_2183);
nand U4661 (N_4661,N_1464,N_2092);
and U4662 (N_4662,N_2084,N_2368);
or U4663 (N_4663,N_286,N_2269);
xnor U4664 (N_4664,N_1966,N_837);
nand U4665 (N_4665,N_655,N_1808);
nand U4666 (N_4666,N_758,N_2166);
xnor U4667 (N_4667,N_1742,N_157);
or U4668 (N_4668,N_1891,N_1898);
nand U4669 (N_4669,N_1164,N_49);
or U4670 (N_4670,N_584,N_226);
xor U4671 (N_4671,N_672,N_2376);
nor U4672 (N_4672,N_1110,N_1428);
xnor U4673 (N_4673,N_217,N_460);
or U4674 (N_4674,N_1797,N_2458);
nand U4675 (N_4675,N_1488,N_2283);
nor U4676 (N_4676,N_1058,N_1253);
and U4677 (N_4677,N_1822,N_990);
nor U4678 (N_4678,N_2037,N_1396);
and U4679 (N_4679,N_1249,N_510);
or U4680 (N_4680,N_776,N_90);
nor U4681 (N_4681,N_833,N_1744);
nor U4682 (N_4682,N_2470,N_1438);
nor U4683 (N_4683,N_1080,N_241);
and U4684 (N_4684,N_1504,N_2085);
and U4685 (N_4685,N_1553,N_2273);
nor U4686 (N_4686,N_1662,N_1001);
and U4687 (N_4687,N_1045,N_1522);
nor U4688 (N_4688,N_2448,N_600);
nor U4689 (N_4689,N_1831,N_1026);
and U4690 (N_4690,N_457,N_1988);
or U4691 (N_4691,N_681,N_1437);
nand U4692 (N_4692,N_1208,N_2374);
nor U4693 (N_4693,N_2000,N_2105);
xor U4694 (N_4694,N_174,N_1220);
and U4695 (N_4695,N_626,N_2499);
and U4696 (N_4696,N_1213,N_370);
or U4697 (N_4697,N_873,N_2020);
nand U4698 (N_4698,N_221,N_76);
nor U4699 (N_4699,N_2416,N_645);
and U4700 (N_4700,N_594,N_540);
and U4701 (N_4701,N_1590,N_64);
and U4702 (N_4702,N_1756,N_404);
nor U4703 (N_4703,N_1019,N_1260);
or U4704 (N_4704,N_1282,N_1027);
nand U4705 (N_4705,N_1575,N_2175);
nand U4706 (N_4706,N_1311,N_652);
nor U4707 (N_4707,N_99,N_846);
nor U4708 (N_4708,N_286,N_1618);
nor U4709 (N_4709,N_242,N_1187);
nor U4710 (N_4710,N_2033,N_1935);
xor U4711 (N_4711,N_2142,N_1872);
and U4712 (N_4712,N_1376,N_1363);
or U4713 (N_4713,N_1313,N_987);
and U4714 (N_4714,N_1147,N_1099);
and U4715 (N_4715,N_1294,N_1727);
or U4716 (N_4716,N_1073,N_2369);
nor U4717 (N_4717,N_167,N_2226);
nor U4718 (N_4718,N_1962,N_1021);
xor U4719 (N_4719,N_842,N_296);
nor U4720 (N_4720,N_482,N_525);
nand U4721 (N_4721,N_1720,N_124);
nor U4722 (N_4722,N_1445,N_695);
nand U4723 (N_4723,N_1936,N_2393);
and U4724 (N_4724,N_2415,N_2139);
nor U4725 (N_4725,N_502,N_2309);
nor U4726 (N_4726,N_990,N_551);
nor U4727 (N_4727,N_1899,N_759);
nor U4728 (N_4728,N_1191,N_2267);
and U4729 (N_4729,N_1509,N_332);
nor U4730 (N_4730,N_1053,N_2297);
and U4731 (N_4731,N_1091,N_94);
and U4732 (N_4732,N_151,N_1762);
and U4733 (N_4733,N_620,N_1662);
and U4734 (N_4734,N_2041,N_1651);
and U4735 (N_4735,N_67,N_666);
nor U4736 (N_4736,N_1291,N_2381);
or U4737 (N_4737,N_2000,N_974);
or U4738 (N_4738,N_1484,N_2444);
or U4739 (N_4739,N_990,N_1372);
and U4740 (N_4740,N_1475,N_2376);
or U4741 (N_4741,N_38,N_1979);
nand U4742 (N_4742,N_2239,N_1771);
and U4743 (N_4743,N_1621,N_92);
nor U4744 (N_4744,N_860,N_103);
or U4745 (N_4745,N_293,N_664);
nand U4746 (N_4746,N_523,N_218);
xnor U4747 (N_4747,N_2467,N_1143);
nor U4748 (N_4748,N_547,N_1117);
nor U4749 (N_4749,N_2257,N_1484);
and U4750 (N_4750,N_2148,N_707);
nand U4751 (N_4751,N_2437,N_1598);
nand U4752 (N_4752,N_707,N_1980);
xor U4753 (N_4753,N_495,N_426);
nor U4754 (N_4754,N_129,N_1948);
and U4755 (N_4755,N_2458,N_143);
nor U4756 (N_4756,N_1892,N_980);
nand U4757 (N_4757,N_1037,N_1309);
and U4758 (N_4758,N_510,N_1743);
and U4759 (N_4759,N_2196,N_2041);
nor U4760 (N_4760,N_291,N_1963);
nor U4761 (N_4761,N_1337,N_32);
nor U4762 (N_4762,N_2363,N_1652);
and U4763 (N_4763,N_394,N_572);
and U4764 (N_4764,N_1141,N_1158);
and U4765 (N_4765,N_1851,N_77);
or U4766 (N_4766,N_213,N_1604);
nor U4767 (N_4767,N_615,N_881);
or U4768 (N_4768,N_2312,N_1679);
and U4769 (N_4769,N_2056,N_1044);
xor U4770 (N_4770,N_1195,N_387);
nor U4771 (N_4771,N_336,N_1895);
nor U4772 (N_4772,N_1943,N_803);
nor U4773 (N_4773,N_801,N_568);
or U4774 (N_4774,N_2005,N_18);
or U4775 (N_4775,N_362,N_2458);
xor U4776 (N_4776,N_1066,N_725);
and U4777 (N_4777,N_626,N_2024);
or U4778 (N_4778,N_2269,N_1165);
or U4779 (N_4779,N_287,N_452);
nor U4780 (N_4780,N_1660,N_1057);
nand U4781 (N_4781,N_586,N_285);
nor U4782 (N_4782,N_1334,N_1580);
xnor U4783 (N_4783,N_541,N_33);
or U4784 (N_4784,N_1987,N_248);
and U4785 (N_4785,N_1246,N_304);
nand U4786 (N_4786,N_1408,N_1622);
and U4787 (N_4787,N_1100,N_324);
nor U4788 (N_4788,N_1416,N_2028);
nor U4789 (N_4789,N_1432,N_1180);
nor U4790 (N_4790,N_124,N_2363);
nand U4791 (N_4791,N_2167,N_682);
nor U4792 (N_4792,N_827,N_2384);
and U4793 (N_4793,N_2463,N_298);
nand U4794 (N_4794,N_599,N_1337);
nand U4795 (N_4795,N_1153,N_1752);
nor U4796 (N_4796,N_439,N_1111);
nand U4797 (N_4797,N_1721,N_271);
and U4798 (N_4798,N_1844,N_1966);
nand U4799 (N_4799,N_997,N_344);
or U4800 (N_4800,N_614,N_1213);
or U4801 (N_4801,N_2177,N_444);
and U4802 (N_4802,N_105,N_1696);
or U4803 (N_4803,N_51,N_1241);
nand U4804 (N_4804,N_1597,N_281);
nor U4805 (N_4805,N_1278,N_1433);
xnor U4806 (N_4806,N_1975,N_1243);
and U4807 (N_4807,N_281,N_1691);
xor U4808 (N_4808,N_349,N_722);
nand U4809 (N_4809,N_753,N_2316);
and U4810 (N_4810,N_1191,N_2022);
nand U4811 (N_4811,N_47,N_812);
nor U4812 (N_4812,N_1364,N_1161);
and U4813 (N_4813,N_2006,N_1297);
and U4814 (N_4814,N_1778,N_815);
and U4815 (N_4815,N_443,N_2167);
or U4816 (N_4816,N_850,N_2261);
and U4817 (N_4817,N_1331,N_1853);
and U4818 (N_4818,N_1157,N_92);
xnor U4819 (N_4819,N_559,N_1311);
nor U4820 (N_4820,N_2340,N_608);
or U4821 (N_4821,N_1028,N_297);
nor U4822 (N_4822,N_650,N_2279);
and U4823 (N_4823,N_2274,N_689);
nor U4824 (N_4824,N_652,N_1141);
nand U4825 (N_4825,N_1161,N_100);
nand U4826 (N_4826,N_1477,N_1793);
nor U4827 (N_4827,N_834,N_2058);
or U4828 (N_4828,N_817,N_163);
nor U4829 (N_4829,N_160,N_1858);
nor U4830 (N_4830,N_1004,N_2432);
and U4831 (N_4831,N_2051,N_924);
or U4832 (N_4832,N_516,N_2318);
xor U4833 (N_4833,N_1191,N_70);
or U4834 (N_4834,N_341,N_2478);
nor U4835 (N_4835,N_930,N_250);
nand U4836 (N_4836,N_715,N_2348);
nand U4837 (N_4837,N_1391,N_2169);
or U4838 (N_4838,N_538,N_117);
or U4839 (N_4839,N_1033,N_214);
xnor U4840 (N_4840,N_1925,N_132);
nand U4841 (N_4841,N_1603,N_1599);
or U4842 (N_4842,N_309,N_2085);
and U4843 (N_4843,N_56,N_1800);
nand U4844 (N_4844,N_120,N_671);
nor U4845 (N_4845,N_1630,N_499);
nand U4846 (N_4846,N_2315,N_1723);
or U4847 (N_4847,N_607,N_1774);
nor U4848 (N_4848,N_848,N_939);
and U4849 (N_4849,N_2499,N_652);
nand U4850 (N_4850,N_642,N_941);
nand U4851 (N_4851,N_2357,N_220);
nor U4852 (N_4852,N_1014,N_2373);
nor U4853 (N_4853,N_1557,N_1713);
nor U4854 (N_4854,N_299,N_1015);
nand U4855 (N_4855,N_252,N_40);
nand U4856 (N_4856,N_2450,N_2196);
or U4857 (N_4857,N_938,N_1991);
nand U4858 (N_4858,N_1550,N_1134);
nor U4859 (N_4859,N_820,N_1845);
nand U4860 (N_4860,N_1312,N_1796);
or U4861 (N_4861,N_462,N_1451);
or U4862 (N_4862,N_81,N_1703);
xor U4863 (N_4863,N_1160,N_2228);
nand U4864 (N_4864,N_518,N_279);
or U4865 (N_4865,N_1648,N_293);
nor U4866 (N_4866,N_741,N_2147);
or U4867 (N_4867,N_927,N_193);
and U4868 (N_4868,N_1427,N_743);
or U4869 (N_4869,N_2257,N_541);
or U4870 (N_4870,N_1049,N_415);
or U4871 (N_4871,N_2425,N_2030);
nand U4872 (N_4872,N_77,N_2315);
nor U4873 (N_4873,N_905,N_780);
or U4874 (N_4874,N_2444,N_579);
nor U4875 (N_4875,N_1467,N_779);
nand U4876 (N_4876,N_384,N_2186);
xnor U4877 (N_4877,N_2073,N_2015);
and U4878 (N_4878,N_393,N_709);
nor U4879 (N_4879,N_997,N_257);
and U4880 (N_4880,N_69,N_788);
and U4881 (N_4881,N_1778,N_2334);
nand U4882 (N_4882,N_1431,N_1026);
nand U4883 (N_4883,N_981,N_1612);
and U4884 (N_4884,N_1876,N_1433);
nand U4885 (N_4885,N_2033,N_797);
nor U4886 (N_4886,N_1754,N_2202);
xnor U4887 (N_4887,N_901,N_633);
nor U4888 (N_4888,N_2295,N_1329);
and U4889 (N_4889,N_338,N_546);
nor U4890 (N_4890,N_2279,N_351);
nor U4891 (N_4891,N_823,N_1197);
nand U4892 (N_4892,N_2267,N_1749);
nor U4893 (N_4893,N_2140,N_1582);
nand U4894 (N_4894,N_1409,N_367);
nor U4895 (N_4895,N_864,N_1149);
and U4896 (N_4896,N_2333,N_164);
or U4897 (N_4897,N_1254,N_118);
nand U4898 (N_4898,N_2118,N_2224);
nand U4899 (N_4899,N_896,N_43);
and U4900 (N_4900,N_1460,N_354);
nand U4901 (N_4901,N_705,N_2270);
xor U4902 (N_4902,N_1119,N_4);
or U4903 (N_4903,N_1885,N_1751);
nor U4904 (N_4904,N_1473,N_500);
nor U4905 (N_4905,N_655,N_2162);
nand U4906 (N_4906,N_1682,N_158);
and U4907 (N_4907,N_2467,N_699);
nand U4908 (N_4908,N_585,N_2068);
nor U4909 (N_4909,N_1206,N_48);
nor U4910 (N_4910,N_1028,N_2086);
xor U4911 (N_4911,N_2119,N_2328);
and U4912 (N_4912,N_2394,N_826);
xnor U4913 (N_4913,N_1989,N_557);
or U4914 (N_4914,N_2035,N_2186);
nand U4915 (N_4915,N_80,N_1357);
and U4916 (N_4916,N_242,N_194);
nand U4917 (N_4917,N_2154,N_1134);
or U4918 (N_4918,N_300,N_239);
and U4919 (N_4919,N_1286,N_181);
and U4920 (N_4920,N_1602,N_901);
nand U4921 (N_4921,N_1187,N_884);
nand U4922 (N_4922,N_1290,N_2085);
nand U4923 (N_4923,N_1413,N_364);
and U4924 (N_4924,N_522,N_1460);
xnor U4925 (N_4925,N_975,N_1379);
xor U4926 (N_4926,N_1668,N_1914);
or U4927 (N_4927,N_199,N_2403);
and U4928 (N_4928,N_138,N_715);
and U4929 (N_4929,N_1133,N_324);
nand U4930 (N_4930,N_1680,N_780);
and U4931 (N_4931,N_1401,N_1885);
or U4932 (N_4932,N_773,N_955);
nor U4933 (N_4933,N_1979,N_1858);
or U4934 (N_4934,N_1897,N_2364);
or U4935 (N_4935,N_1616,N_401);
nand U4936 (N_4936,N_2355,N_2482);
and U4937 (N_4937,N_1656,N_175);
nand U4938 (N_4938,N_301,N_103);
nand U4939 (N_4939,N_1170,N_1029);
nand U4940 (N_4940,N_1417,N_1081);
xor U4941 (N_4941,N_262,N_1290);
nor U4942 (N_4942,N_2481,N_1621);
xor U4943 (N_4943,N_1500,N_1940);
nor U4944 (N_4944,N_28,N_610);
nor U4945 (N_4945,N_626,N_2228);
nand U4946 (N_4946,N_203,N_1066);
or U4947 (N_4947,N_1973,N_1692);
nand U4948 (N_4948,N_16,N_400);
nand U4949 (N_4949,N_1077,N_59);
xor U4950 (N_4950,N_517,N_1032);
or U4951 (N_4951,N_421,N_1013);
nor U4952 (N_4952,N_2115,N_730);
xor U4953 (N_4953,N_1647,N_914);
xor U4954 (N_4954,N_54,N_1169);
nand U4955 (N_4955,N_2424,N_1036);
nand U4956 (N_4956,N_2237,N_504);
nor U4957 (N_4957,N_632,N_1360);
nand U4958 (N_4958,N_1682,N_115);
nand U4959 (N_4959,N_2258,N_563);
nor U4960 (N_4960,N_686,N_584);
nand U4961 (N_4961,N_1575,N_966);
and U4962 (N_4962,N_1498,N_1582);
nand U4963 (N_4963,N_717,N_2392);
and U4964 (N_4964,N_140,N_385);
and U4965 (N_4965,N_2281,N_730);
and U4966 (N_4966,N_1149,N_1890);
nor U4967 (N_4967,N_1135,N_2189);
nand U4968 (N_4968,N_1112,N_1333);
nor U4969 (N_4969,N_550,N_24);
xnor U4970 (N_4970,N_1153,N_1422);
or U4971 (N_4971,N_1993,N_37);
or U4972 (N_4972,N_487,N_1655);
nor U4973 (N_4973,N_1458,N_927);
xor U4974 (N_4974,N_2006,N_2005);
and U4975 (N_4975,N_2046,N_149);
or U4976 (N_4976,N_1387,N_1816);
and U4977 (N_4977,N_1455,N_148);
and U4978 (N_4978,N_2165,N_274);
nand U4979 (N_4979,N_121,N_1153);
or U4980 (N_4980,N_1508,N_215);
or U4981 (N_4981,N_1738,N_1627);
and U4982 (N_4982,N_682,N_749);
or U4983 (N_4983,N_1180,N_800);
xor U4984 (N_4984,N_1985,N_2396);
or U4985 (N_4985,N_89,N_60);
or U4986 (N_4986,N_1366,N_1836);
and U4987 (N_4987,N_1313,N_2269);
xnor U4988 (N_4988,N_2145,N_149);
nand U4989 (N_4989,N_520,N_359);
nor U4990 (N_4990,N_1863,N_2325);
and U4991 (N_4991,N_989,N_142);
xor U4992 (N_4992,N_80,N_1505);
or U4993 (N_4993,N_931,N_726);
or U4994 (N_4994,N_973,N_2119);
nand U4995 (N_4995,N_2257,N_1397);
nand U4996 (N_4996,N_116,N_2234);
and U4997 (N_4997,N_2232,N_1932);
or U4998 (N_4998,N_2091,N_83);
or U4999 (N_4999,N_2019,N_1783);
and UO_0 (O_0,N_4889,N_3901);
nor UO_1 (O_1,N_3393,N_3221);
nor UO_2 (O_2,N_3321,N_4563);
nand UO_3 (O_3,N_4219,N_2675);
and UO_4 (O_4,N_4894,N_3669);
nor UO_5 (O_5,N_3892,N_2938);
nand UO_6 (O_6,N_4963,N_4533);
or UO_7 (O_7,N_3605,N_3546);
and UO_8 (O_8,N_2505,N_3325);
and UO_9 (O_9,N_3530,N_3150);
or UO_10 (O_10,N_3702,N_3448);
nor UO_11 (O_11,N_3711,N_3346);
and UO_12 (O_12,N_4129,N_2891);
nor UO_13 (O_13,N_4372,N_4237);
or UO_14 (O_14,N_3257,N_4893);
nand UO_15 (O_15,N_3703,N_4742);
nor UO_16 (O_16,N_3939,N_4689);
nor UO_17 (O_17,N_3042,N_4439);
and UO_18 (O_18,N_2716,N_3262);
or UO_19 (O_19,N_2669,N_4674);
or UO_20 (O_20,N_4047,N_4247);
nor UO_21 (O_21,N_3662,N_4686);
or UO_22 (O_22,N_3633,N_4437);
nor UO_23 (O_23,N_3493,N_4862);
nor UO_24 (O_24,N_4763,N_4859);
nand UO_25 (O_25,N_4141,N_4462);
and UO_26 (O_26,N_4778,N_4155);
nand UO_27 (O_27,N_3640,N_4080);
nor UO_28 (O_28,N_4407,N_2911);
nand UO_29 (O_29,N_3426,N_4594);
or UO_30 (O_30,N_3488,N_4978);
and UO_31 (O_31,N_3549,N_3418);
and UO_32 (O_32,N_2915,N_2872);
nor UO_33 (O_33,N_2865,N_2862);
nor UO_34 (O_34,N_2981,N_3130);
xor UO_35 (O_35,N_2689,N_3718);
and UO_36 (O_36,N_4195,N_4341);
or UO_37 (O_37,N_2856,N_3720);
and UO_38 (O_38,N_4553,N_4428);
nor UO_39 (O_39,N_4849,N_2925);
nand UO_40 (O_40,N_4732,N_3364);
xor UO_41 (O_41,N_3726,N_2984);
xnor UO_42 (O_42,N_4157,N_4024);
nand UO_43 (O_43,N_2806,N_3974);
and UO_44 (O_44,N_4401,N_2558);
and UO_45 (O_45,N_3473,N_4250);
nor UO_46 (O_46,N_4440,N_2534);
nor UO_47 (O_47,N_4881,N_4322);
nand UO_48 (O_48,N_3193,N_2711);
nand UO_49 (O_49,N_2590,N_2724);
nand UO_50 (O_50,N_2584,N_4333);
nand UO_51 (O_51,N_3139,N_2539);
nand UO_52 (O_52,N_4063,N_4925);
xnor UO_53 (O_53,N_4227,N_3240);
or UO_54 (O_54,N_4004,N_2900);
nand UO_55 (O_55,N_3397,N_2947);
nand UO_56 (O_56,N_4025,N_2685);
nand UO_57 (O_57,N_3353,N_4556);
xnor UO_58 (O_58,N_3784,N_4860);
nand UO_59 (O_59,N_4617,N_3300);
or UO_60 (O_60,N_3615,N_3832);
and UO_61 (O_61,N_4233,N_2813);
and UO_62 (O_62,N_4018,N_4127);
and UO_63 (O_63,N_4998,N_4040);
or UO_64 (O_64,N_2751,N_2730);
nand UO_65 (O_65,N_2566,N_4676);
nor UO_66 (O_66,N_3158,N_4957);
nor UO_67 (O_67,N_2957,N_3661);
or UO_68 (O_68,N_3636,N_3996);
and UO_69 (O_69,N_3502,N_4658);
nor UO_70 (O_70,N_4918,N_3308);
nor UO_71 (O_71,N_2846,N_3445);
and UO_72 (O_72,N_3285,N_4644);
nor UO_73 (O_73,N_2823,N_3781);
and UO_74 (O_74,N_3376,N_3752);
nand UO_75 (O_75,N_3555,N_4485);
and UO_76 (O_76,N_4972,N_4745);
or UO_77 (O_77,N_4604,N_3101);
nor UO_78 (O_78,N_4131,N_3153);
nor UO_79 (O_79,N_3867,N_3414);
or UO_80 (O_80,N_4202,N_3663);
and UO_81 (O_81,N_4021,N_4379);
and UO_82 (O_82,N_3843,N_2552);
xor UO_83 (O_83,N_2598,N_2512);
nand UO_84 (O_84,N_3891,N_2962);
and UO_85 (O_85,N_3174,N_3877);
nor UO_86 (O_86,N_3014,N_4959);
nand UO_87 (O_87,N_3046,N_4558);
xnor UO_88 (O_88,N_3675,N_4320);
nand UO_89 (O_89,N_3865,N_2754);
or UO_90 (O_90,N_4163,N_2781);
nand UO_91 (O_91,N_3383,N_4703);
and UO_92 (O_92,N_2824,N_3269);
xnor UO_93 (O_93,N_3307,N_2560);
or UO_94 (O_94,N_4182,N_4135);
and UO_95 (O_95,N_3911,N_2670);
nor UO_96 (O_96,N_2994,N_4082);
or UO_97 (O_97,N_4713,N_3099);
nand UO_98 (O_98,N_4145,N_3978);
xor UO_99 (O_99,N_4376,N_4993);
or UO_100 (O_100,N_2744,N_3075);
or UO_101 (O_101,N_3273,N_3433);
xnor UO_102 (O_102,N_2561,N_4788);
nand UO_103 (O_103,N_3694,N_2686);
nand UO_104 (O_104,N_4632,N_4944);
nand UO_105 (O_105,N_2701,N_4152);
or UO_106 (O_106,N_3647,N_3519);
nor UO_107 (O_107,N_2960,N_2913);
nand UO_108 (O_108,N_4242,N_4693);
and UO_109 (O_109,N_4646,N_3229);
or UO_110 (O_110,N_4431,N_2531);
nand UO_111 (O_111,N_2919,N_4349);
or UO_112 (O_112,N_4651,N_4191);
xor UO_113 (O_113,N_3791,N_3618);
xor UO_114 (O_114,N_3952,N_4920);
nor UO_115 (O_115,N_3734,N_3776);
nor UO_116 (O_116,N_3856,N_3186);
or UO_117 (O_117,N_2710,N_3635);
nand UO_118 (O_118,N_3271,N_3244);
nand UO_119 (O_119,N_4273,N_3085);
and UO_120 (O_120,N_4159,N_2948);
nor UO_121 (O_121,N_3217,N_2559);
xor UO_122 (O_122,N_3505,N_2732);
or UO_123 (O_123,N_4694,N_4261);
and UO_124 (O_124,N_3523,N_2811);
or UO_125 (O_125,N_3077,N_3517);
or UO_126 (O_126,N_2547,N_3591);
nand UO_127 (O_127,N_2639,N_2506);
xor UO_128 (O_128,N_2897,N_2654);
xnor UO_129 (O_129,N_3476,N_4169);
and UO_130 (O_130,N_4297,N_4013);
nor UO_131 (O_131,N_3379,N_2804);
nand UO_132 (O_132,N_4373,N_2757);
nand UO_133 (O_133,N_3278,N_4675);
or UO_134 (O_134,N_4698,N_3685);
or UO_135 (O_135,N_4608,N_4568);
nor UO_136 (O_136,N_3929,N_4422);
xnor UO_137 (O_137,N_4805,N_4123);
or UO_138 (O_138,N_3252,N_2963);
nand UO_139 (O_139,N_2624,N_3303);
nor UO_140 (O_140,N_3746,N_4058);
nand UO_141 (O_141,N_2604,N_3668);
nor UO_142 (O_142,N_3255,N_4965);
nand UO_143 (O_143,N_4335,N_3622);
xor UO_144 (O_144,N_4610,N_4907);
nand UO_145 (O_145,N_2568,N_3169);
or UO_146 (O_146,N_2904,N_2507);
nor UO_147 (O_147,N_3880,N_3888);
and UO_148 (O_148,N_4387,N_4807);
nand UO_149 (O_149,N_3848,N_4678);
or UO_150 (O_150,N_4890,N_3806);
or UO_151 (O_151,N_3080,N_4601);
and UO_152 (O_152,N_3587,N_3741);
nand UO_153 (O_153,N_2935,N_3770);
nand UO_154 (O_154,N_3037,N_3029);
and UO_155 (O_155,N_2735,N_3601);
nor UO_156 (O_156,N_4648,N_3567);
and UO_157 (O_157,N_3611,N_4098);
nor UO_158 (O_158,N_3179,N_3422);
nand UO_159 (O_159,N_4170,N_4491);
or UO_160 (O_160,N_4101,N_3511);
xnor UO_161 (O_161,N_4724,N_4270);
or UO_162 (O_162,N_3864,N_3884);
and UO_163 (O_163,N_2799,N_3462);
xor UO_164 (O_164,N_4011,N_2971);
and UO_165 (O_165,N_4043,N_3919);
nor UO_166 (O_166,N_4915,N_2623);
or UO_167 (O_167,N_3574,N_2642);
or UO_168 (O_168,N_4314,N_4464);
nor UO_169 (O_169,N_3040,N_2700);
nor UO_170 (O_170,N_4748,N_3686);
or UO_171 (O_171,N_3831,N_4355);
nand UO_172 (O_172,N_3171,N_2793);
or UO_173 (O_173,N_2819,N_2660);
nor UO_174 (O_174,N_4128,N_4706);
and UO_175 (O_175,N_4891,N_4292);
or UO_176 (O_176,N_3276,N_4587);
or UO_177 (O_177,N_4543,N_4909);
nor UO_178 (O_178,N_3156,N_3041);
and UO_179 (O_179,N_4573,N_4806);
nor UO_180 (O_180,N_4663,N_4629);
nor UO_181 (O_181,N_3090,N_3145);
nand UO_182 (O_182,N_3081,N_4985);
nand UO_183 (O_183,N_4512,N_4991);
and UO_184 (O_184,N_4666,N_3194);
and UO_185 (O_185,N_3354,N_3190);
nand UO_186 (O_186,N_2662,N_4221);
nand UO_187 (O_187,N_4330,N_4076);
or UO_188 (O_188,N_3132,N_2929);
and UO_189 (O_189,N_2576,N_2708);
or UO_190 (O_190,N_3007,N_4690);
xnor UO_191 (O_191,N_3026,N_4623);
xnor UO_192 (O_192,N_4150,N_3123);
and UO_193 (O_193,N_2516,N_2525);
nand UO_194 (O_194,N_2653,N_2922);
and UO_195 (O_195,N_4096,N_3411);
xor UO_196 (O_196,N_3748,N_2659);
nand UO_197 (O_197,N_3800,N_4750);
nor UO_198 (O_198,N_3167,N_3682);
or UO_199 (O_199,N_4790,N_2875);
nand UO_200 (O_200,N_2821,N_4901);
nand UO_201 (O_201,N_3482,N_3655);
and UO_202 (O_202,N_2645,N_4786);
nand UO_203 (O_203,N_2609,N_2830);
and UO_204 (O_204,N_4739,N_3958);
nand UO_205 (O_205,N_4821,N_2916);
nand UO_206 (O_206,N_2614,N_2779);
nor UO_207 (O_207,N_3700,N_4412);
nand UO_208 (O_208,N_2556,N_3282);
nor UO_209 (O_209,N_3071,N_3362);
nand UO_210 (O_210,N_3286,N_3573);
nor UO_211 (O_211,N_2648,N_4995);
nor UO_212 (O_212,N_3289,N_3842);
and UO_213 (O_213,N_3117,N_2895);
xor UO_214 (O_214,N_4118,N_2827);
or UO_215 (O_215,N_3201,N_3897);
or UO_216 (O_216,N_4019,N_3225);
and UO_217 (O_217,N_2863,N_4682);
nand UO_218 (O_218,N_3950,N_4243);
and UO_219 (O_219,N_4103,N_4091);
nor UO_220 (O_220,N_3425,N_3947);
nor UO_221 (O_221,N_2762,N_4133);
and UO_222 (O_222,N_3423,N_2546);
and UO_223 (O_223,N_2973,N_4356);
nand UO_224 (O_224,N_4621,N_4125);
nor UO_225 (O_225,N_3003,N_3997);
nor UO_226 (O_226,N_3559,N_4386);
and UO_227 (O_227,N_4905,N_4911);
xor UO_228 (O_228,N_3665,N_4229);
xnor UO_229 (O_229,N_3359,N_4490);
nand UO_230 (O_230,N_4184,N_2557);
or UO_231 (O_231,N_4442,N_2652);
nor UO_232 (O_232,N_3973,N_2553);
xnor UO_233 (O_233,N_3480,N_4837);
nor UO_234 (O_234,N_4461,N_4359);
nand UO_235 (O_235,N_4639,N_3520);
nor UO_236 (O_236,N_4855,N_2840);
nand UO_237 (O_237,N_4649,N_3582);
and UO_238 (O_238,N_4824,N_4005);
nor UO_239 (O_239,N_4463,N_2765);
nand UO_240 (O_240,N_4307,N_4677);
or UO_241 (O_241,N_3641,N_3056);
nor UO_242 (O_242,N_4968,N_3428);
nand UO_243 (O_243,N_4916,N_2647);
or UO_244 (O_244,N_3142,N_3609);
nor UO_245 (O_245,N_4754,N_3575);
nor UO_246 (O_246,N_4215,N_3027);
and UO_247 (O_247,N_3310,N_2788);
or UO_248 (O_248,N_3219,N_4506);
or UO_249 (O_249,N_3373,N_4519);
nand UO_250 (O_250,N_3730,N_3485);
or UO_251 (O_251,N_3808,N_3597);
and UO_252 (O_252,N_4873,N_4257);
and UO_253 (O_253,N_3930,N_3385);
nand UO_254 (O_254,N_2745,N_3438);
and UO_255 (O_255,N_4939,N_4983);
nor UO_256 (O_256,N_4725,N_3413);
nor UO_257 (O_257,N_2691,N_3468);
nand UO_258 (O_258,N_3094,N_2555);
and UO_259 (O_259,N_3501,N_3088);
and UO_260 (O_260,N_3756,N_4210);
nand UO_261 (O_261,N_4033,N_3568);
or UO_262 (O_262,N_4926,N_3136);
nand UO_263 (O_263,N_2894,N_4728);
and UO_264 (O_264,N_4458,N_4628);
or UO_265 (O_265,N_4220,N_2709);
and UO_266 (O_266,N_3785,N_4028);
and UO_267 (O_267,N_4650,N_4833);
nor UO_268 (O_268,N_3002,N_2883);
or UO_269 (O_269,N_2734,N_3104);
nor UO_270 (O_270,N_4271,N_2888);
and UO_271 (O_271,N_3280,N_4929);
nor UO_272 (O_272,N_4717,N_3751);
or UO_273 (O_273,N_4979,N_4704);
or UO_274 (O_274,N_4245,N_2635);
and UO_275 (O_275,N_4472,N_2787);
and UO_276 (O_276,N_4761,N_2597);
nand UO_277 (O_277,N_4715,N_4953);
nor UO_278 (O_278,N_3098,N_4664);
and UO_279 (O_279,N_4367,N_2780);
xnor UO_280 (O_280,N_3926,N_4535);
and UO_281 (O_281,N_2727,N_2812);
and UO_282 (O_282,N_4090,N_3616);
or UO_283 (O_283,N_2847,N_4352);
nor UO_284 (O_284,N_3933,N_4945);
nand UO_285 (O_285,N_3021,N_3034);
or UO_286 (O_286,N_4630,N_3713);
nor UO_287 (O_287,N_3747,N_3788);
nor UO_288 (O_288,N_2853,N_3982);
nand UO_289 (O_289,N_3889,N_3382);
nor UO_290 (O_290,N_4117,N_3122);
xor UO_291 (O_291,N_4039,N_3813);
and UO_292 (O_292,N_4696,N_4012);
nor UO_293 (O_293,N_4999,N_3890);
nand UO_294 (O_294,N_3613,N_4814);
or UO_295 (O_295,N_4546,N_3696);
and UO_296 (O_296,N_4228,N_4008);
nand UO_297 (O_297,N_3358,N_4771);
xor UO_298 (O_298,N_3768,N_2968);
nand UO_299 (O_299,N_3994,N_3722);
and UO_300 (O_300,N_3484,N_3909);
and UO_301 (O_301,N_3012,N_2785);
and UO_302 (O_302,N_3922,N_3671);
nand UO_303 (O_303,N_2725,N_3779);
nand UO_304 (O_304,N_4108,N_2743);
xnor UO_305 (O_305,N_3610,N_3338);
and UO_306 (O_306,N_3670,N_3323);
nand UO_307 (O_307,N_4218,N_4501);
and UO_308 (O_308,N_2718,N_4138);
and UO_309 (O_309,N_2796,N_4389);
and UO_310 (O_310,N_4812,N_4508);
nor UO_311 (O_311,N_3465,N_3216);
nand UO_312 (O_312,N_4026,N_4374);
nand UO_313 (O_313,N_3175,N_4204);
nor UO_314 (O_314,N_3138,N_3115);
xor UO_315 (O_315,N_4903,N_4347);
and UO_316 (O_316,N_3566,N_4528);
and UO_317 (O_317,N_3691,N_3653);
nor UO_318 (O_318,N_2589,N_4902);
xor UO_319 (O_319,N_3263,N_3695);
nand UO_320 (O_320,N_3769,N_3805);
nor UO_321 (O_321,N_3883,N_2671);
or UO_322 (O_322,N_2607,N_2949);
and UO_323 (O_323,N_3232,N_2773);
nand UO_324 (O_324,N_4569,N_4255);
or UO_325 (O_325,N_4549,N_4942);
nand UO_326 (O_326,N_3869,N_3849);
nor UO_327 (O_327,N_3729,N_2975);
nand UO_328 (O_328,N_2707,N_4884);
or UO_329 (O_329,N_3833,N_3860);
or UO_330 (O_330,N_4764,N_3823);
and UO_331 (O_331,N_2921,N_2985);
or UO_332 (O_332,N_3052,N_4712);
and UO_333 (O_333,N_3623,N_4060);
and UO_334 (O_334,N_3450,N_2839);
or UO_335 (O_335,N_4055,N_4647);
and UO_336 (O_336,N_2632,N_4162);
nand UO_337 (O_337,N_2837,N_3267);
or UO_338 (O_338,N_3799,N_3008);
nor UO_339 (O_339,N_3822,N_4829);
xnor UO_340 (O_340,N_4923,N_2829);
or UO_341 (O_341,N_3689,N_3536);
and UO_342 (O_342,N_2931,N_4510);
or UO_343 (O_343,N_4223,N_4857);
and UO_344 (O_344,N_3927,N_4364);
nand UO_345 (O_345,N_4430,N_3336);
and UO_346 (O_346,N_4611,N_4029);
or UO_347 (O_347,N_3375,N_3006);
nand UO_348 (O_348,N_4588,N_4323);
or UO_349 (O_349,N_4190,N_4643);
or UO_350 (O_350,N_4800,N_4310);
and UO_351 (O_351,N_4231,N_3246);
nand UO_352 (O_352,N_3427,N_3116);
nor UO_353 (O_353,N_4074,N_4226);
nand UO_354 (O_354,N_4536,N_4969);
nor UO_355 (O_355,N_4934,N_4484);
and UO_356 (O_356,N_3506,N_4346);
nand UO_357 (O_357,N_3558,N_3494);
nand UO_358 (O_358,N_4544,N_4151);
nand UO_359 (O_359,N_4752,N_4615);
nor UO_360 (O_360,N_3957,N_4395);
nand UO_361 (O_361,N_3816,N_4415);
or UO_362 (O_362,N_4357,N_3590);
nor UO_363 (O_363,N_3538,N_4010);
nand UO_364 (O_364,N_3872,N_3062);
nand UO_365 (O_365,N_2617,N_3178);
and UO_366 (O_366,N_4887,N_4813);
or UO_367 (O_367,N_3233,N_3055);
nand UO_368 (O_368,N_3648,N_2777);
or UO_369 (O_369,N_2563,N_4147);
xor UO_370 (O_370,N_4877,N_3614);
nand UO_371 (O_371,N_4105,N_4216);
nand UO_372 (O_372,N_3421,N_2684);
and UO_373 (O_373,N_3925,N_3224);
and UO_374 (O_374,N_4614,N_3654);
nor UO_375 (O_375,N_3699,N_4470);
nand UO_376 (O_376,N_3908,N_3328);
nand UO_377 (O_377,N_2509,N_4432);
or UO_378 (O_378,N_4071,N_4200);
nor UO_379 (O_379,N_4345,N_3078);
nor UO_380 (O_380,N_4636,N_3773);
or UO_381 (O_381,N_3985,N_4433);
nor UO_382 (O_382,N_4403,N_2936);
xnor UO_383 (O_383,N_2574,N_3405);
nand UO_384 (O_384,N_4207,N_2995);
nor UO_385 (O_385,N_2712,N_3643);
nor UO_386 (O_386,N_3552,N_3940);
or UO_387 (O_387,N_3329,N_4197);
or UO_388 (O_388,N_2966,N_4937);
or UO_389 (O_389,N_4460,N_3410);
nor UO_390 (O_390,N_4478,N_3586);
nand UO_391 (O_391,N_2884,N_4548);
and UO_392 (O_392,N_4079,N_3395);
nor UO_393 (O_393,N_4507,N_4921);
or UO_394 (O_394,N_2564,N_4511);
and UO_395 (O_395,N_4052,N_2603);
nand UO_396 (O_396,N_3250,N_4048);
and UO_397 (O_397,N_3107,N_4593);
or UO_398 (O_398,N_4592,N_4538);
nor UO_399 (O_399,N_2668,N_3830);
nor UO_400 (O_400,N_3378,N_4022);
nand UO_401 (O_401,N_4795,N_3228);
nand UO_402 (O_402,N_4034,N_2852);
nand UO_403 (O_403,N_4050,N_3499);
xnor UO_404 (O_404,N_3858,N_2914);
nor UO_405 (O_405,N_3327,N_4001);
or UO_406 (O_406,N_3431,N_3065);
nor UO_407 (O_407,N_2620,N_4360);
nand UO_408 (O_408,N_2881,N_3048);
and UO_409 (O_409,N_4279,N_3133);
or UO_410 (O_410,N_2808,N_4225);
and UO_411 (O_411,N_4411,N_4827);
nand UO_412 (O_412,N_4093,N_3659);
or UO_413 (O_413,N_4932,N_4196);
nor UO_414 (O_414,N_3563,N_4987);
nand UO_415 (O_415,N_4494,N_4171);
or UO_416 (O_416,N_3828,N_4688);
and UO_417 (O_417,N_3164,N_4154);
or UO_418 (O_418,N_3798,N_3507);
or UO_419 (O_419,N_4875,N_4952);
nand UO_420 (O_420,N_2991,N_4851);
and UO_421 (O_421,N_4518,N_4695);
nor UO_422 (O_422,N_4880,N_4595);
and UO_423 (O_423,N_2513,N_4612);
nor UO_424 (O_424,N_3264,N_2521);
nand UO_425 (O_425,N_3258,N_4622);
and UO_426 (O_426,N_3988,N_4044);
nor UO_427 (O_427,N_4590,N_4733);
and UO_428 (O_428,N_4282,N_3245);
nand UO_429 (O_429,N_4404,N_3172);
nand UO_430 (O_430,N_3656,N_3357);
nand UO_431 (O_431,N_2771,N_3592);
nor UO_432 (O_432,N_3604,N_3914);
xor UO_433 (O_433,N_3322,N_3020);
or UO_434 (O_434,N_2517,N_3429);
and UO_435 (O_435,N_2946,N_2690);
nand UO_436 (O_436,N_4616,N_2600);
or UO_437 (O_437,N_3016,N_4051);
nand UO_438 (O_438,N_4700,N_3451);
or UO_439 (O_439,N_4469,N_2738);
or UO_440 (O_440,N_4808,N_3624);
nand UO_441 (O_441,N_3059,N_3820);
or UO_442 (O_442,N_4872,N_3495);
nand UO_443 (O_443,N_2523,N_2767);
and UO_444 (O_444,N_4235,N_2851);
nand UO_445 (O_445,N_4815,N_4789);
and UO_446 (O_446,N_4818,N_4868);
and UO_447 (O_447,N_4803,N_4002);
xnor UO_448 (O_448,N_4318,N_4289);
and UO_449 (O_449,N_3369,N_3345);
or UO_450 (O_450,N_3963,N_2575);
and UO_451 (O_451,N_4239,N_3355);
nand UO_452 (O_452,N_3334,N_3570);
xnor UO_453 (O_453,N_4496,N_3199);
and UO_454 (O_454,N_3771,N_4417);
or UO_455 (O_455,N_4094,N_3299);
xor UO_456 (O_456,N_4278,N_2703);
and UO_457 (O_457,N_4637,N_3089);
xnor UO_458 (O_458,N_4955,N_4720);
xnor UO_459 (O_459,N_3564,N_2694);
or UO_460 (O_460,N_3038,N_4084);
and UO_461 (O_461,N_4502,N_3991);
xor UO_462 (O_462,N_4941,N_3625);
or UO_463 (O_463,N_2550,N_3110);
and UO_464 (O_464,N_3868,N_2901);
and UO_465 (O_465,N_4111,N_4804);
nand UO_466 (O_466,N_3907,N_4656);
or UO_467 (O_467,N_4075,N_3441);
nor UO_468 (O_468,N_3166,N_3143);
nand UO_469 (O_469,N_4455,N_2972);
nand UO_470 (O_470,N_3817,N_4311);
xor UO_471 (O_471,N_2783,N_4280);
or UO_472 (O_472,N_2896,N_2818);
xnor UO_473 (O_473,N_2562,N_3954);
xnor UO_474 (O_474,N_3335,N_3057);
nand UO_475 (O_475,N_4366,N_3508);
or UO_476 (O_476,N_3560,N_3434);
and UO_477 (O_477,N_4874,N_2842);
nor UO_478 (O_478,N_4418,N_4468);
and UO_479 (O_479,N_3518,N_2540);
and UO_480 (O_480,N_4185,N_4962);
nor UO_481 (O_481,N_3019,N_4272);
nand UO_482 (O_482,N_4627,N_4557);
nor UO_483 (O_483,N_2702,N_3238);
nand UO_484 (O_484,N_4817,N_2582);
nor UO_485 (O_485,N_2979,N_2705);
and UO_486 (O_486,N_4448,N_4681);
and UO_487 (O_487,N_3073,N_2680);
or UO_488 (O_488,N_3235,N_4583);
nor UO_489 (O_489,N_2776,N_3898);
nor UO_490 (O_490,N_2892,N_4825);
and UO_491 (O_491,N_4095,N_4578);
nor UO_492 (O_492,N_4187,N_3758);
nand UO_493 (O_493,N_4259,N_3443);
xnor UO_494 (O_494,N_3902,N_3966);
nor UO_495 (O_495,N_4505,N_2510);
nor UO_496 (O_496,N_4236,N_3732);
nand UO_497 (O_497,N_4722,N_3176);
and UO_498 (O_498,N_4930,N_4876);
or UO_499 (O_499,N_2739,N_4577);
nor UO_500 (O_500,N_4246,N_4107);
and UO_501 (O_501,N_4038,N_4912);
and UO_502 (O_502,N_3572,N_4435);
nor UO_503 (O_503,N_4423,N_4365);
or UO_504 (O_504,N_4336,N_3363);
or UO_505 (O_505,N_4222,N_2588);
xnor UO_506 (O_506,N_4560,N_3440);
nor UO_507 (O_507,N_3727,N_4797);
nand UO_508 (O_508,N_3857,N_2970);
nand UO_509 (O_509,N_2591,N_2737);
xor UO_510 (O_510,N_4059,N_4416);
and UO_511 (O_511,N_2907,N_3096);
nor UO_512 (O_512,N_3672,N_2616);
or UO_513 (O_513,N_4148,N_3878);
nor UO_514 (O_514,N_4746,N_4238);
nor UO_515 (O_515,N_4267,N_3544);
nand UO_516 (O_516,N_4582,N_3128);
xor UO_517 (O_517,N_2527,N_3969);
nor UO_518 (O_518,N_4757,N_3188);
nor UO_519 (O_519,N_4447,N_3795);
nor UO_520 (O_520,N_3483,N_3854);
nor UO_521 (O_521,N_3399,N_4657);
or UO_522 (O_522,N_3881,N_4492);
or UO_523 (O_523,N_3010,N_3211);
nand UO_524 (O_524,N_4041,N_2822);
and UO_525 (O_525,N_4793,N_4654);
or UO_526 (O_526,N_4989,N_2859);
or UO_527 (O_527,N_2939,N_3737);
nand UO_528 (O_528,N_3131,N_4115);
xor UO_529 (O_529,N_2665,N_3102);
nand UO_530 (O_530,N_4756,N_4158);
or UO_531 (O_531,N_2601,N_4547);
or UO_532 (O_532,N_4679,N_4205);
nor UO_533 (O_533,N_4810,N_4343);
nor UO_534 (O_534,N_3742,N_4120);
nor UO_535 (O_535,N_3984,N_3755);
and UO_536 (O_536,N_3070,N_2683);
xor UO_537 (O_537,N_3305,N_4277);
and UO_538 (O_538,N_3948,N_3015);
nor UO_539 (O_539,N_4449,N_3230);
nand UO_540 (O_540,N_3960,N_3384);
and UO_541 (O_541,N_2959,N_3287);
nor UO_542 (O_542,N_4716,N_3844);
nand UO_543 (O_543,N_3667,N_3472);
or UO_544 (O_544,N_3017,N_4758);
nor UO_545 (O_545,N_2522,N_3709);
and UO_546 (O_546,N_2927,N_2944);
or UO_547 (O_547,N_3458,N_2651);
or UO_548 (O_548,N_4284,N_3237);
nor UO_549 (O_549,N_3904,N_3955);
or UO_550 (O_550,N_3923,N_4530);
and UO_551 (O_551,N_4863,N_4069);
or UO_552 (O_552,N_4371,N_3543);
and UO_553 (O_553,N_3548,N_4067);
nor UO_554 (O_554,N_4392,N_3840);
and UO_555 (O_555,N_3220,N_4275);
or UO_556 (O_556,N_2759,N_4329);
nand UO_557 (O_557,N_4014,N_4268);
xnor UO_558 (O_558,N_3887,N_3419);
or UO_559 (O_559,N_2950,N_3067);
nor UO_560 (O_560,N_4785,N_3753);
and UO_561 (O_561,N_3314,N_3717);
nor UO_562 (O_562,N_3896,N_2674);
or UO_563 (O_563,N_2768,N_3550);
or UO_564 (O_564,N_4400,N_4701);
xor UO_565 (O_565,N_3497,N_2833);
or UO_566 (O_566,N_2719,N_2693);
and UO_567 (O_567,N_4714,N_4620);
and UO_568 (O_568,N_2885,N_2636);
nor UO_569 (O_569,N_3850,N_3621);
and UO_570 (O_570,N_4232,N_3851);
nand UO_571 (O_571,N_4459,N_3704);
nor UO_572 (O_572,N_2814,N_2658);
nor UO_573 (O_573,N_3594,N_4721);
xor UO_574 (O_574,N_3053,N_2887);
nand UO_575 (O_575,N_4296,N_4609);
nand UO_576 (O_576,N_4377,N_3213);
xnor UO_577 (O_577,N_4475,N_3524);
or UO_578 (O_578,N_2764,N_3526);
or UO_579 (O_579,N_4525,N_4179);
nand UO_580 (O_580,N_3197,N_2990);
nand UO_581 (O_581,N_3396,N_2952);
nand UO_582 (O_582,N_4886,N_4444);
nand UO_583 (O_583,N_4668,N_3917);
nor UO_584 (O_584,N_3740,N_4865);
or UO_585 (O_585,N_4199,N_3212);
and UO_586 (O_586,N_4673,N_2876);
nand UO_587 (O_587,N_4122,N_4954);
and UO_588 (O_588,N_4509,N_4826);
or UO_589 (O_589,N_3478,N_3639);
nor UO_590 (O_590,N_4705,N_4178);
nand UO_591 (O_591,N_4426,N_4328);
nor UO_592 (O_592,N_2774,N_3204);
nand UO_593 (O_593,N_4498,N_4542);
nand UO_594 (O_594,N_4413,N_3324);
nor UO_595 (O_595,N_2594,N_4838);
nor UO_596 (O_596,N_3074,N_4769);
nor UO_597 (O_597,N_2596,N_4181);
nor UO_598 (O_598,N_3242,N_2926);
or UO_599 (O_599,N_3436,N_3146);
xor UO_600 (O_600,N_4112,N_4143);
nor UO_601 (O_601,N_3975,N_3388);
and UO_602 (O_602,N_3979,N_4904);
or UO_603 (O_603,N_2967,N_4741);
and UO_604 (O_604,N_3565,N_4943);
and UO_605 (O_605,N_2815,N_3477);
or UO_606 (O_606,N_2746,N_4309);
and UO_607 (O_607,N_4126,N_3964);
nor UO_608 (O_608,N_4189,N_4281);
nand UO_609 (O_609,N_4283,N_3206);
and UO_610 (O_610,N_2993,N_4503);
or UO_611 (O_611,N_2578,N_2772);
nor UO_612 (O_612,N_3972,N_4326);
or UO_613 (O_613,N_3666,N_3970);
and UO_614 (O_614,N_4856,N_3578);
nand UO_615 (O_615,N_3804,N_2845);
or UO_616 (O_616,N_4928,N_2637);
nand UO_617 (O_617,N_4217,N_4802);
and UO_618 (O_618,N_4065,N_3811);
nand UO_619 (O_619,N_4208,N_2508);
or UO_620 (O_620,N_4454,N_4619);
nor UO_621 (O_621,N_3693,N_4816);
nand UO_622 (O_622,N_4669,N_3871);
nand UO_623 (O_623,N_4290,N_2592);
or UO_624 (O_624,N_4531,N_4529);
xor UO_625 (O_625,N_3910,N_4753);
nor UO_626 (O_626,N_3380,N_4847);
or UO_627 (O_627,N_4089,N_3852);
or UO_628 (O_628,N_3024,N_3541);
nand UO_629 (O_629,N_2961,N_2866);
nand UO_630 (O_630,N_4244,N_4085);
xnor UO_631 (O_631,N_3853,N_3608);
and UO_632 (O_632,N_4994,N_4697);
and UO_633 (O_633,N_4212,N_3214);
nor UO_634 (O_634,N_4097,N_3990);
and UO_635 (O_635,N_4109,N_3159);
or UO_636 (O_636,N_3545,N_3439);
nor UO_637 (O_637,N_3231,N_4144);
or UO_638 (O_638,N_2810,N_2682);
or UO_639 (O_639,N_2630,N_4635);
and UO_640 (O_640,N_4765,N_3792);
nand UO_641 (O_641,N_2676,N_3452);
nor UO_642 (O_642,N_3976,N_2673);
nor UO_643 (O_643,N_3215,N_4308);
nor UO_644 (O_644,N_2677,N_2943);
nor UO_645 (O_645,N_3801,N_4369);
nand UO_646 (O_646,N_3292,N_2657);
or UO_647 (O_647,N_3777,N_4385);
nand UO_648 (O_648,N_3404,N_4950);
nand UO_649 (O_649,N_3521,N_4390);
and UO_650 (O_650,N_3372,N_4319);
xnor UO_651 (O_651,N_4613,N_4394);
nor UO_652 (O_652,N_4397,N_3481);
or UO_653 (O_653,N_2729,N_3129);
and UO_654 (O_654,N_4325,N_4175);
nor UO_655 (O_655,N_4834,N_4843);
and UO_656 (O_656,N_3637,N_3254);
or UO_657 (O_657,N_3905,N_4906);
and UO_658 (O_658,N_3588,N_2873);
and UO_659 (O_659,N_3706,N_2924);
and UO_660 (O_660,N_3602,N_2664);
and UO_661 (O_661,N_3941,N_4869);
nand UO_662 (O_662,N_4438,N_2502);
or UO_663 (O_663,N_4086,N_4031);
or UO_664 (O_664,N_4633,N_4316);
nor UO_665 (O_665,N_2749,N_4766);
or UO_666 (O_666,N_3148,N_3205);
or UO_667 (O_667,N_4564,N_3249);
or UO_668 (O_668,N_2969,N_3681);
nor UO_669 (O_669,N_3774,N_3810);
or UO_670 (O_670,N_4665,N_4457);
nor UO_671 (O_671,N_2820,N_4850);
xor UO_672 (O_672,N_3125,N_3084);
and UO_673 (O_673,N_3196,N_3093);
nor UO_674 (O_674,N_3351,N_4780);
and UO_675 (O_675,N_4956,N_4465);
nand UO_676 (O_676,N_4574,N_2752);
nor UO_677 (O_677,N_4361,N_3063);
xnor UO_678 (O_678,N_4393,N_4513);
xor UO_679 (O_679,N_4762,N_3934);
xnor UO_680 (O_680,N_2753,N_4719);
or UO_681 (O_681,N_3961,N_4249);
nand UO_682 (O_682,N_3942,N_4809);
nand UO_683 (O_683,N_4452,N_4738);
or UO_684 (O_684,N_3514,N_4760);
nor UO_685 (O_685,N_2519,N_2501);
and UO_686 (O_686,N_3617,N_3886);
nor UO_687 (O_687,N_4164,N_4344);
or UO_688 (O_688,N_2918,N_3736);
nor UO_689 (O_689,N_4211,N_4783);
nand UO_690 (O_690,N_3463,N_3525);
and UO_691 (O_691,N_4794,N_3218);
and UO_692 (O_692,N_4541,N_2836);
nor UO_693 (O_693,N_2878,N_3182);
and UO_694 (O_694,N_3453,N_3049);
nand UO_695 (O_695,N_4035,N_2698);
nand UO_696 (O_696,N_2720,N_3028);
or UO_697 (O_697,N_4726,N_4420);
nor UO_698 (O_698,N_3435,N_3302);
or UO_699 (O_699,N_4049,N_2537);
and UO_700 (O_700,N_4730,N_4552);
and UO_701 (O_701,N_3874,N_3715);
nand UO_702 (O_702,N_4897,N_4980);
xor UO_703 (O_703,N_3983,N_2855);
or UO_704 (O_704,N_4709,N_2890);
or UO_705 (O_705,N_2870,N_3556);
or UO_706 (O_706,N_3398,N_4399);
xor UO_707 (O_707,N_4521,N_4092);
nand UO_708 (O_708,N_3424,N_3119);
nand UO_709 (O_709,N_3248,N_3112);
and UO_710 (O_710,N_3004,N_2756);
or UO_711 (O_711,N_2956,N_2880);
nand UO_712 (O_712,N_3415,N_3680);
and UO_713 (O_713,N_2529,N_4382);
or UO_714 (O_714,N_2638,N_3386);
nor UO_715 (O_715,N_3509,N_3980);
nor UO_716 (O_716,N_4294,N_3298);
or UO_717 (O_717,N_2544,N_3993);
or UO_718 (O_718,N_3009,N_4153);
and UO_719 (O_719,N_4384,N_2551);
nand UO_720 (O_720,N_4192,N_3714);
nor UO_721 (O_721,N_2569,N_4870);
nand UO_722 (O_722,N_3534,N_3030);
nor UO_723 (O_723,N_2704,N_3745);
nor UO_724 (O_724,N_4410,N_2974);
and UO_725 (O_725,N_3407,N_3701);
nand UO_726 (O_726,N_4878,N_4338);
and UO_727 (O_727,N_4378,N_4571);
xor UO_728 (O_728,N_3977,N_3469);
xnor UO_729 (O_729,N_3834,N_4274);
nand UO_730 (O_730,N_3120,N_4388);
nor UO_731 (O_731,N_4683,N_3342);
xnor UO_732 (O_732,N_4819,N_2696);
xor UO_733 (O_733,N_2807,N_3068);
or UO_734 (O_734,N_4596,N_2937);
nor UO_735 (O_735,N_2728,N_2530);
or UO_736 (O_736,N_4691,N_3539);
nor UO_737 (O_737,N_3243,N_2666);
xnor UO_738 (O_738,N_4302,N_4895);
nor UO_739 (O_739,N_2536,N_3295);
or UO_740 (O_740,N_3023,N_4618);
nand UO_741 (O_741,N_4276,N_2526);
nand UO_742 (O_742,N_3189,N_2541);
and UO_743 (O_743,N_4489,N_2579);
or UO_744 (O_744,N_4671,N_4971);
nand UO_745 (O_745,N_2655,N_2733);
nand UO_746 (O_746,N_4032,N_3862);
or UO_747 (O_747,N_3442,N_4493);
nor UO_748 (O_748,N_3108,N_4792);
and UO_749 (O_749,N_4537,N_3583);
or UO_750 (O_750,N_4919,N_4899);
and UO_751 (O_751,N_4861,N_3906);
and UO_752 (O_752,N_2581,N_3839);
or UO_753 (O_753,N_4625,N_2798);
nand UO_754 (O_754,N_4303,N_2726);
and UO_755 (O_755,N_2714,N_4298);
xor UO_756 (O_756,N_3261,N_4940);
nor UO_757 (O_757,N_4327,N_4835);
nor UO_758 (O_758,N_3819,N_3121);
or UO_759 (O_759,N_3782,N_4600);
and UO_760 (O_760,N_4711,N_2825);
and UO_761 (O_761,N_3420,N_3165);
nand UO_762 (O_762,N_3492,N_2766);
nor UO_763 (O_763,N_4759,N_3787);
and UO_764 (O_764,N_3750,N_4931);
nor UO_765 (O_765,N_3912,N_3306);
and UO_766 (O_766,N_2554,N_3728);
xor UO_767 (O_767,N_3836,N_3368);
or UO_768 (O_768,N_4476,N_4136);
nor UO_769 (O_769,N_4023,N_2999);
or UO_770 (O_770,N_3490,N_4605);
nor UO_771 (O_771,N_3537,N_2794);
and UO_772 (O_772,N_3885,N_3515);
or UO_773 (O_773,N_4598,N_4473);
and UO_774 (O_774,N_4099,N_3620);
nand UO_775 (O_775,N_4348,N_3512);
nor UO_776 (O_776,N_2750,N_2747);
or UO_777 (O_777,N_4584,N_4006);
and UO_778 (O_778,N_3127,N_2763);
or UO_779 (O_779,N_3162,N_4110);
nor UO_780 (O_780,N_3796,N_2964);
nand UO_781 (O_781,N_3134,N_3790);
or UO_782 (O_782,N_3879,N_4286);
nand UO_783 (O_783,N_3203,N_2672);
nor UO_784 (O_784,N_4269,N_4495);
or UO_785 (O_785,N_3658,N_3841);
and UO_786 (O_786,N_4176,N_4871);
and UO_787 (O_787,N_3348,N_3113);
or UO_788 (O_788,N_4551,N_3083);
nor UO_789 (O_789,N_4077,N_3370);
or UO_790 (O_790,N_4522,N_2634);
or UO_791 (O_791,N_3486,N_3013);
nor UO_792 (O_792,N_3082,N_3971);
nand UO_793 (O_793,N_3724,N_4996);
nand UO_794 (O_794,N_3044,N_3835);
xor UO_795 (O_795,N_4396,N_2834);
and UO_796 (O_796,N_4853,N_2920);
nand UO_797 (O_797,N_3838,N_3809);
nor UO_798 (O_798,N_3814,N_2945);
nor UO_799 (O_799,N_3152,N_3222);
or UO_800 (O_800,N_4791,N_2848);
or UO_801 (O_801,N_3577,N_3347);
or UO_802 (O_802,N_4471,N_3938);
nor UO_803 (O_803,N_4935,N_3554);
nor UO_804 (O_804,N_3634,N_3444);
and UO_805 (O_805,N_3824,N_2755);
nand UO_806 (O_806,N_3607,N_4554);
and UO_807 (O_807,N_3783,N_4603);
nor UO_808 (O_808,N_2567,N_2679);
nand UO_809 (O_809,N_4140,N_4027);
nand UO_810 (O_810,N_3060,N_4852);
nor UO_811 (O_811,N_3283,N_3638);
nand UO_812 (O_812,N_4240,N_2577);
nand UO_813 (O_813,N_3999,N_3580);
nor UO_814 (O_814,N_4796,N_3596);
xor UO_815 (O_815,N_3688,N_2511);
or UO_816 (O_816,N_4828,N_3504);
nor UO_817 (O_817,N_2923,N_3223);
nand UO_818 (O_818,N_2742,N_3291);
or UO_819 (O_819,N_4203,N_2867);
or UO_820 (O_820,N_3920,N_4121);
or UO_821 (O_821,N_3340,N_3344);
nand UO_822 (O_822,N_4653,N_3712);
xor UO_823 (O_823,N_4456,N_3786);
nor UO_824 (O_824,N_2621,N_4003);
xnor UO_825 (O_825,N_2903,N_3687);
nand UO_826 (O_826,N_2633,N_4070);
nor UO_827 (O_827,N_4350,N_4427);
and UO_828 (O_828,N_4188,N_4293);
nor UO_829 (O_829,N_3061,N_4183);
xor UO_830 (O_830,N_4007,N_3333);
and UO_831 (O_831,N_2954,N_4602);
and UO_832 (O_832,N_4398,N_3766);
nor UO_833 (O_833,N_3097,N_4624);
nor UO_834 (O_834,N_2841,N_3646);
nand UO_835 (O_835,N_3381,N_3163);
nor UO_836 (O_836,N_4230,N_4315);
and UO_837 (O_837,N_4687,N_3406);
nor UO_838 (O_838,N_3270,N_4831);
and UO_839 (O_839,N_2661,N_3457);
nand UO_840 (O_840,N_3759,N_3916);
and UO_841 (O_841,N_4177,N_3412);
and UO_842 (O_842,N_4287,N_3066);
or UO_843 (O_843,N_3050,N_4036);
and UO_844 (O_844,N_2619,N_4362);
nor UO_845 (O_845,N_3551,N_4474);
and UO_846 (O_846,N_4254,N_2514);
xor UO_847 (O_847,N_2800,N_3631);
nor UO_848 (O_848,N_2857,N_3200);
nor UO_849 (O_849,N_4990,N_4451);
xnor UO_850 (O_850,N_4168,N_3793);
and UO_851 (O_851,N_3366,N_3474);
nand UO_852 (O_852,N_3676,N_4487);
nor UO_853 (O_853,N_3239,N_2687);
and UO_854 (O_854,N_4527,N_3437);
or UO_855 (O_855,N_3330,N_3959);
nand UO_856 (O_856,N_3294,N_4515);
or UO_857 (O_857,N_3987,N_4139);
nor UO_858 (O_858,N_2997,N_3487);
nand UO_859 (O_859,N_4146,N_4288);
or UO_860 (O_860,N_3677,N_3899);
nor UO_861 (O_861,N_3394,N_2986);
and UO_862 (O_862,N_3679,N_4030);
nand UO_863 (O_863,N_3496,N_4380);
or UO_864 (O_864,N_2826,N_3825);
or UO_865 (O_865,N_4224,N_3039);
nor UO_866 (O_866,N_4570,N_4301);
xor UO_867 (O_867,N_3360,N_3087);
nor UO_868 (O_868,N_4477,N_3095);
nand UO_869 (O_869,N_3837,N_3598);
and UO_870 (O_870,N_3387,N_3047);
nand UO_871 (O_871,N_3664,N_2912);
xor UO_872 (O_872,N_3749,N_3692);
nor UO_873 (O_873,N_4655,N_3893);
nor UO_874 (O_874,N_3180,N_3995);
or UO_875 (O_875,N_4626,N_4770);
or UO_876 (O_876,N_3725,N_4068);
and UO_877 (O_877,N_2608,N_3735);
or UO_878 (O_878,N_4408,N_3863);
nor UO_879 (O_879,N_3447,N_4172);
and UO_880 (O_880,N_2640,N_3589);
nor UO_881 (O_881,N_4241,N_4142);
nor UO_882 (O_882,N_2879,N_2681);
nor UO_883 (O_883,N_4830,N_2625);
xnor UO_884 (O_884,N_4391,N_3789);
and UO_885 (O_885,N_4054,N_4988);
nor UO_886 (O_886,N_3829,N_3846);
or UO_887 (O_887,N_4516,N_3202);
and UO_888 (O_888,N_4981,N_3198);
xnor UO_889 (O_889,N_4822,N_3106);
and UO_890 (O_890,N_3226,N_4370);
xor UO_891 (O_891,N_3967,N_4087);
xor UO_892 (O_892,N_2941,N_3069);
and UO_893 (O_893,N_2549,N_4198);
nand UO_894 (O_894,N_4575,N_3349);
nand UO_895 (O_895,N_4811,N_3593);
xnor UO_896 (O_896,N_3542,N_3210);
or UO_897 (O_897,N_2543,N_4723);
xnor UO_898 (O_898,N_3802,N_2988);
nand UO_899 (O_899,N_4672,N_3767);
and UO_900 (O_900,N_3140,N_4896);
nor UO_901 (O_901,N_3690,N_3928);
or UO_902 (O_902,N_3491,N_3876);
xor UO_903 (O_903,N_4061,N_4832);
or UO_904 (O_904,N_4645,N_2626);
nor UO_905 (O_905,N_3937,N_3826);
and UO_906 (O_906,N_3032,N_4846);
nand UO_907 (O_907,N_3764,N_4334);
and UO_908 (O_908,N_3522,N_3827);
nand UO_909 (O_909,N_4586,N_4017);
nor UO_910 (O_910,N_3170,N_4982);
nand UO_911 (O_911,N_2740,N_2809);
xnor UO_912 (O_912,N_4262,N_4734);
and UO_913 (O_913,N_2602,N_2722);
and UO_914 (O_914,N_4045,N_4520);
and UO_915 (O_915,N_2998,N_4479);
or UO_916 (O_916,N_2789,N_3247);
xnor UO_917 (O_917,N_4137,N_4798);
nor UO_918 (O_918,N_3459,N_3946);
and UO_919 (O_919,N_2906,N_3337);
xor UO_920 (O_920,N_4992,N_4331);
xnor UO_921 (O_921,N_4866,N_2611);
xor UO_922 (O_922,N_4562,N_3859);
or UO_923 (O_923,N_4161,N_2982);
and UO_924 (O_924,N_2978,N_2736);
nor UO_925 (O_925,N_4160,N_4782);
or UO_926 (O_926,N_4167,N_2649);
nor UO_927 (O_927,N_4295,N_4363);
nand UO_928 (O_928,N_2504,N_2524);
nor UO_929 (O_929,N_4332,N_4727);
nor UO_930 (O_930,N_3058,N_3932);
and UO_931 (O_931,N_3595,N_2928);
or UO_932 (O_932,N_3391,N_3409);
or UO_933 (O_933,N_3576,N_4652);
nor UO_934 (O_934,N_2613,N_2528);
nor UO_935 (O_935,N_4300,N_3744);
and UO_936 (O_936,N_4066,N_4291);
nor UO_937 (O_937,N_4670,N_3339);
nand UO_938 (O_938,N_3168,N_4132);
nand UO_939 (O_939,N_2586,N_2909);
nand UO_940 (O_940,N_3710,N_2533);
nor UO_941 (O_941,N_2641,N_2930);
and UO_942 (O_942,N_3754,N_2706);
nor UO_943 (O_943,N_3281,N_4539);
or UO_944 (O_944,N_2650,N_3652);
nor UO_945 (O_945,N_4264,N_4638);
xnor UO_946 (O_946,N_4707,N_2643);
or UO_947 (O_947,N_2965,N_4938);
nand UO_948 (O_948,N_4589,N_4898);
and UO_949 (O_949,N_4799,N_4597);
xnor UO_950 (O_950,N_2934,N_2629);
and UO_951 (O_951,N_4888,N_4445);
xor UO_952 (O_952,N_4504,N_2520);
nor UO_953 (O_953,N_3390,N_2595);
xor UO_954 (O_954,N_2902,N_4975);
nand UO_955 (O_955,N_4836,N_2571);
nor UO_956 (O_956,N_4317,N_3931);
nand UO_957 (O_957,N_2532,N_3173);
and UO_958 (O_958,N_4787,N_2580);
and UO_959 (O_959,N_3921,N_4053);
nand UO_960 (O_960,N_4692,N_4917);
xor UO_961 (O_961,N_3001,N_4599);
nand UO_962 (O_962,N_3998,N_3361);
nand UO_963 (O_963,N_3684,N_3584);
nand UO_964 (O_964,N_3956,N_3141);
nand UO_965 (O_965,N_3894,N_3227);
and UO_966 (O_966,N_2951,N_4662);
or UO_967 (O_967,N_4124,N_3875);
nor UO_968 (O_968,N_3924,N_3092);
nand UO_969 (O_969,N_2515,N_3821);
nor UO_970 (O_970,N_4046,N_3992);
xor UO_971 (O_971,N_2882,N_2538);
and UO_972 (O_972,N_3627,N_4421);
and UO_973 (O_973,N_3630,N_3772);
and UO_974 (O_974,N_3272,N_4984);
or UO_975 (O_975,N_2838,N_3678);
nand UO_976 (O_976,N_3628,N_3035);
nand UO_977 (O_977,N_2688,N_4193);
or UO_978 (O_978,N_3500,N_3571);
and UO_979 (O_979,N_3260,N_4801);
or UO_980 (O_980,N_4523,N_4532);
and UO_981 (O_981,N_3721,N_3454);
or UO_982 (O_982,N_4747,N_4854);
nor UO_983 (O_983,N_4634,N_3989);
nand UO_984 (O_984,N_3557,N_2874);
nor UO_985 (O_985,N_4088,N_2843);
or UO_986 (O_986,N_2955,N_2989);
and UO_987 (O_987,N_4436,N_4767);
or UO_988 (O_988,N_2980,N_4156);
nor UO_989 (O_989,N_4699,N_3318);
nand UO_990 (O_990,N_4337,N_3953);
nand UO_991 (O_991,N_4755,N_3708);
nand UO_992 (O_992,N_4848,N_4951);
or UO_993 (O_993,N_3794,N_4306);
or UO_994 (O_994,N_3861,N_3352);
nor UO_995 (O_995,N_3350,N_4480);
nor UO_996 (O_996,N_3644,N_4581);
or UO_997 (O_997,N_3408,N_3619);
and UO_998 (O_998,N_2905,N_3311);
nor UO_999 (O_999,N_3532,N_3629);
endmodule