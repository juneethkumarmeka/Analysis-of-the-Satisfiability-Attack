module basic_500_3000_500_30_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_113,In_21);
nand U1 (N_1,In_482,In_495);
nand U2 (N_2,In_467,In_297);
nor U3 (N_3,In_3,In_180);
xor U4 (N_4,In_497,In_314);
and U5 (N_5,In_192,In_289);
nor U6 (N_6,In_84,In_191);
nor U7 (N_7,In_353,In_278);
nor U8 (N_8,In_169,In_105);
nor U9 (N_9,In_351,In_398);
nor U10 (N_10,In_262,In_446);
nor U11 (N_11,In_315,In_494);
nand U12 (N_12,In_20,In_32);
or U13 (N_13,In_340,In_111);
nor U14 (N_14,In_442,In_496);
and U15 (N_15,In_368,In_190);
and U16 (N_16,In_292,In_52);
nor U17 (N_17,In_293,In_498);
or U18 (N_18,In_316,In_490);
nor U19 (N_19,In_261,In_11);
or U20 (N_20,In_233,In_164);
nand U21 (N_21,In_59,In_361);
or U22 (N_22,In_13,In_188);
nand U23 (N_23,In_265,In_218);
or U24 (N_24,In_165,In_109);
nand U25 (N_25,In_324,In_88);
nand U26 (N_26,In_147,In_350);
nand U27 (N_27,In_7,In_44);
or U28 (N_28,In_43,In_499);
nor U29 (N_29,In_267,In_156);
nand U30 (N_30,In_15,In_187);
nor U31 (N_31,In_341,In_214);
and U32 (N_32,In_372,In_354);
nand U33 (N_33,In_250,In_357);
or U34 (N_34,In_79,In_37);
nor U35 (N_35,In_19,In_390);
or U36 (N_36,In_27,In_256);
or U37 (N_37,In_260,In_428);
nand U38 (N_38,In_308,In_312);
and U39 (N_39,In_142,In_396);
nand U40 (N_40,In_42,In_17);
and U41 (N_41,In_334,In_458);
nand U42 (N_42,In_376,In_290);
or U43 (N_43,In_210,In_269);
nor U44 (N_44,In_223,In_444);
and U45 (N_45,In_206,In_374);
nand U46 (N_46,In_101,In_33);
nand U47 (N_47,In_159,In_434);
nor U48 (N_48,In_182,In_384);
nand U49 (N_49,In_46,In_65);
nand U50 (N_50,In_411,In_453);
nor U51 (N_51,In_451,In_115);
nand U52 (N_52,In_108,In_454);
nand U53 (N_53,In_204,In_323);
or U54 (N_54,In_440,In_282);
or U55 (N_55,In_415,In_221);
nand U56 (N_56,In_227,In_201);
and U57 (N_57,In_141,In_209);
or U58 (N_58,In_380,In_254);
and U59 (N_59,In_53,In_18);
or U60 (N_60,In_72,In_386);
nor U61 (N_61,In_75,In_445);
nor U62 (N_62,In_177,In_421);
nor U63 (N_63,In_220,In_329);
and U64 (N_64,In_345,In_270);
and U65 (N_65,In_419,In_364);
or U66 (N_66,In_60,In_122);
and U67 (N_67,In_279,In_58);
or U68 (N_68,In_130,In_34);
and U69 (N_69,In_51,In_479);
or U70 (N_70,In_45,In_459);
or U71 (N_71,In_333,In_68);
nor U72 (N_72,In_346,In_127);
nand U73 (N_73,In_143,In_394);
nor U74 (N_74,In_28,In_248);
nand U75 (N_75,In_62,In_129);
nor U76 (N_76,In_197,In_242);
nor U77 (N_77,In_36,In_401);
nor U78 (N_78,In_429,In_41);
nand U79 (N_79,In_66,In_366);
nor U80 (N_80,In_311,In_492);
nor U81 (N_81,In_12,In_480);
or U82 (N_82,In_230,In_234);
and U83 (N_83,In_2,In_4);
nor U84 (N_84,In_47,In_54);
and U85 (N_85,In_456,In_275);
nand U86 (N_86,In_400,In_94);
nand U87 (N_87,In_304,In_22);
or U88 (N_88,In_14,In_322);
xor U89 (N_89,In_483,In_102);
nand U90 (N_90,In_76,In_395);
and U91 (N_91,In_306,In_356);
or U92 (N_92,In_154,In_119);
nand U93 (N_93,In_493,In_291);
or U94 (N_94,In_186,In_399);
or U95 (N_95,In_121,In_245);
or U96 (N_96,In_131,In_416);
nor U97 (N_97,In_420,In_126);
and U98 (N_98,In_358,In_484);
or U99 (N_99,In_303,In_287);
nor U100 (N_100,N_57,In_77);
nand U101 (N_101,N_44,In_157);
nand U102 (N_102,N_73,In_486);
nand U103 (N_103,In_388,In_447);
and U104 (N_104,N_9,In_194);
nand U105 (N_105,In_202,In_26);
nand U106 (N_106,In_410,In_295);
nor U107 (N_107,In_99,In_475);
or U108 (N_108,N_58,In_48);
nor U109 (N_109,In_104,In_81);
nand U110 (N_110,In_403,N_69);
nor U111 (N_111,In_189,In_407);
or U112 (N_112,In_163,In_235);
and U113 (N_113,In_307,In_213);
or U114 (N_114,In_240,N_16);
or U115 (N_115,In_405,In_120);
and U116 (N_116,In_472,In_63);
nor U117 (N_117,N_80,In_413);
and U118 (N_118,N_22,In_418);
nor U119 (N_119,In_298,N_40);
or U120 (N_120,In_8,In_320);
or U121 (N_121,In_309,In_431);
nand U122 (N_122,In_302,N_28);
xor U123 (N_123,N_63,In_263);
or U124 (N_124,N_99,In_425);
nor U125 (N_125,In_69,In_408);
nor U126 (N_126,In_469,In_125);
nand U127 (N_127,In_424,In_31);
nor U128 (N_128,In_319,In_225);
or U129 (N_129,In_412,In_171);
or U130 (N_130,In_463,In_117);
nor U131 (N_131,In_237,N_43);
nand U132 (N_132,In_266,In_73);
nand U133 (N_133,N_96,In_488);
or U134 (N_134,In_461,In_193);
or U135 (N_135,In_236,In_82);
nor U136 (N_136,In_56,In_93);
and U137 (N_137,In_359,In_100);
and U138 (N_138,In_369,N_30);
nand U139 (N_139,In_228,In_352);
nand U140 (N_140,In_133,In_149);
nand U141 (N_141,N_86,In_466);
nand U142 (N_142,In_160,In_229);
nand U143 (N_143,In_150,In_325);
or U144 (N_144,N_52,N_68);
or U145 (N_145,In_216,N_98);
or U146 (N_146,In_281,In_86);
and U147 (N_147,In_478,In_35);
or U148 (N_148,In_310,In_183);
or U149 (N_149,In_387,N_77);
nor U150 (N_150,In_389,N_27);
nor U151 (N_151,In_55,N_78);
and U152 (N_152,In_299,In_30);
nor U153 (N_153,In_208,In_199);
nor U154 (N_154,In_371,In_367);
or U155 (N_155,N_39,In_70);
and U156 (N_156,In_327,In_383);
nor U157 (N_157,In_116,N_76);
or U158 (N_158,In_326,N_53);
or U159 (N_159,N_26,In_378);
nand U160 (N_160,In_257,In_140);
and U161 (N_161,N_11,N_70);
nand U162 (N_162,In_264,In_243);
and U163 (N_163,N_2,In_404);
or U164 (N_164,In_487,In_476);
nor U165 (N_165,In_460,In_244);
nand U166 (N_166,In_450,In_335);
or U167 (N_167,In_377,In_96);
nand U168 (N_168,In_226,In_285);
nand U169 (N_169,In_222,In_328);
xnor U170 (N_170,In_184,In_74);
or U171 (N_171,N_23,In_370);
or U172 (N_172,In_249,In_238);
and U173 (N_173,In_144,N_64);
nor U174 (N_174,N_97,N_21);
nand U175 (N_175,In_426,N_0);
nor U176 (N_176,In_16,N_41);
nor U177 (N_177,N_14,In_112);
or U178 (N_178,In_300,N_1);
nand U179 (N_179,In_132,In_146);
nand U180 (N_180,In_305,N_34);
or U181 (N_181,In_318,N_61);
nand U182 (N_182,In_332,In_6);
nand U183 (N_183,N_45,In_203);
or U184 (N_184,N_38,N_84);
nor U185 (N_185,In_83,In_465);
and U186 (N_186,In_135,In_462);
or U187 (N_187,In_385,In_107);
xnor U188 (N_188,In_301,In_471);
nand U189 (N_189,In_241,In_381);
and U190 (N_190,N_42,In_178);
nor U191 (N_191,N_49,In_71);
and U192 (N_192,In_137,In_284);
and U193 (N_193,In_61,In_153);
nor U194 (N_194,In_283,N_95);
nor U195 (N_195,N_19,In_215);
and U196 (N_196,In_491,In_170);
nor U197 (N_197,In_24,N_79);
nand U198 (N_198,In_80,In_106);
or U199 (N_199,N_51,In_176);
nand U200 (N_200,In_118,In_355);
and U201 (N_201,N_180,N_66);
nor U202 (N_202,N_54,N_102);
and U203 (N_203,In_9,In_406);
nand U204 (N_204,N_48,N_132);
nor U205 (N_205,In_155,N_156);
and U206 (N_206,In_198,N_128);
or U207 (N_207,In_375,In_441);
nor U208 (N_208,N_159,In_255);
nand U209 (N_209,N_101,In_64);
and U210 (N_210,In_414,In_246);
nor U211 (N_211,N_186,N_117);
and U212 (N_212,N_130,N_91);
or U213 (N_213,In_391,In_252);
nand U214 (N_214,N_164,In_481);
and U215 (N_215,In_151,N_124);
nor U216 (N_216,N_151,In_457);
nand U217 (N_217,N_111,In_138);
nor U218 (N_218,In_449,N_174);
or U219 (N_219,N_137,In_172);
nand U220 (N_220,In_392,N_47);
or U221 (N_221,N_182,N_170);
nor U222 (N_222,In_436,N_192);
and U223 (N_223,In_379,In_67);
or U224 (N_224,In_336,In_87);
and U225 (N_225,In_470,N_140);
and U226 (N_226,In_338,In_273);
nor U227 (N_227,N_158,N_37);
and U228 (N_228,In_342,In_339);
and U229 (N_229,In_435,In_474);
nor U230 (N_230,In_212,N_110);
nor U231 (N_231,In_331,In_162);
or U232 (N_232,N_176,N_100);
nor U233 (N_233,N_75,In_224);
or U234 (N_234,In_253,In_288);
nor U235 (N_235,N_33,N_104);
nor U236 (N_236,N_74,In_468);
nand U237 (N_237,N_29,In_57);
nor U238 (N_238,N_36,N_162);
or U239 (N_239,N_108,N_152);
or U240 (N_240,In_373,In_1);
nand U241 (N_241,In_433,N_173);
nand U242 (N_242,N_15,In_485);
nand U243 (N_243,N_184,N_187);
and U244 (N_244,In_409,In_97);
and U245 (N_245,N_146,N_87);
and U246 (N_246,In_181,In_382);
nand U247 (N_247,In_473,In_402);
or U248 (N_248,N_185,N_177);
nor U249 (N_249,N_120,N_35);
or U250 (N_250,In_231,N_149);
nor U251 (N_251,N_82,N_179);
nand U252 (N_252,N_31,N_60);
or U253 (N_253,In_423,N_13);
and U254 (N_254,N_134,N_183);
nand U255 (N_255,N_90,In_29);
and U256 (N_256,In_128,N_93);
and U257 (N_257,N_168,In_437);
or U258 (N_258,In_274,In_179);
and U259 (N_259,N_190,N_167);
and U260 (N_260,In_232,N_7);
and U261 (N_261,In_175,In_438);
nand U262 (N_262,N_171,In_38);
nand U263 (N_263,In_167,N_178);
and U264 (N_264,In_271,In_337);
nor U265 (N_265,N_138,In_25);
and U266 (N_266,N_67,In_259);
or U267 (N_267,In_95,In_39);
nand U268 (N_268,In_123,N_160);
and U269 (N_269,N_144,N_165);
nor U270 (N_270,N_8,In_78);
nand U271 (N_271,In_363,In_348);
and U272 (N_272,In_349,N_3);
or U273 (N_273,In_360,N_195);
nand U274 (N_274,In_10,N_6);
nand U275 (N_275,In_85,N_143);
and U276 (N_276,N_103,N_71);
nand U277 (N_277,In_49,In_422);
and U278 (N_278,N_88,N_56);
nor U279 (N_279,In_313,In_5);
nor U280 (N_280,In_280,N_81);
nand U281 (N_281,N_199,In_239);
nor U282 (N_282,N_17,N_5);
or U283 (N_283,In_219,N_20);
nor U284 (N_284,In_343,In_152);
and U285 (N_285,N_94,In_452);
nand U286 (N_286,N_65,In_134);
nor U287 (N_287,N_25,In_397);
nor U288 (N_288,N_121,In_432);
nand U289 (N_289,In_455,N_119);
nand U290 (N_290,In_347,In_110);
nor U291 (N_291,In_330,N_59);
and U292 (N_292,N_188,In_92);
and U293 (N_293,In_195,In_148);
and U294 (N_294,In_98,In_443);
nor U295 (N_295,N_163,In_196);
nand U296 (N_296,N_112,In_251);
and U297 (N_297,N_145,In_344);
or U298 (N_298,In_489,In_174);
and U299 (N_299,N_12,In_40);
or U300 (N_300,N_268,N_92);
or U301 (N_301,N_212,N_166);
and U302 (N_302,N_105,N_267);
nand U303 (N_303,N_200,N_155);
or U304 (N_304,In_317,N_250);
or U305 (N_305,N_270,N_215);
nand U306 (N_306,N_32,N_229);
or U307 (N_307,N_225,N_283);
nor U308 (N_308,In_448,N_271);
nor U309 (N_309,N_246,N_169);
nand U310 (N_310,N_50,N_213);
and U311 (N_311,N_263,N_154);
and U312 (N_312,N_197,N_109);
nor U313 (N_313,N_266,N_290);
and U314 (N_314,N_289,N_247);
or U315 (N_315,N_115,N_224);
and U316 (N_316,In_417,In_427);
and U317 (N_317,In_136,In_91);
and U318 (N_318,In_430,N_211);
and U319 (N_319,N_237,In_124);
nor U320 (N_320,N_295,In_294);
nor U321 (N_321,N_280,In_145);
nand U322 (N_322,N_214,N_258);
or U323 (N_323,N_249,N_253);
nand U324 (N_324,N_234,N_85);
nor U325 (N_325,N_122,N_259);
or U326 (N_326,N_296,N_281);
or U327 (N_327,N_18,N_248);
nor U328 (N_328,In_166,N_286);
or U329 (N_329,N_228,N_265);
and U330 (N_330,N_125,N_298);
and U331 (N_331,N_208,In_286);
and U332 (N_332,In_114,N_216);
nor U333 (N_333,N_191,N_175);
and U334 (N_334,In_362,N_209);
and U335 (N_335,In_217,In_139);
nor U336 (N_336,N_113,N_181);
and U337 (N_337,N_89,N_218);
or U338 (N_338,In_365,N_141);
nor U339 (N_339,In_477,N_172);
nand U340 (N_340,N_157,N_142);
nor U341 (N_341,In_50,N_284);
nand U342 (N_342,N_232,In_321);
nand U343 (N_343,N_217,In_439);
nand U344 (N_344,N_219,N_133);
nand U345 (N_345,N_24,N_148);
and U346 (N_346,N_193,N_261);
or U347 (N_347,N_251,N_278);
and U348 (N_348,N_226,N_83);
or U349 (N_349,N_243,In_90);
or U350 (N_350,N_254,In_89);
xor U351 (N_351,N_221,N_131);
nand U352 (N_352,N_127,N_239);
or U353 (N_353,N_294,In_211);
nand U354 (N_354,N_252,N_257);
nor U355 (N_355,N_236,N_288);
nand U356 (N_356,N_279,N_126);
and U357 (N_357,N_231,N_244);
and U358 (N_358,N_272,In_268);
or U359 (N_359,N_287,N_72);
and U360 (N_360,N_241,N_136);
or U361 (N_361,N_118,N_260);
nand U362 (N_362,N_206,N_275);
nand U363 (N_363,In_161,N_238);
nand U364 (N_364,In_205,N_205);
or U365 (N_365,In_173,N_242);
xnor U366 (N_366,In_272,N_114);
and U367 (N_367,In_276,N_204);
nand U368 (N_368,N_222,N_153);
or U369 (N_369,N_240,N_46);
nand U370 (N_370,N_227,In_103);
and U371 (N_371,In_258,N_233);
nand U372 (N_372,N_256,N_223);
nand U373 (N_373,N_220,N_196);
nor U374 (N_374,N_189,N_264);
nand U375 (N_375,N_282,N_269);
nand U376 (N_376,N_292,N_62);
nor U377 (N_377,In_247,N_161);
nand U378 (N_378,In_158,N_150);
nand U379 (N_379,In_207,In_23);
and U380 (N_380,In_0,N_147);
nand U381 (N_381,N_230,N_129);
nand U382 (N_382,N_107,In_277);
nor U383 (N_383,N_194,N_135);
or U384 (N_384,N_299,N_55);
and U385 (N_385,N_203,N_273);
or U386 (N_386,N_235,N_274);
and U387 (N_387,N_291,In_296);
and U388 (N_388,N_276,N_207);
and U389 (N_389,N_255,N_139);
or U390 (N_390,In_168,In_393);
nor U391 (N_391,N_285,N_262);
nor U392 (N_392,N_123,N_116);
or U393 (N_393,N_202,In_464);
nand U394 (N_394,N_10,N_293);
nand U395 (N_395,N_201,N_210);
and U396 (N_396,N_297,N_245);
nor U397 (N_397,N_4,N_198);
and U398 (N_398,N_106,In_185);
nor U399 (N_399,N_277,In_200);
and U400 (N_400,N_354,N_314);
nor U401 (N_401,N_323,N_332);
nand U402 (N_402,N_322,N_360);
or U403 (N_403,N_316,N_315);
nor U404 (N_404,N_309,N_356);
nand U405 (N_405,N_374,N_306);
nand U406 (N_406,N_398,N_383);
and U407 (N_407,N_329,N_325);
or U408 (N_408,N_328,N_326);
or U409 (N_409,N_357,N_385);
nor U410 (N_410,N_376,N_351);
nand U411 (N_411,N_352,N_367);
nor U412 (N_412,N_393,N_361);
or U413 (N_413,N_342,N_386);
and U414 (N_414,N_304,N_395);
or U415 (N_415,N_381,N_391);
and U416 (N_416,N_305,N_303);
or U417 (N_417,N_380,N_349);
or U418 (N_418,N_327,N_343);
and U419 (N_419,N_339,N_301);
nand U420 (N_420,N_390,N_344);
nor U421 (N_421,N_338,N_370);
nand U422 (N_422,N_377,N_369);
or U423 (N_423,N_336,N_384);
nor U424 (N_424,N_397,N_366);
nand U425 (N_425,N_312,N_313);
or U426 (N_426,N_330,N_368);
and U427 (N_427,N_379,N_371);
nand U428 (N_428,N_307,N_387);
and U429 (N_429,N_355,N_375);
and U430 (N_430,N_302,N_363);
nand U431 (N_431,N_321,N_319);
nand U432 (N_432,N_324,N_348);
nand U433 (N_433,N_362,N_341);
or U434 (N_434,N_317,N_347);
nand U435 (N_435,N_373,N_353);
nor U436 (N_436,N_320,N_333);
nor U437 (N_437,N_345,N_318);
nor U438 (N_438,N_340,N_394);
or U439 (N_439,N_364,N_310);
and U440 (N_440,N_372,N_382);
or U441 (N_441,N_334,N_365);
nand U442 (N_442,N_346,N_335);
or U443 (N_443,N_396,N_399);
or U444 (N_444,N_308,N_392);
and U445 (N_445,N_331,N_378);
or U446 (N_446,N_359,N_300);
and U447 (N_447,N_389,N_358);
or U448 (N_448,N_350,N_311);
nand U449 (N_449,N_337,N_388);
and U450 (N_450,N_301,N_359);
or U451 (N_451,N_326,N_388);
and U452 (N_452,N_342,N_395);
nand U453 (N_453,N_309,N_307);
nor U454 (N_454,N_333,N_330);
nand U455 (N_455,N_371,N_303);
and U456 (N_456,N_353,N_305);
nand U457 (N_457,N_374,N_359);
nor U458 (N_458,N_388,N_385);
nand U459 (N_459,N_331,N_395);
and U460 (N_460,N_388,N_375);
or U461 (N_461,N_342,N_371);
nand U462 (N_462,N_385,N_372);
nand U463 (N_463,N_350,N_372);
and U464 (N_464,N_390,N_341);
nor U465 (N_465,N_362,N_336);
or U466 (N_466,N_310,N_379);
nand U467 (N_467,N_359,N_368);
nand U468 (N_468,N_311,N_371);
nand U469 (N_469,N_323,N_380);
or U470 (N_470,N_378,N_379);
nand U471 (N_471,N_345,N_382);
and U472 (N_472,N_325,N_381);
nor U473 (N_473,N_370,N_353);
nand U474 (N_474,N_389,N_363);
nor U475 (N_475,N_372,N_369);
nor U476 (N_476,N_374,N_347);
nor U477 (N_477,N_391,N_363);
nand U478 (N_478,N_381,N_346);
or U479 (N_479,N_357,N_345);
and U480 (N_480,N_341,N_373);
nor U481 (N_481,N_302,N_309);
or U482 (N_482,N_363,N_349);
and U483 (N_483,N_352,N_346);
and U484 (N_484,N_358,N_365);
and U485 (N_485,N_399,N_360);
nand U486 (N_486,N_308,N_342);
or U487 (N_487,N_317,N_386);
nand U488 (N_488,N_342,N_353);
and U489 (N_489,N_355,N_328);
nand U490 (N_490,N_372,N_379);
nor U491 (N_491,N_366,N_314);
nor U492 (N_492,N_384,N_333);
nor U493 (N_493,N_399,N_317);
or U494 (N_494,N_394,N_304);
nor U495 (N_495,N_359,N_364);
nor U496 (N_496,N_329,N_345);
nand U497 (N_497,N_336,N_369);
nand U498 (N_498,N_336,N_312);
nand U499 (N_499,N_366,N_339);
and U500 (N_500,N_449,N_475);
and U501 (N_501,N_433,N_445);
nand U502 (N_502,N_409,N_410);
nand U503 (N_503,N_420,N_468);
nor U504 (N_504,N_426,N_477);
and U505 (N_505,N_481,N_456);
and U506 (N_506,N_499,N_432);
nand U507 (N_507,N_446,N_440);
or U508 (N_508,N_494,N_462);
or U509 (N_509,N_415,N_439);
and U510 (N_510,N_427,N_438);
nor U511 (N_511,N_469,N_478);
nand U512 (N_512,N_464,N_428);
or U513 (N_513,N_425,N_453);
and U514 (N_514,N_421,N_455);
or U515 (N_515,N_490,N_492);
nand U516 (N_516,N_422,N_495);
or U517 (N_517,N_473,N_488);
nor U518 (N_518,N_487,N_401);
nand U519 (N_519,N_450,N_454);
nand U520 (N_520,N_457,N_480);
or U521 (N_521,N_461,N_436);
or U522 (N_522,N_402,N_491);
and U523 (N_523,N_448,N_443);
nand U524 (N_524,N_463,N_465);
nand U525 (N_525,N_431,N_498);
or U526 (N_526,N_419,N_485);
nor U527 (N_527,N_400,N_437);
and U528 (N_528,N_496,N_403);
nand U529 (N_529,N_412,N_406);
or U530 (N_530,N_486,N_405);
nand U531 (N_531,N_470,N_417);
nand U532 (N_532,N_458,N_424);
nand U533 (N_533,N_467,N_484);
nor U534 (N_534,N_479,N_460);
nor U535 (N_535,N_447,N_483);
nand U536 (N_536,N_416,N_435);
nand U537 (N_537,N_423,N_418);
nand U538 (N_538,N_459,N_493);
nand U539 (N_539,N_472,N_404);
nand U540 (N_540,N_497,N_474);
nor U541 (N_541,N_441,N_476);
nand U542 (N_542,N_452,N_407);
and U543 (N_543,N_444,N_408);
or U544 (N_544,N_451,N_482);
nand U545 (N_545,N_442,N_413);
and U546 (N_546,N_489,N_471);
and U547 (N_547,N_429,N_430);
nand U548 (N_548,N_466,N_411);
and U549 (N_549,N_414,N_434);
nor U550 (N_550,N_441,N_408);
nand U551 (N_551,N_419,N_454);
or U552 (N_552,N_411,N_467);
or U553 (N_553,N_442,N_454);
nand U554 (N_554,N_464,N_451);
nand U555 (N_555,N_426,N_432);
and U556 (N_556,N_402,N_424);
xnor U557 (N_557,N_429,N_441);
nor U558 (N_558,N_432,N_429);
nor U559 (N_559,N_404,N_471);
nand U560 (N_560,N_407,N_439);
or U561 (N_561,N_460,N_411);
or U562 (N_562,N_458,N_462);
nand U563 (N_563,N_453,N_427);
nor U564 (N_564,N_430,N_408);
nor U565 (N_565,N_443,N_498);
and U566 (N_566,N_481,N_497);
or U567 (N_567,N_438,N_477);
and U568 (N_568,N_483,N_497);
and U569 (N_569,N_486,N_491);
and U570 (N_570,N_496,N_409);
nor U571 (N_571,N_417,N_486);
or U572 (N_572,N_474,N_417);
and U573 (N_573,N_463,N_479);
and U574 (N_574,N_415,N_443);
or U575 (N_575,N_465,N_455);
and U576 (N_576,N_480,N_494);
or U577 (N_577,N_465,N_499);
nand U578 (N_578,N_464,N_445);
nor U579 (N_579,N_499,N_449);
and U580 (N_580,N_458,N_402);
and U581 (N_581,N_433,N_407);
and U582 (N_582,N_429,N_409);
or U583 (N_583,N_455,N_498);
nor U584 (N_584,N_452,N_451);
nand U585 (N_585,N_429,N_417);
nor U586 (N_586,N_462,N_463);
nor U587 (N_587,N_402,N_414);
nor U588 (N_588,N_416,N_467);
and U589 (N_589,N_467,N_455);
nor U590 (N_590,N_460,N_496);
nand U591 (N_591,N_486,N_404);
or U592 (N_592,N_433,N_458);
nor U593 (N_593,N_442,N_485);
nand U594 (N_594,N_431,N_425);
nand U595 (N_595,N_463,N_403);
nor U596 (N_596,N_419,N_409);
or U597 (N_597,N_410,N_404);
and U598 (N_598,N_460,N_476);
nor U599 (N_599,N_400,N_492);
nor U600 (N_600,N_572,N_516);
or U601 (N_601,N_569,N_584);
and U602 (N_602,N_534,N_506);
and U603 (N_603,N_573,N_541);
nand U604 (N_604,N_591,N_528);
or U605 (N_605,N_564,N_545);
and U606 (N_606,N_514,N_589);
and U607 (N_607,N_505,N_550);
nand U608 (N_608,N_592,N_561);
nand U609 (N_609,N_533,N_570);
nand U610 (N_610,N_518,N_594);
and U611 (N_611,N_511,N_542);
nand U612 (N_612,N_537,N_504);
nand U613 (N_613,N_515,N_595);
or U614 (N_614,N_520,N_508);
and U615 (N_615,N_576,N_500);
or U616 (N_616,N_563,N_574);
or U617 (N_617,N_587,N_560);
and U618 (N_618,N_517,N_598);
nand U619 (N_619,N_543,N_524);
nor U620 (N_620,N_531,N_548);
nand U621 (N_621,N_580,N_581);
nand U622 (N_622,N_513,N_549);
nand U623 (N_623,N_551,N_544);
nand U624 (N_624,N_510,N_582);
nor U625 (N_625,N_559,N_502);
nand U626 (N_626,N_540,N_583);
or U627 (N_627,N_554,N_535);
and U628 (N_628,N_536,N_512);
or U629 (N_629,N_590,N_503);
nor U630 (N_630,N_597,N_553);
nand U631 (N_631,N_562,N_526);
nor U632 (N_632,N_565,N_523);
and U633 (N_633,N_530,N_577);
or U634 (N_634,N_555,N_519);
nor U635 (N_635,N_556,N_552);
and U636 (N_636,N_507,N_571);
or U637 (N_637,N_566,N_575);
nand U638 (N_638,N_547,N_579);
nor U639 (N_639,N_522,N_585);
or U640 (N_640,N_568,N_501);
nor U641 (N_641,N_593,N_586);
nor U642 (N_642,N_532,N_596);
or U643 (N_643,N_527,N_599);
or U644 (N_644,N_578,N_538);
or U645 (N_645,N_525,N_529);
nor U646 (N_646,N_567,N_558);
nand U647 (N_647,N_557,N_539);
and U648 (N_648,N_509,N_546);
nand U649 (N_649,N_588,N_521);
and U650 (N_650,N_521,N_556);
nor U651 (N_651,N_566,N_541);
nand U652 (N_652,N_543,N_587);
nand U653 (N_653,N_529,N_503);
nor U654 (N_654,N_518,N_556);
nor U655 (N_655,N_511,N_585);
and U656 (N_656,N_595,N_522);
nand U657 (N_657,N_569,N_553);
and U658 (N_658,N_515,N_555);
nand U659 (N_659,N_583,N_572);
nand U660 (N_660,N_525,N_522);
and U661 (N_661,N_577,N_529);
and U662 (N_662,N_500,N_521);
and U663 (N_663,N_557,N_598);
nand U664 (N_664,N_576,N_508);
nor U665 (N_665,N_501,N_534);
or U666 (N_666,N_511,N_535);
and U667 (N_667,N_517,N_530);
or U668 (N_668,N_528,N_552);
nand U669 (N_669,N_553,N_534);
and U670 (N_670,N_563,N_567);
and U671 (N_671,N_554,N_536);
nand U672 (N_672,N_568,N_571);
nor U673 (N_673,N_549,N_568);
nor U674 (N_674,N_532,N_539);
nor U675 (N_675,N_511,N_517);
nor U676 (N_676,N_595,N_511);
nor U677 (N_677,N_573,N_556);
nor U678 (N_678,N_501,N_550);
or U679 (N_679,N_537,N_519);
nand U680 (N_680,N_522,N_530);
nand U681 (N_681,N_508,N_545);
nor U682 (N_682,N_510,N_553);
nand U683 (N_683,N_590,N_509);
nor U684 (N_684,N_569,N_517);
or U685 (N_685,N_534,N_503);
nand U686 (N_686,N_567,N_555);
nor U687 (N_687,N_513,N_581);
nand U688 (N_688,N_567,N_595);
nand U689 (N_689,N_554,N_524);
or U690 (N_690,N_557,N_500);
nand U691 (N_691,N_528,N_547);
nand U692 (N_692,N_568,N_557);
nor U693 (N_693,N_594,N_500);
nand U694 (N_694,N_545,N_540);
or U695 (N_695,N_588,N_585);
or U696 (N_696,N_533,N_500);
nor U697 (N_697,N_537,N_542);
nor U698 (N_698,N_556,N_563);
or U699 (N_699,N_562,N_566);
or U700 (N_700,N_651,N_630);
nand U701 (N_701,N_628,N_637);
xor U702 (N_702,N_690,N_622);
nand U703 (N_703,N_634,N_666);
and U704 (N_704,N_633,N_624);
nand U705 (N_705,N_686,N_638);
and U706 (N_706,N_604,N_656);
nand U707 (N_707,N_611,N_613);
and U708 (N_708,N_639,N_606);
and U709 (N_709,N_674,N_645);
nor U710 (N_710,N_697,N_664);
and U711 (N_711,N_657,N_626);
and U712 (N_712,N_643,N_654);
and U713 (N_713,N_629,N_625);
nor U714 (N_714,N_678,N_688);
or U715 (N_715,N_670,N_675);
nand U716 (N_716,N_648,N_682);
or U717 (N_717,N_641,N_698);
nand U718 (N_718,N_607,N_658);
and U719 (N_719,N_677,N_696);
nor U720 (N_720,N_650,N_621);
or U721 (N_721,N_640,N_644);
or U722 (N_722,N_659,N_687);
or U723 (N_723,N_676,N_627);
or U724 (N_724,N_691,N_681);
nor U725 (N_725,N_695,N_636);
nor U726 (N_726,N_608,N_673);
or U727 (N_727,N_679,N_684);
nor U728 (N_728,N_623,N_601);
nor U729 (N_729,N_694,N_620);
or U730 (N_730,N_662,N_665);
nor U731 (N_731,N_647,N_689);
nor U732 (N_732,N_663,N_699);
nand U733 (N_733,N_680,N_610);
nand U734 (N_734,N_660,N_602);
and U735 (N_735,N_652,N_631);
nand U736 (N_736,N_619,N_632);
and U737 (N_737,N_671,N_661);
or U738 (N_738,N_612,N_617);
nand U739 (N_739,N_603,N_600);
and U740 (N_740,N_667,N_605);
nand U741 (N_741,N_693,N_683);
and U742 (N_742,N_672,N_685);
and U743 (N_743,N_655,N_635);
nand U744 (N_744,N_616,N_668);
nor U745 (N_745,N_642,N_609);
and U746 (N_746,N_618,N_653);
and U747 (N_747,N_692,N_649);
or U748 (N_748,N_669,N_614);
nor U749 (N_749,N_615,N_646);
and U750 (N_750,N_658,N_699);
nor U751 (N_751,N_688,N_639);
nor U752 (N_752,N_625,N_634);
nor U753 (N_753,N_603,N_640);
nor U754 (N_754,N_627,N_655);
and U755 (N_755,N_657,N_654);
and U756 (N_756,N_638,N_637);
and U757 (N_757,N_685,N_639);
nor U758 (N_758,N_617,N_697);
nor U759 (N_759,N_676,N_629);
nand U760 (N_760,N_682,N_615);
and U761 (N_761,N_601,N_667);
nand U762 (N_762,N_600,N_660);
nor U763 (N_763,N_644,N_623);
or U764 (N_764,N_698,N_673);
nand U765 (N_765,N_668,N_620);
or U766 (N_766,N_632,N_622);
or U767 (N_767,N_688,N_611);
or U768 (N_768,N_679,N_681);
nand U769 (N_769,N_684,N_635);
nor U770 (N_770,N_675,N_630);
or U771 (N_771,N_626,N_644);
nand U772 (N_772,N_680,N_675);
nand U773 (N_773,N_639,N_682);
nor U774 (N_774,N_665,N_616);
nand U775 (N_775,N_679,N_600);
nor U776 (N_776,N_679,N_696);
or U777 (N_777,N_665,N_683);
nor U778 (N_778,N_615,N_668);
or U779 (N_779,N_638,N_612);
or U780 (N_780,N_643,N_667);
or U781 (N_781,N_663,N_600);
and U782 (N_782,N_631,N_633);
nand U783 (N_783,N_606,N_619);
nor U784 (N_784,N_684,N_657);
nor U785 (N_785,N_634,N_607);
and U786 (N_786,N_652,N_607);
nand U787 (N_787,N_624,N_626);
nand U788 (N_788,N_647,N_638);
nand U789 (N_789,N_640,N_668);
nand U790 (N_790,N_656,N_694);
or U791 (N_791,N_665,N_659);
nand U792 (N_792,N_688,N_658);
nand U793 (N_793,N_651,N_696);
or U794 (N_794,N_621,N_674);
or U795 (N_795,N_664,N_694);
and U796 (N_796,N_664,N_657);
and U797 (N_797,N_623,N_621);
nor U798 (N_798,N_653,N_690);
nor U799 (N_799,N_659,N_675);
or U800 (N_800,N_759,N_730);
nor U801 (N_801,N_768,N_796);
nor U802 (N_802,N_760,N_720);
nand U803 (N_803,N_704,N_703);
or U804 (N_804,N_795,N_773);
and U805 (N_805,N_749,N_755);
or U806 (N_806,N_788,N_753);
xor U807 (N_807,N_729,N_706);
or U808 (N_808,N_734,N_797);
and U809 (N_809,N_792,N_743);
or U810 (N_810,N_772,N_751);
nor U811 (N_811,N_722,N_791);
nor U812 (N_812,N_745,N_779);
nand U813 (N_813,N_765,N_783);
or U814 (N_814,N_776,N_762);
and U815 (N_815,N_787,N_711);
nor U816 (N_816,N_769,N_732);
or U817 (N_817,N_798,N_780);
nor U818 (N_818,N_712,N_728);
and U819 (N_819,N_746,N_715);
nand U820 (N_820,N_747,N_721);
or U821 (N_821,N_713,N_758);
and U822 (N_822,N_754,N_710);
nand U823 (N_823,N_750,N_742);
nor U824 (N_824,N_719,N_764);
xnor U825 (N_825,N_735,N_785);
or U826 (N_826,N_786,N_702);
nand U827 (N_827,N_744,N_741);
nand U828 (N_828,N_716,N_774);
nand U829 (N_829,N_714,N_718);
or U830 (N_830,N_731,N_723);
and U831 (N_831,N_733,N_717);
or U832 (N_832,N_738,N_782);
or U833 (N_833,N_790,N_736);
and U834 (N_834,N_727,N_705);
nand U835 (N_835,N_781,N_766);
or U836 (N_836,N_793,N_748);
and U837 (N_837,N_700,N_739);
and U838 (N_838,N_771,N_757);
nor U839 (N_839,N_752,N_756);
nand U840 (N_840,N_737,N_709);
nand U841 (N_841,N_707,N_740);
and U842 (N_842,N_799,N_761);
and U843 (N_843,N_708,N_770);
and U844 (N_844,N_726,N_775);
nand U845 (N_845,N_724,N_789);
and U846 (N_846,N_763,N_725);
or U847 (N_847,N_794,N_767);
and U848 (N_848,N_777,N_701);
or U849 (N_849,N_784,N_778);
and U850 (N_850,N_711,N_773);
nor U851 (N_851,N_727,N_754);
nor U852 (N_852,N_727,N_747);
and U853 (N_853,N_718,N_797);
or U854 (N_854,N_791,N_741);
nor U855 (N_855,N_735,N_701);
and U856 (N_856,N_786,N_797);
nor U857 (N_857,N_761,N_723);
or U858 (N_858,N_783,N_738);
and U859 (N_859,N_741,N_796);
and U860 (N_860,N_711,N_734);
nand U861 (N_861,N_721,N_755);
nand U862 (N_862,N_766,N_755);
or U863 (N_863,N_717,N_766);
and U864 (N_864,N_735,N_787);
and U865 (N_865,N_779,N_703);
nand U866 (N_866,N_709,N_718);
nand U867 (N_867,N_792,N_736);
and U868 (N_868,N_745,N_750);
or U869 (N_869,N_782,N_704);
and U870 (N_870,N_747,N_728);
and U871 (N_871,N_743,N_731);
nand U872 (N_872,N_736,N_795);
nor U873 (N_873,N_767,N_736);
nand U874 (N_874,N_782,N_722);
and U875 (N_875,N_741,N_780);
and U876 (N_876,N_726,N_793);
and U877 (N_877,N_792,N_793);
or U878 (N_878,N_743,N_740);
nand U879 (N_879,N_754,N_738);
nand U880 (N_880,N_730,N_726);
nand U881 (N_881,N_738,N_798);
and U882 (N_882,N_798,N_719);
and U883 (N_883,N_709,N_731);
nand U884 (N_884,N_715,N_784);
and U885 (N_885,N_737,N_797);
or U886 (N_886,N_786,N_716);
nor U887 (N_887,N_771,N_729);
nand U888 (N_888,N_714,N_715);
and U889 (N_889,N_789,N_747);
nand U890 (N_890,N_738,N_766);
and U891 (N_891,N_790,N_758);
nor U892 (N_892,N_778,N_776);
and U893 (N_893,N_739,N_776);
and U894 (N_894,N_767,N_766);
and U895 (N_895,N_778,N_733);
nand U896 (N_896,N_771,N_790);
nor U897 (N_897,N_761,N_750);
nand U898 (N_898,N_768,N_737);
and U899 (N_899,N_726,N_766);
nand U900 (N_900,N_844,N_859);
nand U901 (N_901,N_848,N_874);
nor U902 (N_902,N_864,N_866);
nor U903 (N_903,N_876,N_807);
or U904 (N_904,N_825,N_818);
and U905 (N_905,N_860,N_875);
nor U906 (N_906,N_853,N_899);
nor U907 (N_907,N_879,N_808);
and U908 (N_908,N_854,N_823);
nand U909 (N_909,N_885,N_819);
nand U910 (N_910,N_824,N_805);
and U911 (N_911,N_845,N_842);
nor U912 (N_912,N_894,N_852);
and U913 (N_913,N_858,N_802);
nor U914 (N_914,N_813,N_811);
nand U915 (N_915,N_889,N_816);
or U916 (N_916,N_809,N_868);
and U917 (N_917,N_861,N_806);
nand U918 (N_918,N_878,N_887);
nand U919 (N_919,N_877,N_826);
or U920 (N_920,N_814,N_800);
xor U921 (N_921,N_890,N_888);
or U922 (N_922,N_839,N_822);
or U923 (N_923,N_886,N_863);
and U924 (N_924,N_855,N_873);
nor U925 (N_925,N_830,N_891);
or U926 (N_926,N_893,N_827);
nand U927 (N_927,N_829,N_812);
or U928 (N_928,N_835,N_862);
nor U929 (N_929,N_801,N_831);
nor U930 (N_930,N_838,N_850);
and U931 (N_931,N_872,N_832);
nor U932 (N_932,N_897,N_865);
nor U933 (N_933,N_836,N_841);
nand U934 (N_934,N_851,N_810);
or U935 (N_935,N_834,N_898);
nor U936 (N_936,N_815,N_833);
nor U937 (N_937,N_846,N_870);
or U938 (N_938,N_871,N_880);
and U939 (N_939,N_820,N_881);
nor U940 (N_940,N_803,N_843);
nand U941 (N_941,N_869,N_837);
or U942 (N_942,N_883,N_817);
or U943 (N_943,N_882,N_856);
nor U944 (N_944,N_896,N_849);
nand U945 (N_945,N_804,N_828);
nor U946 (N_946,N_840,N_892);
nand U947 (N_947,N_884,N_895);
nor U948 (N_948,N_821,N_857);
nor U949 (N_949,N_867,N_847);
nor U950 (N_950,N_864,N_899);
and U951 (N_951,N_889,N_884);
nor U952 (N_952,N_883,N_875);
nor U953 (N_953,N_869,N_817);
or U954 (N_954,N_838,N_830);
and U955 (N_955,N_854,N_842);
or U956 (N_956,N_828,N_826);
nor U957 (N_957,N_889,N_818);
or U958 (N_958,N_859,N_831);
and U959 (N_959,N_871,N_893);
or U960 (N_960,N_872,N_804);
and U961 (N_961,N_882,N_845);
or U962 (N_962,N_822,N_876);
and U963 (N_963,N_872,N_890);
nand U964 (N_964,N_823,N_893);
nor U965 (N_965,N_829,N_890);
nor U966 (N_966,N_886,N_816);
and U967 (N_967,N_870,N_827);
nand U968 (N_968,N_826,N_889);
and U969 (N_969,N_809,N_869);
nor U970 (N_970,N_874,N_881);
or U971 (N_971,N_881,N_816);
and U972 (N_972,N_872,N_825);
or U973 (N_973,N_881,N_889);
or U974 (N_974,N_882,N_804);
and U975 (N_975,N_872,N_843);
nand U976 (N_976,N_801,N_804);
nor U977 (N_977,N_843,N_822);
nand U978 (N_978,N_860,N_851);
nor U979 (N_979,N_882,N_809);
or U980 (N_980,N_895,N_854);
or U981 (N_981,N_808,N_876);
nand U982 (N_982,N_839,N_883);
nor U983 (N_983,N_829,N_811);
or U984 (N_984,N_844,N_881);
or U985 (N_985,N_845,N_889);
and U986 (N_986,N_860,N_838);
nand U987 (N_987,N_877,N_866);
or U988 (N_988,N_817,N_889);
nand U989 (N_989,N_849,N_821);
xnor U990 (N_990,N_841,N_881);
nor U991 (N_991,N_858,N_861);
nand U992 (N_992,N_837,N_843);
or U993 (N_993,N_808,N_856);
or U994 (N_994,N_833,N_877);
nor U995 (N_995,N_898,N_895);
or U996 (N_996,N_866,N_850);
nor U997 (N_997,N_803,N_833);
or U998 (N_998,N_848,N_817);
nand U999 (N_999,N_860,N_845);
nor U1000 (N_1000,N_999,N_973);
or U1001 (N_1001,N_927,N_906);
and U1002 (N_1002,N_970,N_985);
xor U1003 (N_1003,N_902,N_943);
nor U1004 (N_1004,N_916,N_904);
nor U1005 (N_1005,N_963,N_921);
and U1006 (N_1006,N_991,N_928);
xor U1007 (N_1007,N_926,N_956);
nand U1008 (N_1008,N_961,N_930);
and U1009 (N_1009,N_944,N_932);
and U1010 (N_1010,N_912,N_974);
nand U1011 (N_1011,N_957,N_938);
or U1012 (N_1012,N_942,N_900);
nand U1013 (N_1013,N_982,N_946);
nor U1014 (N_1014,N_964,N_952);
and U1015 (N_1015,N_978,N_992);
and U1016 (N_1016,N_975,N_920);
nor U1017 (N_1017,N_979,N_922);
nor U1018 (N_1018,N_993,N_987);
or U1019 (N_1019,N_937,N_905);
or U1020 (N_1020,N_955,N_996);
and U1021 (N_1021,N_924,N_949);
and U1022 (N_1022,N_910,N_909);
and U1023 (N_1023,N_951,N_994);
and U1024 (N_1024,N_933,N_977);
and U1025 (N_1025,N_984,N_936);
and U1026 (N_1026,N_998,N_959);
and U1027 (N_1027,N_929,N_931);
nor U1028 (N_1028,N_969,N_947);
nand U1029 (N_1029,N_948,N_903);
and U1030 (N_1030,N_950,N_935);
nor U1031 (N_1031,N_953,N_995);
or U1032 (N_1032,N_986,N_983);
nand U1033 (N_1033,N_917,N_989);
or U1034 (N_1034,N_967,N_976);
and U1035 (N_1035,N_919,N_962);
nand U1036 (N_1036,N_923,N_907);
nor U1037 (N_1037,N_945,N_980);
or U1038 (N_1038,N_925,N_997);
nor U1039 (N_1039,N_988,N_913);
nand U1040 (N_1040,N_966,N_908);
nand U1041 (N_1041,N_981,N_990);
nand U1042 (N_1042,N_940,N_901);
nand U1043 (N_1043,N_965,N_918);
nand U1044 (N_1044,N_939,N_972);
and U1045 (N_1045,N_960,N_914);
nor U1046 (N_1046,N_915,N_968);
nand U1047 (N_1047,N_954,N_911);
nor U1048 (N_1048,N_934,N_971);
and U1049 (N_1049,N_941,N_958);
nand U1050 (N_1050,N_970,N_924);
or U1051 (N_1051,N_945,N_914);
nor U1052 (N_1052,N_957,N_934);
nor U1053 (N_1053,N_943,N_921);
nor U1054 (N_1054,N_901,N_930);
nand U1055 (N_1055,N_902,N_942);
nand U1056 (N_1056,N_970,N_998);
nor U1057 (N_1057,N_927,N_972);
or U1058 (N_1058,N_939,N_996);
nor U1059 (N_1059,N_962,N_986);
or U1060 (N_1060,N_943,N_993);
nor U1061 (N_1061,N_924,N_991);
or U1062 (N_1062,N_982,N_969);
or U1063 (N_1063,N_921,N_924);
nand U1064 (N_1064,N_904,N_996);
nand U1065 (N_1065,N_979,N_991);
and U1066 (N_1066,N_979,N_963);
or U1067 (N_1067,N_956,N_996);
nand U1068 (N_1068,N_936,N_950);
and U1069 (N_1069,N_939,N_905);
nor U1070 (N_1070,N_984,N_951);
nand U1071 (N_1071,N_978,N_988);
or U1072 (N_1072,N_954,N_936);
nand U1073 (N_1073,N_984,N_966);
and U1074 (N_1074,N_905,N_993);
or U1075 (N_1075,N_978,N_972);
or U1076 (N_1076,N_936,N_905);
xor U1077 (N_1077,N_982,N_955);
nand U1078 (N_1078,N_997,N_944);
nor U1079 (N_1079,N_961,N_955);
nand U1080 (N_1080,N_970,N_978);
or U1081 (N_1081,N_949,N_973);
or U1082 (N_1082,N_927,N_925);
or U1083 (N_1083,N_909,N_991);
nor U1084 (N_1084,N_934,N_940);
nor U1085 (N_1085,N_924,N_951);
nor U1086 (N_1086,N_981,N_924);
or U1087 (N_1087,N_908,N_995);
or U1088 (N_1088,N_999,N_946);
and U1089 (N_1089,N_952,N_947);
nand U1090 (N_1090,N_997,N_990);
and U1091 (N_1091,N_916,N_987);
nor U1092 (N_1092,N_932,N_982);
nor U1093 (N_1093,N_937,N_948);
and U1094 (N_1094,N_982,N_936);
or U1095 (N_1095,N_941,N_910);
and U1096 (N_1096,N_955,N_991);
nand U1097 (N_1097,N_912,N_978);
nand U1098 (N_1098,N_924,N_939);
nand U1099 (N_1099,N_905,N_972);
and U1100 (N_1100,N_1091,N_1048);
nor U1101 (N_1101,N_1028,N_1098);
nand U1102 (N_1102,N_1031,N_1090);
and U1103 (N_1103,N_1050,N_1002);
nand U1104 (N_1104,N_1088,N_1063);
and U1105 (N_1105,N_1055,N_1067);
xor U1106 (N_1106,N_1081,N_1046);
nand U1107 (N_1107,N_1058,N_1013);
and U1108 (N_1108,N_1042,N_1009);
and U1109 (N_1109,N_1059,N_1017);
or U1110 (N_1110,N_1086,N_1078);
or U1111 (N_1111,N_1073,N_1043);
and U1112 (N_1112,N_1052,N_1023);
or U1113 (N_1113,N_1062,N_1076);
nand U1114 (N_1114,N_1030,N_1071);
nand U1115 (N_1115,N_1053,N_1094);
or U1116 (N_1116,N_1039,N_1047);
nand U1117 (N_1117,N_1003,N_1000);
and U1118 (N_1118,N_1065,N_1049);
nand U1119 (N_1119,N_1001,N_1034);
nand U1120 (N_1120,N_1012,N_1096);
nor U1121 (N_1121,N_1082,N_1064);
nor U1122 (N_1122,N_1041,N_1054);
nor U1123 (N_1123,N_1021,N_1040);
nor U1124 (N_1124,N_1015,N_1026);
or U1125 (N_1125,N_1056,N_1087);
and U1126 (N_1126,N_1070,N_1080);
or U1127 (N_1127,N_1085,N_1024);
nor U1128 (N_1128,N_1038,N_1079);
or U1129 (N_1129,N_1016,N_1025);
or U1130 (N_1130,N_1092,N_1032);
and U1131 (N_1131,N_1060,N_1008);
nand U1132 (N_1132,N_1097,N_1036);
or U1133 (N_1133,N_1084,N_1019);
and U1134 (N_1134,N_1004,N_1011);
or U1135 (N_1135,N_1044,N_1075);
and U1136 (N_1136,N_1057,N_1029);
nand U1137 (N_1137,N_1099,N_1006);
nand U1138 (N_1138,N_1033,N_1061);
nand U1139 (N_1139,N_1093,N_1037);
nor U1140 (N_1140,N_1020,N_1068);
or U1141 (N_1141,N_1018,N_1083);
and U1142 (N_1142,N_1077,N_1089);
and U1143 (N_1143,N_1007,N_1005);
nand U1144 (N_1144,N_1051,N_1072);
nand U1145 (N_1145,N_1074,N_1022);
and U1146 (N_1146,N_1014,N_1095);
and U1147 (N_1147,N_1045,N_1066);
nor U1148 (N_1148,N_1010,N_1027);
nand U1149 (N_1149,N_1035,N_1069);
or U1150 (N_1150,N_1085,N_1019);
nand U1151 (N_1151,N_1005,N_1015);
nand U1152 (N_1152,N_1042,N_1019);
or U1153 (N_1153,N_1041,N_1015);
nand U1154 (N_1154,N_1030,N_1059);
nand U1155 (N_1155,N_1066,N_1018);
nand U1156 (N_1156,N_1048,N_1096);
nand U1157 (N_1157,N_1060,N_1006);
and U1158 (N_1158,N_1019,N_1076);
or U1159 (N_1159,N_1029,N_1070);
or U1160 (N_1160,N_1046,N_1088);
nand U1161 (N_1161,N_1022,N_1075);
nor U1162 (N_1162,N_1084,N_1080);
or U1163 (N_1163,N_1009,N_1021);
or U1164 (N_1164,N_1012,N_1018);
and U1165 (N_1165,N_1079,N_1056);
or U1166 (N_1166,N_1050,N_1038);
nand U1167 (N_1167,N_1017,N_1022);
nand U1168 (N_1168,N_1063,N_1037);
or U1169 (N_1169,N_1033,N_1041);
xnor U1170 (N_1170,N_1063,N_1034);
and U1171 (N_1171,N_1037,N_1061);
nor U1172 (N_1172,N_1053,N_1054);
and U1173 (N_1173,N_1083,N_1027);
or U1174 (N_1174,N_1094,N_1082);
nand U1175 (N_1175,N_1038,N_1036);
or U1176 (N_1176,N_1010,N_1066);
nor U1177 (N_1177,N_1056,N_1028);
and U1178 (N_1178,N_1005,N_1023);
nor U1179 (N_1179,N_1039,N_1077);
nor U1180 (N_1180,N_1023,N_1082);
or U1181 (N_1181,N_1055,N_1033);
nand U1182 (N_1182,N_1090,N_1072);
or U1183 (N_1183,N_1006,N_1018);
and U1184 (N_1184,N_1031,N_1034);
nor U1185 (N_1185,N_1033,N_1058);
nand U1186 (N_1186,N_1032,N_1056);
and U1187 (N_1187,N_1085,N_1066);
or U1188 (N_1188,N_1005,N_1071);
or U1189 (N_1189,N_1049,N_1007);
nor U1190 (N_1190,N_1069,N_1011);
or U1191 (N_1191,N_1063,N_1056);
nand U1192 (N_1192,N_1091,N_1018);
nand U1193 (N_1193,N_1000,N_1053);
nor U1194 (N_1194,N_1011,N_1032);
and U1195 (N_1195,N_1003,N_1069);
or U1196 (N_1196,N_1043,N_1008);
and U1197 (N_1197,N_1014,N_1033);
nand U1198 (N_1198,N_1026,N_1065);
nor U1199 (N_1199,N_1046,N_1079);
or U1200 (N_1200,N_1111,N_1129);
nor U1201 (N_1201,N_1141,N_1150);
or U1202 (N_1202,N_1145,N_1155);
nor U1203 (N_1203,N_1149,N_1159);
nor U1204 (N_1204,N_1184,N_1146);
or U1205 (N_1205,N_1119,N_1126);
nor U1206 (N_1206,N_1198,N_1185);
and U1207 (N_1207,N_1144,N_1168);
nand U1208 (N_1208,N_1164,N_1107);
and U1209 (N_1209,N_1113,N_1140);
nor U1210 (N_1210,N_1188,N_1151);
nor U1211 (N_1211,N_1163,N_1137);
nand U1212 (N_1212,N_1131,N_1166);
nand U1213 (N_1213,N_1192,N_1101);
nand U1214 (N_1214,N_1123,N_1172);
nor U1215 (N_1215,N_1118,N_1193);
nor U1216 (N_1216,N_1143,N_1197);
nor U1217 (N_1217,N_1152,N_1124);
and U1218 (N_1218,N_1153,N_1139);
nor U1219 (N_1219,N_1102,N_1196);
and U1220 (N_1220,N_1154,N_1173);
or U1221 (N_1221,N_1132,N_1183);
and U1222 (N_1222,N_1156,N_1178);
nor U1223 (N_1223,N_1104,N_1186);
or U1224 (N_1224,N_1105,N_1117);
nor U1225 (N_1225,N_1180,N_1100);
and U1226 (N_1226,N_1109,N_1170);
and U1227 (N_1227,N_1121,N_1116);
nor U1228 (N_1228,N_1157,N_1127);
nand U1229 (N_1229,N_1176,N_1165);
or U1230 (N_1230,N_1182,N_1138);
and U1231 (N_1231,N_1161,N_1158);
and U1232 (N_1232,N_1114,N_1110);
nor U1233 (N_1233,N_1133,N_1120);
and U1234 (N_1234,N_1174,N_1167);
nor U1235 (N_1235,N_1115,N_1103);
or U1236 (N_1236,N_1142,N_1125);
or U1237 (N_1237,N_1147,N_1195);
nand U1238 (N_1238,N_1108,N_1136);
xor U1239 (N_1239,N_1134,N_1171);
nand U1240 (N_1240,N_1199,N_1181);
nand U1241 (N_1241,N_1190,N_1112);
nor U1242 (N_1242,N_1177,N_1162);
and U1243 (N_1243,N_1189,N_1179);
nand U1244 (N_1244,N_1175,N_1128);
nor U1245 (N_1245,N_1135,N_1194);
nor U1246 (N_1246,N_1191,N_1169);
or U1247 (N_1247,N_1130,N_1122);
nand U1248 (N_1248,N_1148,N_1106);
or U1249 (N_1249,N_1187,N_1160);
and U1250 (N_1250,N_1199,N_1131);
or U1251 (N_1251,N_1112,N_1104);
or U1252 (N_1252,N_1160,N_1155);
or U1253 (N_1253,N_1133,N_1183);
or U1254 (N_1254,N_1196,N_1182);
and U1255 (N_1255,N_1135,N_1127);
or U1256 (N_1256,N_1153,N_1195);
or U1257 (N_1257,N_1128,N_1139);
nand U1258 (N_1258,N_1182,N_1108);
or U1259 (N_1259,N_1127,N_1164);
and U1260 (N_1260,N_1157,N_1185);
or U1261 (N_1261,N_1164,N_1131);
or U1262 (N_1262,N_1183,N_1126);
nor U1263 (N_1263,N_1116,N_1143);
nand U1264 (N_1264,N_1129,N_1159);
nand U1265 (N_1265,N_1149,N_1134);
and U1266 (N_1266,N_1164,N_1126);
and U1267 (N_1267,N_1164,N_1122);
nand U1268 (N_1268,N_1143,N_1127);
or U1269 (N_1269,N_1111,N_1162);
or U1270 (N_1270,N_1116,N_1157);
or U1271 (N_1271,N_1118,N_1150);
nor U1272 (N_1272,N_1196,N_1197);
nand U1273 (N_1273,N_1166,N_1139);
and U1274 (N_1274,N_1145,N_1139);
nand U1275 (N_1275,N_1185,N_1153);
and U1276 (N_1276,N_1198,N_1128);
nor U1277 (N_1277,N_1103,N_1164);
nor U1278 (N_1278,N_1147,N_1151);
nor U1279 (N_1279,N_1144,N_1122);
nand U1280 (N_1280,N_1198,N_1120);
and U1281 (N_1281,N_1121,N_1175);
or U1282 (N_1282,N_1125,N_1120);
nand U1283 (N_1283,N_1124,N_1114);
nand U1284 (N_1284,N_1167,N_1169);
nor U1285 (N_1285,N_1169,N_1183);
nor U1286 (N_1286,N_1109,N_1130);
and U1287 (N_1287,N_1112,N_1137);
and U1288 (N_1288,N_1152,N_1156);
nor U1289 (N_1289,N_1106,N_1104);
and U1290 (N_1290,N_1174,N_1191);
nand U1291 (N_1291,N_1143,N_1189);
and U1292 (N_1292,N_1144,N_1152);
and U1293 (N_1293,N_1132,N_1143);
nand U1294 (N_1294,N_1174,N_1131);
and U1295 (N_1295,N_1152,N_1138);
or U1296 (N_1296,N_1124,N_1162);
and U1297 (N_1297,N_1178,N_1132);
nand U1298 (N_1298,N_1157,N_1163);
and U1299 (N_1299,N_1175,N_1182);
nor U1300 (N_1300,N_1285,N_1214);
nand U1301 (N_1301,N_1276,N_1211);
and U1302 (N_1302,N_1228,N_1215);
nor U1303 (N_1303,N_1289,N_1297);
and U1304 (N_1304,N_1263,N_1246);
nor U1305 (N_1305,N_1227,N_1238);
and U1306 (N_1306,N_1281,N_1222);
or U1307 (N_1307,N_1232,N_1288);
and U1308 (N_1308,N_1226,N_1266);
nor U1309 (N_1309,N_1219,N_1207);
nor U1310 (N_1310,N_1242,N_1223);
or U1311 (N_1311,N_1230,N_1251);
or U1312 (N_1312,N_1259,N_1254);
and U1313 (N_1313,N_1241,N_1255);
nor U1314 (N_1314,N_1204,N_1256);
nor U1315 (N_1315,N_1200,N_1293);
nand U1316 (N_1316,N_1291,N_1239);
or U1317 (N_1317,N_1220,N_1249);
or U1318 (N_1318,N_1234,N_1244);
nand U1319 (N_1319,N_1265,N_1257);
or U1320 (N_1320,N_1235,N_1210);
and U1321 (N_1321,N_1299,N_1217);
nor U1322 (N_1322,N_1264,N_1233);
nor U1323 (N_1323,N_1286,N_1274);
and U1324 (N_1324,N_1279,N_1272);
or U1325 (N_1325,N_1203,N_1296);
nand U1326 (N_1326,N_1282,N_1284);
or U1327 (N_1327,N_1271,N_1270);
nand U1328 (N_1328,N_1205,N_1201);
nand U1329 (N_1329,N_1248,N_1261);
nor U1330 (N_1330,N_1206,N_1225);
and U1331 (N_1331,N_1237,N_1252);
and U1332 (N_1332,N_1277,N_1262);
and U1333 (N_1333,N_1298,N_1290);
nor U1334 (N_1334,N_1212,N_1269);
xnor U1335 (N_1335,N_1243,N_1213);
nor U1336 (N_1336,N_1229,N_1273);
or U1337 (N_1337,N_1202,N_1283);
nand U1338 (N_1338,N_1236,N_1292);
nor U1339 (N_1339,N_1253,N_1240);
nand U1340 (N_1340,N_1258,N_1275);
nand U1341 (N_1341,N_1268,N_1295);
nand U1342 (N_1342,N_1250,N_1224);
nand U1343 (N_1343,N_1209,N_1260);
nor U1344 (N_1344,N_1216,N_1208);
or U1345 (N_1345,N_1287,N_1294);
nor U1346 (N_1346,N_1245,N_1278);
and U1347 (N_1347,N_1280,N_1267);
or U1348 (N_1348,N_1221,N_1231);
nand U1349 (N_1349,N_1247,N_1218);
nor U1350 (N_1350,N_1240,N_1265);
nor U1351 (N_1351,N_1238,N_1261);
nor U1352 (N_1352,N_1233,N_1270);
nor U1353 (N_1353,N_1284,N_1291);
nor U1354 (N_1354,N_1230,N_1243);
or U1355 (N_1355,N_1221,N_1211);
nand U1356 (N_1356,N_1299,N_1231);
and U1357 (N_1357,N_1297,N_1245);
or U1358 (N_1358,N_1210,N_1283);
nor U1359 (N_1359,N_1288,N_1290);
nor U1360 (N_1360,N_1242,N_1255);
and U1361 (N_1361,N_1283,N_1274);
and U1362 (N_1362,N_1230,N_1244);
nand U1363 (N_1363,N_1237,N_1226);
or U1364 (N_1364,N_1226,N_1256);
nand U1365 (N_1365,N_1261,N_1274);
nand U1366 (N_1366,N_1234,N_1286);
nand U1367 (N_1367,N_1204,N_1221);
and U1368 (N_1368,N_1252,N_1299);
nor U1369 (N_1369,N_1254,N_1221);
nor U1370 (N_1370,N_1203,N_1205);
and U1371 (N_1371,N_1202,N_1224);
nand U1372 (N_1372,N_1269,N_1271);
and U1373 (N_1373,N_1229,N_1277);
or U1374 (N_1374,N_1245,N_1273);
nand U1375 (N_1375,N_1249,N_1291);
nor U1376 (N_1376,N_1226,N_1275);
nand U1377 (N_1377,N_1222,N_1234);
or U1378 (N_1378,N_1205,N_1269);
nor U1379 (N_1379,N_1296,N_1225);
nand U1380 (N_1380,N_1225,N_1264);
or U1381 (N_1381,N_1266,N_1221);
nor U1382 (N_1382,N_1252,N_1251);
nand U1383 (N_1383,N_1209,N_1278);
or U1384 (N_1384,N_1256,N_1250);
or U1385 (N_1385,N_1234,N_1203);
or U1386 (N_1386,N_1278,N_1286);
or U1387 (N_1387,N_1255,N_1259);
or U1388 (N_1388,N_1219,N_1298);
and U1389 (N_1389,N_1297,N_1223);
and U1390 (N_1390,N_1273,N_1284);
and U1391 (N_1391,N_1250,N_1204);
or U1392 (N_1392,N_1286,N_1233);
nand U1393 (N_1393,N_1222,N_1233);
nor U1394 (N_1394,N_1285,N_1241);
and U1395 (N_1395,N_1224,N_1215);
nand U1396 (N_1396,N_1225,N_1275);
nand U1397 (N_1397,N_1287,N_1222);
or U1398 (N_1398,N_1242,N_1240);
and U1399 (N_1399,N_1224,N_1292);
nor U1400 (N_1400,N_1363,N_1320);
or U1401 (N_1401,N_1378,N_1360);
or U1402 (N_1402,N_1355,N_1335);
or U1403 (N_1403,N_1380,N_1377);
nand U1404 (N_1404,N_1328,N_1385);
and U1405 (N_1405,N_1395,N_1382);
or U1406 (N_1406,N_1301,N_1332);
or U1407 (N_1407,N_1351,N_1352);
or U1408 (N_1408,N_1367,N_1373);
nand U1409 (N_1409,N_1396,N_1312);
or U1410 (N_1410,N_1305,N_1383);
and U1411 (N_1411,N_1311,N_1323);
and U1412 (N_1412,N_1309,N_1322);
nor U1413 (N_1413,N_1321,N_1303);
nor U1414 (N_1414,N_1313,N_1310);
nand U1415 (N_1415,N_1381,N_1343);
nand U1416 (N_1416,N_1329,N_1386);
nor U1417 (N_1417,N_1336,N_1338);
nor U1418 (N_1418,N_1318,N_1370);
or U1419 (N_1419,N_1344,N_1349);
nor U1420 (N_1420,N_1327,N_1362);
nor U1421 (N_1421,N_1326,N_1307);
and U1422 (N_1422,N_1398,N_1334);
and U1423 (N_1423,N_1356,N_1353);
nand U1424 (N_1424,N_1348,N_1333);
and U1425 (N_1425,N_1388,N_1390);
nor U1426 (N_1426,N_1316,N_1399);
nor U1427 (N_1427,N_1337,N_1372);
nand U1428 (N_1428,N_1317,N_1308);
or U1429 (N_1429,N_1315,N_1319);
nor U1430 (N_1430,N_1341,N_1325);
nand U1431 (N_1431,N_1371,N_1364);
nand U1432 (N_1432,N_1366,N_1339);
and U1433 (N_1433,N_1314,N_1342);
or U1434 (N_1434,N_1330,N_1379);
nand U1435 (N_1435,N_1387,N_1306);
nand U1436 (N_1436,N_1347,N_1391);
and U1437 (N_1437,N_1392,N_1304);
and U1438 (N_1438,N_1350,N_1302);
and U1439 (N_1439,N_1345,N_1358);
and U1440 (N_1440,N_1369,N_1324);
and U1441 (N_1441,N_1340,N_1393);
and U1442 (N_1442,N_1300,N_1365);
or U1443 (N_1443,N_1376,N_1331);
nand U1444 (N_1444,N_1361,N_1346);
nor U1445 (N_1445,N_1394,N_1375);
nand U1446 (N_1446,N_1374,N_1384);
or U1447 (N_1447,N_1354,N_1397);
nor U1448 (N_1448,N_1357,N_1368);
nand U1449 (N_1449,N_1359,N_1389);
nand U1450 (N_1450,N_1382,N_1374);
and U1451 (N_1451,N_1348,N_1374);
or U1452 (N_1452,N_1325,N_1345);
nor U1453 (N_1453,N_1329,N_1355);
nand U1454 (N_1454,N_1322,N_1371);
or U1455 (N_1455,N_1348,N_1388);
or U1456 (N_1456,N_1322,N_1348);
and U1457 (N_1457,N_1349,N_1341);
nor U1458 (N_1458,N_1380,N_1339);
nor U1459 (N_1459,N_1368,N_1335);
and U1460 (N_1460,N_1388,N_1313);
nand U1461 (N_1461,N_1381,N_1332);
nor U1462 (N_1462,N_1339,N_1361);
nand U1463 (N_1463,N_1315,N_1337);
or U1464 (N_1464,N_1382,N_1348);
nor U1465 (N_1465,N_1395,N_1330);
nor U1466 (N_1466,N_1326,N_1317);
xor U1467 (N_1467,N_1327,N_1349);
nor U1468 (N_1468,N_1376,N_1347);
or U1469 (N_1469,N_1362,N_1380);
nand U1470 (N_1470,N_1330,N_1303);
nor U1471 (N_1471,N_1383,N_1318);
nand U1472 (N_1472,N_1367,N_1383);
or U1473 (N_1473,N_1329,N_1396);
xnor U1474 (N_1474,N_1348,N_1366);
and U1475 (N_1475,N_1354,N_1344);
nor U1476 (N_1476,N_1312,N_1379);
xnor U1477 (N_1477,N_1316,N_1308);
or U1478 (N_1478,N_1344,N_1310);
nand U1479 (N_1479,N_1367,N_1372);
or U1480 (N_1480,N_1335,N_1308);
nor U1481 (N_1481,N_1366,N_1335);
and U1482 (N_1482,N_1344,N_1335);
or U1483 (N_1483,N_1335,N_1317);
nor U1484 (N_1484,N_1370,N_1350);
nor U1485 (N_1485,N_1311,N_1362);
and U1486 (N_1486,N_1357,N_1313);
and U1487 (N_1487,N_1348,N_1395);
nor U1488 (N_1488,N_1303,N_1343);
or U1489 (N_1489,N_1342,N_1310);
and U1490 (N_1490,N_1386,N_1356);
nor U1491 (N_1491,N_1380,N_1357);
or U1492 (N_1492,N_1301,N_1348);
or U1493 (N_1493,N_1395,N_1356);
or U1494 (N_1494,N_1338,N_1319);
and U1495 (N_1495,N_1318,N_1369);
nor U1496 (N_1496,N_1315,N_1394);
and U1497 (N_1497,N_1344,N_1395);
nand U1498 (N_1498,N_1367,N_1313);
nand U1499 (N_1499,N_1357,N_1342);
or U1500 (N_1500,N_1496,N_1405);
nand U1501 (N_1501,N_1474,N_1456);
nor U1502 (N_1502,N_1445,N_1483);
nor U1503 (N_1503,N_1420,N_1413);
nand U1504 (N_1504,N_1434,N_1455);
nand U1505 (N_1505,N_1416,N_1460);
nand U1506 (N_1506,N_1424,N_1427);
or U1507 (N_1507,N_1442,N_1495);
nor U1508 (N_1508,N_1418,N_1476);
or U1509 (N_1509,N_1459,N_1446);
or U1510 (N_1510,N_1473,N_1431);
or U1511 (N_1511,N_1480,N_1410);
and U1512 (N_1512,N_1419,N_1436);
xor U1513 (N_1513,N_1406,N_1440);
and U1514 (N_1514,N_1449,N_1429);
nor U1515 (N_1515,N_1485,N_1407);
nor U1516 (N_1516,N_1494,N_1428);
or U1517 (N_1517,N_1452,N_1443);
nand U1518 (N_1518,N_1477,N_1461);
nand U1519 (N_1519,N_1402,N_1403);
nand U1520 (N_1520,N_1411,N_1422);
or U1521 (N_1521,N_1448,N_1464);
or U1522 (N_1522,N_1438,N_1453);
nor U1523 (N_1523,N_1491,N_1475);
and U1524 (N_1524,N_1486,N_1426);
nand U1525 (N_1525,N_1417,N_1421);
nand U1526 (N_1526,N_1482,N_1490);
nand U1527 (N_1527,N_1470,N_1484);
nor U1528 (N_1528,N_1404,N_1454);
and U1529 (N_1529,N_1415,N_1412);
and U1530 (N_1530,N_1466,N_1463);
or U1531 (N_1531,N_1499,N_1457);
and U1532 (N_1532,N_1401,N_1472);
or U1533 (N_1533,N_1432,N_1469);
nand U1534 (N_1534,N_1487,N_1468);
nand U1535 (N_1535,N_1414,N_1492);
or U1536 (N_1536,N_1498,N_1451);
or U1537 (N_1537,N_1430,N_1425);
nor U1538 (N_1538,N_1435,N_1467);
or U1539 (N_1539,N_1493,N_1433);
or U1540 (N_1540,N_1400,N_1423);
nand U1541 (N_1541,N_1444,N_1437);
nor U1542 (N_1542,N_1489,N_1450);
nand U1543 (N_1543,N_1478,N_1409);
nand U1544 (N_1544,N_1471,N_1479);
and U1545 (N_1545,N_1497,N_1447);
nand U1546 (N_1546,N_1481,N_1441);
and U1547 (N_1547,N_1488,N_1408);
and U1548 (N_1548,N_1458,N_1465);
or U1549 (N_1549,N_1462,N_1439);
or U1550 (N_1550,N_1417,N_1468);
nor U1551 (N_1551,N_1424,N_1463);
nor U1552 (N_1552,N_1419,N_1491);
or U1553 (N_1553,N_1484,N_1487);
nand U1554 (N_1554,N_1450,N_1491);
nor U1555 (N_1555,N_1455,N_1493);
nand U1556 (N_1556,N_1413,N_1477);
nand U1557 (N_1557,N_1479,N_1415);
or U1558 (N_1558,N_1422,N_1479);
or U1559 (N_1559,N_1444,N_1464);
nand U1560 (N_1560,N_1459,N_1409);
or U1561 (N_1561,N_1463,N_1445);
nor U1562 (N_1562,N_1409,N_1486);
or U1563 (N_1563,N_1476,N_1412);
or U1564 (N_1564,N_1466,N_1408);
or U1565 (N_1565,N_1422,N_1488);
or U1566 (N_1566,N_1484,N_1495);
xor U1567 (N_1567,N_1497,N_1465);
nand U1568 (N_1568,N_1460,N_1420);
nand U1569 (N_1569,N_1463,N_1480);
nand U1570 (N_1570,N_1425,N_1471);
or U1571 (N_1571,N_1476,N_1407);
nand U1572 (N_1572,N_1419,N_1438);
nand U1573 (N_1573,N_1486,N_1438);
nand U1574 (N_1574,N_1438,N_1417);
or U1575 (N_1575,N_1470,N_1454);
or U1576 (N_1576,N_1437,N_1481);
nor U1577 (N_1577,N_1493,N_1411);
and U1578 (N_1578,N_1473,N_1478);
nor U1579 (N_1579,N_1434,N_1498);
nor U1580 (N_1580,N_1495,N_1468);
or U1581 (N_1581,N_1436,N_1464);
or U1582 (N_1582,N_1445,N_1490);
nor U1583 (N_1583,N_1438,N_1458);
or U1584 (N_1584,N_1449,N_1417);
or U1585 (N_1585,N_1415,N_1449);
and U1586 (N_1586,N_1461,N_1457);
and U1587 (N_1587,N_1469,N_1464);
and U1588 (N_1588,N_1461,N_1468);
and U1589 (N_1589,N_1462,N_1451);
xnor U1590 (N_1590,N_1434,N_1412);
nor U1591 (N_1591,N_1408,N_1461);
nor U1592 (N_1592,N_1489,N_1423);
nor U1593 (N_1593,N_1417,N_1446);
or U1594 (N_1594,N_1443,N_1465);
or U1595 (N_1595,N_1465,N_1413);
or U1596 (N_1596,N_1453,N_1454);
nor U1597 (N_1597,N_1440,N_1433);
nor U1598 (N_1598,N_1400,N_1403);
nand U1599 (N_1599,N_1469,N_1429);
nor U1600 (N_1600,N_1547,N_1590);
nor U1601 (N_1601,N_1517,N_1548);
nand U1602 (N_1602,N_1542,N_1586);
nand U1603 (N_1603,N_1555,N_1593);
nand U1604 (N_1604,N_1516,N_1582);
and U1605 (N_1605,N_1502,N_1562);
or U1606 (N_1606,N_1507,N_1559);
nand U1607 (N_1607,N_1558,N_1587);
or U1608 (N_1608,N_1513,N_1510);
or U1609 (N_1609,N_1581,N_1579);
and U1610 (N_1610,N_1574,N_1566);
and U1611 (N_1611,N_1543,N_1525);
nand U1612 (N_1612,N_1594,N_1556);
or U1613 (N_1613,N_1541,N_1589);
nor U1614 (N_1614,N_1505,N_1526);
nand U1615 (N_1615,N_1568,N_1580);
or U1616 (N_1616,N_1503,N_1588);
nand U1617 (N_1617,N_1506,N_1557);
or U1618 (N_1618,N_1592,N_1528);
or U1619 (N_1619,N_1572,N_1561);
or U1620 (N_1620,N_1584,N_1514);
nand U1621 (N_1621,N_1535,N_1597);
nor U1622 (N_1622,N_1571,N_1583);
nor U1623 (N_1623,N_1504,N_1550);
and U1624 (N_1624,N_1520,N_1578);
nand U1625 (N_1625,N_1533,N_1538);
and U1626 (N_1626,N_1569,N_1595);
nor U1627 (N_1627,N_1570,N_1529);
or U1628 (N_1628,N_1524,N_1522);
nand U1629 (N_1629,N_1536,N_1501);
and U1630 (N_1630,N_1523,N_1527);
and U1631 (N_1631,N_1560,N_1515);
nand U1632 (N_1632,N_1540,N_1553);
nand U1633 (N_1633,N_1532,N_1554);
nor U1634 (N_1634,N_1549,N_1546);
and U1635 (N_1635,N_1509,N_1534);
and U1636 (N_1636,N_1565,N_1521);
or U1637 (N_1637,N_1596,N_1519);
or U1638 (N_1638,N_1531,N_1508);
or U1639 (N_1639,N_1544,N_1518);
or U1640 (N_1640,N_1512,N_1576);
nor U1641 (N_1641,N_1567,N_1545);
nor U1642 (N_1642,N_1598,N_1537);
nand U1643 (N_1643,N_1577,N_1500);
nand U1644 (N_1644,N_1591,N_1585);
or U1645 (N_1645,N_1573,N_1551);
or U1646 (N_1646,N_1530,N_1599);
or U1647 (N_1647,N_1511,N_1552);
nand U1648 (N_1648,N_1575,N_1564);
nand U1649 (N_1649,N_1563,N_1539);
nor U1650 (N_1650,N_1541,N_1510);
or U1651 (N_1651,N_1567,N_1580);
and U1652 (N_1652,N_1507,N_1519);
nand U1653 (N_1653,N_1532,N_1565);
or U1654 (N_1654,N_1549,N_1510);
and U1655 (N_1655,N_1523,N_1575);
and U1656 (N_1656,N_1560,N_1587);
and U1657 (N_1657,N_1521,N_1529);
nor U1658 (N_1658,N_1531,N_1579);
nor U1659 (N_1659,N_1513,N_1523);
nand U1660 (N_1660,N_1598,N_1542);
and U1661 (N_1661,N_1503,N_1560);
nor U1662 (N_1662,N_1551,N_1515);
and U1663 (N_1663,N_1530,N_1566);
nand U1664 (N_1664,N_1560,N_1553);
nand U1665 (N_1665,N_1543,N_1546);
and U1666 (N_1666,N_1561,N_1541);
nor U1667 (N_1667,N_1570,N_1542);
nand U1668 (N_1668,N_1552,N_1542);
nor U1669 (N_1669,N_1554,N_1542);
or U1670 (N_1670,N_1537,N_1576);
or U1671 (N_1671,N_1515,N_1502);
nor U1672 (N_1672,N_1599,N_1554);
nand U1673 (N_1673,N_1540,N_1572);
or U1674 (N_1674,N_1570,N_1597);
and U1675 (N_1675,N_1595,N_1578);
nor U1676 (N_1676,N_1517,N_1544);
or U1677 (N_1677,N_1518,N_1538);
nor U1678 (N_1678,N_1566,N_1547);
and U1679 (N_1679,N_1526,N_1569);
or U1680 (N_1680,N_1593,N_1562);
nor U1681 (N_1681,N_1564,N_1510);
nor U1682 (N_1682,N_1552,N_1599);
or U1683 (N_1683,N_1566,N_1536);
and U1684 (N_1684,N_1569,N_1522);
or U1685 (N_1685,N_1555,N_1575);
nor U1686 (N_1686,N_1573,N_1572);
or U1687 (N_1687,N_1577,N_1522);
and U1688 (N_1688,N_1530,N_1518);
and U1689 (N_1689,N_1561,N_1535);
nor U1690 (N_1690,N_1554,N_1566);
and U1691 (N_1691,N_1527,N_1559);
or U1692 (N_1692,N_1588,N_1582);
nor U1693 (N_1693,N_1505,N_1515);
nand U1694 (N_1694,N_1504,N_1591);
nor U1695 (N_1695,N_1580,N_1535);
nand U1696 (N_1696,N_1521,N_1593);
or U1697 (N_1697,N_1529,N_1576);
nor U1698 (N_1698,N_1531,N_1551);
and U1699 (N_1699,N_1518,N_1578);
and U1700 (N_1700,N_1600,N_1633);
and U1701 (N_1701,N_1624,N_1651);
and U1702 (N_1702,N_1611,N_1694);
and U1703 (N_1703,N_1654,N_1605);
or U1704 (N_1704,N_1658,N_1696);
and U1705 (N_1705,N_1681,N_1621);
and U1706 (N_1706,N_1648,N_1671);
nor U1707 (N_1707,N_1620,N_1609);
or U1708 (N_1708,N_1666,N_1629);
or U1709 (N_1709,N_1634,N_1606);
nand U1710 (N_1710,N_1673,N_1643);
nor U1711 (N_1711,N_1663,N_1684);
and U1712 (N_1712,N_1623,N_1695);
or U1713 (N_1713,N_1678,N_1653);
nor U1714 (N_1714,N_1677,N_1638);
and U1715 (N_1715,N_1693,N_1646);
nor U1716 (N_1716,N_1676,N_1698);
or U1717 (N_1717,N_1637,N_1647);
and U1718 (N_1718,N_1699,N_1618);
nor U1719 (N_1719,N_1692,N_1685);
nor U1720 (N_1720,N_1674,N_1639);
and U1721 (N_1721,N_1645,N_1625);
and U1722 (N_1722,N_1683,N_1660);
or U1723 (N_1723,N_1612,N_1622);
or U1724 (N_1724,N_1614,N_1601);
nor U1725 (N_1725,N_1630,N_1613);
nand U1726 (N_1726,N_1615,N_1616);
nand U1727 (N_1727,N_1655,N_1627);
or U1728 (N_1728,N_1662,N_1679);
xor U1729 (N_1729,N_1604,N_1670);
or U1730 (N_1730,N_1686,N_1602);
nor U1731 (N_1731,N_1665,N_1640);
or U1732 (N_1732,N_1691,N_1617);
nand U1733 (N_1733,N_1675,N_1659);
or U1734 (N_1734,N_1668,N_1644);
and U1735 (N_1735,N_1669,N_1631);
nor U1736 (N_1736,N_1687,N_1628);
nor U1737 (N_1737,N_1607,N_1619);
or U1738 (N_1738,N_1610,N_1635);
nand U1739 (N_1739,N_1652,N_1636);
or U1740 (N_1740,N_1672,N_1649);
nand U1741 (N_1741,N_1656,N_1664);
or U1742 (N_1742,N_1650,N_1608);
and U1743 (N_1743,N_1641,N_1680);
and U1744 (N_1744,N_1690,N_1642);
or U1745 (N_1745,N_1626,N_1661);
nor U1746 (N_1746,N_1667,N_1603);
nor U1747 (N_1747,N_1689,N_1688);
nor U1748 (N_1748,N_1697,N_1682);
nor U1749 (N_1749,N_1657,N_1632);
nor U1750 (N_1750,N_1646,N_1699);
and U1751 (N_1751,N_1699,N_1611);
nor U1752 (N_1752,N_1613,N_1607);
nor U1753 (N_1753,N_1674,N_1620);
or U1754 (N_1754,N_1654,N_1641);
nor U1755 (N_1755,N_1601,N_1684);
or U1756 (N_1756,N_1681,N_1643);
and U1757 (N_1757,N_1693,N_1606);
nor U1758 (N_1758,N_1662,N_1603);
xor U1759 (N_1759,N_1685,N_1649);
nand U1760 (N_1760,N_1647,N_1660);
nand U1761 (N_1761,N_1699,N_1633);
and U1762 (N_1762,N_1629,N_1607);
nor U1763 (N_1763,N_1672,N_1635);
nand U1764 (N_1764,N_1637,N_1656);
nor U1765 (N_1765,N_1674,N_1623);
nor U1766 (N_1766,N_1649,N_1642);
nor U1767 (N_1767,N_1643,N_1609);
or U1768 (N_1768,N_1662,N_1690);
nand U1769 (N_1769,N_1619,N_1601);
nand U1770 (N_1770,N_1658,N_1602);
and U1771 (N_1771,N_1621,N_1628);
nor U1772 (N_1772,N_1606,N_1639);
and U1773 (N_1773,N_1640,N_1664);
or U1774 (N_1774,N_1653,N_1673);
nand U1775 (N_1775,N_1625,N_1695);
nand U1776 (N_1776,N_1689,N_1657);
and U1777 (N_1777,N_1610,N_1609);
and U1778 (N_1778,N_1674,N_1610);
and U1779 (N_1779,N_1675,N_1676);
and U1780 (N_1780,N_1685,N_1609);
nor U1781 (N_1781,N_1697,N_1696);
nand U1782 (N_1782,N_1670,N_1641);
nand U1783 (N_1783,N_1635,N_1629);
nand U1784 (N_1784,N_1657,N_1651);
and U1785 (N_1785,N_1601,N_1602);
or U1786 (N_1786,N_1688,N_1608);
nor U1787 (N_1787,N_1650,N_1610);
nand U1788 (N_1788,N_1620,N_1652);
nor U1789 (N_1789,N_1674,N_1677);
nor U1790 (N_1790,N_1660,N_1651);
nor U1791 (N_1791,N_1625,N_1666);
nand U1792 (N_1792,N_1685,N_1668);
nor U1793 (N_1793,N_1629,N_1656);
nand U1794 (N_1794,N_1695,N_1674);
or U1795 (N_1795,N_1690,N_1650);
nor U1796 (N_1796,N_1620,N_1605);
or U1797 (N_1797,N_1686,N_1681);
and U1798 (N_1798,N_1663,N_1607);
nand U1799 (N_1799,N_1634,N_1620);
nor U1800 (N_1800,N_1709,N_1785);
nand U1801 (N_1801,N_1799,N_1745);
nor U1802 (N_1802,N_1798,N_1716);
nand U1803 (N_1803,N_1703,N_1790);
and U1804 (N_1804,N_1765,N_1764);
nand U1805 (N_1805,N_1786,N_1737);
nand U1806 (N_1806,N_1705,N_1754);
nand U1807 (N_1807,N_1721,N_1746);
nand U1808 (N_1808,N_1796,N_1775);
nor U1809 (N_1809,N_1701,N_1713);
and U1810 (N_1810,N_1782,N_1741);
nand U1811 (N_1811,N_1788,N_1760);
or U1812 (N_1812,N_1763,N_1733);
and U1813 (N_1813,N_1724,N_1718);
nor U1814 (N_1814,N_1723,N_1762);
and U1815 (N_1815,N_1759,N_1726);
nor U1816 (N_1816,N_1711,N_1780);
nor U1817 (N_1817,N_1797,N_1784);
nor U1818 (N_1818,N_1751,N_1758);
and U1819 (N_1819,N_1715,N_1767);
nor U1820 (N_1820,N_1712,N_1710);
or U1821 (N_1821,N_1795,N_1734);
nor U1822 (N_1822,N_1757,N_1719);
nand U1823 (N_1823,N_1750,N_1781);
and U1824 (N_1824,N_1727,N_1739);
nand U1825 (N_1825,N_1779,N_1720);
nand U1826 (N_1826,N_1771,N_1728);
nand U1827 (N_1827,N_1704,N_1770);
and U1828 (N_1828,N_1768,N_1747);
nand U1829 (N_1829,N_1735,N_1702);
nor U1830 (N_1830,N_1783,N_1725);
nor U1831 (N_1831,N_1700,N_1749);
and U1832 (N_1832,N_1787,N_1740);
or U1833 (N_1833,N_1766,N_1732);
or U1834 (N_1834,N_1778,N_1714);
nor U1835 (N_1835,N_1777,N_1769);
and U1836 (N_1836,N_1772,N_1792);
or U1837 (N_1837,N_1791,N_1789);
and U1838 (N_1838,N_1722,N_1729);
nand U1839 (N_1839,N_1793,N_1743);
and U1840 (N_1840,N_1706,N_1717);
nor U1841 (N_1841,N_1736,N_1707);
nand U1842 (N_1842,N_1731,N_1755);
and U1843 (N_1843,N_1753,N_1761);
nor U1844 (N_1844,N_1794,N_1752);
and U1845 (N_1845,N_1774,N_1730);
and U1846 (N_1846,N_1744,N_1756);
and U1847 (N_1847,N_1748,N_1773);
nand U1848 (N_1848,N_1742,N_1776);
or U1849 (N_1849,N_1738,N_1708);
or U1850 (N_1850,N_1734,N_1714);
or U1851 (N_1851,N_1783,N_1734);
and U1852 (N_1852,N_1729,N_1788);
or U1853 (N_1853,N_1799,N_1739);
and U1854 (N_1854,N_1711,N_1778);
and U1855 (N_1855,N_1719,N_1787);
or U1856 (N_1856,N_1701,N_1796);
nor U1857 (N_1857,N_1791,N_1782);
nand U1858 (N_1858,N_1767,N_1793);
nand U1859 (N_1859,N_1717,N_1703);
and U1860 (N_1860,N_1770,N_1786);
or U1861 (N_1861,N_1753,N_1749);
and U1862 (N_1862,N_1712,N_1790);
nor U1863 (N_1863,N_1711,N_1745);
nor U1864 (N_1864,N_1721,N_1745);
nor U1865 (N_1865,N_1746,N_1701);
and U1866 (N_1866,N_1715,N_1701);
or U1867 (N_1867,N_1748,N_1747);
or U1868 (N_1868,N_1710,N_1713);
or U1869 (N_1869,N_1739,N_1740);
nand U1870 (N_1870,N_1745,N_1747);
nor U1871 (N_1871,N_1741,N_1717);
and U1872 (N_1872,N_1709,N_1758);
xor U1873 (N_1873,N_1738,N_1736);
or U1874 (N_1874,N_1748,N_1771);
nor U1875 (N_1875,N_1720,N_1789);
nand U1876 (N_1876,N_1735,N_1749);
nor U1877 (N_1877,N_1751,N_1786);
nand U1878 (N_1878,N_1756,N_1798);
nor U1879 (N_1879,N_1727,N_1758);
and U1880 (N_1880,N_1725,N_1780);
nor U1881 (N_1881,N_1744,N_1777);
or U1882 (N_1882,N_1770,N_1707);
nor U1883 (N_1883,N_1719,N_1756);
and U1884 (N_1884,N_1718,N_1786);
and U1885 (N_1885,N_1713,N_1704);
and U1886 (N_1886,N_1722,N_1713);
nor U1887 (N_1887,N_1788,N_1742);
or U1888 (N_1888,N_1732,N_1721);
nor U1889 (N_1889,N_1730,N_1719);
or U1890 (N_1890,N_1713,N_1765);
nand U1891 (N_1891,N_1734,N_1779);
or U1892 (N_1892,N_1734,N_1750);
nand U1893 (N_1893,N_1714,N_1773);
nor U1894 (N_1894,N_1785,N_1739);
nand U1895 (N_1895,N_1753,N_1779);
and U1896 (N_1896,N_1713,N_1769);
nand U1897 (N_1897,N_1755,N_1781);
nor U1898 (N_1898,N_1765,N_1777);
and U1899 (N_1899,N_1793,N_1701);
nor U1900 (N_1900,N_1808,N_1822);
nor U1901 (N_1901,N_1801,N_1864);
nor U1902 (N_1902,N_1831,N_1840);
nand U1903 (N_1903,N_1860,N_1890);
nand U1904 (N_1904,N_1862,N_1867);
nand U1905 (N_1905,N_1881,N_1811);
and U1906 (N_1906,N_1813,N_1879);
nand U1907 (N_1907,N_1882,N_1810);
nor U1908 (N_1908,N_1854,N_1869);
and U1909 (N_1909,N_1868,N_1844);
or U1910 (N_1910,N_1877,N_1828);
or U1911 (N_1911,N_1898,N_1875);
or U1912 (N_1912,N_1836,N_1852);
nor U1913 (N_1913,N_1816,N_1825);
or U1914 (N_1914,N_1821,N_1865);
nor U1915 (N_1915,N_1835,N_1846);
and U1916 (N_1916,N_1870,N_1829);
and U1917 (N_1917,N_1804,N_1885);
and U1918 (N_1918,N_1830,N_1842);
nand U1919 (N_1919,N_1800,N_1814);
and U1920 (N_1920,N_1807,N_1851);
or U1921 (N_1921,N_1809,N_1883);
and U1922 (N_1922,N_1863,N_1850);
or U1923 (N_1923,N_1833,N_1826);
nor U1924 (N_1924,N_1861,N_1892);
nor U1925 (N_1925,N_1812,N_1848);
nor U1926 (N_1926,N_1872,N_1876);
nor U1927 (N_1927,N_1843,N_1891);
nor U1928 (N_1928,N_1858,N_1847);
nor U1929 (N_1929,N_1815,N_1806);
nor U1930 (N_1930,N_1837,N_1874);
nor U1931 (N_1931,N_1827,N_1859);
nand U1932 (N_1932,N_1887,N_1873);
and U1933 (N_1933,N_1895,N_1805);
and U1934 (N_1934,N_1838,N_1839);
nor U1935 (N_1935,N_1820,N_1878);
and U1936 (N_1936,N_1853,N_1889);
or U1937 (N_1937,N_1803,N_1888);
and U1938 (N_1938,N_1817,N_1849);
nor U1939 (N_1939,N_1823,N_1857);
and U1940 (N_1940,N_1818,N_1880);
nand U1941 (N_1941,N_1886,N_1841);
nand U1942 (N_1942,N_1855,N_1884);
nand U1943 (N_1943,N_1897,N_1856);
nand U1944 (N_1944,N_1899,N_1819);
or U1945 (N_1945,N_1802,N_1834);
nand U1946 (N_1946,N_1824,N_1894);
and U1947 (N_1947,N_1896,N_1866);
or U1948 (N_1948,N_1893,N_1832);
or U1949 (N_1949,N_1845,N_1871);
nor U1950 (N_1950,N_1878,N_1829);
xnor U1951 (N_1951,N_1827,N_1893);
and U1952 (N_1952,N_1865,N_1800);
or U1953 (N_1953,N_1819,N_1884);
and U1954 (N_1954,N_1812,N_1832);
nand U1955 (N_1955,N_1804,N_1833);
nand U1956 (N_1956,N_1884,N_1811);
or U1957 (N_1957,N_1882,N_1808);
or U1958 (N_1958,N_1888,N_1821);
and U1959 (N_1959,N_1823,N_1826);
nand U1960 (N_1960,N_1858,N_1824);
nand U1961 (N_1961,N_1852,N_1855);
nand U1962 (N_1962,N_1897,N_1842);
or U1963 (N_1963,N_1897,N_1850);
or U1964 (N_1964,N_1879,N_1848);
nand U1965 (N_1965,N_1869,N_1885);
and U1966 (N_1966,N_1863,N_1877);
or U1967 (N_1967,N_1850,N_1871);
or U1968 (N_1968,N_1881,N_1829);
and U1969 (N_1969,N_1859,N_1872);
nand U1970 (N_1970,N_1844,N_1832);
and U1971 (N_1971,N_1868,N_1884);
nand U1972 (N_1972,N_1886,N_1801);
or U1973 (N_1973,N_1868,N_1801);
nand U1974 (N_1974,N_1810,N_1871);
nor U1975 (N_1975,N_1884,N_1842);
nand U1976 (N_1976,N_1899,N_1882);
and U1977 (N_1977,N_1850,N_1831);
nand U1978 (N_1978,N_1808,N_1855);
and U1979 (N_1979,N_1825,N_1855);
nor U1980 (N_1980,N_1815,N_1888);
nor U1981 (N_1981,N_1887,N_1843);
or U1982 (N_1982,N_1847,N_1866);
and U1983 (N_1983,N_1882,N_1826);
and U1984 (N_1984,N_1849,N_1857);
and U1985 (N_1985,N_1802,N_1879);
nor U1986 (N_1986,N_1850,N_1836);
nand U1987 (N_1987,N_1801,N_1856);
or U1988 (N_1988,N_1821,N_1889);
nand U1989 (N_1989,N_1889,N_1870);
and U1990 (N_1990,N_1800,N_1823);
nor U1991 (N_1991,N_1882,N_1864);
and U1992 (N_1992,N_1825,N_1823);
nand U1993 (N_1993,N_1848,N_1857);
nand U1994 (N_1994,N_1830,N_1873);
and U1995 (N_1995,N_1860,N_1867);
nor U1996 (N_1996,N_1812,N_1874);
and U1997 (N_1997,N_1895,N_1825);
or U1998 (N_1998,N_1859,N_1884);
nand U1999 (N_1999,N_1863,N_1856);
nor U2000 (N_2000,N_1953,N_1929);
or U2001 (N_2001,N_1951,N_1932);
xor U2002 (N_2002,N_1908,N_1981);
nor U2003 (N_2003,N_1962,N_1945);
or U2004 (N_2004,N_1907,N_1974);
nor U2005 (N_2005,N_1920,N_1931);
or U2006 (N_2006,N_1933,N_1971);
or U2007 (N_2007,N_1988,N_1991);
nor U2008 (N_2008,N_1949,N_1977);
nand U2009 (N_2009,N_1930,N_1995);
nor U2010 (N_2010,N_1984,N_1987);
nor U2011 (N_2011,N_1943,N_1902);
nand U2012 (N_2012,N_1969,N_1927);
nand U2013 (N_2013,N_1964,N_1967);
and U2014 (N_2014,N_1989,N_1922);
xnor U2015 (N_2015,N_1923,N_1968);
and U2016 (N_2016,N_1982,N_1924);
and U2017 (N_2017,N_1985,N_1959);
nor U2018 (N_2018,N_1990,N_1935);
nand U2019 (N_2019,N_1910,N_1939);
nand U2020 (N_2020,N_1948,N_1954);
and U2021 (N_2021,N_1998,N_1992);
nor U2022 (N_2022,N_1938,N_1913);
and U2023 (N_2023,N_1950,N_1905);
nor U2024 (N_2024,N_1958,N_1996);
and U2025 (N_2025,N_1957,N_1956);
or U2026 (N_2026,N_1946,N_1952);
nand U2027 (N_2027,N_1941,N_1961);
and U2028 (N_2028,N_1942,N_1936);
nor U2029 (N_2029,N_1921,N_1973);
nor U2030 (N_2030,N_1997,N_1978);
and U2031 (N_2031,N_1970,N_1955);
nand U2032 (N_2032,N_1906,N_1917);
and U2033 (N_2033,N_1944,N_1914);
and U2034 (N_2034,N_1918,N_1966);
nand U2035 (N_2035,N_1915,N_1940);
and U2036 (N_2036,N_1916,N_1993);
or U2037 (N_2037,N_1980,N_1909);
nor U2038 (N_2038,N_1928,N_1963);
and U2039 (N_2039,N_1972,N_1937);
or U2040 (N_2040,N_1901,N_1999);
or U2041 (N_2041,N_1986,N_1979);
xnor U2042 (N_2042,N_1983,N_1934);
or U2043 (N_2043,N_1994,N_1975);
or U2044 (N_2044,N_1926,N_1976);
nor U2045 (N_2045,N_1903,N_1904);
and U2046 (N_2046,N_1912,N_1900);
xnor U2047 (N_2047,N_1919,N_1947);
nand U2048 (N_2048,N_1960,N_1911);
or U2049 (N_2049,N_1925,N_1965);
and U2050 (N_2050,N_1921,N_1938);
nand U2051 (N_2051,N_1982,N_1920);
xnor U2052 (N_2052,N_1935,N_1955);
and U2053 (N_2053,N_1985,N_1978);
nand U2054 (N_2054,N_1948,N_1999);
nor U2055 (N_2055,N_1953,N_1912);
nand U2056 (N_2056,N_1956,N_1997);
nor U2057 (N_2057,N_1916,N_1939);
or U2058 (N_2058,N_1934,N_1907);
and U2059 (N_2059,N_1906,N_1999);
nor U2060 (N_2060,N_1935,N_1976);
and U2061 (N_2061,N_1982,N_1938);
and U2062 (N_2062,N_1987,N_1988);
or U2063 (N_2063,N_1962,N_1966);
or U2064 (N_2064,N_1938,N_1951);
or U2065 (N_2065,N_1937,N_1909);
and U2066 (N_2066,N_1973,N_1951);
xnor U2067 (N_2067,N_1961,N_1927);
nor U2068 (N_2068,N_1929,N_1967);
and U2069 (N_2069,N_1981,N_1958);
or U2070 (N_2070,N_1954,N_1952);
or U2071 (N_2071,N_1998,N_1938);
and U2072 (N_2072,N_1922,N_1936);
and U2073 (N_2073,N_1945,N_1915);
nand U2074 (N_2074,N_1908,N_1993);
nand U2075 (N_2075,N_1905,N_1922);
nor U2076 (N_2076,N_1951,N_1925);
and U2077 (N_2077,N_1958,N_1940);
and U2078 (N_2078,N_1980,N_1944);
and U2079 (N_2079,N_1935,N_1989);
or U2080 (N_2080,N_1983,N_1939);
or U2081 (N_2081,N_1956,N_1925);
and U2082 (N_2082,N_1973,N_1923);
or U2083 (N_2083,N_1947,N_1904);
and U2084 (N_2084,N_1946,N_1983);
nand U2085 (N_2085,N_1932,N_1966);
and U2086 (N_2086,N_1914,N_1961);
or U2087 (N_2087,N_1936,N_1910);
and U2088 (N_2088,N_1973,N_1999);
or U2089 (N_2089,N_1922,N_1951);
or U2090 (N_2090,N_1938,N_1986);
nand U2091 (N_2091,N_1946,N_1951);
nand U2092 (N_2092,N_1906,N_1934);
nor U2093 (N_2093,N_1979,N_1936);
or U2094 (N_2094,N_1917,N_1980);
nand U2095 (N_2095,N_1985,N_1934);
and U2096 (N_2096,N_1918,N_1983);
or U2097 (N_2097,N_1904,N_1918);
nand U2098 (N_2098,N_1988,N_1901);
and U2099 (N_2099,N_1986,N_1927);
nand U2100 (N_2100,N_2096,N_2075);
and U2101 (N_2101,N_2034,N_2081);
or U2102 (N_2102,N_2077,N_2062);
nand U2103 (N_2103,N_2095,N_2045);
nor U2104 (N_2104,N_2080,N_2059);
nor U2105 (N_2105,N_2052,N_2082);
and U2106 (N_2106,N_2030,N_2067);
or U2107 (N_2107,N_2025,N_2056);
and U2108 (N_2108,N_2029,N_2069);
xor U2109 (N_2109,N_2003,N_2011);
nand U2110 (N_2110,N_2055,N_2074);
nand U2111 (N_2111,N_2057,N_2016);
nor U2112 (N_2112,N_2061,N_2068);
nor U2113 (N_2113,N_2024,N_2043);
or U2114 (N_2114,N_2021,N_2065);
or U2115 (N_2115,N_2054,N_2039);
or U2116 (N_2116,N_2000,N_2088);
nand U2117 (N_2117,N_2058,N_2037);
nor U2118 (N_2118,N_2071,N_2026);
nor U2119 (N_2119,N_2006,N_2084);
and U2120 (N_2120,N_2091,N_2064);
nor U2121 (N_2121,N_2083,N_2040);
or U2122 (N_2122,N_2020,N_2099);
or U2123 (N_2123,N_2035,N_2093);
nor U2124 (N_2124,N_2009,N_2060);
nor U2125 (N_2125,N_2027,N_2038);
nor U2126 (N_2126,N_2094,N_2090);
nand U2127 (N_2127,N_2007,N_2018);
nor U2128 (N_2128,N_2085,N_2036);
nor U2129 (N_2129,N_2023,N_2028);
or U2130 (N_2130,N_2049,N_2041);
nand U2131 (N_2131,N_2010,N_2070);
or U2132 (N_2132,N_2087,N_2089);
nand U2133 (N_2133,N_2013,N_2063);
or U2134 (N_2134,N_2004,N_2053);
nand U2135 (N_2135,N_2079,N_2044);
or U2136 (N_2136,N_2019,N_2002);
and U2137 (N_2137,N_2050,N_2042);
nor U2138 (N_2138,N_2046,N_2098);
nand U2139 (N_2139,N_2073,N_2031);
or U2140 (N_2140,N_2015,N_2008);
or U2141 (N_2141,N_2086,N_2066);
and U2142 (N_2142,N_2022,N_2092);
nand U2143 (N_2143,N_2012,N_2076);
nand U2144 (N_2144,N_2017,N_2033);
or U2145 (N_2145,N_2005,N_2078);
nand U2146 (N_2146,N_2014,N_2001);
and U2147 (N_2147,N_2047,N_2072);
nand U2148 (N_2148,N_2097,N_2051);
nand U2149 (N_2149,N_2048,N_2032);
nand U2150 (N_2150,N_2062,N_2040);
and U2151 (N_2151,N_2064,N_2059);
and U2152 (N_2152,N_2041,N_2012);
and U2153 (N_2153,N_2057,N_2084);
and U2154 (N_2154,N_2035,N_2080);
nand U2155 (N_2155,N_2006,N_2001);
or U2156 (N_2156,N_2075,N_2031);
nand U2157 (N_2157,N_2014,N_2099);
and U2158 (N_2158,N_2004,N_2090);
nor U2159 (N_2159,N_2095,N_2005);
nand U2160 (N_2160,N_2047,N_2071);
and U2161 (N_2161,N_2037,N_2008);
nand U2162 (N_2162,N_2092,N_2037);
and U2163 (N_2163,N_2044,N_2083);
nand U2164 (N_2164,N_2084,N_2095);
nand U2165 (N_2165,N_2075,N_2072);
nand U2166 (N_2166,N_2052,N_2080);
nor U2167 (N_2167,N_2088,N_2050);
and U2168 (N_2168,N_2077,N_2001);
or U2169 (N_2169,N_2050,N_2057);
and U2170 (N_2170,N_2094,N_2031);
nor U2171 (N_2171,N_2048,N_2003);
nand U2172 (N_2172,N_2038,N_2036);
or U2173 (N_2173,N_2018,N_2025);
nor U2174 (N_2174,N_2063,N_2002);
or U2175 (N_2175,N_2043,N_2004);
nand U2176 (N_2176,N_2072,N_2041);
nor U2177 (N_2177,N_2010,N_2002);
or U2178 (N_2178,N_2094,N_2037);
nor U2179 (N_2179,N_2065,N_2003);
nand U2180 (N_2180,N_2011,N_2054);
or U2181 (N_2181,N_2074,N_2073);
or U2182 (N_2182,N_2090,N_2070);
and U2183 (N_2183,N_2026,N_2017);
or U2184 (N_2184,N_2074,N_2063);
nor U2185 (N_2185,N_2097,N_2070);
or U2186 (N_2186,N_2074,N_2087);
or U2187 (N_2187,N_2006,N_2016);
nand U2188 (N_2188,N_2066,N_2036);
and U2189 (N_2189,N_2006,N_2072);
and U2190 (N_2190,N_2055,N_2051);
or U2191 (N_2191,N_2057,N_2069);
nand U2192 (N_2192,N_2053,N_2010);
or U2193 (N_2193,N_2068,N_2028);
nand U2194 (N_2194,N_2089,N_2034);
and U2195 (N_2195,N_2099,N_2004);
or U2196 (N_2196,N_2086,N_2060);
and U2197 (N_2197,N_2023,N_2063);
nand U2198 (N_2198,N_2056,N_2061);
or U2199 (N_2199,N_2014,N_2095);
or U2200 (N_2200,N_2106,N_2135);
nand U2201 (N_2201,N_2115,N_2114);
or U2202 (N_2202,N_2157,N_2193);
and U2203 (N_2203,N_2181,N_2107);
nor U2204 (N_2204,N_2171,N_2197);
nand U2205 (N_2205,N_2190,N_2155);
nand U2206 (N_2206,N_2180,N_2188);
or U2207 (N_2207,N_2102,N_2101);
or U2208 (N_2208,N_2141,N_2196);
nand U2209 (N_2209,N_2116,N_2187);
nand U2210 (N_2210,N_2129,N_2140);
xnor U2211 (N_2211,N_2185,N_2151);
or U2212 (N_2212,N_2112,N_2110);
nor U2213 (N_2213,N_2169,N_2182);
or U2214 (N_2214,N_2119,N_2111);
and U2215 (N_2215,N_2184,N_2125);
nand U2216 (N_2216,N_2154,N_2124);
nor U2217 (N_2217,N_2108,N_2145);
and U2218 (N_2218,N_2192,N_2132);
and U2219 (N_2219,N_2130,N_2126);
nor U2220 (N_2220,N_2118,N_2136);
or U2221 (N_2221,N_2173,N_2161);
nand U2222 (N_2222,N_2104,N_2142);
or U2223 (N_2223,N_2189,N_2167);
or U2224 (N_2224,N_2177,N_2150);
or U2225 (N_2225,N_2137,N_2121);
nor U2226 (N_2226,N_2195,N_2143);
and U2227 (N_2227,N_2191,N_2186);
nor U2228 (N_2228,N_2146,N_2127);
and U2229 (N_2229,N_2144,N_2179);
nor U2230 (N_2230,N_2138,N_2170);
nand U2231 (N_2231,N_2123,N_2149);
or U2232 (N_2232,N_2164,N_2128);
nor U2233 (N_2233,N_2139,N_2183);
and U2234 (N_2234,N_2120,N_2168);
or U2235 (N_2235,N_2194,N_2117);
xor U2236 (N_2236,N_2198,N_2147);
nand U2237 (N_2237,N_2176,N_2159);
or U2238 (N_2238,N_2178,N_2100);
and U2239 (N_2239,N_2172,N_2153);
and U2240 (N_2240,N_2122,N_2160);
or U2241 (N_2241,N_2148,N_2152);
nand U2242 (N_2242,N_2134,N_2162);
nand U2243 (N_2243,N_2156,N_2158);
or U2244 (N_2244,N_2165,N_2166);
and U2245 (N_2245,N_2163,N_2199);
or U2246 (N_2246,N_2109,N_2175);
and U2247 (N_2247,N_2103,N_2131);
nor U2248 (N_2248,N_2174,N_2105);
nor U2249 (N_2249,N_2133,N_2113);
or U2250 (N_2250,N_2103,N_2155);
or U2251 (N_2251,N_2191,N_2194);
nor U2252 (N_2252,N_2157,N_2180);
nand U2253 (N_2253,N_2184,N_2185);
and U2254 (N_2254,N_2190,N_2164);
nand U2255 (N_2255,N_2174,N_2155);
nor U2256 (N_2256,N_2134,N_2191);
nand U2257 (N_2257,N_2149,N_2115);
and U2258 (N_2258,N_2176,N_2101);
or U2259 (N_2259,N_2168,N_2196);
or U2260 (N_2260,N_2192,N_2197);
nand U2261 (N_2261,N_2192,N_2191);
and U2262 (N_2262,N_2184,N_2193);
nor U2263 (N_2263,N_2119,N_2181);
or U2264 (N_2264,N_2183,N_2117);
and U2265 (N_2265,N_2136,N_2115);
or U2266 (N_2266,N_2165,N_2106);
and U2267 (N_2267,N_2110,N_2109);
nand U2268 (N_2268,N_2113,N_2140);
and U2269 (N_2269,N_2184,N_2100);
xor U2270 (N_2270,N_2110,N_2125);
nor U2271 (N_2271,N_2197,N_2190);
nand U2272 (N_2272,N_2149,N_2192);
nor U2273 (N_2273,N_2164,N_2196);
nor U2274 (N_2274,N_2118,N_2166);
nand U2275 (N_2275,N_2195,N_2198);
and U2276 (N_2276,N_2132,N_2175);
and U2277 (N_2277,N_2126,N_2195);
nand U2278 (N_2278,N_2162,N_2125);
nand U2279 (N_2279,N_2128,N_2177);
nand U2280 (N_2280,N_2157,N_2145);
nand U2281 (N_2281,N_2179,N_2115);
or U2282 (N_2282,N_2183,N_2147);
nor U2283 (N_2283,N_2196,N_2119);
nor U2284 (N_2284,N_2123,N_2158);
nand U2285 (N_2285,N_2152,N_2188);
nand U2286 (N_2286,N_2122,N_2110);
nor U2287 (N_2287,N_2120,N_2129);
nand U2288 (N_2288,N_2182,N_2104);
and U2289 (N_2289,N_2100,N_2107);
nor U2290 (N_2290,N_2193,N_2135);
nand U2291 (N_2291,N_2180,N_2168);
nor U2292 (N_2292,N_2138,N_2112);
or U2293 (N_2293,N_2145,N_2134);
nor U2294 (N_2294,N_2124,N_2121);
nand U2295 (N_2295,N_2173,N_2185);
nor U2296 (N_2296,N_2195,N_2122);
and U2297 (N_2297,N_2177,N_2155);
nand U2298 (N_2298,N_2149,N_2145);
nor U2299 (N_2299,N_2197,N_2172);
and U2300 (N_2300,N_2297,N_2253);
and U2301 (N_2301,N_2243,N_2231);
nand U2302 (N_2302,N_2286,N_2293);
or U2303 (N_2303,N_2210,N_2289);
nand U2304 (N_2304,N_2240,N_2205);
nand U2305 (N_2305,N_2221,N_2279);
nor U2306 (N_2306,N_2299,N_2298);
or U2307 (N_2307,N_2201,N_2238);
nor U2308 (N_2308,N_2282,N_2208);
nand U2309 (N_2309,N_2245,N_2285);
nor U2310 (N_2310,N_2236,N_2291);
and U2311 (N_2311,N_2233,N_2249);
or U2312 (N_2312,N_2264,N_2232);
and U2313 (N_2313,N_2220,N_2287);
nand U2314 (N_2314,N_2214,N_2206);
nor U2315 (N_2315,N_2218,N_2260);
and U2316 (N_2316,N_2266,N_2251);
nor U2317 (N_2317,N_2246,N_2235);
nor U2318 (N_2318,N_2250,N_2257);
or U2319 (N_2319,N_2252,N_2224);
or U2320 (N_2320,N_2215,N_2269);
and U2321 (N_2321,N_2277,N_2226);
nor U2322 (N_2322,N_2222,N_2268);
and U2323 (N_2323,N_2278,N_2284);
nand U2324 (N_2324,N_2242,N_2207);
or U2325 (N_2325,N_2209,N_2273);
nor U2326 (N_2326,N_2203,N_2234);
nor U2327 (N_2327,N_2256,N_2272);
and U2328 (N_2328,N_2288,N_2241);
or U2329 (N_2329,N_2254,N_2270);
and U2330 (N_2330,N_2259,N_2216);
or U2331 (N_2331,N_2227,N_2280);
nor U2332 (N_2332,N_2290,N_2219);
or U2333 (N_2333,N_2261,N_2223);
nand U2334 (N_2334,N_2239,N_2200);
nor U2335 (N_2335,N_2244,N_2211);
nor U2336 (N_2336,N_2265,N_2274);
or U2337 (N_2337,N_2255,N_2295);
or U2338 (N_2338,N_2212,N_2258);
and U2339 (N_2339,N_2248,N_2247);
and U2340 (N_2340,N_2275,N_2271);
nand U2341 (N_2341,N_2225,N_2276);
or U2342 (N_2342,N_2267,N_2230);
nand U2343 (N_2343,N_2292,N_2204);
nor U2344 (N_2344,N_2213,N_2237);
or U2345 (N_2345,N_2283,N_2202);
and U2346 (N_2346,N_2296,N_2281);
nand U2347 (N_2347,N_2229,N_2263);
nand U2348 (N_2348,N_2294,N_2228);
and U2349 (N_2349,N_2217,N_2262);
or U2350 (N_2350,N_2258,N_2228);
nand U2351 (N_2351,N_2263,N_2217);
or U2352 (N_2352,N_2240,N_2278);
nor U2353 (N_2353,N_2223,N_2285);
and U2354 (N_2354,N_2255,N_2247);
nand U2355 (N_2355,N_2213,N_2214);
or U2356 (N_2356,N_2272,N_2200);
or U2357 (N_2357,N_2237,N_2296);
or U2358 (N_2358,N_2201,N_2292);
nand U2359 (N_2359,N_2292,N_2202);
and U2360 (N_2360,N_2299,N_2243);
nor U2361 (N_2361,N_2222,N_2225);
nor U2362 (N_2362,N_2276,N_2200);
nand U2363 (N_2363,N_2249,N_2242);
nand U2364 (N_2364,N_2211,N_2214);
or U2365 (N_2365,N_2207,N_2290);
nand U2366 (N_2366,N_2207,N_2278);
nor U2367 (N_2367,N_2277,N_2289);
nor U2368 (N_2368,N_2259,N_2290);
and U2369 (N_2369,N_2262,N_2264);
and U2370 (N_2370,N_2284,N_2250);
or U2371 (N_2371,N_2260,N_2228);
nand U2372 (N_2372,N_2281,N_2282);
nand U2373 (N_2373,N_2235,N_2236);
or U2374 (N_2374,N_2231,N_2210);
and U2375 (N_2375,N_2286,N_2204);
nor U2376 (N_2376,N_2249,N_2275);
or U2377 (N_2377,N_2235,N_2273);
nand U2378 (N_2378,N_2298,N_2237);
and U2379 (N_2379,N_2229,N_2205);
nand U2380 (N_2380,N_2218,N_2281);
nand U2381 (N_2381,N_2223,N_2204);
and U2382 (N_2382,N_2244,N_2263);
nor U2383 (N_2383,N_2287,N_2280);
nor U2384 (N_2384,N_2292,N_2275);
nor U2385 (N_2385,N_2242,N_2247);
nor U2386 (N_2386,N_2276,N_2233);
xor U2387 (N_2387,N_2297,N_2272);
and U2388 (N_2388,N_2230,N_2296);
nand U2389 (N_2389,N_2208,N_2224);
nand U2390 (N_2390,N_2244,N_2200);
xnor U2391 (N_2391,N_2236,N_2255);
or U2392 (N_2392,N_2226,N_2286);
nor U2393 (N_2393,N_2267,N_2282);
nand U2394 (N_2394,N_2237,N_2209);
or U2395 (N_2395,N_2259,N_2236);
or U2396 (N_2396,N_2237,N_2212);
and U2397 (N_2397,N_2204,N_2224);
or U2398 (N_2398,N_2298,N_2258);
or U2399 (N_2399,N_2272,N_2281);
nor U2400 (N_2400,N_2369,N_2323);
nor U2401 (N_2401,N_2336,N_2322);
or U2402 (N_2402,N_2366,N_2381);
nand U2403 (N_2403,N_2302,N_2378);
or U2404 (N_2404,N_2309,N_2346);
or U2405 (N_2405,N_2389,N_2396);
nor U2406 (N_2406,N_2351,N_2317);
nand U2407 (N_2407,N_2305,N_2363);
and U2408 (N_2408,N_2388,N_2315);
nor U2409 (N_2409,N_2313,N_2367);
and U2410 (N_2410,N_2370,N_2326);
nand U2411 (N_2411,N_2379,N_2365);
or U2412 (N_2412,N_2373,N_2318);
nand U2413 (N_2413,N_2382,N_2301);
and U2414 (N_2414,N_2356,N_2359);
or U2415 (N_2415,N_2348,N_2394);
and U2416 (N_2416,N_2368,N_2357);
and U2417 (N_2417,N_2387,N_2306);
or U2418 (N_2418,N_2339,N_2333);
nand U2419 (N_2419,N_2300,N_2371);
nor U2420 (N_2420,N_2385,N_2353);
nor U2421 (N_2421,N_2324,N_2304);
or U2422 (N_2422,N_2358,N_2399);
or U2423 (N_2423,N_2349,N_2344);
nand U2424 (N_2424,N_2319,N_2320);
nor U2425 (N_2425,N_2390,N_2310);
nand U2426 (N_2426,N_2391,N_2395);
and U2427 (N_2427,N_2337,N_2354);
nand U2428 (N_2428,N_2311,N_2338);
nand U2429 (N_2429,N_2355,N_2364);
nand U2430 (N_2430,N_2376,N_2308);
nand U2431 (N_2431,N_2345,N_2372);
and U2432 (N_2432,N_2386,N_2380);
or U2433 (N_2433,N_2361,N_2314);
and U2434 (N_2434,N_2343,N_2327);
nor U2435 (N_2435,N_2321,N_2312);
nand U2436 (N_2436,N_2398,N_2397);
nand U2437 (N_2437,N_2350,N_2316);
nor U2438 (N_2438,N_2375,N_2342);
and U2439 (N_2439,N_2383,N_2374);
nor U2440 (N_2440,N_2335,N_2303);
nand U2441 (N_2441,N_2332,N_2331);
nand U2442 (N_2442,N_2377,N_2328);
nor U2443 (N_2443,N_2334,N_2330);
nor U2444 (N_2444,N_2307,N_2362);
and U2445 (N_2445,N_2325,N_2340);
or U2446 (N_2446,N_2392,N_2352);
nand U2447 (N_2447,N_2384,N_2360);
or U2448 (N_2448,N_2393,N_2329);
nand U2449 (N_2449,N_2347,N_2341);
or U2450 (N_2450,N_2302,N_2313);
and U2451 (N_2451,N_2369,N_2302);
or U2452 (N_2452,N_2324,N_2362);
or U2453 (N_2453,N_2393,N_2368);
or U2454 (N_2454,N_2385,N_2386);
or U2455 (N_2455,N_2362,N_2329);
and U2456 (N_2456,N_2377,N_2303);
nor U2457 (N_2457,N_2358,N_2353);
and U2458 (N_2458,N_2340,N_2306);
nand U2459 (N_2459,N_2340,N_2332);
or U2460 (N_2460,N_2344,N_2379);
or U2461 (N_2461,N_2385,N_2306);
or U2462 (N_2462,N_2396,N_2324);
nor U2463 (N_2463,N_2369,N_2347);
and U2464 (N_2464,N_2332,N_2345);
and U2465 (N_2465,N_2340,N_2398);
and U2466 (N_2466,N_2357,N_2335);
nand U2467 (N_2467,N_2313,N_2388);
or U2468 (N_2468,N_2347,N_2352);
nand U2469 (N_2469,N_2378,N_2398);
and U2470 (N_2470,N_2319,N_2388);
and U2471 (N_2471,N_2374,N_2384);
or U2472 (N_2472,N_2335,N_2376);
or U2473 (N_2473,N_2376,N_2364);
nand U2474 (N_2474,N_2348,N_2328);
nor U2475 (N_2475,N_2324,N_2336);
nor U2476 (N_2476,N_2348,N_2397);
or U2477 (N_2477,N_2345,N_2382);
and U2478 (N_2478,N_2313,N_2301);
or U2479 (N_2479,N_2310,N_2376);
and U2480 (N_2480,N_2391,N_2301);
and U2481 (N_2481,N_2345,N_2324);
or U2482 (N_2482,N_2394,N_2302);
and U2483 (N_2483,N_2371,N_2362);
or U2484 (N_2484,N_2337,N_2364);
and U2485 (N_2485,N_2395,N_2302);
nor U2486 (N_2486,N_2376,N_2392);
or U2487 (N_2487,N_2300,N_2352);
or U2488 (N_2488,N_2325,N_2343);
xor U2489 (N_2489,N_2313,N_2386);
nor U2490 (N_2490,N_2353,N_2367);
and U2491 (N_2491,N_2306,N_2301);
nand U2492 (N_2492,N_2301,N_2365);
nor U2493 (N_2493,N_2321,N_2381);
and U2494 (N_2494,N_2323,N_2336);
and U2495 (N_2495,N_2393,N_2398);
and U2496 (N_2496,N_2379,N_2366);
or U2497 (N_2497,N_2369,N_2346);
nand U2498 (N_2498,N_2395,N_2362);
or U2499 (N_2499,N_2332,N_2390);
nand U2500 (N_2500,N_2485,N_2405);
nand U2501 (N_2501,N_2467,N_2412);
or U2502 (N_2502,N_2468,N_2460);
nand U2503 (N_2503,N_2492,N_2474);
nor U2504 (N_2504,N_2495,N_2469);
nand U2505 (N_2505,N_2450,N_2487);
nor U2506 (N_2506,N_2421,N_2496);
nor U2507 (N_2507,N_2453,N_2428);
and U2508 (N_2508,N_2409,N_2435);
nand U2509 (N_2509,N_2401,N_2400);
or U2510 (N_2510,N_2480,N_2486);
and U2511 (N_2511,N_2461,N_2423);
and U2512 (N_2512,N_2406,N_2438);
and U2513 (N_2513,N_2430,N_2448);
nand U2514 (N_2514,N_2440,N_2493);
nor U2515 (N_2515,N_2481,N_2439);
or U2516 (N_2516,N_2410,N_2449);
nand U2517 (N_2517,N_2478,N_2452);
or U2518 (N_2518,N_2414,N_2484);
and U2519 (N_2519,N_2404,N_2475);
and U2520 (N_2520,N_2443,N_2498);
nand U2521 (N_2521,N_2402,N_2429);
nand U2522 (N_2522,N_2491,N_2419);
xor U2523 (N_2523,N_2456,N_2417);
nand U2524 (N_2524,N_2472,N_2442);
or U2525 (N_2525,N_2408,N_2477);
nand U2526 (N_2526,N_2462,N_2494);
nand U2527 (N_2527,N_2463,N_2407);
or U2528 (N_2528,N_2424,N_2489);
and U2529 (N_2529,N_2403,N_2488);
and U2530 (N_2530,N_2451,N_2427);
nand U2531 (N_2531,N_2482,N_2416);
nor U2532 (N_2532,N_2445,N_2411);
and U2533 (N_2533,N_2454,N_2465);
nand U2534 (N_2534,N_2459,N_2464);
or U2535 (N_2535,N_2499,N_2470);
nand U2536 (N_2536,N_2457,N_2466);
and U2537 (N_2537,N_2420,N_2490);
or U2538 (N_2538,N_2426,N_2415);
and U2539 (N_2539,N_2458,N_2473);
and U2540 (N_2540,N_2497,N_2436);
or U2541 (N_2541,N_2425,N_2476);
nand U2542 (N_2542,N_2432,N_2479);
or U2543 (N_2543,N_2444,N_2418);
or U2544 (N_2544,N_2437,N_2455);
nand U2545 (N_2545,N_2483,N_2431);
nand U2546 (N_2546,N_2471,N_2413);
nor U2547 (N_2547,N_2433,N_2446);
or U2548 (N_2548,N_2434,N_2422);
or U2549 (N_2549,N_2447,N_2441);
and U2550 (N_2550,N_2477,N_2482);
or U2551 (N_2551,N_2429,N_2431);
or U2552 (N_2552,N_2477,N_2488);
nor U2553 (N_2553,N_2458,N_2433);
nor U2554 (N_2554,N_2434,N_2432);
or U2555 (N_2555,N_2494,N_2460);
nor U2556 (N_2556,N_2452,N_2404);
nor U2557 (N_2557,N_2424,N_2410);
or U2558 (N_2558,N_2438,N_2463);
nand U2559 (N_2559,N_2493,N_2495);
nand U2560 (N_2560,N_2421,N_2459);
and U2561 (N_2561,N_2461,N_2437);
or U2562 (N_2562,N_2480,N_2400);
nand U2563 (N_2563,N_2450,N_2493);
nand U2564 (N_2564,N_2401,N_2457);
and U2565 (N_2565,N_2413,N_2450);
nor U2566 (N_2566,N_2471,N_2415);
nor U2567 (N_2567,N_2477,N_2478);
and U2568 (N_2568,N_2492,N_2451);
and U2569 (N_2569,N_2498,N_2426);
nor U2570 (N_2570,N_2491,N_2417);
nor U2571 (N_2571,N_2414,N_2402);
nor U2572 (N_2572,N_2448,N_2478);
nand U2573 (N_2573,N_2488,N_2453);
nor U2574 (N_2574,N_2484,N_2466);
nand U2575 (N_2575,N_2448,N_2481);
and U2576 (N_2576,N_2452,N_2490);
nor U2577 (N_2577,N_2487,N_2467);
nor U2578 (N_2578,N_2414,N_2424);
and U2579 (N_2579,N_2479,N_2472);
nand U2580 (N_2580,N_2486,N_2484);
or U2581 (N_2581,N_2410,N_2473);
or U2582 (N_2582,N_2472,N_2447);
nand U2583 (N_2583,N_2441,N_2425);
or U2584 (N_2584,N_2459,N_2466);
or U2585 (N_2585,N_2481,N_2437);
and U2586 (N_2586,N_2403,N_2430);
or U2587 (N_2587,N_2400,N_2466);
and U2588 (N_2588,N_2402,N_2491);
or U2589 (N_2589,N_2440,N_2433);
or U2590 (N_2590,N_2439,N_2475);
or U2591 (N_2591,N_2445,N_2423);
and U2592 (N_2592,N_2487,N_2494);
nor U2593 (N_2593,N_2470,N_2480);
nand U2594 (N_2594,N_2486,N_2400);
nand U2595 (N_2595,N_2418,N_2480);
nor U2596 (N_2596,N_2414,N_2498);
nor U2597 (N_2597,N_2442,N_2463);
nand U2598 (N_2598,N_2402,N_2482);
nor U2599 (N_2599,N_2487,N_2411);
or U2600 (N_2600,N_2524,N_2525);
nand U2601 (N_2601,N_2544,N_2543);
or U2602 (N_2602,N_2501,N_2532);
nor U2603 (N_2603,N_2581,N_2589);
and U2604 (N_2604,N_2548,N_2550);
and U2605 (N_2605,N_2553,N_2515);
nand U2606 (N_2606,N_2552,N_2547);
and U2607 (N_2607,N_2564,N_2570);
nand U2608 (N_2608,N_2565,N_2514);
nor U2609 (N_2609,N_2500,N_2588);
nor U2610 (N_2610,N_2507,N_2587);
nor U2611 (N_2611,N_2556,N_2591);
nand U2612 (N_2612,N_2572,N_2577);
nand U2613 (N_2613,N_2545,N_2502);
or U2614 (N_2614,N_2546,N_2529);
and U2615 (N_2615,N_2539,N_2578);
or U2616 (N_2616,N_2509,N_2518);
and U2617 (N_2617,N_2516,N_2574);
nand U2618 (N_2618,N_2560,N_2521);
and U2619 (N_2619,N_2562,N_2557);
nand U2620 (N_2620,N_2585,N_2511);
nor U2621 (N_2621,N_2510,N_2541);
or U2622 (N_2622,N_2536,N_2520);
or U2623 (N_2623,N_2527,N_2594);
nand U2624 (N_2624,N_2586,N_2526);
nand U2625 (N_2625,N_2566,N_2505);
or U2626 (N_2626,N_2571,N_2579);
nand U2627 (N_2627,N_2568,N_2595);
and U2628 (N_2628,N_2596,N_2569);
nor U2629 (N_2629,N_2559,N_2558);
nand U2630 (N_2630,N_2573,N_2504);
nor U2631 (N_2631,N_2561,N_2583);
or U2632 (N_2632,N_2575,N_2537);
or U2633 (N_2633,N_2555,N_2563);
nand U2634 (N_2634,N_2567,N_2512);
and U2635 (N_2635,N_2592,N_2519);
and U2636 (N_2636,N_2554,N_2503);
or U2637 (N_2637,N_2534,N_2540);
or U2638 (N_2638,N_2508,N_2533);
xor U2639 (N_2639,N_2551,N_2576);
nand U2640 (N_2640,N_2593,N_2522);
nor U2641 (N_2641,N_2523,N_2580);
and U2642 (N_2642,N_2582,N_2538);
and U2643 (N_2643,N_2513,N_2542);
nor U2644 (N_2644,N_2584,N_2530);
and U2645 (N_2645,N_2599,N_2517);
nor U2646 (N_2646,N_2590,N_2528);
or U2647 (N_2647,N_2597,N_2535);
nand U2648 (N_2648,N_2549,N_2598);
or U2649 (N_2649,N_2531,N_2506);
nor U2650 (N_2650,N_2530,N_2591);
nand U2651 (N_2651,N_2500,N_2565);
nand U2652 (N_2652,N_2555,N_2552);
and U2653 (N_2653,N_2533,N_2565);
or U2654 (N_2654,N_2567,N_2595);
or U2655 (N_2655,N_2532,N_2522);
nand U2656 (N_2656,N_2583,N_2531);
and U2657 (N_2657,N_2575,N_2570);
nand U2658 (N_2658,N_2560,N_2597);
or U2659 (N_2659,N_2502,N_2541);
or U2660 (N_2660,N_2530,N_2541);
and U2661 (N_2661,N_2501,N_2593);
nand U2662 (N_2662,N_2527,N_2569);
nand U2663 (N_2663,N_2551,N_2557);
and U2664 (N_2664,N_2590,N_2559);
nand U2665 (N_2665,N_2588,N_2544);
nor U2666 (N_2666,N_2540,N_2586);
nor U2667 (N_2667,N_2545,N_2574);
and U2668 (N_2668,N_2562,N_2525);
and U2669 (N_2669,N_2565,N_2505);
nor U2670 (N_2670,N_2592,N_2508);
and U2671 (N_2671,N_2593,N_2578);
nand U2672 (N_2672,N_2570,N_2576);
nand U2673 (N_2673,N_2530,N_2597);
and U2674 (N_2674,N_2507,N_2543);
nand U2675 (N_2675,N_2552,N_2577);
and U2676 (N_2676,N_2560,N_2578);
nand U2677 (N_2677,N_2546,N_2568);
nor U2678 (N_2678,N_2526,N_2560);
and U2679 (N_2679,N_2533,N_2545);
nand U2680 (N_2680,N_2524,N_2569);
or U2681 (N_2681,N_2547,N_2562);
and U2682 (N_2682,N_2540,N_2544);
or U2683 (N_2683,N_2541,N_2572);
nor U2684 (N_2684,N_2543,N_2502);
nand U2685 (N_2685,N_2546,N_2589);
and U2686 (N_2686,N_2557,N_2539);
nor U2687 (N_2687,N_2500,N_2593);
nor U2688 (N_2688,N_2539,N_2506);
nor U2689 (N_2689,N_2521,N_2557);
nor U2690 (N_2690,N_2563,N_2579);
and U2691 (N_2691,N_2510,N_2581);
nand U2692 (N_2692,N_2520,N_2528);
nor U2693 (N_2693,N_2554,N_2518);
and U2694 (N_2694,N_2596,N_2502);
and U2695 (N_2695,N_2572,N_2540);
or U2696 (N_2696,N_2576,N_2510);
and U2697 (N_2697,N_2531,N_2548);
and U2698 (N_2698,N_2566,N_2575);
and U2699 (N_2699,N_2547,N_2572);
or U2700 (N_2700,N_2666,N_2628);
and U2701 (N_2701,N_2623,N_2654);
or U2702 (N_2702,N_2691,N_2676);
nand U2703 (N_2703,N_2604,N_2613);
nor U2704 (N_2704,N_2614,N_2645);
xnor U2705 (N_2705,N_2617,N_2658);
and U2706 (N_2706,N_2675,N_2649);
nor U2707 (N_2707,N_2609,N_2626);
and U2708 (N_2708,N_2674,N_2684);
and U2709 (N_2709,N_2660,N_2632);
nand U2710 (N_2710,N_2622,N_2651);
or U2711 (N_2711,N_2681,N_2692);
nor U2712 (N_2712,N_2610,N_2616);
nor U2713 (N_2713,N_2693,N_2653);
or U2714 (N_2714,N_2690,N_2688);
nor U2715 (N_2715,N_2605,N_2668);
and U2716 (N_2716,N_2669,N_2615);
nand U2717 (N_2717,N_2663,N_2689);
and U2718 (N_2718,N_2656,N_2694);
nand U2719 (N_2719,N_2673,N_2621);
nor U2720 (N_2720,N_2601,N_2625);
xnor U2721 (N_2721,N_2655,N_2667);
nor U2722 (N_2722,N_2677,N_2606);
nor U2723 (N_2723,N_2665,N_2685);
nand U2724 (N_2724,N_2641,N_2607);
and U2725 (N_2725,N_2630,N_2608);
nand U2726 (N_2726,N_2648,N_2679);
nand U2727 (N_2727,N_2646,N_2687);
nor U2728 (N_2728,N_2631,N_2603);
and U2729 (N_2729,N_2624,N_2671);
nand U2730 (N_2730,N_2697,N_2636);
and U2731 (N_2731,N_2652,N_2659);
or U2732 (N_2732,N_2643,N_2638);
or U2733 (N_2733,N_2633,N_2642);
and U2734 (N_2734,N_2612,N_2695);
nand U2735 (N_2735,N_2634,N_2678);
nand U2736 (N_2736,N_2657,N_2672);
and U2737 (N_2737,N_2618,N_2662);
nor U2738 (N_2738,N_2680,N_2637);
or U2739 (N_2739,N_2670,N_2635);
and U2740 (N_2740,N_2650,N_2600);
nor U2741 (N_2741,N_2629,N_2639);
nor U2742 (N_2742,N_2664,N_2640);
and U2743 (N_2743,N_2699,N_2682);
and U2744 (N_2744,N_2698,N_2647);
nand U2745 (N_2745,N_2683,N_2686);
or U2746 (N_2746,N_2644,N_2611);
and U2747 (N_2747,N_2620,N_2602);
and U2748 (N_2748,N_2696,N_2619);
nand U2749 (N_2749,N_2661,N_2627);
and U2750 (N_2750,N_2632,N_2674);
nand U2751 (N_2751,N_2676,N_2669);
and U2752 (N_2752,N_2680,N_2628);
and U2753 (N_2753,N_2641,N_2613);
nand U2754 (N_2754,N_2652,N_2685);
nor U2755 (N_2755,N_2676,N_2682);
nand U2756 (N_2756,N_2685,N_2616);
nor U2757 (N_2757,N_2627,N_2618);
nor U2758 (N_2758,N_2690,N_2659);
nand U2759 (N_2759,N_2603,N_2662);
nand U2760 (N_2760,N_2608,N_2632);
nor U2761 (N_2761,N_2643,N_2619);
nor U2762 (N_2762,N_2657,N_2678);
and U2763 (N_2763,N_2695,N_2694);
nand U2764 (N_2764,N_2683,N_2655);
and U2765 (N_2765,N_2632,N_2623);
nand U2766 (N_2766,N_2642,N_2678);
and U2767 (N_2767,N_2615,N_2608);
and U2768 (N_2768,N_2675,N_2613);
and U2769 (N_2769,N_2602,N_2648);
nand U2770 (N_2770,N_2600,N_2631);
or U2771 (N_2771,N_2668,N_2615);
and U2772 (N_2772,N_2691,N_2682);
and U2773 (N_2773,N_2670,N_2606);
or U2774 (N_2774,N_2690,N_2665);
and U2775 (N_2775,N_2699,N_2683);
nor U2776 (N_2776,N_2652,N_2693);
nand U2777 (N_2777,N_2681,N_2694);
nor U2778 (N_2778,N_2631,N_2674);
nand U2779 (N_2779,N_2679,N_2696);
nor U2780 (N_2780,N_2629,N_2608);
nand U2781 (N_2781,N_2614,N_2698);
and U2782 (N_2782,N_2676,N_2608);
or U2783 (N_2783,N_2614,N_2621);
and U2784 (N_2784,N_2656,N_2622);
nor U2785 (N_2785,N_2627,N_2652);
and U2786 (N_2786,N_2614,N_2690);
nand U2787 (N_2787,N_2634,N_2646);
nor U2788 (N_2788,N_2678,N_2610);
or U2789 (N_2789,N_2662,N_2631);
nor U2790 (N_2790,N_2692,N_2607);
nand U2791 (N_2791,N_2633,N_2634);
nand U2792 (N_2792,N_2632,N_2628);
or U2793 (N_2793,N_2673,N_2662);
or U2794 (N_2794,N_2642,N_2693);
nor U2795 (N_2795,N_2619,N_2654);
nand U2796 (N_2796,N_2629,N_2683);
and U2797 (N_2797,N_2640,N_2632);
and U2798 (N_2798,N_2629,N_2652);
or U2799 (N_2799,N_2683,N_2613);
or U2800 (N_2800,N_2775,N_2754);
nor U2801 (N_2801,N_2755,N_2782);
nor U2802 (N_2802,N_2781,N_2723);
nand U2803 (N_2803,N_2774,N_2709);
nor U2804 (N_2804,N_2795,N_2797);
nand U2805 (N_2805,N_2794,N_2768);
nor U2806 (N_2806,N_2771,N_2776);
and U2807 (N_2807,N_2714,N_2791);
or U2808 (N_2808,N_2779,N_2746);
nand U2809 (N_2809,N_2785,N_2735);
and U2810 (N_2810,N_2784,N_2741);
nor U2811 (N_2811,N_2748,N_2701);
nand U2812 (N_2812,N_2716,N_2772);
or U2813 (N_2813,N_2793,N_2733);
nand U2814 (N_2814,N_2749,N_2719);
and U2815 (N_2815,N_2712,N_2777);
nand U2816 (N_2816,N_2770,N_2713);
nor U2817 (N_2817,N_2758,N_2773);
nand U2818 (N_2818,N_2710,N_2727);
nand U2819 (N_2819,N_2750,N_2769);
and U2820 (N_2820,N_2762,N_2706);
nand U2821 (N_2821,N_2757,N_2765);
nor U2822 (N_2822,N_2729,N_2708);
nand U2823 (N_2823,N_2792,N_2742);
and U2824 (N_2824,N_2778,N_2767);
and U2825 (N_2825,N_2720,N_2730);
nand U2826 (N_2826,N_2752,N_2780);
nor U2827 (N_2827,N_2707,N_2722);
nand U2828 (N_2828,N_2761,N_2798);
nand U2829 (N_2829,N_2799,N_2740);
or U2830 (N_2830,N_2738,N_2744);
nor U2831 (N_2831,N_2724,N_2711);
or U2832 (N_2832,N_2715,N_2783);
and U2833 (N_2833,N_2736,N_2725);
xnor U2834 (N_2834,N_2796,N_2700);
nand U2835 (N_2835,N_2788,N_2728);
nand U2836 (N_2836,N_2702,N_2745);
nand U2837 (N_2837,N_2760,N_2766);
nor U2838 (N_2838,N_2790,N_2717);
xor U2839 (N_2839,N_2786,N_2739);
nor U2840 (N_2840,N_2787,N_2704);
nand U2841 (N_2841,N_2743,N_2734);
and U2842 (N_2842,N_2751,N_2747);
or U2843 (N_2843,N_2763,N_2732);
nor U2844 (N_2844,N_2756,N_2789);
nor U2845 (N_2845,N_2753,N_2703);
nor U2846 (N_2846,N_2737,N_2764);
nor U2847 (N_2847,N_2726,N_2705);
or U2848 (N_2848,N_2721,N_2731);
nor U2849 (N_2849,N_2718,N_2759);
and U2850 (N_2850,N_2766,N_2776);
nand U2851 (N_2851,N_2741,N_2760);
or U2852 (N_2852,N_2754,N_2764);
nand U2853 (N_2853,N_2730,N_2761);
and U2854 (N_2854,N_2756,N_2743);
or U2855 (N_2855,N_2728,N_2740);
nand U2856 (N_2856,N_2717,N_2770);
or U2857 (N_2857,N_2702,N_2747);
and U2858 (N_2858,N_2703,N_2775);
nand U2859 (N_2859,N_2732,N_2791);
nand U2860 (N_2860,N_2759,N_2728);
and U2861 (N_2861,N_2729,N_2792);
nand U2862 (N_2862,N_2740,N_2718);
nand U2863 (N_2863,N_2755,N_2701);
nor U2864 (N_2864,N_2777,N_2769);
nor U2865 (N_2865,N_2785,N_2739);
nand U2866 (N_2866,N_2785,N_2709);
and U2867 (N_2867,N_2786,N_2794);
nand U2868 (N_2868,N_2791,N_2793);
or U2869 (N_2869,N_2746,N_2726);
nor U2870 (N_2870,N_2722,N_2751);
and U2871 (N_2871,N_2754,N_2724);
or U2872 (N_2872,N_2791,N_2759);
nand U2873 (N_2873,N_2765,N_2747);
or U2874 (N_2874,N_2715,N_2781);
nand U2875 (N_2875,N_2733,N_2758);
nor U2876 (N_2876,N_2708,N_2701);
or U2877 (N_2877,N_2761,N_2760);
and U2878 (N_2878,N_2716,N_2784);
nor U2879 (N_2879,N_2782,N_2775);
nor U2880 (N_2880,N_2734,N_2786);
nand U2881 (N_2881,N_2745,N_2758);
nand U2882 (N_2882,N_2781,N_2725);
nand U2883 (N_2883,N_2769,N_2703);
or U2884 (N_2884,N_2717,N_2756);
and U2885 (N_2885,N_2794,N_2778);
or U2886 (N_2886,N_2755,N_2770);
nand U2887 (N_2887,N_2726,N_2744);
or U2888 (N_2888,N_2781,N_2729);
or U2889 (N_2889,N_2793,N_2789);
nor U2890 (N_2890,N_2731,N_2743);
nor U2891 (N_2891,N_2732,N_2762);
nand U2892 (N_2892,N_2703,N_2738);
nor U2893 (N_2893,N_2750,N_2714);
or U2894 (N_2894,N_2774,N_2729);
or U2895 (N_2895,N_2708,N_2733);
and U2896 (N_2896,N_2786,N_2779);
nand U2897 (N_2897,N_2747,N_2724);
or U2898 (N_2898,N_2728,N_2784);
nor U2899 (N_2899,N_2784,N_2759);
and U2900 (N_2900,N_2814,N_2882);
or U2901 (N_2901,N_2849,N_2894);
and U2902 (N_2902,N_2840,N_2818);
nand U2903 (N_2903,N_2846,N_2823);
nor U2904 (N_2904,N_2830,N_2809);
nor U2905 (N_2905,N_2839,N_2880);
nor U2906 (N_2906,N_2811,N_2884);
nand U2907 (N_2907,N_2820,N_2881);
or U2908 (N_2908,N_2890,N_2843);
nor U2909 (N_2909,N_2803,N_2850);
or U2910 (N_2910,N_2885,N_2805);
nand U2911 (N_2911,N_2853,N_2871);
nor U2912 (N_2912,N_2868,N_2808);
or U2913 (N_2913,N_2867,N_2841);
xor U2914 (N_2914,N_2817,N_2876);
nor U2915 (N_2915,N_2842,N_2821);
and U2916 (N_2916,N_2801,N_2832);
nor U2917 (N_2917,N_2896,N_2870);
nand U2918 (N_2918,N_2813,N_2855);
and U2919 (N_2919,N_2831,N_2858);
or U2920 (N_2920,N_2854,N_2852);
xnor U2921 (N_2921,N_2826,N_2861);
and U2922 (N_2922,N_2806,N_2822);
nand U2923 (N_2923,N_2834,N_2833);
nor U2924 (N_2924,N_2895,N_2845);
nor U2925 (N_2925,N_2878,N_2857);
and U2926 (N_2926,N_2835,N_2800);
and U2927 (N_2927,N_2838,N_2825);
nor U2928 (N_2928,N_2812,N_2802);
or U2929 (N_2929,N_2899,N_2828);
nor U2930 (N_2930,N_2887,N_2893);
and U2931 (N_2931,N_2877,N_2829);
nand U2932 (N_2932,N_2847,N_2810);
nand U2933 (N_2933,N_2898,N_2866);
and U2934 (N_2934,N_2824,N_2836);
nor U2935 (N_2935,N_2807,N_2873);
and U2936 (N_2936,N_2892,N_2860);
xnor U2937 (N_2937,N_2883,N_2886);
nand U2938 (N_2938,N_2875,N_2862);
nor U2939 (N_2939,N_2819,N_2865);
or U2940 (N_2940,N_2837,N_2897);
nand U2941 (N_2941,N_2872,N_2863);
nor U2942 (N_2942,N_2815,N_2889);
nor U2943 (N_2943,N_2874,N_2816);
nand U2944 (N_2944,N_2888,N_2891);
nand U2945 (N_2945,N_2856,N_2864);
or U2946 (N_2946,N_2848,N_2844);
nand U2947 (N_2947,N_2827,N_2879);
nor U2948 (N_2948,N_2869,N_2859);
nand U2949 (N_2949,N_2804,N_2851);
nand U2950 (N_2950,N_2828,N_2891);
or U2951 (N_2951,N_2841,N_2872);
or U2952 (N_2952,N_2888,N_2897);
xor U2953 (N_2953,N_2845,N_2827);
nand U2954 (N_2954,N_2808,N_2845);
nor U2955 (N_2955,N_2832,N_2812);
nand U2956 (N_2956,N_2871,N_2879);
and U2957 (N_2957,N_2896,N_2861);
nor U2958 (N_2958,N_2874,N_2807);
nor U2959 (N_2959,N_2818,N_2845);
or U2960 (N_2960,N_2868,N_2838);
nand U2961 (N_2961,N_2888,N_2828);
and U2962 (N_2962,N_2894,N_2802);
or U2963 (N_2963,N_2898,N_2837);
nor U2964 (N_2964,N_2839,N_2812);
or U2965 (N_2965,N_2856,N_2841);
nand U2966 (N_2966,N_2838,N_2830);
nand U2967 (N_2967,N_2829,N_2887);
nor U2968 (N_2968,N_2811,N_2879);
or U2969 (N_2969,N_2853,N_2856);
nand U2970 (N_2970,N_2828,N_2858);
and U2971 (N_2971,N_2858,N_2867);
and U2972 (N_2972,N_2835,N_2897);
and U2973 (N_2973,N_2833,N_2890);
and U2974 (N_2974,N_2816,N_2825);
nand U2975 (N_2975,N_2833,N_2826);
and U2976 (N_2976,N_2831,N_2876);
and U2977 (N_2977,N_2894,N_2896);
and U2978 (N_2978,N_2874,N_2886);
nand U2979 (N_2979,N_2801,N_2830);
nand U2980 (N_2980,N_2837,N_2835);
nor U2981 (N_2981,N_2892,N_2843);
nand U2982 (N_2982,N_2881,N_2828);
nand U2983 (N_2983,N_2888,N_2839);
or U2984 (N_2984,N_2899,N_2888);
nor U2985 (N_2985,N_2809,N_2824);
and U2986 (N_2986,N_2843,N_2881);
nor U2987 (N_2987,N_2882,N_2895);
or U2988 (N_2988,N_2809,N_2882);
xnor U2989 (N_2989,N_2821,N_2848);
or U2990 (N_2990,N_2897,N_2809);
nor U2991 (N_2991,N_2837,N_2841);
nand U2992 (N_2992,N_2831,N_2877);
nand U2993 (N_2993,N_2897,N_2827);
or U2994 (N_2994,N_2848,N_2830);
nand U2995 (N_2995,N_2843,N_2852);
nand U2996 (N_2996,N_2862,N_2843);
or U2997 (N_2997,N_2890,N_2855);
nor U2998 (N_2998,N_2865,N_2848);
and U2999 (N_2999,N_2884,N_2837);
nand UO_0 (O_0,N_2928,N_2922);
nor UO_1 (O_1,N_2949,N_2965);
nand UO_2 (O_2,N_2931,N_2902);
nor UO_3 (O_3,N_2907,N_2956);
or UO_4 (O_4,N_2979,N_2984);
nor UO_5 (O_5,N_2978,N_2955);
and UO_6 (O_6,N_2992,N_2975);
and UO_7 (O_7,N_2939,N_2990);
nor UO_8 (O_8,N_2901,N_2926);
nor UO_9 (O_9,N_2910,N_2927);
or UO_10 (O_10,N_2969,N_2974);
nand UO_11 (O_11,N_2905,N_2976);
or UO_12 (O_12,N_2913,N_2929);
nand UO_13 (O_13,N_2967,N_2982);
or UO_14 (O_14,N_2914,N_2997);
nor UO_15 (O_15,N_2917,N_2964);
nand UO_16 (O_16,N_2942,N_2930);
or UO_17 (O_17,N_2957,N_2953);
nand UO_18 (O_18,N_2985,N_2934);
nand UO_19 (O_19,N_2971,N_2989);
or UO_20 (O_20,N_2912,N_2948);
nand UO_21 (O_21,N_2911,N_2958);
nor UO_22 (O_22,N_2983,N_2909);
nand UO_23 (O_23,N_2998,N_2915);
or UO_24 (O_24,N_2943,N_2945);
and UO_25 (O_25,N_2924,N_2951);
or UO_26 (O_26,N_2986,N_2973);
nand UO_27 (O_27,N_2937,N_2921);
or UO_28 (O_28,N_2968,N_2987);
nor UO_29 (O_29,N_2954,N_2996);
nand UO_30 (O_30,N_2944,N_2991);
or UO_31 (O_31,N_2946,N_2963);
or UO_32 (O_32,N_2960,N_2977);
or UO_33 (O_33,N_2933,N_2904);
and UO_34 (O_34,N_2993,N_2966);
or UO_35 (O_35,N_2938,N_2900);
or UO_36 (O_36,N_2947,N_2919);
and UO_37 (O_37,N_2972,N_2950);
or UO_38 (O_38,N_2961,N_2941);
and UO_39 (O_39,N_2920,N_2988);
and UO_40 (O_40,N_2981,N_2916);
nor UO_41 (O_41,N_2923,N_2970);
or UO_42 (O_42,N_2995,N_2940);
and UO_43 (O_43,N_2906,N_2952);
or UO_44 (O_44,N_2903,N_2959);
nand UO_45 (O_45,N_2908,N_2918);
nand UO_46 (O_46,N_2925,N_2980);
nor UO_47 (O_47,N_2999,N_2936);
nor UO_48 (O_48,N_2932,N_2935);
nand UO_49 (O_49,N_2962,N_2994);
and UO_50 (O_50,N_2968,N_2967);
and UO_51 (O_51,N_2946,N_2988);
nor UO_52 (O_52,N_2942,N_2991);
nor UO_53 (O_53,N_2932,N_2969);
nand UO_54 (O_54,N_2951,N_2996);
or UO_55 (O_55,N_2943,N_2907);
nand UO_56 (O_56,N_2983,N_2938);
nor UO_57 (O_57,N_2932,N_2971);
nor UO_58 (O_58,N_2937,N_2927);
or UO_59 (O_59,N_2954,N_2935);
nor UO_60 (O_60,N_2990,N_2945);
nand UO_61 (O_61,N_2961,N_2900);
nand UO_62 (O_62,N_2925,N_2908);
and UO_63 (O_63,N_2901,N_2995);
and UO_64 (O_64,N_2924,N_2982);
and UO_65 (O_65,N_2957,N_2965);
and UO_66 (O_66,N_2928,N_2943);
nand UO_67 (O_67,N_2940,N_2984);
and UO_68 (O_68,N_2986,N_2988);
nand UO_69 (O_69,N_2956,N_2932);
nor UO_70 (O_70,N_2988,N_2951);
nand UO_71 (O_71,N_2975,N_2950);
nand UO_72 (O_72,N_2904,N_2912);
or UO_73 (O_73,N_2930,N_2985);
nor UO_74 (O_74,N_2946,N_2907);
and UO_75 (O_75,N_2936,N_2979);
or UO_76 (O_76,N_2923,N_2922);
nand UO_77 (O_77,N_2917,N_2901);
or UO_78 (O_78,N_2963,N_2952);
nand UO_79 (O_79,N_2929,N_2924);
or UO_80 (O_80,N_2922,N_2979);
or UO_81 (O_81,N_2989,N_2900);
and UO_82 (O_82,N_2944,N_2976);
or UO_83 (O_83,N_2996,N_2994);
and UO_84 (O_84,N_2907,N_2982);
or UO_85 (O_85,N_2937,N_2934);
nand UO_86 (O_86,N_2910,N_2955);
and UO_87 (O_87,N_2924,N_2978);
and UO_88 (O_88,N_2971,N_2996);
and UO_89 (O_89,N_2908,N_2932);
or UO_90 (O_90,N_2958,N_2968);
and UO_91 (O_91,N_2904,N_2986);
nor UO_92 (O_92,N_2996,N_2988);
nor UO_93 (O_93,N_2911,N_2999);
nand UO_94 (O_94,N_2992,N_2917);
nand UO_95 (O_95,N_2917,N_2981);
and UO_96 (O_96,N_2932,N_2902);
nor UO_97 (O_97,N_2924,N_2925);
or UO_98 (O_98,N_2945,N_2927);
nor UO_99 (O_99,N_2937,N_2983);
nor UO_100 (O_100,N_2923,N_2926);
and UO_101 (O_101,N_2917,N_2928);
and UO_102 (O_102,N_2983,N_2959);
nand UO_103 (O_103,N_2952,N_2944);
nor UO_104 (O_104,N_2920,N_2939);
nand UO_105 (O_105,N_2979,N_2961);
and UO_106 (O_106,N_2989,N_2904);
nor UO_107 (O_107,N_2960,N_2983);
nor UO_108 (O_108,N_2993,N_2960);
xnor UO_109 (O_109,N_2952,N_2972);
or UO_110 (O_110,N_2939,N_2962);
nand UO_111 (O_111,N_2912,N_2940);
nor UO_112 (O_112,N_2959,N_2972);
nand UO_113 (O_113,N_2934,N_2909);
nand UO_114 (O_114,N_2936,N_2983);
and UO_115 (O_115,N_2922,N_2910);
nand UO_116 (O_116,N_2949,N_2958);
or UO_117 (O_117,N_2946,N_2910);
or UO_118 (O_118,N_2934,N_2914);
nor UO_119 (O_119,N_2973,N_2951);
and UO_120 (O_120,N_2962,N_2960);
nor UO_121 (O_121,N_2966,N_2957);
and UO_122 (O_122,N_2960,N_2992);
nand UO_123 (O_123,N_2995,N_2956);
nand UO_124 (O_124,N_2927,N_2993);
and UO_125 (O_125,N_2931,N_2911);
nand UO_126 (O_126,N_2979,N_2952);
or UO_127 (O_127,N_2920,N_2963);
or UO_128 (O_128,N_2969,N_2978);
and UO_129 (O_129,N_2998,N_2903);
or UO_130 (O_130,N_2985,N_2978);
nor UO_131 (O_131,N_2957,N_2902);
nor UO_132 (O_132,N_2993,N_2909);
and UO_133 (O_133,N_2920,N_2969);
and UO_134 (O_134,N_2979,N_2924);
nand UO_135 (O_135,N_2915,N_2966);
or UO_136 (O_136,N_2981,N_2929);
and UO_137 (O_137,N_2930,N_2966);
or UO_138 (O_138,N_2931,N_2919);
and UO_139 (O_139,N_2934,N_2995);
nor UO_140 (O_140,N_2925,N_2910);
nor UO_141 (O_141,N_2982,N_2938);
or UO_142 (O_142,N_2912,N_2966);
or UO_143 (O_143,N_2923,N_2908);
nor UO_144 (O_144,N_2977,N_2932);
nor UO_145 (O_145,N_2916,N_2965);
and UO_146 (O_146,N_2990,N_2986);
nand UO_147 (O_147,N_2991,N_2962);
nand UO_148 (O_148,N_2954,N_2923);
and UO_149 (O_149,N_2949,N_2959);
nor UO_150 (O_150,N_2996,N_2926);
nand UO_151 (O_151,N_2950,N_2910);
or UO_152 (O_152,N_2918,N_2967);
or UO_153 (O_153,N_2986,N_2979);
or UO_154 (O_154,N_2996,N_2997);
or UO_155 (O_155,N_2966,N_2974);
nor UO_156 (O_156,N_2948,N_2902);
nor UO_157 (O_157,N_2914,N_2990);
nor UO_158 (O_158,N_2954,N_2949);
nor UO_159 (O_159,N_2941,N_2907);
or UO_160 (O_160,N_2933,N_2938);
nor UO_161 (O_161,N_2942,N_2980);
nor UO_162 (O_162,N_2925,N_2934);
and UO_163 (O_163,N_2910,N_2937);
or UO_164 (O_164,N_2957,N_2911);
or UO_165 (O_165,N_2902,N_2901);
or UO_166 (O_166,N_2987,N_2938);
and UO_167 (O_167,N_2975,N_2900);
or UO_168 (O_168,N_2929,N_2919);
nand UO_169 (O_169,N_2987,N_2920);
and UO_170 (O_170,N_2986,N_2956);
nor UO_171 (O_171,N_2900,N_2955);
nor UO_172 (O_172,N_2926,N_2964);
nor UO_173 (O_173,N_2969,N_2941);
nor UO_174 (O_174,N_2929,N_2979);
nand UO_175 (O_175,N_2955,N_2992);
nand UO_176 (O_176,N_2982,N_2916);
nor UO_177 (O_177,N_2983,N_2988);
or UO_178 (O_178,N_2918,N_2952);
and UO_179 (O_179,N_2966,N_2918);
or UO_180 (O_180,N_2976,N_2922);
xor UO_181 (O_181,N_2978,N_2990);
nand UO_182 (O_182,N_2927,N_2930);
or UO_183 (O_183,N_2910,N_2914);
nand UO_184 (O_184,N_2939,N_2946);
nand UO_185 (O_185,N_2957,N_2973);
nor UO_186 (O_186,N_2941,N_2942);
or UO_187 (O_187,N_2952,N_2962);
and UO_188 (O_188,N_2984,N_2982);
nor UO_189 (O_189,N_2921,N_2976);
nor UO_190 (O_190,N_2936,N_2903);
nand UO_191 (O_191,N_2909,N_2941);
or UO_192 (O_192,N_2945,N_2941);
nor UO_193 (O_193,N_2916,N_2992);
and UO_194 (O_194,N_2902,N_2959);
and UO_195 (O_195,N_2903,N_2924);
and UO_196 (O_196,N_2989,N_2914);
or UO_197 (O_197,N_2923,N_2933);
nor UO_198 (O_198,N_2990,N_2983);
and UO_199 (O_199,N_2935,N_2928);
nor UO_200 (O_200,N_2942,N_2900);
or UO_201 (O_201,N_2959,N_2901);
or UO_202 (O_202,N_2958,N_2935);
nand UO_203 (O_203,N_2930,N_2960);
nor UO_204 (O_204,N_2952,N_2933);
nor UO_205 (O_205,N_2925,N_2937);
and UO_206 (O_206,N_2914,N_2905);
or UO_207 (O_207,N_2997,N_2926);
nand UO_208 (O_208,N_2943,N_2953);
or UO_209 (O_209,N_2978,N_2930);
or UO_210 (O_210,N_2979,N_2944);
or UO_211 (O_211,N_2925,N_2922);
and UO_212 (O_212,N_2977,N_2954);
nor UO_213 (O_213,N_2935,N_2940);
and UO_214 (O_214,N_2919,N_2923);
and UO_215 (O_215,N_2952,N_2954);
and UO_216 (O_216,N_2963,N_2923);
nand UO_217 (O_217,N_2919,N_2932);
or UO_218 (O_218,N_2997,N_2972);
or UO_219 (O_219,N_2935,N_2951);
or UO_220 (O_220,N_2901,N_2940);
nand UO_221 (O_221,N_2983,N_2972);
nor UO_222 (O_222,N_2970,N_2935);
nand UO_223 (O_223,N_2933,N_2934);
and UO_224 (O_224,N_2980,N_2927);
nand UO_225 (O_225,N_2969,N_2998);
and UO_226 (O_226,N_2920,N_2999);
and UO_227 (O_227,N_2907,N_2934);
and UO_228 (O_228,N_2906,N_2996);
nor UO_229 (O_229,N_2911,N_2929);
and UO_230 (O_230,N_2940,N_2989);
nand UO_231 (O_231,N_2983,N_2968);
and UO_232 (O_232,N_2991,N_2900);
and UO_233 (O_233,N_2939,N_2921);
or UO_234 (O_234,N_2970,N_2931);
or UO_235 (O_235,N_2945,N_2974);
xnor UO_236 (O_236,N_2995,N_2992);
nor UO_237 (O_237,N_2921,N_2969);
or UO_238 (O_238,N_2991,N_2957);
nor UO_239 (O_239,N_2947,N_2927);
or UO_240 (O_240,N_2982,N_2949);
or UO_241 (O_241,N_2989,N_2950);
and UO_242 (O_242,N_2902,N_2978);
nor UO_243 (O_243,N_2996,N_2944);
nor UO_244 (O_244,N_2987,N_2982);
and UO_245 (O_245,N_2997,N_2944);
nand UO_246 (O_246,N_2974,N_2906);
or UO_247 (O_247,N_2905,N_2959);
nor UO_248 (O_248,N_2986,N_2960);
or UO_249 (O_249,N_2939,N_2985);
nor UO_250 (O_250,N_2928,N_2946);
nor UO_251 (O_251,N_2955,N_2973);
and UO_252 (O_252,N_2951,N_2905);
nor UO_253 (O_253,N_2920,N_2909);
nand UO_254 (O_254,N_2989,N_2963);
and UO_255 (O_255,N_2998,N_2962);
and UO_256 (O_256,N_2922,N_2930);
or UO_257 (O_257,N_2932,N_2942);
xnor UO_258 (O_258,N_2932,N_2960);
nand UO_259 (O_259,N_2922,N_2963);
nand UO_260 (O_260,N_2992,N_2948);
or UO_261 (O_261,N_2947,N_2989);
nor UO_262 (O_262,N_2970,N_2955);
or UO_263 (O_263,N_2975,N_2977);
nor UO_264 (O_264,N_2930,N_2970);
or UO_265 (O_265,N_2936,N_2900);
nor UO_266 (O_266,N_2906,N_2919);
or UO_267 (O_267,N_2911,N_2927);
or UO_268 (O_268,N_2938,N_2998);
nand UO_269 (O_269,N_2976,N_2993);
and UO_270 (O_270,N_2909,N_2998);
and UO_271 (O_271,N_2922,N_2991);
nor UO_272 (O_272,N_2997,N_2984);
and UO_273 (O_273,N_2937,N_2966);
and UO_274 (O_274,N_2993,N_2958);
nor UO_275 (O_275,N_2977,N_2934);
or UO_276 (O_276,N_2909,N_2936);
and UO_277 (O_277,N_2934,N_2981);
nor UO_278 (O_278,N_2919,N_2988);
and UO_279 (O_279,N_2973,N_2962);
and UO_280 (O_280,N_2903,N_2919);
xor UO_281 (O_281,N_2908,N_2931);
nand UO_282 (O_282,N_2977,N_2979);
and UO_283 (O_283,N_2938,N_2961);
and UO_284 (O_284,N_2936,N_2924);
nor UO_285 (O_285,N_2972,N_2909);
nor UO_286 (O_286,N_2978,N_2947);
nor UO_287 (O_287,N_2957,N_2924);
or UO_288 (O_288,N_2994,N_2933);
nand UO_289 (O_289,N_2928,N_2913);
and UO_290 (O_290,N_2925,N_2956);
nand UO_291 (O_291,N_2945,N_2906);
and UO_292 (O_292,N_2986,N_2908);
nand UO_293 (O_293,N_2937,N_2931);
and UO_294 (O_294,N_2937,N_2978);
and UO_295 (O_295,N_2972,N_2995);
nor UO_296 (O_296,N_2944,N_2929);
and UO_297 (O_297,N_2932,N_2927);
and UO_298 (O_298,N_2960,N_2917);
or UO_299 (O_299,N_2905,N_2950);
and UO_300 (O_300,N_2954,N_2927);
or UO_301 (O_301,N_2938,N_2995);
or UO_302 (O_302,N_2908,N_2984);
nor UO_303 (O_303,N_2988,N_2998);
or UO_304 (O_304,N_2979,N_2972);
and UO_305 (O_305,N_2944,N_2984);
and UO_306 (O_306,N_2934,N_2966);
nor UO_307 (O_307,N_2913,N_2915);
xor UO_308 (O_308,N_2970,N_2947);
nor UO_309 (O_309,N_2967,N_2963);
or UO_310 (O_310,N_2951,N_2900);
nor UO_311 (O_311,N_2987,N_2943);
nor UO_312 (O_312,N_2974,N_2999);
and UO_313 (O_313,N_2985,N_2905);
nor UO_314 (O_314,N_2943,N_2934);
or UO_315 (O_315,N_2984,N_2995);
or UO_316 (O_316,N_2972,N_2914);
nor UO_317 (O_317,N_2921,N_2918);
or UO_318 (O_318,N_2916,N_2978);
nand UO_319 (O_319,N_2926,N_2999);
nor UO_320 (O_320,N_2959,N_2952);
nor UO_321 (O_321,N_2952,N_2946);
and UO_322 (O_322,N_2949,N_2922);
or UO_323 (O_323,N_2961,N_2937);
nand UO_324 (O_324,N_2908,N_2912);
nand UO_325 (O_325,N_2936,N_2963);
and UO_326 (O_326,N_2947,N_2959);
nand UO_327 (O_327,N_2988,N_2930);
nor UO_328 (O_328,N_2908,N_2903);
nand UO_329 (O_329,N_2979,N_2976);
or UO_330 (O_330,N_2999,N_2962);
nor UO_331 (O_331,N_2940,N_2900);
and UO_332 (O_332,N_2952,N_2941);
or UO_333 (O_333,N_2960,N_2971);
nand UO_334 (O_334,N_2921,N_2931);
or UO_335 (O_335,N_2903,N_2934);
nand UO_336 (O_336,N_2908,N_2994);
nor UO_337 (O_337,N_2980,N_2932);
or UO_338 (O_338,N_2972,N_2907);
or UO_339 (O_339,N_2956,N_2928);
or UO_340 (O_340,N_2938,N_2984);
nor UO_341 (O_341,N_2988,N_2943);
nor UO_342 (O_342,N_2997,N_2915);
or UO_343 (O_343,N_2994,N_2965);
nand UO_344 (O_344,N_2953,N_2952);
and UO_345 (O_345,N_2905,N_2981);
or UO_346 (O_346,N_2949,N_2977);
and UO_347 (O_347,N_2926,N_2995);
and UO_348 (O_348,N_2972,N_2968);
or UO_349 (O_349,N_2939,N_2978);
and UO_350 (O_350,N_2925,N_2930);
nor UO_351 (O_351,N_2929,N_2959);
nor UO_352 (O_352,N_2913,N_2905);
or UO_353 (O_353,N_2934,N_2973);
or UO_354 (O_354,N_2947,N_2974);
nor UO_355 (O_355,N_2982,N_2956);
nor UO_356 (O_356,N_2965,N_2958);
nand UO_357 (O_357,N_2956,N_2911);
and UO_358 (O_358,N_2987,N_2971);
or UO_359 (O_359,N_2988,N_2985);
or UO_360 (O_360,N_2990,N_2951);
or UO_361 (O_361,N_2936,N_2914);
nor UO_362 (O_362,N_2918,N_2924);
or UO_363 (O_363,N_2916,N_2976);
nand UO_364 (O_364,N_2990,N_2913);
or UO_365 (O_365,N_2959,N_2958);
or UO_366 (O_366,N_2959,N_2937);
and UO_367 (O_367,N_2968,N_2986);
or UO_368 (O_368,N_2989,N_2941);
or UO_369 (O_369,N_2970,N_2908);
nand UO_370 (O_370,N_2955,N_2982);
nand UO_371 (O_371,N_2972,N_2935);
or UO_372 (O_372,N_2919,N_2937);
nand UO_373 (O_373,N_2925,N_2926);
and UO_374 (O_374,N_2931,N_2950);
and UO_375 (O_375,N_2957,N_2938);
and UO_376 (O_376,N_2930,N_2963);
and UO_377 (O_377,N_2913,N_2909);
nor UO_378 (O_378,N_2929,N_2937);
and UO_379 (O_379,N_2979,N_2985);
nor UO_380 (O_380,N_2992,N_2967);
nand UO_381 (O_381,N_2971,N_2942);
or UO_382 (O_382,N_2965,N_2982);
nand UO_383 (O_383,N_2942,N_2966);
nand UO_384 (O_384,N_2986,N_2911);
nor UO_385 (O_385,N_2938,N_2929);
or UO_386 (O_386,N_2909,N_2924);
or UO_387 (O_387,N_2964,N_2974);
nor UO_388 (O_388,N_2908,N_2982);
or UO_389 (O_389,N_2916,N_2914);
nor UO_390 (O_390,N_2908,N_2919);
and UO_391 (O_391,N_2917,N_2909);
nor UO_392 (O_392,N_2987,N_2980);
nor UO_393 (O_393,N_2917,N_2978);
and UO_394 (O_394,N_2955,N_2917);
or UO_395 (O_395,N_2916,N_2975);
and UO_396 (O_396,N_2975,N_2921);
nand UO_397 (O_397,N_2919,N_2957);
or UO_398 (O_398,N_2902,N_2967);
and UO_399 (O_399,N_2964,N_2943);
xnor UO_400 (O_400,N_2983,N_2945);
and UO_401 (O_401,N_2900,N_2928);
nand UO_402 (O_402,N_2907,N_2987);
nand UO_403 (O_403,N_2978,N_2960);
nor UO_404 (O_404,N_2912,N_2924);
nor UO_405 (O_405,N_2979,N_2909);
and UO_406 (O_406,N_2927,N_2917);
or UO_407 (O_407,N_2939,N_2955);
and UO_408 (O_408,N_2991,N_2987);
nand UO_409 (O_409,N_2956,N_2974);
and UO_410 (O_410,N_2925,N_2923);
and UO_411 (O_411,N_2993,N_2933);
or UO_412 (O_412,N_2949,N_2998);
or UO_413 (O_413,N_2984,N_2972);
nand UO_414 (O_414,N_2966,N_2917);
nand UO_415 (O_415,N_2925,N_2957);
and UO_416 (O_416,N_2954,N_2932);
nand UO_417 (O_417,N_2919,N_2948);
nand UO_418 (O_418,N_2912,N_2981);
or UO_419 (O_419,N_2983,N_2971);
or UO_420 (O_420,N_2976,N_2978);
and UO_421 (O_421,N_2943,N_2981);
and UO_422 (O_422,N_2904,N_2982);
nand UO_423 (O_423,N_2932,N_2930);
nand UO_424 (O_424,N_2902,N_2922);
nor UO_425 (O_425,N_2936,N_2961);
nor UO_426 (O_426,N_2959,N_2922);
and UO_427 (O_427,N_2954,N_2969);
nand UO_428 (O_428,N_2912,N_2955);
and UO_429 (O_429,N_2914,N_2929);
and UO_430 (O_430,N_2955,N_2906);
or UO_431 (O_431,N_2962,N_2982);
nor UO_432 (O_432,N_2950,N_2938);
or UO_433 (O_433,N_2974,N_2929);
nor UO_434 (O_434,N_2956,N_2934);
and UO_435 (O_435,N_2934,N_2942);
nor UO_436 (O_436,N_2960,N_2931);
and UO_437 (O_437,N_2972,N_2989);
or UO_438 (O_438,N_2966,N_2927);
nor UO_439 (O_439,N_2942,N_2954);
xor UO_440 (O_440,N_2954,N_2940);
and UO_441 (O_441,N_2960,N_2995);
and UO_442 (O_442,N_2945,N_2967);
nor UO_443 (O_443,N_2995,N_2997);
or UO_444 (O_444,N_2942,N_2994);
nand UO_445 (O_445,N_2971,N_2933);
or UO_446 (O_446,N_2966,N_2997);
nor UO_447 (O_447,N_2962,N_2919);
and UO_448 (O_448,N_2955,N_2998);
nand UO_449 (O_449,N_2940,N_2915);
and UO_450 (O_450,N_2953,N_2910);
nor UO_451 (O_451,N_2982,N_2953);
and UO_452 (O_452,N_2952,N_2947);
and UO_453 (O_453,N_2929,N_2916);
nand UO_454 (O_454,N_2938,N_2932);
nor UO_455 (O_455,N_2939,N_2952);
nor UO_456 (O_456,N_2958,N_2936);
nor UO_457 (O_457,N_2994,N_2957);
or UO_458 (O_458,N_2910,N_2999);
nand UO_459 (O_459,N_2944,N_2969);
nand UO_460 (O_460,N_2910,N_2934);
or UO_461 (O_461,N_2936,N_2976);
and UO_462 (O_462,N_2934,N_2950);
and UO_463 (O_463,N_2935,N_2938);
nand UO_464 (O_464,N_2930,N_2917);
nor UO_465 (O_465,N_2981,N_2930);
and UO_466 (O_466,N_2967,N_2970);
nand UO_467 (O_467,N_2988,N_2900);
and UO_468 (O_468,N_2951,N_2961);
and UO_469 (O_469,N_2931,N_2983);
nand UO_470 (O_470,N_2996,N_2952);
and UO_471 (O_471,N_2946,N_2964);
or UO_472 (O_472,N_2990,N_2992);
or UO_473 (O_473,N_2907,N_2904);
nand UO_474 (O_474,N_2975,N_2961);
nand UO_475 (O_475,N_2909,N_2976);
or UO_476 (O_476,N_2946,N_2927);
nand UO_477 (O_477,N_2983,N_2910);
or UO_478 (O_478,N_2948,N_2913);
and UO_479 (O_479,N_2991,N_2970);
or UO_480 (O_480,N_2971,N_2940);
nor UO_481 (O_481,N_2983,N_2950);
and UO_482 (O_482,N_2934,N_2901);
or UO_483 (O_483,N_2942,N_2922);
and UO_484 (O_484,N_2950,N_2933);
or UO_485 (O_485,N_2945,N_2950);
nand UO_486 (O_486,N_2901,N_2964);
and UO_487 (O_487,N_2966,N_2946);
nand UO_488 (O_488,N_2970,N_2957);
or UO_489 (O_489,N_2942,N_2929);
and UO_490 (O_490,N_2995,N_2935);
nor UO_491 (O_491,N_2992,N_2905);
and UO_492 (O_492,N_2967,N_2985);
nand UO_493 (O_493,N_2976,N_2953);
nand UO_494 (O_494,N_2928,N_2901);
nand UO_495 (O_495,N_2997,N_2954);
nor UO_496 (O_496,N_2929,N_2932);
nor UO_497 (O_497,N_2933,N_2951);
and UO_498 (O_498,N_2944,N_2916);
and UO_499 (O_499,N_2998,N_2919);
endmodule