module basic_2500_25000_3000_5_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_2103,In_688);
nor U1 (N_1,In_1365,In_1910);
or U2 (N_2,In_597,In_525);
nor U3 (N_3,In_1085,In_589);
nor U4 (N_4,In_1514,In_1699);
and U5 (N_5,In_1371,In_1171);
nor U6 (N_6,In_2183,In_738);
and U7 (N_7,In_1788,In_2086);
nor U8 (N_8,In_1813,In_224);
xnor U9 (N_9,In_1036,In_2264);
and U10 (N_10,In_1299,In_1223);
and U11 (N_11,In_2300,In_2393);
nand U12 (N_12,In_1951,In_148);
or U13 (N_13,In_423,In_2322);
and U14 (N_14,In_1852,In_674);
nor U15 (N_15,In_686,In_230);
or U16 (N_16,In_1193,In_1262);
and U17 (N_17,In_790,In_1661);
nor U18 (N_18,In_1793,In_1157);
or U19 (N_19,In_1521,In_664);
nor U20 (N_20,In_2464,In_784);
nor U21 (N_21,In_870,In_2447);
and U22 (N_22,In_1434,In_1055);
and U23 (N_23,In_1833,In_94);
or U24 (N_24,In_89,In_1447);
nand U25 (N_25,In_207,In_2313);
nor U26 (N_26,In_563,In_2198);
and U27 (N_27,In_1058,In_1473);
and U28 (N_28,In_438,In_275);
and U29 (N_29,In_1470,In_1240);
xor U30 (N_30,In_1501,In_454);
nand U31 (N_31,In_985,In_2437);
and U32 (N_32,In_1758,In_977);
nand U33 (N_33,In_278,In_2360);
nand U34 (N_34,In_994,In_2054);
or U35 (N_35,In_1149,In_1934);
nand U36 (N_36,In_1021,In_183);
nand U37 (N_37,In_86,In_893);
nand U38 (N_38,In_173,In_840);
and U39 (N_39,In_1771,In_1639);
and U40 (N_40,In_1052,In_2058);
and U41 (N_41,In_25,In_73);
or U42 (N_42,In_691,In_1790);
and U43 (N_43,In_2175,In_1257);
nand U44 (N_44,In_1696,In_759);
nor U45 (N_45,In_1125,In_960);
or U46 (N_46,In_2482,In_1814);
nor U47 (N_47,In_1121,In_622);
and U48 (N_48,In_2170,In_2476);
nor U49 (N_49,In_1566,In_1953);
and U50 (N_50,In_2239,In_1837);
nand U51 (N_51,In_2024,In_21);
or U52 (N_52,In_1358,In_270);
or U53 (N_53,In_1380,In_1682);
and U54 (N_54,In_1166,In_1153);
nand U55 (N_55,In_2108,In_2152);
or U56 (N_56,In_846,In_888);
xor U57 (N_57,In_1641,In_1264);
nor U58 (N_58,In_549,In_2295);
and U59 (N_59,In_1369,In_1513);
or U60 (N_60,In_699,In_1263);
nor U61 (N_61,In_1307,In_370);
xor U62 (N_62,In_1712,In_2299);
or U63 (N_63,In_1973,In_1030);
or U64 (N_64,In_1418,In_2163);
or U65 (N_65,In_1656,In_832);
nand U66 (N_66,In_1573,In_596);
or U67 (N_67,In_1607,In_872);
xor U68 (N_68,In_1700,In_1575);
and U69 (N_69,In_23,In_718);
nand U70 (N_70,In_277,In_49);
nand U71 (N_71,In_1714,In_584);
and U72 (N_72,In_1744,In_1594);
or U73 (N_73,In_740,In_1693);
or U74 (N_74,In_1342,In_1232);
or U75 (N_75,In_151,In_2235);
or U76 (N_76,In_624,In_179);
or U77 (N_77,In_1192,In_608);
nor U78 (N_78,In_407,In_362);
nand U79 (N_79,In_2277,In_1533);
nor U80 (N_80,In_783,In_1584);
nand U81 (N_81,In_2391,In_472);
nor U82 (N_82,In_159,In_2135);
or U83 (N_83,In_1968,In_2211);
nor U84 (N_84,In_511,In_1721);
and U85 (N_85,In_464,In_623);
or U86 (N_86,In_1912,In_1069);
or U87 (N_87,In_2387,In_2061);
or U88 (N_88,In_1853,In_1482);
or U89 (N_89,In_2439,In_1517);
and U90 (N_90,In_1260,In_786);
or U91 (N_91,In_1618,In_1511);
or U92 (N_92,In_1271,In_1003);
or U93 (N_93,In_1830,In_1590);
and U94 (N_94,In_1529,In_164);
xor U95 (N_95,In_1207,In_2319);
and U96 (N_96,In_2237,In_243);
or U97 (N_97,In_1218,In_1161);
nand U98 (N_98,In_1826,In_96);
or U99 (N_99,In_2094,In_765);
or U100 (N_100,In_105,In_1255);
nor U101 (N_101,In_2244,In_1976);
or U102 (N_102,In_1824,In_1905);
nor U103 (N_103,In_510,In_399);
or U104 (N_104,In_2029,In_487);
and U105 (N_105,In_1165,In_1914);
nor U106 (N_106,In_1659,In_2402);
xnor U107 (N_107,In_630,In_1298);
nor U108 (N_108,In_1782,In_926);
or U109 (N_109,In_530,In_273);
nand U110 (N_110,In_2017,In_614);
nand U111 (N_111,In_294,In_1624);
xnor U112 (N_112,In_848,In_1215);
nor U113 (N_113,In_1505,In_2261);
nor U114 (N_114,In_1010,In_601);
or U115 (N_115,In_282,In_1838);
and U116 (N_116,In_1295,In_489);
and U117 (N_117,In_1550,In_643);
nand U118 (N_118,In_1160,In_1754);
nor U119 (N_119,In_567,In_1448);
or U120 (N_120,In_1820,In_2341);
and U121 (N_121,In_1370,In_2310);
or U122 (N_122,In_353,In_514);
and U123 (N_123,In_1375,In_681);
nand U124 (N_124,In_1004,In_1679);
and U125 (N_125,In_861,In_2);
nor U126 (N_126,In_636,In_2263);
and U127 (N_127,In_1316,In_637);
or U128 (N_128,In_2499,In_1582);
and U129 (N_129,In_2106,In_2012);
nor U130 (N_130,In_390,In_2098);
and U131 (N_131,In_70,In_1797);
xor U132 (N_132,In_1416,In_42);
and U133 (N_133,In_760,In_857);
and U134 (N_134,In_312,In_989);
nor U135 (N_135,In_2425,In_196);
nor U136 (N_136,In_2355,In_283);
nor U137 (N_137,In_19,In_1775);
nand U138 (N_138,In_873,In_2326);
or U139 (N_139,In_2160,In_2398);
or U140 (N_140,In_695,In_1390);
xnor U141 (N_141,In_1178,In_112);
nand U142 (N_142,In_2129,In_359);
nor U143 (N_143,In_2265,In_1731);
nand U144 (N_144,In_949,In_225);
and U145 (N_145,In_1544,In_2035);
nor U146 (N_146,In_298,In_1631);
nor U147 (N_147,In_247,In_754);
nor U148 (N_148,In_841,In_1955);
and U149 (N_149,In_1426,In_1078);
nor U150 (N_150,In_743,In_1664);
and U151 (N_151,In_2060,In_1565);
nand U152 (N_152,In_2492,In_693);
or U153 (N_153,In_414,In_371);
nor U154 (N_154,In_2463,In_1620);
nand U155 (N_155,In_1488,In_1733);
and U156 (N_156,In_397,In_168);
nor U157 (N_157,In_2433,In_449);
nor U158 (N_158,In_2087,In_2409);
xnor U159 (N_159,In_2490,In_367);
nand U160 (N_160,In_280,In_1143);
or U161 (N_161,In_1174,In_2445);
and U162 (N_162,In_588,In_1972);
or U163 (N_163,In_2288,In_484);
nor U164 (N_164,In_2206,In_1116);
nor U165 (N_165,In_912,In_268);
nand U166 (N_166,In_1043,In_1847);
or U167 (N_167,In_331,In_1842);
nand U168 (N_168,In_809,In_1167);
or U169 (N_169,In_1547,In_385);
and U170 (N_170,In_866,In_2357);
or U171 (N_171,In_1431,In_1930);
xor U172 (N_172,In_130,In_1660);
and U173 (N_173,In_758,In_1858);
or U174 (N_174,In_160,In_658);
and U175 (N_175,In_742,In_1974);
nor U176 (N_176,In_188,In_1519);
nand U177 (N_177,In_2117,In_217);
nor U178 (N_178,In_1348,In_1466);
nor U179 (N_179,In_482,In_733);
nand U180 (N_180,In_36,In_2053);
and U181 (N_181,In_772,In_984);
nor U182 (N_182,In_381,In_248);
nand U183 (N_183,In_966,In_867);
or U184 (N_184,In_1610,In_1795);
and U185 (N_185,In_2291,In_2431);
nor U186 (N_186,In_97,In_1845);
nor U187 (N_187,In_2328,In_739);
nand U188 (N_188,In_1928,In_2189);
or U189 (N_189,In_1611,In_1224);
or U190 (N_190,In_1780,In_1366);
nor U191 (N_191,In_1132,In_1638);
xnor U192 (N_192,In_633,In_1635);
or U193 (N_193,In_405,In_1749);
or U194 (N_194,In_2336,In_1957);
nand U195 (N_195,In_120,In_1405);
nor U196 (N_196,In_137,In_1735);
nor U197 (N_197,In_1850,In_542);
nor U198 (N_198,In_2041,In_1381);
nor U199 (N_199,In_2411,In_43);
and U200 (N_200,In_1056,In_1927);
nor U201 (N_201,In_2259,In_1334);
nand U202 (N_202,In_1282,In_2217);
nand U203 (N_203,In_1233,In_1979);
and U204 (N_204,In_1269,In_1873);
or U205 (N_205,In_2469,In_2373);
nand U206 (N_206,In_1480,In_2304);
nor U207 (N_207,In_647,In_369);
nand U208 (N_208,In_1204,In_895);
xnor U209 (N_209,In_1322,In_950);
nor U210 (N_210,In_1290,In_610);
nor U211 (N_211,In_671,In_980);
or U212 (N_212,In_2050,In_347);
and U213 (N_213,In_1241,In_1146);
nor U214 (N_214,In_1015,In_1831);
nand U215 (N_215,In_1285,In_750);
or U216 (N_216,In_2231,In_1064);
and U217 (N_217,In_1076,In_901);
or U218 (N_218,In_198,In_1843);
or U219 (N_219,In_2361,In_1807);
and U220 (N_220,In_1595,In_890);
nand U221 (N_221,In_879,In_1008);
and U222 (N_222,In_138,In_1303);
and U223 (N_223,In_1092,In_1868);
nand U224 (N_224,In_92,In_2181);
xnor U225 (N_225,In_939,In_1190);
and U226 (N_226,In_2044,In_1516);
or U227 (N_227,In_85,In_2171);
nand U228 (N_228,In_2203,In_1235);
and U229 (N_229,In_1546,In_264);
nand U230 (N_230,In_1188,In_2009);
nor U231 (N_231,In_1420,In_2225);
nor U232 (N_232,In_690,In_561);
nor U233 (N_233,In_1561,In_330);
or U234 (N_234,In_2334,In_1162);
nand U235 (N_235,In_1701,In_654);
and U236 (N_236,In_1410,In_755);
or U237 (N_237,In_2455,In_1219);
nand U238 (N_238,In_1281,In_194);
nand U239 (N_239,In_1982,In_402);
or U240 (N_240,In_953,In_1096);
and U241 (N_241,In_2456,In_2333);
nor U242 (N_242,In_340,In_2089);
nor U243 (N_243,In_125,In_748);
or U244 (N_244,In_1892,In_779);
or U245 (N_245,In_1527,In_291);
or U246 (N_246,In_506,In_1343);
nor U247 (N_247,In_792,In_2369);
nand U248 (N_248,In_1265,In_618);
nor U249 (N_249,In_2283,In_1104);
or U250 (N_250,In_927,In_1086);
nand U251 (N_251,In_1574,In_1805);
nor U252 (N_252,In_613,In_579);
nand U253 (N_253,In_811,In_206);
nand U254 (N_254,In_887,In_925);
nand U255 (N_255,In_1267,In_673);
and U256 (N_256,In_805,In_1242);
and U257 (N_257,In_969,In_1942);
xor U258 (N_258,In_2120,In_37);
and U259 (N_259,In_2159,In_2424);
nand U260 (N_260,In_1960,In_982);
nand U261 (N_261,In_1177,In_426);
nand U262 (N_262,In_1938,In_413);
nand U263 (N_263,In_2475,In_1999);
and U264 (N_264,In_680,In_1323);
nor U265 (N_265,In_649,In_706);
nor U266 (N_266,In_851,In_1083);
and U267 (N_267,In_1238,In_1919);
nand U268 (N_268,In_2438,In_350);
and U269 (N_269,In_2386,In_136);
nor U270 (N_270,In_190,In_1836);
nand U271 (N_271,In_1159,In_1662);
and U272 (N_272,In_1998,In_1877);
or U273 (N_273,In_52,In_1601);
nand U274 (N_274,In_2247,In_1774);
and U275 (N_275,In_807,In_305);
nand U276 (N_276,In_1301,In_835);
or U277 (N_277,In_2119,In_10);
nor U278 (N_278,In_1861,In_1337);
nor U279 (N_279,In_1062,In_382);
nand U280 (N_280,In_2468,In_1201);
nor U281 (N_281,In_572,In_553);
or U282 (N_282,In_481,In_1804);
nor U283 (N_283,In_2276,In_383);
or U284 (N_284,In_826,In_2007);
and U285 (N_285,In_1170,In_1090);
nand U286 (N_286,In_1646,In_523);
nand U287 (N_287,In_463,In_1433);
nor U288 (N_288,In_1479,In_246);
nand U289 (N_289,In_274,In_725);
nor U290 (N_290,In_2250,In_239);
nor U291 (N_291,In_737,In_1231);
nand U292 (N_292,In_167,In_1136);
nand U293 (N_293,In_2208,In_1913);
nand U294 (N_294,In_1275,In_1593);
and U295 (N_295,In_1113,In_1073);
nor U296 (N_296,In_971,In_163);
or U297 (N_297,In_1692,In_2118);
nor U298 (N_298,In_1925,In_1980);
and U299 (N_299,In_915,In_1724);
and U300 (N_300,In_797,In_1455);
or U301 (N_301,In_1562,In_1716);
nand U302 (N_302,In_2180,In_2407);
nand U303 (N_303,In_524,In_2200);
nor U304 (N_304,In_2262,In_2219);
or U305 (N_305,In_1407,In_492);
nand U306 (N_306,In_1779,In_434);
nor U307 (N_307,In_1228,In_1306);
nand U308 (N_308,In_1216,In_1522);
and U309 (N_309,In_1985,In_1675);
nand U310 (N_310,In_2462,In_2335);
and U311 (N_311,In_1894,In_116);
nor U312 (N_312,In_1227,In_337);
nor U313 (N_313,In_2075,In_31);
nand U314 (N_314,In_659,In_1670);
and U315 (N_315,In_2116,In_896);
and U316 (N_316,In_2470,In_2216);
nand U317 (N_317,In_2067,In_2389);
and U318 (N_318,In_2176,In_285);
nand U319 (N_319,In_1567,In_308);
nor U320 (N_320,In_2136,In_916);
nor U321 (N_321,In_2144,In_1537);
or U322 (N_322,In_1869,In_900);
and U323 (N_323,In_1308,In_507);
or U324 (N_324,In_1667,In_81);
xor U325 (N_325,In_155,In_2421);
or U326 (N_326,In_2082,In_1332);
nand U327 (N_327,In_1939,In_1866);
nand U328 (N_328,In_1671,In_398);
xor U329 (N_329,In_2002,In_1074);
nand U330 (N_330,In_942,In_392);
and U331 (N_331,In_1324,In_394);
and U332 (N_332,In_493,In_1684);
nand U333 (N_333,In_1128,In_2214);
or U334 (N_334,In_829,In_1251);
nor U335 (N_335,In_2370,In_615);
or U336 (N_336,In_27,In_854);
nand U337 (N_337,In_1630,In_1765);
nor U338 (N_338,In_304,In_2133);
or U339 (N_339,In_1619,In_2394);
and U340 (N_340,In_1849,In_2441);
nor U341 (N_341,In_1551,In_545);
nand U342 (N_342,In_60,In_2122);
nand U343 (N_343,In_1045,In_2454);
nor U344 (N_344,In_1647,In_751);
and U345 (N_345,In_1506,In_48);
and U346 (N_346,In_2459,In_2286);
nor U347 (N_347,In_1643,In_1135);
and U348 (N_348,In_18,In_1183);
nor U349 (N_349,In_2091,In_201);
and U350 (N_350,In_1773,In_1829);
nand U351 (N_351,In_475,In_1821);
nor U352 (N_352,In_338,In_490);
and U353 (N_353,In_1734,In_1457);
nand U354 (N_354,In_995,In_1888);
and U355 (N_355,In_1082,In_427);
and U356 (N_356,In_2320,In_773);
xor U357 (N_357,In_1526,In_696);
xnor U358 (N_358,In_358,In_301);
nand U359 (N_359,In_1451,In_319);
and U360 (N_360,In_761,In_263);
nor U361 (N_361,In_2260,In_1732);
nor U362 (N_362,In_1937,In_197);
or U363 (N_363,In_1564,In_957);
nor U364 (N_364,In_528,In_1037);
xor U365 (N_365,In_2209,In_1810);
nor U366 (N_366,In_2487,In_456);
or U367 (N_367,In_1500,In_2385);
nand U368 (N_368,In_271,In_2045);
and U369 (N_369,In_1195,In_1668);
nand U370 (N_370,In_2197,In_2240);
and U371 (N_371,In_1540,In_2329);
or U372 (N_372,In_1024,In_485);
xor U373 (N_373,In_1512,In_728);
nor U374 (N_374,In_2381,In_1490);
and U375 (N_375,In_335,In_603);
and U376 (N_376,In_1249,In_2070);
nor U377 (N_377,In_2281,In_886);
and U378 (N_378,In_828,In_500);
and U379 (N_379,In_1289,In_1477);
xor U380 (N_380,In_95,In_79);
xor U381 (N_381,In_1983,In_1932);
nor U382 (N_382,In_868,In_2037);
nor U383 (N_383,In_747,In_1509);
nand U384 (N_384,In_2048,In_2268);
nor U385 (N_385,In_1032,In_389);
or U386 (N_386,In_2173,In_952);
and U387 (N_387,In_1389,In_787);
nor U388 (N_388,In_2042,In_2342);
nor U389 (N_389,In_1304,In_1553);
or U390 (N_390,In_1377,In_757);
or U391 (N_391,In_1632,In_1578);
nand U392 (N_392,In_598,In_93);
nand U393 (N_393,In_1007,In_2392);
nor U394 (N_394,In_2210,In_2365);
nor U395 (N_395,In_1243,In_1393);
nor U396 (N_396,In_570,In_1502);
nand U397 (N_397,In_1175,In_632);
or U398 (N_398,In_213,In_1379);
and U399 (N_399,In_2316,In_1552);
nand U400 (N_400,In_1066,In_1012);
nand U401 (N_401,In_1368,In_1966);
and U402 (N_402,In_599,In_2096);
and U403 (N_403,In_1728,In_491);
nand U404 (N_404,In_1181,In_1060);
nand U405 (N_405,In_1936,In_540);
nor U406 (N_406,In_1962,In_1621);
nand U407 (N_407,In_2236,In_816);
nand U408 (N_408,In_635,In_1363);
or U409 (N_409,In_1239,In_1746);
nor U410 (N_410,In_2450,In_602);
or U411 (N_411,In_824,In_1528);
nand U412 (N_412,In_22,In_1669);
and U413 (N_413,In_1769,In_344);
nor U414 (N_414,In_140,In_419);
nor U415 (N_415,In_232,In_2348);
xor U416 (N_416,In_1252,In_1729);
nor U417 (N_417,In_71,In_2016);
nand U418 (N_418,In_117,In_126);
nor U419 (N_419,In_1122,In_65);
nor U420 (N_420,In_2390,In_1534);
and U421 (N_421,In_692,In_1504);
xnor U422 (N_422,In_2494,In_101);
nor U423 (N_423,In_1680,In_941);
nor U424 (N_424,In_2057,In_592);
nand U425 (N_425,In_2253,In_2298);
or U426 (N_426,In_1856,In_714);
or U427 (N_427,In_50,In_106);
nand U428 (N_428,In_1835,In_856);
or U429 (N_429,In_1666,In_2275);
nand U430 (N_430,In_587,In_391);
nand U431 (N_431,In_1860,In_2130);
nand U432 (N_432,In_1725,In_109);
nand U433 (N_433,In_591,In_1191);
and U434 (N_434,In_852,In_2429);
and U435 (N_435,In_59,In_1268);
and U436 (N_436,In_1523,In_934);
nor U437 (N_437,In_1213,In_864);
nor U438 (N_438,In_993,In_1419);
and U439 (N_439,In_2014,In_1198);
nor U440 (N_440,In_1445,In_802);
nand U441 (N_441,In_147,In_33);
nand U442 (N_442,In_1704,In_259);
nor U443 (N_443,In_90,In_2422);
nor U444 (N_444,In_279,In_499);
or U445 (N_445,In_1441,In_919);
or U446 (N_446,In_1319,In_1870);
or U447 (N_447,In_16,In_191);
nand U448 (N_448,In_1587,In_2324);
or U449 (N_449,In_166,In_2488);
and U450 (N_450,In_1194,In_497);
nand U451 (N_451,In_2148,In_9);
and U452 (N_452,In_918,In_2156);
and U453 (N_453,In_1350,In_1446);
and U454 (N_454,In_653,In_2444);
nand U455 (N_455,In_2372,In_2257);
nor U456 (N_456,In_1053,In_1690);
or U457 (N_457,In_365,In_1600);
and U458 (N_458,In_1283,In_775);
nand U459 (N_459,In_689,In_41);
nand U460 (N_460,In_111,In_1710);
and U461 (N_461,In_1339,In_1697);
and U462 (N_462,In_988,In_2289);
nand U463 (N_463,In_1395,In_1663);
nor U464 (N_464,In_462,In_1878);
nand U465 (N_465,In_914,In_2193);
nor U466 (N_466,In_534,In_715);
and U467 (N_467,In_1210,In_1398);
nand U468 (N_468,In_1815,In_1145);
nor U469 (N_469,In_2036,In_2222);
nor U470 (N_470,In_260,In_128);
and U471 (N_471,In_735,In_257);
or U472 (N_472,In_1467,In_1946);
nand U473 (N_473,In_564,In_823);
nand U474 (N_474,In_242,In_1672);
nand U475 (N_475,In_1855,In_1640);
nor U476 (N_476,In_1352,In_682);
or U477 (N_477,In_470,In_1944);
or U478 (N_478,In_1711,In_1876);
nor U479 (N_479,In_1730,In_1627);
nand U480 (N_480,In_1689,In_1687);
or U481 (N_481,In_2434,In_938);
nand U482 (N_482,In_35,In_1781);
and U483 (N_483,In_1846,In_1444);
nand U484 (N_484,In_1653,In_2399);
nand U485 (N_485,In_878,In_2147);
nand U486 (N_486,In_2230,In_5);
nor U487 (N_487,In_1278,In_1717);
nor U488 (N_488,In_1503,In_1387);
nor U489 (N_489,In_1212,In_1080);
or U490 (N_490,In_621,In_1462);
nor U491 (N_491,In_327,In_286);
xor U492 (N_492,In_1067,In_1456);
nor U493 (N_493,In_818,In_645);
and U494 (N_494,In_384,In_904);
or U495 (N_495,In_2228,In_2432);
or U496 (N_496,In_1637,In_1718);
nor U497 (N_497,In_313,In_1475);
nand U498 (N_498,In_237,In_1994);
or U499 (N_499,In_1465,In_2430);
or U500 (N_500,In_1485,In_208);
and U501 (N_501,In_1759,In_2443);
or U502 (N_502,In_1542,In_1209);
and U503 (N_503,In_2179,In_2080);
and U504 (N_504,In_1768,In_2218);
or U505 (N_505,In_2107,In_2081);
and U506 (N_506,In_1357,In_1154);
and U507 (N_507,In_626,In_53);
and U508 (N_508,In_1476,In_2287);
or U509 (N_509,In_314,In_1006);
and U510 (N_510,In_1556,In_1474);
and U511 (N_511,In_2124,In_850);
and U512 (N_512,In_2150,In_845);
and U513 (N_513,In_2331,In_366);
or U514 (N_514,In_533,In_898);
nand U515 (N_515,In_474,In_1150);
or U516 (N_516,In_193,In_1000);
and U517 (N_517,In_1918,In_766);
or U518 (N_518,In_393,In_316);
nor U519 (N_519,In_26,In_778);
nand U520 (N_520,In_2229,In_874);
or U521 (N_521,In_544,In_74);
xor U522 (N_522,In_1591,In_2325);
or U523 (N_523,In_297,In_2374);
and U524 (N_524,In_1226,In_1291);
or U525 (N_525,In_720,In_1580);
and U526 (N_526,In_1811,In_150);
and U527 (N_527,In_675,In_1427);
or U528 (N_528,In_1134,In_2383);
nand U529 (N_529,In_1148,In_1374);
xor U530 (N_530,In_461,In_1406);
or U531 (N_531,In_1075,In_672);
and U532 (N_532,In_17,In_2353);
and U533 (N_533,In_1650,In_1172);
nor U534 (N_534,In_1214,In_1492);
xnor U535 (N_535,In_374,In_1935);
or U536 (N_536,In_15,In_986);
or U537 (N_537,In_552,In_2069);
or U538 (N_538,In_1107,In_1606);
nand U539 (N_539,In_947,In_2347);
nand U540 (N_540,In_1900,In_299);
or U541 (N_541,In_2292,In_883);
nor U542 (N_542,In_334,In_1453);
nand U543 (N_543,In_2140,In_386);
or U544 (N_544,In_973,In_1187);
or U545 (N_545,In_983,In_2363);
nand U546 (N_546,In_627,In_1196);
and U547 (N_547,In_569,In_707);
nand U548 (N_548,In_262,In_1628);
or U549 (N_549,In_2023,In_1137);
or U550 (N_550,In_1346,In_1592);
nand U551 (N_551,In_2241,In_292);
nor U552 (N_552,In_2185,In_2296);
nand U553 (N_553,In_432,In_1284);
xnor U554 (N_554,In_457,In_1099);
and U555 (N_555,In_377,In_730);
nor U556 (N_556,In_2395,In_1276);
and U557 (N_557,In_2154,In_403);
and U558 (N_558,In_749,In_556);
and U559 (N_559,In_219,In_1616);
nor U560 (N_560,In_1312,In_1844);
nor U561 (N_561,In_2059,In_465);
xor U562 (N_562,In_685,In_1225);
nand U563 (N_563,In_300,In_1723);
nand U564 (N_564,In_800,In_767);
nand U565 (N_565,In_1051,In_373);
xor U566 (N_566,In_1354,In_625);
nor U567 (N_567,In_2034,In_1338);
and U568 (N_568,In_1220,In_1098);
nand U569 (N_569,In_2076,In_2481);
and U570 (N_570,In_1698,In_211);
nand U571 (N_571,In_1014,In_2251);
or U572 (N_572,In_238,In_2314);
or U573 (N_573,In_827,In_1382);
nor U574 (N_574,In_77,In_251);
xnor U575 (N_575,In_2155,In_1123);
nand U576 (N_576,In_858,In_1629);
and U577 (N_577,In_1545,In_2177);
nand U578 (N_578,In_2191,In_98);
nand U579 (N_579,In_1802,In_1155);
or U580 (N_580,In_1924,In_501);
or U581 (N_581,In_1997,In_476);
or U582 (N_582,In_795,In_2420);
nand U583 (N_583,In_1655,In_2238);
nand U584 (N_584,In_322,In_1536);
or U585 (N_585,In_1454,In_2332);
nand U586 (N_586,In_1532,In_508);
and U587 (N_587,In_899,In_2205);
or U588 (N_588,In_944,In_2088);
nor U589 (N_589,In_352,In_2138);
and U590 (N_590,In_181,In_882);
and U591 (N_591,In_859,In_891);
or U592 (N_592,In_149,In_2109);
or U593 (N_593,In_585,In_2378);
nor U594 (N_594,In_1748,In_968);
and U595 (N_595,In_162,In_2397);
or U596 (N_596,In_1050,In_2020);
xor U597 (N_597,In_1880,In_646);
xor U598 (N_598,In_2485,In_326);
nor U599 (N_599,In_2477,In_1356);
and U600 (N_600,In_2005,In_182);
nor U601 (N_601,In_1277,In_1950);
nand U602 (N_602,In_480,In_541);
nor U603 (N_603,In_2479,In_1179);
nor U604 (N_604,In_1920,In_1840);
nor U605 (N_605,In_2297,In_1422);
nor U606 (N_606,In_1141,In_1579);
nand U607 (N_607,In_1109,In_415);
or U608 (N_608,In_573,In_1739);
nor U609 (N_609,In_287,In_2452);
nand U610 (N_610,In_1140,In_1495);
nor U611 (N_611,In_152,In_1246);
nand U612 (N_612,In_1531,In_1555);
or U613 (N_613,In_113,In_1617);
or U614 (N_614,In_124,In_1906);
or U615 (N_615,In_1200,In_221);
and U616 (N_616,In_932,In_180);
nor U617 (N_617,In_192,In_2368);
nor U618 (N_618,In_1176,In_1158);
or U619 (N_619,In_494,In_1515);
nor U620 (N_620,In_1156,In_992);
and U621 (N_621,In_1525,In_67);
nor U622 (N_622,In_1569,In_516);
nand U623 (N_623,In_814,In_2497);
or U624 (N_624,In_342,In_1385);
or U625 (N_625,In_307,In_2317);
nand U626 (N_626,In_2293,In_1077);
nor U627 (N_627,In_69,In_847);
and U628 (N_628,In_789,In_911);
nand U629 (N_629,In_108,In_909);
or U630 (N_630,In_2457,In_2484);
and U631 (N_631,In_1756,In_897);
nand U632 (N_632,In_2182,In_1173);
nand U633 (N_633,In_928,In_2337);
or U634 (N_634,In_1042,In_756);
nor U635 (N_635,In_2196,In_590);
nand U636 (N_636,In_791,In_1349);
nor U637 (N_637,In_1803,In_1054);
and U638 (N_638,In_2001,In_1583);
nor U639 (N_639,In_1023,In_543);
or U640 (N_640,In_56,In_2382);
or U641 (N_641,In_907,In_1559);
or U642 (N_642,In_2125,In_1112);
nand U643 (N_643,In_638,In_803);
nand U644 (N_644,In_404,In_1776);
nand U645 (N_645,In_1421,In_965);
nand U646 (N_646,In_844,In_1926);
and U647 (N_647,In_679,In_479);
xor U648 (N_648,In_240,In_2233);
nor U649 (N_649,In_1891,In_935);
nor U650 (N_650,In_2158,In_2039);
nand U651 (N_651,In_894,In_1199);
or U652 (N_652,In_1321,In_1596);
nand U653 (N_653,In_801,In_1720);
nand U654 (N_654,In_661,In_1881);
nand U655 (N_655,In_2451,In_2418);
nand U656 (N_656,In_1164,In_431);
or U657 (N_657,In_1040,In_252);
xor U658 (N_658,In_2004,In_32);
or U659 (N_659,In_88,In_1254);
xor U660 (N_660,In_946,In_2428);
nor U661 (N_661,In_1707,In_68);
and U662 (N_662,In_571,In_703);
nand U663 (N_663,In_1430,In_448);
nand U664 (N_664,In_2384,In_171);
nand U665 (N_665,In_1987,In_1737);
and U666 (N_666,In_1169,In_1088);
or U667 (N_667,In_30,In_2306);
or U668 (N_668,In_1376,In_1615);
nand U669 (N_669,In_1991,In_595);
or U670 (N_670,In_363,In_2227);
or U671 (N_671,In_974,In_2141);
nand U672 (N_672,In_782,In_650);
nand U673 (N_673,In_1948,In_1921);
and U674 (N_674,In_1703,In_84);
or U675 (N_675,In_1989,In_1317);
or U676 (N_676,In_1424,In_831);
and U677 (N_677,In_1459,In_2448);
nand U678 (N_678,In_640,In_1986);
and U679 (N_679,In_1851,In_2068);
nor U680 (N_680,In_158,In_134);
nor U681 (N_681,In_1816,In_2423);
and U682 (N_682,In_560,In_2356);
or U683 (N_683,In_1763,In_2090);
nor U684 (N_684,In_1677,In_1995);
or U685 (N_685,In_1244,In_303);
nand U686 (N_686,In_295,In_1828);
and U687 (N_687,In_2290,In_2414);
and U688 (N_688,In_1413,In_336);
and U689 (N_689,In_453,In_641);
and U690 (N_690,In_1882,In_1002);
and U691 (N_691,In_998,In_2032);
and U692 (N_692,In_1722,In_2346);
or U693 (N_693,In_1801,In_2194);
or U694 (N_694,In_1893,In_2266);
nor U695 (N_695,In_1772,In_1353);
nand U696 (N_696,In_174,In_1336);
and U697 (N_697,In_255,In_1678);
nand U698 (N_698,In_548,In_2095);
nor U699 (N_699,In_2212,In_1005);
or U700 (N_700,In_1458,In_657);
nand U701 (N_701,In_1839,In_2153);
nand U702 (N_702,In_102,In_1612);
or U703 (N_703,In_100,In_447);
nor U704 (N_704,In_905,In_1203);
or U705 (N_705,In_233,In_1373);
and U706 (N_706,In_1464,In_2396);
nor U707 (N_707,In_813,In_115);
or U708 (N_708,In_639,In_1614);
and U709 (N_709,In_997,In_315);
nor U710 (N_710,In_1131,In_2110);
nor U711 (N_711,In_651,In_970);
nor U712 (N_712,In_498,In_471);
nand U713 (N_713,In_1794,In_2489);
or U714 (N_714,In_1245,In_1144);
and U715 (N_715,In_267,In_667);
or U716 (N_716,In_1394,In_1626);
or U717 (N_717,In_1423,In_554);
or U718 (N_718,In_1038,In_1415);
or U719 (N_719,In_2486,In_1084);
and U720 (N_720,In_1903,In_131);
and U721 (N_721,In_2149,In_1114);
and U722 (N_722,In_1035,In_1401);
nor U723 (N_723,In_364,In_346);
and U724 (N_724,In_2128,In_1604);
xnor U725 (N_725,In_1068,In_1990);
or U726 (N_726,In_593,In_1996);
nand U727 (N_727,In_1287,In_289);
nor U728 (N_728,In_1691,In_810);
and U729 (N_729,In_517,In_576);
nand U730 (N_730,In_1065,In_1549);
nand U731 (N_731,In_1411,In_473);
and U732 (N_732,In_1709,In_47);
and U733 (N_733,In_380,In_808);
or U734 (N_734,In_265,In_1019);
nand U735 (N_735,In_189,In_1783);
nor U736 (N_736,In_1327,In_28);
or U737 (N_737,In_1822,In_1463);
and U738 (N_738,In_1229,In_607);
or U739 (N_739,In_199,In_1013);
nor U740 (N_740,In_1510,In_321);
nand U741 (N_741,In_400,In_2164);
nor U742 (N_742,In_406,In_1890);
xor U743 (N_743,In_1577,In_933);
and U744 (N_744,In_2367,In_55);
nor U745 (N_745,In_1897,In_156);
nand U746 (N_746,In_44,In_1817);
nor U747 (N_747,In_924,In_2366);
nand U748 (N_748,In_24,In_1605);
nor U749 (N_749,In_435,In_139);
nand U750 (N_750,In_849,In_662);
and U751 (N_751,In_798,In_780);
or U752 (N_752,In_2278,In_1305);
and U753 (N_753,In_1063,In_1361);
and U754 (N_754,In_1333,In_694);
or U755 (N_755,In_13,In_1872);
nor U756 (N_756,In_1685,In_2254);
or U757 (N_757,In_2388,In_1750);
and U758 (N_758,In_1028,In_1025);
nor U759 (N_759,In_860,In_1120);
nand U760 (N_760,In_348,In_356);
nor U761 (N_761,In_1530,In_7);
or U762 (N_762,In_709,In_215);
or U763 (N_763,In_1644,In_1372);
nor U764 (N_764,In_1309,In_1106);
nor U765 (N_765,In_881,In_446);
and U766 (N_766,In_2000,In_1741);
xnor U767 (N_767,In_1743,In_368);
nor U768 (N_768,In_2162,In_114);
xor U769 (N_769,In_34,In_311);
nand U770 (N_770,In_1087,In_1742);
and U771 (N_771,In_1493,In_129);
and U772 (N_772,In_721,In_1943);
nor U773 (N_773,In_1819,In_976);
nor U774 (N_774,In_1402,In_619);
and U775 (N_775,In_1883,In_75);
nor U776 (N_776,In_504,In_1895);
nor U777 (N_777,In_1081,In_843);
or U778 (N_778,In_2498,In_520);
or U779 (N_779,In_1818,In_1665);
or U780 (N_780,In_2309,In_2132);
or U781 (N_781,In_226,In_1072);
nor U782 (N_782,In_296,In_1091);
nor U783 (N_783,In_1089,In_1884);
nor U784 (N_784,In_1020,In_670);
nand U785 (N_785,In_2019,In_455);
or U786 (N_786,In_611,In_2400);
and U787 (N_787,In_2204,In_2471);
and U788 (N_788,In_1543,In_216);
or U789 (N_789,In_0,In_642);
xnor U790 (N_790,In_568,In_332);
or U791 (N_791,In_885,In_1438);
nor U792 (N_792,In_2221,In_796);
xor U793 (N_793,In_1362,In_812);
and U794 (N_794,In_355,In_1142);
nand U795 (N_795,In_799,In_1570);
or U796 (N_796,In_2040,In_145);
and U797 (N_797,In_266,In_170);
nand U798 (N_798,In_1548,In_1211);
nand U799 (N_799,In_1293,In_600);
nand U800 (N_800,In_1800,In_1520);
nand U801 (N_801,In_46,In_817);
xor U802 (N_802,In_962,In_440);
nand U803 (N_803,In_987,In_1396);
or U804 (N_804,In_2272,In_557);
or U805 (N_805,In_2282,In_1335);
nor U806 (N_806,In_1778,In_1094);
or U807 (N_807,In_991,In_1253);
nand U808 (N_808,In_2495,In_2305);
nand U809 (N_809,In_2224,In_1412);
or U810 (N_810,In_1963,In_1806);
or U811 (N_811,In_2199,In_1648);
and U812 (N_812,In_1297,In_959);
nor U813 (N_813,In_66,In_1341);
and U814 (N_814,In_2435,In_323);
nand U815 (N_815,In_220,In_702);
and U816 (N_816,In_1956,In_354);
and U817 (N_817,In_430,In_1184);
or U818 (N_818,In_1496,In_2114);
and U819 (N_819,In_1889,In_655);
and U820 (N_820,In_562,In_1832);
or U821 (N_821,In_1100,In_1439);
and U822 (N_822,In_1409,In_1294);
nand U823 (N_823,In_2062,In_855);
nand U824 (N_824,In_871,In_734);
and U825 (N_825,In_2273,In_2011);
nand U826 (N_826,In_2105,In_417);
nand U827 (N_827,In_1571,In_1127);
nand U828 (N_828,In_1568,In_1180);
nor U829 (N_829,In_2100,In_1557);
nor U830 (N_830,In_2362,In_1208);
nor U831 (N_831,In_2352,In_920);
nor U832 (N_832,In_2093,In_2046);
or U833 (N_833,In_2195,In_1952);
nor U834 (N_834,In_269,In_1217);
or U835 (N_835,In_1623,In_1747);
nor U836 (N_836,In_1598,In_40);
and U837 (N_837,In_2043,In_2052);
nor U838 (N_838,In_2047,In_184);
nand U839 (N_839,In_318,In_1101);
and U840 (N_840,In_2351,In_700);
or U841 (N_841,In_175,In_704);
or U842 (N_842,In_1383,In_723);
nor U843 (N_843,In_2405,In_930);
nand U844 (N_844,In_408,In_1428);
and U845 (N_845,In_2349,In_76);
and U846 (N_846,In_1130,In_1189);
nor U847 (N_847,In_837,In_2157);
nand U848 (N_848,In_774,In_2343);
nor U849 (N_849,In_146,In_1328);
or U850 (N_850,In_1791,In_187);
nor U851 (N_851,In_2493,In_478);
or U852 (N_852,In_2056,In_604);
nand U853 (N_853,In_764,In_375);
nand U854 (N_854,In_422,In_776);
or U855 (N_855,In_2097,In_458);
nand U856 (N_856,In_2131,In_227);
and U857 (N_857,In_819,In_1755);
or U858 (N_858,In_726,In_2327);
nor U859 (N_859,In_2021,In_701);
and U860 (N_860,In_1879,In_2079);
nor U861 (N_861,In_1139,In_1885);
nand U862 (N_862,In_1118,In_2249);
and U863 (N_863,In_1404,In_1535);
nor U864 (N_864,In_185,In_1658);
and U865 (N_865,In_668,In_1391);
nand U866 (N_866,In_1908,In_2252);
nand U867 (N_867,In_1929,In_1151);
or U868 (N_868,In_1507,In_1001);
xnor U869 (N_869,In_2145,In_1777);
xnor U870 (N_870,In_99,In_2280);
and U871 (N_871,In_1468,In_2055);
nor U872 (N_872,In_1787,In_2354);
nand U873 (N_873,In_923,In_2234);
or U874 (N_874,In_536,In_762);
or U875 (N_875,In_121,In_317);
nor U876 (N_876,In_379,In_1634);
and U877 (N_877,In_1886,In_2274);
and U878 (N_878,In_1489,In_421);
and U879 (N_879,In_746,In_1857);
and U880 (N_880,In_1310,In_2165);
or U881 (N_881,In_1554,In_1364);
or U882 (N_882,In_1796,In_1110);
nor U883 (N_883,In_1070,In_1274);
nand U884 (N_884,In_1236,In_529);
xor U885 (N_885,In_1702,In_744);
nor U886 (N_886,In_62,In_401);
nor U887 (N_887,In_157,In_2071);
or U888 (N_888,In_2015,In_204);
and U889 (N_889,In_1922,In_1442);
or U890 (N_890,In_1518,In_1812);
nor U891 (N_891,In_63,In_122);
nor U892 (N_892,In_1585,In_488);
and U893 (N_893,In_729,In_1034);
and U894 (N_894,In_1706,In_1602);
nand U895 (N_895,In_2338,In_2123);
nand U896 (N_896,In_794,In_981);
nor U897 (N_897,In_1331,In_990);
or U898 (N_898,In_724,In_2344);
xor U899 (N_899,In_1288,In_1958);
nor U900 (N_900,In_2466,In_996);
nand U901 (N_901,In_2270,In_1673);
nor U902 (N_902,In_708,In_1392);
nand U903 (N_903,In_1133,In_1039);
nor U904 (N_904,In_1499,In_169);
or U905 (N_905,In_1688,In_1940);
or U906 (N_906,In_1597,In_1061);
and U907 (N_907,In_722,In_1862);
nand U908 (N_908,In_1472,In_290);
nand U909 (N_909,In_1115,In_118);
and U910 (N_910,In_967,In_1736);
and U911 (N_911,In_2078,In_582);
or U912 (N_912,In_1992,In_2350);
nand U913 (N_913,In_1484,In_1726);
nand U914 (N_914,In_1386,In_12);
nand U915 (N_915,In_1674,In_1625);
nand U916 (N_916,In_503,In_1182);
or U917 (N_917,In_763,In_411);
nor U918 (N_918,In_2101,In_429);
or U919 (N_919,In_2190,In_777);
nand U920 (N_920,In_45,In_1009);
nor U921 (N_921,In_110,In_727);
nand U922 (N_922,In_1033,In_20);
nand U923 (N_923,In_29,In_2168);
and U924 (N_924,In_1766,In_1247);
and U925 (N_925,In_502,In_2340);
and U926 (N_926,In_186,In_1168);
nor U927 (N_927,In_1461,In_1126);
nand U928 (N_928,In_581,In_1011);
and U929 (N_929,In_1708,In_1206);
and U930 (N_930,In_177,In_1770);
nor U931 (N_931,In_2371,In_889);
nand U932 (N_932,In_1345,In_172);
or U933 (N_933,In_612,In_2285);
and U934 (N_934,In_1259,In_1785);
and U935 (N_935,In_2142,In_178);
xor U936 (N_936,In_2174,In_1347);
or U937 (N_937,In_2339,In_1941);
nor U938 (N_938,In_1471,In_1138);
nand U939 (N_939,In_752,In_1915);
nor U940 (N_940,In_822,In_666);
and U941 (N_941,In_495,In_1902);
or U942 (N_942,In_1437,In_11);
nand U943 (N_943,In_1286,In_357);
nand U944 (N_944,In_1654,In_1563);
nor U945 (N_945,In_256,In_820);
xnor U946 (N_946,In_2166,In_2465);
nand U947 (N_947,In_1969,In_2453);
nor U948 (N_948,In_2248,In_978);
nor U949 (N_949,In_1834,In_272);
and U950 (N_950,In_964,In_1280);
or U951 (N_951,In_2074,In_869);
nand U952 (N_952,In_235,In_1344);
and U953 (N_953,In_1497,In_677);
or U954 (N_954,In_956,In_467);
or U955 (N_955,In_2271,In_341);
and U956 (N_956,In_1026,In_420);
nand U957 (N_957,In_1745,In_1163);
nor U958 (N_958,In_1384,In_2031);
nand U959 (N_959,In_2025,In_788);
nand U960 (N_960,In_328,In_1988);
nand U961 (N_961,In_91,In_566);
and U962 (N_962,In_2022,In_793);
nand U963 (N_963,In_2033,In_320);
or U964 (N_964,In_441,In_1486);
or U965 (N_965,In_142,In_769);
nor U966 (N_966,In_512,In_1854);
nor U967 (N_967,In_2178,In_2379);
or U968 (N_968,In_937,In_2064);
and U969 (N_969,In_522,In_214);
nand U970 (N_970,In_2115,In_1705);
nand U971 (N_971,In_1234,In_880);
nor U972 (N_972,In_678,In_1417);
nand U973 (N_973,In_1657,In_940);
or U974 (N_974,In_1272,In_8);
nand U975 (N_975,In_2279,In_2406);
nor U976 (N_976,In_2006,In_574);
or U977 (N_977,In_1576,In_2027);
nor U978 (N_978,In_2188,In_2461);
nand U979 (N_979,In_1947,In_1481);
nor U980 (N_980,In_1786,In_1539);
nor U981 (N_981,In_785,In_2330);
nand U982 (N_982,In_1713,In_628);
nand U983 (N_983,In_535,In_1360);
nor U984 (N_984,In_2483,In_578);
nor U985 (N_985,In_2201,In_1975);
or U986 (N_986,In_424,In_1799);
nand U987 (N_987,In_1949,In_2102);
and U988 (N_988,In_906,In_955);
and U989 (N_989,In_361,In_2267);
nand U990 (N_990,In_2167,In_665);
or U991 (N_991,In_2478,In_1871);
and U992 (N_992,In_372,In_1);
and U993 (N_993,In_2084,In_954);
nor U994 (N_994,In_261,In_519);
nand U995 (N_995,In_127,In_1859);
and U996 (N_996,In_2480,In_2215);
and U997 (N_997,In_1355,In_1945);
nor U998 (N_998,In_1508,In_469);
xnor U999 (N_999,In_917,In_1108);
nor U1000 (N_1000,In_2376,In_1111);
and U1001 (N_1001,In_443,In_876);
and U1002 (N_1002,In_1686,In_1917);
nand U1003 (N_1003,In_1320,In_310);
xnor U1004 (N_1004,In_2112,In_521);
or U1005 (N_1005,In_410,In_1414);
or U1006 (N_1006,In_1097,In_2243);
nand U1007 (N_1007,In_1792,In_345);
and U1008 (N_1008,In_2085,In_2192);
and U1009 (N_1009,In_2187,In_1436);
or U1010 (N_1010,In_351,In_1978);
and U1011 (N_1011,In_2003,In_1095);
or U1012 (N_1012,In_2440,In_360);
nor U1013 (N_1013,In_2301,In_617);
nor U1014 (N_1014,In_2412,In_1904);
or U1015 (N_1015,In_218,In_719);
or U1016 (N_1016,In_1761,In_1399);
nand U1017 (N_1017,In_293,In_1622);
or U1018 (N_1018,In_460,In_51);
and U1019 (N_1019,In_2121,In_83);
nand U1020 (N_1020,In_594,In_1901);
and U1021 (N_1021,In_1197,In_104);
or U1022 (N_1022,In_1027,In_1964);
and U1023 (N_1023,In_1017,In_839);
and U1024 (N_1024,In_176,In_2172);
and U1025 (N_1025,In_711,In_683);
nor U1026 (N_1026,In_195,In_652);
and U1027 (N_1027,In_1124,In_2308);
and U1028 (N_1028,In_1538,In_143);
and U1029 (N_1029,In_325,In_2028);
or U1030 (N_1030,In_1809,In_1429);
nand U1031 (N_1031,In_842,In_1270);
nand U1032 (N_1032,In_712,In_1105);
nor U1033 (N_1033,In_781,In_825);
or U1034 (N_1034,In_1652,In_1916);
nand U1035 (N_1035,In_1588,In_1524);
nor U1036 (N_1036,In_2345,In_2066);
and U1037 (N_1037,In_732,In_515);
and U1038 (N_1038,In_1031,In_2030);
nand U1039 (N_1039,In_2311,In_103);
and U1040 (N_1040,In_329,In_663);
and U1041 (N_1041,In_1185,In_2083);
or U1042 (N_1042,In_606,In_205);
or U1043 (N_1043,In_1981,In_551);
nor U1044 (N_1044,In_877,In_1292);
or U1045 (N_1045,In_559,In_2051);
nand U1046 (N_1046,In_388,In_1613);
nand U1047 (N_1047,In_459,In_1460);
and U1048 (N_1048,In_1367,In_884);
nor U1049 (N_1049,In_1119,In_2436);
and U1050 (N_1050,In_1340,In_509);
or U1051 (N_1051,In_676,In_1315);
nor U1052 (N_1052,In_753,In_2258);
or U1053 (N_1053,In_1642,In_1046);
and U1054 (N_1054,In_1603,In_378);
or U1055 (N_1055,In_1222,In_948);
xor U1056 (N_1056,In_2063,In_538);
or U1057 (N_1057,In_1760,In_921);
nor U1058 (N_1058,In_349,In_439);
nor U1059 (N_1059,In_2472,In_1911);
nor U1060 (N_1060,In_1147,In_731);
xor U1061 (N_1061,In_2496,In_806);
nand U1062 (N_1062,In_444,In_387);
nand U1063 (N_1063,In_705,In_768);
nand U1064 (N_1064,In_1403,In_979);
or U1065 (N_1065,In_2072,In_1589);
nand U1066 (N_1066,In_1965,In_1313);
nor U1067 (N_1067,In_1923,In_1318);
nor U1068 (N_1068,In_2302,In_1314);
or U1069 (N_1069,In_1636,In_1266);
nand U1070 (N_1070,In_2220,In_1044);
and U1071 (N_1071,In_2255,In_135);
and U1072 (N_1072,In_258,In_2312);
nor U1073 (N_1073,In_1425,In_580);
and U1074 (N_1074,In_539,In_1221);
or U1075 (N_1075,In_2038,In_428);
or U1076 (N_1076,In_1230,In_1397);
nor U1077 (N_1077,In_1993,In_1681);
and U1078 (N_1078,In_1907,In_1875);
nand U1079 (N_1079,In_153,In_1450);
nor U1080 (N_1080,In_309,In_838);
and U1081 (N_1081,In_1740,In_241);
or U1082 (N_1082,In_1753,In_586);
nor U1083 (N_1083,In_892,In_141);
nand U1084 (N_1084,In_1874,In_1494);
nand U1085 (N_1085,In_2403,In_648);
nor U1086 (N_1086,In_288,In_1478);
and U1087 (N_1087,In_532,In_376);
and U1088 (N_1088,In_1469,In_1971);
and U1089 (N_1089,In_1435,In_698);
nand U1090 (N_1090,In_1898,In_2073);
nand U1091 (N_1091,In_324,In_2294);
nand U1092 (N_1092,In_736,In_577);
and U1093 (N_1093,In_1359,In_1967);
or U1094 (N_1094,In_2242,In_1825);
nand U1095 (N_1095,In_903,In_2303);
or U1096 (N_1096,In_1757,In_2213);
or U1097 (N_1097,In_821,In_61);
or U1098 (N_1098,In_1440,In_281);
and U1099 (N_1099,In_1599,In_1608);
and U1100 (N_1100,In_2111,In_922);
nor U1101 (N_1101,In_1302,In_620);
and U1102 (N_1102,In_2413,In_1695);
nand U1103 (N_1103,In_396,In_1764);
nor U1104 (N_1104,In_2018,In_1784);
and U1105 (N_1105,In_902,In_1931);
nor U1106 (N_1106,In_2099,In_2202);
or U1107 (N_1107,In_513,In_107);
nand U1108 (N_1108,In_425,In_1738);
nor U1109 (N_1109,In_1572,In_229);
or U1110 (N_1110,In_1296,In_1808);
nor U1111 (N_1111,In_486,In_412);
and U1112 (N_1112,In_2426,In_717);
and U1113 (N_1113,In_931,In_254);
nor U1114 (N_1114,In_1057,In_1047);
nand U1115 (N_1115,In_526,In_2417);
xor U1116 (N_1116,In_339,In_80);
or U1117 (N_1117,In_710,In_1449);
or U1118 (N_1118,In_975,In_1586);
nand U1119 (N_1119,In_477,In_1609);
nor U1120 (N_1120,In_395,In_4);
nor U1121 (N_1121,In_200,In_1959);
nand U1122 (N_1122,In_450,In_132);
and U1123 (N_1123,In_558,In_1899);
nand U1124 (N_1124,In_2245,In_1727);
nand U1125 (N_1125,In_2256,In_1022);
or U1126 (N_1126,In_202,In_2377);
or U1127 (N_1127,In_1400,In_875);
or U1128 (N_1128,In_203,In_656);
and U1129 (N_1129,In_1408,In_6);
and U1130 (N_1130,In_2410,In_684);
and U1131 (N_1131,In_2223,In_862);
and U1132 (N_1132,In_687,In_1909);
nand U1133 (N_1133,In_644,In_1041);
nand U1134 (N_1134,In_575,In_2151);
or U1135 (N_1135,In_306,In_72);
nor U1136 (N_1136,In_2169,In_1977);
or U1137 (N_1137,In_1330,In_771);
nand U1138 (N_1138,In_669,In_583);
nor U1139 (N_1139,In_119,In_555);
and U1140 (N_1140,In_1719,In_1048);
and U1141 (N_1141,In_436,In_38);
and U1142 (N_1142,In_609,In_804);
and U1143 (N_1143,In_951,In_1798);
nor U1144 (N_1144,In_1498,In_2013);
or U1145 (N_1145,In_1752,In_2416);
nand U1146 (N_1146,In_913,In_1117);
nand U1147 (N_1147,In_1432,In_209);
nand U1148 (N_1148,In_1237,In_1651);
nor U1149 (N_1149,In_2404,In_1079);
nor U1150 (N_1150,In_1093,In_78);
or U1151 (N_1151,In_57,In_963);
and U1152 (N_1152,In_929,In_1649);
nand U1153 (N_1153,In_945,In_1633);
nor U1154 (N_1154,In_1848,In_770);
or U1155 (N_1155,In_745,In_1059);
nand U1156 (N_1156,In_961,In_302);
and U1157 (N_1157,In_2359,In_2408);
nor U1158 (N_1158,In_2419,In_1694);
and U1159 (N_1159,In_1388,In_1273);
nor U1160 (N_1160,In_2113,In_1841);
nand U1161 (N_1161,In_2010,In_2127);
nor U1162 (N_1162,In_1984,In_1896);
or U1163 (N_1163,In_2467,In_527);
or U1164 (N_1164,In_999,In_445);
or U1165 (N_1165,In_2358,In_1541);
nor U1166 (N_1166,In_1202,In_1279);
and U1167 (N_1167,In_1261,In_212);
or U1168 (N_1168,In_836,In_1715);
nand U1169 (N_1169,In_629,In_2077);
or U1170 (N_1170,In_144,In_2049);
nand U1171 (N_1171,In_2364,In_1049);
nand U1172 (N_1172,In_1762,In_418);
and U1173 (N_1173,In_161,In_865);
and U1174 (N_1174,In_2161,In_1205);
and U1175 (N_1175,In_1311,In_2008);
or U1176 (N_1176,In_1676,In_223);
or U1177 (N_1177,In_833,In_716);
nand U1178 (N_1178,In_972,In_2226);
and U1179 (N_1179,In_1258,In_1645);
nor U1180 (N_1180,In_222,In_14);
nor U1181 (N_1181,In_3,In_1767);
xnor U1182 (N_1182,In_1102,In_1351);
nor U1183 (N_1183,In_2460,In_1152);
nand U1184 (N_1184,In_616,In_1103);
or U1185 (N_1185,In_2104,In_1863);
nand U1186 (N_1186,In_1250,In_2139);
and U1187 (N_1187,In_1071,In_697);
nor U1188 (N_1188,In_343,In_1954);
and U1189 (N_1189,In_834,In_451);
or U1190 (N_1190,In_1867,In_1186);
or U1191 (N_1191,In_2491,In_2092);
or U1192 (N_1192,In_2449,In_87);
and U1193 (N_1193,In_741,In_1558);
or U1194 (N_1194,In_228,In_244);
nor U1195 (N_1195,In_1256,In_253);
and U1196 (N_1196,In_1933,In_1581);
nand U1197 (N_1197,In_1452,In_2232);
nand U1198 (N_1198,In_2146,In_2427);
nand U1199 (N_1199,In_1129,In_231);
nor U1200 (N_1200,In_496,In_210);
and U1201 (N_1201,In_518,In_437);
and U1202 (N_1202,In_39,In_82);
nor U1203 (N_1203,In_605,In_853);
nand U1204 (N_1204,In_660,In_1970);
and U1205 (N_1205,In_713,In_505);
and U1206 (N_1206,In_2315,In_2318);
or U1207 (N_1207,In_2026,In_1491);
or U1208 (N_1208,In_1961,In_64);
and U1209 (N_1209,In_133,In_234);
or U1210 (N_1210,In_943,In_416);
xor U1211 (N_1211,In_1560,In_1248);
and U1212 (N_1212,In_2284,In_531);
and U1213 (N_1213,In_863,In_537);
nor U1214 (N_1214,In_2458,In_1865);
and U1215 (N_1215,In_2246,In_1487);
or U1216 (N_1216,In_433,In_2269);
or U1217 (N_1217,In_1683,In_830);
and U1218 (N_1218,In_958,In_631);
and U1219 (N_1219,In_165,In_1325);
and U1220 (N_1220,In_2126,In_2143);
nand U1221 (N_1221,In_2186,In_468);
and U1222 (N_1222,In_815,In_236);
nand U1223 (N_1223,In_333,In_2474);
nand U1224 (N_1224,In_1016,In_1823);
nand U1225 (N_1225,In_1018,In_2473);
and U1226 (N_1226,In_466,In_1827);
nand U1227 (N_1227,In_123,In_54);
nand U1228 (N_1228,In_2375,In_483);
nor U1229 (N_1229,In_1300,In_2401);
nand U1230 (N_1230,In_1029,In_2307);
and U1231 (N_1231,In_634,In_2134);
and U1232 (N_1232,In_2380,In_565);
nand U1233 (N_1233,In_276,In_2415);
or U1234 (N_1234,In_1378,In_1751);
nor U1235 (N_1235,In_250,In_442);
and U1236 (N_1236,In_58,In_550);
nand U1237 (N_1237,In_936,In_409);
nor U1238 (N_1238,In_910,In_908);
nor U1239 (N_1239,In_2137,In_1443);
or U1240 (N_1240,In_1329,In_1789);
and U1241 (N_1241,In_2065,In_1326);
or U1242 (N_1242,In_2442,In_547);
and U1243 (N_1243,In_1483,In_1887);
nor U1244 (N_1244,In_284,In_2184);
nor U1245 (N_1245,In_1864,In_2323);
or U1246 (N_1246,In_2207,In_245);
nor U1247 (N_1247,In_452,In_249);
nand U1248 (N_1248,In_2446,In_546);
and U1249 (N_1249,In_154,In_2321);
xnor U1250 (N_1250,In_1874,In_1651);
nand U1251 (N_1251,In_1474,In_1837);
nor U1252 (N_1252,In_1449,In_1806);
or U1253 (N_1253,In_708,In_613);
and U1254 (N_1254,In_2023,In_2261);
and U1255 (N_1255,In_1379,In_1921);
and U1256 (N_1256,In_731,In_677);
xor U1257 (N_1257,In_1663,In_1304);
nor U1258 (N_1258,In_480,In_1458);
or U1259 (N_1259,In_1902,In_225);
nor U1260 (N_1260,In_1412,In_1136);
and U1261 (N_1261,In_2415,In_2095);
xnor U1262 (N_1262,In_617,In_108);
nor U1263 (N_1263,In_1011,In_1523);
nand U1264 (N_1264,In_167,In_2063);
and U1265 (N_1265,In_109,In_1968);
and U1266 (N_1266,In_1067,In_130);
and U1267 (N_1267,In_423,In_2021);
nand U1268 (N_1268,In_444,In_1929);
and U1269 (N_1269,In_1438,In_1252);
and U1270 (N_1270,In_2202,In_1605);
nor U1271 (N_1271,In_810,In_623);
nand U1272 (N_1272,In_594,In_1764);
or U1273 (N_1273,In_1827,In_200);
nand U1274 (N_1274,In_90,In_1088);
nor U1275 (N_1275,In_1395,In_2336);
or U1276 (N_1276,In_2233,In_1264);
nand U1277 (N_1277,In_38,In_487);
or U1278 (N_1278,In_735,In_439);
nor U1279 (N_1279,In_1731,In_215);
nor U1280 (N_1280,In_945,In_644);
or U1281 (N_1281,In_1711,In_1942);
or U1282 (N_1282,In_1216,In_1660);
xnor U1283 (N_1283,In_1019,In_2247);
and U1284 (N_1284,In_722,In_202);
nor U1285 (N_1285,In_432,In_1208);
nor U1286 (N_1286,In_2491,In_2043);
and U1287 (N_1287,In_1503,In_2111);
nor U1288 (N_1288,In_1490,In_286);
nand U1289 (N_1289,In_1161,In_1669);
or U1290 (N_1290,In_1777,In_2380);
nand U1291 (N_1291,In_2212,In_491);
or U1292 (N_1292,In_2104,In_1624);
nand U1293 (N_1293,In_71,In_219);
or U1294 (N_1294,In_258,In_881);
and U1295 (N_1295,In_2058,In_1173);
and U1296 (N_1296,In_31,In_915);
or U1297 (N_1297,In_1148,In_1581);
nor U1298 (N_1298,In_1104,In_1345);
nor U1299 (N_1299,In_2304,In_1062);
nand U1300 (N_1300,In_1642,In_1728);
and U1301 (N_1301,In_1495,In_989);
and U1302 (N_1302,In_1096,In_1034);
and U1303 (N_1303,In_856,In_1683);
nand U1304 (N_1304,In_2236,In_1175);
or U1305 (N_1305,In_562,In_158);
xor U1306 (N_1306,In_645,In_2428);
xnor U1307 (N_1307,In_578,In_332);
or U1308 (N_1308,In_2334,In_938);
and U1309 (N_1309,In_311,In_2365);
and U1310 (N_1310,In_1743,In_1101);
or U1311 (N_1311,In_859,In_2485);
or U1312 (N_1312,In_866,In_1044);
or U1313 (N_1313,In_2464,In_1135);
xnor U1314 (N_1314,In_2243,In_369);
nand U1315 (N_1315,In_2276,In_459);
and U1316 (N_1316,In_14,In_432);
and U1317 (N_1317,In_813,In_1186);
nor U1318 (N_1318,In_1223,In_1709);
and U1319 (N_1319,In_44,In_2083);
nand U1320 (N_1320,In_624,In_1767);
nand U1321 (N_1321,In_2192,In_308);
and U1322 (N_1322,In_950,In_2066);
and U1323 (N_1323,In_542,In_301);
and U1324 (N_1324,In_1627,In_94);
xor U1325 (N_1325,In_2257,In_1101);
and U1326 (N_1326,In_1572,In_62);
or U1327 (N_1327,In_731,In_564);
nand U1328 (N_1328,In_1702,In_635);
nand U1329 (N_1329,In_773,In_1804);
nor U1330 (N_1330,In_2413,In_640);
or U1331 (N_1331,In_980,In_2185);
and U1332 (N_1332,In_897,In_1319);
nor U1333 (N_1333,In_711,In_685);
and U1334 (N_1334,In_1473,In_2435);
or U1335 (N_1335,In_2065,In_673);
nor U1336 (N_1336,In_1504,In_1204);
or U1337 (N_1337,In_2290,In_305);
and U1338 (N_1338,In_513,In_2443);
and U1339 (N_1339,In_2405,In_646);
nand U1340 (N_1340,In_1445,In_1047);
or U1341 (N_1341,In_1714,In_526);
nand U1342 (N_1342,In_774,In_1513);
nand U1343 (N_1343,In_1335,In_676);
nor U1344 (N_1344,In_937,In_1056);
nand U1345 (N_1345,In_1958,In_866);
nor U1346 (N_1346,In_1042,In_498);
nor U1347 (N_1347,In_1339,In_693);
or U1348 (N_1348,In_1598,In_336);
or U1349 (N_1349,In_2115,In_916);
nor U1350 (N_1350,In_881,In_1307);
nor U1351 (N_1351,In_122,In_1337);
nor U1352 (N_1352,In_1440,In_39);
nor U1353 (N_1353,In_963,In_802);
nor U1354 (N_1354,In_722,In_1694);
nor U1355 (N_1355,In_1745,In_1113);
nand U1356 (N_1356,In_1005,In_354);
or U1357 (N_1357,In_1077,In_69);
and U1358 (N_1358,In_36,In_752);
nor U1359 (N_1359,In_809,In_2478);
or U1360 (N_1360,In_1475,In_1860);
nand U1361 (N_1361,In_245,In_172);
or U1362 (N_1362,In_1356,In_148);
nand U1363 (N_1363,In_127,In_1439);
and U1364 (N_1364,In_2192,In_2231);
nor U1365 (N_1365,In_1137,In_372);
nor U1366 (N_1366,In_487,In_2390);
nand U1367 (N_1367,In_1135,In_1533);
or U1368 (N_1368,In_430,In_2157);
nand U1369 (N_1369,In_1593,In_390);
and U1370 (N_1370,In_383,In_801);
and U1371 (N_1371,In_1013,In_1282);
or U1372 (N_1372,In_1277,In_2353);
nor U1373 (N_1373,In_938,In_2485);
and U1374 (N_1374,In_1459,In_803);
or U1375 (N_1375,In_2026,In_698);
nor U1376 (N_1376,In_2310,In_1544);
nor U1377 (N_1377,In_2001,In_1254);
xor U1378 (N_1378,In_459,In_2483);
nand U1379 (N_1379,In_953,In_2003);
nor U1380 (N_1380,In_2082,In_949);
nor U1381 (N_1381,In_833,In_531);
nor U1382 (N_1382,In_985,In_314);
nor U1383 (N_1383,In_197,In_1458);
and U1384 (N_1384,In_220,In_1798);
nor U1385 (N_1385,In_33,In_1926);
and U1386 (N_1386,In_2475,In_2309);
and U1387 (N_1387,In_1205,In_1052);
nand U1388 (N_1388,In_1292,In_862);
and U1389 (N_1389,In_1655,In_216);
or U1390 (N_1390,In_677,In_525);
nand U1391 (N_1391,In_1187,In_719);
or U1392 (N_1392,In_2210,In_1419);
nor U1393 (N_1393,In_2252,In_91);
and U1394 (N_1394,In_965,In_691);
nand U1395 (N_1395,In_60,In_784);
nor U1396 (N_1396,In_849,In_580);
nand U1397 (N_1397,In_2095,In_1408);
or U1398 (N_1398,In_1652,In_395);
nand U1399 (N_1399,In_422,In_248);
nand U1400 (N_1400,In_122,In_1297);
and U1401 (N_1401,In_2310,In_2325);
nor U1402 (N_1402,In_972,In_1379);
and U1403 (N_1403,In_2433,In_328);
nand U1404 (N_1404,In_808,In_165);
and U1405 (N_1405,In_2362,In_413);
and U1406 (N_1406,In_20,In_345);
nor U1407 (N_1407,In_775,In_2093);
xnor U1408 (N_1408,In_2052,In_615);
and U1409 (N_1409,In_375,In_1815);
or U1410 (N_1410,In_562,In_951);
and U1411 (N_1411,In_1844,In_1358);
nand U1412 (N_1412,In_419,In_1925);
and U1413 (N_1413,In_201,In_1764);
and U1414 (N_1414,In_794,In_303);
and U1415 (N_1415,In_1794,In_1810);
nand U1416 (N_1416,In_2100,In_1717);
and U1417 (N_1417,In_927,In_88);
and U1418 (N_1418,In_984,In_1451);
nand U1419 (N_1419,In_1261,In_102);
or U1420 (N_1420,In_271,In_1292);
or U1421 (N_1421,In_662,In_2060);
and U1422 (N_1422,In_1376,In_1489);
or U1423 (N_1423,In_256,In_372);
nand U1424 (N_1424,In_2318,In_358);
or U1425 (N_1425,In_358,In_1407);
and U1426 (N_1426,In_2100,In_1756);
or U1427 (N_1427,In_764,In_1);
or U1428 (N_1428,In_2397,In_389);
nor U1429 (N_1429,In_1178,In_739);
nor U1430 (N_1430,In_1929,In_2462);
nand U1431 (N_1431,In_2321,In_1291);
nor U1432 (N_1432,In_1921,In_45);
nand U1433 (N_1433,In_776,In_2491);
nand U1434 (N_1434,In_912,In_709);
and U1435 (N_1435,In_1048,In_2093);
nor U1436 (N_1436,In_908,In_2188);
or U1437 (N_1437,In_876,In_1941);
and U1438 (N_1438,In_2231,In_1104);
or U1439 (N_1439,In_777,In_887);
or U1440 (N_1440,In_741,In_873);
nor U1441 (N_1441,In_1394,In_1254);
and U1442 (N_1442,In_239,In_797);
nand U1443 (N_1443,In_309,In_1177);
or U1444 (N_1444,In_1115,In_23);
and U1445 (N_1445,In_814,In_2109);
nor U1446 (N_1446,In_923,In_1665);
nor U1447 (N_1447,In_1596,In_725);
and U1448 (N_1448,In_681,In_1560);
and U1449 (N_1449,In_2331,In_188);
nand U1450 (N_1450,In_2245,In_477);
nor U1451 (N_1451,In_930,In_1764);
and U1452 (N_1452,In_1459,In_1901);
and U1453 (N_1453,In_2265,In_1123);
or U1454 (N_1454,In_1412,In_518);
and U1455 (N_1455,In_1369,In_610);
nor U1456 (N_1456,In_2087,In_1547);
and U1457 (N_1457,In_1099,In_2458);
xnor U1458 (N_1458,In_321,In_2497);
or U1459 (N_1459,In_184,In_482);
or U1460 (N_1460,In_487,In_253);
nand U1461 (N_1461,In_1576,In_668);
nand U1462 (N_1462,In_590,In_1094);
nor U1463 (N_1463,In_572,In_422);
or U1464 (N_1464,In_1050,In_548);
nand U1465 (N_1465,In_897,In_1359);
and U1466 (N_1466,In_99,In_301);
and U1467 (N_1467,In_1981,In_298);
and U1468 (N_1468,In_397,In_87);
or U1469 (N_1469,In_2109,In_112);
or U1470 (N_1470,In_1130,In_2186);
or U1471 (N_1471,In_1764,In_2311);
and U1472 (N_1472,In_1176,In_555);
nor U1473 (N_1473,In_903,In_1113);
nor U1474 (N_1474,In_13,In_144);
nand U1475 (N_1475,In_127,In_1337);
nand U1476 (N_1476,In_900,In_2133);
and U1477 (N_1477,In_1148,In_1556);
or U1478 (N_1478,In_94,In_1971);
and U1479 (N_1479,In_2047,In_293);
or U1480 (N_1480,In_289,In_1050);
nor U1481 (N_1481,In_623,In_1722);
and U1482 (N_1482,In_2272,In_1723);
nand U1483 (N_1483,In_487,In_1988);
nor U1484 (N_1484,In_1744,In_1682);
or U1485 (N_1485,In_1392,In_2276);
or U1486 (N_1486,In_2162,In_854);
nand U1487 (N_1487,In_2311,In_394);
nand U1488 (N_1488,In_423,In_71);
and U1489 (N_1489,In_89,In_1507);
or U1490 (N_1490,In_1614,In_816);
or U1491 (N_1491,In_1120,In_904);
and U1492 (N_1492,In_1644,In_2284);
nand U1493 (N_1493,In_1039,In_1828);
nand U1494 (N_1494,In_802,In_670);
or U1495 (N_1495,In_847,In_1892);
or U1496 (N_1496,In_1692,In_169);
and U1497 (N_1497,In_1912,In_435);
or U1498 (N_1498,In_1443,In_1676);
or U1499 (N_1499,In_42,In_15);
or U1500 (N_1500,In_726,In_1832);
nor U1501 (N_1501,In_2373,In_2130);
nor U1502 (N_1502,In_22,In_1177);
nand U1503 (N_1503,In_376,In_309);
and U1504 (N_1504,In_701,In_467);
or U1505 (N_1505,In_1873,In_1237);
nand U1506 (N_1506,In_1637,In_384);
nand U1507 (N_1507,In_789,In_778);
nand U1508 (N_1508,In_308,In_25);
or U1509 (N_1509,In_2210,In_333);
nor U1510 (N_1510,In_1000,In_1928);
nor U1511 (N_1511,In_2281,In_1637);
or U1512 (N_1512,In_2259,In_1050);
or U1513 (N_1513,In_1195,In_1887);
and U1514 (N_1514,In_761,In_228);
or U1515 (N_1515,In_1407,In_1617);
and U1516 (N_1516,In_1871,In_1820);
nor U1517 (N_1517,In_139,In_732);
and U1518 (N_1518,In_296,In_1155);
nand U1519 (N_1519,In_1253,In_194);
nand U1520 (N_1520,In_1500,In_1384);
nand U1521 (N_1521,In_1079,In_2277);
nand U1522 (N_1522,In_2440,In_1994);
or U1523 (N_1523,In_675,In_1650);
or U1524 (N_1524,In_498,In_1240);
nor U1525 (N_1525,In_1381,In_2326);
nor U1526 (N_1526,In_324,In_1556);
nand U1527 (N_1527,In_45,In_15);
nor U1528 (N_1528,In_642,In_660);
nand U1529 (N_1529,In_1454,In_197);
and U1530 (N_1530,In_466,In_847);
nor U1531 (N_1531,In_136,In_698);
nor U1532 (N_1532,In_729,In_1320);
and U1533 (N_1533,In_340,In_984);
and U1534 (N_1534,In_2091,In_2000);
or U1535 (N_1535,In_1622,In_2033);
and U1536 (N_1536,In_1223,In_739);
nand U1537 (N_1537,In_615,In_2471);
nor U1538 (N_1538,In_2355,In_469);
nor U1539 (N_1539,In_1229,In_1899);
or U1540 (N_1540,In_1841,In_140);
and U1541 (N_1541,In_106,In_1217);
and U1542 (N_1542,In_1950,In_654);
nor U1543 (N_1543,In_1170,In_5);
nor U1544 (N_1544,In_1652,In_48);
and U1545 (N_1545,In_2448,In_1708);
nor U1546 (N_1546,In_574,In_1746);
and U1547 (N_1547,In_1457,In_1998);
nor U1548 (N_1548,In_339,In_2362);
or U1549 (N_1549,In_170,In_1702);
nor U1550 (N_1550,In_2301,In_398);
nand U1551 (N_1551,In_1417,In_2203);
and U1552 (N_1552,In_579,In_766);
nor U1553 (N_1553,In_2235,In_1066);
or U1554 (N_1554,In_845,In_2050);
and U1555 (N_1555,In_2471,In_1927);
nor U1556 (N_1556,In_2140,In_275);
nand U1557 (N_1557,In_2451,In_1244);
and U1558 (N_1558,In_1014,In_940);
and U1559 (N_1559,In_701,In_2272);
nor U1560 (N_1560,In_874,In_2481);
nor U1561 (N_1561,In_402,In_2438);
and U1562 (N_1562,In_1424,In_2407);
and U1563 (N_1563,In_670,In_1288);
or U1564 (N_1564,In_1569,In_2253);
nand U1565 (N_1565,In_2194,In_2187);
or U1566 (N_1566,In_540,In_1262);
and U1567 (N_1567,In_1417,In_530);
nor U1568 (N_1568,In_75,In_2396);
nor U1569 (N_1569,In_2175,In_2339);
or U1570 (N_1570,In_1912,In_1650);
nor U1571 (N_1571,In_781,In_891);
nor U1572 (N_1572,In_2054,In_231);
or U1573 (N_1573,In_1182,In_2138);
xor U1574 (N_1574,In_1703,In_695);
nor U1575 (N_1575,In_935,In_2311);
and U1576 (N_1576,In_1721,In_1507);
nand U1577 (N_1577,In_917,In_1929);
and U1578 (N_1578,In_1510,In_206);
and U1579 (N_1579,In_2022,In_469);
or U1580 (N_1580,In_846,In_1939);
nand U1581 (N_1581,In_400,In_2069);
nor U1582 (N_1582,In_1848,In_964);
or U1583 (N_1583,In_1807,In_1079);
nor U1584 (N_1584,In_2202,In_108);
and U1585 (N_1585,In_1891,In_343);
or U1586 (N_1586,In_346,In_2366);
or U1587 (N_1587,In_1997,In_1625);
and U1588 (N_1588,In_2186,In_1122);
nand U1589 (N_1589,In_1583,In_2232);
and U1590 (N_1590,In_157,In_24);
nor U1591 (N_1591,In_644,In_1137);
and U1592 (N_1592,In_1150,In_2264);
nor U1593 (N_1593,In_1870,In_406);
and U1594 (N_1594,In_234,In_1589);
nand U1595 (N_1595,In_1784,In_269);
nand U1596 (N_1596,In_1166,In_1764);
xnor U1597 (N_1597,In_1226,In_1312);
and U1598 (N_1598,In_1242,In_126);
xnor U1599 (N_1599,In_503,In_1167);
nor U1600 (N_1600,In_1775,In_1062);
or U1601 (N_1601,In_1924,In_567);
or U1602 (N_1602,In_1457,In_1580);
and U1603 (N_1603,In_605,In_784);
and U1604 (N_1604,In_1906,In_90);
nand U1605 (N_1605,In_974,In_1329);
or U1606 (N_1606,In_1124,In_1600);
nand U1607 (N_1607,In_2331,In_720);
or U1608 (N_1608,In_1664,In_1789);
or U1609 (N_1609,In_472,In_2303);
and U1610 (N_1610,In_608,In_794);
nand U1611 (N_1611,In_2221,In_1181);
nand U1612 (N_1612,In_484,In_947);
nand U1613 (N_1613,In_203,In_649);
nand U1614 (N_1614,In_1735,In_2417);
or U1615 (N_1615,In_1447,In_1283);
nand U1616 (N_1616,In_57,In_25);
or U1617 (N_1617,In_56,In_1152);
xnor U1618 (N_1618,In_1394,In_1185);
and U1619 (N_1619,In_1670,In_707);
xor U1620 (N_1620,In_1617,In_1582);
nand U1621 (N_1621,In_2141,In_1927);
nor U1622 (N_1622,In_2283,In_1499);
or U1623 (N_1623,In_477,In_472);
or U1624 (N_1624,In_2077,In_1266);
and U1625 (N_1625,In_280,In_1403);
and U1626 (N_1626,In_288,In_110);
nor U1627 (N_1627,In_610,In_1890);
and U1628 (N_1628,In_669,In_2419);
nor U1629 (N_1629,In_912,In_758);
and U1630 (N_1630,In_237,In_1141);
nor U1631 (N_1631,In_234,In_681);
or U1632 (N_1632,In_2201,In_2227);
and U1633 (N_1633,In_1299,In_1323);
nor U1634 (N_1634,In_1336,In_2214);
nand U1635 (N_1635,In_360,In_643);
nor U1636 (N_1636,In_2327,In_1197);
and U1637 (N_1637,In_2440,In_1011);
or U1638 (N_1638,In_189,In_856);
nor U1639 (N_1639,In_679,In_1048);
and U1640 (N_1640,In_2195,In_1387);
nand U1641 (N_1641,In_190,In_1641);
xnor U1642 (N_1642,In_1533,In_2403);
and U1643 (N_1643,In_1720,In_1511);
and U1644 (N_1644,In_1659,In_2158);
nor U1645 (N_1645,In_1717,In_741);
and U1646 (N_1646,In_547,In_281);
and U1647 (N_1647,In_1462,In_73);
or U1648 (N_1648,In_355,In_140);
and U1649 (N_1649,In_2045,In_2101);
or U1650 (N_1650,In_382,In_1896);
nand U1651 (N_1651,In_750,In_1210);
or U1652 (N_1652,In_1853,In_1391);
nand U1653 (N_1653,In_16,In_195);
or U1654 (N_1654,In_496,In_2233);
and U1655 (N_1655,In_2304,In_1927);
or U1656 (N_1656,In_998,In_1217);
and U1657 (N_1657,In_1028,In_1528);
or U1658 (N_1658,In_388,In_811);
nand U1659 (N_1659,In_2374,In_351);
nor U1660 (N_1660,In_474,In_1669);
and U1661 (N_1661,In_402,In_810);
nand U1662 (N_1662,In_806,In_821);
or U1663 (N_1663,In_1334,In_741);
nor U1664 (N_1664,In_2463,In_1249);
or U1665 (N_1665,In_2036,In_1248);
and U1666 (N_1666,In_1516,In_2235);
nor U1667 (N_1667,In_859,In_1761);
and U1668 (N_1668,In_920,In_1878);
or U1669 (N_1669,In_2144,In_292);
or U1670 (N_1670,In_1804,In_1637);
nor U1671 (N_1671,In_208,In_856);
nand U1672 (N_1672,In_366,In_1170);
nor U1673 (N_1673,In_15,In_1806);
nor U1674 (N_1674,In_1059,In_559);
and U1675 (N_1675,In_1903,In_1913);
nand U1676 (N_1676,In_1543,In_2001);
or U1677 (N_1677,In_1044,In_2328);
or U1678 (N_1678,In_52,In_195);
nor U1679 (N_1679,In_1674,In_1337);
nor U1680 (N_1680,In_1916,In_879);
nand U1681 (N_1681,In_1303,In_251);
and U1682 (N_1682,In_1618,In_1156);
nand U1683 (N_1683,In_1214,In_821);
nor U1684 (N_1684,In_1727,In_1157);
nand U1685 (N_1685,In_87,In_2007);
or U1686 (N_1686,In_111,In_135);
or U1687 (N_1687,In_479,In_976);
nand U1688 (N_1688,In_1385,In_1720);
xnor U1689 (N_1689,In_2223,In_2227);
nand U1690 (N_1690,In_951,In_763);
nor U1691 (N_1691,In_1368,In_2078);
and U1692 (N_1692,In_2450,In_26);
and U1693 (N_1693,In_432,In_2055);
and U1694 (N_1694,In_1990,In_529);
nand U1695 (N_1695,In_714,In_473);
nand U1696 (N_1696,In_1616,In_2135);
or U1697 (N_1697,In_1190,In_2218);
and U1698 (N_1698,In_436,In_2323);
nor U1699 (N_1699,In_924,In_1369);
nand U1700 (N_1700,In_133,In_1540);
or U1701 (N_1701,In_1713,In_2424);
or U1702 (N_1702,In_1337,In_620);
or U1703 (N_1703,In_917,In_1381);
or U1704 (N_1704,In_280,In_1763);
xnor U1705 (N_1705,In_2224,In_871);
and U1706 (N_1706,In_1224,In_1756);
and U1707 (N_1707,In_1567,In_1899);
xnor U1708 (N_1708,In_910,In_126);
and U1709 (N_1709,In_429,In_334);
nand U1710 (N_1710,In_1191,In_261);
or U1711 (N_1711,In_2051,In_872);
nor U1712 (N_1712,In_636,In_1835);
and U1713 (N_1713,In_1832,In_2445);
nand U1714 (N_1714,In_2272,In_2219);
nor U1715 (N_1715,In_189,In_714);
and U1716 (N_1716,In_124,In_1184);
or U1717 (N_1717,In_1795,In_1670);
xor U1718 (N_1718,In_2411,In_864);
or U1719 (N_1719,In_823,In_253);
nand U1720 (N_1720,In_56,In_1934);
nand U1721 (N_1721,In_1683,In_2068);
or U1722 (N_1722,In_342,In_2490);
and U1723 (N_1723,In_1209,In_16);
and U1724 (N_1724,In_432,In_2201);
nand U1725 (N_1725,In_1280,In_2015);
nand U1726 (N_1726,In_1809,In_1778);
and U1727 (N_1727,In_1471,In_2162);
and U1728 (N_1728,In_1150,In_155);
nor U1729 (N_1729,In_909,In_1654);
nor U1730 (N_1730,In_1375,In_734);
nor U1731 (N_1731,In_62,In_577);
or U1732 (N_1732,In_1039,In_1459);
nand U1733 (N_1733,In_840,In_1285);
nor U1734 (N_1734,In_1085,In_665);
nand U1735 (N_1735,In_185,In_1920);
or U1736 (N_1736,In_2261,In_270);
and U1737 (N_1737,In_2472,In_2185);
nand U1738 (N_1738,In_1036,In_1265);
nor U1739 (N_1739,In_2492,In_1641);
nand U1740 (N_1740,In_683,In_763);
nand U1741 (N_1741,In_1271,In_1306);
or U1742 (N_1742,In_1610,In_1230);
nand U1743 (N_1743,In_982,In_2250);
or U1744 (N_1744,In_876,In_1303);
nand U1745 (N_1745,In_150,In_1009);
nand U1746 (N_1746,In_2065,In_1201);
nor U1747 (N_1747,In_2109,In_215);
nand U1748 (N_1748,In_99,In_2307);
or U1749 (N_1749,In_1862,In_1913);
and U1750 (N_1750,In_173,In_2176);
nor U1751 (N_1751,In_412,In_1693);
or U1752 (N_1752,In_839,In_925);
nor U1753 (N_1753,In_874,In_2014);
nor U1754 (N_1754,In_2102,In_2419);
nor U1755 (N_1755,In_1867,In_1442);
nor U1756 (N_1756,In_2417,In_1030);
nand U1757 (N_1757,In_1933,In_144);
or U1758 (N_1758,In_1332,In_631);
or U1759 (N_1759,In_1821,In_1131);
nand U1760 (N_1760,In_1498,In_329);
nor U1761 (N_1761,In_1629,In_141);
or U1762 (N_1762,In_450,In_1044);
or U1763 (N_1763,In_540,In_8);
and U1764 (N_1764,In_427,In_442);
nor U1765 (N_1765,In_2152,In_353);
or U1766 (N_1766,In_1199,In_1534);
and U1767 (N_1767,In_1538,In_1393);
and U1768 (N_1768,In_1707,In_1890);
nor U1769 (N_1769,In_64,In_1510);
and U1770 (N_1770,In_2269,In_1192);
nor U1771 (N_1771,In_1726,In_393);
and U1772 (N_1772,In_2487,In_2044);
and U1773 (N_1773,In_1674,In_1793);
or U1774 (N_1774,In_14,In_2046);
and U1775 (N_1775,In_27,In_2352);
and U1776 (N_1776,In_1662,In_2140);
nor U1777 (N_1777,In_393,In_130);
nor U1778 (N_1778,In_243,In_946);
and U1779 (N_1779,In_644,In_1182);
or U1780 (N_1780,In_2361,In_984);
xor U1781 (N_1781,In_1943,In_400);
or U1782 (N_1782,In_1976,In_572);
nor U1783 (N_1783,In_1564,In_1616);
nand U1784 (N_1784,In_318,In_2339);
or U1785 (N_1785,In_2156,In_1398);
nand U1786 (N_1786,In_2119,In_2079);
or U1787 (N_1787,In_1485,In_22);
nor U1788 (N_1788,In_1312,In_1363);
or U1789 (N_1789,In_1066,In_629);
or U1790 (N_1790,In_778,In_1744);
and U1791 (N_1791,In_2395,In_768);
and U1792 (N_1792,In_1197,In_289);
nor U1793 (N_1793,In_1673,In_1956);
nor U1794 (N_1794,In_469,In_423);
nor U1795 (N_1795,In_2332,In_824);
and U1796 (N_1796,In_1019,In_1677);
nor U1797 (N_1797,In_1983,In_1910);
nor U1798 (N_1798,In_846,In_868);
or U1799 (N_1799,In_1309,In_1110);
and U1800 (N_1800,In_2296,In_1718);
and U1801 (N_1801,In_1560,In_2177);
and U1802 (N_1802,In_967,In_304);
nand U1803 (N_1803,In_1875,In_961);
nand U1804 (N_1804,In_1211,In_1391);
nand U1805 (N_1805,In_2050,In_1593);
nor U1806 (N_1806,In_745,In_1195);
xnor U1807 (N_1807,In_1998,In_93);
or U1808 (N_1808,In_1907,In_615);
or U1809 (N_1809,In_2080,In_1786);
nor U1810 (N_1810,In_736,In_673);
or U1811 (N_1811,In_2490,In_1103);
nor U1812 (N_1812,In_1760,In_1844);
nand U1813 (N_1813,In_1815,In_1710);
or U1814 (N_1814,In_1667,In_223);
and U1815 (N_1815,In_163,In_1396);
nor U1816 (N_1816,In_950,In_85);
and U1817 (N_1817,In_2084,In_1982);
nand U1818 (N_1818,In_2216,In_2150);
nand U1819 (N_1819,In_177,In_745);
and U1820 (N_1820,In_335,In_1531);
or U1821 (N_1821,In_1902,In_790);
or U1822 (N_1822,In_372,In_1458);
nand U1823 (N_1823,In_1174,In_1444);
or U1824 (N_1824,In_2184,In_124);
nand U1825 (N_1825,In_1283,In_1920);
and U1826 (N_1826,In_1614,In_1930);
or U1827 (N_1827,In_1287,In_53);
nand U1828 (N_1828,In_1730,In_2194);
nand U1829 (N_1829,In_55,In_711);
nor U1830 (N_1830,In_227,In_1311);
xor U1831 (N_1831,In_74,In_2048);
xor U1832 (N_1832,In_578,In_550);
or U1833 (N_1833,In_433,In_1806);
nor U1834 (N_1834,In_1843,In_1229);
or U1835 (N_1835,In_1261,In_512);
or U1836 (N_1836,In_357,In_293);
and U1837 (N_1837,In_1606,In_648);
nand U1838 (N_1838,In_1306,In_1762);
and U1839 (N_1839,In_426,In_2491);
nor U1840 (N_1840,In_358,In_491);
nand U1841 (N_1841,In_1454,In_2196);
xnor U1842 (N_1842,In_642,In_2064);
nand U1843 (N_1843,In_2051,In_746);
nor U1844 (N_1844,In_1202,In_1831);
nor U1845 (N_1845,In_2080,In_1706);
and U1846 (N_1846,In_1883,In_599);
nand U1847 (N_1847,In_1737,In_1144);
and U1848 (N_1848,In_2281,In_1376);
and U1849 (N_1849,In_767,In_1343);
nor U1850 (N_1850,In_501,In_938);
nor U1851 (N_1851,In_2280,In_635);
nand U1852 (N_1852,In_834,In_2460);
nor U1853 (N_1853,In_2273,In_1331);
nor U1854 (N_1854,In_1901,In_1921);
nand U1855 (N_1855,In_1306,In_202);
or U1856 (N_1856,In_1844,In_1842);
nor U1857 (N_1857,In_1818,In_1816);
or U1858 (N_1858,In_1772,In_1684);
nand U1859 (N_1859,In_305,In_1498);
nor U1860 (N_1860,In_1694,In_2365);
nand U1861 (N_1861,In_1779,In_1437);
nor U1862 (N_1862,In_242,In_851);
and U1863 (N_1863,In_778,In_269);
and U1864 (N_1864,In_721,In_438);
or U1865 (N_1865,In_241,In_1211);
nor U1866 (N_1866,In_880,In_678);
nor U1867 (N_1867,In_1752,In_1533);
or U1868 (N_1868,In_2332,In_2146);
nor U1869 (N_1869,In_1605,In_1552);
nor U1870 (N_1870,In_592,In_1461);
and U1871 (N_1871,In_1916,In_752);
or U1872 (N_1872,In_249,In_1831);
nor U1873 (N_1873,In_1243,In_782);
nand U1874 (N_1874,In_444,In_1299);
and U1875 (N_1875,In_517,In_573);
or U1876 (N_1876,In_113,In_1577);
nor U1877 (N_1877,In_1360,In_894);
and U1878 (N_1878,In_1602,In_2409);
nand U1879 (N_1879,In_1109,In_2011);
nand U1880 (N_1880,In_107,In_55);
nor U1881 (N_1881,In_234,In_303);
nor U1882 (N_1882,In_91,In_123);
and U1883 (N_1883,In_174,In_1815);
or U1884 (N_1884,In_724,In_1472);
nand U1885 (N_1885,In_2075,In_338);
or U1886 (N_1886,In_1187,In_1652);
nor U1887 (N_1887,In_1000,In_499);
nor U1888 (N_1888,In_2112,In_2334);
nor U1889 (N_1889,In_173,In_2193);
nor U1890 (N_1890,In_1079,In_2486);
nor U1891 (N_1891,In_99,In_1691);
and U1892 (N_1892,In_1343,In_1095);
nand U1893 (N_1893,In_1043,In_2192);
or U1894 (N_1894,In_200,In_2346);
nor U1895 (N_1895,In_1101,In_681);
nor U1896 (N_1896,In_984,In_1924);
nand U1897 (N_1897,In_696,In_1197);
nand U1898 (N_1898,In_1370,In_570);
nor U1899 (N_1899,In_1147,In_1833);
or U1900 (N_1900,In_199,In_1202);
or U1901 (N_1901,In_1847,In_1892);
or U1902 (N_1902,In_1141,In_1852);
nor U1903 (N_1903,In_1631,In_1377);
and U1904 (N_1904,In_1125,In_1273);
or U1905 (N_1905,In_540,In_1786);
or U1906 (N_1906,In_988,In_22);
and U1907 (N_1907,In_856,In_222);
nand U1908 (N_1908,In_2113,In_2346);
nor U1909 (N_1909,In_1540,In_1301);
and U1910 (N_1910,In_389,In_873);
nor U1911 (N_1911,In_2461,In_289);
nand U1912 (N_1912,In_2102,In_191);
and U1913 (N_1913,In_1923,In_1189);
or U1914 (N_1914,In_716,In_479);
nor U1915 (N_1915,In_1001,In_453);
nor U1916 (N_1916,In_1821,In_2485);
and U1917 (N_1917,In_1000,In_2062);
nand U1918 (N_1918,In_722,In_864);
nor U1919 (N_1919,In_2494,In_96);
nand U1920 (N_1920,In_1797,In_184);
and U1921 (N_1921,In_1933,In_10);
or U1922 (N_1922,In_1679,In_1092);
nand U1923 (N_1923,In_1461,In_848);
or U1924 (N_1924,In_1003,In_2001);
nand U1925 (N_1925,In_473,In_580);
nor U1926 (N_1926,In_2443,In_395);
or U1927 (N_1927,In_668,In_1635);
nand U1928 (N_1928,In_1501,In_799);
and U1929 (N_1929,In_194,In_284);
nor U1930 (N_1930,In_1363,In_2418);
nor U1931 (N_1931,In_1573,In_2192);
nor U1932 (N_1932,In_390,In_1897);
and U1933 (N_1933,In_1764,In_989);
nand U1934 (N_1934,In_1063,In_455);
nor U1935 (N_1935,In_1061,In_287);
or U1936 (N_1936,In_2024,In_1441);
nand U1937 (N_1937,In_1023,In_452);
or U1938 (N_1938,In_1083,In_803);
nand U1939 (N_1939,In_146,In_1815);
or U1940 (N_1940,In_1490,In_469);
and U1941 (N_1941,In_1055,In_1596);
nand U1942 (N_1942,In_2132,In_986);
or U1943 (N_1943,In_1457,In_1648);
and U1944 (N_1944,In_1984,In_2383);
nand U1945 (N_1945,In_2061,In_399);
and U1946 (N_1946,In_2118,In_1284);
and U1947 (N_1947,In_601,In_66);
nor U1948 (N_1948,In_603,In_348);
or U1949 (N_1949,In_1182,In_455);
nand U1950 (N_1950,In_1938,In_2119);
nand U1951 (N_1951,In_1731,In_2405);
nand U1952 (N_1952,In_2380,In_594);
or U1953 (N_1953,In_2326,In_2389);
nor U1954 (N_1954,In_2066,In_2071);
nand U1955 (N_1955,In_1915,In_1079);
xnor U1956 (N_1956,In_1926,In_1815);
nand U1957 (N_1957,In_184,In_412);
nor U1958 (N_1958,In_1389,In_1042);
nor U1959 (N_1959,In_713,In_2146);
nor U1960 (N_1960,In_1006,In_528);
or U1961 (N_1961,In_1765,In_797);
nor U1962 (N_1962,In_1489,In_1984);
nand U1963 (N_1963,In_872,In_1286);
nand U1964 (N_1964,In_1961,In_1863);
nor U1965 (N_1965,In_1525,In_2050);
xnor U1966 (N_1966,In_960,In_2371);
nor U1967 (N_1967,In_454,In_604);
or U1968 (N_1968,In_1513,In_405);
nand U1969 (N_1969,In_2219,In_1897);
and U1970 (N_1970,In_838,In_832);
or U1971 (N_1971,In_2128,In_244);
nand U1972 (N_1972,In_1480,In_2470);
nor U1973 (N_1973,In_1056,In_1823);
or U1974 (N_1974,In_548,In_1339);
nor U1975 (N_1975,In_1711,In_2215);
or U1976 (N_1976,In_640,In_1789);
or U1977 (N_1977,In_835,In_1314);
or U1978 (N_1978,In_2200,In_1905);
and U1979 (N_1979,In_1632,In_2019);
nor U1980 (N_1980,In_1437,In_1074);
nor U1981 (N_1981,In_145,In_1066);
and U1982 (N_1982,In_2362,In_1513);
nor U1983 (N_1983,In_168,In_2488);
or U1984 (N_1984,In_2149,In_2451);
xnor U1985 (N_1985,In_1076,In_1535);
nand U1986 (N_1986,In_761,In_602);
nand U1987 (N_1987,In_2262,In_509);
or U1988 (N_1988,In_1923,In_2290);
nor U1989 (N_1989,In_1227,In_1822);
nand U1990 (N_1990,In_1118,In_1759);
and U1991 (N_1991,In_1092,In_117);
nand U1992 (N_1992,In_548,In_121);
and U1993 (N_1993,In_824,In_2061);
or U1994 (N_1994,In_1010,In_1445);
and U1995 (N_1995,In_2289,In_286);
or U1996 (N_1996,In_1163,In_515);
nor U1997 (N_1997,In_754,In_347);
nor U1998 (N_1998,In_2089,In_454);
nor U1999 (N_1999,In_1333,In_1766);
nand U2000 (N_2000,In_754,In_2129);
nand U2001 (N_2001,In_1832,In_1858);
nor U2002 (N_2002,In_1645,In_1902);
or U2003 (N_2003,In_909,In_1532);
nor U2004 (N_2004,In_1020,In_2071);
xor U2005 (N_2005,In_1148,In_1535);
nor U2006 (N_2006,In_1829,In_419);
or U2007 (N_2007,In_1362,In_1550);
or U2008 (N_2008,In_321,In_1319);
nand U2009 (N_2009,In_2305,In_1918);
xnor U2010 (N_2010,In_355,In_525);
nand U2011 (N_2011,In_1020,In_296);
nor U2012 (N_2012,In_1640,In_1838);
nor U2013 (N_2013,In_408,In_853);
and U2014 (N_2014,In_1257,In_2472);
and U2015 (N_2015,In_1972,In_2098);
or U2016 (N_2016,In_2464,In_1194);
nor U2017 (N_2017,In_2088,In_2139);
xnor U2018 (N_2018,In_2218,In_2464);
and U2019 (N_2019,In_2479,In_2481);
nand U2020 (N_2020,In_460,In_251);
nand U2021 (N_2021,In_1410,In_1956);
nor U2022 (N_2022,In_1969,In_505);
nor U2023 (N_2023,In_1928,In_2022);
or U2024 (N_2024,In_1125,In_292);
and U2025 (N_2025,In_135,In_2472);
nand U2026 (N_2026,In_317,In_987);
nand U2027 (N_2027,In_1738,In_1458);
and U2028 (N_2028,In_914,In_1919);
nor U2029 (N_2029,In_688,In_1128);
and U2030 (N_2030,In_402,In_221);
nor U2031 (N_2031,In_1131,In_689);
xor U2032 (N_2032,In_2457,In_1815);
nor U2033 (N_2033,In_1038,In_1069);
nand U2034 (N_2034,In_2181,In_1419);
or U2035 (N_2035,In_869,In_2126);
and U2036 (N_2036,In_1616,In_783);
nand U2037 (N_2037,In_1383,In_977);
or U2038 (N_2038,In_841,In_1222);
or U2039 (N_2039,In_1558,In_2459);
and U2040 (N_2040,In_351,In_124);
nand U2041 (N_2041,In_674,In_1708);
or U2042 (N_2042,In_2048,In_564);
and U2043 (N_2043,In_711,In_2171);
and U2044 (N_2044,In_17,In_2463);
or U2045 (N_2045,In_1360,In_13);
and U2046 (N_2046,In_378,In_2137);
nor U2047 (N_2047,In_701,In_1543);
nand U2048 (N_2048,In_2360,In_2124);
and U2049 (N_2049,In_332,In_874);
and U2050 (N_2050,In_1222,In_1974);
nor U2051 (N_2051,In_592,In_2484);
and U2052 (N_2052,In_2052,In_2358);
nand U2053 (N_2053,In_1273,In_848);
nand U2054 (N_2054,In_724,In_1518);
or U2055 (N_2055,In_157,In_1620);
nor U2056 (N_2056,In_1730,In_1583);
nand U2057 (N_2057,In_1471,In_1468);
or U2058 (N_2058,In_921,In_2042);
or U2059 (N_2059,In_2036,In_1830);
or U2060 (N_2060,In_1786,In_591);
and U2061 (N_2061,In_1186,In_305);
nor U2062 (N_2062,In_2128,In_1241);
nand U2063 (N_2063,In_1074,In_1654);
nor U2064 (N_2064,In_175,In_772);
or U2065 (N_2065,In_1533,In_1965);
and U2066 (N_2066,In_432,In_95);
or U2067 (N_2067,In_2211,In_1297);
or U2068 (N_2068,In_2134,In_2216);
or U2069 (N_2069,In_2083,In_1572);
nand U2070 (N_2070,In_2439,In_666);
and U2071 (N_2071,In_2149,In_1076);
nor U2072 (N_2072,In_582,In_607);
or U2073 (N_2073,In_2421,In_787);
or U2074 (N_2074,In_475,In_2267);
or U2075 (N_2075,In_2115,In_1427);
nor U2076 (N_2076,In_1535,In_2144);
nor U2077 (N_2077,In_1903,In_415);
or U2078 (N_2078,In_2499,In_1264);
nand U2079 (N_2079,In_1393,In_1327);
xor U2080 (N_2080,In_2496,In_909);
or U2081 (N_2081,In_1777,In_2343);
nand U2082 (N_2082,In_1392,In_233);
nor U2083 (N_2083,In_2008,In_1172);
nor U2084 (N_2084,In_643,In_1884);
nand U2085 (N_2085,In_2203,In_796);
nor U2086 (N_2086,In_2411,In_1788);
or U2087 (N_2087,In_672,In_1321);
nor U2088 (N_2088,In_331,In_1761);
xor U2089 (N_2089,In_556,In_530);
nand U2090 (N_2090,In_1408,In_1850);
or U2091 (N_2091,In_1535,In_127);
nor U2092 (N_2092,In_553,In_1798);
or U2093 (N_2093,In_363,In_688);
and U2094 (N_2094,In_280,In_1365);
nand U2095 (N_2095,In_803,In_172);
or U2096 (N_2096,In_1694,In_317);
and U2097 (N_2097,In_697,In_2086);
nand U2098 (N_2098,In_1182,In_885);
or U2099 (N_2099,In_2402,In_1252);
and U2100 (N_2100,In_1832,In_1220);
nand U2101 (N_2101,In_451,In_1262);
nand U2102 (N_2102,In_189,In_988);
nor U2103 (N_2103,In_2458,In_1284);
and U2104 (N_2104,In_1264,In_1747);
or U2105 (N_2105,In_975,In_871);
nand U2106 (N_2106,In_2393,In_1138);
nand U2107 (N_2107,In_2289,In_9);
and U2108 (N_2108,In_301,In_1547);
or U2109 (N_2109,In_855,In_1398);
nand U2110 (N_2110,In_376,In_1125);
xnor U2111 (N_2111,In_714,In_14);
and U2112 (N_2112,In_179,In_2219);
nand U2113 (N_2113,In_586,In_925);
and U2114 (N_2114,In_2361,In_823);
or U2115 (N_2115,In_1211,In_630);
and U2116 (N_2116,In_157,In_175);
nand U2117 (N_2117,In_2390,In_1065);
nand U2118 (N_2118,In_1898,In_1184);
or U2119 (N_2119,In_1858,In_138);
and U2120 (N_2120,In_65,In_96);
nand U2121 (N_2121,In_2114,In_7);
nor U2122 (N_2122,In_1099,In_348);
nor U2123 (N_2123,In_2191,In_1986);
nand U2124 (N_2124,In_1229,In_2415);
nor U2125 (N_2125,In_1172,In_596);
nor U2126 (N_2126,In_11,In_1235);
and U2127 (N_2127,In_767,In_2360);
nor U2128 (N_2128,In_1890,In_1658);
nand U2129 (N_2129,In_2394,In_1516);
nor U2130 (N_2130,In_1199,In_1969);
nand U2131 (N_2131,In_1464,In_27);
xor U2132 (N_2132,In_1057,In_1918);
or U2133 (N_2133,In_2208,In_1885);
or U2134 (N_2134,In_1611,In_1874);
or U2135 (N_2135,In_365,In_344);
nand U2136 (N_2136,In_987,In_2339);
xnor U2137 (N_2137,In_107,In_337);
nor U2138 (N_2138,In_2204,In_2315);
or U2139 (N_2139,In_771,In_2434);
nand U2140 (N_2140,In_1441,In_1142);
or U2141 (N_2141,In_2430,In_434);
nand U2142 (N_2142,In_397,In_1799);
nand U2143 (N_2143,In_509,In_1559);
nand U2144 (N_2144,In_1736,In_2057);
and U2145 (N_2145,In_302,In_895);
and U2146 (N_2146,In_2,In_1375);
nor U2147 (N_2147,In_2349,In_808);
nor U2148 (N_2148,In_1528,In_2278);
nand U2149 (N_2149,In_2416,In_1667);
nor U2150 (N_2150,In_653,In_1091);
nand U2151 (N_2151,In_497,In_2005);
or U2152 (N_2152,In_447,In_433);
and U2153 (N_2153,In_752,In_925);
or U2154 (N_2154,In_590,In_1579);
or U2155 (N_2155,In_265,In_375);
and U2156 (N_2156,In_392,In_1331);
nand U2157 (N_2157,In_2160,In_1661);
nand U2158 (N_2158,In_841,In_2334);
nor U2159 (N_2159,In_1627,In_544);
and U2160 (N_2160,In_1456,In_945);
and U2161 (N_2161,In_1081,In_1916);
nand U2162 (N_2162,In_1174,In_2430);
nand U2163 (N_2163,In_747,In_566);
nand U2164 (N_2164,In_66,In_549);
nor U2165 (N_2165,In_152,In_89);
and U2166 (N_2166,In_770,In_1054);
and U2167 (N_2167,In_138,In_1935);
and U2168 (N_2168,In_1595,In_1352);
and U2169 (N_2169,In_1768,In_979);
nand U2170 (N_2170,In_478,In_1382);
nand U2171 (N_2171,In_1617,In_147);
or U2172 (N_2172,In_255,In_873);
and U2173 (N_2173,In_1618,In_304);
or U2174 (N_2174,In_1840,In_2025);
or U2175 (N_2175,In_1464,In_1507);
nand U2176 (N_2176,In_2074,In_935);
or U2177 (N_2177,In_287,In_2096);
and U2178 (N_2178,In_54,In_1040);
nand U2179 (N_2179,In_1353,In_13);
nand U2180 (N_2180,In_1547,In_388);
or U2181 (N_2181,In_1300,In_1911);
nand U2182 (N_2182,In_1707,In_629);
or U2183 (N_2183,In_2277,In_1573);
xnor U2184 (N_2184,In_181,In_1792);
nor U2185 (N_2185,In_1520,In_570);
nand U2186 (N_2186,In_2392,In_230);
nor U2187 (N_2187,In_2253,In_1760);
and U2188 (N_2188,In_217,In_1798);
or U2189 (N_2189,In_714,In_2256);
nand U2190 (N_2190,In_157,In_1473);
nor U2191 (N_2191,In_1951,In_1401);
nand U2192 (N_2192,In_1682,In_603);
or U2193 (N_2193,In_1126,In_1303);
or U2194 (N_2194,In_1451,In_1318);
and U2195 (N_2195,In_2012,In_1280);
nand U2196 (N_2196,In_428,In_1326);
or U2197 (N_2197,In_1963,In_1849);
nand U2198 (N_2198,In_166,In_2174);
nand U2199 (N_2199,In_198,In_1439);
nor U2200 (N_2200,In_46,In_1877);
or U2201 (N_2201,In_1578,In_2310);
nor U2202 (N_2202,In_1255,In_243);
nor U2203 (N_2203,In_118,In_1935);
nor U2204 (N_2204,In_1825,In_41);
or U2205 (N_2205,In_1808,In_614);
or U2206 (N_2206,In_1353,In_1840);
and U2207 (N_2207,In_2112,In_224);
nand U2208 (N_2208,In_109,In_606);
nor U2209 (N_2209,In_2035,In_2235);
and U2210 (N_2210,In_134,In_1927);
or U2211 (N_2211,In_1802,In_1173);
or U2212 (N_2212,In_1167,In_781);
and U2213 (N_2213,In_101,In_2165);
nor U2214 (N_2214,In_1859,In_2256);
nor U2215 (N_2215,In_949,In_743);
and U2216 (N_2216,In_1405,In_34);
or U2217 (N_2217,In_710,In_1115);
nand U2218 (N_2218,In_2045,In_774);
and U2219 (N_2219,In_1006,In_385);
nor U2220 (N_2220,In_2180,In_777);
and U2221 (N_2221,In_607,In_228);
and U2222 (N_2222,In_2243,In_1716);
nand U2223 (N_2223,In_1548,In_755);
nand U2224 (N_2224,In_10,In_2301);
nand U2225 (N_2225,In_2135,In_1563);
nand U2226 (N_2226,In_438,In_1869);
nand U2227 (N_2227,In_64,In_54);
or U2228 (N_2228,In_2397,In_870);
or U2229 (N_2229,In_2245,In_1052);
nor U2230 (N_2230,In_822,In_398);
nor U2231 (N_2231,In_909,In_942);
nand U2232 (N_2232,In_1040,In_1359);
or U2233 (N_2233,In_2255,In_669);
nand U2234 (N_2234,In_1803,In_696);
nor U2235 (N_2235,In_1552,In_1539);
nor U2236 (N_2236,In_1157,In_2334);
nand U2237 (N_2237,In_606,In_2047);
or U2238 (N_2238,In_2412,In_1650);
or U2239 (N_2239,In_263,In_698);
nand U2240 (N_2240,In_1532,In_2276);
nor U2241 (N_2241,In_1227,In_1930);
or U2242 (N_2242,In_1286,In_914);
and U2243 (N_2243,In_1662,In_2308);
and U2244 (N_2244,In_721,In_958);
and U2245 (N_2245,In_962,In_513);
nand U2246 (N_2246,In_998,In_989);
nand U2247 (N_2247,In_2035,In_526);
nor U2248 (N_2248,In_1000,In_1584);
xnor U2249 (N_2249,In_707,In_301);
xor U2250 (N_2250,In_413,In_390);
nand U2251 (N_2251,In_915,In_301);
nand U2252 (N_2252,In_681,In_858);
or U2253 (N_2253,In_2002,In_346);
or U2254 (N_2254,In_1875,In_2498);
nand U2255 (N_2255,In_1634,In_1448);
and U2256 (N_2256,In_1253,In_1065);
or U2257 (N_2257,In_1443,In_2330);
nor U2258 (N_2258,In_1632,In_529);
nor U2259 (N_2259,In_1655,In_241);
nor U2260 (N_2260,In_7,In_94);
nand U2261 (N_2261,In_2005,In_1073);
nor U2262 (N_2262,In_599,In_669);
or U2263 (N_2263,In_1095,In_758);
or U2264 (N_2264,In_2009,In_160);
and U2265 (N_2265,In_1265,In_116);
or U2266 (N_2266,In_813,In_1084);
nand U2267 (N_2267,In_36,In_2480);
nand U2268 (N_2268,In_245,In_460);
and U2269 (N_2269,In_2256,In_1130);
or U2270 (N_2270,In_1900,In_812);
nand U2271 (N_2271,In_2333,In_2059);
nand U2272 (N_2272,In_2106,In_2269);
nor U2273 (N_2273,In_826,In_2184);
nor U2274 (N_2274,In_923,In_1559);
nand U2275 (N_2275,In_614,In_260);
and U2276 (N_2276,In_271,In_1909);
nand U2277 (N_2277,In_477,In_939);
nand U2278 (N_2278,In_1966,In_1782);
nor U2279 (N_2279,In_733,In_1916);
or U2280 (N_2280,In_1678,In_2329);
or U2281 (N_2281,In_907,In_1286);
nor U2282 (N_2282,In_510,In_91);
nand U2283 (N_2283,In_1166,In_1473);
nor U2284 (N_2284,In_520,In_235);
and U2285 (N_2285,In_1819,In_1171);
and U2286 (N_2286,In_2440,In_1944);
and U2287 (N_2287,In_2423,In_2297);
nor U2288 (N_2288,In_1960,In_1167);
xor U2289 (N_2289,In_588,In_2150);
and U2290 (N_2290,In_1271,In_2153);
or U2291 (N_2291,In_1192,In_2078);
nand U2292 (N_2292,In_2273,In_2171);
or U2293 (N_2293,In_1836,In_915);
or U2294 (N_2294,In_1124,In_1956);
nand U2295 (N_2295,In_221,In_1178);
nand U2296 (N_2296,In_173,In_2182);
and U2297 (N_2297,In_625,In_870);
nor U2298 (N_2298,In_289,In_1879);
and U2299 (N_2299,In_1348,In_962);
nand U2300 (N_2300,In_1298,In_2489);
nand U2301 (N_2301,In_435,In_259);
xnor U2302 (N_2302,In_1610,In_250);
and U2303 (N_2303,In_1859,In_1183);
nand U2304 (N_2304,In_106,In_254);
nand U2305 (N_2305,In_539,In_194);
or U2306 (N_2306,In_1038,In_609);
or U2307 (N_2307,In_2159,In_824);
or U2308 (N_2308,In_1081,In_1214);
nand U2309 (N_2309,In_1608,In_1742);
and U2310 (N_2310,In_802,In_1667);
or U2311 (N_2311,In_2452,In_2217);
nor U2312 (N_2312,In_2431,In_2018);
nand U2313 (N_2313,In_1276,In_2382);
nand U2314 (N_2314,In_940,In_1352);
nor U2315 (N_2315,In_1813,In_1456);
nand U2316 (N_2316,In_733,In_1281);
or U2317 (N_2317,In_489,In_1595);
and U2318 (N_2318,In_453,In_1023);
nand U2319 (N_2319,In_341,In_144);
nor U2320 (N_2320,In_1369,In_1854);
nor U2321 (N_2321,In_1052,In_1166);
nor U2322 (N_2322,In_1009,In_2023);
and U2323 (N_2323,In_585,In_2369);
nand U2324 (N_2324,In_1228,In_1248);
or U2325 (N_2325,In_1320,In_2169);
nor U2326 (N_2326,In_1318,In_1618);
nor U2327 (N_2327,In_2223,In_720);
and U2328 (N_2328,In_335,In_1139);
nor U2329 (N_2329,In_2104,In_1085);
or U2330 (N_2330,In_2129,In_2269);
and U2331 (N_2331,In_885,In_987);
and U2332 (N_2332,In_1890,In_2320);
and U2333 (N_2333,In_460,In_2202);
and U2334 (N_2334,In_1074,In_83);
nand U2335 (N_2335,In_1446,In_1915);
nand U2336 (N_2336,In_1132,In_1197);
nand U2337 (N_2337,In_2401,In_1984);
or U2338 (N_2338,In_1302,In_337);
nor U2339 (N_2339,In_39,In_470);
nand U2340 (N_2340,In_791,In_2361);
and U2341 (N_2341,In_971,In_1271);
nand U2342 (N_2342,In_2488,In_377);
xor U2343 (N_2343,In_373,In_445);
and U2344 (N_2344,In_582,In_519);
nand U2345 (N_2345,In_98,In_900);
and U2346 (N_2346,In_961,In_1610);
nand U2347 (N_2347,In_656,In_1714);
and U2348 (N_2348,In_1004,In_248);
nand U2349 (N_2349,In_1904,In_354);
nand U2350 (N_2350,In_550,In_109);
nand U2351 (N_2351,In_1307,In_1696);
xnor U2352 (N_2352,In_1363,In_831);
and U2353 (N_2353,In_1255,In_74);
and U2354 (N_2354,In_1210,In_1566);
and U2355 (N_2355,In_1450,In_1004);
nand U2356 (N_2356,In_2373,In_2353);
or U2357 (N_2357,In_803,In_41);
and U2358 (N_2358,In_1075,In_2080);
nor U2359 (N_2359,In_929,In_2276);
and U2360 (N_2360,In_1764,In_1677);
or U2361 (N_2361,In_790,In_1989);
nor U2362 (N_2362,In_924,In_525);
nand U2363 (N_2363,In_1929,In_717);
nor U2364 (N_2364,In_1583,In_478);
or U2365 (N_2365,In_1827,In_1829);
nor U2366 (N_2366,In_1078,In_1098);
or U2367 (N_2367,In_1698,In_1983);
nor U2368 (N_2368,In_566,In_1139);
or U2369 (N_2369,In_62,In_1580);
or U2370 (N_2370,In_860,In_2084);
or U2371 (N_2371,In_2498,In_1620);
and U2372 (N_2372,In_2215,In_60);
xnor U2373 (N_2373,In_446,In_1261);
nand U2374 (N_2374,In_306,In_1498);
nor U2375 (N_2375,In_43,In_2183);
and U2376 (N_2376,In_482,In_1665);
nor U2377 (N_2377,In_2123,In_1413);
nand U2378 (N_2378,In_2230,In_1162);
or U2379 (N_2379,In_815,In_1888);
nand U2380 (N_2380,In_1752,In_1590);
xor U2381 (N_2381,In_1047,In_2184);
xor U2382 (N_2382,In_1265,In_2084);
or U2383 (N_2383,In_966,In_841);
and U2384 (N_2384,In_2429,In_809);
or U2385 (N_2385,In_1225,In_521);
nor U2386 (N_2386,In_652,In_65);
nor U2387 (N_2387,In_2416,In_1750);
nor U2388 (N_2388,In_2129,In_1317);
nand U2389 (N_2389,In_40,In_419);
nand U2390 (N_2390,In_1334,In_1732);
nand U2391 (N_2391,In_1858,In_1774);
and U2392 (N_2392,In_116,In_198);
nand U2393 (N_2393,In_279,In_1299);
nand U2394 (N_2394,In_1258,In_776);
nand U2395 (N_2395,In_2381,In_345);
and U2396 (N_2396,In_266,In_1409);
or U2397 (N_2397,In_1847,In_1448);
or U2398 (N_2398,In_1307,In_1059);
or U2399 (N_2399,In_2448,In_2417);
nand U2400 (N_2400,In_773,In_451);
nor U2401 (N_2401,In_1023,In_2068);
nand U2402 (N_2402,In_1152,In_1252);
or U2403 (N_2403,In_1313,In_2119);
and U2404 (N_2404,In_1417,In_1427);
or U2405 (N_2405,In_805,In_1582);
nand U2406 (N_2406,In_1939,In_421);
nand U2407 (N_2407,In_2316,In_813);
and U2408 (N_2408,In_2165,In_1111);
and U2409 (N_2409,In_1004,In_2095);
nand U2410 (N_2410,In_1747,In_361);
nor U2411 (N_2411,In_1254,In_2139);
nand U2412 (N_2412,In_364,In_2454);
or U2413 (N_2413,In_2245,In_20);
and U2414 (N_2414,In_1273,In_2184);
and U2415 (N_2415,In_1868,In_2408);
and U2416 (N_2416,In_868,In_149);
or U2417 (N_2417,In_1800,In_1238);
or U2418 (N_2418,In_293,In_71);
or U2419 (N_2419,In_2239,In_1949);
nor U2420 (N_2420,In_469,In_1140);
or U2421 (N_2421,In_2392,In_548);
or U2422 (N_2422,In_2157,In_435);
and U2423 (N_2423,In_867,In_2405);
and U2424 (N_2424,In_2194,In_800);
and U2425 (N_2425,In_775,In_2031);
xnor U2426 (N_2426,In_1032,In_2026);
and U2427 (N_2427,In_1631,In_584);
nand U2428 (N_2428,In_343,In_1132);
and U2429 (N_2429,In_335,In_1502);
and U2430 (N_2430,In_289,In_718);
nor U2431 (N_2431,In_120,In_700);
nor U2432 (N_2432,In_1327,In_394);
nand U2433 (N_2433,In_529,In_2028);
nor U2434 (N_2434,In_1822,In_460);
or U2435 (N_2435,In_794,In_897);
or U2436 (N_2436,In_819,In_2498);
nand U2437 (N_2437,In_210,In_553);
and U2438 (N_2438,In_1629,In_773);
or U2439 (N_2439,In_2378,In_73);
xnor U2440 (N_2440,In_2060,In_651);
nor U2441 (N_2441,In_180,In_937);
nand U2442 (N_2442,In_422,In_13);
and U2443 (N_2443,In_580,In_2422);
or U2444 (N_2444,In_2211,In_673);
nor U2445 (N_2445,In_398,In_653);
or U2446 (N_2446,In_82,In_1246);
nor U2447 (N_2447,In_1767,In_1513);
nand U2448 (N_2448,In_2169,In_911);
and U2449 (N_2449,In_96,In_1440);
nand U2450 (N_2450,In_1416,In_366);
nor U2451 (N_2451,In_2073,In_553);
or U2452 (N_2452,In_1607,In_215);
nor U2453 (N_2453,In_1699,In_1864);
and U2454 (N_2454,In_848,In_887);
nand U2455 (N_2455,In_1163,In_1605);
and U2456 (N_2456,In_523,In_416);
nand U2457 (N_2457,In_2235,In_27);
or U2458 (N_2458,In_376,In_765);
nand U2459 (N_2459,In_2238,In_2160);
nor U2460 (N_2460,In_935,In_576);
xnor U2461 (N_2461,In_80,In_2303);
and U2462 (N_2462,In_63,In_1627);
nor U2463 (N_2463,In_1380,In_1856);
nor U2464 (N_2464,In_2430,In_1326);
or U2465 (N_2465,In_1419,In_2207);
or U2466 (N_2466,In_2079,In_2142);
and U2467 (N_2467,In_599,In_297);
xnor U2468 (N_2468,In_2358,In_1806);
nor U2469 (N_2469,In_2008,In_1075);
nor U2470 (N_2470,In_2198,In_1959);
or U2471 (N_2471,In_1708,In_1775);
or U2472 (N_2472,In_1128,In_2230);
and U2473 (N_2473,In_550,In_1092);
or U2474 (N_2474,In_350,In_2338);
and U2475 (N_2475,In_32,In_2188);
or U2476 (N_2476,In_559,In_1956);
or U2477 (N_2477,In_465,In_1973);
and U2478 (N_2478,In_2103,In_2131);
or U2479 (N_2479,In_717,In_2137);
and U2480 (N_2480,In_1049,In_2170);
nor U2481 (N_2481,In_2434,In_2143);
and U2482 (N_2482,In_563,In_1914);
nand U2483 (N_2483,In_109,In_629);
and U2484 (N_2484,In_2114,In_672);
and U2485 (N_2485,In_638,In_440);
or U2486 (N_2486,In_591,In_2158);
and U2487 (N_2487,In_2197,In_2370);
nor U2488 (N_2488,In_1932,In_2220);
and U2489 (N_2489,In_623,In_489);
nor U2490 (N_2490,In_200,In_2136);
nor U2491 (N_2491,In_231,In_1941);
nand U2492 (N_2492,In_2286,In_534);
or U2493 (N_2493,In_166,In_1094);
or U2494 (N_2494,In_1046,In_2310);
nand U2495 (N_2495,In_1744,In_1640);
or U2496 (N_2496,In_2201,In_231);
nor U2497 (N_2497,In_1824,In_1875);
and U2498 (N_2498,In_882,In_2076);
nand U2499 (N_2499,In_958,In_874);
nor U2500 (N_2500,In_1203,In_1572);
xor U2501 (N_2501,In_1111,In_859);
xor U2502 (N_2502,In_786,In_937);
and U2503 (N_2503,In_1085,In_1000);
nor U2504 (N_2504,In_1446,In_1752);
and U2505 (N_2505,In_1141,In_1998);
nor U2506 (N_2506,In_846,In_955);
nor U2507 (N_2507,In_2333,In_1088);
nor U2508 (N_2508,In_645,In_2343);
or U2509 (N_2509,In_1099,In_275);
and U2510 (N_2510,In_1837,In_408);
nor U2511 (N_2511,In_1422,In_1816);
nand U2512 (N_2512,In_2215,In_1137);
nor U2513 (N_2513,In_39,In_1294);
or U2514 (N_2514,In_1836,In_105);
nor U2515 (N_2515,In_50,In_789);
or U2516 (N_2516,In_728,In_807);
nand U2517 (N_2517,In_1660,In_2419);
nand U2518 (N_2518,In_1043,In_674);
and U2519 (N_2519,In_1578,In_803);
nand U2520 (N_2520,In_1674,In_386);
or U2521 (N_2521,In_873,In_1173);
and U2522 (N_2522,In_493,In_2230);
nor U2523 (N_2523,In_14,In_1050);
nand U2524 (N_2524,In_1495,In_509);
or U2525 (N_2525,In_1897,In_1723);
and U2526 (N_2526,In_1924,In_1909);
and U2527 (N_2527,In_1938,In_1526);
and U2528 (N_2528,In_2443,In_1104);
and U2529 (N_2529,In_2417,In_605);
and U2530 (N_2530,In_833,In_1992);
nor U2531 (N_2531,In_1290,In_696);
nand U2532 (N_2532,In_1971,In_2403);
and U2533 (N_2533,In_362,In_616);
nand U2534 (N_2534,In_89,In_1810);
nor U2535 (N_2535,In_2396,In_1607);
nor U2536 (N_2536,In_1351,In_970);
nand U2537 (N_2537,In_456,In_1139);
or U2538 (N_2538,In_1802,In_1);
nand U2539 (N_2539,In_1141,In_2115);
nor U2540 (N_2540,In_1743,In_629);
and U2541 (N_2541,In_696,In_2497);
and U2542 (N_2542,In_1612,In_36);
nand U2543 (N_2543,In_1889,In_2306);
or U2544 (N_2544,In_769,In_756);
nor U2545 (N_2545,In_1630,In_1010);
nand U2546 (N_2546,In_1798,In_1673);
nor U2547 (N_2547,In_549,In_1395);
and U2548 (N_2548,In_234,In_1178);
nand U2549 (N_2549,In_1225,In_650);
nand U2550 (N_2550,In_1000,In_333);
or U2551 (N_2551,In_1618,In_526);
and U2552 (N_2552,In_2233,In_446);
or U2553 (N_2553,In_2238,In_1633);
nand U2554 (N_2554,In_133,In_458);
and U2555 (N_2555,In_1813,In_407);
nor U2556 (N_2556,In_159,In_1495);
or U2557 (N_2557,In_2014,In_912);
or U2558 (N_2558,In_1768,In_1070);
and U2559 (N_2559,In_2040,In_1790);
nand U2560 (N_2560,In_1562,In_629);
and U2561 (N_2561,In_487,In_1274);
nor U2562 (N_2562,In_467,In_1541);
and U2563 (N_2563,In_1599,In_1053);
nor U2564 (N_2564,In_624,In_690);
nor U2565 (N_2565,In_521,In_1248);
nand U2566 (N_2566,In_2494,In_512);
nand U2567 (N_2567,In_449,In_300);
nand U2568 (N_2568,In_2050,In_1342);
or U2569 (N_2569,In_1942,In_2156);
and U2570 (N_2570,In_669,In_2265);
nand U2571 (N_2571,In_1496,In_285);
or U2572 (N_2572,In_1481,In_1016);
nor U2573 (N_2573,In_1365,In_2039);
and U2574 (N_2574,In_1060,In_1111);
nand U2575 (N_2575,In_986,In_1791);
or U2576 (N_2576,In_353,In_352);
and U2577 (N_2577,In_686,In_1283);
nor U2578 (N_2578,In_2130,In_2030);
and U2579 (N_2579,In_241,In_2231);
nor U2580 (N_2580,In_2383,In_1266);
and U2581 (N_2581,In_123,In_665);
nor U2582 (N_2582,In_1386,In_907);
and U2583 (N_2583,In_949,In_1347);
or U2584 (N_2584,In_1435,In_1992);
and U2585 (N_2585,In_2408,In_2481);
and U2586 (N_2586,In_18,In_1665);
and U2587 (N_2587,In_1276,In_2422);
nor U2588 (N_2588,In_1371,In_1773);
or U2589 (N_2589,In_1736,In_2249);
nand U2590 (N_2590,In_1392,In_835);
and U2591 (N_2591,In_10,In_1997);
or U2592 (N_2592,In_131,In_1901);
and U2593 (N_2593,In_721,In_1861);
nor U2594 (N_2594,In_544,In_511);
and U2595 (N_2595,In_1309,In_1592);
nor U2596 (N_2596,In_2108,In_529);
or U2597 (N_2597,In_1426,In_2154);
and U2598 (N_2598,In_1584,In_2333);
or U2599 (N_2599,In_90,In_250);
nor U2600 (N_2600,In_380,In_204);
nor U2601 (N_2601,In_1165,In_799);
or U2602 (N_2602,In_761,In_1276);
nand U2603 (N_2603,In_1011,In_1032);
nor U2604 (N_2604,In_878,In_599);
and U2605 (N_2605,In_2087,In_438);
nor U2606 (N_2606,In_1748,In_415);
or U2607 (N_2607,In_1762,In_1390);
or U2608 (N_2608,In_830,In_1457);
and U2609 (N_2609,In_1210,In_1922);
and U2610 (N_2610,In_2482,In_587);
and U2611 (N_2611,In_2428,In_2016);
nor U2612 (N_2612,In_2448,In_1958);
nor U2613 (N_2613,In_947,In_2039);
nand U2614 (N_2614,In_1788,In_412);
and U2615 (N_2615,In_1109,In_516);
xnor U2616 (N_2616,In_139,In_1746);
nand U2617 (N_2617,In_1473,In_2370);
nand U2618 (N_2618,In_5,In_1434);
nor U2619 (N_2619,In_1837,In_726);
nand U2620 (N_2620,In_1886,In_1309);
nand U2621 (N_2621,In_1611,In_366);
or U2622 (N_2622,In_1217,In_994);
or U2623 (N_2623,In_2458,In_1232);
nand U2624 (N_2624,In_1897,In_1982);
xor U2625 (N_2625,In_1982,In_371);
nor U2626 (N_2626,In_2093,In_317);
or U2627 (N_2627,In_2433,In_1125);
nand U2628 (N_2628,In_676,In_1812);
nand U2629 (N_2629,In_949,In_663);
or U2630 (N_2630,In_1112,In_853);
and U2631 (N_2631,In_353,In_606);
and U2632 (N_2632,In_2349,In_297);
nor U2633 (N_2633,In_1503,In_1881);
or U2634 (N_2634,In_1377,In_703);
and U2635 (N_2635,In_171,In_1012);
nor U2636 (N_2636,In_710,In_73);
or U2637 (N_2637,In_422,In_1973);
nand U2638 (N_2638,In_654,In_1810);
and U2639 (N_2639,In_1759,In_1134);
and U2640 (N_2640,In_1495,In_2279);
nand U2641 (N_2641,In_1761,In_1302);
or U2642 (N_2642,In_209,In_1093);
and U2643 (N_2643,In_1881,In_369);
and U2644 (N_2644,In_1947,In_53);
nor U2645 (N_2645,In_1659,In_2070);
and U2646 (N_2646,In_93,In_1731);
and U2647 (N_2647,In_1967,In_2272);
nor U2648 (N_2648,In_853,In_91);
nor U2649 (N_2649,In_1802,In_1917);
and U2650 (N_2650,In_595,In_478);
and U2651 (N_2651,In_2197,In_1436);
nand U2652 (N_2652,In_2352,In_162);
or U2653 (N_2653,In_1202,In_1027);
or U2654 (N_2654,In_1809,In_1927);
and U2655 (N_2655,In_1367,In_1405);
or U2656 (N_2656,In_523,In_981);
or U2657 (N_2657,In_2174,In_2251);
nand U2658 (N_2658,In_1316,In_550);
and U2659 (N_2659,In_1111,In_2467);
nand U2660 (N_2660,In_2038,In_1798);
or U2661 (N_2661,In_2022,In_715);
nor U2662 (N_2662,In_2272,In_2421);
nand U2663 (N_2663,In_1904,In_1516);
or U2664 (N_2664,In_563,In_2441);
nor U2665 (N_2665,In_322,In_204);
nor U2666 (N_2666,In_326,In_1664);
xnor U2667 (N_2667,In_1025,In_850);
or U2668 (N_2668,In_2210,In_1120);
and U2669 (N_2669,In_1682,In_2172);
and U2670 (N_2670,In_451,In_1599);
nand U2671 (N_2671,In_1743,In_2215);
nor U2672 (N_2672,In_2207,In_215);
and U2673 (N_2673,In_1155,In_1711);
and U2674 (N_2674,In_387,In_1206);
or U2675 (N_2675,In_381,In_1905);
nor U2676 (N_2676,In_186,In_2157);
nor U2677 (N_2677,In_1283,In_1855);
and U2678 (N_2678,In_662,In_1111);
nand U2679 (N_2679,In_1684,In_523);
nand U2680 (N_2680,In_904,In_418);
and U2681 (N_2681,In_1151,In_1613);
nor U2682 (N_2682,In_801,In_509);
nand U2683 (N_2683,In_1611,In_1833);
xnor U2684 (N_2684,In_2406,In_491);
nand U2685 (N_2685,In_2316,In_2308);
or U2686 (N_2686,In_125,In_238);
nor U2687 (N_2687,In_605,In_2326);
and U2688 (N_2688,In_1689,In_299);
nor U2689 (N_2689,In_2413,In_1290);
or U2690 (N_2690,In_320,In_1312);
or U2691 (N_2691,In_292,In_432);
and U2692 (N_2692,In_2350,In_1693);
nand U2693 (N_2693,In_1610,In_2453);
nor U2694 (N_2694,In_1009,In_1887);
or U2695 (N_2695,In_1542,In_648);
nand U2696 (N_2696,In_2422,In_1656);
and U2697 (N_2697,In_2425,In_764);
nand U2698 (N_2698,In_2485,In_1347);
xor U2699 (N_2699,In_901,In_1258);
nor U2700 (N_2700,In_2468,In_2133);
and U2701 (N_2701,In_1915,In_1123);
nand U2702 (N_2702,In_633,In_703);
or U2703 (N_2703,In_381,In_1585);
and U2704 (N_2704,In_1462,In_1857);
nor U2705 (N_2705,In_2029,In_1027);
and U2706 (N_2706,In_45,In_508);
nand U2707 (N_2707,In_1144,In_1695);
nor U2708 (N_2708,In_773,In_2075);
or U2709 (N_2709,In_2294,In_2057);
or U2710 (N_2710,In_340,In_1273);
and U2711 (N_2711,In_962,In_1495);
and U2712 (N_2712,In_1591,In_530);
nor U2713 (N_2713,In_2184,In_217);
or U2714 (N_2714,In_1131,In_614);
nand U2715 (N_2715,In_1143,In_1443);
nand U2716 (N_2716,In_594,In_2444);
nand U2717 (N_2717,In_2078,In_822);
and U2718 (N_2718,In_444,In_320);
and U2719 (N_2719,In_1107,In_161);
nor U2720 (N_2720,In_2379,In_2450);
nor U2721 (N_2721,In_1195,In_1908);
nand U2722 (N_2722,In_1269,In_1393);
and U2723 (N_2723,In_83,In_504);
nand U2724 (N_2724,In_2310,In_1559);
xnor U2725 (N_2725,In_653,In_770);
nor U2726 (N_2726,In_515,In_1588);
nor U2727 (N_2727,In_1240,In_1353);
nor U2728 (N_2728,In_2241,In_1548);
or U2729 (N_2729,In_453,In_1616);
nand U2730 (N_2730,In_712,In_1811);
or U2731 (N_2731,In_721,In_1932);
or U2732 (N_2732,In_2341,In_2253);
or U2733 (N_2733,In_1526,In_1721);
and U2734 (N_2734,In_1990,In_219);
nor U2735 (N_2735,In_2172,In_1745);
nand U2736 (N_2736,In_2468,In_364);
or U2737 (N_2737,In_1818,In_1603);
and U2738 (N_2738,In_2097,In_1424);
nand U2739 (N_2739,In_2205,In_784);
and U2740 (N_2740,In_339,In_1533);
nand U2741 (N_2741,In_2464,In_2355);
or U2742 (N_2742,In_783,In_712);
and U2743 (N_2743,In_2237,In_1748);
nor U2744 (N_2744,In_2306,In_778);
and U2745 (N_2745,In_1586,In_625);
and U2746 (N_2746,In_1793,In_1689);
and U2747 (N_2747,In_2288,In_644);
nor U2748 (N_2748,In_1296,In_1568);
nand U2749 (N_2749,In_2298,In_1770);
and U2750 (N_2750,In_1866,In_788);
and U2751 (N_2751,In_133,In_1012);
and U2752 (N_2752,In_359,In_1721);
nand U2753 (N_2753,In_1456,In_1231);
and U2754 (N_2754,In_2057,In_1489);
nor U2755 (N_2755,In_968,In_208);
or U2756 (N_2756,In_91,In_2088);
nand U2757 (N_2757,In_2241,In_2315);
or U2758 (N_2758,In_1151,In_530);
and U2759 (N_2759,In_761,In_1946);
and U2760 (N_2760,In_788,In_467);
nor U2761 (N_2761,In_1738,In_1578);
nor U2762 (N_2762,In_2267,In_155);
and U2763 (N_2763,In_2314,In_1988);
or U2764 (N_2764,In_2381,In_1518);
and U2765 (N_2765,In_1201,In_1582);
or U2766 (N_2766,In_2392,In_1332);
nor U2767 (N_2767,In_1853,In_1578);
nand U2768 (N_2768,In_2124,In_1284);
and U2769 (N_2769,In_2474,In_1690);
or U2770 (N_2770,In_1008,In_708);
nand U2771 (N_2771,In_1405,In_157);
and U2772 (N_2772,In_2017,In_503);
nor U2773 (N_2773,In_2443,In_2176);
nor U2774 (N_2774,In_1506,In_96);
nor U2775 (N_2775,In_542,In_1568);
nor U2776 (N_2776,In_525,In_902);
and U2777 (N_2777,In_1951,In_1901);
or U2778 (N_2778,In_1060,In_626);
or U2779 (N_2779,In_2471,In_82);
and U2780 (N_2780,In_939,In_769);
nor U2781 (N_2781,In_1361,In_94);
nor U2782 (N_2782,In_1891,In_1084);
nand U2783 (N_2783,In_2235,In_382);
nand U2784 (N_2784,In_2079,In_1647);
nor U2785 (N_2785,In_107,In_1427);
nor U2786 (N_2786,In_1791,In_2434);
or U2787 (N_2787,In_1133,In_1293);
nor U2788 (N_2788,In_270,In_2069);
nor U2789 (N_2789,In_1224,In_1937);
nor U2790 (N_2790,In_1516,In_6);
or U2791 (N_2791,In_2011,In_2101);
or U2792 (N_2792,In_85,In_1369);
nor U2793 (N_2793,In_231,In_1030);
nor U2794 (N_2794,In_2122,In_2080);
nand U2795 (N_2795,In_1161,In_2383);
and U2796 (N_2796,In_929,In_165);
nor U2797 (N_2797,In_68,In_2400);
nand U2798 (N_2798,In_2147,In_2289);
xnor U2799 (N_2799,In_614,In_413);
xor U2800 (N_2800,In_771,In_953);
xnor U2801 (N_2801,In_400,In_946);
nand U2802 (N_2802,In_513,In_476);
and U2803 (N_2803,In_1876,In_433);
nor U2804 (N_2804,In_1198,In_1840);
and U2805 (N_2805,In_1499,In_2259);
and U2806 (N_2806,In_2155,In_1921);
nor U2807 (N_2807,In_589,In_319);
nor U2808 (N_2808,In_230,In_2361);
and U2809 (N_2809,In_1567,In_2000);
nand U2810 (N_2810,In_355,In_935);
nor U2811 (N_2811,In_2109,In_1445);
nand U2812 (N_2812,In_235,In_2167);
nor U2813 (N_2813,In_2271,In_1283);
or U2814 (N_2814,In_1374,In_901);
and U2815 (N_2815,In_717,In_2114);
nand U2816 (N_2816,In_1303,In_1527);
nand U2817 (N_2817,In_601,In_978);
nand U2818 (N_2818,In_179,In_1078);
nand U2819 (N_2819,In_202,In_2322);
nor U2820 (N_2820,In_1810,In_1855);
and U2821 (N_2821,In_694,In_1515);
nor U2822 (N_2822,In_1726,In_1416);
nand U2823 (N_2823,In_1457,In_2280);
or U2824 (N_2824,In_1321,In_968);
or U2825 (N_2825,In_532,In_1915);
or U2826 (N_2826,In_2485,In_608);
and U2827 (N_2827,In_1498,In_778);
and U2828 (N_2828,In_2241,In_761);
or U2829 (N_2829,In_116,In_723);
nor U2830 (N_2830,In_4,In_1146);
or U2831 (N_2831,In_180,In_2066);
nor U2832 (N_2832,In_880,In_1372);
or U2833 (N_2833,In_2302,In_337);
and U2834 (N_2834,In_1624,In_54);
or U2835 (N_2835,In_1467,In_1670);
nand U2836 (N_2836,In_2409,In_546);
nand U2837 (N_2837,In_1070,In_1174);
and U2838 (N_2838,In_2309,In_545);
and U2839 (N_2839,In_175,In_1958);
nor U2840 (N_2840,In_52,In_1408);
nor U2841 (N_2841,In_451,In_179);
nand U2842 (N_2842,In_1313,In_348);
nand U2843 (N_2843,In_293,In_52);
or U2844 (N_2844,In_245,In_1215);
and U2845 (N_2845,In_2,In_432);
nand U2846 (N_2846,In_164,In_75);
and U2847 (N_2847,In_1149,In_1383);
nand U2848 (N_2848,In_197,In_649);
nand U2849 (N_2849,In_386,In_1331);
nor U2850 (N_2850,In_1556,In_2269);
or U2851 (N_2851,In_2449,In_1346);
nor U2852 (N_2852,In_1974,In_1838);
nand U2853 (N_2853,In_2324,In_991);
xnor U2854 (N_2854,In_896,In_1020);
nand U2855 (N_2855,In_2092,In_286);
nor U2856 (N_2856,In_828,In_1822);
nand U2857 (N_2857,In_1755,In_1708);
nand U2858 (N_2858,In_1458,In_1133);
or U2859 (N_2859,In_83,In_1805);
and U2860 (N_2860,In_65,In_2187);
nor U2861 (N_2861,In_359,In_47);
nand U2862 (N_2862,In_88,In_2049);
or U2863 (N_2863,In_1966,In_1988);
or U2864 (N_2864,In_1722,In_1925);
or U2865 (N_2865,In_314,In_556);
nor U2866 (N_2866,In_1254,In_2368);
nor U2867 (N_2867,In_1435,In_1256);
and U2868 (N_2868,In_547,In_12);
or U2869 (N_2869,In_453,In_1460);
nor U2870 (N_2870,In_2442,In_790);
nor U2871 (N_2871,In_741,In_2292);
nand U2872 (N_2872,In_2471,In_1128);
or U2873 (N_2873,In_80,In_973);
or U2874 (N_2874,In_335,In_1003);
nor U2875 (N_2875,In_1488,In_118);
or U2876 (N_2876,In_1222,In_813);
and U2877 (N_2877,In_14,In_1328);
nand U2878 (N_2878,In_2323,In_2149);
nor U2879 (N_2879,In_886,In_1998);
or U2880 (N_2880,In_2477,In_2087);
or U2881 (N_2881,In_1661,In_159);
xnor U2882 (N_2882,In_347,In_544);
or U2883 (N_2883,In_590,In_1149);
nor U2884 (N_2884,In_2144,In_1514);
and U2885 (N_2885,In_1689,In_658);
nand U2886 (N_2886,In_2428,In_2244);
nor U2887 (N_2887,In_1508,In_1114);
nor U2888 (N_2888,In_1381,In_88);
nand U2889 (N_2889,In_988,In_178);
nand U2890 (N_2890,In_1042,In_1544);
nor U2891 (N_2891,In_413,In_645);
nand U2892 (N_2892,In_622,In_398);
nand U2893 (N_2893,In_1105,In_1115);
or U2894 (N_2894,In_2128,In_1671);
nand U2895 (N_2895,In_137,In_887);
and U2896 (N_2896,In_1425,In_2087);
nand U2897 (N_2897,In_971,In_1655);
and U2898 (N_2898,In_1614,In_2134);
or U2899 (N_2899,In_2095,In_1376);
nor U2900 (N_2900,In_2193,In_2001);
and U2901 (N_2901,In_2449,In_1943);
or U2902 (N_2902,In_1568,In_2108);
nor U2903 (N_2903,In_986,In_806);
or U2904 (N_2904,In_1215,In_494);
nand U2905 (N_2905,In_926,In_2400);
nor U2906 (N_2906,In_864,In_533);
nand U2907 (N_2907,In_1306,In_383);
nand U2908 (N_2908,In_1722,In_261);
nor U2909 (N_2909,In_613,In_2252);
nor U2910 (N_2910,In_634,In_2000);
and U2911 (N_2911,In_2454,In_95);
nor U2912 (N_2912,In_1476,In_1333);
nor U2913 (N_2913,In_121,In_1417);
nor U2914 (N_2914,In_20,In_143);
or U2915 (N_2915,In_2271,In_1183);
nor U2916 (N_2916,In_1600,In_2401);
and U2917 (N_2917,In_1469,In_2495);
and U2918 (N_2918,In_276,In_2050);
xor U2919 (N_2919,In_985,In_389);
nand U2920 (N_2920,In_1785,In_377);
or U2921 (N_2921,In_433,In_110);
and U2922 (N_2922,In_2058,In_172);
and U2923 (N_2923,In_1314,In_548);
or U2924 (N_2924,In_612,In_2272);
nand U2925 (N_2925,In_1122,In_577);
nor U2926 (N_2926,In_444,In_1109);
and U2927 (N_2927,In_2228,In_1878);
or U2928 (N_2928,In_1794,In_706);
nand U2929 (N_2929,In_425,In_1796);
nand U2930 (N_2930,In_1652,In_805);
nand U2931 (N_2931,In_1489,In_954);
nand U2932 (N_2932,In_1930,In_1082);
or U2933 (N_2933,In_2142,In_2370);
and U2934 (N_2934,In_2436,In_2360);
nand U2935 (N_2935,In_583,In_445);
or U2936 (N_2936,In_2246,In_354);
nand U2937 (N_2937,In_1761,In_2017);
or U2938 (N_2938,In_1788,In_1921);
nor U2939 (N_2939,In_1644,In_850);
nor U2940 (N_2940,In_2063,In_1401);
or U2941 (N_2941,In_805,In_81);
or U2942 (N_2942,In_1890,In_1849);
or U2943 (N_2943,In_2396,In_44);
or U2944 (N_2944,In_418,In_590);
nand U2945 (N_2945,In_1495,In_1650);
nand U2946 (N_2946,In_610,In_1591);
nand U2947 (N_2947,In_1359,In_1886);
nand U2948 (N_2948,In_1345,In_1264);
nand U2949 (N_2949,In_2122,In_2366);
xnor U2950 (N_2950,In_1241,In_235);
xor U2951 (N_2951,In_2383,In_1229);
nor U2952 (N_2952,In_227,In_282);
or U2953 (N_2953,In_1790,In_382);
and U2954 (N_2954,In_816,In_369);
nor U2955 (N_2955,In_2404,In_1725);
or U2956 (N_2956,In_1505,In_1438);
and U2957 (N_2957,In_973,In_1284);
and U2958 (N_2958,In_123,In_2160);
and U2959 (N_2959,In_611,In_124);
nand U2960 (N_2960,In_1816,In_766);
and U2961 (N_2961,In_2196,In_795);
nor U2962 (N_2962,In_1401,In_1288);
and U2963 (N_2963,In_1238,In_1029);
xor U2964 (N_2964,In_377,In_2423);
or U2965 (N_2965,In_1830,In_1621);
nor U2966 (N_2966,In_1649,In_1168);
nand U2967 (N_2967,In_570,In_468);
nor U2968 (N_2968,In_276,In_1724);
or U2969 (N_2969,In_1513,In_829);
nand U2970 (N_2970,In_1783,In_903);
or U2971 (N_2971,In_2125,In_1773);
nand U2972 (N_2972,In_39,In_644);
or U2973 (N_2973,In_1489,In_2033);
and U2974 (N_2974,In_405,In_1842);
nor U2975 (N_2975,In_1159,In_1992);
nor U2976 (N_2976,In_404,In_145);
nand U2977 (N_2977,In_1599,In_1475);
xnor U2978 (N_2978,In_511,In_300);
nand U2979 (N_2979,In_806,In_1951);
nand U2980 (N_2980,In_791,In_1150);
or U2981 (N_2981,In_1784,In_433);
or U2982 (N_2982,In_681,In_617);
nand U2983 (N_2983,In_804,In_497);
or U2984 (N_2984,In_1439,In_2003);
nand U2985 (N_2985,In_692,In_2239);
nand U2986 (N_2986,In_302,In_268);
nor U2987 (N_2987,In_1691,In_2421);
nor U2988 (N_2988,In_2082,In_756);
and U2989 (N_2989,In_1772,In_629);
or U2990 (N_2990,In_1147,In_2193);
nand U2991 (N_2991,In_1581,In_2446);
and U2992 (N_2992,In_1681,In_1844);
nor U2993 (N_2993,In_824,In_184);
nor U2994 (N_2994,In_1601,In_290);
nand U2995 (N_2995,In_1988,In_2300);
nor U2996 (N_2996,In_913,In_1073);
or U2997 (N_2997,In_1957,In_2238);
nor U2998 (N_2998,In_1742,In_2462);
and U2999 (N_2999,In_307,In_1934);
nor U3000 (N_3000,In_1419,In_1444);
or U3001 (N_3001,In_465,In_1618);
or U3002 (N_3002,In_1003,In_1083);
or U3003 (N_3003,In_1421,In_190);
and U3004 (N_3004,In_75,In_1816);
xor U3005 (N_3005,In_2198,In_1168);
nand U3006 (N_3006,In_301,In_2330);
and U3007 (N_3007,In_856,In_1008);
and U3008 (N_3008,In_183,In_1731);
nand U3009 (N_3009,In_2237,In_1936);
or U3010 (N_3010,In_1219,In_2265);
or U3011 (N_3011,In_1275,In_1107);
xor U3012 (N_3012,In_1695,In_2361);
or U3013 (N_3013,In_2462,In_1192);
and U3014 (N_3014,In_1049,In_2260);
nor U3015 (N_3015,In_1301,In_803);
and U3016 (N_3016,In_2208,In_1930);
nand U3017 (N_3017,In_199,In_216);
or U3018 (N_3018,In_128,In_1148);
and U3019 (N_3019,In_197,In_1115);
nand U3020 (N_3020,In_798,In_1915);
nand U3021 (N_3021,In_430,In_1069);
nor U3022 (N_3022,In_143,In_265);
and U3023 (N_3023,In_1679,In_657);
and U3024 (N_3024,In_823,In_1948);
or U3025 (N_3025,In_903,In_320);
or U3026 (N_3026,In_1861,In_81);
and U3027 (N_3027,In_1248,In_1159);
nor U3028 (N_3028,In_554,In_1345);
nand U3029 (N_3029,In_2226,In_525);
or U3030 (N_3030,In_361,In_762);
nor U3031 (N_3031,In_1646,In_171);
nor U3032 (N_3032,In_2018,In_1301);
or U3033 (N_3033,In_711,In_821);
nor U3034 (N_3034,In_1133,In_1788);
nand U3035 (N_3035,In_813,In_708);
nor U3036 (N_3036,In_506,In_2473);
or U3037 (N_3037,In_28,In_142);
nor U3038 (N_3038,In_636,In_373);
xnor U3039 (N_3039,In_766,In_1908);
and U3040 (N_3040,In_1571,In_2311);
and U3041 (N_3041,In_2495,In_1181);
nor U3042 (N_3042,In_635,In_1570);
nor U3043 (N_3043,In_1564,In_1445);
or U3044 (N_3044,In_1254,In_1919);
and U3045 (N_3045,In_238,In_2024);
or U3046 (N_3046,In_641,In_2411);
nand U3047 (N_3047,In_1556,In_1678);
nand U3048 (N_3048,In_7,In_1741);
and U3049 (N_3049,In_107,In_2476);
nand U3050 (N_3050,In_1834,In_1925);
nand U3051 (N_3051,In_443,In_1774);
nor U3052 (N_3052,In_1215,In_539);
and U3053 (N_3053,In_500,In_154);
nand U3054 (N_3054,In_302,In_1399);
and U3055 (N_3055,In_1046,In_1502);
nor U3056 (N_3056,In_1681,In_688);
or U3057 (N_3057,In_1455,In_2356);
nor U3058 (N_3058,In_715,In_854);
and U3059 (N_3059,In_1978,In_1476);
or U3060 (N_3060,In_2003,In_798);
or U3061 (N_3061,In_934,In_210);
and U3062 (N_3062,In_778,In_138);
and U3063 (N_3063,In_918,In_1070);
nor U3064 (N_3064,In_571,In_1420);
nor U3065 (N_3065,In_596,In_592);
nor U3066 (N_3066,In_1610,In_1107);
xor U3067 (N_3067,In_582,In_2431);
or U3068 (N_3068,In_2446,In_1295);
nand U3069 (N_3069,In_983,In_1188);
nor U3070 (N_3070,In_687,In_1866);
and U3071 (N_3071,In_1623,In_207);
or U3072 (N_3072,In_114,In_1782);
nor U3073 (N_3073,In_1285,In_359);
or U3074 (N_3074,In_2262,In_1526);
nor U3075 (N_3075,In_2321,In_256);
and U3076 (N_3076,In_2400,In_1225);
nor U3077 (N_3077,In_1478,In_1512);
nor U3078 (N_3078,In_1916,In_589);
nor U3079 (N_3079,In_2107,In_1907);
nand U3080 (N_3080,In_1017,In_804);
nor U3081 (N_3081,In_1577,In_2455);
and U3082 (N_3082,In_1998,In_36);
and U3083 (N_3083,In_917,In_1715);
and U3084 (N_3084,In_488,In_829);
nor U3085 (N_3085,In_231,In_94);
and U3086 (N_3086,In_1281,In_1825);
or U3087 (N_3087,In_895,In_2402);
or U3088 (N_3088,In_603,In_2104);
nor U3089 (N_3089,In_1831,In_1382);
and U3090 (N_3090,In_1112,In_843);
nand U3091 (N_3091,In_1342,In_1985);
and U3092 (N_3092,In_2232,In_2164);
and U3093 (N_3093,In_1370,In_2254);
and U3094 (N_3094,In_1514,In_1541);
nand U3095 (N_3095,In_229,In_1370);
xnor U3096 (N_3096,In_881,In_870);
and U3097 (N_3097,In_1004,In_1413);
nand U3098 (N_3098,In_192,In_1806);
nor U3099 (N_3099,In_1895,In_366);
xor U3100 (N_3100,In_726,In_2116);
nor U3101 (N_3101,In_35,In_1465);
or U3102 (N_3102,In_1744,In_963);
nand U3103 (N_3103,In_2169,In_1231);
nor U3104 (N_3104,In_1743,In_1114);
nand U3105 (N_3105,In_1037,In_393);
or U3106 (N_3106,In_1670,In_1923);
or U3107 (N_3107,In_86,In_683);
nand U3108 (N_3108,In_274,In_451);
or U3109 (N_3109,In_901,In_2103);
and U3110 (N_3110,In_489,In_1203);
and U3111 (N_3111,In_2166,In_630);
or U3112 (N_3112,In_746,In_709);
or U3113 (N_3113,In_1600,In_511);
nand U3114 (N_3114,In_712,In_363);
nor U3115 (N_3115,In_1688,In_763);
nand U3116 (N_3116,In_2252,In_292);
nor U3117 (N_3117,In_2480,In_1901);
nor U3118 (N_3118,In_1261,In_1798);
nand U3119 (N_3119,In_1147,In_121);
nor U3120 (N_3120,In_1813,In_2282);
and U3121 (N_3121,In_1222,In_382);
and U3122 (N_3122,In_1092,In_892);
and U3123 (N_3123,In_1467,In_1280);
and U3124 (N_3124,In_1313,In_2374);
nor U3125 (N_3125,In_1023,In_1856);
nand U3126 (N_3126,In_2377,In_989);
or U3127 (N_3127,In_62,In_447);
or U3128 (N_3128,In_1709,In_699);
nand U3129 (N_3129,In_1434,In_525);
or U3130 (N_3130,In_175,In_1730);
nand U3131 (N_3131,In_1848,In_1775);
xnor U3132 (N_3132,In_2052,In_403);
nand U3133 (N_3133,In_783,In_1049);
nand U3134 (N_3134,In_1008,In_1847);
nor U3135 (N_3135,In_2402,In_1359);
and U3136 (N_3136,In_1410,In_2453);
and U3137 (N_3137,In_477,In_1164);
nand U3138 (N_3138,In_2297,In_1176);
nand U3139 (N_3139,In_812,In_1031);
nor U3140 (N_3140,In_1455,In_668);
and U3141 (N_3141,In_1636,In_320);
or U3142 (N_3142,In_616,In_2227);
nand U3143 (N_3143,In_1311,In_757);
nand U3144 (N_3144,In_1113,In_24);
nor U3145 (N_3145,In_1162,In_796);
nor U3146 (N_3146,In_1343,In_665);
and U3147 (N_3147,In_50,In_1326);
or U3148 (N_3148,In_2009,In_1485);
nand U3149 (N_3149,In_1409,In_1346);
nand U3150 (N_3150,In_612,In_482);
nor U3151 (N_3151,In_2428,In_1500);
nand U3152 (N_3152,In_1999,In_466);
and U3153 (N_3153,In_2209,In_2215);
or U3154 (N_3154,In_1492,In_809);
nor U3155 (N_3155,In_460,In_2046);
and U3156 (N_3156,In_752,In_547);
and U3157 (N_3157,In_2196,In_1735);
nor U3158 (N_3158,In_855,In_412);
nand U3159 (N_3159,In_408,In_1423);
and U3160 (N_3160,In_244,In_2009);
nor U3161 (N_3161,In_446,In_325);
or U3162 (N_3162,In_267,In_2294);
and U3163 (N_3163,In_797,In_2299);
nor U3164 (N_3164,In_1391,In_2097);
or U3165 (N_3165,In_514,In_2488);
nor U3166 (N_3166,In_1647,In_656);
nand U3167 (N_3167,In_597,In_575);
nand U3168 (N_3168,In_54,In_986);
or U3169 (N_3169,In_503,In_780);
nand U3170 (N_3170,In_1732,In_2229);
nand U3171 (N_3171,In_286,In_889);
and U3172 (N_3172,In_963,In_1253);
nand U3173 (N_3173,In_1215,In_193);
nor U3174 (N_3174,In_650,In_1448);
nand U3175 (N_3175,In_288,In_587);
or U3176 (N_3176,In_1450,In_1955);
and U3177 (N_3177,In_1593,In_637);
and U3178 (N_3178,In_1003,In_1022);
nand U3179 (N_3179,In_2062,In_764);
or U3180 (N_3180,In_1554,In_1993);
or U3181 (N_3181,In_1386,In_1023);
nor U3182 (N_3182,In_1179,In_1823);
and U3183 (N_3183,In_933,In_1080);
nand U3184 (N_3184,In_1858,In_835);
and U3185 (N_3185,In_1133,In_987);
nor U3186 (N_3186,In_39,In_1332);
and U3187 (N_3187,In_2101,In_527);
and U3188 (N_3188,In_1706,In_1572);
and U3189 (N_3189,In_1848,In_1285);
and U3190 (N_3190,In_1574,In_2030);
nand U3191 (N_3191,In_2390,In_2438);
or U3192 (N_3192,In_980,In_178);
nor U3193 (N_3193,In_136,In_1393);
or U3194 (N_3194,In_610,In_834);
and U3195 (N_3195,In_1472,In_703);
nand U3196 (N_3196,In_1227,In_2197);
nand U3197 (N_3197,In_1652,In_2483);
nand U3198 (N_3198,In_1009,In_2064);
or U3199 (N_3199,In_104,In_501);
or U3200 (N_3200,In_1205,In_2373);
or U3201 (N_3201,In_1599,In_1523);
and U3202 (N_3202,In_2095,In_2053);
nor U3203 (N_3203,In_2347,In_2091);
nor U3204 (N_3204,In_1809,In_111);
nor U3205 (N_3205,In_345,In_2346);
nand U3206 (N_3206,In_2454,In_1074);
nand U3207 (N_3207,In_1121,In_589);
and U3208 (N_3208,In_963,In_1920);
and U3209 (N_3209,In_1800,In_2288);
nand U3210 (N_3210,In_1903,In_2310);
and U3211 (N_3211,In_1615,In_5);
nand U3212 (N_3212,In_1494,In_2474);
nand U3213 (N_3213,In_951,In_522);
nand U3214 (N_3214,In_683,In_1490);
nor U3215 (N_3215,In_1662,In_1759);
or U3216 (N_3216,In_2484,In_1073);
or U3217 (N_3217,In_2452,In_2275);
and U3218 (N_3218,In_323,In_1383);
nor U3219 (N_3219,In_31,In_625);
nand U3220 (N_3220,In_1548,In_1804);
or U3221 (N_3221,In_825,In_873);
and U3222 (N_3222,In_2030,In_1628);
or U3223 (N_3223,In_180,In_1429);
or U3224 (N_3224,In_2139,In_112);
nand U3225 (N_3225,In_1732,In_2107);
nor U3226 (N_3226,In_7,In_1331);
and U3227 (N_3227,In_1955,In_802);
xor U3228 (N_3228,In_2266,In_1378);
and U3229 (N_3229,In_895,In_2493);
or U3230 (N_3230,In_1906,In_842);
nor U3231 (N_3231,In_2449,In_1855);
and U3232 (N_3232,In_2068,In_1692);
and U3233 (N_3233,In_706,In_479);
or U3234 (N_3234,In_2018,In_1871);
xor U3235 (N_3235,In_1325,In_890);
nor U3236 (N_3236,In_1434,In_953);
and U3237 (N_3237,In_2164,In_923);
xnor U3238 (N_3238,In_1711,In_1923);
nand U3239 (N_3239,In_1296,In_815);
nor U3240 (N_3240,In_1062,In_149);
nand U3241 (N_3241,In_1161,In_2482);
nand U3242 (N_3242,In_482,In_5);
or U3243 (N_3243,In_2171,In_1957);
nand U3244 (N_3244,In_2320,In_2060);
nand U3245 (N_3245,In_847,In_2115);
nor U3246 (N_3246,In_1585,In_946);
nor U3247 (N_3247,In_1571,In_2179);
and U3248 (N_3248,In_1595,In_2323);
nand U3249 (N_3249,In_750,In_472);
nand U3250 (N_3250,In_1448,In_2188);
or U3251 (N_3251,In_1469,In_1502);
and U3252 (N_3252,In_759,In_970);
xor U3253 (N_3253,In_1684,In_719);
nand U3254 (N_3254,In_2257,In_1074);
and U3255 (N_3255,In_2325,In_923);
or U3256 (N_3256,In_957,In_2357);
nand U3257 (N_3257,In_1291,In_459);
nor U3258 (N_3258,In_1855,In_2410);
or U3259 (N_3259,In_282,In_1051);
nand U3260 (N_3260,In_47,In_2013);
nor U3261 (N_3261,In_1847,In_831);
or U3262 (N_3262,In_260,In_1376);
or U3263 (N_3263,In_445,In_2031);
and U3264 (N_3264,In_218,In_2399);
and U3265 (N_3265,In_97,In_2027);
or U3266 (N_3266,In_2445,In_1058);
or U3267 (N_3267,In_1944,In_963);
and U3268 (N_3268,In_133,In_643);
nor U3269 (N_3269,In_2208,In_1759);
or U3270 (N_3270,In_1548,In_1234);
nor U3271 (N_3271,In_1446,In_842);
or U3272 (N_3272,In_948,In_929);
nand U3273 (N_3273,In_746,In_2496);
nor U3274 (N_3274,In_170,In_1861);
and U3275 (N_3275,In_1905,In_1138);
and U3276 (N_3276,In_898,In_1691);
nor U3277 (N_3277,In_934,In_1478);
nor U3278 (N_3278,In_2364,In_2188);
nand U3279 (N_3279,In_443,In_1020);
and U3280 (N_3280,In_196,In_2292);
nor U3281 (N_3281,In_388,In_2296);
nor U3282 (N_3282,In_273,In_482);
nand U3283 (N_3283,In_184,In_2080);
or U3284 (N_3284,In_2324,In_1837);
and U3285 (N_3285,In_927,In_1252);
nand U3286 (N_3286,In_1466,In_1954);
and U3287 (N_3287,In_1157,In_244);
nand U3288 (N_3288,In_855,In_328);
nor U3289 (N_3289,In_2207,In_93);
or U3290 (N_3290,In_1098,In_1699);
or U3291 (N_3291,In_897,In_283);
or U3292 (N_3292,In_1904,In_679);
nor U3293 (N_3293,In_297,In_778);
nor U3294 (N_3294,In_1444,In_2062);
nand U3295 (N_3295,In_1796,In_109);
nand U3296 (N_3296,In_724,In_1767);
nor U3297 (N_3297,In_54,In_1607);
or U3298 (N_3298,In_2465,In_1576);
or U3299 (N_3299,In_2333,In_2482);
or U3300 (N_3300,In_291,In_984);
or U3301 (N_3301,In_1667,In_1910);
and U3302 (N_3302,In_325,In_1800);
and U3303 (N_3303,In_1388,In_1578);
and U3304 (N_3304,In_2317,In_1308);
nor U3305 (N_3305,In_62,In_572);
nand U3306 (N_3306,In_1396,In_2461);
or U3307 (N_3307,In_2025,In_1869);
nand U3308 (N_3308,In_2017,In_2310);
nor U3309 (N_3309,In_1061,In_986);
nor U3310 (N_3310,In_613,In_1534);
nor U3311 (N_3311,In_607,In_536);
nor U3312 (N_3312,In_1015,In_1793);
or U3313 (N_3313,In_35,In_1196);
nor U3314 (N_3314,In_820,In_2049);
or U3315 (N_3315,In_1852,In_2172);
nand U3316 (N_3316,In_404,In_914);
and U3317 (N_3317,In_1015,In_1618);
and U3318 (N_3318,In_1778,In_2447);
or U3319 (N_3319,In_397,In_1879);
nand U3320 (N_3320,In_1123,In_1933);
nor U3321 (N_3321,In_1910,In_1739);
or U3322 (N_3322,In_1652,In_2453);
nor U3323 (N_3323,In_1980,In_434);
and U3324 (N_3324,In_19,In_1307);
nand U3325 (N_3325,In_106,In_1783);
nor U3326 (N_3326,In_536,In_331);
nor U3327 (N_3327,In_297,In_883);
or U3328 (N_3328,In_110,In_1665);
nand U3329 (N_3329,In_1944,In_1618);
and U3330 (N_3330,In_2482,In_1557);
or U3331 (N_3331,In_252,In_1987);
and U3332 (N_3332,In_2166,In_2102);
nor U3333 (N_3333,In_483,In_1019);
or U3334 (N_3334,In_1787,In_414);
nand U3335 (N_3335,In_629,In_678);
nor U3336 (N_3336,In_1447,In_2203);
or U3337 (N_3337,In_129,In_1377);
and U3338 (N_3338,In_272,In_1828);
nor U3339 (N_3339,In_621,In_622);
and U3340 (N_3340,In_1035,In_546);
nand U3341 (N_3341,In_2449,In_1700);
and U3342 (N_3342,In_444,In_1997);
nand U3343 (N_3343,In_952,In_1219);
nor U3344 (N_3344,In_1516,In_774);
nor U3345 (N_3345,In_699,In_1660);
and U3346 (N_3346,In_902,In_2018);
and U3347 (N_3347,In_2282,In_956);
and U3348 (N_3348,In_983,In_1654);
nor U3349 (N_3349,In_1433,In_1676);
nand U3350 (N_3350,In_771,In_1770);
nand U3351 (N_3351,In_849,In_2033);
nand U3352 (N_3352,In_1243,In_1397);
or U3353 (N_3353,In_1083,In_483);
nand U3354 (N_3354,In_631,In_1479);
and U3355 (N_3355,In_1609,In_219);
and U3356 (N_3356,In_850,In_573);
nand U3357 (N_3357,In_1467,In_646);
nand U3358 (N_3358,In_245,In_1397);
nand U3359 (N_3359,In_1209,In_466);
nand U3360 (N_3360,In_265,In_2009);
or U3361 (N_3361,In_922,In_541);
and U3362 (N_3362,In_1587,In_618);
nand U3363 (N_3363,In_7,In_1812);
and U3364 (N_3364,In_2292,In_2148);
nor U3365 (N_3365,In_2275,In_1524);
and U3366 (N_3366,In_892,In_241);
nor U3367 (N_3367,In_2348,In_1741);
and U3368 (N_3368,In_1654,In_1692);
nand U3369 (N_3369,In_1906,In_1268);
xnor U3370 (N_3370,In_68,In_1220);
or U3371 (N_3371,In_2273,In_440);
nor U3372 (N_3372,In_701,In_1945);
nand U3373 (N_3373,In_1422,In_910);
nand U3374 (N_3374,In_643,In_2016);
nand U3375 (N_3375,In_1049,In_632);
or U3376 (N_3376,In_1798,In_1263);
or U3377 (N_3377,In_617,In_1835);
nand U3378 (N_3378,In_828,In_421);
and U3379 (N_3379,In_116,In_59);
or U3380 (N_3380,In_366,In_848);
or U3381 (N_3381,In_2228,In_1038);
and U3382 (N_3382,In_160,In_1557);
nand U3383 (N_3383,In_2295,In_2103);
or U3384 (N_3384,In_769,In_1219);
or U3385 (N_3385,In_992,In_855);
nor U3386 (N_3386,In_1644,In_2091);
and U3387 (N_3387,In_1272,In_324);
nand U3388 (N_3388,In_1150,In_391);
nor U3389 (N_3389,In_1499,In_1705);
nor U3390 (N_3390,In_1436,In_2065);
and U3391 (N_3391,In_1456,In_2049);
nor U3392 (N_3392,In_1934,In_1347);
nand U3393 (N_3393,In_402,In_1927);
or U3394 (N_3394,In_738,In_535);
or U3395 (N_3395,In_545,In_846);
nor U3396 (N_3396,In_677,In_1113);
and U3397 (N_3397,In_1415,In_2427);
nor U3398 (N_3398,In_893,In_220);
xnor U3399 (N_3399,In_10,In_1118);
nor U3400 (N_3400,In_355,In_2101);
and U3401 (N_3401,In_1855,In_255);
nand U3402 (N_3402,In_537,In_1235);
nand U3403 (N_3403,In_470,In_943);
and U3404 (N_3404,In_223,In_1203);
and U3405 (N_3405,In_1536,In_2475);
or U3406 (N_3406,In_1937,In_661);
nor U3407 (N_3407,In_2317,In_1604);
and U3408 (N_3408,In_1241,In_1929);
and U3409 (N_3409,In_1890,In_630);
nor U3410 (N_3410,In_864,In_726);
and U3411 (N_3411,In_301,In_1941);
and U3412 (N_3412,In_618,In_186);
or U3413 (N_3413,In_2007,In_364);
nor U3414 (N_3414,In_1131,In_2304);
nand U3415 (N_3415,In_289,In_466);
nor U3416 (N_3416,In_2052,In_1633);
nor U3417 (N_3417,In_383,In_789);
or U3418 (N_3418,In_747,In_164);
or U3419 (N_3419,In_997,In_1135);
and U3420 (N_3420,In_1008,In_1188);
nor U3421 (N_3421,In_59,In_1652);
and U3422 (N_3422,In_1196,In_441);
and U3423 (N_3423,In_556,In_1209);
nor U3424 (N_3424,In_1067,In_486);
nand U3425 (N_3425,In_1662,In_2239);
or U3426 (N_3426,In_55,In_1651);
and U3427 (N_3427,In_1268,In_2262);
and U3428 (N_3428,In_85,In_1601);
nand U3429 (N_3429,In_1078,In_1970);
nor U3430 (N_3430,In_10,In_1653);
and U3431 (N_3431,In_986,In_2271);
or U3432 (N_3432,In_2369,In_2185);
nor U3433 (N_3433,In_340,In_1907);
and U3434 (N_3434,In_1690,In_1178);
nor U3435 (N_3435,In_2179,In_1919);
or U3436 (N_3436,In_1292,In_7);
and U3437 (N_3437,In_2060,In_637);
nand U3438 (N_3438,In_1136,In_96);
and U3439 (N_3439,In_2169,In_883);
nor U3440 (N_3440,In_43,In_1264);
nand U3441 (N_3441,In_1670,In_1634);
xnor U3442 (N_3442,In_1471,In_2215);
nor U3443 (N_3443,In_645,In_1321);
and U3444 (N_3444,In_1319,In_1038);
and U3445 (N_3445,In_922,In_2383);
nor U3446 (N_3446,In_102,In_2495);
or U3447 (N_3447,In_577,In_2447);
and U3448 (N_3448,In_2187,In_199);
or U3449 (N_3449,In_714,In_428);
nor U3450 (N_3450,In_1127,In_980);
nand U3451 (N_3451,In_603,In_588);
or U3452 (N_3452,In_1421,In_2436);
nor U3453 (N_3453,In_2030,In_700);
or U3454 (N_3454,In_1348,In_1938);
and U3455 (N_3455,In_2367,In_1417);
nand U3456 (N_3456,In_2172,In_707);
nand U3457 (N_3457,In_215,In_790);
or U3458 (N_3458,In_214,In_2351);
and U3459 (N_3459,In_2297,In_2432);
or U3460 (N_3460,In_847,In_307);
and U3461 (N_3461,In_95,In_1791);
nor U3462 (N_3462,In_231,In_2348);
xnor U3463 (N_3463,In_41,In_1955);
and U3464 (N_3464,In_1787,In_2335);
nor U3465 (N_3465,In_2457,In_326);
and U3466 (N_3466,In_1604,In_568);
and U3467 (N_3467,In_613,In_1477);
or U3468 (N_3468,In_2279,In_1202);
or U3469 (N_3469,In_119,In_692);
and U3470 (N_3470,In_438,In_2010);
or U3471 (N_3471,In_1341,In_1117);
nor U3472 (N_3472,In_2197,In_1980);
xnor U3473 (N_3473,In_1799,In_1915);
or U3474 (N_3474,In_1279,In_2314);
and U3475 (N_3475,In_1522,In_1323);
nand U3476 (N_3476,In_2235,In_1235);
and U3477 (N_3477,In_811,In_322);
xnor U3478 (N_3478,In_524,In_1619);
nor U3479 (N_3479,In_2235,In_1984);
nand U3480 (N_3480,In_1792,In_1660);
nand U3481 (N_3481,In_2222,In_490);
and U3482 (N_3482,In_1939,In_807);
and U3483 (N_3483,In_2423,In_1101);
nor U3484 (N_3484,In_120,In_481);
or U3485 (N_3485,In_2072,In_192);
nand U3486 (N_3486,In_897,In_242);
nand U3487 (N_3487,In_1329,In_1909);
and U3488 (N_3488,In_2086,In_595);
nor U3489 (N_3489,In_2468,In_1678);
and U3490 (N_3490,In_2267,In_1984);
nor U3491 (N_3491,In_1337,In_2462);
nand U3492 (N_3492,In_1204,In_1997);
nand U3493 (N_3493,In_115,In_1694);
nand U3494 (N_3494,In_989,In_1861);
nand U3495 (N_3495,In_1106,In_1762);
nand U3496 (N_3496,In_1851,In_1325);
and U3497 (N_3497,In_774,In_306);
xor U3498 (N_3498,In_1064,In_2030);
nand U3499 (N_3499,In_1985,In_2288);
nor U3500 (N_3500,In_1053,In_2473);
or U3501 (N_3501,In_1344,In_540);
nor U3502 (N_3502,In_1126,In_1174);
nand U3503 (N_3503,In_852,In_553);
nand U3504 (N_3504,In_633,In_1339);
or U3505 (N_3505,In_1773,In_1539);
nor U3506 (N_3506,In_694,In_543);
nor U3507 (N_3507,In_1941,In_2206);
or U3508 (N_3508,In_1302,In_1024);
nor U3509 (N_3509,In_193,In_2286);
and U3510 (N_3510,In_1897,In_1435);
and U3511 (N_3511,In_1250,In_80);
or U3512 (N_3512,In_2317,In_644);
nand U3513 (N_3513,In_1806,In_2030);
nand U3514 (N_3514,In_1427,In_1414);
and U3515 (N_3515,In_1553,In_1613);
nor U3516 (N_3516,In_874,In_1409);
nor U3517 (N_3517,In_1364,In_1708);
nand U3518 (N_3518,In_2325,In_2150);
and U3519 (N_3519,In_1228,In_558);
nor U3520 (N_3520,In_1620,In_187);
and U3521 (N_3521,In_1148,In_1921);
nor U3522 (N_3522,In_551,In_1882);
nor U3523 (N_3523,In_1262,In_33);
and U3524 (N_3524,In_420,In_971);
and U3525 (N_3525,In_2150,In_2219);
nor U3526 (N_3526,In_1918,In_775);
xnor U3527 (N_3527,In_1204,In_1604);
nand U3528 (N_3528,In_328,In_9);
nor U3529 (N_3529,In_466,In_1546);
or U3530 (N_3530,In_1949,In_1883);
nand U3531 (N_3531,In_2103,In_2408);
nand U3532 (N_3532,In_1683,In_2476);
nand U3533 (N_3533,In_1377,In_1013);
nand U3534 (N_3534,In_307,In_1385);
nand U3535 (N_3535,In_1867,In_108);
nand U3536 (N_3536,In_2340,In_2190);
or U3537 (N_3537,In_485,In_1963);
or U3538 (N_3538,In_2363,In_1538);
nor U3539 (N_3539,In_1466,In_1083);
or U3540 (N_3540,In_817,In_2347);
or U3541 (N_3541,In_2300,In_1900);
and U3542 (N_3542,In_708,In_2179);
or U3543 (N_3543,In_1702,In_472);
nand U3544 (N_3544,In_1681,In_882);
xor U3545 (N_3545,In_1684,In_901);
and U3546 (N_3546,In_2341,In_1667);
and U3547 (N_3547,In_332,In_1779);
nand U3548 (N_3548,In_435,In_1519);
nand U3549 (N_3549,In_115,In_678);
nand U3550 (N_3550,In_675,In_2272);
nor U3551 (N_3551,In_2058,In_2336);
or U3552 (N_3552,In_439,In_1016);
and U3553 (N_3553,In_2163,In_834);
or U3554 (N_3554,In_561,In_825);
and U3555 (N_3555,In_1481,In_1443);
and U3556 (N_3556,In_1463,In_1239);
or U3557 (N_3557,In_2123,In_1002);
nand U3558 (N_3558,In_1935,In_1698);
nor U3559 (N_3559,In_96,In_1770);
and U3560 (N_3560,In_26,In_1898);
or U3561 (N_3561,In_1946,In_542);
and U3562 (N_3562,In_503,In_1283);
or U3563 (N_3563,In_1736,In_1555);
and U3564 (N_3564,In_739,In_1381);
and U3565 (N_3565,In_955,In_1285);
nor U3566 (N_3566,In_422,In_536);
nor U3567 (N_3567,In_1071,In_2013);
or U3568 (N_3568,In_132,In_390);
or U3569 (N_3569,In_1680,In_354);
and U3570 (N_3570,In_1398,In_2220);
xnor U3571 (N_3571,In_803,In_1390);
or U3572 (N_3572,In_2440,In_2045);
or U3573 (N_3573,In_1523,In_1292);
nor U3574 (N_3574,In_1338,In_2026);
and U3575 (N_3575,In_422,In_210);
or U3576 (N_3576,In_1201,In_655);
nor U3577 (N_3577,In_1652,In_1494);
or U3578 (N_3578,In_1916,In_2285);
and U3579 (N_3579,In_540,In_2270);
nor U3580 (N_3580,In_1420,In_1750);
nor U3581 (N_3581,In_1422,In_1322);
and U3582 (N_3582,In_377,In_1888);
nor U3583 (N_3583,In_526,In_402);
nor U3584 (N_3584,In_87,In_269);
nand U3585 (N_3585,In_1012,In_367);
nand U3586 (N_3586,In_80,In_200);
and U3587 (N_3587,In_1778,In_1122);
and U3588 (N_3588,In_1598,In_1052);
or U3589 (N_3589,In_60,In_1214);
nand U3590 (N_3590,In_1141,In_2012);
nand U3591 (N_3591,In_2444,In_2099);
and U3592 (N_3592,In_392,In_2128);
nand U3593 (N_3593,In_1184,In_756);
nor U3594 (N_3594,In_1187,In_671);
nor U3595 (N_3595,In_1905,In_2000);
or U3596 (N_3596,In_473,In_2338);
and U3597 (N_3597,In_1857,In_504);
and U3598 (N_3598,In_2346,In_2246);
nor U3599 (N_3599,In_722,In_384);
nand U3600 (N_3600,In_1802,In_291);
nor U3601 (N_3601,In_1288,In_1070);
and U3602 (N_3602,In_2055,In_1857);
or U3603 (N_3603,In_1870,In_1413);
nor U3604 (N_3604,In_337,In_192);
nand U3605 (N_3605,In_85,In_1960);
or U3606 (N_3606,In_1731,In_559);
and U3607 (N_3607,In_1003,In_626);
and U3608 (N_3608,In_2353,In_307);
nor U3609 (N_3609,In_2357,In_729);
nand U3610 (N_3610,In_627,In_1391);
nand U3611 (N_3611,In_1335,In_1205);
and U3612 (N_3612,In_625,In_92);
nor U3613 (N_3613,In_2287,In_495);
nand U3614 (N_3614,In_1378,In_1614);
nor U3615 (N_3615,In_946,In_1052);
or U3616 (N_3616,In_495,In_1947);
and U3617 (N_3617,In_40,In_953);
or U3618 (N_3618,In_397,In_1276);
nand U3619 (N_3619,In_2109,In_397);
xor U3620 (N_3620,In_827,In_1710);
nand U3621 (N_3621,In_48,In_37);
nor U3622 (N_3622,In_2122,In_1782);
or U3623 (N_3623,In_1579,In_1667);
nand U3624 (N_3624,In_1709,In_2135);
or U3625 (N_3625,In_2208,In_1394);
and U3626 (N_3626,In_790,In_2097);
and U3627 (N_3627,In_1113,In_1831);
nor U3628 (N_3628,In_55,In_319);
and U3629 (N_3629,In_2196,In_381);
nor U3630 (N_3630,In_717,In_1198);
nand U3631 (N_3631,In_913,In_580);
nand U3632 (N_3632,In_1817,In_947);
or U3633 (N_3633,In_2038,In_1726);
and U3634 (N_3634,In_595,In_1133);
and U3635 (N_3635,In_2476,In_444);
nor U3636 (N_3636,In_495,In_2135);
nand U3637 (N_3637,In_2254,In_1022);
nor U3638 (N_3638,In_250,In_1094);
or U3639 (N_3639,In_2419,In_749);
nand U3640 (N_3640,In_990,In_2023);
nor U3641 (N_3641,In_1374,In_1531);
and U3642 (N_3642,In_2372,In_3);
or U3643 (N_3643,In_1,In_1091);
and U3644 (N_3644,In_514,In_2081);
and U3645 (N_3645,In_688,In_1366);
or U3646 (N_3646,In_2372,In_1655);
xnor U3647 (N_3647,In_1241,In_447);
nor U3648 (N_3648,In_1806,In_1177);
nand U3649 (N_3649,In_1330,In_158);
and U3650 (N_3650,In_1805,In_269);
or U3651 (N_3651,In_1066,In_2477);
nor U3652 (N_3652,In_1650,In_2259);
nor U3653 (N_3653,In_874,In_962);
or U3654 (N_3654,In_1535,In_2400);
nand U3655 (N_3655,In_1497,In_1081);
or U3656 (N_3656,In_2349,In_2438);
nand U3657 (N_3657,In_1070,In_261);
and U3658 (N_3658,In_2208,In_1236);
nand U3659 (N_3659,In_1153,In_1117);
and U3660 (N_3660,In_2442,In_692);
and U3661 (N_3661,In_1154,In_1668);
xor U3662 (N_3662,In_2481,In_171);
nand U3663 (N_3663,In_1822,In_574);
or U3664 (N_3664,In_283,In_1064);
or U3665 (N_3665,In_260,In_546);
nor U3666 (N_3666,In_2257,In_655);
nand U3667 (N_3667,In_426,In_1604);
or U3668 (N_3668,In_2327,In_1281);
nor U3669 (N_3669,In_2305,In_494);
nor U3670 (N_3670,In_1639,In_661);
nand U3671 (N_3671,In_1461,In_1884);
or U3672 (N_3672,In_1044,In_1501);
or U3673 (N_3673,In_2334,In_355);
and U3674 (N_3674,In_1641,In_2244);
nand U3675 (N_3675,In_19,In_2322);
nand U3676 (N_3676,In_521,In_1902);
nor U3677 (N_3677,In_1761,In_1994);
nand U3678 (N_3678,In_1871,In_740);
nor U3679 (N_3679,In_1923,In_20);
nand U3680 (N_3680,In_2445,In_1888);
and U3681 (N_3681,In_2263,In_82);
nor U3682 (N_3682,In_1590,In_1475);
nor U3683 (N_3683,In_405,In_785);
xnor U3684 (N_3684,In_305,In_355);
nor U3685 (N_3685,In_1029,In_2033);
and U3686 (N_3686,In_1135,In_911);
nor U3687 (N_3687,In_1397,In_315);
nand U3688 (N_3688,In_1440,In_997);
or U3689 (N_3689,In_1958,In_1950);
or U3690 (N_3690,In_610,In_619);
nor U3691 (N_3691,In_935,In_124);
nand U3692 (N_3692,In_1701,In_447);
nand U3693 (N_3693,In_863,In_2492);
nand U3694 (N_3694,In_1595,In_1764);
and U3695 (N_3695,In_2262,In_2107);
and U3696 (N_3696,In_143,In_934);
and U3697 (N_3697,In_1691,In_909);
or U3698 (N_3698,In_883,In_1594);
and U3699 (N_3699,In_1841,In_1260);
nand U3700 (N_3700,In_542,In_1181);
or U3701 (N_3701,In_1570,In_1914);
nor U3702 (N_3702,In_665,In_2395);
nor U3703 (N_3703,In_1549,In_1461);
nor U3704 (N_3704,In_127,In_2292);
and U3705 (N_3705,In_2252,In_2347);
or U3706 (N_3706,In_810,In_1204);
and U3707 (N_3707,In_1467,In_476);
or U3708 (N_3708,In_95,In_1647);
nand U3709 (N_3709,In_655,In_45);
and U3710 (N_3710,In_942,In_2434);
xor U3711 (N_3711,In_1178,In_1060);
nor U3712 (N_3712,In_731,In_1239);
and U3713 (N_3713,In_1437,In_567);
nor U3714 (N_3714,In_1036,In_2127);
nor U3715 (N_3715,In_497,In_1385);
nand U3716 (N_3716,In_2363,In_1179);
nor U3717 (N_3717,In_1267,In_2409);
and U3718 (N_3718,In_1017,In_1666);
nand U3719 (N_3719,In_386,In_2290);
or U3720 (N_3720,In_1468,In_1584);
and U3721 (N_3721,In_339,In_1183);
and U3722 (N_3722,In_596,In_1905);
nand U3723 (N_3723,In_2400,In_681);
nor U3724 (N_3724,In_2318,In_1361);
nand U3725 (N_3725,In_2319,In_2405);
and U3726 (N_3726,In_1118,In_669);
and U3727 (N_3727,In_2482,In_2070);
or U3728 (N_3728,In_1452,In_1260);
or U3729 (N_3729,In_1883,In_317);
nand U3730 (N_3730,In_270,In_443);
and U3731 (N_3731,In_221,In_53);
and U3732 (N_3732,In_1280,In_190);
nand U3733 (N_3733,In_2379,In_2363);
nand U3734 (N_3734,In_2425,In_1103);
nand U3735 (N_3735,In_2322,In_1897);
xor U3736 (N_3736,In_391,In_1054);
and U3737 (N_3737,In_749,In_248);
xnor U3738 (N_3738,In_2465,In_1245);
nor U3739 (N_3739,In_1939,In_1743);
and U3740 (N_3740,In_129,In_2074);
nor U3741 (N_3741,In_1056,In_1633);
or U3742 (N_3742,In_471,In_2281);
nand U3743 (N_3743,In_1492,In_65);
nor U3744 (N_3744,In_2391,In_934);
or U3745 (N_3745,In_1052,In_699);
nand U3746 (N_3746,In_30,In_465);
nand U3747 (N_3747,In_1905,In_1080);
or U3748 (N_3748,In_428,In_1462);
or U3749 (N_3749,In_1578,In_381);
or U3750 (N_3750,In_722,In_1661);
nor U3751 (N_3751,In_624,In_2214);
nor U3752 (N_3752,In_867,In_2135);
and U3753 (N_3753,In_1107,In_837);
and U3754 (N_3754,In_415,In_2010);
nand U3755 (N_3755,In_832,In_2378);
and U3756 (N_3756,In_1378,In_1480);
nand U3757 (N_3757,In_1745,In_965);
or U3758 (N_3758,In_1967,In_1631);
xnor U3759 (N_3759,In_2105,In_717);
and U3760 (N_3760,In_1840,In_2250);
and U3761 (N_3761,In_696,In_1809);
or U3762 (N_3762,In_2422,In_1744);
or U3763 (N_3763,In_2153,In_910);
nand U3764 (N_3764,In_2024,In_2388);
or U3765 (N_3765,In_1631,In_2435);
nand U3766 (N_3766,In_2496,In_591);
and U3767 (N_3767,In_1985,In_1313);
and U3768 (N_3768,In_938,In_2020);
or U3769 (N_3769,In_2295,In_517);
nand U3770 (N_3770,In_476,In_140);
or U3771 (N_3771,In_1861,In_1515);
and U3772 (N_3772,In_252,In_1670);
and U3773 (N_3773,In_138,In_1821);
nor U3774 (N_3774,In_1344,In_2499);
or U3775 (N_3775,In_90,In_2166);
and U3776 (N_3776,In_487,In_1547);
nor U3777 (N_3777,In_101,In_762);
and U3778 (N_3778,In_1795,In_1629);
nor U3779 (N_3779,In_460,In_134);
and U3780 (N_3780,In_2040,In_254);
nor U3781 (N_3781,In_923,In_1545);
nor U3782 (N_3782,In_1760,In_134);
nor U3783 (N_3783,In_911,In_36);
or U3784 (N_3784,In_630,In_1715);
or U3785 (N_3785,In_2033,In_58);
nand U3786 (N_3786,In_1429,In_1650);
nand U3787 (N_3787,In_642,In_1436);
nand U3788 (N_3788,In_1362,In_1142);
or U3789 (N_3789,In_169,In_1973);
xnor U3790 (N_3790,In_1384,In_2028);
and U3791 (N_3791,In_2186,In_1486);
or U3792 (N_3792,In_165,In_677);
nand U3793 (N_3793,In_302,In_1480);
nand U3794 (N_3794,In_2251,In_1446);
and U3795 (N_3795,In_572,In_941);
nand U3796 (N_3796,In_1878,In_2127);
nor U3797 (N_3797,In_2343,In_1996);
nor U3798 (N_3798,In_2354,In_397);
and U3799 (N_3799,In_962,In_373);
and U3800 (N_3800,In_1904,In_2462);
or U3801 (N_3801,In_781,In_1942);
xor U3802 (N_3802,In_1548,In_93);
or U3803 (N_3803,In_1229,In_1343);
or U3804 (N_3804,In_1587,In_1773);
xnor U3805 (N_3805,In_105,In_2287);
nand U3806 (N_3806,In_572,In_537);
nand U3807 (N_3807,In_2485,In_1017);
nand U3808 (N_3808,In_1653,In_1761);
nand U3809 (N_3809,In_238,In_462);
nor U3810 (N_3810,In_1105,In_59);
xnor U3811 (N_3811,In_2465,In_1151);
nor U3812 (N_3812,In_601,In_1765);
nand U3813 (N_3813,In_98,In_303);
nand U3814 (N_3814,In_2352,In_1677);
nand U3815 (N_3815,In_2327,In_682);
or U3816 (N_3816,In_899,In_1347);
and U3817 (N_3817,In_1604,In_2383);
xnor U3818 (N_3818,In_144,In_106);
or U3819 (N_3819,In_862,In_1798);
nor U3820 (N_3820,In_1015,In_1635);
nand U3821 (N_3821,In_2374,In_1264);
nor U3822 (N_3822,In_487,In_2476);
or U3823 (N_3823,In_1477,In_403);
or U3824 (N_3824,In_900,In_2145);
or U3825 (N_3825,In_714,In_589);
or U3826 (N_3826,In_2393,In_2314);
nand U3827 (N_3827,In_1997,In_1413);
or U3828 (N_3828,In_1136,In_623);
or U3829 (N_3829,In_612,In_345);
or U3830 (N_3830,In_588,In_2127);
and U3831 (N_3831,In_2050,In_1718);
and U3832 (N_3832,In_1411,In_1753);
xnor U3833 (N_3833,In_1396,In_2246);
nand U3834 (N_3834,In_1884,In_221);
nor U3835 (N_3835,In_134,In_967);
or U3836 (N_3836,In_679,In_2337);
nand U3837 (N_3837,In_1366,In_1171);
nand U3838 (N_3838,In_1087,In_437);
and U3839 (N_3839,In_2416,In_1479);
nor U3840 (N_3840,In_1623,In_1556);
and U3841 (N_3841,In_1848,In_2291);
and U3842 (N_3842,In_654,In_950);
or U3843 (N_3843,In_1665,In_925);
or U3844 (N_3844,In_2292,In_519);
and U3845 (N_3845,In_2273,In_1056);
and U3846 (N_3846,In_92,In_1526);
nand U3847 (N_3847,In_1055,In_2231);
or U3848 (N_3848,In_1318,In_366);
nor U3849 (N_3849,In_2199,In_1496);
and U3850 (N_3850,In_1508,In_1163);
nand U3851 (N_3851,In_1019,In_1690);
nand U3852 (N_3852,In_989,In_2118);
nor U3853 (N_3853,In_1207,In_2124);
or U3854 (N_3854,In_2,In_2180);
and U3855 (N_3855,In_1695,In_153);
nor U3856 (N_3856,In_1292,In_953);
nand U3857 (N_3857,In_2146,In_1497);
and U3858 (N_3858,In_26,In_1232);
nand U3859 (N_3859,In_261,In_1053);
or U3860 (N_3860,In_230,In_1867);
nor U3861 (N_3861,In_373,In_430);
nand U3862 (N_3862,In_2240,In_1738);
and U3863 (N_3863,In_1206,In_2237);
nand U3864 (N_3864,In_114,In_536);
and U3865 (N_3865,In_1462,In_1366);
or U3866 (N_3866,In_546,In_1963);
nand U3867 (N_3867,In_902,In_1569);
nand U3868 (N_3868,In_2156,In_2244);
and U3869 (N_3869,In_427,In_1764);
nor U3870 (N_3870,In_655,In_270);
nor U3871 (N_3871,In_2300,In_2116);
nor U3872 (N_3872,In_744,In_2432);
and U3873 (N_3873,In_1851,In_641);
nand U3874 (N_3874,In_2089,In_1964);
and U3875 (N_3875,In_2203,In_1277);
nor U3876 (N_3876,In_1255,In_1858);
and U3877 (N_3877,In_338,In_422);
xnor U3878 (N_3878,In_803,In_844);
nand U3879 (N_3879,In_799,In_854);
and U3880 (N_3880,In_2370,In_1734);
and U3881 (N_3881,In_1688,In_80);
and U3882 (N_3882,In_1258,In_1666);
nand U3883 (N_3883,In_1305,In_179);
nand U3884 (N_3884,In_305,In_1013);
and U3885 (N_3885,In_1780,In_749);
and U3886 (N_3886,In_1435,In_374);
or U3887 (N_3887,In_1005,In_171);
and U3888 (N_3888,In_73,In_2313);
and U3889 (N_3889,In_806,In_516);
nor U3890 (N_3890,In_1719,In_1127);
and U3891 (N_3891,In_794,In_28);
nor U3892 (N_3892,In_943,In_993);
or U3893 (N_3893,In_160,In_56);
nor U3894 (N_3894,In_595,In_366);
nor U3895 (N_3895,In_1247,In_1251);
nor U3896 (N_3896,In_1313,In_35);
nor U3897 (N_3897,In_342,In_776);
or U3898 (N_3898,In_1849,In_417);
and U3899 (N_3899,In_684,In_933);
nand U3900 (N_3900,In_1943,In_1986);
or U3901 (N_3901,In_47,In_478);
and U3902 (N_3902,In_1769,In_1721);
and U3903 (N_3903,In_2484,In_1429);
nor U3904 (N_3904,In_2069,In_1846);
nor U3905 (N_3905,In_2177,In_302);
or U3906 (N_3906,In_1627,In_869);
nor U3907 (N_3907,In_1683,In_1705);
nor U3908 (N_3908,In_88,In_205);
or U3909 (N_3909,In_1182,In_179);
nor U3910 (N_3910,In_1929,In_1426);
or U3911 (N_3911,In_840,In_308);
nand U3912 (N_3912,In_494,In_1754);
nor U3913 (N_3913,In_1763,In_1551);
nand U3914 (N_3914,In_1059,In_1452);
and U3915 (N_3915,In_554,In_1459);
xnor U3916 (N_3916,In_1009,In_116);
nand U3917 (N_3917,In_645,In_504);
nand U3918 (N_3918,In_464,In_281);
and U3919 (N_3919,In_867,In_1313);
nand U3920 (N_3920,In_2017,In_1985);
nand U3921 (N_3921,In_10,In_2171);
nor U3922 (N_3922,In_2112,In_1971);
or U3923 (N_3923,In_2440,In_683);
or U3924 (N_3924,In_1156,In_2311);
or U3925 (N_3925,In_1621,In_1874);
and U3926 (N_3926,In_1108,In_313);
or U3927 (N_3927,In_1895,In_2186);
or U3928 (N_3928,In_248,In_2327);
nor U3929 (N_3929,In_1949,In_814);
nand U3930 (N_3930,In_1653,In_1694);
xnor U3931 (N_3931,In_2028,In_2227);
nor U3932 (N_3932,In_2335,In_439);
nand U3933 (N_3933,In_378,In_2299);
nor U3934 (N_3934,In_1038,In_1288);
or U3935 (N_3935,In_2365,In_845);
nand U3936 (N_3936,In_2085,In_930);
nor U3937 (N_3937,In_2450,In_1523);
or U3938 (N_3938,In_831,In_1979);
nor U3939 (N_3939,In_156,In_1137);
or U3940 (N_3940,In_380,In_583);
nor U3941 (N_3941,In_179,In_817);
nand U3942 (N_3942,In_385,In_1675);
nand U3943 (N_3943,In_2011,In_1366);
and U3944 (N_3944,In_470,In_369);
nor U3945 (N_3945,In_1155,In_857);
and U3946 (N_3946,In_2176,In_2446);
and U3947 (N_3947,In_338,In_1475);
nand U3948 (N_3948,In_161,In_2076);
or U3949 (N_3949,In_1234,In_242);
nand U3950 (N_3950,In_342,In_2042);
nor U3951 (N_3951,In_2197,In_824);
xor U3952 (N_3952,In_168,In_2209);
nor U3953 (N_3953,In_1415,In_865);
nand U3954 (N_3954,In_317,In_1958);
nand U3955 (N_3955,In_1031,In_352);
nor U3956 (N_3956,In_1489,In_36);
nand U3957 (N_3957,In_1462,In_547);
or U3958 (N_3958,In_519,In_2428);
nor U3959 (N_3959,In_488,In_434);
or U3960 (N_3960,In_524,In_593);
and U3961 (N_3961,In_1981,In_1924);
nand U3962 (N_3962,In_1733,In_257);
nor U3963 (N_3963,In_1558,In_2027);
or U3964 (N_3964,In_1166,In_2214);
nand U3965 (N_3965,In_1348,In_819);
nor U3966 (N_3966,In_1592,In_2196);
or U3967 (N_3967,In_826,In_2166);
and U3968 (N_3968,In_37,In_160);
nor U3969 (N_3969,In_1897,In_435);
nand U3970 (N_3970,In_897,In_1628);
nor U3971 (N_3971,In_1265,In_1050);
nor U3972 (N_3972,In_1808,In_1354);
or U3973 (N_3973,In_1520,In_2479);
nand U3974 (N_3974,In_2008,In_2073);
nand U3975 (N_3975,In_348,In_1393);
nand U3976 (N_3976,In_275,In_1367);
nand U3977 (N_3977,In_878,In_2088);
or U3978 (N_3978,In_1782,In_2034);
nand U3979 (N_3979,In_239,In_2465);
nand U3980 (N_3980,In_898,In_1179);
xor U3981 (N_3981,In_1943,In_1690);
and U3982 (N_3982,In_2312,In_1370);
nor U3983 (N_3983,In_1368,In_2018);
nand U3984 (N_3984,In_2376,In_1349);
or U3985 (N_3985,In_350,In_2169);
or U3986 (N_3986,In_37,In_1673);
nor U3987 (N_3987,In_1237,In_1249);
nand U3988 (N_3988,In_620,In_638);
nand U3989 (N_3989,In_1044,In_2294);
nand U3990 (N_3990,In_2143,In_18);
nor U3991 (N_3991,In_68,In_1051);
nand U3992 (N_3992,In_31,In_1039);
or U3993 (N_3993,In_477,In_1985);
nor U3994 (N_3994,In_502,In_2377);
and U3995 (N_3995,In_1828,In_610);
xor U3996 (N_3996,In_2246,In_234);
or U3997 (N_3997,In_1715,In_1211);
and U3998 (N_3998,In_1034,In_1577);
or U3999 (N_3999,In_2246,In_14);
or U4000 (N_4000,In_1839,In_1092);
nor U4001 (N_4001,In_564,In_336);
nand U4002 (N_4002,In_160,In_1702);
and U4003 (N_4003,In_1136,In_1087);
xor U4004 (N_4004,In_75,In_1806);
or U4005 (N_4005,In_428,In_1425);
nor U4006 (N_4006,In_493,In_2323);
and U4007 (N_4007,In_2310,In_1079);
nand U4008 (N_4008,In_2037,In_886);
xor U4009 (N_4009,In_595,In_1114);
nor U4010 (N_4010,In_907,In_238);
or U4011 (N_4011,In_207,In_1885);
or U4012 (N_4012,In_2357,In_324);
and U4013 (N_4013,In_1388,In_39);
or U4014 (N_4014,In_1297,In_1636);
and U4015 (N_4015,In_202,In_199);
and U4016 (N_4016,In_1853,In_1171);
nor U4017 (N_4017,In_793,In_2156);
nand U4018 (N_4018,In_1452,In_1317);
or U4019 (N_4019,In_1945,In_950);
or U4020 (N_4020,In_1315,In_816);
nor U4021 (N_4021,In_193,In_1560);
nand U4022 (N_4022,In_446,In_482);
nor U4023 (N_4023,In_1182,In_88);
nand U4024 (N_4024,In_644,In_8);
nor U4025 (N_4025,In_2431,In_524);
nor U4026 (N_4026,In_1414,In_588);
and U4027 (N_4027,In_1959,In_508);
and U4028 (N_4028,In_793,In_261);
and U4029 (N_4029,In_2175,In_313);
nor U4030 (N_4030,In_467,In_670);
and U4031 (N_4031,In_1167,In_1984);
and U4032 (N_4032,In_573,In_627);
nor U4033 (N_4033,In_883,In_53);
or U4034 (N_4034,In_2274,In_2361);
or U4035 (N_4035,In_496,In_247);
or U4036 (N_4036,In_2287,In_48);
xnor U4037 (N_4037,In_1114,In_437);
nand U4038 (N_4038,In_1903,In_53);
nor U4039 (N_4039,In_1505,In_1327);
nor U4040 (N_4040,In_988,In_2499);
nor U4041 (N_4041,In_1594,In_434);
xor U4042 (N_4042,In_1934,In_1526);
nand U4043 (N_4043,In_1755,In_2422);
nor U4044 (N_4044,In_1650,In_720);
or U4045 (N_4045,In_6,In_531);
nor U4046 (N_4046,In_2467,In_2092);
nor U4047 (N_4047,In_2001,In_480);
and U4048 (N_4048,In_746,In_2057);
and U4049 (N_4049,In_345,In_411);
nor U4050 (N_4050,In_866,In_1449);
and U4051 (N_4051,In_2118,In_975);
and U4052 (N_4052,In_118,In_610);
and U4053 (N_4053,In_31,In_1681);
nor U4054 (N_4054,In_775,In_1984);
nand U4055 (N_4055,In_1348,In_2037);
or U4056 (N_4056,In_424,In_995);
xor U4057 (N_4057,In_1652,In_1586);
nor U4058 (N_4058,In_729,In_2441);
xnor U4059 (N_4059,In_561,In_2188);
nor U4060 (N_4060,In_2455,In_609);
or U4061 (N_4061,In_1916,In_430);
or U4062 (N_4062,In_948,In_1097);
xor U4063 (N_4063,In_2427,In_839);
nor U4064 (N_4064,In_1734,In_1380);
nand U4065 (N_4065,In_1309,In_2435);
and U4066 (N_4066,In_1085,In_319);
nor U4067 (N_4067,In_2389,In_2233);
nor U4068 (N_4068,In_1604,In_2207);
nand U4069 (N_4069,In_2032,In_791);
nand U4070 (N_4070,In_1330,In_1842);
nor U4071 (N_4071,In_1327,In_1301);
nor U4072 (N_4072,In_79,In_2088);
nand U4073 (N_4073,In_1703,In_1480);
nor U4074 (N_4074,In_883,In_684);
or U4075 (N_4075,In_47,In_1236);
or U4076 (N_4076,In_379,In_2190);
or U4077 (N_4077,In_1465,In_1658);
nor U4078 (N_4078,In_2090,In_122);
and U4079 (N_4079,In_943,In_1670);
nor U4080 (N_4080,In_665,In_379);
and U4081 (N_4081,In_1861,In_419);
nand U4082 (N_4082,In_1797,In_1272);
and U4083 (N_4083,In_1331,In_230);
nor U4084 (N_4084,In_797,In_1842);
xor U4085 (N_4085,In_1141,In_346);
nand U4086 (N_4086,In_2118,In_1242);
and U4087 (N_4087,In_289,In_1928);
nand U4088 (N_4088,In_707,In_24);
nand U4089 (N_4089,In_1731,In_1855);
nand U4090 (N_4090,In_726,In_552);
and U4091 (N_4091,In_92,In_1040);
nand U4092 (N_4092,In_1569,In_1638);
and U4093 (N_4093,In_136,In_1757);
nand U4094 (N_4094,In_1940,In_526);
nor U4095 (N_4095,In_1975,In_2372);
and U4096 (N_4096,In_312,In_2035);
or U4097 (N_4097,In_442,In_382);
xnor U4098 (N_4098,In_1917,In_1224);
nor U4099 (N_4099,In_853,In_2487);
and U4100 (N_4100,In_2381,In_2211);
and U4101 (N_4101,In_467,In_923);
and U4102 (N_4102,In_498,In_1302);
or U4103 (N_4103,In_1569,In_72);
nor U4104 (N_4104,In_2310,In_420);
and U4105 (N_4105,In_126,In_1251);
nand U4106 (N_4106,In_2078,In_1575);
nand U4107 (N_4107,In_862,In_1614);
or U4108 (N_4108,In_1953,In_2040);
nor U4109 (N_4109,In_884,In_1183);
or U4110 (N_4110,In_124,In_2428);
nor U4111 (N_4111,In_2234,In_2197);
nand U4112 (N_4112,In_1064,In_2264);
or U4113 (N_4113,In_2442,In_2454);
or U4114 (N_4114,In_1539,In_2457);
nor U4115 (N_4115,In_742,In_510);
nor U4116 (N_4116,In_1283,In_170);
nor U4117 (N_4117,In_1703,In_2116);
and U4118 (N_4118,In_598,In_1467);
and U4119 (N_4119,In_333,In_647);
nor U4120 (N_4120,In_951,In_1530);
nor U4121 (N_4121,In_93,In_8);
or U4122 (N_4122,In_961,In_2277);
nand U4123 (N_4123,In_32,In_328);
or U4124 (N_4124,In_1635,In_2176);
and U4125 (N_4125,In_1416,In_271);
and U4126 (N_4126,In_2150,In_1187);
nand U4127 (N_4127,In_391,In_490);
nor U4128 (N_4128,In_1461,In_1380);
and U4129 (N_4129,In_1567,In_712);
and U4130 (N_4130,In_2367,In_1836);
nand U4131 (N_4131,In_2310,In_436);
nor U4132 (N_4132,In_2030,In_1809);
nand U4133 (N_4133,In_1343,In_1555);
or U4134 (N_4134,In_1075,In_1427);
nor U4135 (N_4135,In_754,In_388);
xor U4136 (N_4136,In_1817,In_228);
nor U4137 (N_4137,In_1811,In_1637);
or U4138 (N_4138,In_726,In_1304);
nor U4139 (N_4139,In_377,In_418);
or U4140 (N_4140,In_2097,In_942);
nor U4141 (N_4141,In_555,In_849);
and U4142 (N_4142,In_8,In_1571);
or U4143 (N_4143,In_1642,In_1913);
and U4144 (N_4144,In_1942,In_1287);
and U4145 (N_4145,In_713,In_2391);
and U4146 (N_4146,In_1849,In_835);
and U4147 (N_4147,In_156,In_1571);
or U4148 (N_4148,In_2428,In_1412);
nor U4149 (N_4149,In_1895,In_347);
or U4150 (N_4150,In_1806,In_1659);
nor U4151 (N_4151,In_1096,In_2292);
xnor U4152 (N_4152,In_33,In_2108);
xnor U4153 (N_4153,In_1057,In_1575);
and U4154 (N_4154,In_1795,In_1239);
nor U4155 (N_4155,In_2411,In_2057);
or U4156 (N_4156,In_890,In_2140);
nand U4157 (N_4157,In_2017,In_1855);
nand U4158 (N_4158,In_612,In_153);
or U4159 (N_4159,In_1900,In_723);
xnor U4160 (N_4160,In_1471,In_1037);
and U4161 (N_4161,In_1160,In_1962);
or U4162 (N_4162,In_901,In_907);
nor U4163 (N_4163,In_2422,In_856);
and U4164 (N_4164,In_2346,In_1050);
or U4165 (N_4165,In_1695,In_1410);
nand U4166 (N_4166,In_1202,In_1906);
nand U4167 (N_4167,In_656,In_2239);
or U4168 (N_4168,In_1107,In_55);
nand U4169 (N_4169,In_1135,In_467);
nor U4170 (N_4170,In_1178,In_959);
nor U4171 (N_4171,In_1394,In_217);
or U4172 (N_4172,In_760,In_1784);
nand U4173 (N_4173,In_2285,In_1333);
xor U4174 (N_4174,In_1841,In_2106);
nand U4175 (N_4175,In_501,In_334);
nand U4176 (N_4176,In_39,In_1335);
and U4177 (N_4177,In_1812,In_28);
or U4178 (N_4178,In_726,In_929);
and U4179 (N_4179,In_2451,In_8);
and U4180 (N_4180,In_2453,In_1078);
and U4181 (N_4181,In_882,In_1061);
or U4182 (N_4182,In_1703,In_1064);
nand U4183 (N_4183,In_1482,In_452);
and U4184 (N_4184,In_2240,In_536);
nand U4185 (N_4185,In_1999,In_1142);
xnor U4186 (N_4186,In_418,In_937);
nor U4187 (N_4187,In_674,In_1063);
or U4188 (N_4188,In_1607,In_2097);
nand U4189 (N_4189,In_2049,In_1330);
nand U4190 (N_4190,In_146,In_345);
or U4191 (N_4191,In_334,In_2491);
or U4192 (N_4192,In_2012,In_888);
nand U4193 (N_4193,In_734,In_537);
or U4194 (N_4194,In_496,In_2066);
nor U4195 (N_4195,In_105,In_1192);
nor U4196 (N_4196,In_10,In_376);
and U4197 (N_4197,In_1171,In_1217);
nand U4198 (N_4198,In_1071,In_1920);
nor U4199 (N_4199,In_1638,In_700);
nand U4200 (N_4200,In_2279,In_1086);
or U4201 (N_4201,In_748,In_1754);
nand U4202 (N_4202,In_839,In_2198);
nand U4203 (N_4203,In_1356,In_388);
and U4204 (N_4204,In_88,In_735);
nor U4205 (N_4205,In_674,In_810);
and U4206 (N_4206,In_2347,In_507);
or U4207 (N_4207,In_1434,In_1596);
nor U4208 (N_4208,In_1235,In_227);
nand U4209 (N_4209,In_1945,In_1413);
xor U4210 (N_4210,In_1320,In_375);
nand U4211 (N_4211,In_1635,In_960);
and U4212 (N_4212,In_1079,In_973);
nand U4213 (N_4213,In_908,In_1393);
or U4214 (N_4214,In_166,In_899);
or U4215 (N_4215,In_480,In_908);
and U4216 (N_4216,In_2118,In_2232);
nand U4217 (N_4217,In_385,In_2406);
and U4218 (N_4218,In_731,In_1678);
or U4219 (N_4219,In_1438,In_330);
or U4220 (N_4220,In_795,In_1410);
nor U4221 (N_4221,In_2034,In_549);
nor U4222 (N_4222,In_1879,In_279);
and U4223 (N_4223,In_920,In_598);
and U4224 (N_4224,In_2346,In_726);
xnor U4225 (N_4225,In_191,In_1609);
nand U4226 (N_4226,In_1887,In_2270);
nand U4227 (N_4227,In_1213,In_293);
nor U4228 (N_4228,In_2382,In_2453);
and U4229 (N_4229,In_213,In_1174);
nor U4230 (N_4230,In_455,In_1595);
and U4231 (N_4231,In_906,In_1701);
and U4232 (N_4232,In_1033,In_1237);
nor U4233 (N_4233,In_626,In_1372);
nor U4234 (N_4234,In_2012,In_1184);
and U4235 (N_4235,In_2232,In_2108);
or U4236 (N_4236,In_1450,In_1159);
or U4237 (N_4237,In_791,In_546);
nor U4238 (N_4238,In_2097,In_961);
nor U4239 (N_4239,In_199,In_109);
nor U4240 (N_4240,In_295,In_1820);
nand U4241 (N_4241,In_2126,In_872);
nand U4242 (N_4242,In_859,In_1414);
nor U4243 (N_4243,In_2408,In_1197);
or U4244 (N_4244,In_178,In_679);
or U4245 (N_4245,In_679,In_1047);
and U4246 (N_4246,In_1410,In_1292);
or U4247 (N_4247,In_1851,In_1054);
or U4248 (N_4248,In_1381,In_24);
nor U4249 (N_4249,In_1091,In_627);
nand U4250 (N_4250,In_1940,In_2067);
or U4251 (N_4251,In_2398,In_1920);
nand U4252 (N_4252,In_1942,In_1494);
or U4253 (N_4253,In_1794,In_718);
nor U4254 (N_4254,In_233,In_2388);
or U4255 (N_4255,In_2179,In_1366);
and U4256 (N_4256,In_694,In_1116);
nor U4257 (N_4257,In_1414,In_1462);
and U4258 (N_4258,In_1650,In_217);
and U4259 (N_4259,In_1682,In_398);
and U4260 (N_4260,In_633,In_1057);
or U4261 (N_4261,In_2290,In_803);
and U4262 (N_4262,In_2365,In_1123);
and U4263 (N_4263,In_661,In_710);
nand U4264 (N_4264,In_1226,In_1528);
nand U4265 (N_4265,In_2132,In_1178);
nor U4266 (N_4266,In_1062,In_1860);
and U4267 (N_4267,In_1302,In_189);
nor U4268 (N_4268,In_531,In_267);
and U4269 (N_4269,In_1295,In_833);
or U4270 (N_4270,In_382,In_2312);
nand U4271 (N_4271,In_2209,In_1077);
or U4272 (N_4272,In_1625,In_263);
or U4273 (N_4273,In_1060,In_1056);
and U4274 (N_4274,In_1434,In_532);
nor U4275 (N_4275,In_732,In_1728);
or U4276 (N_4276,In_141,In_55);
or U4277 (N_4277,In_1133,In_1183);
nor U4278 (N_4278,In_1738,In_2113);
or U4279 (N_4279,In_260,In_645);
nand U4280 (N_4280,In_1827,In_2334);
xor U4281 (N_4281,In_2314,In_381);
or U4282 (N_4282,In_2456,In_341);
xnor U4283 (N_4283,In_838,In_1561);
and U4284 (N_4284,In_969,In_2435);
nand U4285 (N_4285,In_551,In_529);
and U4286 (N_4286,In_333,In_1023);
nor U4287 (N_4287,In_363,In_1150);
or U4288 (N_4288,In_106,In_1542);
xor U4289 (N_4289,In_1334,In_2186);
nor U4290 (N_4290,In_764,In_2122);
or U4291 (N_4291,In_1364,In_2432);
nor U4292 (N_4292,In_1902,In_2350);
nor U4293 (N_4293,In_589,In_1039);
nand U4294 (N_4294,In_964,In_1463);
nor U4295 (N_4295,In_1195,In_11);
and U4296 (N_4296,In_1331,In_1060);
and U4297 (N_4297,In_859,In_1711);
nand U4298 (N_4298,In_75,In_738);
nor U4299 (N_4299,In_309,In_2044);
or U4300 (N_4300,In_453,In_1614);
nand U4301 (N_4301,In_867,In_2057);
and U4302 (N_4302,In_1630,In_178);
nand U4303 (N_4303,In_1799,In_107);
and U4304 (N_4304,In_46,In_1821);
or U4305 (N_4305,In_1097,In_116);
and U4306 (N_4306,In_2403,In_1587);
nor U4307 (N_4307,In_143,In_761);
nor U4308 (N_4308,In_503,In_246);
and U4309 (N_4309,In_975,In_766);
nor U4310 (N_4310,In_1607,In_295);
and U4311 (N_4311,In_997,In_966);
nand U4312 (N_4312,In_753,In_656);
or U4313 (N_4313,In_880,In_1674);
nor U4314 (N_4314,In_1410,In_1442);
or U4315 (N_4315,In_1338,In_404);
and U4316 (N_4316,In_1234,In_694);
and U4317 (N_4317,In_111,In_2156);
nand U4318 (N_4318,In_1431,In_812);
nand U4319 (N_4319,In_2289,In_594);
nor U4320 (N_4320,In_1537,In_233);
and U4321 (N_4321,In_150,In_2056);
or U4322 (N_4322,In_2226,In_1651);
and U4323 (N_4323,In_474,In_2306);
nor U4324 (N_4324,In_1211,In_1424);
and U4325 (N_4325,In_2442,In_1409);
nand U4326 (N_4326,In_1597,In_2257);
or U4327 (N_4327,In_2220,In_2008);
nand U4328 (N_4328,In_982,In_1675);
or U4329 (N_4329,In_1206,In_1009);
and U4330 (N_4330,In_826,In_1580);
and U4331 (N_4331,In_391,In_2154);
nor U4332 (N_4332,In_2245,In_1708);
nor U4333 (N_4333,In_905,In_498);
or U4334 (N_4334,In_1733,In_940);
nor U4335 (N_4335,In_1521,In_1016);
nand U4336 (N_4336,In_1556,In_1044);
or U4337 (N_4337,In_1188,In_1663);
nand U4338 (N_4338,In_1389,In_1674);
xor U4339 (N_4339,In_854,In_1707);
nor U4340 (N_4340,In_1573,In_679);
and U4341 (N_4341,In_829,In_1427);
nand U4342 (N_4342,In_2319,In_1548);
xnor U4343 (N_4343,In_961,In_867);
nor U4344 (N_4344,In_689,In_1270);
nor U4345 (N_4345,In_2436,In_1182);
nand U4346 (N_4346,In_84,In_429);
nand U4347 (N_4347,In_1097,In_1204);
or U4348 (N_4348,In_1993,In_1977);
nor U4349 (N_4349,In_2319,In_1609);
or U4350 (N_4350,In_1606,In_1972);
and U4351 (N_4351,In_1224,In_490);
and U4352 (N_4352,In_1390,In_1974);
and U4353 (N_4353,In_1964,In_1843);
nor U4354 (N_4354,In_165,In_241);
nand U4355 (N_4355,In_1347,In_981);
and U4356 (N_4356,In_1600,In_802);
nor U4357 (N_4357,In_1247,In_1423);
nand U4358 (N_4358,In_434,In_773);
nor U4359 (N_4359,In_2048,In_2286);
nor U4360 (N_4360,In_1035,In_1165);
nand U4361 (N_4361,In_484,In_439);
and U4362 (N_4362,In_1356,In_1726);
nor U4363 (N_4363,In_1564,In_1401);
or U4364 (N_4364,In_923,In_1094);
or U4365 (N_4365,In_2431,In_1826);
or U4366 (N_4366,In_1463,In_1873);
and U4367 (N_4367,In_2360,In_1031);
nor U4368 (N_4368,In_2210,In_2236);
nand U4369 (N_4369,In_80,In_1568);
xor U4370 (N_4370,In_556,In_598);
or U4371 (N_4371,In_1246,In_1022);
and U4372 (N_4372,In_829,In_2091);
or U4373 (N_4373,In_1225,In_2051);
nand U4374 (N_4374,In_1688,In_48);
nor U4375 (N_4375,In_1873,In_703);
nor U4376 (N_4376,In_1327,In_1250);
and U4377 (N_4377,In_1642,In_337);
and U4378 (N_4378,In_1787,In_866);
nor U4379 (N_4379,In_1217,In_2306);
nor U4380 (N_4380,In_1457,In_1073);
or U4381 (N_4381,In_2205,In_1462);
and U4382 (N_4382,In_66,In_2440);
nor U4383 (N_4383,In_1443,In_2488);
nand U4384 (N_4384,In_2450,In_85);
nand U4385 (N_4385,In_2226,In_1519);
or U4386 (N_4386,In_2328,In_242);
or U4387 (N_4387,In_312,In_922);
nor U4388 (N_4388,In_713,In_817);
or U4389 (N_4389,In_2128,In_39);
or U4390 (N_4390,In_1495,In_607);
or U4391 (N_4391,In_78,In_1701);
and U4392 (N_4392,In_1845,In_2223);
nand U4393 (N_4393,In_483,In_2133);
or U4394 (N_4394,In_1723,In_184);
nor U4395 (N_4395,In_1263,In_1082);
nor U4396 (N_4396,In_687,In_699);
nor U4397 (N_4397,In_896,In_1411);
or U4398 (N_4398,In_868,In_2451);
and U4399 (N_4399,In_564,In_2463);
or U4400 (N_4400,In_864,In_568);
nand U4401 (N_4401,In_626,In_2316);
xnor U4402 (N_4402,In_991,In_148);
and U4403 (N_4403,In_1299,In_519);
nand U4404 (N_4404,In_2051,In_911);
and U4405 (N_4405,In_2199,In_2179);
xor U4406 (N_4406,In_1647,In_365);
nand U4407 (N_4407,In_1616,In_83);
or U4408 (N_4408,In_1229,In_777);
nand U4409 (N_4409,In_1780,In_1684);
nor U4410 (N_4410,In_1798,In_781);
or U4411 (N_4411,In_1266,In_1268);
nor U4412 (N_4412,In_2452,In_2131);
or U4413 (N_4413,In_2183,In_2332);
or U4414 (N_4414,In_1302,In_2216);
or U4415 (N_4415,In_1576,In_258);
and U4416 (N_4416,In_222,In_2120);
nor U4417 (N_4417,In_800,In_971);
or U4418 (N_4418,In_963,In_2005);
nor U4419 (N_4419,In_741,In_1361);
or U4420 (N_4420,In_1817,In_1190);
and U4421 (N_4421,In_999,In_1678);
nand U4422 (N_4422,In_2078,In_995);
nand U4423 (N_4423,In_1466,In_1926);
nand U4424 (N_4424,In_892,In_678);
or U4425 (N_4425,In_1415,In_981);
nor U4426 (N_4426,In_876,In_1206);
or U4427 (N_4427,In_1163,In_1703);
nand U4428 (N_4428,In_2244,In_967);
nor U4429 (N_4429,In_1783,In_737);
nor U4430 (N_4430,In_529,In_1058);
xnor U4431 (N_4431,In_1529,In_1916);
and U4432 (N_4432,In_1064,In_385);
and U4433 (N_4433,In_71,In_371);
or U4434 (N_4434,In_1357,In_558);
and U4435 (N_4435,In_2442,In_1366);
or U4436 (N_4436,In_11,In_70);
and U4437 (N_4437,In_2049,In_390);
xor U4438 (N_4438,In_2041,In_806);
and U4439 (N_4439,In_41,In_1089);
nor U4440 (N_4440,In_1550,In_2333);
or U4441 (N_4441,In_905,In_476);
or U4442 (N_4442,In_669,In_1131);
nor U4443 (N_4443,In_1357,In_663);
xor U4444 (N_4444,In_560,In_1466);
nor U4445 (N_4445,In_2239,In_868);
and U4446 (N_4446,In_1603,In_2100);
or U4447 (N_4447,In_2053,In_2046);
nand U4448 (N_4448,In_2356,In_624);
nand U4449 (N_4449,In_2066,In_1933);
nand U4450 (N_4450,In_2306,In_1926);
or U4451 (N_4451,In_479,In_804);
and U4452 (N_4452,In_1442,In_475);
xor U4453 (N_4453,In_1199,In_530);
and U4454 (N_4454,In_2426,In_862);
nand U4455 (N_4455,In_979,In_811);
nand U4456 (N_4456,In_50,In_2238);
nand U4457 (N_4457,In_1122,In_2171);
or U4458 (N_4458,In_1167,In_2021);
or U4459 (N_4459,In_139,In_1157);
or U4460 (N_4460,In_1613,In_1495);
nor U4461 (N_4461,In_2187,In_1383);
nor U4462 (N_4462,In_562,In_500);
nand U4463 (N_4463,In_232,In_1272);
nor U4464 (N_4464,In_1858,In_1177);
or U4465 (N_4465,In_1930,In_1706);
nor U4466 (N_4466,In_1661,In_1033);
and U4467 (N_4467,In_857,In_1364);
nor U4468 (N_4468,In_1633,In_605);
nand U4469 (N_4469,In_1385,In_1879);
nand U4470 (N_4470,In_2454,In_2407);
and U4471 (N_4471,In_1457,In_1270);
nand U4472 (N_4472,In_236,In_592);
or U4473 (N_4473,In_1480,In_2103);
nor U4474 (N_4474,In_1580,In_306);
nor U4475 (N_4475,In_1621,In_1488);
or U4476 (N_4476,In_1604,In_2362);
nor U4477 (N_4477,In_1777,In_1200);
or U4478 (N_4478,In_1780,In_1392);
or U4479 (N_4479,In_679,In_1975);
nand U4480 (N_4480,In_697,In_2466);
nor U4481 (N_4481,In_1658,In_322);
nand U4482 (N_4482,In_1434,In_2332);
or U4483 (N_4483,In_686,In_242);
nor U4484 (N_4484,In_731,In_199);
nand U4485 (N_4485,In_14,In_2036);
or U4486 (N_4486,In_1588,In_903);
nand U4487 (N_4487,In_1891,In_763);
nor U4488 (N_4488,In_984,In_535);
or U4489 (N_4489,In_1658,In_1887);
or U4490 (N_4490,In_2459,In_2278);
and U4491 (N_4491,In_1009,In_635);
nor U4492 (N_4492,In_2246,In_995);
and U4493 (N_4493,In_1953,In_1961);
and U4494 (N_4494,In_663,In_1191);
nor U4495 (N_4495,In_1003,In_2279);
or U4496 (N_4496,In_154,In_1172);
and U4497 (N_4497,In_1872,In_471);
and U4498 (N_4498,In_208,In_390);
nand U4499 (N_4499,In_1679,In_2443);
or U4500 (N_4500,In_1283,In_1726);
nand U4501 (N_4501,In_1251,In_1918);
xnor U4502 (N_4502,In_601,In_828);
nand U4503 (N_4503,In_958,In_1652);
nand U4504 (N_4504,In_19,In_74);
and U4505 (N_4505,In_322,In_356);
or U4506 (N_4506,In_966,In_1236);
and U4507 (N_4507,In_549,In_1699);
or U4508 (N_4508,In_2325,In_167);
and U4509 (N_4509,In_1302,In_509);
or U4510 (N_4510,In_829,In_1055);
nor U4511 (N_4511,In_521,In_120);
nor U4512 (N_4512,In_341,In_60);
or U4513 (N_4513,In_2406,In_372);
nand U4514 (N_4514,In_2385,In_1119);
and U4515 (N_4515,In_13,In_271);
and U4516 (N_4516,In_1613,In_1564);
nand U4517 (N_4517,In_1519,In_256);
nor U4518 (N_4518,In_621,In_1390);
xnor U4519 (N_4519,In_1589,In_652);
nor U4520 (N_4520,In_1115,In_1080);
nand U4521 (N_4521,In_698,In_2364);
nor U4522 (N_4522,In_72,In_2348);
or U4523 (N_4523,In_236,In_1725);
nand U4524 (N_4524,In_911,In_524);
or U4525 (N_4525,In_402,In_2392);
nor U4526 (N_4526,In_1657,In_2373);
and U4527 (N_4527,In_68,In_2139);
or U4528 (N_4528,In_81,In_1379);
and U4529 (N_4529,In_206,In_2233);
xnor U4530 (N_4530,In_55,In_1374);
nand U4531 (N_4531,In_2206,In_1293);
nand U4532 (N_4532,In_2262,In_2382);
nand U4533 (N_4533,In_416,In_1575);
or U4534 (N_4534,In_2190,In_818);
or U4535 (N_4535,In_2360,In_1965);
or U4536 (N_4536,In_1992,In_150);
and U4537 (N_4537,In_1409,In_2487);
nor U4538 (N_4538,In_545,In_706);
or U4539 (N_4539,In_1697,In_2088);
nand U4540 (N_4540,In_1187,In_682);
nor U4541 (N_4541,In_1727,In_2276);
and U4542 (N_4542,In_1199,In_799);
nand U4543 (N_4543,In_1560,In_1190);
or U4544 (N_4544,In_435,In_6);
and U4545 (N_4545,In_767,In_2040);
or U4546 (N_4546,In_1086,In_1047);
nand U4547 (N_4547,In_1128,In_1837);
nor U4548 (N_4548,In_2412,In_792);
nor U4549 (N_4549,In_1460,In_2108);
nand U4550 (N_4550,In_1425,In_1956);
nand U4551 (N_4551,In_1373,In_958);
nor U4552 (N_4552,In_2240,In_621);
nor U4553 (N_4553,In_196,In_189);
and U4554 (N_4554,In_758,In_1215);
nand U4555 (N_4555,In_2138,In_266);
and U4556 (N_4556,In_1718,In_1928);
nor U4557 (N_4557,In_494,In_480);
or U4558 (N_4558,In_250,In_1688);
and U4559 (N_4559,In_2041,In_2297);
and U4560 (N_4560,In_738,In_316);
nand U4561 (N_4561,In_1334,In_922);
nor U4562 (N_4562,In_2064,In_420);
nor U4563 (N_4563,In_2029,In_1677);
and U4564 (N_4564,In_256,In_1940);
nor U4565 (N_4565,In_1472,In_1249);
nor U4566 (N_4566,In_116,In_218);
or U4567 (N_4567,In_1023,In_1564);
or U4568 (N_4568,In_2099,In_1332);
nand U4569 (N_4569,In_452,In_427);
or U4570 (N_4570,In_296,In_187);
or U4571 (N_4571,In_1263,In_151);
nand U4572 (N_4572,In_147,In_1869);
nor U4573 (N_4573,In_1985,In_1639);
or U4574 (N_4574,In_2480,In_2224);
or U4575 (N_4575,In_607,In_1278);
xor U4576 (N_4576,In_726,In_2095);
nor U4577 (N_4577,In_544,In_1692);
nand U4578 (N_4578,In_1499,In_434);
and U4579 (N_4579,In_1068,In_1111);
xor U4580 (N_4580,In_859,In_326);
or U4581 (N_4581,In_2483,In_667);
xor U4582 (N_4582,In_2466,In_731);
nand U4583 (N_4583,In_1225,In_394);
nor U4584 (N_4584,In_870,In_2056);
and U4585 (N_4585,In_410,In_1023);
nand U4586 (N_4586,In_1502,In_2107);
nor U4587 (N_4587,In_965,In_2343);
nand U4588 (N_4588,In_2073,In_1223);
or U4589 (N_4589,In_560,In_2262);
nor U4590 (N_4590,In_381,In_1197);
nor U4591 (N_4591,In_1333,In_676);
nand U4592 (N_4592,In_369,In_1523);
or U4593 (N_4593,In_337,In_2044);
nand U4594 (N_4594,In_2252,In_2063);
nand U4595 (N_4595,In_1311,In_1128);
nand U4596 (N_4596,In_271,In_2212);
nand U4597 (N_4597,In_123,In_2124);
and U4598 (N_4598,In_1995,In_460);
nand U4599 (N_4599,In_2246,In_1412);
or U4600 (N_4600,In_1865,In_431);
or U4601 (N_4601,In_482,In_994);
and U4602 (N_4602,In_2127,In_959);
nand U4603 (N_4603,In_1166,In_276);
and U4604 (N_4604,In_91,In_1700);
nor U4605 (N_4605,In_135,In_157);
nand U4606 (N_4606,In_2403,In_2092);
or U4607 (N_4607,In_214,In_945);
and U4608 (N_4608,In_1482,In_1942);
or U4609 (N_4609,In_1897,In_608);
and U4610 (N_4610,In_325,In_293);
xor U4611 (N_4611,In_509,In_894);
and U4612 (N_4612,In_1342,In_688);
nor U4613 (N_4613,In_1637,In_282);
nor U4614 (N_4614,In_421,In_2481);
and U4615 (N_4615,In_819,In_686);
nand U4616 (N_4616,In_377,In_1054);
and U4617 (N_4617,In_1287,In_1283);
or U4618 (N_4618,In_739,In_1359);
nand U4619 (N_4619,In_1985,In_245);
and U4620 (N_4620,In_822,In_1785);
nand U4621 (N_4621,In_152,In_1037);
nand U4622 (N_4622,In_1153,In_848);
nand U4623 (N_4623,In_1146,In_413);
nand U4624 (N_4624,In_1695,In_1706);
nand U4625 (N_4625,In_174,In_1059);
nor U4626 (N_4626,In_628,In_1213);
or U4627 (N_4627,In_2288,In_2083);
nand U4628 (N_4628,In_647,In_1878);
nand U4629 (N_4629,In_1429,In_81);
nor U4630 (N_4630,In_1281,In_394);
or U4631 (N_4631,In_684,In_1049);
and U4632 (N_4632,In_2384,In_121);
and U4633 (N_4633,In_1479,In_899);
and U4634 (N_4634,In_924,In_356);
nand U4635 (N_4635,In_1784,In_2136);
nor U4636 (N_4636,In_59,In_2250);
nor U4637 (N_4637,In_210,In_1330);
nand U4638 (N_4638,In_2012,In_2465);
and U4639 (N_4639,In_2268,In_928);
nand U4640 (N_4640,In_1566,In_1213);
nor U4641 (N_4641,In_1721,In_1350);
and U4642 (N_4642,In_1239,In_332);
nand U4643 (N_4643,In_197,In_1665);
nor U4644 (N_4644,In_2477,In_84);
and U4645 (N_4645,In_2404,In_468);
nor U4646 (N_4646,In_2077,In_2156);
nor U4647 (N_4647,In_1613,In_1208);
nand U4648 (N_4648,In_1780,In_73);
nand U4649 (N_4649,In_809,In_511);
nand U4650 (N_4650,In_1190,In_2375);
nand U4651 (N_4651,In_990,In_2025);
or U4652 (N_4652,In_2378,In_2089);
nor U4653 (N_4653,In_2451,In_2300);
or U4654 (N_4654,In_174,In_1867);
nand U4655 (N_4655,In_1935,In_2102);
nand U4656 (N_4656,In_2293,In_1067);
and U4657 (N_4657,In_1566,In_571);
nand U4658 (N_4658,In_2482,In_2122);
nand U4659 (N_4659,In_786,In_2166);
nand U4660 (N_4660,In_2018,In_1478);
nand U4661 (N_4661,In_529,In_1850);
nor U4662 (N_4662,In_1821,In_808);
xor U4663 (N_4663,In_400,In_1528);
nand U4664 (N_4664,In_306,In_1255);
nand U4665 (N_4665,In_1452,In_1054);
and U4666 (N_4666,In_370,In_2061);
or U4667 (N_4667,In_1289,In_772);
nor U4668 (N_4668,In_1806,In_1669);
nor U4669 (N_4669,In_1256,In_1490);
nand U4670 (N_4670,In_1151,In_1605);
or U4671 (N_4671,In_1604,In_2031);
nor U4672 (N_4672,In_1765,In_44);
nor U4673 (N_4673,In_1260,In_942);
and U4674 (N_4674,In_2253,In_2121);
nor U4675 (N_4675,In_343,In_2207);
nand U4676 (N_4676,In_1554,In_1932);
and U4677 (N_4677,In_2237,In_2180);
nand U4678 (N_4678,In_2109,In_1733);
and U4679 (N_4679,In_1628,In_1076);
nand U4680 (N_4680,In_83,In_231);
nand U4681 (N_4681,In_2270,In_2143);
nand U4682 (N_4682,In_266,In_2496);
and U4683 (N_4683,In_437,In_982);
nand U4684 (N_4684,In_1629,In_223);
nor U4685 (N_4685,In_228,In_1064);
nand U4686 (N_4686,In_1608,In_1316);
or U4687 (N_4687,In_1739,In_1919);
nor U4688 (N_4688,In_2267,In_368);
nand U4689 (N_4689,In_736,In_574);
nor U4690 (N_4690,In_1653,In_1645);
nand U4691 (N_4691,In_2176,In_1361);
nand U4692 (N_4692,In_2035,In_1827);
or U4693 (N_4693,In_278,In_587);
and U4694 (N_4694,In_811,In_59);
or U4695 (N_4695,In_320,In_517);
nand U4696 (N_4696,In_1952,In_288);
nor U4697 (N_4697,In_1371,In_8);
and U4698 (N_4698,In_2094,In_1734);
nor U4699 (N_4699,In_1839,In_1405);
nand U4700 (N_4700,In_1884,In_484);
and U4701 (N_4701,In_768,In_1146);
nor U4702 (N_4702,In_1065,In_1803);
and U4703 (N_4703,In_1056,In_470);
or U4704 (N_4704,In_1083,In_2358);
and U4705 (N_4705,In_2485,In_2484);
nand U4706 (N_4706,In_2368,In_30);
or U4707 (N_4707,In_2131,In_1218);
and U4708 (N_4708,In_653,In_767);
and U4709 (N_4709,In_2131,In_1183);
nand U4710 (N_4710,In_1182,In_1449);
nor U4711 (N_4711,In_1294,In_2415);
or U4712 (N_4712,In_398,In_726);
nor U4713 (N_4713,In_1091,In_408);
or U4714 (N_4714,In_561,In_893);
and U4715 (N_4715,In_2145,In_875);
or U4716 (N_4716,In_1670,In_1246);
and U4717 (N_4717,In_1216,In_2212);
and U4718 (N_4718,In_28,In_426);
and U4719 (N_4719,In_1604,In_729);
nor U4720 (N_4720,In_442,In_1359);
nor U4721 (N_4721,In_178,In_87);
and U4722 (N_4722,In_582,In_179);
or U4723 (N_4723,In_2042,In_2450);
and U4724 (N_4724,In_1152,In_2396);
or U4725 (N_4725,In_127,In_2339);
or U4726 (N_4726,In_1590,In_830);
nand U4727 (N_4727,In_567,In_2081);
nor U4728 (N_4728,In_630,In_1618);
or U4729 (N_4729,In_1707,In_713);
and U4730 (N_4730,In_2258,In_1989);
or U4731 (N_4731,In_1613,In_215);
or U4732 (N_4732,In_1109,In_1034);
or U4733 (N_4733,In_1194,In_2318);
or U4734 (N_4734,In_1171,In_821);
xnor U4735 (N_4735,In_2146,In_580);
nor U4736 (N_4736,In_1050,In_1944);
and U4737 (N_4737,In_81,In_1705);
nand U4738 (N_4738,In_945,In_263);
or U4739 (N_4739,In_713,In_1631);
nor U4740 (N_4740,In_677,In_2366);
and U4741 (N_4741,In_1673,In_1706);
nand U4742 (N_4742,In_978,In_81);
nor U4743 (N_4743,In_2142,In_66);
nand U4744 (N_4744,In_1460,In_1461);
nor U4745 (N_4745,In_1099,In_1001);
or U4746 (N_4746,In_781,In_1175);
and U4747 (N_4747,In_1887,In_638);
and U4748 (N_4748,In_457,In_778);
nor U4749 (N_4749,In_2263,In_1621);
nor U4750 (N_4750,In_1316,In_985);
and U4751 (N_4751,In_2462,In_2188);
and U4752 (N_4752,In_2244,In_568);
nor U4753 (N_4753,In_1591,In_114);
or U4754 (N_4754,In_1744,In_511);
nand U4755 (N_4755,In_197,In_1625);
nor U4756 (N_4756,In_2146,In_1993);
xor U4757 (N_4757,In_2223,In_1135);
or U4758 (N_4758,In_1098,In_1471);
or U4759 (N_4759,In_325,In_833);
nor U4760 (N_4760,In_2336,In_2156);
nand U4761 (N_4761,In_512,In_770);
nand U4762 (N_4762,In_1419,In_489);
and U4763 (N_4763,In_2209,In_67);
or U4764 (N_4764,In_1511,In_1733);
and U4765 (N_4765,In_1162,In_2396);
nor U4766 (N_4766,In_240,In_1631);
nor U4767 (N_4767,In_1825,In_524);
and U4768 (N_4768,In_2067,In_1150);
and U4769 (N_4769,In_611,In_1554);
or U4770 (N_4770,In_2250,In_2060);
or U4771 (N_4771,In_1880,In_1513);
and U4772 (N_4772,In_1996,In_1297);
nor U4773 (N_4773,In_1778,In_1508);
or U4774 (N_4774,In_1847,In_370);
nor U4775 (N_4775,In_1001,In_1803);
or U4776 (N_4776,In_809,In_325);
nand U4777 (N_4777,In_1617,In_945);
nand U4778 (N_4778,In_1395,In_424);
nand U4779 (N_4779,In_2445,In_327);
and U4780 (N_4780,In_2254,In_821);
nor U4781 (N_4781,In_2123,In_460);
or U4782 (N_4782,In_1597,In_2263);
nand U4783 (N_4783,In_2272,In_154);
and U4784 (N_4784,In_2181,In_2025);
nor U4785 (N_4785,In_1378,In_472);
nor U4786 (N_4786,In_1195,In_218);
or U4787 (N_4787,In_246,In_187);
nor U4788 (N_4788,In_998,In_1258);
and U4789 (N_4789,In_2087,In_263);
nor U4790 (N_4790,In_1199,In_405);
or U4791 (N_4791,In_1741,In_1495);
xnor U4792 (N_4792,In_2353,In_2314);
nand U4793 (N_4793,In_940,In_1479);
or U4794 (N_4794,In_701,In_1801);
nor U4795 (N_4795,In_99,In_848);
or U4796 (N_4796,In_1901,In_592);
nand U4797 (N_4797,In_1606,In_242);
nor U4798 (N_4798,In_1034,In_1503);
nand U4799 (N_4799,In_2161,In_1646);
and U4800 (N_4800,In_1851,In_2186);
nand U4801 (N_4801,In_1239,In_881);
and U4802 (N_4802,In_559,In_408);
or U4803 (N_4803,In_695,In_2116);
or U4804 (N_4804,In_807,In_2288);
nand U4805 (N_4805,In_399,In_155);
nor U4806 (N_4806,In_1629,In_2160);
or U4807 (N_4807,In_562,In_723);
nand U4808 (N_4808,In_2142,In_628);
nor U4809 (N_4809,In_743,In_1567);
or U4810 (N_4810,In_1263,In_230);
or U4811 (N_4811,In_2424,In_1001);
nor U4812 (N_4812,In_2280,In_228);
or U4813 (N_4813,In_1040,In_1808);
nor U4814 (N_4814,In_1877,In_725);
nor U4815 (N_4815,In_1812,In_1027);
or U4816 (N_4816,In_157,In_2353);
nand U4817 (N_4817,In_1811,In_325);
and U4818 (N_4818,In_1690,In_227);
nand U4819 (N_4819,In_1801,In_1097);
nand U4820 (N_4820,In_1469,In_2494);
or U4821 (N_4821,In_1387,In_1136);
nor U4822 (N_4822,In_1908,In_1778);
and U4823 (N_4823,In_1344,In_2210);
nand U4824 (N_4824,In_1377,In_1902);
or U4825 (N_4825,In_557,In_311);
and U4826 (N_4826,In_798,In_1476);
and U4827 (N_4827,In_1188,In_747);
nor U4828 (N_4828,In_1549,In_2232);
nor U4829 (N_4829,In_60,In_2271);
nor U4830 (N_4830,In_2233,In_714);
or U4831 (N_4831,In_1450,In_288);
or U4832 (N_4832,In_2320,In_1661);
and U4833 (N_4833,In_372,In_2136);
nand U4834 (N_4834,In_759,In_185);
or U4835 (N_4835,In_1407,In_1683);
or U4836 (N_4836,In_859,In_28);
nor U4837 (N_4837,In_1882,In_733);
and U4838 (N_4838,In_788,In_1747);
nor U4839 (N_4839,In_1817,In_109);
nor U4840 (N_4840,In_944,In_46);
nand U4841 (N_4841,In_1257,In_2294);
or U4842 (N_4842,In_1996,In_823);
or U4843 (N_4843,In_1055,In_1015);
or U4844 (N_4844,In_1779,In_1628);
nand U4845 (N_4845,In_1460,In_881);
and U4846 (N_4846,In_1313,In_941);
nand U4847 (N_4847,In_1270,In_759);
nor U4848 (N_4848,In_1553,In_1023);
or U4849 (N_4849,In_2074,In_381);
and U4850 (N_4850,In_1562,In_1050);
nor U4851 (N_4851,In_510,In_1771);
nor U4852 (N_4852,In_1380,In_1116);
or U4853 (N_4853,In_2481,In_1125);
and U4854 (N_4854,In_512,In_958);
and U4855 (N_4855,In_386,In_1555);
nand U4856 (N_4856,In_120,In_1551);
or U4857 (N_4857,In_1446,In_2289);
nand U4858 (N_4858,In_1965,In_674);
nor U4859 (N_4859,In_1992,In_1947);
or U4860 (N_4860,In_117,In_2328);
nor U4861 (N_4861,In_1270,In_1700);
or U4862 (N_4862,In_2163,In_203);
and U4863 (N_4863,In_1057,In_1787);
nor U4864 (N_4864,In_1398,In_998);
and U4865 (N_4865,In_2199,In_1342);
or U4866 (N_4866,In_2355,In_2021);
or U4867 (N_4867,In_2150,In_632);
or U4868 (N_4868,In_126,In_1852);
or U4869 (N_4869,In_1721,In_1992);
and U4870 (N_4870,In_513,In_2470);
and U4871 (N_4871,In_1864,In_1624);
nand U4872 (N_4872,In_1470,In_1010);
nor U4873 (N_4873,In_846,In_211);
xnor U4874 (N_4874,In_158,In_1691);
nor U4875 (N_4875,In_1062,In_1584);
xor U4876 (N_4876,In_535,In_1927);
nand U4877 (N_4877,In_584,In_2006);
nand U4878 (N_4878,In_2244,In_155);
nor U4879 (N_4879,In_1784,In_1851);
and U4880 (N_4880,In_2155,In_1369);
xor U4881 (N_4881,In_200,In_1553);
nand U4882 (N_4882,In_388,In_319);
or U4883 (N_4883,In_1224,In_835);
and U4884 (N_4884,In_1051,In_1730);
or U4885 (N_4885,In_2233,In_2490);
nand U4886 (N_4886,In_1543,In_1350);
nor U4887 (N_4887,In_2136,In_2204);
or U4888 (N_4888,In_335,In_915);
nand U4889 (N_4889,In_1292,In_1883);
and U4890 (N_4890,In_517,In_54);
nor U4891 (N_4891,In_531,In_1528);
nand U4892 (N_4892,In_1301,In_427);
nand U4893 (N_4893,In_2331,In_1645);
nand U4894 (N_4894,In_1975,In_477);
and U4895 (N_4895,In_2263,In_1835);
and U4896 (N_4896,In_2396,In_42);
and U4897 (N_4897,In_2330,In_2229);
or U4898 (N_4898,In_1827,In_937);
and U4899 (N_4899,In_727,In_770);
or U4900 (N_4900,In_1634,In_2466);
or U4901 (N_4901,In_881,In_1402);
nor U4902 (N_4902,In_995,In_1710);
nor U4903 (N_4903,In_731,In_2399);
nor U4904 (N_4904,In_828,In_1493);
nand U4905 (N_4905,In_1637,In_1201);
nand U4906 (N_4906,In_1440,In_429);
and U4907 (N_4907,In_2008,In_2397);
or U4908 (N_4908,In_524,In_1706);
or U4909 (N_4909,In_1505,In_795);
nand U4910 (N_4910,In_996,In_197);
or U4911 (N_4911,In_294,In_1401);
or U4912 (N_4912,In_40,In_92);
nand U4913 (N_4913,In_2009,In_2127);
or U4914 (N_4914,In_708,In_1597);
or U4915 (N_4915,In_2131,In_258);
nand U4916 (N_4916,In_1477,In_1392);
nand U4917 (N_4917,In_852,In_874);
or U4918 (N_4918,In_1575,In_1946);
xor U4919 (N_4919,In_1819,In_1575);
nand U4920 (N_4920,In_8,In_643);
or U4921 (N_4921,In_1094,In_1704);
nand U4922 (N_4922,In_1711,In_1304);
or U4923 (N_4923,In_1340,In_29);
and U4924 (N_4924,In_1748,In_2139);
and U4925 (N_4925,In_1618,In_396);
nand U4926 (N_4926,In_443,In_2024);
or U4927 (N_4927,In_1896,In_1733);
or U4928 (N_4928,In_1966,In_189);
nor U4929 (N_4929,In_2048,In_1769);
nand U4930 (N_4930,In_804,In_2413);
nor U4931 (N_4931,In_408,In_1596);
and U4932 (N_4932,In_90,In_24);
and U4933 (N_4933,In_812,In_244);
nand U4934 (N_4934,In_1331,In_2037);
and U4935 (N_4935,In_1986,In_567);
nor U4936 (N_4936,In_782,In_1131);
or U4937 (N_4937,In_2338,In_972);
or U4938 (N_4938,In_684,In_2091);
nand U4939 (N_4939,In_1015,In_619);
or U4940 (N_4940,In_1686,In_2410);
nand U4941 (N_4941,In_2174,In_2041);
nor U4942 (N_4942,In_1862,In_923);
and U4943 (N_4943,In_261,In_1956);
nor U4944 (N_4944,In_947,In_1157);
nand U4945 (N_4945,In_979,In_848);
nor U4946 (N_4946,In_651,In_2449);
or U4947 (N_4947,In_1076,In_1895);
and U4948 (N_4948,In_699,In_946);
or U4949 (N_4949,In_677,In_1822);
nand U4950 (N_4950,In_1339,In_1567);
nor U4951 (N_4951,In_706,In_2331);
or U4952 (N_4952,In_663,In_2068);
nand U4953 (N_4953,In_734,In_1099);
xor U4954 (N_4954,In_2134,In_2337);
nand U4955 (N_4955,In_951,In_804);
and U4956 (N_4956,In_2294,In_1938);
nor U4957 (N_4957,In_2054,In_2317);
and U4958 (N_4958,In_1645,In_503);
nor U4959 (N_4959,In_1018,In_1282);
nand U4960 (N_4960,In_1093,In_1532);
nand U4961 (N_4961,In_680,In_293);
or U4962 (N_4962,In_2356,In_721);
or U4963 (N_4963,In_1555,In_1381);
or U4964 (N_4964,In_2354,In_1912);
nor U4965 (N_4965,In_1221,In_347);
xnor U4966 (N_4966,In_418,In_625);
or U4967 (N_4967,In_1684,In_232);
nor U4968 (N_4968,In_1114,In_238);
or U4969 (N_4969,In_994,In_1370);
or U4970 (N_4970,In_175,In_929);
or U4971 (N_4971,In_1352,In_1436);
and U4972 (N_4972,In_1501,In_1519);
xnor U4973 (N_4973,In_1368,In_1058);
nand U4974 (N_4974,In_1089,In_765);
or U4975 (N_4975,In_51,In_116);
or U4976 (N_4976,In_595,In_2029);
nand U4977 (N_4977,In_461,In_2014);
and U4978 (N_4978,In_1769,In_1398);
or U4979 (N_4979,In_1581,In_1994);
and U4980 (N_4980,In_2319,In_1664);
or U4981 (N_4981,In_440,In_842);
nand U4982 (N_4982,In_1057,In_1169);
nand U4983 (N_4983,In_1842,In_2300);
xor U4984 (N_4984,In_157,In_228);
and U4985 (N_4985,In_2170,In_344);
or U4986 (N_4986,In_54,In_1997);
xor U4987 (N_4987,In_1363,In_263);
nor U4988 (N_4988,In_640,In_1368);
or U4989 (N_4989,In_1538,In_495);
or U4990 (N_4990,In_1558,In_1347);
and U4991 (N_4991,In_1612,In_2073);
and U4992 (N_4992,In_342,In_1625);
nor U4993 (N_4993,In_1494,In_1596);
and U4994 (N_4994,In_578,In_908);
nor U4995 (N_4995,In_364,In_1738);
nand U4996 (N_4996,In_1042,In_267);
and U4997 (N_4997,In_433,In_1915);
nor U4998 (N_4998,In_445,In_201);
nor U4999 (N_4999,In_2101,In_2037);
nor U5000 (N_5000,N_2116,N_302);
and U5001 (N_5001,N_2940,N_4821);
nor U5002 (N_5002,N_137,N_3881);
nor U5003 (N_5003,N_2976,N_2577);
and U5004 (N_5004,N_2344,N_734);
nor U5005 (N_5005,N_3178,N_632);
and U5006 (N_5006,N_1317,N_2161);
and U5007 (N_5007,N_3296,N_4656);
nor U5008 (N_5008,N_70,N_605);
nor U5009 (N_5009,N_1713,N_2469);
nand U5010 (N_5010,N_3283,N_4599);
or U5011 (N_5011,N_1564,N_206);
nor U5012 (N_5012,N_2311,N_2417);
nand U5013 (N_5013,N_3015,N_2167);
and U5014 (N_5014,N_2025,N_1014);
nor U5015 (N_5015,N_1722,N_4775);
xor U5016 (N_5016,N_701,N_3917);
or U5017 (N_5017,N_1211,N_4046);
nor U5018 (N_5018,N_1562,N_1786);
and U5019 (N_5019,N_2157,N_1436);
and U5020 (N_5020,N_894,N_4432);
or U5021 (N_5021,N_1382,N_2759);
nor U5022 (N_5022,N_3447,N_3575);
and U5023 (N_5023,N_4238,N_167);
nand U5024 (N_5024,N_2140,N_4163);
nor U5025 (N_5025,N_1956,N_3517);
nand U5026 (N_5026,N_2018,N_3840);
nand U5027 (N_5027,N_843,N_4928);
or U5028 (N_5028,N_2009,N_1172);
nand U5029 (N_5029,N_313,N_1711);
xor U5030 (N_5030,N_3603,N_1648);
or U5031 (N_5031,N_4191,N_3003);
nor U5032 (N_5032,N_2591,N_2388);
nor U5033 (N_5033,N_986,N_3953);
or U5034 (N_5034,N_1576,N_456);
xor U5035 (N_5035,N_2557,N_2599);
and U5036 (N_5036,N_4883,N_3698);
nor U5037 (N_5037,N_2284,N_4858);
and U5038 (N_5038,N_3272,N_3353);
or U5039 (N_5039,N_1838,N_1578);
and U5040 (N_5040,N_3251,N_4183);
nor U5041 (N_5041,N_3907,N_1961);
and U5042 (N_5042,N_4275,N_3045);
and U5043 (N_5043,N_3910,N_2463);
or U5044 (N_5044,N_3487,N_3906);
nor U5045 (N_5045,N_3853,N_4882);
or U5046 (N_5046,N_3723,N_2154);
or U5047 (N_5047,N_882,N_1470);
and U5048 (N_5048,N_4819,N_4353);
nand U5049 (N_5049,N_2912,N_176);
nand U5050 (N_5050,N_985,N_2088);
nor U5051 (N_5051,N_1764,N_328);
nand U5052 (N_5052,N_2455,N_284);
or U5053 (N_5053,N_980,N_4859);
nor U5054 (N_5054,N_612,N_2673);
nand U5055 (N_5055,N_2805,N_3512);
or U5056 (N_5056,N_267,N_2792);
nand U5057 (N_5057,N_4936,N_2176);
nand U5058 (N_5058,N_3266,N_2510);
and U5059 (N_5059,N_2272,N_1738);
nor U5060 (N_5060,N_4388,N_3809);
nand U5061 (N_5061,N_1502,N_3959);
nor U5062 (N_5062,N_3616,N_4184);
nor U5063 (N_5063,N_1015,N_3792);
and U5064 (N_5064,N_4422,N_2137);
and U5065 (N_5065,N_1141,N_1773);
nand U5066 (N_5066,N_1131,N_3529);
and U5067 (N_5067,N_2627,N_3510);
and U5068 (N_5068,N_3882,N_2499);
nand U5069 (N_5069,N_2521,N_3238);
nor U5070 (N_5070,N_2776,N_4547);
or U5071 (N_5071,N_4538,N_1928);
or U5072 (N_5072,N_1695,N_433);
or U5073 (N_5073,N_4055,N_3531);
nor U5074 (N_5074,N_752,N_2808);
nor U5075 (N_5075,N_4808,N_1352);
and U5076 (N_5076,N_3685,N_144);
and U5077 (N_5077,N_3320,N_178);
and U5078 (N_5078,N_3765,N_4109);
or U5079 (N_5079,N_2551,N_1124);
nor U5080 (N_5080,N_3502,N_4826);
or U5081 (N_5081,N_2346,N_1781);
nor U5082 (N_5082,N_604,N_3795);
nand U5083 (N_5083,N_4169,N_368);
or U5084 (N_5084,N_3637,N_2078);
nor U5085 (N_5085,N_50,N_124);
nand U5086 (N_5086,N_3051,N_2429);
or U5087 (N_5087,N_510,N_647);
nor U5088 (N_5088,N_4241,N_2491);
nand U5089 (N_5089,N_2714,N_3684);
or U5090 (N_5090,N_2538,N_2489);
nor U5091 (N_5091,N_3337,N_1278);
nor U5092 (N_5092,N_3576,N_3965);
nand U5093 (N_5093,N_1453,N_3035);
or U5094 (N_5094,N_1539,N_3639);
or U5095 (N_5095,N_3432,N_3362);
nand U5096 (N_5096,N_3008,N_264);
and U5097 (N_5097,N_4701,N_4968);
xnor U5098 (N_5098,N_1255,N_1431);
nor U5099 (N_5099,N_1637,N_3268);
nor U5100 (N_5100,N_4799,N_4279);
and U5101 (N_5101,N_4494,N_3503);
nand U5102 (N_5102,N_2664,N_3781);
nand U5103 (N_5103,N_1831,N_3478);
and U5104 (N_5104,N_4822,N_3636);
nand U5105 (N_5105,N_3799,N_2563);
and U5106 (N_5106,N_1231,N_3562);
or U5107 (N_5107,N_4631,N_1173);
nor U5108 (N_5108,N_3345,N_2804);
nor U5109 (N_5109,N_2782,N_1684);
nor U5110 (N_5110,N_4291,N_785);
or U5111 (N_5111,N_873,N_4651);
nor U5112 (N_5112,N_4919,N_1507);
nand U5113 (N_5113,N_1816,N_3434);
nand U5114 (N_5114,N_3674,N_2688);
nor U5115 (N_5115,N_991,N_4776);
nand U5116 (N_5116,N_746,N_3845);
and U5117 (N_5117,N_3108,N_1440);
nand U5118 (N_5118,N_1777,N_2820);
nand U5119 (N_5119,N_690,N_697);
and U5120 (N_5120,N_2327,N_1366);
nand U5121 (N_5121,N_641,N_591);
or U5122 (N_5122,N_1282,N_3394);
nor U5123 (N_5123,N_3229,N_324);
and U5124 (N_5124,N_1441,N_3941);
nor U5125 (N_5125,N_4188,N_1088);
and U5126 (N_5126,N_3293,N_3679);
or U5127 (N_5127,N_1159,N_721);
nor U5128 (N_5128,N_4827,N_4528);
nand U5129 (N_5129,N_2197,N_3821);
and U5130 (N_5130,N_447,N_2106);
or U5131 (N_5131,N_1027,N_4354);
and U5132 (N_5132,N_2317,N_3729);
and U5133 (N_5133,N_2210,N_3547);
nor U5134 (N_5134,N_2155,N_374);
and U5135 (N_5135,N_891,N_2692);
and U5136 (N_5136,N_2486,N_3996);
nor U5137 (N_5137,N_4125,N_2244);
or U5138 (N_5138,N_966,N_2497);
and U5139 (N_5139,N_2373,N_1292);
or U5140 (N_5140,N_2592,N_4932);
nor U5141 (N_5141,N_3280,N_2370);
nand U5142 (N_5142,N_4645,N_2836);
nor U5143 (N_5143,N_1257,N_12);
nand U5144 (N_5144,N_2614,N_1752);
and U5145 (N_5145,N_4954,N_3314);
xnor U5146 (N_5146,N_55,N_2515);
nor U5147 (N_5147,N_2462,N_3618);
nor U5148 (N_5148,N_3905,N_552);
nor U5149 (N_5149,N_2293,N_2694);
nand U5150 (N_5150,N_4802,N_3082);
nand U5151 (N_5151,N_3085,N_2606);
nand U5152 (N_5152,N_2775,N_326);
or U5153 (N_5153,N_3165,N_1508);
xnor U5154 (N_5154,N_1300,N_2299);
and U5155 (N_5155,N_805,N_4282);
and U5156 (N_5156,N_1647,N_45);
and U5157 (N_5157,N_2477,N_10);
and U5158 (N_5158,N_3683,N_476);
and U5159 (N_5159,N_2956,N_4722);
and U5160 (N_5160,N_1705,N_1817);
nor U5161 (N_5161,N_2934,N_1858);
and U5162 (N_5162,N_2487,N_1936);
and U5163 (N_5163,N_4490,N_2230);
or U5164 (N_5164,N_3744,N_3405);
nor U5165 (N_5165,N_3805,N_502);
and U5166 (N_5166,N_1630,N_4708);
and U5167 (N_5167,N_4863,N_3895);
nand U5168 (N_5168,N_3756,N_2132);
nor U5169 (N_5169,N_2642,N_530);
nand U5170 (N_5170,N_1567,N_2800);
and U5171 (N_5171,N_4004,N_3484);
and U5172 (N_5172,N_4330,N_2020);
or U5173 (N_5173,N_3156,N_3014);
or U5174 (N_5174,N_297,N_14);
or U5175 (N_5175,N_25,N_2412);
or U5176 (N_5176,N_1718,N_883);
or U5177 (N_5177,N_3589,N_835);
and U5178 (N_5178,N_4262,N_2849);
nor U5179 (N_5179,N_881,N_2000);
nor U5180 (N_5180,N_2198,N_32);
nand U5181 (N_5181,N_4710,N_3220);
or U5182 (N_5182,N_3592,N_1566);
nor U5183 (N_5183,N_3587,N_1560);
nor U5184 (N_5184,N_3339,N_2022);
nand U5185 (N_5185,N_4966,N_2646);
and U5186 (N_5186,N_2368,N_2689);
and U5187 (N_5187,N_3469,N_546);
and U5188 (N_5188,N_2514,N_3284);
nand U5189 (N_5189,N_846,N_3368);
or U5190 (N_5190,N_1809,N_1298);
or U5191 (N_5191,N_2962,N_379);
and U5192 (N_5192,N_3520,N_3292);
xnor U5193 (N_5193,N_3951,N_3412);
nand U5194 (N_5194,N_1391,N_4982);
xor U5195 (N_5195,N_3149,N_3141);
nand U5196 (N_5196,N_2335,N_1098);
or U5197 (N_5197,N_2558,N_973);
nand U5198 (N_5198,N_1519,N_2982);
nor U5199 (N_5199,N_4771,N_1148);
and U5200 (N_5200,N_3753,N_1156);
xor U5201 (N_5201,N_1602,N_3931);
and U5202 (N_5202,N_4894,N_1247);
nor U5203 (N_5203,N_4495,N_4187);
or U5204 (N_5204,N_4349,N_1716);
nand U5205 (N_5205,N_2798,N_2286);
nor U5206 (N_5206,N_4663,N_2325);
nand U5207 (N_5207,N_4769,N_2861);
and U5208 (N_5208,N_1673,N_2602);
or U5209 (N_5209,N_4890,N_889);
nor U5210 (N_5210,N_4669,N_2064);
or U5211 (N_5211,N_2439,N_4694);
nand U5212 (N_5212,N_2931,N_2677);
and U5213 (N_5213,N_3159,N_2447);
nand U5214 (N_5214,N_2850,N_4586);
nor U5215 (N_5215,N_2493,N_1772);
and U5216 (N_5216,N_3092,N_662);
or U5217 (N_5217,N_4854,N_917);
nor U5218 (N_5218,N_1360,N_1422);
and U5219 (N_5219,N_2616,N_3103);
nand U5220 (N_5220,N_4329,N_2651);
or U5221 (N_5221,N_961,N_1108);
nand U5222 (N_5222,N_2250,N_316);
or U5223 (N_5223,N_2179,N_2188);
nor U5224 (N_5224,N_3312,N_1070);
nor U5225 (N_5225,N_2217,N_1723);
and U5226 (N_5226,N_808,N_3173);
or U5227 (N_5227,N_4247,N_2997);
and U5228 (N_5228,N_4094,N_4480);
nor U5229 (N_5229,N_4618,N_4611);
nor U5230 (N_5230,N_4502,N_2552);
nand U5231 (N_5231,N_1877,N_4934);
nand U5232 (N_5232,N_4491,N_926);
or U5233 (N_5233,N_3209,N_250);
nor U5234 (N_5234,N_1586,N_892);
and U5235 (N_5235,N_4104,N_3902);
nor U5236 (N_5236,N_1275,N_953);
or U5237 (N_5237,N_4174,N_3114);
nor U5238 (N_5238,N_1209,N_3979);
nor U5239 (N_5239,N_1009,N_3399);
or U5240 (N_5240,N_3939,N_971);
xor U5241 (N_5241,N_1867,N_668);
and U5242 (N_5242,N_3331,N_575);
or U5243 (N_5243,N_2669,N_249);
nand U5244 (N_5244,N_3676,N_4462);
and U5245 (N_5245,N_1756,N_908);
nor U5246 (N_5246,N_1934,N_3742);
nor U5247 (N_5247,N_3052,N_3814);
and U5248 (N_5248,N_3946,N_3525);
nand U5249 (N_5249,N_511,N_3461);
or U5250 (N_5250,N_79,N_1324);
nor U5251 (N_5251,N_794,N_3303);
nor U5252 (N_5252,N_1251,N_394);
nor U5253 (N_5253,N_2726,N_312);
or U5254 (N_5254,N_3214,N_941);
or U5255 (N_5255,N_1910,N_4851);
and U5256 (N_5256,N_547,N_4395);
and U5257 (N_5257,N_2619,N_560);
nor U5258 (N_5258,N_3380,N_3010);
or U5259 (N_5259,N_3697,N_4469);
or U5260 (N_5260,N_899,N_221);
and U5261 (N_5261,N_1994,N_2957);
nor U5262 (N_5262,N_1952,N_2095);
nand U5263 (N_5263,N_2833,N_1557);
and U5264 (N_5264,N_3334,N_764);
or U5265 (N_5265,N_2522,N_3803);
nand U5266 (N_5266,N_1907,N_350);
or U5267 (N_5267,N_4182,N_4561);
nand U5268 (N_5268,N_1672,N_1457);
nor U5269 (N_5269,N_938,N_1375);
xor U5270 (N_5270,N_2754,N_253);
nand U5271 (N_5271,N_758,N_2475);
and U5272 (N_5272,N_1397,N_367);
or U5273 (N_5273,N_4552,N_2948);
nand U5274 (N_5274,N_85,N_2605);
and U5275 (N_5275,N_900,N_2452);
or U5276 (N_5276,N_2911,N_2654);
or U5277 (N_5277,N_3271,N_3187);
nor U5278 (N_5278,N_2995,N_4584);
or U5279 (N_5279,N_2513,N_3068);
and U5280 (N_5280,N_3908,N_1398);
xor U5281 (N_5281,N_2548,N_2334);
nand U5282 (N_5282,N_4804,N_4481);
and U5283 (N_5283,N_2693,N_1524);
nor U5284 (N_5284,N_1083,N_673);
and U5285 (N_5285,N_3059,N_3648);
and U5286 (N_5286,N_4419,N_3629);
or U5287 (N_5287,N_755,N_2525);
or U5288 (N_5288,N_2432,N_1686);
nor U5289 (N_5289,N_509,N_431);
nand U5290 (N_5290,N_1693,N_335);
nand U5291 (N_5291,N_2363,N_3340);
or U5292 (N_5292,N_887,N_3160);
or U5293 (N_5293,N_3100,N_3501);
and U5294 (N_5294,N_2937,N_308);
and U5295 (N_5295,N_2969,N_1212);
and U5296 (N_5296,N_2291,N_3689);
nor U5297 (N_5297,N_2001,N_845);
nand U5298 (N_5298,N_698,N_597);
and U5299 (N_5299,N_4306,N_1265);
or U5300 (N_5300,N_2853,N_3956);
nor U5301 (N_5301,N_1077,N_3568);
nor U5302 (N_5302,N_3414,N_566);
and U5303 (N_5303,N_291,N_2947);
nor U5304 (N_5304,N_4199,N_4497);
nand U5305 (N_5305,N_1370,N_563);
nand U5306 (N_5306,N_1343,N_1926);
or U5307 (N_5307,N_1549,N_4766);
nor U5308 (N_5308,N_4088,N_2319);
nand U5309 (N_5309,N_271,N_2738);
nand U5310 (N_5310,N_3577,N_4782);
nand U5311 (N_5311,N_2013,N_1622);
nand U5312 (N_5312,N_2361,N_2277);
or U5313 (N_5313,N_1978,N_40);
or U5314 (N_5314,N_4844,N_2594);
nor U5315 (N_5315,N_2015,N_3384);
and U5316 (N_5316,N_3675,N_2952);
nand U5317 (N_5317,N_2090,N_163);
nor U5318 (N_5318,N_133,N_1226);
xnor U5319 (N_5319,N_4704,N_3087);
and U5320 (N_5320,N_204,N_714);
and U5321 (N_5321,N_1061,N_2946);
and U5322 (N_5322,N_2415,N_4849);
nor U5323 (N_5323,N_1848,N_1101);
or U5324 (N_5324,N_3890,N_4325);
nor U5325 (N_5325,N_1902,N_2381);
nor U5326 (N_5326,N_4718,N_2281);
nor U5327 (N_5327,N_469,N_4272);
or U5328 (N_5328,N_381,N_2129);
nor U5329 (N_5329,N_3217,N_4042);
nand U5330 (N_5330,N_1921,N_1719);
nor U5331 (N_5331,N_342,N_1168);
nand U5332 (N_5332,N_4452,N_2348);
nor U5333 (N_5333,N_3395,N_988);
nand U5334 (N_5334,N_3761,N_2019);
and U5335 (N_5335,N_130,N_2035);
or U5336 (N_5336,N_2970,N_4794);
or U5337 (N_5337,N_4970,N_3573);
or U5338 (N_5338,N_4758,N_161);
nor U5339 (N_5339,N_3826,N_3772);
and U5340 (N_5340,N_3535,N_460);
and U5341 (N_5341,N_531,N_4433);
nor U5342 (N_5342,N_2148,N_3766);
nor U5343 (N_5343,N_299,N_489);
and U5344 (N_5344,N_4671,N_1914);
nand U5345 (N_5345,N_3474,N_548);
xnor U5346 (N_5346,N_730,N_88);
and U5347 (N_5347,N_118,N_2332);
and U5348 (N_5348,N_4106,N_2668);
and U5349 (N_5349,N_377,N_1019);
nor U5350 (N_5350,N_3570,N_3633);
and U5351 (N_5351,N_1183,N_4783);
or U5352 (N_5352,N_2186,N_4043);
nand U5353 (N_5353,N_2908,N_3888);
and U5354 (N_5354,N_4909,N_4439);
or U5355 (N_5355,N_3600,N_1332);
nand U5356 (N_5356,N_4472,N_702);
nor U5357 (N_5357,N_3724,N_1891);
or U5358 (N_5358,N_3594,N_4870);
nor U5359 (N_5359,N_98,N_1214);
and U5360 (N_5360,N_2187,N_3126);
nand U5361 (N_5361,N_1469,N_4348);
and U5362 (N_5362,N_3006,N_454);
and U5363 (N_5363,N_3460,N_4172);
nand U5364 (N_5364,N_4999,N_4972);
or U5365 (N_5365,N_67,N_2678);
nor U5366 (N_5366,N_1444,N_3228);
nand U5367 (N_5367,N_363,N_1644);
xnor U5368 (N_5368,N_658,N_387);
and U5369 (N_5369,N_2769,N_2181);
or U5370 (N_5370,N_2285,N_1465);
and U5371 (N_5371,N_2834,N_4421);
and U5372 (N_5372,N_2533,N_3976);
nand U5373 (N_5373,N_4546,N_3690);
nand U5374 (N_5374,N_169,N_3222);
nor U5375 (N_5375,N_611,N_617);
nor U5376 (N_5376,N_4655,N_4166);
or U5377 (N_5377,N_3523,N_432);
nor U5378 (N_5378,N_4099,N_196);
or U5379 (N_5379,N_3071,N_457);
xor U5380 (N_5380,N_4990,N_2943);
nand U5381 (N_5381,N_666,N_3133);
and U5382 (N_5382,N_2802,N_1030);
nor U5383 (N_5383,N_4114,N_2162);
and U5384 (N_5384,N_417,N_2556);
and U5385 (N_5385,N_871,N_492);
nand U5386 (N_5386,N_1002,N_3347);
and U5387 (N_5387,N_772,N_2199);
nor U5388 (N_5388,N_4813,N_1732);
and U5389 (N_5389,N_3192,N_1966);
nor U5390 (N_5390,N_4406,N_2454);
or U5391 (N_5391,N_3248,N_844);
or U5392 (N_5392,N_4730,N_4324);
nor U5393 (N_5393,N_3877,N_1948);
and U5394 (N_5394,N_3249,N_42);
or U5395 (N_5395,N_1830,N_1859);
or U5396 (N_5396,N_4378,N_107);
or U5397 (N_5397,N_896,N_3104);
or U5398 (N_5398,N_315,N_2502);
and U5399 (N_5399,N_4624,N_4877);
nand U5400 (N_5400,N_754,N_1822);
or U5401 (N_5401,N_2876,N_2519);
or U5402 (N_5402,N_4597,N_4654);
and U5403 (N_5403,N_784,N_3958);
and U5404 (N_5404,N_3370,N_4012);
xnor U5405 (N_5405,N_2691,N_713);
nor U5406 (N_5406,N_3163,N_1774);
or U5407 (N_5407,N_2227,N_4386);
or U5408 (N_5408,N_868,N_352);
nor U5409 (N_5409,N_287,N_3274);
and U5410 (N_5410,N_4375,N_2017);
and U5411 (N_5411,N_2953,N_3921);
or U5412 (N_5412,N_4759,N_652);
or U5413 (N_5413,N_1771,N_2053);
and U5414 (N_5414,N_2892,N_4953);
and U5415 (N_5415,N_1526,N_2965);
and U5416 (N_5416,N_4818,N_1601);
or U5417 (N_5417,N_728,N_4603);
nand U5418 (N_5418,N_2667,N_19);
nor U5419 (N_5419,N_864,N_614);
nor U5420 (N_5420,N_2873,N_227);
and U5421 (N_5421,N_4872,N_1536);
nor U5422 (N_5422,N_2471,N_849);
nand U5423 (N_5423,N_2607,N_2930);
xor U5424 (N_5424,N_1048,N_1091);
nor U5425 (N_5425,N_4665,N_202);
nand U5426 (N_5426,N_3123,N_3208);
and U5427 (N_5427,N_885,N_2909);
and U5428 (N_5428,N_2567,N_3672);
and U5429 (N_5429,N_3566,N_2003);
nand U5430 (N_5430,N_2821,N_990);
and U5431 (N_5431,N_4788,N_4196);
nand U5432 (N_5432,N_3657,N_1260);
nor U5433 (N_5433,N_2219,N_570);
and U5434 (N_5434,N_1748,N_4786);
or U5435 (N_5435,N_2404,N_4357);
and U5436 (N_5436,N_924,N_4261);
nor U5437 (N_5437,N_4344,N_3210);
nor U5438 (N_5438,N_4724,N_403);
nand U5439 (N_5439,N_3865,N_185);
nor U5440 (N_5440,N_1938,N_654);
xor U5441 (N_5441,N_4642,N_4628);
and U5442 (N_5442,N_15,N_4503);
or U5443 (N_5443,N_3462,N_3021);
or U5444 (N_5444,N_1186,N_3360);
nor U5445 (N_5445,N_427,N_3140);
and U5446 (N_5446,N_1592,N_2774);
or U5447 (N_5447,N_1074,N_272);
nand U5448 (N_5448,N_593,N_4307);
and U5449 (N_5449,N_2762,N_2818);
or U5450 (N_5450,N_2643,N_3327);
or U5451 (N_5451,N_4500,N_4956);
and U5452 (N_5452,N_4684,N_3367);
nor U5453 (N_5453,N_1242,N_435);
nand U5454 (N_5454,N_4937,N_481);
or U5455 (N_5455,N_4984,N_832);
nand U5456 (N_5456,N_4373,N_709);
and U5457 (N_5457,N_1374,N_397);
and U5458 (N_5458,N_3544,N_4699);
nand U5459 (N_5459,N_1707,N_708);
and U5460 (N_5460,N_2245,N_1708);
or U5461 (N_5461,N_1862,N_3704);
nor U5462 (N_5462,N_418,N_886);
or U5463 (N_5463,N_465,N_3654);
nor U5464 (N_5464,N_1217,N_4607);
nor U5465 (N_5465,N_2099,N_4218);
nor U5466 (N_5466,N_464,N_4935);
or U5467 (N_5467,N_1449,N_321);
nor U5468 (N_5468,N_4234,N_3851);
and U5469 (N_5469,N_1663,N_16);
or U5470 (N_5470,N_4554,N_2604);
nand U5471 (N_5471,N_1483,N_2215);
and U5472 (N_5472,N_4466,N_1633);
and U5473 (N_5473,N_1339,N_4152);
nand U5474 (N_5474,N_34,N_4311);
nand U5475 (N_5475,N_1906,N_841);
and U5476 (N_5476,N_4839,N_3746);
and U5477 (N_5477,N_3244,N_1059);
or U5478 (N_5478,N_179,N_2758);
nand U5479 (N_5479,N_4942,N_2724);
nor U5480 (N_5480,N_1221,N_1426);
and U5481 (N_5481,N_416,N_1826);
and U5482 (N_5482,N_1581,N_4728);
nor U5483 (N_5483,N_750,N_288);
and U5484 (N_5484,N_4248,N_2270);
or U5485 (N_5485,N_4393,N_4342);
nor U5486 (N_5486,N_1827,N_1500);
and U5487 (N_5487,N_3709,N_1006);
and U5488 (N_5488,N_2712,N_1294);
nor U5489 (N_5489,N_2838,N_1428);
xor U5490 (N_5490,N_2460,N_1573);
nand U5491 (N_5491,N_1204,N_2742);
nor U5492 (N_5492,N_914,N_3144);
nand U5493 (N_5493,N_1041,N_1999);
nor U5494 (N_5494,N_164,N_2052);
or U5495 (N_5495,N_482,N_4750);
and U5496 (N_5496,N_1338,N_4916);
nand U5497 (N_5497,N_289,N_4626);
or U5498 (N_5498,N_2260,N_4292);
nor U5499 (N_5499,N_2222,N_4719);
or U5500 (N_5500,N_3253,N_3233);
or U5501 (N_5501,N_4992,N_49);
or U5502 (N_5502,N_2047,N_2496);
and U5503 (N_5503,N_3352,N_4835);
nor U5504 (N_5504,N_770,N_4154);
nand U5505 (N_5505,N_4873,N_2968);
and U5506 (N_5506,N_4581,N_2073);
and U5507 (N_5507,N_2964,N_1724);
nand U5508 (N_5508,N_2505,N_1314);
and U5509 (N_5509,N_4425,N_3972);
nand U5510 (N_5510,N_1527,N_4170);
and U5511 (N_5511,N_3017,N_2634);
or U5512 (N_5512,N_2376,N_323);
nand U5513 (N_5513,N_4428,N_3801);
nand U5514 (N_5514,N_3341,N_3034);
nand U5515 (N_5515,N_1829,N_1788);
nor U5516 (N_5516,N_4723,N_1692);
or U5517 (N_5517,N_4662,N_4753);
nand U5518 (N_5518,N_2183,N_4267);
nor U5519 (N_5519,N_648,N_1433);
and U5520 (N_5520,N_3670,N_4505);
nand U5521 (N_5521,N_2986,N_1636);
and U5522 (N_5522,N_2784,N_4440);
nand U5523 (N_5523,N_943,N_1776);
nor U5524 (N_5524,N_2587,N_4945);
nand U5525 (N_5525,N_4293,N_3671);
and U5526 (N_5526,N_4738,N_1662);
nand U5527 (N_5527,N_1399,N_1393);
nor U5528 (N_5528,N_2789,N_629);
or U5529 (N_5529,N_2766,N_303);
or U5530 (N_5530,N_4801,N_2296);
or U5531 (N_5531,N_4105,N_2459);
nand U5532 (N_5532,N_1596,N_1997);
nand U5533 (N_5533,N_4674,N_1322);
nor U5534 (N_5534,N_4430,N_2733);
and U5535 (N_5535,N_1065,N_140);
nor U5536 (N_5536,N_4326,N_4039);
nor U5537 (N_5537,N_4098,N_3962);
nor U5538 (N_5538,N_4679,N_3993);
nor U5539 (N_5539,N_2887,N_2872);
nand U5540 (N_5540,N_4764,N_2589);
and U5541 (N_5541,N_4461,N_1749);
and U5542 (N_5542,N_4498,N_3847);
nor U5543 (N_5543,N_3749,N_4841);
and U5544 (N_5544,N_4361,N_2801);
and U5545 (N_5545,N_1658,N_2029);
nand U5546 (N_5546,N_1086,N_3815);
and U5547 (N_5547,N_4486,N_2274);
nor U5548 (N_5548,N_2048,N_682);
or U5549 (N_5549,N_4779,N_1544);
and U5550 (N_5550,N_834,N_166);
xnor U5551 (N_5551,N_3128,N_4424);
nor U5552 (N_5552,N_1797,N_1767);
nand U5553 (N_5553,N_4059,N_829);
nor U5554 (N_5554,N_4637,N_2457);
nor U5555 (N_5555,N_4506,N_372);
and U5556 (N_5556,N_2859,N_2623);
nor U5557 (N_5557,N_3282,N_4785);
and U5558 (N_5558,N_3298,N_2094);
and U5559 (N_5559,N_3361,N_610);
nor U5560 (N_5560,N_2787,N_290);
nand U5561 (N_5561,N_1276,N_4400);
nor U5562 (N_5562,N_2403,N_1710);
or U5563 (N_5563,N_3199,N_2147);
nand U5564 (N_5564,N_1983,N_3830);
nor U5565 (N_5565,N_3752,N_711);
nand U5566 (N_5566,N_4681,N_1402);
and U5567 (N_5567,N_4958,N_2501);
and U5568 (N_5568,N_4925,N_1964);
nand U5569 (N_5569,N_670,N_994);
or U5570 (N_5570,N_1523,N_4852);
and U5571 (N_5571,N_4997,N_1965);
nor U5572 (N_5572,N_964,N_376);
or U5573 (N_5573,N_3376,N_4327);
or U5574 (N_5574,N_3800,N_851);
and U5575 (N_5575,N_3094,N_3287);
and U5576 (N_5576,N_1079,N_1401);
and U5577 (N_5577,N_622,N_329);
and U5578 (N_5578,N_4093,N_1087);
and U5579 (N_5579,N_3596,N_4295);
nand U5580 (N_5580,N_3860,N_3932);
or U5581 (N_5581,N_602,N_4111);
and U5582 (N_5582,N_2727,N_638);
nor U5583 (N_5583,N_850,N_4024);
or U5584 (N_5584,N_3291,N_3528);
nand U5585 (N_5585,N_3348,N_2321);
nor U5586 (N_5586,N_4384,N_3669);
or U5587 (N_5587,N_3755,N_2430);
or U5588 (N_5588,N_3164,N_3707);
or U5589 (N_5589,N_2559,N_4117);
or U5590 (N_5590,N_3063,N_1337);
nand U5591 (N_5591,N_2256,N_1972);
nor U5592 (N_5592,N_1815,N_1166);
and U5593 (N_5593,N_703,N_3236);
or U5594 (N_5594,N_37,N_2647);
nor U5595 (N_5595,N_732,N_3571);
or U5596 (N_5596,N_1750,N_621);
and U5597 (N_5597,N_3393,N_28);
nor U5598 (N_5598,N_997,N_3027);
nor U5599 (N_5599,N_2298,N_4601);
or U5600 (N_5600,N_1555,N_4305);
nor U5601 (N_5601,N_2652,N_3404);
or U5602 (N_5602,N_3967,N_4845);
nor U5603 (N_5603,N_1747,N_2631);
nand U5604 (N_5604,N_421,N_576);
or U5605 (N_5605,N_2959,N_353);
nor U5606 (N_5606,N_4933,N_4565);
or U5607 (N_5607,N_3563,N_2144);
and U5608 (N_5608,N_561,N_3927);
and U5609 (N_5609,N_3617,N_848);
nand U5610 (N_5610,N_1291,N_2406);
or U5611 (N_5611,N_2797,N_545);
or U5612 (N_5612,N_3867,N_1600);
and U5613 (N_5613,N_1514,N_1857);
nor U5614 (N_5614,N_1656,N_4463);
xnor U5615 (N_5615,N_365,N_4855);
and U5616 (N_5616,N_3856,N_491);
nand U5617 (N_5617,N_2889,N_4310);
and U5618 (N_5618,N_3557,N_3829);
nor U5619 (N_5619,N_2936,N_1135);
and U5620 (N_5620,N_967,N_4380);
and U5621 (N_5621,N_3013,N_4058);
nand U5622 (N_5622,N_2212,N_1787);
and U5623 (N_5623,N_2919,N_3869);
nand U5624 (N_5624,N_3161,N_4483);
nor U5625 (N_5625,N_1677,N_1084);
and U5626 (N_5626,N_968,N_2663);
and U5627 (N_5627,N_3306,N_1668);
or U5628 (N_5628,N_1082,N_586);
nand U5629 (N_5629,N_4762,N_4389);
nor U5630 (N_5630,N_2687,N_1890);
or U5631 (N_5631,N_1661,N_1900);
nand U5632 (N_5632,N_1800,N_541);
or U5633 (N_5633,N_1432,N_4897);
or U5634 (N_5634,N_1942,N_1116);
and U5635 (N_5635,N_2338,N_4652);
or U5636 (N_5636,N_1261,N_3301);
and U5637 (N_5637,N_2405,N_558);
nand U5638 (N_5638,N_1880,N_4539);
nor U5639 (N_5639,N_2049,N_2079);
or U5640 (N_5640,N_2612,N_1248);
xor U5641 (N_5641,N_2715,N_1473);
and U5642 (N_5642,N_2295,N_528);
or U5643 (N_5643,N_1240,N_2303);
or U5644 (N_5644,N_1512,N_4436);
xnor U5645 (N_5645,N_1912,N_2150);
or U5646 (N_5646,N_2568,N_3433);
or U5647 (N_5647,N_500,N_279);
nand U5648 (N_5648,N_660,N_4787);
nor U5649 (N_5649,N_2736,N_3049);
and U5650 (N_5650,N_3553,N_4902);
or U5651 (N_5651,N_810,N_2490);
or U5652 (N_5652,N_823,N_4733);
and U5653 (N_5653,N_2927,N_2353);
and U5654 (N_5654,N_2610,N_1147);
nand U5655 (N_5655,N_1290,N_4233);
nand U5656 (N_5656,N_1144,N_4271);
or U5657 (N_5657,N_2435,N_3791);
or U5658 (N_5658,N_3398,N_2699);
nand U5659 (N_5659,N_1023,N_935);
nand U5660 (N_5660,N_4853,N_3099);
nand U5661 (N_5661,N_1712,N_2832);
or U5662 (N_5662,N_743,N_3446);
xor U5663 (N_5663,N_2231,N_4559);
nand U5664 (N_5664,N_817,N_1273);
nor U5665 (N_5665,N_4355,N_927);
nand U5666 (N_5666,N_2067,N_1957);
or U5667 (N_5667,N_1510,N_2749);
and U5668 (N_5668,N_2958,N_1207);
or U5669 (N_5669,N_2397,N_1157);
nand U5670 (N_5670,N_1753,N_340);
nor U5671 (N_5671,N_1413,N_824);
nand U5672 (N_5672,N_2939,N_3152);
and U5673 (N_5673,N_1215,N_4101);
and U5674 (N_5674,N_479,N_3719);
nor U5675 (N_5675,N_11,N_4450);
or U5676 (N_5676,N_819,N_2280);
nand U5677 (N_5677,N_1986,N_2991);
nor U5678 (N_5678,N_4341,N_322);
or U5679 (N_5679,N_4833,N_3113);
or U5680 (N_5680,N_1933,N_3497);
and U5681 (N_5681,N_3254,N_2683);
nor U5682 (N_5682,N_1482,N_1281);
and U5683 (N_5683,N_601,N_4673);
nor U5684 (N_5684,N_4939,N_62);
and U5685 (N_5685,N_2779,N_4115);
and U5686 (N_5686,N_4986,N_4041);
and U5687 (N_5687,N_3005,N_1100);
nor U5688 (N_5688,N_3203,N_1898);
or U5689 (N_5689,N_4073,N_1143);
nor U5690 (N_5690,N_3490,N_3498);
nand U5691 (N_5691,N_360,N_3142);
nand U5692 (N_5692,N_2967,N_618);
or U5693 (N_5693,N_2572,N_4431);
nor U5694 (N_5694,N_183,N_590);
and U5695 (N_5695,N_3473,N_2575);
nor U5696 (N_5696,N_2184,N_2881);
and U5697 (N_5697,N_856,N_2225);
nand U5698 (N_5698,N_3441,N_4198);
nand U5699 (N_5699,N_170,N_759);
and U5700 (N_5700,N_3451,N_634);
or U5701 (N_5701,N_4917,N_1000);
and U5702 (N_5702,N_3224,N_20);
and U5703 (N_5703,N_1554,N_224);
nor U5704 (N_5704,N_4398,N_4834);
nor U5705 (N_5705,N_675,N_485);
nor U5706 (N_5706,N_4437,N_3396);
and U5707 (N_5707,N_695,N_3688);
or U5708 (N_5708,N_4752,N_2998);
and U5709 (N_5709,N_677,N_2509);
or U5710 (N_5710,N_3409,N_2845);
and U5711 (N_5711,N_3667,N_3621);
nand U5712 (N_5712,N_4377,N_2037);
and U5713 (N_5713,N_3053,N_9);
nor U5714 (N_5714,N_2924,N_556);
nand U5715 (N_5715,N_4300,N_207);
nand U5716 (N_5716,N_1923,N_788);
nor U5717 (N_5717,N_1452,N_3770);
or U5718 (N_5718,N_3785,N_2810);
nor U5719 (N_5719,N_2372,N_3950);
and U5720 (N_5720,N_1028,N_2772);
nor U5721 (N_5721,N_2815,N_2);
nor U5722 (N_5722,N_2343,N_226);
and U5723 (N_5723,N_4625,N_3836);
nor U5724 (N_5724,N_3262,N_1970);
or U5725 (N_5725,N_1799,N_3721);
nor U5726 (N_5726,N_223,N_145);
nand U5727 (N_5727,N_2474,N_958);
nor U5728 (N_5728,N_1365,N_1798);
and U5729 (N_5729,N_4593,N_244);
nor U5730 (N_5730,N_2767,N_4121);
nor U5731 (N_5731,N_2237,N_4053);
nand U5732 (N_5732,N_4455,N_3107);
nor U5733 (N_5733,N_818,N_111);
xnor U5734 (N_5734,N_4850,N_2822);
or U5735 (N_5735,N_3453,N_1851);
nand U5736 (N_5736,N_661,N_916);
and U5737 (N_5737,N_2114,N_4768);
nor U5738 (N_5738,N_3922,N_1495);
nand U5739 (N_5739,N_3515,N_4967);
or U5740 (N_5740,N_884,N_1714);
or U5741 (N_5741,N_1595,N_2618);
and U5742 (N_5742,N_4582,N_3537);
or U5743 (N_5743,N_521,N_2629);
and U5744 (N_5744,N_2825,N_2266);
nand U5745 (N_5745,N_386,N_4369);
nor U5746 (N_5746,N_1381,N_3556);
or U5747 (N_5747,N_2300,N_1377);
and U5748 (N_5748,N_3762,N_4901);
and U5749 (N_5749,N_4413,N_3841);
and U5750 (N_5750,N_3852,N_1454);
nand U5751 (N_5751,N_4809,N_4071);
and U5752 (N_5752,N_1804,N_1669);
or U5753 (N_5753,N_3355,N_274);
and U5754 (N_5754,N_4866,N_311);
nand U5755 (N_5755,N_1176,N_930);
nand U5756 (N_5756,N_2941,N_4633);
nand U5757 (N_5757,N_3022,N_362);
nand U5758 (N_5758,N_104,N_2306);
or U5759 (N_5759,N_1843,N_2470);
and U5760 (N_5760,N_4345,N_2852);
and U5761 (N_5761,N_2865,N_4781);
nand U5762 (N_5762,N_1356,N_486);
and U5763 (N_5763,N_203,N_95);
or U5764 (N_5764,N_4757,N_283);
nor U5765 (N_5765,N_1760,N_3640);
nand U5766 (N_5766,N_1863,N_1531);
and U5767 (N_5767,N_1540,N_2516);
or U5768 (N_5768,N_1238,N_659);
or U5769 (N_5769,N_4221,N_2464);
nor U5770 (N_5770,N_97,N_2275);
and U5771 (N_5771,N_1227,N_1163);
nor U5772 (N_5772,N_2074,N_1384);
or U5773 (N_5773,N_2626,N_963);
nand U5774 (N_5774,N_1990,N_4533);
and U5775 (N_5775,N_2422,N_1670);
or U5776 (N_5776,N_1197,N_1613);
and U5777 (N_5777,N_4442,N_4190);
nand U5778 (N_5778,N_3763,N_2292);
and U5779 (N_5779,N_4396,N_3481);
nor U5780 (N_5780,N_689,N_3227);
nor U5781 (N_5781,N_3387,N_4672);
nand U5782 (N_5782,N_2315,N_2110);
and U5783 (N_5783,N_2142,N_4996);
nor U5784 (N_5784,N_3550,N_606);
or U5785 (N_5785,N_932,N_2428);
and U5786 (N_5786,N_2146,N_1054);
nand U5787 (N_5787,N_4445,N_270);
nor U5788 (N_5788,N_1119,N_2786);
nand U5789 (N_5789,N_1739,N_2811);
nor U5790 (N_5790,N_1599,N_2640);
nand U5791 (N_5791,N_3645,N_3263);
and U5792 (N_5792,N_3782,N_1878);
nor U5793 (N_5793,N_1080,N_2590);
nand U5794 (N_5794,N_645,N_643);
nand U5795 (N_5795,N_3130,N_1188);
and U5796 (N_5796,N_4613,N_1114);
nor U5797 (N_5797,N_1796,N_1085);
and U5798 (N_5798,N_2550,N_4717);
or U5799 (N_5799,N_2021,N_1060);
nand U5800 (N_5800,N_2200,N_2287);
or U5801 (N_5801,N_2914,N_2662);
or U5802 (N_5802,N_2910,N_2989);
xor U5803 (N_5803,N_44,N_4688);
or U5804 (N_5804,N_2290,N_2051);
or U5805 (N_5805,N_3514,N_2745);
and U5806 (N_5806,N_429,N_2921);
or U5807 (N_5807,N_3538,N_1477);
and U5808 (N_5808,N_948,N_1055);
and U5809 (N_5809,N_2751,N_1580);
nor U5810 (N_5810,N_3310,N_4230);
nor U5811 (N_5811,N_1140,N_2310);
and U5812 (N_5812,N_978,N_1805);
nor U5813 (N_5813,N_1813,N_2333);
nor U5814 (N_5814,N_3030,N_3041);
and U5815 (N_5815,N_1743,N_4596);
or U5816 (N_5816,N_977,N_1844);
and U5817 (N_5817,N_4739,N_2520);
nand U5818 (N_5818,N_3886,N_1618);
or U5819 (N_5819,N_2273,N_3868);
nor U5820 (N_5820,N_796,N_355);
or U5821 (N_5821,N_4510,N_862);
and U5822 (N_5822,N_1538,N_1224);
and U5823 (N_5823,N_1126,N_4456);
nand U5824 (N_5824,N_2190,N_4382);
nor U5825 (N_5825,N_2324,N_1089);
nor U5826 (N_5826,N_4840,N_3887);
and U5827 (N_5827,N_1625,N_504);
nand U5828 (N_5828,N_3610,N_127);
nand U5829 (N_5829,N_3884,N_4138);
nor U5830 (N_5830,N_75,N_2416);
nor U5831 (N_5831,N_1715,N_4525);
nand U5832 (N_5832,N_4194,N_3169);
nand U5833 (N_5833,N_343,N_676);
nand U5834 (N_5834,N_3424,N_4861);
nand U5835 (N_5835,N_23,N_2529);
nand U5836 (N_5836,N_799,N_4124);
nand U5837 (N_5837,N_1546,N_3970);
nand U5838 (N_5838,N_257,N_2111);
and U5839 (N_5839,N_1492,N_3585);
and U5840 (N_5840,N_2441,N_4256);
nor U5841 (N_5841,N_3036,N_587);
nor U5842 (N_5842,N_47,N_4367);
nand U5843 (N_5843,N_2121,N_94);
nand U5844 (N_5844,N_2523,N_2660);
nor U5845 (N_5845,N_4885,N_525);
and U5846 (N_5846,N_4632,N_3046);
nand U5847 (N_5847,N_4016,N_2598);
nor U5848 (N_5848,N_1325,N_4040);
nor U5849 (N_5849,N_1958,N_2863);
nand U5850 (N_5850,N_4881,N_4368);
or U5851 (N_5851,N_1346,N_102);
nand U5852 (N_5852,N_1123,N_1690);
and U5853 (N_5853,N_26,N_1939);
and U5854 (N_5854,N_1913,N_3075);
nand U5855 (N_5855,N_1390,N_4692);
and U5856 (N_5856,N_1593,N_2842);
and U5857 (N_5857,N_4973,N_657);
and U5858 (N_5858,N_2573,N_2711);
and U5859 (N_5859,N_1770,N_3465);
xor U5860 (N_5860,N_2145,N_3143);
nand U5861 (N_5861,N_4910,N_3505);
nor U5862 (N_5862,N_1769,N_4742);
nor U5863 (N_5863,N_1569,N_2877);
xnor U5864 (N_5864,N_630,N_3696);
or U5865 (N_5865,N_2096,N_3825);
or U5866 (N_5866,N_1272,N_906);
or U5867 (N_5867,N_3835,N_3545);
and U5868 (N_5868,N_3893,N_230);
xnor U5869 (N_5869,N_3904,N_2350);
or U5870 (N_5870,N_443,N_3936);
nand U5871 (N_5871,N_1142,N_4317);
or U5872 (N_5872,N_4438,N_1761);
nand U5873 (N_5873,N_807,N_1697);
or U5874 (N_5874,N_1050,N_1881);
nor U5875 (N_5875,N_194,N_2761);
nor U5876 (N_5876,N_1814,N_3270);
or U5877 (N_5877,N_2044,N_636);
or U5878 (N_5878,N_4475,N_4880);
or U5879 (N_5879,N_3062,N_1745);
and U5880 (N_5880,N_1210,N_325);
nor U5881 (N_5881,N_3864,N_237);
nand U5882 (N_5882,N_4260,N_3191);
xor U5883 (N_5883,N_3466,N_2314);
nand U5884 (N_5884,N_3354,N_1922);
and U5885 (N_5885,N_2109,N_2100);
nand U5886 (N_5886,N_1194,N_3492);
nand U5887 (N_5887,N_1062,N_987);
nor U5888 (N_5888,N_1256,N_1960);
or U5889 (N_5889,N_256,N_753);
nor U5890 (N_5890,N_4713,N_184);
nor U5891 (N_5891,N_615,N_2024);
nor U5892 (N_5892,N_3273,N_946);
xor U5893 (N_5893,N_4900,N_4789);
nand U5894 (N_5894,N_2524,N_2868);
nor U5895 (N_5895,N_2764,N_2732);
nor U5896 (N_5896,N_1998,N_1920);
nand U5897 (N_5897,N_4676,N_285);
and U5898 (N_5898,N_699,N_1892);
nand U5899 (N_5899,N_565,N_4049);
nor U5900 (N_5900,N_4515,N_4884);
and U5901 (N_5901,N_3666,N_1459);
nand U5902 (N_5902,N_1924,N_4703);
and U5903 (N_5903,N_1481,N_422);
and U5904 (N_5904,N_1403,N_512);
and U5905 (N_5905,N_4133,N_4411);
nand U5906 (N_5906,N_4524,N_4680);
nand U5907 (N_5907,N_2453,N_992);
nor U5908 (N_5908,N_2411,N_2152);
nor U5909 (N_5909,N_1590,N_1847);
nor U5910 (N_5910,N_2066,N_960);
nand U5911 (N_5911,N_3439,N_1927);
and U5912 (N_5912,N_1353,N_4028);
or U5913 (N_5913,N_252,N_236);
nand U5914 (N_5914,N_1149,N_74);
nor U5915 (N_5915,N_580,N_2655);
or U5916 (N_5916,N_276,N_4726);
or U5917 (N_5917,N_1947,N_3650);
nor U5918 (N_5918,N_2696,N_1941);
xnor U5919 (N_5919,N_4843,N_2254);
and U5920 (N_5920,N_1702,N_3822);
or U5921 (N_5921,N_4683,N_4165);
nand U5922 (N_5922,N_77,N_2484);
nand U5923 (N_5923,N_448,N_656);
nor U5924 (N_5924,N_3804,N_2632);
or U5925 (N_5925,N_653,N_1355);
nand U5926 (N_5926,N_923,N_3359);
or U5927 (N_5927,N_1266,N_154);
nor U5928 (N_5928,N_2133,N_1202);
and U5929 (N_5929,N_2955,N_205);
and U5930 (N_5930,N_273,N_1794);
nor U5931 (N_5931,N_1901,N_3582);
nand U5932 (N_5932,N_1334,N_4979);
or U5933 (N_5933,N_1350,N_3275);
or U5934 (N_5934,N_4670,N_1834);
nor U5935 (N_5935,N_2593,N_1854);
and U5936 (N_5936,N_2731,N_3336);
xor U5937 (N_5937,N_1057,N_1323);
nand U5938 (N_5938,N_4731,N_4402);
nor U5939 (N_5939,N_4441,N_4685);
or U5940 (N_5940,N_3420,N_3894);
nor U5941 (N_5941,N_3377,N_897);
and U5942 (N_5942,N_2236,N_320);
and U5943 (N_5943,N_3574,N_4541);
and U5944 (N_5944,N_455,N_3839);
and U5945 (N_5945,N_665,N_4682);
and U5946 (N_5946,N_4846,N_132);
nor U5947 (N_5947,N_3281,N_1751);
nand U5948 (N_5948,N_557,N_3769);
nor U5949 (N_5949,N_2635,N_1742);
or U5950 (N_5950,N_4962,N_1329);
nor U5951 (N_5951,N_2888,N_2671);
and U5952 (N_5952,N_878,N_1335);
nand U5953 (N_5953,N_2414,N_4899);
and U5954 (N_5954,N_1262,N_2172);
nor U5955 (N_5955,N_412,N_4964);
nor U5956 (N_5956,N_4507,N_2625);
or U5957 (N_5957,N_4800,N_1003);
nand U5958 (N_5958,N_53,N_867);
xor U5959 (N_5959,N_1783,N_2407);
nor U5960 (N_5960,N_1737,N_1447);
or U5961 (N_5961,N_3074,N_3925);
and U5962 (N_5962,N_493,N_101);
nand U5963 (N_5963,N_4197,N_1996);
nand U5964 (N_5964,N_2974,N_2923);
nor U5965 (N_5965,N_3928,N_3122);
or U5966 (N_5966,N_4038,N_1701);
nor U5967 (N_5967,N_1036,N_4702);
nand U5968 (N_5968,N_4981,N_4030);
and U5969 (N_5969,N_4575,N_4705);
or U5970 (N_5970,N_105,N_936);
nand U5971 (N_5971,N_4185,N_1380);
nand U5972 (N_5972,N_181,N_438);
and U5973 (N_5973,N_306,N_2545);
or U5974 (N_5974,N_3328,N_1832);
or U5975 (N_5975,N_3039,N_4860);
nand U5976 (N_5976,N_4167,N_2320);
xor U5977 (N_5977,N_4540,N_1811);
nand U5978 (N_5978,N_2951,N_2783);
or U5979 (N_5979,N_3506,N_620);
nand U5980 (N_5980,N_501,N_2083);
and U5981 (N_5981,N_970,N_1522);
or U5982 (N_5982,N_3218,N_4010);
and U5983 (N_5983,N_1051,N_4617);
xnor U5984 (N_5984,N_4168,N_156);
nand U5985 (N_5985,N_3823,N_2949);
and U5986 (N_5986,N_1638,N_3480);
nand U5987 (N_5987,N_1122,N_3552);
and U5988 (N_5988,N_3754,N_3472);
and U5989 (N_5989,N_3019,N_298);
xor U5990 (N_5990,N_1201,N_3105);
nand U5991 (N_5991,N_2208,N_775);
nand U5992 (N_5992,N_925,N_696);
nand U5993 (N_5993,N_1045,N_3708);
and U5994 (N_5994,N_1515,N_2994);
nor U5995 (N_5995,N_3174,N_804);
nand U5996 (N_5996,N_246,N_3947);
nand U5997 (N_5997,N_3663,N_1974);
nand U5998 (N_5998,N_3518,N_2086);
nor U5999 (N_5999,N_6,N_293);
nor U6000 (N_6000,N_2423,N_4025);
or U6001 (N_6001,N_382,N_2582);
nor U6002 (N_6002,N_1488,N_2530);
nand U6003 (N_6003,N_2562,N_4914);
or U6004 (N_6004,N_1793,N_3846);
nand U6005 (N_6005,N_2340,N_3158);
and U6006 (N_6006,N_3190,N_761);
nor U6007 (N_6007,N_1871,N_3876);
nor U6008 (N_6008,N_2261,N_4511);
nand U6009 (N_6009,N_4192,N_3680);
nand U6010 (N_6010,N_4555,N_1404);
or U6011 (N_6011,N_2034,N_333);
nand U6012 (N_6012,N_2382,N_2613);
nor U6013 (N_6013,N_278,N_336);
and U6014 (N_6014,N_3295,N_3069);
nand U6015 (N_6015,N_842,N_2351);
and U6016 (N_6016,N_1579,N_3031);
nor U6017 (N_6017,N_783,N_1823);
nand U6018 (N_6018,N_4830,N_2472);
nand U6019 (N_6019,N_2289,N_3638);
nand U6020 (N_6020,N_2579,N_2304);
and U6021 (N_6021,N_3444,N_4178);
xor U6022 (N_6022,N_2702,N_3117);
nor U6023 (N_6023,N_3954,N_3256);
or U6024 (N_6024,N_4868,N_1090);
or U6025 (N_6025,N_477,N_3167);
and U6026 (N_6026,N_1357,N_3132);
nand U6027 (N_6027,N_3598,N_1175);
xor U6028 (N_6028,N_225,N_2448);
nor U6029 (N_6029,N_3317,N_4119);
and U6030 (N_6030,N_2935,N_1446);
or U6031 (N_6031,N_3900,N_2438);
nand U6032 (N_6032,N_3909,N_3811);
nand U6033 (N_6033,N_3661,N_480);
nand U6034 (N_6034,N_4227,N_865);
nor U6035 (N_6035,N_731,N_4620);
nor U6036 (N_6036,N_2135,N_2893);
nor U6037 (N_6037,N_3475,N_2413);
nor U6038 (N_6038,N_2730,N_1296);
nand U6039 (N_6039,N_4714,N_4280);
or U6040 (N_6040,N_261,N_1721);
nand U6041 (N_6041,N_584,N_2444);
or U6042 (N_6042,N_2819,N_330);
nand U6043 (N_6043,N_4026,N_1945);
or U6044 (N_6044,N_4077,N_667);
nor U6045 (N_6045,N_1700,N_282);
or U6046 (N_6046,N_3338,N_2653);
or U6047 (N_6047,N_2164,N_103);
nor U6048 (N_6048,N_3693,N_3549);
nand U6049 (N_6049,N_2799,N_1869);
or U6050 (N_6050,N_4574,N_866);
or U6051 (N_6051,N_3449,N_4622);
or U6052 (N_6052,N_3417,N_452);
and U6053 (N_6053,N_2684,N_4162);
nor U6054 (N_6054,N_3699,N_522);
nor U6055 (N_6055,N_1915,N_567);
nand U6056 (N_6056,N_870,N_255);
or U6057 (N_6057,N_3009,N_3530);
nor U6058 (N_6058,N_2478,N_809);
nand U6059 (N_6059,N_627,N_423);
nand U6060 (N_6060,N_2046,N_174);
nor U6061 (N_6061,N_3358,N_3365);
xnor U6062 (N_6062,N_1845,N_2103);
nor U6063 (N_6063,N_3265,N_3197);
or U6064 (N_6064,N_767,N_4147);
nor U6065 (N_6065,N_1552,N_4145);
or U6066 (N_6066,N_1367,N_3700);
nor U6067 (N_6067,N_4203,N_1435);
nand U6068 (N_6068,N_3079,N_1363);
nand U6069 (N_6069,N_3180,N_4825);
or U6070 (N_6070,N_430,N_2359);
nand U6071 (N_6071,N_2972,N_2011);
xnor U6072 (N_6072,N_3694,N_1616);
nand U6073 (N_6073,N_1642,N_1137);
nor U6074 (N_6074,N_396,N_3418);
nor U6075 (N_6075,N_4941,N_1929);
nor U6076 (N_6076,N_688,N_1551);
and U6077 (N_6077,N_1369,N_4778);
nand U6078 (N_6078,N_3106,N_1192);
nor U6079 (N_6079,N_4770,N_318);
nor U6080 (N_6080,N_3848,N_633);
nand U6081 (N_6081,N_3246,N_2307);
nor U6082 (N_6082,N_1981,N_3564);
nand U6083 (N_6083,N_2117,N_60);
nand U6084 (N_6084,N_4213,N_3258);
nor U6085 (N_6085,N_68,N_4359);
or U6086 (N_6086,N_2143,N_2364);
nor U6087 (N_6087,N_4479,N_1461);
xor U6088 (N_6088,N_1244,N_177);
nand U6089 (N_6089,N_4924,N_2466);
nor U6090 (N_6090,N_1611,N_4258);
or U6091 (N_6091,N_4286,N_4370);
xor U6092 (N_6092,N_2075,N_1005);
and U6093 (N_6093,N_4107,N_2585);
or U6094 (N_6094,N_189,N_120);
and U6095 (N_6095,N_983,N_4186);
or U6096 (N_6096,N_1351,N_1610);
or U6097 (N_6097,N_910,N_87);
nand U6098 (N_6098,N_607,N_1031);
or U6099 (N_6099,N_2443,N_1299);
or U6100 (N_6100,N_4171,N_4257);
and U6101 (N_6101,N_860,N_1424);
nor U6102 (N_6102,N_762,N_373);
nand U6103 (N_6103,N_4451,N_3389);
or U6104 (N_6104,N_1037,N_2978);
nor U6105 (N_6105,N_859,N_1223);
or U6106 (N_6106,N_1709,N_2482);
and U6107 (N_6107,N_2718,N_234);
nor U6108 (N_6108,N_982,N_3750);
nor U6109 (N_6109,N_4980,N_3660);
nand U6110 (N_6110,N_1572,N_3597);
nand U6111 (N_6111,N_4340,N_0);
or U6112 (N_6112,N_51,N_562);
and U6113 (N_6113,N_1025,N_2495);
or U6114 (N_6114,N_3608,N_1899);
or U6115 (N_6115,N_3168,N_2171);
xor U6116 (N_6116,N_141,N_1321);
or U6117 (N_6117,N_200,N_4051);
or U6118 (N_6118,N_2637,N_2880);
or U6119 (N_6119,N_4712,N_3602);
and U6120 (N_6120,N_1553,N_4175);
nor U6121 (N_6121,N_1967,N_1038);
and U6122 (N_6122,N_1795,N_3177);
and U6123 (N_6123,N_1589,N_121);
or U6124 (N_6124,N_1744,N_4760);
and U6125 (N_6125,N_3425,N_4091);
nand U6126 (N_6126,N_4065,N_251);
nand U6127 (N_6127,N_2806,N_2313);
nand U6128 (N_6128,N_3655,N_3402);
and U6129 (N_6129,N_972,N_4960);
nand U6130 (N_6130,N_1302,N_2008);
and U6131 (N_6131,N_1812,N_4251);
nand U6132 (N_6132,N_1909,N_1758);
nor U6133 (N_6133,N_2005,N_1893);
and U6134 (N_6134,N_4015,N_248);
xor U6135 (N_6135,N_2089,N_4871);
nand U6136 (N_6136,N_3631,N_467);
or U6137 (N_6137,N_4155,N_3952);
nand U6138 (N_6138,N_852,N_3234);
and U6139 (N_6139,N_2966,N_1306);
nor U6140 (N_6140,N_334,N_879);
and U6141 (N_6141,N_56,N_4465);
and U6142 (N_6142,N_693,N_4333);
nand U6143 (N_6143,N_1778,N_4116);
nor U6144 (N_6144,N_3378,N_1930);
and U6145 (N_6145,N_1894,N_1988);
or U6146 (N_6146,N_1545,N_956);
nand U6147 (N_6147,N_3802,N_2700);
and U6148 (N_6148,N_4412,N_2905);
nand U6149 (N_6149,N_3842,N_2257);
nand U6150 (N_6150,N_4211,N_2848);
nand U6151 (N_6151,N_4888,N_4407);
nand U6152 (N_6152,N_4974,N_639);
xnor U6153 (N_6153,N_1792,N_3977);
nand U6154 (N_6154,N_4698,N_2855);
and U6155 (N_6155,N_1855,N_1486);
and U6156 (N_6156,N_3247,N_4504);
nor U6157 (N_6157,N_798,N_3448);
and U6158 (N_6158,N_1841,N_3983);
nor U6159 (N_6159,N_2139,N_2576);
or U6160 (N_6160,N_4664,N_1410);
and U6161 (N_6161,N_1394,N_1313);
or U6162 (N_6162,N_1943,N_1004);
and U6163 (N_6163,N_2087,N_4856);
or U6164 (N_6164,N_2755,N_2658);
nor U6165 (N_6165,N_861,N_4416);
nor U6166 (N_6166,N_4499,N_4220);
nor U6167 (N_6167,N_2115,N_1373);
nor U6168 (N_6168,N_4460,N_2175);
and U6169 (N_6169,N_542,N_3991);
nor U6170 (N_6170,N_2488,N_4067);
and U6171 (N_6171,N_4108,N_3632);
or U6172 (N_6172,N_4564,N_517);
and U6173 (N_6173,N_3857,N_880);
and U6174 (N_6174,N_3850,N_1819);
nor U6175 (N_6175,N_4572,N_3778);
or U6176 (N_6176,N_726,N_4204);
nor U6177 (N_6177,N_3200,N_811);
nand U6178 (N_6178,N_4249,N_3426);
and U6179 (N_6179,N_1471,N_3560);
and U6180 (N_6180,N_4600,N_4903);
and U6181 (N_6181,N_822,N_1627);
or U6182 (N_6182,N_3780,N_1621);
nand U6183 (N_6183,N_4159,N_4033);
and U6184 (N_6184,N_1269,N_3896);
or U6185 (N_6185,N_3579,N_3508);
and U6186 (N_6186,N_1307,N_3734);
nand U6187 (N_6187,N_3419,N_4570);
nor U6188 (N_6188,N_2379,N_1977);
nand U6189 (N_6189,N_71,N_663);
nor U6190 (N_6190,N_4896,N_2061);
and U6191 (N_6191,N_582,N_4591);
and U6192 (N_6192,N_1754,N_488);
or U6193 (N_6193,N_2879,N_13);
or U6194 (N_6194,N_72,N_3125);
and U6195 (N_6195,N_243,N_680);
and U6196 (N_6196,N_4392,N_1170);
nand U6197 (N_6197,N_1230,N_3739);
and U6198 (N_6198,N_2010,N_2672);
or U6199 (N_6199,N_3407,N_3838);
nand U6200 (N_6200,N_4097,N_4696);
and U6201 (N_6201,N_2240,N_2977);
and U6202 (N_6202,N_1239,N_2440);
nor U6203 (N_6203,N_478,N_1130);
or U6204 (N_6204,N_1364,N_3875);
and U6205 (N_6205,N_4075,N_537);
xnor U6206 (N_6206,N_2897,N_4217);
or U6207 (N_6207,N_262,N_3308);
and U6208 (N_6208,N_4434,N_535);
or U6209 (N_6209,N_3175,N_4641);
and U6210 (N_6210,N_3787,N_1782);
nand U6211 (N_6211,N_3471,N_2192);
nand U6212 (N_6212,N_155,N_2903);
or U6213 (N_6213,N_739,N_1010);
or U6214 (N_6214,N_4604,N_4120);
nor U6215 (N_6215,N_2481,N_1591);
and U6216 (N_6216,N_1336,N_1763);
nor U6217 (N_6217,N_2004,N_3540);
nor U6218 (N_6218,N_1614,N_2891);
and U6219 (N_6219,N_1687,N_3494);
nor U6220 (N_6220,N_150,N_1659);
and U6221 (N_6221,N_3155,N_4923);
or U6222 (N_6222,N_4889,N_2104);
nor U6223 (N_6223,N_58,N_1072);
xor U6224 (N_6224,N_3555,N_3101);
nor U6225 (N_6225,N_3619,N_3885);
and U6226 (N_6226,N_624,N_2926);
and U6227 (N_6227,N_1604,N_863);
and U6228 (N_6228,N_4549,N_736);
nand U6229 (N_6229,N_409,N_3898);
and U6230 (N_6230,N_1383,N_109);
nand U6231 (N_6231,N_436,N_579);
and U6232 (N_6232,N_933,N_473);
nand U6233 (N_6233,N_3738,N_4022);
or U6234 (N_6234,N_589,N_4869);
nand U6235 (N_6235,N_296,N_1475);
and U6236 (N_6236,N_1612,N_2527);
nand U6237 (N_6237,N_2512,N_3987);
and U6238 (N_6238,N_1220,N_806);
or U6239 (N_6239,N_780,N_4630);
and U6240 (N_6240,N_550,N_1052);
and U6241 (N_6241,N_407,N_1411);
or U6242 (N_6242,N_3595,N_869);
nand U6243 (N_6243,N_4608,N_4725);
or U6244 (N_6244,N_4921,N_3001);
or U6245 (N_6245,N_2633,N_4792);
nand U6246 (N_6246,N_4206,N_4720);
nor U6247 (N_6247,N_833,N_1499);
nor U6248 (N_6248,N_3381,N_2249);
or U6249 (N_6249,N_1937,N_905);
nand U6250 (N_6250,N_3491,N_2721);
or U6251 (N_6251,N_2870,N_2748);
nor U6252 (N_6252,N_3488,N_2125);
nand U6253 (N_6253,N_1665,N_1026);
and U6254 (N_6254,N_1725,N_3879);
nand U6255 (N_6255,N_2492,N_4083);
or U6256 (N_6256,N_4926,N_2701);
nand U6257 (N_6257,N_1868,N_346);
and U6258 (N_6258,N_1846,N_2371);
nor U6259 (N_6259,N_2537,N_213);
or U6260 (N_6260,N_3020,N_3994);
nor U6261 (N_6261,N_157,N_3583);
nand U6262 (N_6262,N_4212,N_1462);
nor U6263 (N_6263,N_3969,N_4294);
and U6264 (N_6264,N_3757,N_266);
nand U6265 (N_6265,N_1046,N_3934);
and U6266 (N_6266,N_4253,N_3000);
nand U6267 (N_6267,N_1150,N_2717);
or U6268 (N_6268,N_4032,N_3330);
nor U6269 (N_6269,N_646,N_1047);
nand U6270 (N_6270,N_4560,N_3423);
nand U6271 (N_6271,N_609,N_1896);
nor U6272 (N_6272,N_4686,N_4567);
nor U6273 (N_6273,N_3593,N_3504);
nand U6274 (N_6274,N_3728,N_4531);
and U6275 (N_6275,N_4949,N_2235);
and U6276 (N_6276,N_1179,N_4740);
and U6277 (N_6277,N_4001,N_3513);
and U6278 (N_6278,N_1480,N_1963);
and U6279 (N_6279,N_484,N_1949);
nor U6280 (N_6280,N_3824,N_2377);
and U6281 (N_6281,N_4905,N_940);
nor U6282 (N_6282,N_153,N_2392);
nor U6283 (N_6283,N_3912,N_1234);
nand U6284 (N_6284,N_347,N_603);
nand U6285 (N_6285,N_3136,N_3613);
and U6286 (N_6286,N_793,N_3604);
and U6287 (N_6287,N_4151,N_821);
nand U6288 (N_6288,N_1280,N_4276);
and U6289 (N_6289,N_4210,N_1288);
or U6290 (N_6290,N_1680,N_3828);
nand U6291 (N_6291,N_3586,N_2954);
nand U6292 (N_6292,N_2151,N_4773);
nor U6293 (N_6293,N_2597,N_4732);
and U6294 (N_6294,N_1109,N_3344);
nor U6295 (N_6295,N_4927,N_3391);
or U6296 (N_6296,N_655,N_679);
nor U6297 (N_6297,N_2709,N_3148);
nor U6298 (N_6298,N_4426,N_1975);
or U6299 (N_6299,N_35,N_4535);
nand U6300 (N_6300,N_544,N_1017);
or U6301 (N_6301,N_1305,N_4405);
or U6302 (N_6302,N_2813,N_3499);
nand U6303 (N_6303,N_4891,N_812);
nand U6304 (N_6304,N_1487,N_2308);
and U6305 (N_6305,N_2178,N_1007);
or U6306 (N_6306,N_2554,N_86);
nor U6307 (N_6307,N_1330,N_2900);
nand U6308 (N_6308,N_398,N_2193);
or U6309 (N_6309,N_2269,N_3691);
nor U6310 (N_6310,N_114,N_3241);
nor U6311 (N_6311,N_3343,N_2925);
and U6312 (N_6312,N_3102,N_54);
nor U6313 (N_6313,N_4749,N_129);
nor U6314 (N_6314,N_4470,N_3911);
nor U6315 (N_6315,N_4379,N_1733);
nand U6316 (N_6316,N_2288,N_912);
or U6317 (N_6317,N_4142,N_3090);
or U6318 (N_6318,N_588,N_2906);
or U6319 (N_6319,N_69,N_2081);
nand U6320 (N_6320,N_4675,N_3854);
or U6321 (N_6321,N_1379,N_2485);
or U6322 (N_6322,N_344,N_4944);
or U6323 (N_6323,N_4487,N_4086);
nand U6324 (N_6324,N_4219,N_4590);
nand U6325 (N_6325,N_171,N_2342);
and U6326 (N_6326,N_2408,N_1962);
or U6327 (N_6327,N_651,N_4269);
or U6328 (N_6328,N_4784,N_1525);
and U6329 (N_6329,N_3002,N_4874);
or U6330 (N_6330,N_981,N_2973);
and U6331 (N_6331,N_3790,N_4079);
nor U6332 (N_6332,N_4235,N_836);
nand U6333 (N_6333,N_4103,N_717);
and U6334 (N_6334,N_756,N_173);
or U6335 (N_6335,N_513,N_1587);
nor U6336 (N_6336,N_4023,N_4222);
or U6337 (N_6337,N_1245,N_2041);
or U6338 (N_6338,N_199,N_3422);
and U6339 (N_6339,N_877,N_1516);
and U6340 (N_6340,N_4790,N_92);
or U6341 (N_6341,N_4517,N_5);
nand U6342 (N_6342,N_3193,N_1973);
nor U6343 (N_6343,N_3,N_4745);
nor U6344 (N_6344,N_30,N_471);
or U6345 (N_6345,N_1146,N_383);
nor U6346 (N_6346,N_3968,N_275);
or U6347 (N_6347,N_2536,N_4020);
xnor U6348 (N_6348,N_749,N_1071);
nand U6349 (N_6349,N_1439,N_3206);
and U6350 (N_6350,N_3767,N_1496);
xnor U6351 (N_6351,N_3793,N_4649);
nand U6352 (N_6352,N_4207,N_1577);
nor U6353 (N_6353,N_974,N_4711);
nor U6354 (N_6354,N_1509,N_4832);
or U6355 (N_6355,N_674,N_4278);
or U6356 (N_6356,N_4435,N_2763);
or U6357 (N_6357,N_3626,N_1528);
nor U6358 (N_6358,N_1917,N_3055);
nor U6359 (N_6359,N_4063,N_847);
nor U6360 (N_6360,N_2258,N_928);
nand U6361 (N_6361,N_2323,N_4302);
nand U6362 (N_6362,N_2920,N_401);
and U6363 (N_6363,N_1916,N_4748);
nand U6364 (N_6364,N_4284,N_4976);
or U6365 (N_6365,N_2426,N_4772);
nand U6366 (N_6366,N_2386,N_2725);
or U6367 (N_6367,N_505,N_3903);
nor U6368 (N_6368,N_2809,N_962);
or U6369 (N_6369,N_1904,N_3311);
nand U6370 (N_6370,N_2984,N_998);
nor U6371 (N_6371,N_1503,N_2055);
and U6372 (N_6372,N_2398,N_1286);
or U6373 (N_6373,N_233,N_4255);
nor U6374 (N_6374,N_3601,N_2596);
or U6375 (N_6375,N_128,N_954);
nand U6376 (N_6376,N_3789,N_4602);
and U6377 (N_6377,N_2322,N_4743);
and U6378 (N_6378,N_1267,N_2494);
nor U6379 (N_6379,N_2827,N_1520);
and U6380 (N_6380,N_1556,N_4285);
or U6381 (N_6381,N_73,N_1361);
or U6382 (N_6382,N_2229,N_3237);
and U6383 (N_6383,N_1969,N_1835);
and U6384 (N_6384,N_1155,N_3813);
or U6385 (N_6385,N_3058,N_2276);
nor U6386 (N_6386,N_3024,N_1284);
or U6387 (N_6387,N_1277,N_2031);
and U6388 (N_6388,N_700,N_3612);
nor U6389 (N_6389,N_3990,N_4904);
or U6390 (N_6390,N_2153,N_3146);
or U6391 (N_6391,N_1837,N_4612);
nand U6392 (N_6392,N_4920,N_2719);
nand U6393 (N_6393,N_4007,N_3060);
or U6394 (N_6394,N_3477,N_751);
nand U6395 (N_6395,N_2068,N_91);
nand U6396 (N_6396,N_441,N_1533);
and U6397 (N_6397,N_1726,N_280);
or U6398 (N_6398,N_2704,N_378);
nand U6399 (N_6399,N_4780,N_1362);
nor U6400 (N_6400,N_2450,N_4715);
or U6401 (N_6401,N_534,N_3764);
nand U6402 (N_6402,N_2535,N_4544);
nand U6403 (N_6403,N_3539,N_497);
nor U6404 (N_6404,N_2638,N_2279);
or U6405 (N_6405,N_3390,N_2644);
and U6406 (N_6406,N_919,N_3527);
nor U6407 (N_6407,N_790,N_4084);
or U6408 (N_6408,N_4464,N_2620);
or U6409 (N_6409,N_3534,N_577);
nor U6410 (N_6410,N_3076,N_3050);
nand U6411 (N_6411,N_4895,N_4842);
nand U6412 (N_6412,N_4060,N_4229);
nand U6413 (N_6413,N_1603,N_4343);
and U6414 (N_6414,N_1995,N_2427);
and U6415 (N_6415,N_3711,N_745);
nand U6416 (N_6416,N_4006,N_814);
nor U6417 (N_6417,N_1985,N_2682);
or U6418 (N_6418,N_3883,N_3716);
or U6419 (N_6419,N_4816,N_3937);
and U6420 (N_6420,N_3533,N_4459);
xnor U6421 (N_6421,N_4308,N_4492);
and U6422 (N_6422,N_2518,N_4864);
nand U6423 (N_6423,N_3300,N_2177);
nor U6424 (N_6424,N_1171,N_1347);
and U6425 (N_6425,N_2770,N_4989);
nand U6426 (N_6426,N_2239,N_3464);
or U6427 (N_6427,N_1504,N_2302);
or U6428 (N_6428,N_3151,N_1547);
or U6429 (N_6429,N_2309,N_1935);
xor U6430 (N_6430,N_2913,N_3196);
nor U6431 (N_6431,N_1032,N_2246);
or U6432 (N_6432,N_3580,N_2158);
nor U6433 (N_6433,N_685,N_96);
or U6434 (N_6434,N_1232,N_840);
nand U6435 (N_6435,N_2262,N_440);
nand U6436 (N_6436,N_277,N_1550);
and U6437 (N_6437,N_3285,N_222);
or U6438 (N_6438,N_2795,N_2480);
or U6439 (N_6439,N_1420,N_951);
and U6440 (N_6440,N_4573,N_4018);
nor U6441 (N_6441,N_3496,N_4774);
and U6442 (N_6442,N_1154,N_2560);
and U6443 (N_6443,N_4356,N_180);
or U6444 (N_6444,N_3942,N_2817);
and U6445 (N_6445,N_4797,N_4598);
and U6446 (N_6446,N_2062,N_2960);
or U6447 (N_6447,N_1706,N_2301);
and U6448 (N_6448,N_678,N_3542);
or U6449 (N_6449,N_538,N_3964);
nor U6450 (N_6450,N_2695,N_4514);
nor U6451 (N_6451,N_3289,N_4226);
nand U6452 (N_6452,N_1884,N_2247);
nand U6453 (N_6453,N_1044,N_3388);
nor U6454 (N_6454,N_2828,N_2739);
or U6455 (N_6455,N_1584,N_1839);
nand U6456 (N_6456,N_1228,N_3097);
nor U6457 (N_6457,N_508,N_4848);
and U6458 (N_6458,N_1191,N_1505);
and U6459 (N_6459,N_301,N_855);
nor U6460 (N_6460,N_3066,N_813);
or U6461 (N_6461,N_3715,N_516);
or U6462 (N_6462,N_837,N_555);
or U6463 (N_6463,N_247,N_1198);
or U6464 (N_6464,N_1396,N_3411);
nor U6465 (N_6465,N_3442,N_2539);
nor U6466 (N_6466,N_4643,N_3810);
or U6467 (N_6467,N_625,N_1850);
nor U6468 (N_6468,N_779,N_2570);
and U6469 (N_6469,N_462,N_89);
nand U6470 (N_6470,N_2981,N_3454);
nor U6471 (N_6471,N_2318,N_3543);
or U6472 (N_6472,N_146,N_38);
nand U6473 (N_6473,N_540,N_3383);
nor U6474 (N_6474,N_4090,N_2916);
and U6475 (N_6475,N_1583,N_187);
and U6476 (N_6476,N_3084,N_572);
and U6477 (N_6477,N_4754,N_3004);
nand U6478 (N_6478,N_549,N_4644);
nor U6479 (N_6479,N_218,N_934);
nor U6480 (N_6480,N_122,N_748);
nand U6481 (N_6481,N_4811,N_2112);
xnor U6482 (N_6482,N_3933,N_2060);
or U6483 (N_6483,N_201,N_3920);
nand U6484 (N_6484,N_4530,N_487);
xor U6485 (N_6485,N_1810,N_1177);
or U6486 (N_6486,N_3131,N_2038);
nand U6487 (N_6487,N_392,N_3321);
or U6488 (N_6488,N_1484,N_2278);
or U6489 (N_6489,N_815,N_2915);
or U6490 (N_6490,N_384,N_131);
or U6491 (N_6491,N_3872,N_4181);
nand U6492 (N_6492,N_3455,N_2698);
and U6493 (N_6493,N_1303,N_984);
nor U6494 (N_6494,N_2336,N_2988);
and U6495 (N_6495,N_4838,N_345);
or U6496 (N_6496,N_2124,N_1327);
nand U6497 (N_6497,N_408,N_1951);
or U6498 (N_6498,N_4550,N_3221);
and U6499 (N_6499,N_3047,N_3701);
and U6500 (N_6500,N_126,N_2753);
or U6501 (N_6501,N_1691,N_1870);
and U6502 (N_6502,N_3373,N_294);
nand U6503 (N_6503,N_2268,N_1011);
or U6504 (N_6504,N_2993,N_1067);
or U6505 (N_6505,N_3923,N_1833);
xnor U6506 (N_6506,N_3786,N_4536);
nand U6507 (N_6507,N_4677,N_490);
nor U6508 (N_6508,N_159,N_3827);
xor U6509 (N_6509,N_3807,N_2383);
nand U6510 (N_6510,N_1008,N_3452);
nand U6511 (N_6511,N_1879,N_4729);
nor U6512 (N_6512,N_1925,N_2232);
and U6513 (N_6513,N_1190,N_3871);
or U6514 (N_6514,N_281,N_2541);
nor U6515 (N_6515,N_613,N_2056);
nand U6516 (N_6516,N_4553,N_4164);
nor U6517 (N_6517,N_3154,N_2168);
or U6518 (N_6518,N_2216,N_2875);
nor U6519 (N_6519,N_2077,N_3652);
or U6520 (N_6520,N_3400,N_268);
and U6521 (N_6521,N_4401,N_3153);
or U6522 (N_6522,N_4128,N_494);
or U6523 (N_6523,N_2352,N_4448);
nand U6524 (N_6524,N_2706,N_2410);
nor U6525 (N_6525,N_771,N_4263);
or U6526 (N_6526,N_2747,N_3988);
or U6527 (N_6527,N_1671,N_4793);
nand U6528 (N_6528,N_2999,N_1852);
or U6529 (N_6529,N_3201,N_3541);
nand U6530 (N_6530,N_193,N_594);
xnor U6531 (N_6531,N_2737,N_4913);
or U6532 (N_6532,N_3935,N_2896);
xnor U6533 (N_6533,N_2697,N_4634);
nand U6534 (N_6534,N_1318,N_3880);
or U6535 (N_6535,N_76,N_4893);
and U6536 (N_6536,N_3630,N_1779);
or U6537 (N_6537,N_4137,N_4019);
nor U6538 (N_6538,N_3410,N_1476);
and U6539 (N_6539,N_3110,N_3299);
or U6540 (N_6540,N_2990,N_391);
or U6541 (N_6541,N_2345,N_2992);
or U6542 (N_6542,N_331,N_2113);
or U6543 (N_6543,N_2564,N_2883);
nor U6544 (N_6544,N_4011,N_1416);
nand U6545 (N_6545,N_3726,N_3641);
and U6546 (N_6546,N_1105,N_554);
nor U6547 (N_6547,N_4756,N_3302);
nor U6548 (N_6548,N_3548,N_995);
or U6549 (N_6549,N_854,N_238);
nor U6550 (N_6550,N_3794,N_4648);
nor U6551 (N_6551,N_3546,N_3961);
nor U6552 (N_6552,N_2773,N_619);
and U6553 (N_6553,N_2574,N_4482);
and U6554 (N_6554,N_2944,N_989);
or U6555 (N_6555,N_1160,N_4940);
and U6556 (N_6556,N_920,N_7);
nor U6557 (N_6557,N_4144,N_781);
nor U6558 (N_6558,N_3294,N_1931);
nor U6559 (N_6559,N_3668,N_2390);
or U6560 (N_6560,N_4501,N_2105);
and U6561 (N_6561,N_4527,N_1442);
nor U6562 (N_6562,N_543,N_4959);
and U6563 (N_6563,N_4817,N_4957);
xnor U6564 (N_6564,N_4153,N_3476);
and U6565 (N_6565,N_3584,N_4453);
nor U6566 (N_6566,N_2902,N_3350);
and U6567 (N_6567,N_706,N_424);
nand U6568 (N_6568,N_415,N_532);
or U6569 (N_6569,N_4952,N_1458);
or U6570 (N_6570,N_3662,N_3415);
and U6571 (N_6571,N_3205,N_1342);
nor U6572 (N_6572,N_3751,N_1802);
and U6573 (N_6573,N_2189,N_3558);
nand U6574 (N_6574,N_1164,N_1095);
and U6575 (N_6575,N_2356,N_380);
nor U6576 (N_6576,N_2420,N_1468);
nand U6577 (N_6577,N_216,N_2756);
and U6578 (N_6578,N_922,N_1415);
and U6579 (N_6579,N_2617,N_106);
and U6580 (N_6580,N_692,N_4141);
nand U6581 (N_6581,N_3678,N_769);
nor U6582 (N_6582,N_1073,N_1840);
nand U6583 (N_6583,N_3138,N_2622);
nand U6584 (N_6584,N_691,N_3245);
and U6585 (N_6585,N_64,N_1081);
and U6586 (N_6586,N_2128,N_1940);
nand U6587 (N_6587,N_1652,N_944);
or U6588 (N_6588,N_4474,N_4027);
or U6589 (N_6589,N_4316,N_3783);
xor U6590 (N_6590,N_4080,N_2012);
nand U6591 (N_6591,N_3007,N_57);
and U6592 (N_6592,N_348,N_3240);
nand U6593 (N_6593,N_3369,N_519);
and U6594 (N_6594,N_3758,N_4000);
and U6595 (N_6595,N_2014,N_3940);
or U6596 (N_6596,N_4478,N_2220);
xnor U6597 (N_6597,N_466,N_1856);
nor U6598 (N_6598,N_3532,N_2253);
or U6599 (N_6599,N_2757,N_410);
and U6600 (N_6600,N_2107,N_4545);
xor U6601 (N_6601,N_3157,N_1660);
and U6602 (N_6602,N_2072,N_2248);
nand U6603 (N_6603,N_573,N_1400);
nor U6604 (N_6604,N_1293,N_1136);
or U6605 (N_6605,N_1182,N_4735);
nand U6606 (N_6606,N_1167,N_686);
or U6607 (N_6607,N_1623,N_820);
or U6608 (N_6608,N_3862,N_3428);
nor U6609 (N_6609,N_188,N_1467);
nor U6610 (N_6610,N_3073,N_1606);
and U6611 (N_6611,N_411,N_82);
nand U6612 (N_6612,N_1803,N_370);
or U6613 (N_6613,N_2791,N_3335);
or U6614 (N_6614,N_1498,N_4737);
and U6615 (N_6615,N_1094,N_1184);
nand U6616 (N_6616,N_245,N_3771);
nand U6617 (N_6617,N_1174,N_4496);
nand U6618 (N_6618,N_650,N_683);
or U6619 (N_6619,N_2816,N_2027);
nor U6620 (N_6620,N_3025,N_339);
and U6621 (N_6621,N_1728,N_965);
and U6622 (N_6622,N_1617,N_2790);
or U6623 (N_6623,N_2864,N_4193);
xor U6624 (N_6624,N_2621,N_4237);
xnor U6625 (N_6625,N_2807,N_2223);
or U6626 (N_6626,N_2609,N_3279);
nand U6627 (N_6627,N_4556,N_1316);
or U6628 (N_6628,N_3703,N_3960);
nor U6629 (N_6629,N_2656,N_3736);
and U6630 (N_6630,N_2233,N_4467);
nor U6631 (N_6631,N_2716,N_2894);
nand U6632 (N_6632,N_3356,N_1106);
nor U6633 (N_6633,N_3986,N_2378);
nor U6634 (N_6634,N_4319,N_3861);
nand U6635 (N_6635,N_1645,N_3486);
nand U6636 (N_6636,N_671,N_3463);
and U6637 (N_6637,N_2241,N_259);
nand U6638 (N_6638,N_681,N_3086);
nand U6639 (N_6639,N_3182,N_718);
nor U6640 (N_6640,N_4592,N_125);
nor U6641 (N_6641,N_258,N_551);
and U6642 (N_6642,N_1532,N_3207);
and U6643 (N_6643,N_1558,N_195);
nor U6644 (N_6644,N_4403,N_1651);
and U6645 (N_6645,N_4646,N_3382);
nor U6646 (N_6646,N_3083,N_172);
or U6647 (N_6647,N_1605,N_2857);
or U6648 (N_6648,N_1430,N_2963);
or U6649 (N_6649,N_3091,N_608);
and U6650 (N_6650,N_2674,N_4383);
nand U6651 (N_6651,N_254,N_4806);
nand U6652 (N_6652,N_1570,N_2456);
or U6653 (N_6653,N_3818,N_672);
nand U6654 (N_6654,N_3072,N_3718);
and U6655 (N_6655,N_2141,N_3385);
and U6656 (N_6656,N_175,N_3834);
and U6657 (N_6657,N_3870,N_2126);
nor U6658 (N_6658,N_4358,N_4372);
and U6659 (N_6659,N_737,N_4399);
nor U6660 (N_6660,N_1521,N_2649);
and U6661 (N_6661,N_3297,N_959);
nand U6662 (N_6662,N_4876,N_2713);
nand U6663 (N_6663,N_260,N_2846);
and U6664 (N_6664,N_1218,N_3176);
xnor U6665 (N_6665,N_720,N_3088);
and U6666 (N_6666,N_1989,N_4619);
or U6667 (N_6667,N_3250,N_1423);
nor U6668 (N_6668,N_4691,N_1022);
or U6669 (N_6669,N_1043,N_1189);
or U6670 (N_6670,N_3999,N_3018);
or U6671 (N_6671,N_2393,N_1791);
nor U6672 (N_6672,N_2546,N_950);
and U6673 (N_6673,N_215,N_4955);
or U6674 (N_6674,N_3305,N_3260);
and U6675 (N_6675,N_147,N_1392);
nor U6676 (N_6676,N_2534,N_3313);
or U6677 (N_6677,N_2265,N_4047);
nor U6678 (N_6678,N_4447,N_1349);
nand U6679 (N_6679,N_1069,N_1585);
nand U6680 (N_6680,N_3235,N_4148);
nand U6681 (N_6681,N_3067,N_496);
nand U6682 (N_6682,N_2517,N_3955);
nor U6683 (N_6683,N_684,N_3445);
and U6684 (N_6684,N_1666,N_975);
nand U6685 (N_6685,N_3677,N_4157);
nand U6686 (N_6686,N_2093,N_4298);
xnor U6687 (N_6687,N_1058,N_3483);
and U6688 (N_6688,N_3622,N_1864);
xor U6689 (N_6689,N_585,N_3139);
or U6690 (N_6690,N_911,N_3915);
nor U6691 (N_6691,N_3121,N_4948);
nor U6692 (N_6692,N_4415,N_2996);
nor U6693 (N_6693,N_2659,N_2708);
nor U6694 (N_6694,N_1634,N_3109);
nor U6695 (N_6695,N_2549,N_100);
nand U6696 (N_6696,N_3225,N_1807);
or U6697 (N_6697,N_4074,N_3033);
nor U6698 (N_6698,N_4288,N_4488);
nand U6699 (N_6699,N_2347,N_3957);
and U6700 (N_6700,N_3665,N_4522);
nor U6701 (N_6701,N_2119,N_2238);
nand U6702 (N_6702,N_1650,N_2528);
nand U6703 (N_6703,N_61,N_1472);
nor U6704 (N_6704,N_2803,N_3706);
or U6705 (N_6705,N_4044,N_1376);
nor U6706 (N_6706,N_2641,N_4716);
nor U6707 (N_6707,N_1162,N_1535);
nand U6708 (N_6708,N_1861,N_1029);
and U6709 (N_6709,N_4214,N_1565);
nand U6710 (N_6710,N_1491,N_1315);
xor U6711 (N_6711,N_4493,N_4371);
and U6712 (N_6712,N_2728,N_2483);
nor U6713 (N_6713,N_1021,N_4606);
and U6714 (N_6714,N_3216,N_3457);
and U6715 (N_6715,N_3048,N_1388);
or U6716 (N_6716,N_2214,N_1053);
and U6717 (N_6717,N_766,N_4610);
nor U6718 (N_6718,N_2503,N_2829);
nand U6719 (N_6719,N_186,N_2436);
and U6720 (N_6720,N_740,N_3628);
nor U6721 (N_6721,N_3264,N_664);
and U6722 (N_6722,N_3985,N_1200);
and U6723 (N_6723,N_2788,N_337);
or U6724 (N_6724,N_623,N_4374);
nor U6725 (N_6725,N_2768,N_4231);
and U6726 (N_6726,N_2156,N_1785);
nor U6727 (N_6727,N_2744,N_1908);
xor U6728 (N_6728,N_307,N_2419);
and U6729 (N_6729,N_1649,N_3949);
and U6730 (N_6730,N_3189,N_4409);
nand U6731 (N_6731,N_419,N_3832);
nor U6732 (N_6732,N_1236,N_4886);
nor U6733 (N_6733,N_4338,N_533);
and U6734 (N_6734,N_2282,N_292);
nor U6735 (N_6735,N_2070,N_1759);
nor U6736 (N_6736,N_4621,N_2367);
or U6737 (N_6737,N_4347,N_4477);
nor U6738 (N_6738,N_4201,N_3290);
nand U6739 (N_6739,N_795,N_2561);
nor U6740 (N_6740,N_1887,N_4150);
and U6741 (N_6741,N_3185,N_3166);
xnor U6742 (N_6742,N_802,N_3524);
nand U6743 (N_6743,N_1698,N_4085);
or U6744 (N_6744,N_4824,N_2476);
nand U6745 (N_6745,N_4381,N_4578);
or U6746 (N_6746,N_4659,N_3276);
nand U6747 (N_6747,N_2297,N_1225);
or U6748 (N_6748,N_4887,N_1406);
and U6749 (N_6749,N_113,N_2866);
or U6750 (N_6750,N_2785,N_3997);
nand U6751 (N_6751,N_445,N_3722);
nor U6752 (N_6752,N_414,N_3656);
nand U6753 (N_6753,N_3467,N_2899);
and U6754 (N_6754,N_3916,N_4823);
or U6755 (N_6755,N_3681,N_2002);
and U6756 (N_6756,N_4562,N_2645);
nand U6757 (N_6757,N_4577,N_2023);
nand U6758 (N_6758,N_1825,N_4697);
and U6759 (N_6759,N_4239,N_3171);
nor U6760 (N_6760,N_3798,N_2134);
nand U6761 (N_6761,N_468,N_3975);
nor U6762 (N_6762,N_3054,N_4687);
or U6763 (N_6763,N_4489,N_2234);
nand U6764 (N_6764,N_2071,N_4509);
or U6765 (N_6765,N_4519,N_4865);
and U6766 (N_6766,N_1571,N_3430);
and U6767 (N_6767,N_2980,N_942);
nor U6768 (N_6768,N_710,N_3397);
or U6769 (N_6769,N_913,N_149);
and U6770 (N_6770,N_3040,N_644);
nor U6771 (N_6771,N_309,N_2504);
or U6772 (N_6772,N_4837,N_4313);
and U6773 (N_6773,N_4176,N_1421);
nand U6774 (N_6774,N_2895,N_3038);
and U6775 (N_6775,N_2506,N_4112);
nand U6776 (N_6776,N_4320,N_1295);
nand U6777 (N_6777,N_446,N_22);
or U6778 (N_6778,N_4089,N_3551);
nor U6779 (N_6779,N_4123,N_3620);
nand U6780 (N_6780,N_1409,N_3644);
nor U6781 (N_6781,N_2123,N_2740);
nand U6782 (N_6782,N_1485,N_3324);
nor U6783 (N_6783,N_2856,N_1982);
or U6784 (N_6784,N_3819,N_4129);
or U6785 (N_6785,N_1354,N_4287);
and U6786 (N_6786,N_1195,N_119);
nor U6787 (N_6787,N_359,N_3204);
or U6788 (N_6788,N_4410,N_3057);
nor U6789 (N_6789,N_4523,N_3326);
nor U6790 (N_6790,N_228,N_420);
nor U6791 (N_6791,N_4057,N_2874);
nor U6792 (N_6792,N_3733,N_3307);
nand U6793 (N_6793,N_1801,N_915);
or U6794 (N_6794,N_459,N_3837);
or U6795 (N_6795,N_4289,N_1755);
or U6796 (N_6796,N_574,N_2793);
or U6797 (N_6797,N_4216,N_2101);
and U6798 (N_6798,N_4056,N_2365);
and U6799 (N_6799,N_1035,N_4635);
nand U6800 (N_6800,N_4290,N_4245);
and U6801 (N_6801,N_4471,N_1389);
and U6802 (N_6802,N_4589,N_3784);
and U6803 (N_6803,N_3588,N_2305);
and U6804 (N_6804,N_3408,N_1679);
and U6805 (N_6805,N_117,N_3495);
nand U6806 (N_6806,N_235,N_2425);
and U6807 (N_6807,N_3743,N_1253);
nand U6808 (N_6808,N_2710,N_1024);
or U6809 (N_6809,N_2271,N_1443);
nand U6810 (N_6810,N_437,N_2878);
nand U6811 (N_6811,N_3259,N_160);
or U6812 (N_6812,N_2735,N_4994);
or U6813 (N_6813,N_1479,N_4473);
nand U6814 (N_6814,N_1161,N_1609);
or U6815 (N_6815,N_2871,N_803);
nand U6816 (N_6816,N_1746,N_539);
nor U6817 (N_6817,N_3653,N_1107);
and U6818 (N_6818,N_3269,N_2169);
or U6819 (N_6819,N_385,N_1992);
and U6820 (N_6820,N_1717,N_3427);
nor U6821 (N_6821,N_4332,N_304);
nand U6822 (N_6822,N_1372,N_4616);
or U6823 (N_6823,N_4134,N_3329);
nand U6824 (N_6824,N_428,N_4064);
nor U6825 (N_6825,N_4977,N_1328);
nand U6826 (N_6826,N_229,N_2526);
nand U6827 (N_6827,N_2394,N_136);
or U6828 (N_6828,N_2252,N_4350);
nand U6829 (N_6829,N_3379,N_4529);
nor U6830 (N_6830,N_2182,N_2312);
nor U6831 (N_6831,N_148,N_4243);
nand U6832 (N_6832,N_1741,N_393);
nand U6833 (N_6833,N_2401,N_1066);
nor U6834 (N_6834,N_3634,N_4054);
and U6835 (N_6835,N_3226,N_1808);
or U6836 (N_6836,N_2544,N_3526);
and U6837 (N_6837,N_3760,N_39);
nand U6838 (N_6838,N_1824,N_3304);
and U6839 (N_6839,N_4629,N_2898);
or U6840 (N_6840,N_483,N_3181);
nor U6841 (N_6841,N_3500,N_723);
xnor U6842 (N_6842,N_1919,N_458);
xor U6843 (N_6843,N_1345,N_2326);
or U6844 (N_6844,N_3732,N_3971);
and U6845 (N_6845,N_83,N_1115);
or U6846 (N_6846,N_4136,N_4143);
nand U6847 (N_6847,N_1478,N_2581);
or U6848 (N_6848,N_24,N_3817);
nand U6849 (N_6849,N_4946,N_1903);
and U6850 (N_6850,N_1918,N_2283);
nand U6851 (N_6851,N_1543,N_2741);
and U6852 (N_6852,N_143,N_2166);
or U6853 (N_6853,N_3119,N_1129);
nor U6854 (N_6854,N_2036,N_857);
or U6855 (N_6855,N_1437,N_4297);
and U6856 (N_6856,N_4476,N_1113);
or U6857 (N_6857,N_3198,N_4796);
or U6858 (N_6858,N_1387,N_4661);
or U6859 (N_6859,N_3607,N_3243);
and U6860 (N_6860,N_1976,N_2869);
nand U6861 (N_6861,N_2201,N_4557);
nor U6862 (N_6862,N_4127,N_4242);
nor U6863 (N_6863,N_1096,N_3554);
and U6864 (N_6864,N_2185,N_529);
or U6865 (N_6865,N_2360,N_2316);
nor U6866 (N_6866,N_2375,N_2039);
nor U6867 (N_6867,N_1534,N_404);
and U6868 (N_6868,N_4678,N_108);
or U6869 (N_6869,N_1460,N_2202);
or U6870 (N_6870,N_4336,N_2975);
nor U6871 (N_6871,N_1099,N_559);
nor U6872 (N_6872,N_777,N_4950);
nand U6873 (N_6873,N_1263,N_3747);
or U6874 (N_6874,N_858,N_4975);
nand U6875 (N_6875,N_2069,N_1312);
or U6876 (N_6876,N_4334,N_1968);
and U6877 (N_6877,N_2127,N_4002);
or U6878 (N_6878,N_4721,N_3134);
and U6879 (N_6879,N_1740,N_4568);
or U6880 (N_6880,N_2765,N_1598);
and U6881 (N_6881,N_3943,N_1243);
nor U6882 (N_6882,N_999,N_1118);
or U6883 (N_6883,N_463,N_4569);
nor U6884 (N_6884,N_640,N_3963);
nand U6885 (N_6885,N_1731,N_2584);
nor U6886 (N_6886,N_4576,N_2780);
and U6887 (N_6887,N_116,N_1784);
nand U6888 (N_6888,N_220,N_4518);
xnor U6889 (N_6889,N_4700,N_4205);
nand U6890 (N_6890,N_4337,N_2680);
xor U6891 (N_6891,N_3966,N_3435);
and U6892 (N_6892,N_3945,N_4930);
or U6893 (N_6893,N_4454,N_2507);
and U6894 (N_6894,N_3456,N_319);
or U6895 (N_6895,N_1,N_2979);
nor U6896 (N_6896,N_366,N_2583);
nor U6897 (N_6897,N_3215,N_4828);
or U6898 (N_6898,N_4036,N_3702);
and U6899 (N_6899,N_3322,N_2251);
nand U6900 (N_6900,N_4647,N_719);
or U6901 (N_6901,N_1076,N_4364);
nand U6902 (N_6902,N_1427,N_2666);
nand U6903 (N_6903,N_402,N_1429);
nand U6904 (N_6904,N_1412,N_2091);
nand U6905 (N_6905,N_4444,N_4657);
nand U6906 (N_6906,N_4240,N_776);
or U6907 (N_6907,N_3162,N_1828);
nand U6908 (N_6908,N_123,N_400);
and U6909 (N_6909,N_890,N_4879);
or U6910 (N_6910,N_1657,N_425);
and U6911 (N_6911,N_2409,N_1049);
nand U6912 (N_6912,N_2130,N_4139);
and U6913 (N_6913,N_168,N_2330);
and U6914 (N_6914,N_4807,N_1905);
or U6915 (N_6915,N_1954,N_3745);
nor U6916 (N_6916,N_4805,N_3740);
nand U6917 (N_6917,N_903,N_3863);
nand U6918 (N_6918,N_1103,N_2636);
and U6919 (N_6919,N_3914,N_3037);
nor U6920 (N_6920,N_197,N_4005);
nand U6921 (N_6921,N_4266,N_4947);
xnor U6922 (N_6922,N_413,N_338);
and U6923 (N_6923,N_1068,N_1185);
nand U6924 (N_6924,N_4003,N_4965);
nor U6925 (N_6925,N_2479,N_3309);
or U6926 (N_6926,N_4301,N_3223);
nor U6927 (N_6927,N_4512,N_3325);
and U6928 (N_6928,N_1405,N_786);
or U6929 (N_6929,N_4668,N_2547);
nand U6930 (N_6930,N_1955,N_4160);
nand U6931 (N_6931,N_2752,N_41);
xnor U6932 (N_6932,N_1619,N_2603);
nor U6933 (N_6933,N_1517,N_2387);
nor U6934 (N_6934,N_4427,N_1674);
or U6935 (N_6935,N_3682,N_2661);
and U6936 (N_6936,N_3776,N_4690);
nand U6937 (N_6937,N_4767,N_4908);
xnor U6938 (N_6938,N_475,N_2159);
and U6939 (N_6939,N_4315,N_3874);
nand U6940 (N_6940,N_1542,N_2228);
nor U6941 (N_6941,N_3416,N_18);
nand U6942 (N_6942,N_1268,N_3219);
and U6943 (N_6943,N_354,N_1821);
nor U6944 (N_6944,N_3647,N_3741);
xor U6945 (N_6945,N_3319,N_2831);
or U6946 (N_6946,N_1494,N_2945);
and U6947 (N_6947,N_3901,N_4180);
and U6948 (N_6948,N_1237,N_3458);
nor U6949 (N_6949,N_1889,N_4580);
and U6950 (N_6950,N_1727,N_2170);
nand U6951 (N_6951,N_3831,N_3124);
and U6952 (N_6952,N_1734,N_269);
nor U6953 (N_6953,N_898,N_760);
or U6954 (N_6954,N_568,N_2860);
and U6955 (N_6955,N_1818,N_1319);
or U6956 (N_6956,N_4791,N_4878);
nand U6957 (N_6957,N_3777,N_1408);
and U6958 (N_6958,N_4707,N_1235);
nand U6959 (N_6959,N_3521,N_4951);
nor U6960 (N_6960,N_63,N_4076);
and U6961 (N_6961,N_1959,N_2259);
nor U6962 (N_6962,N_3357,N_3695);
and U6963 (N_6963,N_406,N_744);
nor U6964 (N_6964,N_3624,N_564);
or U6965 (N_6965,N_4236,N_722);
and U6966 (N_6966,N_3692,N_1152);
nand U6967 (N_6967,N_4209,N_451);
nand U6968 (N_6968,N_3899,N_4095);
nand U6969 (N_6969,N_4961,N_3468);
and U6970 (N_6970,N_2858,N_4283);
and U6971 (N_6971,N_375,N_872);
nand U6972 (N_6972,N_1911,N_1289);
nor U6973 (N_6973,N_3470,N_715);
or U6974 (N_6974,N_4898,N_2294);
xor U6975 (N_6975,N_929,N_1608);
nand U6976 (N_6976,N_4035,N_4658);
and U6977 (N_6977,N_4309,N_3995);
nand U6978 (N_6978,N_495,N_1395);
nor U6979 (N_6979,N_1358,N_191);
and U6980 (N_6980,N_4252,N_3687);
or U6981 (N_6981,N_2211,N_2854);
or U6982 (N_6982,N_4362,N_4906);
or U6983 (N_6983,N_27,N_2778);
nand U6984 (N_6984,N_2242,N_1643);
or U6985 (N_6985,N_792,N_4246);
nor U6986 (N_6986,N_3386,N_1445);
and U6987 (N_6987,N_2006,N_1187);
or U6988 (N_6988,N_2033,N_2690);
nor U6989 (N_6989,N_3374,N_1886);
xnor U6990 (N_6990,N_3643,N_4918);
or U6991 (N_6991,N_4034,N_2337);
and U6992 (N_6992,N_2929,N_3129);
and U6993 (N_6993,N_571,N_876);
nand U6994 (N_6994,N_3042,N_4365);
nand U6995 (N_6995,N_2531,N_4741);
nor U6996 (N_6996,N_642,N_1110);
nand U6997 (N_6997,N_4543,N_1104);
nand U6998 (N_6998,N_3278,N_265);
or U6999 (N_6999,N_765,N_4605);
or U7000 (N_7000,N_1541,N_3375);
nand U7001 (N_7001,N_3712,N_1206);
and U7002 (N_7002,N_4224,N_4296);
nor U7003 (N_7003,N_4417,N_2624);
or U7004 (N_7004,N_3438,N_4339);
nor U7005 (N_7005,N_4110,N_1865);
nor U7006 (N_7006,N_4931,N_2389);
nand U7007 (N_7007,N_4734,N_4215);
nor U7008 (N_7008,N_3255,N_1872);
nand U7009 (N_7009,N_1953,N_2569);
nand U7010 (N_7010,N_3998,N_3179);
xor U7011 (N_7011,N_507,N_993);
nor U7012 (N_7012,N_3808,N_1574);
and U7013 (N_7013,N_3686,N_3774);
nand U7014 (N_7014,N_358,N_789);
or U7015 (N_7015,N_3493,N_2341);
and U7016 (N_7016,N_3366,N_1016);
or U7017 (N_7017,N_1653,N_2615);
nand U7018 (N_7018,N_3080,N_1696);
nand U7019 (N_7019,N_4423,N_390);
or U7020 (N_7020,N_4366,N_1241);
nand U7021 (N_7021,N_31,N_3333);
nand U7022 (N_7022,N_1689,N_4777);
or U7023 (N_7023,N_1639,N_351);
nor U7024 (N_7024,N_1169,N_4232);
nor U7025 (N_7025,N_2595,N_1582);
xor U7026 (N_7026,N_757,N_2224);
nand U7027 (N_7027,N_2194,N_1768);
nand U7028 (N_7028,N_2907,N_1730);
or U7029 (N_7029,N_472,N_1866);
nor U7030 (N_7030,N_1033,N_439);
nor U7031 (N_7031,N_4122,N_4328);
and U7032 (N_7032,N_2136,N_499);
and U7033 (N_7033,N_4516,N_2434);
nor U7034 (N_7034,N_1806,N_2400);
nand U7035 (N_7035,N_2076,N_3735);
nand U7036 (N_7036,N_600,N_2191);
or U7037 (N_7037,N_2498,N_3731);
nor U7038 (N_7038,N_3929,N_3843);
or U7039 (N_7039,N_2750,N_3135);
nor U7040 (N_7040,N_3599,N_135);
nor U7041 (N_7041,N_1466,N_1628);
nor U7042 (N_7042,N_2578,N_1664);
and U7043 (N_7043,N_631,N_3980);
nand U7044 (N_7044,N_725,N_3646);
and U7045 (N_7045,N_2016,N_2843);
nand U7046 (N_7046,N_2421,N_2823);
and U7047 (N_7047,N_1694,N_3044);
nor U7048 (N_7048,N_2396,N_853);
nor U7049 (N_7049,N_2173,N_1685);
and U7050 (N_7050,N_498,N_2473);
and U7051 (N_7051,N_1249,N_4875);
nand U7052 (N_7052,N_3137,N_1145);
nor U7053 (N_7053,N_2442,N_3891);
and U7054 (N_7054,N_4991,N_1888);
nor U7055 (N_7055,N_4693,N_2445);
and U7056 (N_7056,N_4068,N_2555);
and U7057 (N_7057,N_3172,N_4484);
nand U7058 (N_7058,N_1624,N_2532);
or U7059 (N_7059,N_3098,N_444);
nor U7060 (N_7060,N_2630,N_4650);
and U7061 (N_7061,N_4857,N_461);
xnor U7062 (N_7062,N_3892,N_93);
or U7063 (N_7063,N_3078,N_3938);
and U7064 (N_7064,N_2122,N_2045);
nand U7065 (N_7065,N_3118,N_838);
nor U7066 (N_7066,N_211,N_3982);
nand U7067 (N_7067,N_3516,N_2628);
nor U7068 (N_7068,N_1222,N_4418);
nor U7069 (N_7069,N_4971,N_2950);
nand U7070 (N_7070,N_2508,N_3614);
nor U7071 (N_7071,N_1075,N_3974);
nor U7072 (N_7072,N_1133,N_2796);
nor U7073 (N_7073,N_165,N_4736);
or U7074 (N_7074,N_4653,N_1001);
nand U7075 (N_7075,N_3252,N_4929);
nor U7076 (N_7076,N_1311,N_59);
and U7077 (N_7077,N_4763,N_3992);
nand U7078 (N_7078,N_1259,N_2424);
nor U7079 (N_7079,N_4588,N_1309);
and U7080 (N_7080,N_4915,N_1456);
and U7081 (N_7081,N_1513,N_1151);
or U7082 (N_7082,N_592,N_4408);
and U7083 (N_7083,N_1063,N_4404);
nand U7084 (N_7084,N_3346,N_1252);
nor U7085 (N_7085,N_1326,N_2467);
and U7086 (N_7086,N_1340,N_1842);
or U7087 (N_7087,N_1153,N_4566);
and U7088 (N_7088,N_1213,N_1853);
nor U7089 (N_7089,N_3332,N_4534);
nand U7090 (N_7090,N_286,N_2839);
nand U7091 (N_7091,N_2043,N_1506);
nor U7092 (N_7092,N_1128,N_831);
or U7093 (N_7093,N_3913,N_569);
nor U7094 (N_7094,N_4429,N_707);
nand U7095 (N_7095,N_4113,N_1165);
nand U7096 (N_7096,N_3833,N_2542);
nor U7097 (N_7097,N_4815,N_4795);
and U7098 (N_7098,N_2705,N_2933);
or U7099 (N_7099,N_2391,N_1676);
nand U7100 (N_7100,N_830,N_506);
or U7101 (N_7101,N_3673,N_874);
and U7102 (N_7102,N_3413,N_4706);
and U7103 (N_7103,N_839,N_735);
nor U7104 (N_7104,N_1735,N_3581);
nor U7105 (N_7105,N_1984,N_3779);
nor U7106 (N_7106,N_1434,N_3485);
or U7107 (N_7107,N_4609,N_2209);
and U7108 (N_7108,N_4847,N_1615);
and U7109 (N_7109,N_1093,N_1417);
or U7110 (N_7110,N_2812,N_2851);
nand U7111 (N_7111,N_36,N_2830);
and U7112 (N_7112,N_2082,N_3351);
and U7113 (N_7113,N_357,N_4998);
xnor U7114 (N_7114,N_2771,N_2160);
or U7115 (N_7115,N_4202,N_2665);
or U7116 (N_7116,N_2511,N_1246);
nand U7117 (N_7117,N_2588,N_1678);
or U7118 (N_7118,N_2675,N_4061);
nor U7119 (N_7119,N_4614,N_2040);
or U7120 (N_7120,N_219,N_4627);
and U7121 (N_7121,N_904,N_2395);
nand U7122 (N_7122,N_787,N_3127);
and U7123 (N_7123,N_4087,N_3096);
and U7124 (N_7124,N_3170,N_1683);
nor U7125 (N_7125,N_3572,N_1407);
or U7126 (N_7126,N_2263,N_1125);
and U7127 (N_7127,N_4346,N_2204);
nor U7128 (N_7128,N_2213,N_1178);
nand U7129 (N_7129,N_4867,N_369);
xor U7130 (N_7130,N_1064,N_2120);
nor U7131 (N_7131,N_1139,N_4636);
and U7132 (N_7132,N_3089,N_3844);
or U7133 (N_7133,N_2458,N_4623);
nand U7134 (N_7134,N_2886,N_3859);
and U7135 (N_7135,N_1699,N_1193);
and U7136 (N_7136,N_4363,N_332);
nor U7137 (N_7137,N_2961,N_3717);
and U7138 (N_7138,N_2058,N_4727);
and U7139 (N_7139,N_4223,N_46);
nand U7140 (N_7140,N_341,N_4017);
or U7141 (N_7141,N_3522,N_426);
nor U7142 (N_7142,N_2918,N_4988);
and U7143 (N_7143,N_3511,N_2826);
xnor U7144 (N_7144,N_3093,N_48);
nand U7145 (N_7145,N_3231,N_1895);
nand U7146 (N_7146,N_3820,N_4638);
or U7147 (N_7147,N_909,N_1451);
nand U7148 (N_7148,N_2468,N_1219);
nor U7149 (N_7149,N_1078,N_2328);
or U7150 (N_7150,N_4195,N_1635);
nand U7151 (N_7151,N_581,N_957);
and U7152 (N_7152,N_947,N_4009);
or U7153 (N_7153,N_4299,N_2255);
nor U7154 (N_7154,N_112,N_4268);
or U7155 (N_7155,N_4304,N_3796);
or U7156 (N_7156,N_3768,N_527);
nand U7157 (N_7157,N_4321,N_305);
or U7158 (N_7158,N_1425,N_3710);
nand U7159 (N_7159,N_2543,N_976);
or U7160 (N_7160,N_3849,N_553);
or U7161 (N_7161,N_1682,N_151);
nor U7162 (N_7162,N_773,N_2092);
nor U7163 (N_7163,N_1111,N_190);
nor U7164 (N_7164,N_3812,N_1530);
nor U7165 (N_7165,N_578,N_2243);
or U7166 (N_7166,N_4281,N_1882);
and U7167 (N_7167,N_2600,N_2746);
or U7168 (N_7168,N_2149,N_1180);
nand U7169 (N_7169,N_3043,N_3232);
nor U7170 (N_7170,N_3239,N_635);
and U7171 (N_7171,N_4744,N_1283);
and U7172 (N_7172,N_4391,N_2195);
and U7173 (N_7173,N_4689,N_1588);
nand U7174 (N_7174,N_4303,N_1655);
nand U7175 (N_7175,N_2835,N_361);
or U7176 (N_7176,N_4520,N_3392);
and U7177 (N_7177,N_1820,N_2566);
and U7178 (N_7178,N_687,N_4048);
and U7179 (N_7179,N_583,N_2824);
or U7180 (N_7180,N_2465,N_4537);
nor U7181 (N_7181,N_4014,N_2987);
and U7182 (N_7182,N_763,N_1493);
nor U7183 (N_7183,N_4131,N_3111);
or U7184 (N_7184,N_1897,N_3459);
nor U7185 (N_7185,N_3401,N_1490);
nor U7186 (N_7186,N_2794,N_2901);
or U7187 (N_7187,N_1102,N_1341);
nand U7188 (N_7188,N_1348,N_3372);
nand U7189 (N_7189,N_1419,N_3257);
or U7190 (N_7190,N_3277,N_182);
and U7191 (N_7191,N_3371,N_4911);
nand U7192 (N_7192,N_1873,N_4829);
nand U7193 (N_7193,N_2885,N_4594);
or U7194 (N_7194,N_2841,N_4963);
nand U7195 (N_7195,N_939,N_4161);
or U7196 (N_7196,N_2867,N_2650);
nor U7197 (N_7197,N_4390,N_1127);
nand U7198 (N_7198,N_1270,N_3016);
or U7199 (N_7199,N_4761,N_1640);
and U7200 (N_7200,N_1704,N_2760);
and U7201 (N_7201,N_2385,N_2723);
and U7202 (N_7202,N_1138,N_1181);
and U7203 (N_7203,N_4323,N_3150);
or U7204 (N_7204,N_2433,N_4943);
or U7205 (N_7205,N_2734,N_3878);
and U7206 (N_7206,N_1208,N_4571);
and U7207 (N_7207,N_514,N_2180);
nor U7208 (N_7208,N_1297,N_515);
and U7209 (N_7209,N_4443,N_1950);
and U7210 (N_7210,N_4254,N_4820);
nand U7211 (N_7211,N_3364,N_2059);
nor U7212 (N_7212,N_2685,N_192);
nor U7213 (N_7213,N_4274,N_4803);
nand U7214 (N_7214,N_4836,N_825);
nand U7215 (N_7215,N_4021,N_2097);
or U7216 (N_7216,N_3116,N_1368);
nand U7217 (N_7217,N_4352,N_1199);
nor U7218 (N_7218,N_3064,N_2026);
or U7219 (N_7219,N_3816,N_4273);
or U7220 (N_7220,N_3642,N_2331);
and U7221 (N_7221,N_3978,N_3918);
nand U7222 (N_7222,N_4542,N_4050);
or U7223 (N_7223,N_520,N_4414);
nor U7224 (N_7224,N_1629,N_110);
and U7225 (N_7225,N_52,N_4277);
nor U7226 (N_7226,N_3720,N_4225);
xnor U7227 (N_7227,N_1092,N_2042);
and U7228 (N_7228,N_1720,N_1501);
or U7229 (N_7229,N_4394,N_1056);
or U7230 (N_7230,N_2165,N_1414);
and U7231 (N_7231,N_4052,N_142);
and U7232 (N_7232,N_310,N_388);
or U7233 (N_7233,N_4314,N_1849);
nor U7234 (N_7234,N_3211,N_2431);
and U7235 (N_7235,N_78,N_1875);
or U7236 (N_7236,N_778,N_3775);
or U7237 (N_7237,N_364,N_4387);
and U7238 (N_7238,N_2206,N_921);
and U7239 (N_7239,N_2030,N_209);
nand U7240 (N_7240,N_3077,N_3559);
and U7241 (N_7241,N_4755,N_774);
or U7242 (N_7242,N_1646,N_4862);
and U7243 (N_7243,N_214,N_3737);
nand U7244 (N_7244,N_1775,N_231);
nor U7245 (N_7245,N_3437,N_1497);
nand U7246 (N_7246,N_1040,N_3565);
nor U7247 (N_7247,N_733,N_4468);
xnor U7248 (N_7248,N_1518,N_931);
nor U7249 (N_7249,N_4548,N_3635);
nor U7250 (N_7250,N_3973,N_4360);
nand U7251 (N_7251,N_2085,N_2354);
and U7252 (N_7252,N_300,N_2882);
nor U7253 (N_7253,N_1464,N_955);
or U7254 (N_7254,N_628,N_43);
or U7255 (N_7255,N_4814,N_4100);
nor U7256 (N_7256,N_598,N_450);
and U7257 (N_7257,N_738,N_4335);
xnor U7258 (N_7258,N_2349,N_937);
nand U7259 (N_7259,N_2781,N_3029);
nor U7260 (N_7260,N_371,N_4066);
nor U7261 (N_7261,N_4751,N_2648);
or U7262 (N_7262,N_782,N_3797);
or U7263 (N_7263,N_84,N_2571);
and U7264 (N_7264,N_139,N_1474);
and U7265 (N_7265,N_1883,N_2267);
nor U7266 (N_7266,N_3479,N_240);
and U7267 (N_7267,N_2922,N_4449);
nor U7268 (N_7268,N_158,N_1042);
xnor U7269 (N_7269,N_4126,N_4563);
nor U7270 (N_7270,N_2437,N_3611);
and U7271 (N_7271,N_3773,N_2917);
or U7272 (N_7272,N_3028,N_704);
nand U7273 (N_7273,N_2890,N_3195);
nor U7274 (N_7274,N_4746,N_217);
nor U7275 (N_7275,N_4508,N_4132);
and U7276 (N_7276,N_1681,N_4179);
nand U7277 (N_7277,N_295,N_768);
nand U7278 (N_7278,N_33,N_518);
nor U7279 (N_7279,N_724,N_1993);
nand U7280 (N_7280,N_3230,N_4045);
nand U7281 (N_7281,N_791,N_727);
and U7282 (N_7282,N_1455,N_4264);
and U7283 (N_7283,N_2084,N_4446);
or U7284 (N_7284,N_742,N_1971);
or U7285 (N_7285,N_2500,N_4069);
nand U7286 (N_7286,N_649,N_893);
and U7287 (N_7287,N_4938,N_1511);
and U7288 (N_7288,N_907,N_356);
nor U7289 (N_7289,N_3649,N_3026);
nor U7290 (N_7290,N_2205,N_2446);
nand U7291 (N_7291,N_3115,N_895);
nand U7292 (N_7292,N_2355,N_1860);
nor U7293 (N_7293,N_4013,N_2837);
nand U7294 (N_7294,N_2196,N_1310);
and U7295 (N_7295,N_115,N_1264);
nand U7296 (N_7296,N_3919,N_2339);
nor U7297 (N_7297,N_1489,N_1229);
nor U7298 (N_7298,N_162,N_3120);
nor U7299 (N_7299,N_596,N_3569);
nor U7300 (N_7300,N_138,N_4081);
nand U7301 (N_7301,N_2611,N_3591);
and U7302 (N_7302,N_4102,N_1765);
nor U7303 (N_7303,N_2050,N_3145);
or U7304 (N_7304,N_210,N_1836);
or U7305 (N_7305,N_4660,N_2418);
and U7306 (N_7306,N_1320,N_4513);
nand U7307 (N_7307,N_2639,N_3730);
nand U7308 (N_7308,N_3897,N_828);
and U7309 (N_7309,N_3032,N_1876);
and U7310 (N_7310,N_66,N_4695);
xor U7311 (N_7311,N_4082,N_81);
and U7312 (N_7312,N_1675,N_2904);
or U7313 (N_7313,N_729,N_1438);
and U7314 (N_7314,N_2722,N_2670);
nor U7315 (N_7315,N_327,N_2703);
nand U7316 (N_7316,N_827,N_1537);
nand U7317 (N_7317,N_2369,N_918);
nor U7318 (N_7318,N_90,N_1667);
or U7319 (N_7319,N_4130,N_741);
nor U7320 (N_7320,N_902,N_2586);
nand U7321 (N_7321,N_3443,N_1034);
nor U7322 (N_7322,N_888,N_3705);
or U7323 (N_7323,N_1991,N_1279);
nor U7324 (N_7324,N_3615,N_4907);
nand U7325 (N_7325,N_2032,N_2884);
and U7326 (N_7326,N_3318,N_1013);
nand U7327 (N_7327,N_694,N_4922);
nor U7328 (N_7328,N_1254,N_1780);
or U7329 (N_7329,N_3714,N_21);
or U7330 (N_7330,N_2384,N_2938);
nor U7331 (N_7331,N_2366,N_2681);
and U7332 (N_7332,N_2729,N_945);
nand U7333 (N_7333,N_3056,N_3989);
or U7334 (N_7334,N_3406,N_3984);
nand U7335 (N_7335,N_3606,N_2553);
nor U7336 (N_7336,N_3567,N_2676);
and U7337 (N_7337,N_2971,N_3806);
nand U7338 (N_7338,N_3536,N_2057);
nor U7339 (N_7339,N_3429,N_1233);
nand U7340 (N_7340,N_2461,N_3561);
nor U7341 (N_7341,N_4173,N_949);
and U7342 (N_7342,N_2601,N_232);
nand U7343 (N_7343,N_3261,N_3725);
and U7344 (N_7344,N_1654,N_4595);
or U7345 (N_7345,N_1594,N_1559);
or U7346 (N_7346,N_2942,N_4177);
nor U7347 (N_7347,N_1980,N_3748);
xnor U7348 (N_7348,N_3658,N_595);
and U7349 (N_7349,N_3507,N_29);
nand U7350 (N_7350,N_241,N_4200);
nand U7351 (N_7351,N_2449,N_3519);
and U7352 (N_7352,N_4376,N_3590);
or U7353 (N_7353,N_1932,N_1790);
and U7354 (N_7354,N_1287,N_2203);
or U7355 (N_7355,N_1736,N_526);
nand U7356 (N_7356,N_1359,N_3623);
and U7357 (N_7357,N_4798,N_4579);
or U7358 (N_7358,N_4158,N_1158);
nand U7359 (N_7359,N_2362,N_449);
and U7360 (N_7360,N_4812,N_2932);
and U7361 (N_7361,N_3183,N_1012);
and U7362 (N_7362,N_3866,N_399);
nand U7363 (N_7363,N_3788,N_3242);
or U7364 (N_7364,N_4072,N_3759);
and U7365 (N_7365,N_2565,N_1874);
nor U7366 (N_7366,N_1450,N_3926);
and U7367 (N_7367,N_2608,N_4810);
nand U7368 (N_7368,N_152,N_1216);
nand U7369 (N_7369,N_3873,N_1304);
or U7370 (N_7370,N_4993,N_2264);
nand U7371 (N_7371,N_3403,N_4457);
or U7372 (N_7372,N_3023,N_4318);
and U7373 (N_7373,N_4640,N_4322);
nand U7374 (N_7374,N_1344,N_2707);
nand U7375 (N_7375,N_4351,N_4747);
nor U7376 (N_7376,N_1132,N_314);
nand U7377 (N_7377,N_2743,N_901);
nor U7378 (N_7378,N_1946,N_2108);
nand U7379 (N_7379,N_242,N_716);
nand U7380 (N_7380,N_4031,N_801);
and U7381 (N_7381,N_3609,N_2374);
nand U7382 (N_7382,N_1331,N_536);
nor U7383 (N_7383,N_4583,N_2054);
nand U7384 (N_7384,N_2218,N_4259);
or U7385 (N_7385,N_4985,N_705);
nor U7386 (N_7386,N_3184,N_1196);
and U7387 (N_7387,N_4062,N_2358);
or U7388 (N_7388,N_2118,N_2985);
or U7389 (N_7389,N_2844,N_4558);
nand U7390 (N_7390,N_4,N_1561);
nand U7391 (N_7391,N_3727,N_3188);
nor U7392 (N_7392,N_2063,N_1258);
and U7393 (N_7393,N_4208,N_2814);
or U7394 (N_7394,N_2329,N_2928);
nand U7395 (N_7395,N_2138,N_4331);
nand U7396 (N_7396,N_3625,N_1762);
and U7397 (N_7397,N_2847,N_4397);
nor U7398 (N_7398,N_198,N_3070);
and U7399 (N_7399,N_4244,N_4969);
and U7400 (N_7400,N_979,N_1134);
or U7401 (N_7401,N_1757,N_1631);
nor U7402 (N_7402,N_3436,N_3212);
or U7403 (N_7403,N_317,N_4420);
nand U7404 (N_7404,N_1117,N_2028);
or U7405 (N_7405,N_65,N_1250);
nand U7406 (N_7406,N_3315,N_616);
nor U7407 (N_7407,N_524,N_1607);
and U7408 (N_7408,N_3489,N_4587);
nand U7409 (N_7409,N_2226,N_1097);
and U7410 (N_7410,N_239,N_4312);
and U7411 (N_7411,N_3012,N_1371);
xnor U7412 (N_7412,N_1018,N_263);
nand U7413 (N_7413,N_1463,N_4667);
xnor U7414 (N_7414,N_1378,N_4585);
or U7415 (N_7415,N_1688,N_4092);
and U7416 (N_7416,N_4485,N_2657);
nand U7417 (N_7417,N_1308,N_1563);
nor U7418 (N_7418,N_349,N_4140);
and U7419 (N_7419,N_4008,N_3450);
and U7420 (N_7420,N_3924,N_3482);
and U7421 (N_7421,N_1729,N_3011);
nor U7422 (N_7422,N_4639,N_1529);
and U7423 (N_7423,N_1632,N_4189);
or U7424 (N_7424,N_4987,N_4149);
or U7425 (N_7425,N_1205,N_4983);
and U7426 (N_7426,N_1766,N_4037);
and U7427 (N_7427,N_2131,N_389);
or U7428 (N_7428,N_3081,N_3186);
and U7429 (N_7429,N_1301,N_969);
and U7430 (N_7430,N_1039,N_3431);
or U7431 (N_7431,N_1203,N_669);
nor U7432 (N_7432,N_3421,N_4156);
nor U7433 (N_7433,N_3286,N_1641);
nor U7434 (N_7434,N_4118,N_2098);
nand U7435 (N_7435,N_2686,N_3930);
nand U7436 (N_7436,N_1112,N_1597);
nand U7437 (N_7437,N_4709,N_4228);
and U7438 (N_7438,N_4765,N_3440);
or U7439 (N_7439,N_3509,N_4029);
and U7440 (N_7440,N_599,N_3981);
or U7441 (N_7441,N_4831,N_3889);
nor U7442 (N_7442,N_3213,N_4265);
nand U7443 (N_7443,N_3627,N_442);
or U7444 (N_7444,N_1626,N_1271);
nor U7445 (N_7445,N_523,N_3349);
or U7446 (N_7446,N_3855,N_1568);
xnor U7447 (N_7447,N_2720,N_637);
nand U7448 (N_7448,N_212,N_797);
nor U7449 (N_7449,N_1944,N_1386);
nor U7450 (N_7450,N_2679,N_2357);
nor U7451 (N_7451,N_3659,N_8);
or U7452 (N_7452,N_3342,N_453);
or U7453 (N_7453,N_4551,N_405);
and U7454 (N_7454,N_2580,N_2080);
or U7455 (N_7455,N_1885,N_3112);
nand U7456 (N_7456,N_4146,N_4078);
nand U7457 (N_7457,N_3858,N_1121);
nand U7458 (N_7458,N_4270,N_2402);
and U7459 (N_7459,N_1020,N_4521);
or U7460 (N_7460,N_800,N_3578);
nor U7461 (N_7461,N_2399,N_134);
or U7462 (N_7462,N_1448,N_4912);
nor U7463 (N_7463,N_99,N_1285);
and U7464 (N_7464,N_3194,N_3095);
and U7465 (N_7465,N_4615,N_4532);
nand U7466 (N_7466,N_1548,N_2777);
or U7467 (N_7467,N_434,N_470);
nor U7468 (N_7468,N_3664,N_875);
nand U7469 (N_7469,N_2007,N_80);
or U7470 (N_7470,N_1575,N_4892);
or U7471 (N_7471,N_4250,N_1789);
nor U7472 (N_7472,N_1620,N_712);
and U7473 (N_7473,N_4096,N_2163);
nand U7474 (N_7474,N_996,N_2065);
and U7475 (N_7475,N_3651,N_826);
nor U7476 (N_7476,N_952,N_3267);
nor U7477 (N_7477,N_3316,N_3061);
and U7478 (N_7478,N_3713,N_2540);
nor U7479 (N_7479,N_1703,N_4070);
and U7480 (N_7480,N_3605,N_2102);
or U7481 (N_7481,N_2380,N_2983);
and U7482 (N_7482,N_1385,N_4385);
xor U7483 (N_7483,N_4458,N_4135);
nor U7484 (N_7484,N_3147,N_1333);
or U7485 (N_7485,N_17,N_3065);
and U7486 (N_7486,N_3363,N_3202);
nand U7487 (N_7487,N_4995,N_208);
nand U7488 (N_7488,N_1274,N_626);
or U7489 (N_7489,N_3944,N_2174);
xor U7490 (N_7490,N_3948,N_2451);
or U7491 (N_7491,N_474,N_4978);
nor U7492 (N_7492,N_2840,N_395);
and U7493 (N_7493,N_816,N_2862);
nand U7494 (N_7494,N_747,N_2221);
or U7495 (N_7495,N_1120,N_1979);
nor U7496 (N_7496,N_503,N_1418);
nor U7497 (N_7497,N_2207,N_3288);
or U7498 (N_7498,N_4526,N_4666);
nand U7499 (N_7499,N_1987,N_3323);
and U7500 (N_7500,N_302,N_1828);
nor U7501 (N_7501,N_4796,N_2049);
and U7502 (N_7502,N_1308,N_4323);
nand U7503 (N_7503,N_2040,N_3154);
nand U7504 (N_7504,N_2576,N_2907);
or U7505 (N_7505,N_4318,N_1188);
and U7506 (N_7506,N_4554,N_3564);
nor U7507 (N_7507,N_2416,N_347);
and U7508 (N_7508,N_222,N_1073);
and U7509 (N_7509,N_1770,N_1199);
nor U7510 (N_7510,N_1252,N_2813);
nand U7511 (N_7511,N_1667,N_3392);
or U7512 (N_7512,N_4156,N_2263);
nand U7513 (N_7513,N_2168,N_1556);
and U7514 (N_7514,N_941,N_2707);
and U7515 (N_7515,N_2387,N_2776);
xnor U7516 (N_7516,N_1641,N_3016);
and U7517 (N_7517,N_2536,N_2205);
nand U7518 (N_7518,N_399,N_39);
nand U7519 (N_7519,N_3060,N_411);
or U7520 (N_7520,N_4399,N_828);
nor U7521 (N_7521,N_1866,N_1865);
nand U7522 (N_7522,N_2473,N_1116);
or U7523 (N_7523,N_1581,N_213);
xnor U7524 (N_7524,N_2299,N_2193);
and U7525 (N_7525,N_2691,N_4283);
or U7526 (N_7526,N_2454,N_2787);
nor U7527 (N_7527,N_4662,N_332);
and U7528 (N_7528,N_4971,N_1743);
and U7529 (N_7529,N_119,N_4877);
or U7530 (N_7530,N_1217,N_4284);
and U7531 (N_7531,N_3375,N_3657);
or U7532 (N_7532,N_90,N_4091);
and U7533 (N_7533,N_3815,N_4448);
nand U7534 (N_7534,N_1541,N_2829);
and U7535 (N_7535,N_2428,N_1463);
nand U7536 (N_7536,N_4475,N_773);
nor U7537 (N_7537,N_1169,N_4455);
and U7538 (N_7538,N_3911,N_4632);
nor U7539 (N_7539,N_2588,N_4660);
and U7540 (N_7540,N_3088,N_710);
nand U7541 (N_7541,N_360,N_2257);
nand U7542 (N_7542,N_2435,N_3862);
and U7543 (N_7543,N_2938,N_580);
or U7544 (N_7544,N_3808,N_4741);
and U7545 (N_7545,N_981,N_3503);
nor U7546 (N_7546,N_3554,N_3226);
nor U7547 (N_7547,N_778,N_2217);
and U7548 (N_7548,N_1193,N_3566);
or U7549 (N_7549,N_1196,N_1325);
nand U7550 (N_7550,N_4410,N_1023);
or U7551 (N_7551,N_2633,N_2663);
and U7552 (N_7552,N_1894,N_4395);
or U7553 (N_7553,N_807,N_1589);
or U7554 (N_7554,N_618,N_690);
and U7555 (N_7555,N_2453,N_464);
nand U7556 (N_7556,N_39,N_2195);
or U7557 (N_7557,N_2115,N_4970);
and U7558 (N_7558,N_2493,N_483);
xnor U7559 (N_7559,N_2988,N_490);
nor U7560 (N_7560,N_4759,N_270);
or U7561 (N_7561,N_1258,N_3002);
nor U7562 (N_7562,N_305,N_469);
and U7563 (N_7563,N_2380,N_1041);
nand U7564 (N_7564,N_259,N_2284);
nor U7565 (N_7565,N_2874,N_3019);
and U7566 (N_7566,N_3819,N_714);
nand U7567 (N_7567,N_3191,N_2296);
nor U7568 (N_7568,N_4140,N_208);
and U7569 (N_7569,N_1989,N_1828);
and U7570 (N_7570,N_4180,N_3625);
or U7571 (N_7571,N_3625,N_4937);
nor U7572 (N_7572,N_1581,N_2200);
nand U7573 (N_7573,N_2948,N_1129);
nor U7574 (N_7574,N_3710,N_775);
or U7575 (N_7575,N_1854,N_3972);
nand U7576 (N_7576,N_1662,N_1784);
nand U7577 (N_7577,N_4703,N_1261);
nor U7578 (N_7578,N_4711,N_3282);
or U7579 (N_7579,N_4403,N_497);
and U7580 (N_7580,N_4567,N_2405);
nor U7581 (N_7581,N_305,N_1119);
and U7582 (N_7582,N_318,N_911);
and U7583 (N_7583,N_2864,N_2785);
nor U7584 (N_7584,N_1610,N_3441);
nor U7585 (N_7585,N_2638,N_3935);
and U7586 (N_7586,N_1461,N_898);
nor U7587 (N_7587,N_3257,N_2630);
and U7588 (N_7588,N_1192,N_143);
and U7589 (N_7589,N_4873,N_555);
or U7590 (N_7590,N_1266,N_3327);
nor U7591 (N_7591,N_2140,N_2594);
nor U7592 (N_7592,N_2062,N_828);
nor U7593 (N_7593,N_312,N_1741);
and U7594 (N_7594,N_1928,N_138);
nor U7595 (N_7595,N_2288,N_4729);
nand U7596 (N_7596,N_4741,N_1304);
nor U7597 (N_7597,N_969,N_831);
or U7598 (N_7598,N_4714,N_2449);
or U7599 (N_7599,N_266,N_4615);
xor U7600 (N_7600,N_1288,N_890);
xnor U7601 (N_7601,N_357,N_4933);
and U7602 (N_7602,N_1795,N_4428);
nor U7603 (N_7603,N_4742,N_4270);
and U7604 (N_7604,N_1214,N_758);
or U7605 (N_7605,N_1718,N_4635);
and U7606 (N_7606,N_1091,N_1431);
or U7607 (N_7607,N_3788,N_2930);
or U7608 (N_7608,N_3778,N_2604);
xor U7609 (N_7609,N_3251,N_2004);
or U7610 (N_7610,N_4407,N_2487);
nor U7611 (N_7611,N_785,N_3867);
nand U7612 (N_7612,N_200,N_1912);
nor U7613 (N_7613,N_3822,N_2479);
nor U7614 (N_7614,N_3939,N_4811);
nand U7615 (N_7615,N_1177,N_3214);
nand U7616 (N_7616,N_4845,N_3684);
nor U7617 (N_7617,N_1045,N_2343);
nand U7618 (N_7618,N_3422,N_3458);
or U7619 (N_7619,N_2550,N_31);
or U7620 (N_7620,N_4712,N_909);
or U7621 (N_7621,N_3599,N_989);
nand U7622 (N_7622,N_4199,N_4892);
nand U7623 (N_7623,N_4478,N_1064);
nor U7624 (N_7624,N_4571,N_4715);
nor U7625 (N_7625,N_1908,N_573);
nand U7626 (N_7626,N_176,N_3774);
and U7627 (N_7627,N_4093,N_3087);
nor U7628 (N_7628,N_2618,N_3598);
nor U7629 (N_7629,N_70,N_1154);
or U7630 (N_7630,N_2999,N_895);
nand U7631 (N_7631,N_3075,N_4963);
nor U7632 (N_7632,N_1789,N_3727);
or U7633 (N_7633,N_2932,N_1633);
or U7634 (N_7634,N_887,N_2986);
nor U7635 (N_7635,N_3511,N_510);
and U7636 (N_7636,N_1340,N_1115);
nor U7637 (N_7637,N_2836,N_943);
xnor U7638 (N_7638,N_198,N_362);
nor U7639 (N_7639,N_2022,N_1446);
nand U7640 (N_7640,N_2036,N_1294);
xor U7641 (N_7641,N_303,N_897);
nand U7642 (N_7642,N_848,N_4264);
and U7643 (N_7643,N_992,N_4940);
or U7644 (N_7644,N_3158,N_3201);
nand U7645 (N_7645,N_4433,N_604);
nand U7646 (N_7646,N_1423,N_3026);
nand U7647 (N_7647,N_1670,N_3003);
or U7648 (N_7648,N_3718,N_1343);
nor U7649 (N_7649,N_4318,N_2671);
nand U7650 (N_7650,N_3779,N_1505);
nand U7651 (N_7651,N_507,N_1740);
nor U7652 (N_7652,N_3116,N_1073);
nor U7653 (N_7653,N_343,N_2709);
nor U7654 (N_7654,N_4130,N_3171);
or U7655 (N_7655,N_2208,N_452);
nand U7656 (N_7656,N_1202,N_2819);
or U7657 (N_7657,N_4018,N_890);
and U7658 (N_7658,N_3349,N_3123);
nand U7659 (N_7659,N_935,N_2531);
or U7660 (N_7660,N_2376,N_4388);
nor U7661 (N_7661,N_1069,N_3025);
and U7662 (N_7662,N_4410,N_3935);
nand U7663 (N_7663,N_1495,N_2711);
or U7664 (N_7664,N_4114,N_2584);
nand U7665 (N_7665,N_1520,N_2828);
nor U7666 (N_7666,N_1674,N_3730);
nand U7667 (N_7667,N_2680,N_2464);
nand U7668 (N_7668,N_4514,N_3534);
nand U7669 (N_7669,N_3241,N_638);
or U7670 (N_7670,N_4889,N_601);
and U7671 (N_7671,N_1821,N_2499);
or U7672 (N_7672,N_1933,N_3264);
or U7673 (N_7673,N_859,N_2992);
or U7674 (N_7674,N_1107,N_984);
or U7675 (N_7675,N_207,N_3605);
nor U7676 (N_7676,N_4214,N_4254);
and U7677 (N_7677,N_2181,N_412);
xnor U7678 (N_7678,N_2512,N_948);
nor U7679 (N_7679,N_2785,N_2601);
and U7680 (N_7680,N_4774,N_4068);
xor U7681 (N_7681,N_4147,N_4290);
and U7682 (N_7682,N_4212,N_3786);
nand U7683 (N_7683,N_4815,N_3495);
and U7684 (N_7684,N_3600,N_311);
or U7685 (N_7685,N_4809,N_3661);
nor U7686 (N_7686,N_4133,N_4428);
or U7687 (N_7687,N_1228,N_2164);
and U7688 (N_7688,N_3928,N_3754);
or U7689 (N_7689,N_1694,N_2288);
or U7690 (N_7690,N_1344,N_1103);
and U7691 (N_7691,N_1414,N_199);
and U7692 (N_7692,N_805,N_2012);
and U7693 (N_7693,N_1775,N_3827);
nor U7694 (N_7694,N_1499,N_1268);
and U7695 (N_7695,N_665,N_2927);
nand U7696 (N_7696,N_1729,N_4071);
or U7697 (N_7697,N_3086,N_626);
nand U7698 (N_7698,N_1303,N_4902);
or U7699 (N_7699,N_1892,N_927);
nand U7700 (N_7700,N_2157,N_2345);
nor U7701 (N_7701,N_1798,N_4208);
nand U7702 (N_7702,N_2984,N_3780);
and U7703 (N_7703,N_4786,N_4061);
nor U7704 (N_7704,N_547,N_4676);
nand U7705 (N_7705,N_2255,N_1273);
nand U7706 (N_7706,N_1908,N_2044);
or U7707 (N_7707,N_1742,N_3991);
and U7708 (N_7708,N_4392,N_2490);
nor U7709 (N_7709,N_3773,N_1156);
or U7710 (N_7710,N_3080,N_411);
nor U7711 (N_7711,N_118,N_1056);
and U7712 (N_7712,N_2137,N_1867);
nor U7713 (N_7713,N_2448,N_2366);
or U7714 (N_7714,N_2361,N_839);
or U7715 (N_7715,N_641,N_3312);
or U7716 (N_7716,N_4383,N_3127);
or U7717 (N_7717,N_2539,N_4026);
nor U7718 (N_7718,N_2452,N_4619);
nand U7719 (N_7719,N_431,N_4116);
or U7720 (N_7720,N_2067,N_4468);
nand U7721 (N_7721,N_4038,N_4341);
or U7722 (N_7722,N_3253,N_4320);
or U7723 (N_7723,N_3104,N_3054);
and U7724 (N_7724,N_4231,N_3989);
and U7725 (N_7725,N_1353,N_4880);
and U7726 (N_7726,N_2059,N_4476);
nor U7727 (N_7727,N_4261,N_2794);
nor U7728 (N_7728,N_1928,N_1812);
nor U7729 (N_7729,N_4503,N_655);
or U7730 (N_7730,N_1262,N_3470);
and U7731 (N_7731,N_192,N_4943);
xnor U7732 (N_7732,N_933,N_1678);
nand U7733 (N_7733,N_447,N_3396);
nor U7734 (N_7734,N_4916,N_3212);
and U7735 (N_7735,N_4050,N_853);
and U7736 (N_7736,N_919,N_1853);
and U7737 (N_7737,N_2714,N_271);
or U7738 (N_7738,N_72,N_813);
nor U7739 (N_7739,N_1004,N_4195);
nor U7740 (N_7740,N_573,N_3605);
nand U7741 (N_7741,N_3591,N_2621);
and U7742 (N_7742,N_192,N_650);
nor U7743 (N_7743,N_3853,N_3771);
nand U7744 (N_7744,N_3583,N_2998);
and U7745 (N_7745,N_410,N_4873);
nor U7746 (N_7746,N_1437,N_1404);
nor U7747 (N_7747,N_4032,N_2522);
or U7748 (N_7748,N_4278,N_824);
and U7749 (N_7749,N_722,N_678);
and U7750 (N_7750,N_1536,N_3351);
nand U7751 (N_7751,N_278,N_3863);
and U7752 (N_7752,N_2706,N_26);
nand U7753 (N_7753,N_4835,N_1892);
nand U7754 (N_7754,N_3160,N_3356);
or U7755 (N_7755,N_2996,N_2980);
or U7756 (N_7756,N_3326,N_4039);
nand U7757 (N_7757,N_31,N_2265);
or U7758 (N_7758,N_3390,N_1170);
and U7759 (N_7759,N_4985,N_2142);
or U7760 (N_7760,N_1085,N_983);
or U7761 (N_7761,N_1407,N_1065);
nand U7762 (N_7762,N_3021,N_702);
nand U7763 (N_7763,N_370,N_3469);
nor U7764 (N_7764,N_429,N_4030);
or U7765 (N_7765,N_47,N_1056);
and U7766 (N_7766,N_63,N_2531);
nor U7767 (N_7767,N_736,N_2894);
nand U7768 (N_7768,N_3755,N_2489);
xnor U7769 (N_7769,N_2011,N_4667);
or U7770 (N_7770,N_2835,N_2247);
nor U7771 (N_7771,N_3907,N_1358);
nand U7772 (N_7772,N_4982,N_3409);
nand U7773 (N_7773,N_1375,N_3049);
nor U7774 (N_7774,N_3667,N_1518);
nor U7775 (N_7775,N_4855,N_3531);
and U7776 (N_7776,N_618,N_3550);
nand U7777 (N_7777,N_1173,N_3342);
and U7778 (N_7778,N_4240,N_4716);
and U7779 (N_7779,N_2347,N_4393);
and U7780 (N_7780,N_3009,N_180);
nor U7781 (N_7781,N_4872,N_4503);
nor U7782 (N_7782,N_44,N_1919);
nand U7783 (N_7783,N_992,N_3525);
and U7784 (N_7784,N_366,N_2983);
and U7785 (N_7785,N_4074,N_569);
or U7786 (N_7786,N_1015,N_4015);
nand U7787 (N_7787,N_907,N_2413);
and U7788 (N_7788,N_2805,N_2346);
and U7789 (N_7789,N_1362,N_3096);
nor U7790 (N_7790,N_4579,N_4511);
nor U7791 (N_7791,N_2746,N_1165);
nand U7792 (N_7792,N_2587,N_2600);
nand U7793 (N_7793,N_3105,N_2531);
and U7794 (N_7794,N_2483,N_1614);
xor U7795 (N_7795,N_2103,N_1562);
and U7796 (N_7796,N_491,N_3731);
or U7797 (N_7797,N_1816,N_4751);
nor U7798 (N_7798,N_4802,N_3855);
nand U7799 (N_7799,N_1538,N_4785);
and U7800 (N_7800,N_3208,N_3932);
nor U7801 (N_7801,N_297,N_1497);
or U7802 (N_7802,N_641,N_1009);
nor U7803 (N_7803,N_3938,N_565);
and U7804 (N_7804,N_4542,N_393);
nor U7805 (N_7805,N_1235,N_4259);
nor U7806 (N_7806,N_2784,N_581);
nand U7807 (N_7807,N_3046,N_2122);
xor U7808 (N_7808,N_2286,N_1722);
nand U7809 (N_7809,N_2189,N_4889);
and U7810 (N_7810,N_3829,N_2211);
nor U7811 (N_7811,N_4488,N_3815);
nand U7812 (N_7812,N_1703,N_803);
nor U7813 (N_7813,N_4936,N_4542);
nor U7814 (N_7814,N_2180,N_1536);
nor U7815 (N_7815,N_4374,N_2576);
or U7816 (N_7816,N_4525,N_3949);
nor U7817 (N_7817,N_1242,N_595);
nand U7818 (N_7818,N_4024,N_721);
or U7819 (N_7819,N_2940,N_3216);
or U7820 (N_7820,N_1468,N_1730);
and U7821 (N_7821,N_3929,N_3114);
and U7822 (N_7822,N_484,N_1347);
and U7823 (N_7823,N_3000,N_938);
or U7824 (N_7824,N_4052,N_439);
or U7825 (N_7825,N_3713,N_544);
or U7826 (N_7826,N_3976,N_1700);
nor U7827 (N_7827,N_517,N_4176);
or U7828 (N_7828,N_2963,N_4838);
nand U7829 (N_7829,N_4348,N_2317);
xnor U7830 (N_7830,N_3360,N_4174);
nand U7831 (N_7831,N_4755,N_786);
or U7832 (N_7832,N_4040,N_3628);
nor U7833 (N_7833,N_1142,N_3337);
nor U7834 (N_7834,N_1916,N_2902);
nor U7835 (N_7835,N_400,N_1362);
and U7836 (N_7836,N_1092,N_2088);
or U7837 (N_7837,N_4469,N_2403);
and U7838 (N_7838,N_4853,N_2938);
nor U7839 (N_7839,N_3173,N_2049);
and U7840 (N_7840,N_4150,N_1507);
nand U7841 (N_7841,N_2559,N_2260);
and U7842 (N_7842,N_805,N_4449);
nor U7843 (N_7843,N_888,N_4108);
nand U7844 (N_7844,N_2318,N_1865);
or U7845 (N_7845,N_4949,N_4897);
or U7846 (N_7846,N_4674,N_4161);
and U7847 (N_7847,N_2340,N_225);
and U7848 (N_7848,N_1457,N_2553);
and U7849 (N_7849,N_3819,N_4527);
nor U7850 (N_7850,N_1953,N_2559);
nor U7851 (N_7851,N_3947,N_1802);
nor U7852 (N_7852,N_3567,N_2138);
or U7853 (N_7853,N_4551,N_4368);
nand U7854 (N_7854,N_4310,N_1395);
or U7855 (N_7855,N_3991,N_2915);
and U7856 (N_7856,N_427,N_1127);
nand U7857 (N_7857,N_3297,N_548);
and U7858 (N_7858,N_4465,N_2289);
and U7859 (N_7859,N_2593,N_2093);
nand U7860 (N_7860,N_3640,N_1608);
nand U7861 (N_7861,N_2222,N_4323);
nand U7862 (N_7862,N_389,N_789);
and U7863 (N_7863,N_2666,N_1358);
xnor U7864 (N_7864,N_2333,N_983);
and U7865 (N_7865,N_4785,N_3857);
xor U7866 (N_7866,N_1670,N_2285);
and U7867 (N_7867,N_277,N_4763);
or U7868 (N_7868,N_91,N_1041);
nor U7869 (N_7869,N_981,N_295);
and U7870 (N_7870,N_4141,N_1925);
and U7871 (N_7871,N_2159,N_3033);
or U7872 (N_7872,N_2564,N_811);
and U7873 (N_7873,N_4395,N_3488);
xnor U7874 (N_7874,N_4772,N_1893);
nand U7875 (N_7875,N_3395,N_1106);
or U7876 (N_7876,N_3666,N_3905);
nor U7877 (N_7877,N_577,N_4597);
nor U7878 (N_7878,N_4929,N_350);
nand U7879 (N_7879,N_4717,N_4862);
or U7880 (N_7880,N_1625,N_2799);
nand U7881 (N_7881,N_1307,N_945);
nor U7882 (N_7882,N_2252,N_4594);
nor U7883 (N_7883,N_1731,N_4446);
or U7884 (N_7884,N_1728,N_3484);
nor U7885 (N_7885,N_1043,N_3337);
nor U7886 (N_7886,N_548,N_737);
nor U7887 (N_7887,N_2233,N_951);
nor U7888 (N_7888,N_3936,N_183);
or U7889 (N_7889,N_81,N_4477);
and U7890 (N_7890,N_2361,N_4530);
and U7891 (N_7891,N_4137,N_4871);
and U7892 (N_7892,N_4355,N_688);
or U7893 (N_7893,N_3210,N_1699);
or U7894 (N_7894,N_959,N_3548);
or U7895 (N_7895,N_159,N_4782);
nor U7896 (N_7896,N_2359,N_3394);
nor U7897 (N_7897,N_3922,N_316);
or U7898 (N_7898,N_1494,N_3820);
or U7899 (N_7899,N_4258,N_880);
nand U7900 (N_7900,N_972,N_4396);
nand U7901 (N_7901,N_2273,N_4135);
and U7902 (N_7902,N_1358,N_794);
or U7903 (N_7903,N_550,N_4129);
or U7904 (N_7904,N_330,N_2095);
or U7905 (N_7905,N_3266,N_3648);
nand U7906 (N_7906,N_1592,N_997);
and U7907 (N_7907,N_2584,N_871);
and U7908 (N_7908,N_2268,N_518);
nand U7909 (N_7909,N_3573,N_2045);
nand U7910 (N_7910,N_4598,N_2607);
and U7911 (N_7911,N_1366,N_3526);
and U7912 (N_7912,N_1710,N_1684);
or U7913 (N_7913,N_3047,N_2989);
or U7914 (N_7914,N_3559,N_3890);
nand U7915 (N_7915,N_2046,N_4488);
or U7916 (N_7916,N_39,N_481);
nor U7917 (N_7917,N_4891,N_4033);
xnor U7918 (N_7918,N_556,N_3382);
and U7919 (N_7919,N_2809,N_3479);
or U7920 (N_7920,N_4282,N_2656);
or U7921 (N_7921,N_4350,N_1755);
or U7922 (N_7922,N_121,N_3779);
and U7923 (N_7923,N_3707,N_1806);
nor U7924 (N_7924,N_4609,N_2890);
nand U7925 (N_7925,N_3198,N_380);
or U7926 (N_7926,N_4655,N_4652);
nor U7927 (N_7927,N_968,N_1196);
nand U7928 (N_7928,N_3046,N_3037);
and U7929 (N_7929,N_1111,N_3447);
and U7930 (N_7930,N_3383,N_2590);
nor U7931 (N_7931,N_4864,N_4634);
or U7932 (N_7932,N_2555,N_2227);
and U7933 (N_7933,N_3235,N_4876);
nor U7934 (N_7934,N_567,N_1786);
and U7935 (N_7935,N_1723,N_1008);
nand U7936 (N_7936,N_167,N_3442);
or U7937 (N_7937,N_1006,N_4970);
or U7938 (N_7938,N_4687,N_402);
nand U7939 (N_7939,N_3647,N_3095);
or U7940 (N_7940,N_659,N_3707);
nor U7941 (N_7941,N_4781,N_3313);
nand U7942 (N_7942,N_4311,N_1063);
and U7943 (N_7943,N_2936,N_3848);
nor U7944 (N_7944,N_931,N_2531);
nand U7945 (N_7945,N_2507,N_2965);
or U7946 (N_7946,N_4813,N_467);
xor U7947 (N_7947,N_3640,N_2572);
or U7948 (N_7948,N_3169,N_4430);
and U7949 (N_7949,N_4420,N_3091);
nor U7950 (N_7950,N_321,N_959);
nor U7951 (N_7951,N_2308,N_725);
and U7952 (N_7952,N_2766,N_4173);
and U7953 (N_7953,N_3830,N_800);
or U7954 (N_7954,N_136,N_2084);
nand U7955 (N_7955,N_259,N_1040);
or U7956 (N_7956,N_1829,N_4796);
nor U7957 (N_7957,N_3793,N_3795);
nor U7958 (N_7958,N_1268,N_1731);
nand U7959 (N_7959,N_804,N_351);
and U7960 (N_7960,N_2474,N_3275);
nor U7961 (N_7961,N_4423,N_1017);
nor U7962 (N_7962,N_4828,N_3054);
xnor U7963 (N_7963,N_381,N_3631);
or U7964 (N_7964,N_1506,N_1028);
nand U7965 (N_7965,N_776,N_4089);
nand U7966 (N_7966,N_3350,N_1069);
nor U7967 (N_7967,N_3566,N_2965);
and U7968 (N_7968,N_4892,N_992);
and U7969 (N_7969,N_4905,N_2587);
and U7970 (N_7970,N_3031,N_1386);
and U7971 (N_7971,N_4131,N_1904);
nand U7972 (N_7972,N_1650,N_441);
and U7973 (N_7973,N_2220,N_2588);
or U7974 (N_7974,N_4876,N_428);
or U7975 (N_7975,N_4512,N_1911);
nand U7976 (N_7976,N_1553,N_1172);
nand U7977 (N_7977,N_184,N_1684);
and U7978 (N_7978,N_4436,N_1597);
or U7979 (N_7979,N_1742,N_377);
and U7980 (N_7980,N_788,N_3790);
and U7981 (N_7981,N_2977,N_892);
nor U7982 (N_7982,N_4140,N_2270);
and U7983 (N_7983,N_196,N_914);
or U7984 (N_7984,N_1869,N_874);
or U7985 (N_7985,N_3098,N_1040);
and U7986 (N_7986,N_1740,N_3457);
or U7987 (N_7987,N_4207,N_1821);
nand U7988 (N_7988,N_4449,N_203);
and U7989 (N_7989,N_3938,N_3230);
nand U7990 (N_7990,N_2097,N_4012);
nand U7991 (N_7991,N_4656,N_1207);
and U7992 (N_7992,N_152,N_3925);
and U7993 (N_7993,N_454,N_2151);
nor U7994 (N_7994,N_621,N_3954);
or U7995 (N_7995,N_3296,N_2336);
and U7996 (N_7996,N_2624,N_2389);
nand U7997 (N_7997,N_2053,N_220);
nor U7998 (N_7998,N_3847,N_1893);
nand U7999 (N_7999,N_3493,N_4512);
and U8000 (N_8000,N_2077,N_1516);
nand U8001 (N_8001,N_3119,N_4537);
or U8002 (N_8002,N_4817,N_4719);
nor U8003 (N_8003,N_1890,N_1684);
nor U8004 (N_8004,N_3143,N_1324);
or U8005 (N_8005,N_1548,N_3204);
nor U8006 (N_8006,N_4364,N_1315);
nor U8007 (N_8007,N_1396,N_4792);
nand U8008 (N_8008,N_2164,N_4709);
or U8009 (N_8009,N_3449,N_4629);
nand U8010 (N_8010,N_2261,N_55);
nand U8011 (N_8011,N_3814,N_1953);
or U8012 (N_8012,N_4518,N_1819);
or U8013 (N_8013,N_4216,N_2536);
nor U8014 (N_8014,N_3951,N_3844);
nand U8015 (N_8015,N_2747,N_3349);
nand U8016 (N_8016,N_1031,N_570);
or U8017 (N_8017,N_1417,N_2511);
or U8018 (N_8018,N_2646,N_776);
nor U8019 (N_8019,N_1292,N_1019);
nand U8020 (N_8020,N_1159,N_4055);
and U8021 (N_8021,N_3487,N_4269);
and U8022 (N_8022,N_4140,N_4444);
nand U8023 (N_8023,N_2829,N_4696);
nor U8024 (N_8024,N_1459,N_2663);
nor U8025 (N_8025,N_3561,N_2544);
and U8026 (N_8026,N_1178,N_2500);
nor U8027 (N_8027,N_1179,N_3058);
nor U8028 (N_8028,N_1830,N_980);
and U8029 (N_8029,N_4481,N_3594);
or U8030 (N_8030,N_2768,N_791);
xnor U8031 (N_8031,N_2490,N_4500);
nor U8032 (N_8032,N_4136,N_2752);
or U8033 (N_8033,N_4557,N_3046);
nand U8034 (N_8034,N_2976,N_2126);
or U8035 (N_8035,N_2110,N_2621);
and U8036 (N_8036,N_3952,N_1202);
nor U8037 (N_8037,N_1846,N_4404);
or U8038 (N_8038,N_3740,N_2195);
nand U8039 (N_8039,N_3578,N_469);
nor U8040 (N_8040,N_4684,N_261);
or U8041 (N_8041,N_2331,N_4424);
and U8042 (N_8042,N_216,N_3313);
nor U8043 (N_8043,N_3955,N_2467);
nand U8044 (N_8044,N_4412,N_1744);
nand U8045 (N_8045,N_1754,N_519);
and U8046 (N_8046,N_3433,N_4034);
xor U8047 (N_8047,N_291,N_228);
nor U8048 (N_8048,N_3654,N_4956);
and U8049 (N_8049,N_560,N_260);
or U8050 (N_8050,N_2143,N_925);
and U8051 (N_8051,N_2254,N_2632);
or U8052 (N_8052,N_1783,N_3651);
nand U8053 (N_8053,N_2873,N_3562);
or U8054 (N_8054,N_1252,N_2983);
or U8055 (N_8055,N_33,N_4941);
nor U8056 (N_8056,N_3337,N_3074);
nor U8057 (N_8057,N_3020,N_458);
nor U8058 (N_8058,N_2053,N_548);
xnor U8059 (N_8059,N_2502,N_4024);
or U8060 (N_8060,N_1503,N_4111);
or U8061 (N_8061,N_4466,N_1291);
and U8062 (N_8062,N_1341,N_1406);
nor U8063 (N_8063,N_4423,N_993);
or U8064 (N_8064,N_4577,N_2198);
or U8065 (N_8065,N_2850,N_1346);
nor U8066 (N_8066,N_1505,N_326);
nand U8067 (N_8067,N_1985,N_3770);
or U8068 (N_8068,N_2587,N_3819);
xnor U8069 (N_8069,N_4546,N_3896);
nand U8070 (N_8070,N_2499,N_2677);
or U8071 (N_8071,N_2598,N_3984);
and U8072 (N_8072,N_1854,N_1746);
or U8073 (N_8073,N_1862,N_230);
nand U8074 (N_8074,N_4635,N_2924);
and U8075 (N_8075,N_3816,N_1198);
nor U8076 (N_8076,N_1695,N_2450);
nand U8077 (N_8077,N_508,N_2044);
xor U8078 (N_8078,N_395,N_4242);
nand U8079 (N_8079,N_2596,N_1710);
nor U8080 (N_8080,N_4787,N_3216);
nand U8081 (N_8081,N_4610,N_2530);
nor U8082 (N_8082,N_4397,N_1017);
nand U8083 (N_8083,N_4087,N_3120);
nor U8084 (N_8084,N_4323,N_3680);
nor U8085 (N_8085,N_4261,N_1307);
nor U8086 (N_8086,N_1925,N_306);
and U8087 (N_8087,N_67,N_2584);
nand U8088 (N_8088,N_3909,N_3684);
nand U8089 (N_8089,N_1360,N_808);
and U8090 (N_8090,N_4562,N_3774);
xor U8091 (N_8091,N_3762,N_3429);
or U8092 (N_8092,N_1850,N_564);
or U8093 (N_8093,N_1825,N_4760);
nor U8094 (N_8094,N_2575,N_2717);
or U8095 (N_8095,N_2301,N_3931);
or U8096 (N_8096,N_581,N_3491);
or U8097 (N_8097,N_1754,N_1856);
nor U8098 (N_8098,N_780,N_4104);
nor U8099 (N_8099,N_3609,N_1217);
nor U8100 (N_8100,N_122,N_4636);
nand U8101 (N_8101,N_2943,N_2264);
or U8102 (N_8102,N_2685,N_4365);
or U8103 (N_8103,N_1926,N_4296);
nand U8104 (N_8104,N_1050,N_4891);
nand U8105 (N_8105,N_3770,N_3991);
or U8106 (N_8106,N_4799,N_2078);
xnor U8107 (N_8107,N_2069,N_2706);
nand U8108 (N_8108,N_4826,N_3017);
nor U8109 (N_8109,N_4270,N_4860);
nand U8110 (N_8110,N_1399,N_837);
or U8111 (N_8111,N_1069,N_4114);
nand U8112 (N_8112,N_2953,N_447);
nor U8113 (N_8113,N_974,N_271);
or U8114 (N_8114,N_870,N_3385);
or U8115 (N_8115,N_3769,N_2143);
nor U8116 (N_8116,N_2641,N_43);
or U8117 (N_8117,N_312,N_4739);
nand U8118 (N_8118,N_3149,N_3921);
nand U8119 (N_8119,N_3515,N_4873);
nand U8120 (N_8120,N_1930,N_1431);
nor U8121 (N_8121,N_3470,N_180);
nor U8122 (N_8122,N_1319,N_2748);
or U8123 (N_8123,N_3129,N_3316);
and U8124 (N_8124,N_381,N_663);
and U8125 (N_8125,N_507,N_427);
and U8126 (N_8126,N_951,N_4825);
nand U8127 (N_8127,N_3523,N_1080);
or U8128 (N_8128,N_1140,N_614);
nand U8129 (N_8129,N_662,N_1412);
or U8130 (N_8130,N_2059,N_4983);
xnor U8131 (N_8131,N_3383,N_3348);
nor U8132 (N_8132,N_3074,N_4407);
nor U8133 (N_8133,N_4627,N_2421);
nor U8134 (N_8134,N_2776,N_2651);
nor U8135 (N_8135,N_2976,N_2452);
nand U8136 (N_8136,N_3578,N_4599);
nand U8137 (N_8137,N_3798,N_1023);
nor U8138 (N_8138,N_4089,N_3047);
nand U8139 (N_8139,N_383,N_3447);
and U8140 (N_8140,N_658,N_2667);
nand U8141 (N_8141,N_1359,N_2543);
nor U8142 (N_8142,N_2831,N_4084);
nor U8143 (N_8143,N_718,N_3739);
and U8144 (N_8144,N_4126,N_3737);
nand U8145 (N_8145,N_3469,N_2516);
and U8146 (N_8146,N_3491,N_4001);
nor U8147 (N_8147,N_4117,N_1882);
or U8148 (N_8148,N_1633,N_1012);
or U8149 (N_8149,N_3317,N_94);
nor U8150 (N_8150,N_1314,N_2573);
or U8151 (N_8151,N_179,N_1918);
or U8152 (N_8152,N_1485,N_2874);
or U8153 (N_8153,N_2198,N_2877);
and U8154 (N_8154,N_692,N_4056);
and U8155 (N_8155,N_1099,N_1363);
and U8156 (N_8156,N_3716,N_189);
or U8157 (N_8157,N_847,N_3534);
nor U8158 (N_8158,N_2190,N_4071);
nor U8159 (N_8159,N_1735,N_864);
or U8160 (N_8160,N_3422,N_825);
nand U8161 (N_8161,N_433,N_3013);
or U8162 (N_8162,N_2509,N_315);
nand U8163 (N_8163,N_83,N_4038);
nand U8164 (N_8164,N_1100,N_4196);
nand U8165 (N_8165,N_669,N_2890);
and U8166 (N_8166,N_2859,N_3586);
and U8167 (N_8167,N_3327,N_3709);
nand U8168 (N_8168,N_4636,N_1117);
nand U8169 (N_8169,N_4651,N_152);
nor U8170 (N_8170,N_4148,N_1625);
nand U8171 (N_8171,N_2596,N_3358);
nor U8172 (N_8172,N_3830,N_4655);
nor U8173 (N_8173,N_4521,N_1031);
nor U8174 (N_8174,N_1652,N_3159);
or U8175 (N_8175,N_1240,N_4268);
or U8176 (N_8176,N_1867,N_4177);
or U8177 (N_8177,N_4602,N_4773);
nand U8178 (N_8178,N_4539,N_3367);
nand U8179 (N_8179,N_2252,N_553);
and U8180 (N_8180,N_2369,N_1917);
nor U8181 (N_8181,N_1602,N_1931);
or U8182 (N_8182,N_170,N_3058);
or U8183 (N_8183,N_4307,N_4356);
or U8184 (N_8184,N_3021,N_363);
nor U8185 (N_8185,N_4672,N_1827);
nor U8186 (N_8186,N_1488,N_3110);
nand U8187 (N_8187,N_4170,N_1705);
and U8188 (N_8188,N_4427,N_1320);
nand U8189 (N_8189,N_2657,N_2708);
or U8190 (N_8190,N_902,N_1004);
and U8191 (N_8191,N_4898,N_2893);
nand U8192 (N_8192,N_1013,N_1502);
nor U8193 (N_8193,N_942,N_97);
and U8194 (N_8194,N_3903,N_4369);
and U8195 (N_8195,N_3087,N_1461);
nor U8196 (N_8196,N_355,N_985);
or U8197 (N_8197,N_1079,N_1660);
or U8198 (N_8198,N_685,N_4498);
nand U8199 (N_8199,N_1476,N_2933);
and U8200 (N_8200,N_2255,N_3849);
nand U8201 (N_8201,N_5,N_3775);
and U8202 (N_8202,N_769,N_3292);
nand U8203 (N_8203,N_2482,N_1980);
nor U8204 (N_8204,N_158,N_3350);
and U8205 (N_8205,N_3570,N_3246);
and U8206 (N_8206,N_1578,N_2672);
or U8207 (N_8207,N_4792,N_3187);
and U8208 (N_8208,N_4382,N_3266);
nor U8209 (N_8209,N_1426,N_4488);
nand U8210 (N_8210,N_1474,N_1685);
nor U8211 (N_8211,N_344,N_451);
and U8212 (N_8212,N_4696,N_635);
nand U8213 (N_8213,N_4643,N_3571);
or U8214 (N_8214,N_1772,N_3212);
nor U8215 (N_8215,N_4860,N_3806);
nor U8216 (N_8216,N_1362,N_2236);
and U8217 (N_8217,N_2463,N_3152);
and U8218 (N_8218,N_4207,N_1377);
and U8219 (N_8219,N_4211,N_1724);
and U8220 (N_8220,N_3251,N_1023);
nor U8221 (N_8221,N_2683,N_1336);
or U8222 (N_8222,N_3539,N_272);
nor U8223 (N_8223,N_4343,N_4847);
and U8224 (N_8224,N_1783,N_346);
nor U8225 (N_8225,N_4764,N_1551);
nand U8226 (N_8226,N_4992,N_3590);
or U8227 (N_8227,N_4023,N_1723);
xnor U8228 (N_8228,N_3050,N_2221);
nand U8229 (N_8229,N_283,N_4793);
and U8230 (N_8230,N_4096,N_15);
nand U8231 (N_8231,N_1155,N_3165);
or U8232 (N_8232,N_4258,N_776);
nor U8233 (N_8233,N_4356,N_441);
nand U8234 (N_8234,N_3388,N_4771);
nand U8235 (N_8235,N_2438,N_2686);
nand U8236 (N_8236,N_1095,N_1569);
and U8237 (N_8237,N_618,N_4251);
nand U8238 (N_8238,N_1437,N_2126);
nor U8239 (N_8239,N_451,N_1124);
or U8240 (N_8240,N_887,N_731);
nor U8241 (N_8241,N_2963,N_4753);
and U8242 (N_8242,N_422,N_554);
nor U8243 (N_8243,N_375,N_3020);
or U8244 (N_8244,N_1374,N_3527);
and U8245 (N_8245,N_549,N_3977);
or U8246 (N_8246,N_4777,N_1088);
or U8247 (N_8247,N_854,N_3951);
nor U8248 (N_8248,N_3430,N_4537);
nor U8249 (N_8249,N_1706,N_4980);
nor U8250 (N_8250,N_1040,N_3557);
nor U8251 (N_8251,N_2880,N_276);
nand U8252 (N_8252,N_3319,N_687);
nor U8253 (N_8253,N_3251,N_704);
or U8254 (N_8254,N_2903,N_990);
or U8255 (N_8255,N_4580,N_4424);
nor U8256 (N_8256,N_4295,N_1322);
nand U8257 (N_8257,N_1636,N_4360);
nor U8258 (N_8258,N_3824,N_709);
nor U8259 (N_8259,N_2559,N_3330);
nor U8260 (N_8260,N_1883,N_3227);
and U8261 (N_8261,N_4775,N_2695);
and U8262 (N_8262,N_4886,N_2967);
or U8263 (N_8263,N_3646,N_17);
nand U8264 (N_8264,N_3019,N_2799);
or U8265 (N_8265,N_3639,N_4899);
nand U8266 (N_8266,N_4814,N_507);
or U8267 (N_8267,N_2360,N_36);
and U8268 (N_8268,N_977,N_844);
and U8269 (N_8269,N_181,N_1674);
and U8270 (N_8270,N_2770,N_3155);
nor U8271 (N_8271,N_4678,N_3741);
nor U8272 (N_8272,N_2088,N_4443);
or U8273 (N_8273,N_4468,N_3052);
and U8274 (N_8274,N_3137,N_4553);
and U8275 (N_8275,N_4746,N_1198);
nand U8276 (N_8276,N_876,N_2650);
nand U8277 (N_8277,N_2684,N_2955);
nand U8278 (N_8278,N_32,N_1790);
and U8279 (N_8279,N_904,N_704);
nand U8280 (N_8280,N_1630,N_2557);
nand U8281 (N_8281,N_145,N_3500);
nand U8282 (N_8282,N_3114,N_884);
and U8283 (N_8283,N_2816,N_1551);
or U8284 (N_8284,N_1561,N_3761);
and U8285 (N_8285,N_110,N_487);
xnor U8286 (N_8286,N_1562,N_2787);
nand U8287 (N_8287,N_85,N_3222);
or U8288 (N_8288,N_36,N_752);
nand U8289 (N_8289,N_2333,N_3261);
or U8290 (N_8290,N_3823,N_3078);
nand U8291 (N_8291,N_4564,N_1344);
and U8292 (N_8292,N_4915,N_1703);
nor U8293 (N_8293,N_4171,N_599);
nor U8294 (N_8294,N_1235,N_3068);
nand U8295 (N_8295,N_4294,N_3279);
nand U8296 (N_8296,N_3955,N_2130);
and U8297 (N_8297,N_3473,N_416);
or U8298 (N_8298,N_3217,N_940);
or U8299 (N_8299,N_1555,N_1170);
nor U8300 (N_8300,N_4770,N_4822);
xnor U8301 (N_8301,N_4281,N_1048);
and U8302 (N_8302,N_2966,N_271);
nor U8303 (N_8303,N_4198,N_406);
nor U8304 (N_8304,N_2947,N_4163);
nor U8305 (N_8305,N_3146,N_4717);
or U8306 (N_8306,N_477,N_4243);
and U8307 (N_8307,N_579,N_4926);
nand U8308 (N_8308,N_395,N_3451);
nand U8309 (N_8309,N_4056,N_4083);
or U8310 (N_8310,N_898,N_4587);
nor U8311 (N_8311,N_419,N_2943);
and U8312 (N_8312,N_1142,N_2970);
and U8313 (N_8313,N_2702,N_4510);
or U8314 (N_8314,N_3626,N_4944);
nand U8315 (N_8315,N_1294,N_1878);
nand U8316 (N_8316,N_1852,N_1086);
nand U8317 (N_8317,N_3023,N_1520);
nor U8318 (N_8318,N_2202,N_3704);
nand U8319 (N_8319,N_1900,N_1290);
or U8320 (N_8320,N_3079,N_1233);
nand U8321 (N_8321,N_2987,N_4279);
nand U8322 (N_8322,N_2254,N_3241);
and U8323 (N_8323,N_3147,N_1376);
and U8324 (N_8324,N_2003,N_3782);
xnor U8325 (N_8325,N_2567,N_4108);
and U8326 (N_8326,N_2736,N_4040);
and U8327 (N_8327,N_2762,N_3217);
and U8328 (N_8328,N_3558,N_2549);
nor U8329 (N_8329,N_514,N_2920);
and U8330 (N_8330,N_2795,N_169);
nand U8331 (N_8331,N_4913,N_2922);
nor U8332 (N_8332,N_450,N_1342);
nand U8333 (N_8333,N_1108,N_1583);
or U8334 (N_8334,N_650,N_4651);
and U8335 (N_8335,N_4420,N_4479);
nor U8336 (N_8336,N_3633,N_1713);
nor U8337 (N_8337,N_3777,N_2177);
nand U8338 (N_8338,N_4759,N_2867);
nor U8339 (N_8339,N_2376,N_752);
and U8340 (N_8340,N_3007,N_728);
and U8341 (N_8341,N_1876,N_4392);
xnor U8342 (N_8342,N_4533,N_3557);
nand U8343 (N_8343,N_1595,N_733);
or U8344 (N_8344,N_2098,N_3799);
nand U8345 (N_8345,N_3793,N_9);
and U8346 (N_8346,N_848,N_927);
or U8347 (N_8347,N_4483,N_1199);
nand U8348 (N_8348,N_3359,N_2479);
nand U8349 (N_8349,N_3497,N_431);
or U8350 (N_8350,N_2912,N_734);
nor U8351 (N_8351,N_2943,N_633);
or U8352 (N_8352,N_3186,N_2893);
or U8353 (N_8353,N_493,N_1132);
nor U8354 (N_8354,N_86,N_1429);
nand U8355 (N_8355,N_2375,N_4023);
nand U8356 (N_8356,N_2065,N_2680);
or U8357 (N_8357,N_3313,N_4177);
or U8358 (N_8358,N_33,N_4641);
nand U8359 (N_8359,N_329,N_3418);
nand U8360 (N_8360,N_2253,N_2223);
or U8361 (N_8361,N_4006,N_2514);
xnor U8362 (N_8362,N_333,N_4195);
nor U8363 (N_8363,N_2815,N_3826);
or U8364 (N_8364,N_1133,N_4760);
nand U8365 (N_8365,N_4524,N_2162);
or U8366 (N_8366,N_4783,N_574);
and U8367 (N_8367,N_4139,N_4810);
nor U8368 (N_8368,N_414,N_436);
nand U8369 (N_8369,N_1737,N_3818);
or U8370 (N_8370,N_831,N_3841);
or U8371 (N_8371,N_4406,N_2790);
nor U8372 (N_8372,N_4806,N_934);
and U8373 (N_8373,N_1949,N_1091);
nand U8374 (N_8374,N_4602,N_2556);
nor U8375 (N_8375,N_2797,N_1403);
or U8376 (N_8376,N_2064,N_1840);
and U8377 (N_8377,N_4751,N_1786);
nor U8378 (N_8378,N_4337,N_3028);
nor U8379 (N_8379,N_4252,N_163);
and U8380 (N_8380,N_1621,N_4925);
or U8381 (N_8381,N_3430,N_3597);
nand U8382 (N_8382,N_3553,N_3923);
nor U8383 (N_8383,N_2801,N_4960);
and U8384 (N_8384,N_2268,N_1676);
nand U8385 (N_8385,N_1330,N_164);
nor U8386 (N_8386,N_4188,N_3755);
or U8387 (N_8387,N_2962,N_425);
nor U8388 (N_8388,N_2253,N_705);
nor U8389 (N_8389,N_3412,N_4069);
and U8390 (N_8390,N_1601,N_3962);
nor U8391 (N_8391,N_4656,N_1873);
nand U8392 (N_8392,N_1091,N_1533);
and U8393 (N_8393,N_4932,N_2588);
nor U8394 (N_8394,N_509,N_969);
nor U8395 (N_8395,N_2034,N_222);
or U8396 (N_8396,N_1149,N_2463);
or U8397 (N_8397,N_3128,N_3125);
and U8398 (N_8398,N_2695,N_35);
nor U8399 (N_8399,N_725,N_2651);
or U8400 (N_8400,N_1075,N_2759);
or U8401 (N_8401,N_1338,N_1798);
nor U8402 (N_8402,N_3940,N_1783);
and U8403 (N_8403,N_59,N_4352);
nand U8404 (N_8404,N_3350,N_638);
nor U8405 (N_8405,N_454,N_2735);
and U8406 (N_8406,N_4898,N_2991);
nor U8407 (N_8407,N_2851,N_989);
nand U8408 (N_8408,N_4653,N_4961);
or U8409 (N_8409,N_4594,N_4264);
nor U8410 (N_8410,N_215,N_1695);
or U8411 (N_8411,N_1435,N_4853);
and U8412 (N_8412,N_1667,N_3994);
nand U8413 (N_8413,N_165,N_661);
or U8414 (N_8414,N_2657,N_2488);
nand U8415 (N_8415,N_1817,N_593);
or U8416 (N_8416,N_3290,N_1898);
nand U8417 (N_8417,N_3910,N_1979);
or U8418 (N_8418,N_3229,N_1239);
and U8419 (N_8419,N_3084,N_4263);
or U8420 (N_8420,N_4339,N_380);
nand U8421 (N_8421,N_480,N_2725);
and U8422 (N_8422,N_669,N_1984);
nor U8423 (N_8423,N_1539,N_2271);
nand U8424 (N_8424,N_646,N_4911);
nor U8425 (N_8425,N_4676,N_3641);
nor U8426 (N_8426,N_3888,N_4916);
or U8427 (N_8427,N_504,N_2755);
nand U8428 (N_8428,N_685,N_4505);
and U8429 (N_8429,N_2234,N_993);
and U8430 (N_8430,N_3757,N_4926);
or U8431 (N_8431,N_2524,N_1599);
or U8432 (N_8432,N_2239,N_1078);
nand U8433 (N_8433,N_4903,N_3229);
and U8434 (N_8434,N_3268,N_3105);
nor U8435 (N_8435,N_1307,N_4996);
and U8436 (N_8436,N_832,N_162);
nor U8437 (N_8437,N_494,N_3282);
or U8438 (N_8438,N_3732,N_789);
nor U8439 (N_8439,N_4018,N_1773);
and U8440 (N_8440,N_922,N_3345);
or U8441 (N_8441,N_919,N_2561);
nor U8442 (N_8442,N_968,N_2420);
or U8443 (N_8443,N_4224,N_3764);
nor U8444 (N_8444,N_2365,N_4860);
xor U8445 (N_8445,N_2261,N_3902);
xnor U8446 (N_8446,N_1518,N_2855);
xnor U8447 (N_8447,N_800,N_1744);
and U8448 (N_8448,N_4041,N_3824);
xnor U8449 (N_8449,N_1437,N_2177);
and U8450 (N_8450,N_1712,N_2996);
nor U8451 (N_8451,N_4450,N_3709);
nor U8452 (N_8452,N_4893,N_4327);
nor U8453 (N_8453,N_572,N_3939);
nand U8454 (N_8454,N_491,N_1387);
nand U8455 (N_8455,N_4389,N_3759);
nor U8456 (N_8456,N_2710,N_1694);
nand U8457 (N_8457,N_4679,N_2328);
nand U8458 (N_8458,N_4940,N_959);
nand U8459 (N_8459,N_4095,N_1759);
and U8460 (N_8460,N_80,N_3527);
nor U8461 (N_8461,N_870,N_363);
and U8462 (N_8462,N_260,N_898);
nor U8463 (N_8463,N_4776,N_4265);
or U8464 (N_8464,N_4835,N_158);
and U8465 (N_8465,N_1775,N_4116);
nor U8466 (N_8466,N_907,N_1097);
nor U8467 (N_8467,N_854,N_2730);
nand U8468 (N_8468,N_4094,N_2270);
and U8469 (N_8469,N_86,N_3);
or U8470 (N_8470,N_4139,N_429);
nor U8471 (N_8471,N_2227,N_2096);
nand U8472 (N_8472,N_2777,N_1393);
or U8473 (N_8473,N_4346,N_2370);
nand U8474 (N_8474,N_4831,N_3738);
and U8475 (N_8475,N_1972,N_2699);
or U8476 (N_8476,N_4393,N_3768);
or U8477 (N_8477,N_975,N_621);
nor U8478 (N_8478,N_3824,N_4132);
and U8479 (N_8479,N_2884,N_3343);
nor U8480 (N_8480,N_3555,N_741);
nand U8481 (N_8481,N_2129,N_2228);
or U8482 (N_8482,N_2781,N_3309);
and U8483 (N_8483,N_2838,N_4884);
or U8484 (N_8484,N_3510,N_4560);
nor U8485 (N_8485,N_2351,N_3800);
and U8486 (N_8486,N_4653,N_1410);
and U8487 (N_8487,N_2348,N_1819);
nor U8488 (N_8488,N_1414,N_3091);
nand U8489 (N_8489,N_3846,N_1853);
and U8490 (N_8490,N_3931,N_174);
or U8491 (N_8491,N_3922,N_1965);
nand U8492 (N_8492,N_3400,N_640);
nor U8493 (N_8493,N_1806,N_2949);
nor U8494 (N_8494,N_4413,N_2944);
and U8495 (N_8495,N_644,N_2375);
or U8496 (N_8496,N_14,N_105);
or U8497 (N_8497,N_1399,N_3722);
nand U8498 (N_8498,N_2563,N_1546);
or U8499 (N_8499,N_2361,N_691);
or U8500 (N_8500,N_2177,N_4323);
nand U8501 (N_8501,N_3329,N_4922);
nand U8502 (N_8502,N_1042,N_3556);
nand U8503 (N_8503,N_833,N_1690);
and U8504 (N_8504,N_3460,N_1154);
or U8505 (N_8505,N_4510,N_4677);
and U8506 (N_8506,N_1451,N_43);
xor U8507 (N_8507,N_607,N_3259);
nor U8508 (N_8508,N_27,N_2011);
or U8509 (N_8509,N_612,N_3105);
nor U8510 (N_8510,N_1842,N_1173);
or U8511 (N_8511,N_698,N_3026);
nor U8512 (N_8512,N_3550,N_1246);
or U8513 (N_8513,N_2212,N_4269);
nor U8514 (N_8514,N_4259,N_2608);
nand U8515 (N_8515,N_4624,N_304);
nor U8516 (N_8516,N_2200,N_2150);
or U8517 (N_8517,N_1489,N_3081);
or U8518 (N_8518,N_3432,N_1291);
and U8519 (N_8519,N_4271,N_1082);
or U8520 (N_8520,N_3496,N_1281);
xor U8521 (N_8521,N_3866,N_3886);
nand U8522 (N_8522,N_2548,N_1727);
nand U8523 (N_8523,N_1614,N_1180);
or U8524 (N_8524,N_4861,N_977);
nor U8525 (N_8525,N_196,N_1845);
or U8526 (N_8526,N_2864,N_4600);
nor U8527 (N_8527,N_1426,N_483);
nor U8528 (N_8528,N_713,N_1259);
or U8529 (N_8529,N_459,N_3213);
nor U8530 (N_8530,N_2745,N_4144);
nor U8531 (N_8531,N_4723,N_3555);
nor U8532 (N_8532,N_3590,N_1717);
and U8533 (N_8533,N_4531,N_2792);
nand U8534 (N_8534,N_3165,N_415);
and U8535 (N_8535,N_4659,N_4141);
nand U8536 (N_8536,N_2973,N_3763);
or U8537 (N_8537,N_3375,N_4446);
or U8538 (N_8538,N_2176,N_427);
or U8539 (N_8539,N_3038,N_542);
nor U8540 (N_8540,N_1715,N_1307);
or U8541 (N_8541,N_3795,N_4656);
nor U8542 (N_8542,N_1089,N_2995);
nor U8543 (N_8543,N_2937,N_4995);
nand U8544 (N_8544,N_4931,N_3463);
and U8545 (N_8545,N_2888,N_2348);
nor U8546 (N_8546,N_3269,N_4357);
and U8547 (N_8547,N_1611,N_3845);
and U8548 (N_8548,N_4007,N_2951);
and U8549 (N_8549,N_4462,N_1869);
and U8550 (N_8550,N_1705,N_2806);
and U8551 (N_8551,N_2860,N_2748);
or U8552 (N_8552,N_3602,N_3210);
nor U8553 (N_8553,N_139,N_4724);
nand U8554 (N_8554,N_46,N_4729);
nor U8555 (N_8555,N_4886,N_2676);
nand U8556 (N_8556,N_1965,N_2801);
nand U8557 (N_8557,N_4792,N_2913);
nand U8558 (N_8558,N_1243,N_4401);
nor U8559 (N_8559,N_3717,N_1993);
and U8560 (N_8560,N_4808,N_2114);
nand U8561 (N_8561,N_2071,N_4420);
nand U8562 (N_8562,N_2665,N_3145);
nand U8563 (N_8563,N_803,N_4099);
or U8564 (N_8564,N_240,N_120);
nor U8565 (N_8565,N_4680,N_552);
xor U8566 (N_8566,N_2791,N_1485);
nand U8567 (N_8567,N_2478,N_3847);
nor U8568 (N_8568,N_2568,N_3379);
nor U8569 (N_8569,N_2608,N_264);
nor U8570 (N_8570,N_1571,N_4599);
nand U8571 (N_8571,N_607,N_4210);
nor U8572 (N_8572,N_1454,N_600);
or U8573 (N_8573,N_2530,N_3203);
and U8574 (N_8574,N_1262,N_1711);
and U8575 (N_8575,N_2422,N_2651);
nor U8576 (N_8576,N_2110,N_2948);
nor U8577 (N_8577,N_2026,N_3263);
nor U8578 (N_8578,N_2813,N_1745);
nand U8579 (N_8579,N_2508,N_1201);
nor U8580 (N_8580,N_1850,N_9);
and U8581 (N_8581,N_3731,N_3366);
nor U8582 (N_8582,N_1591,N_45);
or U8583 (N_8583,N_3190,N_221);
or U8584 (N_8584,N_4872,N_2102);
or U8585 (N_8585,N_1716,N_4379);
nand U8586 (N_8586,N_389,N_902);
nor U8587 (N_8587,N_4966,N_2651);
or U8588 (N_8588,N_2917,N_2698);
or U8589 (N_8589,N_284,N_1224);
nor U8590 (N_8590,N_2090,N_70);
and U8591 (N_8591,N_2086,N_95);
or U8592 (N_8592,N_2979,N_2955);
or U8593 (N_8593,N_4287,N_2891);
nand U8594 (N_8594,N_420,N_2963);
or U8595 (N_8595,N_3085,N_101);
nand U8596 (N_8596,N_3302,N_251);
nand U8597 (N_8597,N_2502,N_2873);
nand U8598 (N_8598,N_1198,N_689);
or U8599 (N_8599,N_1314,N_3763);
or U8600 (N_8600,N_4076,N_3917);
nand U8601 (N_8601,N_4347,N_246);
and U8602 (N_8602,N_4920,N_920);
and U8603 (N_8603,N_2953,N_1040);
nand U8604 (N_8604,N_3439,N_3400);
or U8605 (N_8605,N_4776,N_867);
and U8606 (N_8606,N_395,N_471);
or U8607 (N_8607,N_2916,N_1708);
and U8608 (N_8608,N_1028,N_4151);
or U8609 (N_8609,N_279,N_2404);
xnor U8610 (N_8610,N_4715,N_4577);
nand U8611 (N_8611,N_3733,N_3954);
or U8612 (N_8612,N_1331,N_3074);
and U8613 (N_8613,N_3408,N_4981);
or U8614 (N_8614,N_3705,N_4173);
nor U8615 (N_8615,N_2587,N_3177);
or U8616 (N_8616,N_2659,N_1058);
or U8617 (N_8617,N_421,N_1837);
or U8618 (N_8618,N_4199,N_3761);
nor U8619 (N_8619,N_2751,N_600);
nand U8620 (N_8620,N_4858,N_3732);
nor U8621 (N_8621,N_190,N_361);
and U8622 (N_8622,N_2117,N_2539);
nand U8623 (N_8623,N_1733,N_4801);
nand U8624 (N_8624,N_3501,N_3880);
nand U8625 (N_8625,N_4090,N_3758);
nor U8626 (N_8626,N_94,N_1944);
and U8627 (N_8627,N_1487,N_1689);
nand U8628 (N_8628,N_2890,N_4854);
nor U8629 (N_8629,N_1670,N_4208);
or U8630 (N_8630,N_1983,N_2032);
nand U8631 (N_8631,N_1650,N_3744);
or U8632 (N_8632,N_4623,N_4122);
and U8633 (N_8633,N_3368,N_1414);
nor U8634 (N_8634,N_1841,N_4884);
xnor U8635 (N_8635,N_2050,N_2531);
or U8636 (N_8636,N_4743,N_4735);
or U8637 (N_8637,N_2298,N_791);
and U8638 (N_8638,N_2387,N_2919);
nor U8639 (N_8639,N_903,N_1423);
nand U8640 (N_8640,N_746,N_1344);
and U8641 (N_8641,N_3073,N_580);
nand U8642 (N_8642,N_2368,N_4106);
or U8643 (N_8643,N_2824,N_3890);
nand U8644 (N_8644,N_3067,N_2833);
or U8645 (N_8645,N_4826,N_2658);
nand U8646 (N_8646,N_4713,N_3155);
nor U8647 (N_8647,N_1470,N_752);
nor U8648 (N_8648,N_224,N_2457);
nor U8649 (N_8649,N_3706,N_2724);
or U8650 (N_8650,N_3361,N_4494);
or U8651 (N_8651,N_4590,N_2641);
or U8652 (N_8652,N_3273,N_757);
nand U8653 (N_8653,N_1602,N_3492);
nor U8654 (N_8654,N_2431,N_2882);
or U8655 (N_8655,N_1080,N_1391);
and U8656 (N_8656,N_2705,N_96);
and U8657 (N_8657,N_2309,N_3536);
and U8658 (N_8658,N_2574,N_3808);
or U8659 (N_8659,N_2623,N_3770);
or U8660 (N_8660,N_4391,N_3671);
or U8661 (N_8661,N_4350,N_1032);
nand U8662 (N_8662,N_1508,N_4539);
and U8663 (N_8663,N_3867,N_4406);
or U8664 (N_8664,N_331,N_4994);
or U8665 (N_8665,N_2127,N_4136);
nor U8666 (N_8666,N_4388,N_399);
and U8667 (N_8667,N_1328,N_873);
or U8668 (N_8668,N_1998,N_3551);
nand U8669 (N_8669,N_3134,N_2348);
or U8670 (N_8670,N_292,N_961);
nand U8671 (N_8671,N_959,N_447);
nor U8672 (N_8672,N_4202,N_4953);
nand U8673 (N_8673,N_2172,N_1653);
nand U8674 (N_8674,N_391,N_1743);
or U8675 (N_8675,N_1937,N_169);
nor U8676 (N_8676,N_2567,N_3201);
and U8677 (N_8677,N_2248,N_690);
nand U8678 (N_8678,N_2941,N_1306);
and U8679 (N_8679,N_3287,N_205);
nand U8680 (N_8680,N_118,N_294);
nand U8681 (N_8681,N_3518,N_198);
and U8682 (N_8682,N_1334,N_3935);
and U8683 (N_8683,N_4764,N_475);
nor U8684 (N_8684,N_3442,N_4701);
or U8685 (N_8685,N_3200,N_3906);
nor U8686 (N_8686,N_440,N_4397);
nor U8687 (N_8687,N_1648,N_2912);
nor U8688 (N_8688,N_3046,N_3680);
nor U8689 (N_8689,N_1028,N_47);
nor U8690 (N_8690,N_1228,N_1587);
or U8691 (N_8691,N_4013,N_875);
nor U8692 (N_8692,N_4798,N_1289);
nand U8693 (N_8693,N_4850,N_997);
or U8694 (N_8694,N_568,N_973);
nor U8695 (N_8695,N_132,N_1427);
or U8696 (N_8696,N_1893,N_1248);
or U8697 (N_8697,N_3610,N_367);
nor U8698 (N_8698,N_1543,N_1754);
nor U8699 (N_8699,N_3088,N_4219);
nand U8700 (N_8700,N_136,N_3925);
nand U8701 (N_8701,N_4369,N_46);
nand U8702 (N_8702,N_2504,N_1579);
and U8703 (N_8703,N_2481,N_1503);
and U8704 (N_8704,N_3795,N_31);
or U8705 (N_8705,N_754,N_3819);
or U8706 (N_8706,N_130,N_3348);
and U8707 (N_8707,N_1429,N_1736);
nand U8708 (N_8708,N_1997,N_2261);
and U8709 (N_8709,N_1818,N_2750);
and U8710 (N_8710,N_4851,N_1991);
and U8711 (N_8711,N_3990,N_461);
and U8712 (N_8712,N_2604,N_349);
and U8713 (N_8713,N_2390,N_1482);
and U8714 (N_8714,N_2079,N_4301);
nor U8715 (N_8715,N_3724,N_4593);
nor U8716 (N_8716,N_464,N_3929);
and U8717 (N_8717,N_1573,N_2644);
nor U8718 (N_8718,N_87,N_911);
and U8719 (N_8719,N_108,N_4156);
and U8720 (N_8720,N_1048,N_1054);
xnor U8721 (N_8721,N_1175,N_223);
and U8722 (N_8722,N_1055,N_44);
and U8723 (N_8723,N_2839,N_576);
and U8724 (N_8724,N_3688,N_2307);
or U8725 (N_8725,N_2280,N_573);
nand U8726 (N_8726,N_3071,N_4486);
nor U8727 (N_8727,N_2423,N_3059);
or U8728 (N_8728,N_893,N_1531);
and U8729 (N_8729,N_1867,N_3090);
or U8730 (N_8730,N_2097,N_152);
nand U8731 (N_8731,N_4193,N_223);
nor U8732 (N_8732,N_1020,N_1223);
and U8733 (N_8733,N_191,N_2974);
and U8734 (N_8734,N_1979,N_4847);
and U8735 (N_8735,N_2544,N_364);
and U8736 (N_8736,N_1024,N_687);
nand U8737 (N_8737,N_4519,N_3700);
or U8738 (N_8738,N_1158,N_1814);
and U8739 (N_8739,N_4813,N_2401);
or U8740 (N_8740,N_3747,N_415);
nor U8741 (N_8741,N_4006,N_262);
nand U8742 (N_8742,N_391,N_2830);
xor U8743 (N_8743,N_3936,N_2405);
nor U8744 (N_8744,N_3000,N_290);
xnor U8745 (N_8745,N_4767,N_835);
and U8746 (N_8746,N_3075,N_2071);
or U8747 (N_8747,N_1201,N_2489);
and U8748 (N_8748,N_4786,N_741);
nor U8749 (N_8749,N_318,N_1203);
nor U8750 (N_8750,N_2267,N_154);
or U8751 (N_8751,N_4305,N_4194);
nor U8752 (N_8752,N_800,N_840);
nand U8753 (N_8753,N_326,N_2485);
or U8754 (N_8754,N_2261,N_4572);
nand U8755 (N_8755,N_4613,N_1023);
nor U8756 (N_8756,N_1294,N_2430);
nand U8757 (N_8757,N_4922,N_2913);
or U8758 (N_8758,N_587,N_3522);
or U8759 (N_8759,N_3671,N_2872);
nand U8760 (N_8760,N_1988,N_677);
nand U8761 (N_8761,N_1800,N_226);
or U8762 (N_8762,N_2590,N_369);
and U8763 (N_8763,N_658,N_3625);
and U8764 (N_8764,N_1361,N_404);
nor U8765 (N_8765,N_106,N_1752);
or U8766 (N_8766,N_3715,N_1374);
or U8767 (N_8767,N_3118,N_2965);
nand U8768 (N_8768,N_899,N_2358);
nand U8769 (N_8769,N_1229,N_4033);
and U8770 (N_8770,N_2541,N_4106);
nand U8771 (N_8771,N_3427,N_2675);
nand U8772 (N_8772,N_1692,N_4888);
nand U8773 (N_8773,N_4534,N_2468);
nand U8774 (N_8774,N_2739,N_749);
or U8775 (N_8775,N_4155,N_3503);
and U8776 (N_8776,N_4957,N_516);
nor U8777 (N_8777,N_4897,N_2505);
nor U8778 (N_8778,N_4573,N_3239);
and U8779 (N_8779,N_3016,N_4126);
or U8780 (N_8780,N_4896,N_3841);
or U8781 (N_8781,N_4378,N_4931);
nor U8782 (N_8782,N_593,N_634);
nor U8783 (N_8783,N_69,N_1495);
and U8784 (N_8784,N_1596,N_2985);
nand U8785 (N_8785,N_2929,N_743);
and U8786 (N_8786,N_678,N_3291);
xnor U8787 (N_8787,N_987,N_3113);
nand U8788 (N_8788,N_2213,N_802);
nand U8789 (N_8789,N_980,N_97);
or U8790 (N_8790,N_3749,N_1729);
xor U8791 (N_8791,N_1620,N_2648);
nor U8792 (N_8792,N_4932,N_2409);
nand U8793 (N_8793,N_4493,N_3173);
or U8794 (N_8794,N_1958,N_4462);
or U8795 (N_8795,N_2007,N_3680);
and U8796 (N_8796,N_4320,N_325);
and U8797 (N_8797,N_3056,N_1103);
nand U8798 (N_8798,N_1024,N_355);
nor U8799 (N_8799,N_3018,N_2673);
and U8800 (N_8800,N_3986,N_1808);
and U8801 (N_8801,N_2739,N_1227);
or U8802 (N_8802,N_2792,N_1341);
or U8803 (N_8803,N_4646,N_2072);
nand U8804 (N_8804,N_3811,N_1620);
nor U8805 (N_8805,N_3964,N_2457);
or U8806 (N_8806,N_2270,N_4701);
and U8807 (N_8807,N_2079,N_1830);
or U8808 (N_8808,N_2309,N_664);
nor U8809 (N_8809,N_116,N_2666);
nand U8810 (N_8810,N_3456,N_661);
xor U8811 (N_8811,N_2816,N_4187);
or U8812 (N_8812,N_1707,N_560);
nand U8813 (N_8813,N_2613,N_162);
and U8814 (N_8814,N_2718,N_2306);
nand U8815 (N_8815,N_4044,N_1363);
nor U8816 (N_8816,N_1633,N_3932);
or U8817 (N_8817,N_3522,N_4673);
and U8818 (N_8818,N_2998,N_2533);
xor U8819 (N_8819,N_2256,N_1478);
nand U8820 (N_8820,N_712,N_2049);
nor U8821 (N_8821,N_434,N_1837);
nand U8822 (N_8822,N_436,N_2872);
nand U8823 (N_8823,N_4502,N_1188);
nand U8824 (N_8824,N_4235,N_1284);
or U8825 (N_8825,N_1450,N_3451);
nor U8826 (N_8826,N_1404,N_3829);
or U8827 (N_8827,N_116,N_2228);
and U8828 (N_8828,N_1296,N_2361);
and U8829 (N_8829,N_3896,N_3611);
nand U8830 (N_8830,N_2260,N_2482);
nor U8831 (N_8831,N_1552,N_4270);
and U8832 (N_8832,N_140,N_1619);
and U8833 (N_8833,N_1841,N_413);
nand U8834 (N_8834,N_499,N_3865);
nand U8835 (N_8835,N_550,N_4450);
nor U8836 (N_8836,N_4435,N_3127);
nor U8837 (N_8837,N_328,N_1065);
or U8838 (N_8838,N_770,N_4447);
and U8839 (N_8839,N_2947,N_3783);
and U8840 (N_8840,N_1346,N_3166);
and U8841 (N_8841,N_2314,N_4880);
nand U8842 (N_8842,N_3116,N_3946);
nor U8843 (N_8843,N_4275,N_120);
and U8844 (N_8844,N_1896,N_3886);
and U8845 (N_8845,N_233,N_2342);
or U8846 (N_8846,N_2833,N_1687);
and U8847 (N_8847,N_4590,N_663);
nor U8848 (N_8848,N_1346,N_3238);
nand U8849 (N_8849,N_1605,N_505);
or U8850 (N_8850,N_1865,N_3009);
nor U8851 (N_8851,N_376,N_3977);
and U8852 (N_8852,N_2412,N_2141);
or U8853 (N_8853,N_3175,N_369);
xnor U8854 (N_8854,N_4841,N_2836);
nor U8855 (N_8855,N_1746,N_4401);
or U8856 (N_8856,N_4976,N_1763);
or U8857 (N_8857,N_2352,N_1434);
and U8858 (N_8858,N_4244,N_2163);
nand U8859 (N_8859,N_3776,N_364);
and U8860 (N_8860,N_1623,N_4930);
or U8861 (N_8861,N_4977,N_4855);
or U8862 (N_8862,N_4876,N_152);
nand U8863 (N_8863,N_2351,N_4327);
and U8864 (N_8864,N_2152,N_4423);
nor U8865 (N_8865,N_395,N_2219);
or U8866 (N_8866,N_541,N_856);
or U8867 (N_8867,N_4212,N_2725);
xnor U8868 (N_8868,N_1117,N_4646);
and U8869 (N_8869,N_3673,N_3391);
and U8870 (N_8870,N_3793,N_4371);
or U8871 (N_8871,N_375,N_3168);
and U8872 (N_8872,N_3760,N_4743);
nor U8873 (N_8873,N_3575,N_93);
or U8874 (N_8874,N_1006,N_425);
or U8875 (N_8875,N_3346,N_349);
and U8876 (N_8876,N_2925,N_2627);
or U8877 (N_8877,N_4684,N_385);
nand U8878 (N_8878,N_4422,N_4748);
and U8879 (N_8879,N_3270,N_964);
and U8880 (N_8880,N_2057,N_2830);
nand U8881 (N_8881,N_1674,N_2856);
and U8882 (N_8882,N_2721,N_996);
or U8883 (N_8883,N_3205,N_3873);
or U8884 (N_8884,N_2864,N_1799);
or U8885 (N_8885,N_4565,N_2767);
and U8886 (N_8886,N_855,N_996);
and U8887 (N_8887,N_310,N_4276);
or U8888 (N_8888,N_830,N_2642);
nand U8889 (N_8889,N_2825,N_4842);
or U8890 (N_8890,N_1797,N_3915);
nor U8891 (N_8891,N_152,N_3011);
nand U8892 (N_8892,N_4684,N_11);
xor U8893 (N_8893,N_4120,N_1341);
nand U8894 (N_8894,N_1338,N_4876);
nor U8895 (N_8895,N_3111,N_1146);
nand U8896 (N_8896,N_1376,N_1920);
or U8897 (N_8897,N_3410,N_4626);
and U8898 (N_8898,N_4771,N_2014);
nor U8899 (N_8899,N_1887,N_2577);
nand U8900 (N_8900,N_1721,N_4845);
and U8901 (N_8901,N_2384,N_4842);
nand U8902 (N_8902,N_526,N_4809);
nand U8903 (N_8903,N_4804,N_3099);
and U8904 (N_8904,N_3977,N_4011);
and U8905 (N_8905,N_4804,N_973);
and U8906 (N_8906,N_4236,N_1882);
and U8907 (N_8907,N_803,N_1091);
or U8908 (N_8908,N_3869,N_1546);
or U8909 (N_8909,N_4216,N_1511);
or U8910 (N_8910,N_4139,N_2908);
or U8911 (N_8911,N_2000,N_1381);
nor U8912 (N_8912,N_2575,N_2547);
nand U8913 (N_8913,N_2232,N_2361);
or U8914 (N_8914,N_535,N_2442);
nor U8915 (N_8915,N_3494,N_618);
nor U8916 (N_8916,N_4386,N_2193);
and U8917 (N_8917,N_125,N_933);
nand U8918 (N_8918,N_3756,N_2913);
or U8919 (N_8919,N_196,N_1472);
nand U8920 (N_8920,N_1174,N_3651);
nand U8921 (N_8921,N_3654,N_4000);
or U8922 (N_8922,N_3791,N_2539);
or U8923 (N_8923,N_3510,N_939);
or U8924 (N_8924,N_4031,N_4633);
or U8925 (N_8925,N_153,N_3185);
nand U8926 (N_8926,N_2850,N_4185);
and U8927 (N_8927,N_3103,N_4293);
or U8928 (N_8928,N_1141,N_4577);
nor U8929 (N_8929,N_4465,N_1035);
nor U8930 (N_8930,N_4869,N_3578);
nor U8931 (N_8931,N_818,N_4242);
nand U8932 (N_8932,N_4798,N_1745);
nor U8933 (N_8933,N_1674,N_1965);
nor U8934 (N_8934,N_1045,N_949);
nand U8935 (N_8935,N_2498,N_294);
or U8936 (N_8936,N_552,N_893);
or U8937 (N_8937,N_2927,N_4290);
nand U8938 (N_8938,N_3127,N_91);
or U8939 (N_8939,N_2124,N_2480);
nor U8940 (N_8940,N_2129,N_2646);
nand U8941 (N_8941,N_4886,N_1447);
or U8942 (N_8942,N_917,N_2649);
and U8943 (N_8943,N_3410,N_2379);
nand U8944 (N_8944,N_752,N_726);
or U8945 (N_8945,N_3246,N_3020);
nand U8946 (N_8946,N_2425,N_255);
or U8947 (N_8947,N_1459,N_1482);
and U8948 (N_8948,N_2507,N_1545);
and U8949 (N_8949,N_607,N_1301);
and U8950 (N_8950,N_3371,N_1129);
and U8951 (N_8951,N_4974,N_1186);
nand U8952 (N_8952,N_3641,N_52);
nor U8953 (N_8953,N_677,N_3110);
and U8954 (N_8954,N_3233,N_2360);
nor U8955 (N_8955,N_346,N_1966);
or U8956 (N_8956,N_676,N_3220);
nor U8957 (N_8957,N_4153,N_75);
nand U8958 (N_8958,N_2091,N_497);
or U8959 (N_8959,N_74,N_2870);
or U8960 (N_8960,N_3094,N_4075);
and U8961 (N_8961,N_4688,N_956);
or U8962 (N_8962,N_772,N_1998);
nand U8963 (N_8963,N_1547,N_4525);
nor U8964 (N_8964,N_208,N_2667);
or U8965 (N_8965,N_1432,N_194);
or U8966 (N_8966,N_4815,N_4810);
nand U8967 (N_8967,N_3996,N_4204);
and U8968 (N_8968,N_1849,N_1559);
nand U8969 (N_8969,N_3687,N_2858);
nor U8970 (N_8970,N_4181,N_1823);
xnor U8971 (N_8971,N_3954,N_1499);
or U8972 (N_8972,N_4097,N_2076);
or U8973 (N_8973,N_2031,N_314);
or U8974 (N_8974,N_4090,N_1069);
and U8975 (N_8975,N_198,N_237);
nor U8976 (N_8976,N_1420,N_1008);
and U8977 (N_8977,N_2603,N_3603);
and U8978 (N_8978,N_2890,N_2558);
and U8979 (N_8979,N_1930,N_432);
and U8980 (N_8980,N_4988,N_581);
nor U8981 (N_8981,N_4079,N_1377);
or U8982 (N_8982,N_1027,N_380);
or U8983 (N_8983,N_690,N_674);
xor U8984 (N_8984,N_4459,N_1139);
and U8985 (N_8985,N_1135,N_3140);
or U8986 (N_8986,N_1194,N_2863);
nor U8987 (N_8987,N_3440,N_1643);
or U8988 (N_8988,N_4379,N_1254);
nor U8989 (N_8989,N_1644,N_1294);
or U8990 (N_8990,N_1379,N_4639);
nor U8991 (N_8991,N_4425,N_1726);
nor U8992 (N_8992,N_2242,N_2397);
nor U8993 (N_8993,N_1267,N_484);
or U8994 (N_8994,N_3715,N_1389);
and U8995 (N_8995,N_101,N_896);
nor U8996 (N_8996,N_719,N_3886);
nand U8997 (N_8997,N_3633,N_3927);
xnor U8998 (N_8998,N_1693,N_2749);
nand U8999 (N_8999,N_2859,N_3566);
nand U9000 (N_9000,N_2641,N_4970);
nand U9001 (N_9001,N_1488,N_3009);
and U9002 (N_9002,N_1274,N_4935);
or U9003 (N_9003,N_395,N_4230);
nand U9004 (N_9004,N_110,N_4252);
and U9005 (N_9005,N_2053,N_3469);
and U9006 (N_9006,N_368,N_2498);
and U9007 (N_9007,N_1990,N_2830);
and U9008 (N_9008,N_3438,N_2892);
nand U9009 (N_9009,N_1291,N_377);
nand U9010 (N_9010,N_2836,N_3551);
or U9011 (N_9011,N_4553,N_3800);
or U9012 (N_9012,N_56,N_626);
and U9013 (N_9013,N_3635,N_761);
nor U9014 (N_9014,N_22,N_1765);
or U9015 (N_9015,N_1326,N_3097);
or U9016 (N_9016,N_2728,N_4126);
nand U9017 (N_9017,N_1232,N_2422);
nand U9018 (N_9018,N_3567,N_488);
or U9019 (N_9019,N_4234,N_3569);
nor U9020 (N_9020,N_3414,N_3466);
and U9021 (N_9021,N_1853,N_2980);
or U9022 (N_9022,N_1406,N_3090);
and U9023 (N_9023,N_3636,N_3273);
and U9024 (N_9024,N_1963,N_4481);
nand U9025 (N_9025,N_618,N_3660);
or U9026 (N_9026,N_3763,N_4105);
or U9027 (N_9027,N_4690,N_3443);
and U9028 (N_9028,N_259,N_3122);
and U9029 (N_9029,N_4210,N_760);
nand U9030 (N_9030,N_4265,N_1913);
or U9031 (N_9031,N_2715,N_4315);
nor U9032 (N_9032,N_4728,N_1053);
or U9033 (N_9033,N_1982,N_4792);
nand U9034 (N_9034,N_4242,N_3168);
or U9035 (N_9035,N_3513,N_3169);
and U9036 (N_9036,N_4156,N_1956);
nor U9037 (N_9037,N_1421,N_804);
and U9038 (N_9038,N_3320,N_2222);
nand U9039 (N_9039,N_2383,N_4218);
nor U9040 (N_9040,N_4155,N_4219);
or U9041 (N_9041,N_4733,N_4910);
and U9042 (N_9042,N_3010,N_890);
and U9043 (N_9043,N_1557,N_1034);
nand U9044 (N_9044,N_3341,N_3345);
or U9045 (N_9045,N_3140,N_1174);
or U9046 (N_9046,N_844,N_4136);
or U9047 (N_9047,N_2647,N_4905);
or U9048 (N_9048,N_571,N_3932);
or U9049 (N_9049,N_4173,N_4977);
nand U9050 (N_9050,N_1982,N_665);
or U9051 (N_9051,N_48,N_3355);
or U9052 (N_9052,N_545,N_643);
or U9053 (N_9053,N_59,N_3272);
nand U9054 (N_9054,N_3287,N_697);
or U9055 (N_9055,N_1996,N_1016);
xnor U9056 (N_9056,N_3060,N_2982);
nor U9057 (N_9057,N_3345,N_916);
nor U9058 (N_9058,N_1179,N_1067);
xnor U9059 (N_9059,N_2900,N_582);
and U9060 (N_9060,N_1753,N_3746);
nand U9061 (N_9061,N_492,N_4140);
nor U9062 (N_9062,N_3927,N_659);
nor U9063 (N_9063,N_3782,N_605);
nor U9064 (N_9064,N_1915,N_3198);
xor U9065 (N_9065,N_3009,N_4704);
or U9066 (N_9066,N_367,N_3026);
nor U9067 (N_9067,N_3278,N_2658);
xor U9068 (N_9068,N_3641,N_848);
nor U9069 (N_9069,N_3278,N_4636);
or U9070 (N_9070,N_1044,N_4479);
nor U9071 (N_9071,N_1434,N_576);
or U9072 (N_9072,N_2104,N_653);
or U9073 (N_9073,N_3149,N_776);
nor U9074 (N_9074,N_1142,N_66);
and U9075 (N_9075,N_2663,N_2339);
nor U9076 (N_9076,N_2103,N_2837);
nor U9077 (N_9077,N_540,N_2733);
and U9078 (N_9078,N_2091,N_1561);
nor U9079 (N_9079,N_2489,N_4963);
nand U9080 (N_9080,N_2604,N_1679);
nand U9081 (N_9081,N_272,N_3606);
nor U9082 (N_9082,N_4739,N_3284);
nand U9083 (N_9083,N_423,N_1896);
or U9084 (N_9084,N_4566,N_1879);
nand U9085 (N_9085,N_2231,N_1048);
or U9086 (N_9086,N_3359,N_2220);
and U9087 (N_9087,N_303,N_617);
nand U9088 (N_9088,N_3486,N_877);
or U9089 (N_9089,N_2366,N_1214);
nor U9090 (N_9090,N_34,N_4276);
nand U9091 (N_9091,N_2465,N_4101);
and U9092 (N_9092,N_3303,N_1871);
nand U9093 (N_9093,N_4378,N_577);
or U9094 (N_9094,N_3859,N_3955);
nor U9095 (N_9095,N_3297,N_1840);
nand U9096 (N_9096,N_1009,N_63);
nor U9097 (N_9097,N_3207,N_1562);
nor U9098 (N_9098,N_1037,N_4768);
and U9099 (N_9099,N_562,N_4886);
nand U9100 (N_9100,N_681,N_2996);
nand U9101 (N_9101,N_2324,N_3053);
or U9102 (N_9102,N_4563,N_726);
nand U9103 (N_9103,N_1410,N_1320);
nor U9104 (N_9104,N_2910,N_4962);
and U9105 (N_9105,N_2837,N_1071);
and U9106 (N_9106,N_2493,N_1054);
nor U9107 (N_9107,N_394,N_1788);
nor U9108 (N_9108,N_3959,N_4580);
and U9109 (N_9109,N_1626,N_2947);
and U9110 (N_9110,N_72,N_4319);
and U9111 (N_9111,N_102,N_3687);
nor U9112 (N_9112,N_3992,N_4766);
and U9113 (N_9113,N_907,N_675);
nand U9114 (N_9114,N_1422,N_1832);
nand U9115 (N_9115,N_3839,N_1563);
nand U9116 (N_9116,N_2462,N_1110);
or U9117 (N_9117,N_171,N_2056);
and U9118 (N_9118,N_1039,N_4520);
nand U9119 (N_9119,N_1874,N_220);
and U9120 (N_9120,N_2566,N_1973);
nand U9121 (N_9121,N_3929,N_893);
nor U9122 (N_9122,N_875,N_2597);
and U9123 (N_9123,N_3522,N_2845);
or U9124 (N_9124,N_1531,N_1923);
nor U9125 (N_9125,N_2974,N_2416);
nor U9126 (N_9126,N_2015,N_1002);
nand U9127 (N_9127,N_1746,N_3115);
or U9128 (N_9128,N_1123,N_3421);
or U9129 (N_9129,N_3933,N_2813);
or U9130 (N_9130,N_487,N_2358);
and U9131 (N_9131,N_4445,N_3815);
or U9132 (N_9132,N_804,N_2602);
nand U9133 (N_9133,N_4566,N_4425);
and U9134 (N_9134,N_3384,N_2886);
xnor U9135 (N_9135,N_1504,N_2556);
nor U9136 (N_9136,N_1873,N_1703);
and U9137 (N_9137,N_3904,N_4864);
nand U9138 (N_9138,N_3578,N_1637);
nor U9139 (N_9139,N_4176,N_2841);
or U9140 (N_9140,N_1322,N_2484);
nor U9141 (N_9141,N_3206,N_4669);
xor U9142 (N_9142,N_1390,N_1855);
nand U9143 (N_9143,N_4770,N_4868);
nand U9144 (N_9144,N_4007,N_70);
and U9145 (N_9145,N_2618,N_2638);
nand U9146 (N_9146,N_20,N_2516);
and U9147 (N_9147,N_2807,N_3384);
nand U9148 (N_9148,N_1355,N_2452);
and U9149 (N_9149,N_3575,N_3774);
xnor U9150 (N_9150,N_4859,N_1561);
nor U9151 (N_9151,N_2737,N_14);
nor U9152 (N_9152,N_3771,N_3359);
nand U9153 (N_9153,N_2486,N_4591);
and U9154 (N_9154,N_736,N_271);
and U9155 (N_9155,N_1642,N_4347);
nand U9156 (N_9156,N_826,N_4360);
nor U9157 (N_9157,N_4720,N_1237);
nor U9158 (N_9158,N_3884,N_3441);
or U9159 (N_9159,N_3285,N_382);
or U9160 (N_9160,N_2070,N_1629);
nor U9161 (N_9161,N_2368,N_485);
nor U9162 (N_9162,N_4664,N_2807);
nand U9163 (N_9163,N_1762,N_746);
or U9164 (N_9164,N_260,N_3053);
nor U9165 (N_9165,N_2822,N_1605);
or U9166 (N_9166,N_1441,N_68);
nand U9167 (N_9167,N_3383,N_451);
nor U9168 (N_9168,N_1833,N_1668);
xor U9169 (N_9169,N_715,N_4371);
nand U9170 (N_9170,N_2997,N_60);
or U9171 (N_9171,N_4371,N_2407);
or U9172 (N_9172,N_4086,N_746);
nand U9173 (N_9173,N_4031,N_2302);
nand U9174 (N_9174,N_3101,N_1726);
and U9175 (N_9175,N_845,N_2274);
and U9176 (N_9176,N_3604,N_4630);
and U9177 (N_9177,N_761,N_1669);
or U9178 (N_9178,N_2481,N_2222);
nand U9179 (N_9179,N_2615,N_120);
and U9180 (N_9180,N_113,N_1363);
nor U9181 (N_9181,N_992,N_4058);
and U9182 (N_9182,N_3189,N_1082);
nand U9183 (N_9183,N_2021,N_4033);
nand U9184 (N_9184,N_2977,N_4563);
and U9185 (N_9185,N_3463,N_3386);
nor U9186 (N_9186,N_920,N_3426);
nand U9187 (N_9187,N_1143,N_4165);
and U9188 (N_9188,N_1192,N_4098);
nand U9189 (N_9189,N_4545,N_2919);
nor U9190 (N_9190,N_1203,N_1277);
and U9191 (N_9191,N_1838,N_3649);
nor U9192 (N_9192,N_2751,N_3026);
nor U9193 (N_9193,N_3574,N_3672);
or U9194 (N_9194,N_2906,N_2674);
and U9195 (N_9195,N_133,N_4702);
nor U9196 (N_9196,N_860,N_2701);
nor U9197 (N_9197,N_241,N_558);
nand U9198 (N_9198,N_1203,N_4990);
or U9199 (N_9199,N_4658,N_30);
or U9200 (N_9200,N_2882,N_1724);
xnor U9201 (N_9201,N_2321,N_3194);
and U9202 (N_9202,N_1104,N_3999);
and U9203 (N_9203,N_2001,N_3012);
nor U9204 (N_9204,N_2310,N_1940);
and U9205 (N_9205,N_3787,N_2579);
and U9206 (N_9206,N_3138,N_381);
and U9207 (N_9207,N_315,N_2243);
nor U9208 (N_9208,N_3364,N_2916);
nand U9209 (N_9209,N_3509,N_1629);
and U9210 (N_9210,N_1242,N_730);
nand U9211 (N_9211,N_4582,N_650);
and U9212 (N_9212,N_4211,N_3033);
nand U9213 (N_9213,N_1514,N_4172);
and U9214 (N_9214,N_4884,N_87);
or U9215 (N_9215,N_1195,N_2176);
and U9216 (N_9216,N_4488,N_1149);
or U9217 (N_9217,N_2048,N_3083);
and U9218 (N_9218,N_738,N_1548);
or U9219 (N_9219,N_2311,N_2393);
or U9220 (N_9220,N_3979,N_3528);
nand U9221 (N_9221,N_2216,N_1555);
nor U9222 (N_9222,N_1572,N_4590);
and U9223 (N_9223,N_3023,N_4406);
nand U9224 (N_9224,N_4409,N_2073);
nand U9225 (N_9225,N_2686,N_2018);
or U9226 (N_9226,N_4018,N_811);
nand U9227 (N_9227,N_1537,N_3824);
nor U9228 (N_9228,N_4481,N_245);
xnor U9229 (N_9229,N_790,N_3973);
and U9230 (N_9230,N_1409,N_3410);
and U9231 (N_9231,N_2647,N_1843);
nand U9232 (N_9232,N_3758,N_984);
nor U9233 (N_9233,N_1396,N_1390);
or U9234 (N_9234,N_2578,N_1362);
and U9235 (N_9235,N_998,N_2938);
or U9236 (N_9236,N_49,N_1180);
and U9237 (N_9237,N_3006,N_2279);
nor U9238 (N_9238,N_3614,N_4888);
nand U9239 (N_9239,N_3664,N_2452);
nand U9240 (N_9240,N_4203,N_413);
or U9241 (N_9241,N_1040,N_2753);
or U9242 (N_9242,N_2179,N_1240);
nor U9243 (N_9243,N_3156,N_4078);
nand U9244 (N_9244,N_1618,N_727);
xor U9245 (N_9245,N_418,N_3529);
or U9246 (N_9246,N_874,N_1947);
nor U9247 (N_9247,N_82,N_301);
and U9248 (N_9248,N_4161,N_4782);
nor U9249 (N_9249,N_1065,N_4270);
or U9250 (N_9250,N_1934,N_4040);
and U9251 (N_9251,N_414,N_1946);
nor U9252 (N_9252,N_4045,N_4686);
nand U9253 (N_9253,N_2362,N_543);
or U9254 (N_9254,N_3349,N_1642);
nand U9255 (N_9255,N_462,N_4652);
nand U9256 (N_9256,N_3659,N_1175);
nand U9257 (N_9257,N_1157,N_2568);
xnor U9258 (N_9258,N_1058,N_2437);
nor U9259 (N_9259,N_4300,N_510);
and U9260 (N_9260,N_1490,N_3129);
and U9261 (N_9261,N_397,N_4502);
nand U9262 (N_9262,N_4571,N_4168);
or U9263 (N_9263,N_2241,N_3540);
or U9264 (N_9264,N_458,N_1139);
nand U9265 (N_9265,N_4661,N_1617);
nand U9266 (N_9266,N_4954,N_4018);
nand U9267 (N_9267,N_2578,N_3115);
and U9268 (N_9268,N_3441,N_2953);
nor U9269 (N_9269,N_2503,N_851);
nand U9270 (N_9270,N_4827,N_3554);
xnor U9271 (N_9271,N_3995,N_3354);
or U9272 (N_9272,N_1867,N_4515);
nand U9273 (N_9273,N_4629,N_2705);
nand U9274 (N_9274,N_980,N_3577);
xor U9275 (N_9275,N_4888,N_4490);
nand U9276 (N_9276,N_3716,N_2343);
or U9277 (N_9277,N_1475,N_2939);
nand U9278 (N_9278,N_2910,N_436);
nand U9279 (N_9279,N_4545,N_4195);
or U9280 (N_9280,N_4117,N_1041);
nand U9281 (N_9281,N_3780,N_3514);
xnor U9282 (N_9282,N_870,N_1902);
and U9283 (N_9283,N_999,N_918);
nor U9284 (N_9284,N_1276,N_4181);
or U9285 (N_9285,N_2670,N_3165);
and U9286 (N_9286,N_4915,N_907);
and U9287 (N_9287,N_4502,N_716);
and U9288 (N_9288,N_558,N_1102);
and U9289 (N_9289,N_3993,N_2310);
or U9290 (N_9290,N_924,N_2641);
or U9291 (N_9291,N_1241,N_1597);
and U9292 (N_9292,N_3092,N_1339);
nor U9293 (N_9293,N_1705,N_2673);
or U9294 (N_9294,N_3649,N_1353);
xor U9295 (N_9295,N_3922,N_3832);
nand U9296 (N_9296,N_1890,N_3301);
or U9297 (N_9297,N_4105,N_1429);
nand U9298 (N_9298,N_2042,N_1978);
nand U9299 (N_9299,N_3075,N_1891);
nand U9300 (N_9300,N_2612,N_3267);
or U9301 (N_9301,N_2644,N_1688);
nand U9302 (N_9302,N_397,N_1280);
nor U9303 (N_9303,N_379,N_1286);
nand U9304 (N_9304,N_3633,N_636);
or U9305 (N_9305,N_103,N_3348);
nor U9306 (N_9306,N_4146,N_2638);
and U9307 (N_9307,N_634,N_1343);
or U9308 (N_9308,N_4283,N_1654);
nor U9309 (N_9309,N_3009,N_3635);
and U9310 (N_9310,N_3618,N_1352);
or U9311 (N_9311,N_433,N_907);
nand U9312 (N_9312,N_4477,N_2916);
nor U9313 (N_9313,N_4092,N_1731);
nor U9314 (N_9314,N_3941,N_3489);
or U9315 (N_9315,N_3076,N_1687);
nand U9316 (N_9316,N_4004,N_1176);
or U9317 (N_9317,N_1906,N_4720);
and U9318 (N_9318,N_4538,N_88);
nand U9319 (N_9319,N_833,N_4803);
or U9320 (N_9320,N_1702,N_1863);
or U9321 (N_9321,N_47,N_1540);
nand U9322 (N_9322,N_1112,N_3799);
nor U9323 (N_9323,N_4636,N_1058);
nor U9324 (N_9324,N_2160,N_2785);
nand U9325 (N_9325,N_450,N_4898);
nor U9326 (N_9326,N_1151,N_1970);
and U9327 (N_9327,N_3451,N_1873);
nand U9328 (N_9328,N_4860,N_2026);
nand U9329 (N_9329,N_256,N_965);
xor U9330 (N_9330,N_753,N_125);
nand U9331 (N_9331,N_4279,N_4820);
and U9332 (N_9332,N_2422,N_1833);
nand U9333 (N_9333,N_279,N_186);
nand U9334 (N_9334,N_4683,N_179);
nor U9335 (N_9335,N_20,N_3610);
nor U9336 (N_9336,N_1343,N_3583);
nor U9337 (N_9337,N_574,N_4786);
or U9338 (N_9338,N_3993,N_1694);
nand U9339 (N_9339,N_545,N_4051);
or U9340 (N_9340,N_681,N_1590);
and U9341 (N_9341,N_2379,N_2577);
nand U9342 (N_9342,N_4952,N_2543);
xnor U9343 (N_9343,N_3627,N_4451);
nand U9344 (N_9344,N_441,N_4257);
nand U9345 (N_9345,N_1965,N_2512);
and U9346 (N_9346,N_1573,N_339);
and U9347 (N_9347,N_2280,N_100);
nor U9348 (N_9348,N_2764,N_1924);
or U9349 (N_9349,N_3460,N_1261);
nor U9350 (N_9350,N_1804,N_4676);
and U9351 (N_9351,N_2185,N_2931);
nor U9352 (N_9352,N_1769,N_1412);
nor U9353 (N_9353,N_3192,N_2082);
nor U9354 (N_9354,N_1938,N_3456);
and U9355 (N_9355,N_638,N_4553);
nor U9356 (N_9356,N_521,N_381);
and U9357 (N_9357,N_508,N_604);
nand U9358 (N_9358,N_3877,N_4756);
and U9359 (N_9359,N_2323,N_818);
or U9360 (N_9360,N_671,N_44);
and U9361 (N_9361,N_3675,N_3259);
or U9362 (N_9362,N_1597,N_3776);
and U9363 (N_9363,N_1369,N_2671);
and U9364 (N_9364,N_4942,N_2861);
and U9365 (N_9365,N_2233,N_3152);
or U9366 (N_9366,N_1511,N_967);
nor U9367 (N_9367,N_1949,N_1392);
and U9368 (N_9368,N_1304,N_1553);
nand U9369 (N_9369,N_4873,N_1212);
and U9370 (N_9370,N_4194,N_3189);
and U9371 (N_9371,N_2308,N_2960);
and U9372 (N_9372,N_891,N_606);
or U9373 (N_9373,N_3494,N_727);
nand U9374 (N_9374,N_4496,N_3991);
nor U9375 (N_9375,N_1816,N_684);
nor U9376 (N_9376,N_4297,N_3446);
and U9377 (N_9377,N_664,N_2967);
and U9378 (N_9378,N_2591,N_10);
or U9379 (N_9379,N_200,N_4443);
and U9380 (N_9380,N_4186,N_3551);
or U9381 (N_9381,N_1732,N_3082);
or U9382 (N_9382,N_2400,N_3696);
nand U9383 (N_9383,N_559,N_33);
nand U9384 (N_9384,N_2642,N_1463);
nand U9385 (N_9385,N_116,N_528);
nand U9386 (N_9386,N_1332,N_981);
and U9387 (N_9387,N_1943,N_3756);
nand U9388 (N_9388,N_2552,N_231);
nand U9389 (N_9389,N_282,N_2098);
nor U9390 (N_9390,N_599,N_3602);
or U9391 (N_9391,N_1577,N_1015);
or U9392 (N_9392,N_2824,N_1558);
or U9393 (N_9393,N_68,N_3882);
nor U9394 (N_9394,N_2234,N_3098);
nand U9395 (N_9395,N_18,N_3423);
nand U9396 (N_9396,N_3847,N_3110);
nand U9397 (N_9397,N_248,N_1543);
and U9398 (N_9398,N_4178,N_2161);
or U9399 (N_9399,N_907,N_2504);
nor U9400 (N_9400,N_670,N_4791);
nand U9401 (N_9401,N_1243,N_50);
and U9402 (N_9402,N_2631,N_3010);
nand U9403 (N_9403,N_984,N_2663);
nand U9404 (N_9404,N_3715,N_1997);
and U9405 (N_9405,N_4082,N_2245);
nor U9406 (N_9406,N_1129,N_1240);
nand U9407 (N_9407,N_3998,N_2895);
nor U9408 (N_9408,N_1757,N_2658);
nor U9409 (N_9409,N_1403,N_842);
nor U9410 (N_9410,N_3833,N_3305);
or U9411 (N_9411,N_969,N_3425);
and U9412 (N_9412,N_1975,N_533);
nor U9413 (N_9413,N_1762,N_4138);
nor U9414 (N_9414,N_4488,N_4220);
nand U9415 (N_9415,N_517,N_26);
or U9416 (N_9416,N_4563,N_2394);
or U9417 (N_9417,N_3647,N_3386);
xnor U9418 (N_9418,N_2974,N_3910);
or U9419 (N_9419,N_1041,N_4063);
and U9420 (N_9420,N_2653,N_2103);
nor U9421 (N_9421,N_2335,N_987);
nand U9422 (N_9422,N_1367,N_323);
nand U9423 (N_9423,N_3937,N_2997);
and U9424 (N_9424,N_3565,N_3173);
nand U9425 (N_9425,N_174,N_4282);
nor U9426 (N_9426,N_965,N_3991);
nor U9427 (N_9427,N_664,N_1972);
and U9428 (N_9428,N_3229,N_2350);
and U9429 (N_9429,N_3482,N_2039);
or U9430 (N_9430,N_2833,N_48);
or U9431 (N_9431,N_614,N_1979);
or U9432 (N_9432,N_97,N_4716);
and U9433 (N_9433,N_1502,N_3236);
or U9434 (N_9434,N_2546,N_599);
nor U9435 (N_9435,N_4208,N_1496);
nor U9436 (N_9436,N_2855,N_3174);
nor U9437 (N_9437,N_2787,N_2000);
or U9438 (N_9438,N_3183,N_2728);
nor U9439 (N_9439,N_2273,N_929);
nand U9440 (N_9440,N_83,N_3153);
or U9441 (N_9441,N_1776,N_38);
nor U9442 (N_9442,N_1495,N_514);
and U9443 (N_9443,N_2570,N_1284);
nand U9444 (N_9444,N_3808,N_4917);
or U9445 (N_9445,N_4377,N_3529);
or U9446 (N_9446,N_581,N_3658);
and U9447 (N_9447,N_2036,N_4624);
or U9448 (N_9448,N_402,N_3056);
or U9449 (N_9449,N_2012,N_1434);
or U9450 (N_9450,N_3842,N_1536);
nor U9451 (N_9451,N_2396,N_4277);
and U9452 (N_9452,N_2785,N_707);
nand U9453 (N_9453,N_4137,N_188);
or U9454 (N_9454,N_3369,N_1551);
or U9455 (N_9455,N_4634,N_3615);
and U9456 (N_9456,N_106,N_3683);
or U9457 (N_9457,N_878,N_3536);
and U9458 (N_9458,N_261,N_3979);
and U9459 (N_9459,N_3530,N_3402);
or U9460 (N_9460,N_4581,N_912);
nand U9461 (N_9461,N_3629,N_21);
or U9462 (N_9462,N_679,N_562);
nor U9463 (N_9463,N_342,N_3875);
or U9464 (N_9464,N_1510,N_1059);
or U9465 (N_9465,N_4713,N_4786);
or U9466 (N_9466,N_2238,N_3559);
and U9467 (N_9467,N_4958,N_2486);
nand U9468 (N_9468,N_4463,N_2326);
nand U9469 (N_9469,N_3053,N_1698);
or U9470 (N_9470,N_3460,N_4672);
or U9471 (N_9471,N_2072,N_2951);
nor U9472 (N_9472,N_4308,N_2518);
or U9473 (N_9473,N_3602,N_346);
and U9474 (N_9474,N_2562,N_2116);
and U9475 (N_9475,N_4152,N_2927);
nor U9476 (N_9476,N_965,N_1897);
or U9477 (N_9477,N_4181,N_2077);
or U9478 (N_9478,N_1036,N_2798);
nor U9479 (N_9479,N_3557,N_1917);
or U9480 (N_9480,N_410,N_6);
or U9481 (N_9481,N_4404,N_3031);
nor U9482 (N_9482,N_4202,N_1841);
nand U9483 (N_9483,N_1846,N_1004);
nor U9484 (N_9484,N_3354,N_670);
nand U9485 (N_9485,N_4346,N_2413);
or U9486 (N_9486,N_1510,N_33);
nor U9487 (N_9487,N_4412,N_2932);
nand U9488 (N_9488,N_2828,N_2352);
nor U9489 (N_9489,N_2716,N_813);
nand U9490 (N_9490,N_4401,N_4488);
nand U9491 (N_9491,N_832,N_2529);
nor U9492 (N_9492,N_1618,N_4134);
and U9493 (N_9493,N_3357,N_4434);
or U9494 (N_9494,N_4898,N_3976);
nand U9495 (N_9495,N_902,N_2721);
or U9496 (N_9496,N_4227,N_3133);
nor U9497 (N_9497,N_2657,N_680);
or U9498 (N_9498,N_2512,N_3607);
or U9499 (N_9499,N_2680,N_3029);
nor U9500 (N_9500,N_708,N_135);
and U9501 (N_9501,N_3013,N_2812);
nor U9502 (N_9502,N_2238,N_2160);
nand U9503 (N_9503,N_149,N_3524);
or U9504 (N_9504,N_1570,N_1882);
nor U9505 (N_9505,N_1449,N_1670);
and U9506 (N_9506,N_3072,N_770);
xor U9507 (N_9507,N_2092,N_2271);
nor U9508 (N_9508,N_1334,N_953);
nor U9509 (N_9509,N_2922,N_8);
nor U9510 (N_9510,N_2963,N_2465);
nand U9511 (N_9511,N_3738,N_4715);
and U9512 (N_9512,N_1951,N_1906);
nand U9513 (N_9513,N_423,N_543);
nor U9514 (N_9514,N_257,N_3244);
nand U9515 (N_9515,N_560,N_1180);
and U9516 (N_9516,N_1594,N_2945);
and U9517 (N_9517,N_879,N_2872);
and U9518 (N_9518,N_4624,N_1523);
nand U9519 (N_9519,N_3587,N_3040);
and U9520 (N_9520,N_1134,N_2925);
and U9521 (N_9521,N_1260,N_2714);
and U9522 (N_9522,N_4933,N_770);
nand U9523 (N_9523,N_2033,N_4115);
nor U9524 (N_9524,N_2776,N_346);
and U9525 (N_9525,N_890,N_1232);
or U9526 (N_9526,N_2364,N_2805);
nand U9527 (N_9527,N_2668,N_2584);
nor U9528 (N_9528,N_300,N_1170);
nand U9529 (N_9529,N_3051,N_1351);
nor U9530 (N_9530,N_2253,N_3068);
nand U9531 (N_9531,N_2725,N_4264);
nor U9532 (N_9532,N_504,N_566);
or U9533 (N_9533,N_2662,N_4119);
and U9534 (N_9534,N_1225,N_3064);
or U9535 (N_9535,N_2198,N_4631);
and U9536 (N_9536,N_2560,N_1373);
nand U9537 (N_9537,N_449,N_2553);
nand U9538 (N_9538,N_1126,N_141);
nand U9539 (N_9539,N_247,N_2209);
xnor U9540 (N_9540,N_4521,N_3413);
or U9541 (N_9541,N_409,N_4927);
nand U9542 (N_9542,N_3714,N_4306);
nor U9543 (N_9543,N_506,N_4020);
and U9544 (N_9544,N_1467,N_210);
and U9545 (N_9545,N_2364,N_1221);
and U9546 (N_9546,N_4048,N_1081);
and U9547 (N_9547,N_213,N_4541);
nor U9548 (N_9548,N_1325,N_4466);
nor U9549 (N_9549,N_4241,N_2404);
or U9550 (N_9550,N_3938,N_4926);
nor U9551 (N_9551,N_3184,N_3447);
nand U9552 (N_9552,N_1552,N_4971);
nand U9553 (N_9553,N_1286,N_2935);
or U9554 (N_9554,N_2099,N_1721);
and U9555 (N_9555,N_886,N_2517);
or U9556 (N_9556,N_899,N_445);
nor U9557 (N_9557,N_615,N_635);
or U9558 (N_9558,N_1376,N_2757);
nand U9559 (N_9559,N_4869,N_3283);
and U9560 (N_9560,N_116,N_4560);
and U9561 (N_9561,N_1669,N_1847);
or U9562 (N_9562,N_3974,N_4762);
or U9563 (N_9563,N_2925,N_1073);
nand U9564 (N_9564,N_616,N_1760);
nor U9565 (N_9565,N_956,N_4646);
nor U9566 (N_9566,N_2135,N_1815);
nand U9567 (N_9567,N_4029,N_4786);
nor U9568 (N_9568,N_1362,N_900);
or U9569 (N_9569,N_3680,N_3528);
or U9570 (N_9570,N_1671,N_1135);
nand U9571 (N_9571,N_935,N_2036);
xor U9572 (N_9572,N_4526,N_257);
and U9573 (N_9573,N_2376,N_552);
and U9574 (N_9574,N_1185,N_2622);
nor U9575 (N_9575,N_662,N_665);
nor U9576 (N_9576,N_2389,N_3185);
nor U9577 (N_9577,N_1869,N_1745);
and U9578 (N_9578,N_2446,N_2621);
and U9579 (N_9579,N_2265,N_3531);
and U9580 (N_9580,N_854,N_3495);
nand U9581 (N_9581,N_1328,N_1379);
nor U9582 (N_9582,N_3624,N_792);
and U9583 (N_9583,N_2971,N_2122);
or U9584 (N_9584,N_3686,N_4105);
or U9585 (N_9585,N_2642,N_1491);
nand U9586 (N_9586,N_1456,N_391);
and U9587 (N_9587,N_1315,N_1738);
nor U9588 (N_9588,N_1343,N_1811);
or U9589 (N_9589,N_2845,N_3397);
nor U9590 (N_9590,N_3913,N_4057);
nand U9591 (N_9591,N_1766,N_4626);
nor U9592 (N_9592,N_2238,N_3761);
nand U9593 (N_9593,N_998,N_4368);
and U9594 (N_9594,N_476,N_2807);
or U9595 (N_9595,N_1140,N_1697);
and U9596 (N_9596,N_174,N_816);
nand U9597 (N_9597,N_2512,N_681);
or U9598 (N_9598,N_3388,N_626);
and U9599 (N_9599,N_575,N_1074);
or U9600 (N_9600,N_2125,N_3141);
xnor U9601 (N_9601,N_1599,N_4096);
nand U9602 (N_9602,N_997,N_1077);
nor U9603 (N_9603,N_2094,N_1323);
nand U9604 (N_9604,N_4417,N_448);
and U9605 (N_9605,N_2251,N_1322);
or U9606 (N_9606,N_2027,N_711);
or U9607 (N_9607,N_2592,N_2284);
and U9608 (N_9608,N_3671,N_4035);
nand U9609 (N_9609,N_581,N_2000);
and U9610 (N_9610,N_3737,N_129);
nor U9611 (N_9611,N_944,N_1321);
nor U9612 (N_9612,N_1454,N_4085);
nand U9613 (N_9613,N_301,N_704);
and U9614 (N_9614,N_1071,N_3818);
or U9615 (N_9615,N_1956,N_2397);
nor U9616 (N_9616,N_2020,N_2816);
and U9617 (N_9617,N_46,N_57);
or U9618 (N_9618,N_4434,N_3782);
and U9619 (N_9619,N_4513,N_56);
nor U9620 (N_9620,N_2592,N_2096);
nor U9621 (N_9621,N_4972,N_3487);
and U9622 (N_9622,N_3366,N_2423);
nor U9623 (N_9623,N_3520,N_992);
and U9624 (N_9624,N_3429,N_4311);
xnor U9625 (N_9625,N_1299,N_4233);
and U9626 (N_9626,N_2890,N_3557);
nor U9627 (N_9627,N_976,N_4234);
nand U9628 (N_9628,N_327,N_1951);
nand U9629 (N_9629,N_1266,N_4851);
nor U9630 (N_9630,N_58,N_1571);
or U9631 (N_9631,N_3478,N_842);
nand U9632 (N_9632,N_1819,N_4810);
nor U9633 (N_9633,N_3903,N_958);
nor U9634 (N_9634,N_2410,N_4088);
or U9635 (N_9635,N_3176,N_1156);
nor U9636 (N_9636,N_387,N_859);
nor U9637 (N_9637,N_4979,N_4627);
and U9638 (N_9638,N_1136,N_3263);
nor U9639 (N_9639,N_3299,N_2970);
xor U9640 (N_9640,N_566,N_4734);
nand U9641 (N_9641,N_1634,N_2599);
nor U9642 (N_9642,N_2321,N_4293);
or U9643 (N_9643,N_3724,N_2775);
nand U9644 (N_9644,N_3903,N_3976);
nor U9645 (N_9645,N_1830,N_4180);
nand U9646 (N_9646,N_2972,N_2654);
and U9647 (N_9647,N_3389,N_1979);
or U9648 (N_9648,N_1479,N_4218);
and U9649 (N_9649,N_406,N_1143);
xnor U9650 (N_9650,N_1927,N_1140);
and U9651 (N_9651,N_3101,N_141);
or U9652 (N_9652,N_485,N_3024);
or U9653 (N_9653,N_4667,N_1036);
nor U9654 (N_9654,N_2801,N_4323);
nand U9655 (N_9655,N_1654,N_1936);
nor U9656 (N_9656,N_3615,N_3838);
or U9657 (N_9657,N_2583,N_3303);
and U9658 (N_9658,N_2511,N_4011);
nor U9659 (N_9659,N_2597,N_4714);
and U9660 (N_9660,N_4196,N_2535);
nor U9661 (N_9661,N_311,N_635);
or U9662 (N_9662,N_4589,N_217);
nor U9663 (N_9663,N_685,N_1044);
nand U9664 (N_9664,N_1280,N_3846);
and U9665 (N_9665,N_2147,N_2485);
or U9666 (N_9666,N_3723,N_1574);
nor U9667 (N_9667,N_220,N_3256);
or U9668 (N_9668,N_2249,N_46);
and U9669 (N_9669,N_3643,N_1210);
or U9670 (N_9670,N_4257,N_4086);
and U9671 (N_9671,N_3821,N_3843);
nor U9672 (N_9672,N_1253,N_1169);
nand U9673 (N_9673,N_4383,N_3025);
nand U9674 (N_9674,N_2556,N_1761);
nor U9675 (N_9675,N_4058,N_2514);
and U9676 (N_9676,N_4417,N_3211);
or U9677 (N_9677,N_4245,N_1709);
or U9678 (N_9678,N_3736,N_843);
nor U9679 (N_9679,N_2246,N_534);
and U9680 (N_9680,N_1402,N_2158);
nor U9681 (N_9681,N_787,N_1986);
or U9682 (N_9682,N_2908,N_4958);
or U9683 (N_9683,N_3632,N_2458);
or U9684 (N_9684,N_4997,N_4731);
nor U9685 (N_9685,N_321,N_1145);
or U9686 (N_9686,N_4862,N_261);
nand U9687 (N_9687,N_2437,N_4841);
or U9688 (N_9688,N_4039,N_4265);
nand U9689 (N_9689,N_656,N_3290);
nand U9690 (N_9690,N_1311,N_129);
nor U9691 (N_9691,N_1318,N_2247);
nand U9692 (N_9692,N_770,N_935);
nand U9693 (N_9693,N_626,N_2543);
nand U9694 (N_9694,N_925,N_2661);
and U9695 (N_9695,N_3385,N_655);
or U9696 (N_9696,N_2457,N_3505);
nand U9697 (N_9697,N_4089,N_344);
nand U9698 (N_9698,N_3358,N_4520);
nor U9699 (N_9699,N_4674,N_3229);
nor U9700 (N_9700,N_768,N_1101);
and U9701 (N_9701,N_861,N_2391);
nor U9702 (N_9702,N_962,N_932);
and U9703 (N_9703,N_1827,N_635);
or U9704 (N_9704,N_1572,N_3100);
nand U9705 (N_9705,N_3484,N_2279);
or U9706 (N_9706,N_4603,N_3731);
xnor U9707 (N_9707,N_1187,N_3817);
or U9708 (N_9708,N_1159,N_3485);
and U9709 (N_9709,N_3921,N_2136);
nand U9710 (N_9710,N_2442,N_4145);
nand U9711 (N_9711,N_474,N_807);
or U9712 (N_9712,N_1673,N_1668);
nor U9713 (N_9713,N_3944,N_1365);
nand U9714 (N_9714,N_658,N_1726);
or U9715 (N_9715,N_2288,N_196);
or U9716 (N_9716,N_497,N_4908);
nand U9717 (N_9717,N_4696,N_3847);
and U9718 (N_9718,N_2171,N_4256);
or U9719 (N_9719,N_4546,N_3145);
nand U9720 (N_9720,N_1403,N_2478);
or U9721 (N_9721,N_2522,N_3858);
and U9722 (N_9722,N_4317,N_3267);
nor U9723 (N_9723,N_4591,N_199);
nor U9724 (N_9724,N_1781,N_2319);
and U9725 (N_9725,N_3105,N_2438);
nor U9726 (N_9726,N_4067,N_3473);
nor U9727 (N_9727,N_2554,N_2196);
nor U9728 (N_9728,N_3340,N_2287);
or U9729 (N_9729,N_2817,N_4361);
or U9730 (N_9730,N_61,N_4618);
nand U9731 (N_9731,N_2315,N_4791);
nand U9732 (N_9732,N_2675,N_1216);
nor U9733 (N_9733,N_2268,N_1710);
and U9734 (N_9734,N_1556,N_3180);
nor U9735 (N_9735,N_4505,N_1026);
xnor U9736 (N_9736,N_2367,N_143);
nor U9737 (N_9737,N_1113,N_1138);
and U9738 (N_9738,N_3352,N_3171);
nor U9739 (N_9739,N_2787,N_4744);
nor U9740 (N_9740,N_3974,N_171);
or U9741 (N_9741,N_1654,N_897);
or U9742 (N_9742,N_4058,N_3527);
or U9743 (N_9743,N_4687,N_2891);
and U9744 (N_9744,N_3843,N_3689);
and U9745 (N_9745,N_4168,N_4142);
and U9746 (N_9746,N_2312,N_1448);
or U9747 (N_9747,N_4429,N_867);
and U9748 (N_9748,N_1040,N_404);
and U9749 (N_9749,N_914,N_4889);
nor U9750 (N_9750,N_4049,N_4400);
nand U9751 (N_9751,N_1983,N_4697);
nand U9752 (N_9752,N_2599,N_4270);
and U9753 (N_9753,N_199,N_1515);
and U9754 (N_9754,N_1277,N_1893);
or U9755 (N_9755,N_1578,N_4942);
nor U9756 (N_9756,N_4672,N_4668);
and U9757 (N_9757,N_2065,N_3724);
nor U9758 (N_9758,N_3854,N_511);
and U9759 (N_9759,N_1220,N_2328);
nor U9760 (N_9760,N_1712,N_3969);
nand U9761 (N_9761,N_2485,N_995);
or U9762 (N_9762,N_3776,N_583);
nand U9763 (N_9763,N_2037,N_530);
and U9764 (N_9764,N_1884,N_4905);
nor U9765 (N_9765,N_2190,N_4782);
and U9766 (N_9766,N_2454,N_393);
nor U9767 (N_9767,N_1257,N_2795);
nor U9768 (N_9768,N_749,N_2092);
nor U9769 (N_9769,N_1289,N_1374);
and U9770 (N_9770,N_4226,N_238);
nor U9771 (N_9771,N_4255,N_4965);
and U9772 (N_9772,N_4678,N_512);
nand U9773 (N_9773,N_3702,N_3876);
or U9774 (N_9774,N_1578,N_4414);
xor U9775 (N_9775,N_3418,N_409);
and U9776 (N_9776,N_4356,N_1279);
or U9777 (N_9777,N_4643,N_2400);
nand U9778 (N_9778,N_441,N_4467);
nor U9779 (N_9779,N_3632,N_2251);
nand U9780 (N_9780,N_4490,N_221);
nor U9781 (N_9781,N_3560,N_3630);
or U9782 (N_9782,N_677,N_107);
nor U9783 (N_9783,N_1319,N_3178);
or U9784 (N_9784,N_1715,N_103);
or U9785 (N_9785,N_821,N_1927);
and U9786 (N_9786,N_1099,N_2784);
nor U9787 (N_9787,N_4981,N_3560);
nor U9788 (N_9788,N_1571,N_4799);
or U9789 (N_9789,N_4790,N_3418);
or U9790 (N_9790,N_2520,N_2188);
and U9791 (N_9791,N_1953,N_3773);
nor U9792 (N_9792,N_1386,N_2641);
nor U9793 (N_9793,N_2235,N_3935);
and U9794 (N_9794,N_4116,N_3811);
nand U9795 (N_9795,N_4860,N_2952);
or U9796 (N_9796,N_1881,N_4632);
or U9797 (N_9797,N_3487,N_3714);
or U9798 (N_9798,N_3780,N_2621);
and U9799 (N_9799,N_3996,N_1097);
and U9800 (N_9800,N_930,N_2337);
or U9801 (N_9801,N_4963,N_3893);
and U9802 (N_9802,N_2996,N_4946);
or U9803 (N_9803,N_3654,N_2347);
nor U9804 (N_9804,N_2778,N_225);
nand U9805 (N_9805,N_66,N_2459);
or U9806 (N_9806,N_3852,N_4702);
nand U9807 (N_9807,N_3368,N_1007);
or U9808 (N_9808,N_525,N_2532);
xnor U9809 (N_9809,N_3244,N_4552);
nand U9810 (N_9810,N_1229,N_26);
or U9811 (N_9811,N_3316,N_4990);
or U9812 (N_9812,N_3131,N_3751);
nor U9813 (N_9813,N_602,N_2449);
nand U9814 (N_9814,N_1789,N_3145);
and U9815 (N_9815,N_1419,N_2590);
and U9816 (N_9816,N_2725,N_3626);
nor U9817 (N_9817,N_4079,N_2417);
or U9818 (N_9818,N_4032,N_4240);
xnor U9819 (N_9819,N_3954,N_1997);
nor U9820 (N_9820,N_412,N_2107);
and U9821 (N_9821,N_3632,N_920);
and U9822 (N_9822,N_3959,N_1594);
or U9823 (N_9823,N_3202,N_1693);
nor U9824 (N_9824,N_3955,N_985);
and U9825 (N_9825,N_530,N_1319);
and U9826 (N_9826,N_2475,N_1143);
and U9827 (N_9827,N_49,N_4086);
nand U9828 (N_9828,N_2679,N_2535);
nand U9829 (N_9829,N_2513,N_518);
nor U9830 (N_9830,N_2073,N_4862);
nor U9831 (N_9831,N_2122,N_2812);
nor U9832 (N_9832,N_2394,N_2369);
or U9833 (N_9833,N_3621,N_284);
or U9834 (N_9834,N_1759,N_1344);
nand U9835 (N_9835,N_4246,N_3397);
and U9836 (N_9836,N_4133,N_806);
and U9837 (N_9837,N_3439,N_2749);
or U9838 (N_9838,N_2149,N_1706);
nor U9839 (N_9839,N_4547,N_1729);
and U9840 (N_9840,N_714,N_3654);
nand U9841 (N_9841,N_4273,N_2817);
xnor U9842 (N_9842,N_4046,N_167);
or U9843 (N_9843,N_1883,N_4641);
nand U9844 (N_9844,N_1709,N_4567);
or U9845 (N_9845,N_2676,N_2842);
nand U9846 (N_9846,N_4749,N_343);
or U9847 (N_9847,N_1442,N_4868);
nand U9848 (N_9848,N_4215,N_685);
nor U9849 (N_9849,N_2845,N_206);
and U9850 (N_9850,N_4733,N_4041);
and U9851 (N_9851,N_3368,N_2600);
nand U9852 (N_9852,N_340,N_3410);
and U9853 (N_9853,N_120,N_2787);
nor U9854 (N_9854,N_4770,N_1184);
and U9855 (N_9855,N_73,N_3173);
nor U9856 (N_9856,N_2674,N_2340);
or U9857 (N_9857,N_477,N_2463);
or U9858 (N_9858,N_3097,N_593);
or U9859 (N_9859,N_3033,N_2165);
or U9860 (N_9860,N_4220,N_747);
or U9861 (N_9861,N_3422,N_807);
or U9862 (N_9862,N_3373,N_874);
xor U9863 (N_9863,N_1446,N_3349);
and U9864 (N_9864,N_181,N_3618);
nor U9865 (N_9865,N_3199,N_58);
and U9866 (N_9866,N_3492,N_2387);
nor U9867 (N_9867,N_4417,N_4801);
nor U9868 (N_9868,N_2230,N_3765);
and U9869 (N_9869,N_1189,N_2747);
nor U9870 (N_9870,N_1740,N_706);
and U9871 (N_9871,N_4863,N_3498);
and U9872 (N_9872,N_650,N_1018);
or U9873 (N_9873,N_4314,N_4839);
or U9874 (N_9874,N_64,N_1159);
nand U9875 (N_9875,N_1095,N_3145);
or U9876 (N_9876,N_2450,N_3260);
xnor U9877 (N_9877,N_4719,N_1120);
nor U9878 (N_9878,N_3514,N_612);
nand U9879 (N_9879,N_4615,N_3033);
nand U9880 (N_9880,N_4380,N_1203);
and U9881 (N_9881,N_548,N_3125);
nor U9882 (N_9882,N_3742,N_2235);
nor U9883 (N_9883,N_3580,N_3673);
nor U9884 (N_9884,N_1523,N_2339);
nand U9885 (N_9885,N_4027,N_3625);
nor U9886 (N_9886,N_922,N_4671);
or U9887 (N_9887,N_3043,N_4247);
or U9888 (N_9888,N_2068,N_2485);
or U9889 (N_9889,N_4513,N_1419);
and U9890 (N_9890,N_1975,N_1139);
or U9891 (N_9891,N_4050,N_264);
and U9892 (N_9892,N_2789,N_3373);
nand U9893 (N_9893,N_1985,N_4440);
or U9894 (N_9894,N_4673,N_1372);
nor U9895 (N_9895,N_2530,N_2866);
and U9896 (N_9896,N_1278,N_342);
nand U9897 (N_9897,N_1855,N_3463);
nor U9898 (N_9898,N_2799,N_3008);
or U9899 (N_9899,N_1152,N_1048);
nand U9900 (N_9900,N_2198,N_1907);
nor U9901 (N_9901,N_143,N_3175);
and U9902 (N_9902,N_4277,N_522);
or U9903 (N_9903,N_3117,N_4475);
nor U9904 (N_9904,N_2305,N_2495);
and U9905 (N_9905,N_3656,N_3134);
and U9906 (N_9906,N_2904,N_2261);
and U9907 (N_9907,N_2717,N_454);
and U9908 (N_9908,N_3856,N_2660);
nand U9909 (N_9909,N_3955,N_2234);
or U9910 (N_9910,N_879,N_743);
or U9911 (N_9911,N_3693,N_2956);
or U9912 (N_9912,N_4702,N_2310);
or U9913 (N_9913,N_1115,N_4756);
nor U9914 (N_9914,N_413,N_518);
nor U9915 (N_9915,N_4917,N_2496);
or U9916 (N_9916,N_4026,N_332);
nand U9917 (N_9917,N_1879,N_1781);
or U9918 (N_9918,N_1648,N_4153);
nand U9919 (N_9919,N_4702,N_2928);
nor U9920 (N_9920,N_1446,N_1365);
nand U9921 (N_9921,N_3700,N_4156);
or U9922 (N_9922,N_2079,N_4809);
nor U9923 (N_9923,N_3663,N_481);
nor U9924 (N_9924,N_3004,N_1539);
nor U9925 (N_9925,N_2507,N_163);
nand U9926 (N_9926,N_4391,N_3158);
and U9927 (N_9927,N_3322,N_898);
and U9928 (N_9928,N_548,N_4506);
xor U9929 (N_9929,N_4216,N_606);
and U9930 (N_9930,N_216,N_4636);
nor U9931 (N_9931,N_1888,N_1069);
and U9932 (N_9932,N_3131,N_223);
and U9933 (N_9933,N_2315,N_4960);
nand U9934 (N_9934,N_706,N_3452);
or U9935 (N_9935,N_4795,N_2814);
and U9936 (N_9936,N_2893,N_2565);
and U9937 (N_9937,N_106,N_3844);
or U9938 (N_9938,N_1387,N_2482);
or U9939 (N_9939,N_1727,N_3876);
or U9940 (N_9940,N_4645,N_589);
nand U9941 (N_9941,N_1973,N_3664);
or U9942 (N_9942,N_4494,N_2583);
nor U9943 (N_9943,N_4121,N_3694);
or U9944 (N_9944,N_651,N_1302);
or U9945 (N_9945,N_224,N_1363);
and U9946 (N_9946,N_3051,N_2178);
nor U9947 (N_9947,N_4416,N_142);
or U9948 (N_9948,N_3731,N_2566);
nand U9949 (N_9949,N_3357,N_4765);
or U9950 (N_9950,N_3183,N_1380);
nor U9951 (N_9951,N_2463,N_3307);
nand U9952 (N_9952,N_1099,N_4161);
nor U9953 (N_9953,N_1156,N_4210);
nand U9954 (N_9954,N_1826,N_4955);
or U9955 (N_9955,N_2635,N_4346);
or U9956 (N_9956,N_3494,N_4028);
and U9957 (N_9957,N_3639,N_4996);
xnor U9958 (N_9958,N_4743,N_2360);
or U9959 (N_9959,N_4887,N_1521);
xnor U9960 (N_9960,N_4508,N_4775);
and U9961 (N_9961,N_4181,N_865);
nand U9962 (N_9962,N_3031,N_845);
and U9963 (N_9963,N_3529,N_4329);
and U9964 (N_9964,N_4186,N_916);
and U9965 (N_9965,N_3995,N_3555);
or U9966 (N_9966,N_424,N_688);
and U9967 (N_9967,N_3672,N_2362);
nand U9968 (N_9968,N_4238,N_981);
nand U9969 (N_9969,N_2885,N_3153);
nor U9970 (N_9970,N_2927,N_248);
and U9971 (N_9971,N_2282,N_3457);
nor U9972 (N_9972,N_2271,N_1280);
nand U9973 (N_9973,N_2678,N_1893);
or U9974 (N_9974,N_1547,N_542);
or U9975 (N_9975,N_2626,N_4202);
and U9976 (N_9976,N_303,N_4800);
nor U9977 (N_9977,N_1908,N_3617);
nand U9978 (N_9978,N_1439,N_481);
nand U9979 (N_9979,N_3268,N_144);
or U9980 (N_9980,N_1865,N_3778);
xor U9981 (N_9981,N_2876,N_2953);
and U9982 (N_9982,N_2954,N_4290);
and U9983 (N_9983,N_839,N_4882);
nand U9984 (N_9984,N_1780,N_4999);
nor U9985 (N_9985,N_3074,N_3909);
nor U9986 (N_9986,N_3564,N_3273);
nand U9987 (N_9987,N_1002,N_3154);
nor U9988 (N_9988,N_1080,N_1377);
nand U9989 (N_9989,N_2853,N_208);
or U9990 (N_9990,N_184,N_571);
nor U9991 (N_9991,N_4209,N_4505);
nor U9992 (N_9992,N_4711,N_4036);
or U9993 (N_9993,N_1198,N_3710);
nor U9994 (N_9994,N_1600,N_988);
nand U9995 (N_9995,N_4527,N_4396);
and U9996 (N_9996,N_81,N_4143);
nand U9997 (N_9997,N_1773,N_3973);
xnor U9998 (N_9998,N_4220,N_1591);
and U9999 (N_9999,N_3839,N_2015);
nor U10000 (N_10000,N_7285,N_6970);
nand U10001 (N_10001,N_6764,N_6605);
and U10002 (N_10002,N_5928,N_7794);
and U10003 (N_10003,N_8181,N_7309);
nand U10004 (N_10004,N_9920,N_6301);
nand U10005 (N_10005,N_5651,N_6910);
or U10006 (N_10006,N_6164,N_8330);
or U10007 (N_10007,N_9123,N_5958);
or U10008 (N_10008,N_6741,N_7022);
nand U10009 (N_10009,N_8363,N_5657);
nand U10010 (N_10010,N_7833,N_8458);
nor U10011 (N_10011,N_6429,N_5310);
and U10012 (N_10012,N_6510,N_9073);
nor U10013 (N_10013,N_7166,N_8172);
nand U10014 (N_10014,N_9353,N_7547);
nand U10015 (N_10015,N_9784,N_6616);
and U10016 (N_10016,N_6427,N_5685);
nand U10017 (N_10017,N_8326,N_6537);
nor U10018 (N_10018,N_6243,N_7897);
nor U10019 (N_10019,N_6881,N_7327);
and U10020 (N_10020,N_5127,N_7753);
and U10021 (N_10021,N_6481,N_8527);
nor U10022 (N_10022,N_7164,N_7893);
nor U10023 (N_10023,N_8377,N_6543);
nor U10024 (N_10024,N_9650,N_7203);
nor U10025 (N_10025,N_7644,N_5041);
or U10026 (N_10026,N_9805,N_5481);
and U10027 (N_10027,N_6830,N_6604);
nor U10028 (N_10028,N_7548,N_6308);
or U10029 (N_10029,N_8317,N_5272);
xnor U10030 (N_10030,N_8985,N_9846);
and U10031 (N_10031,N_5751,N_6240);
nor U10032 (N_10032,N_5290,N_8255);
nor U10033 (N_10033,N_9514,N_6114);
and U10034 (N_10034,N_8052,N_7000);
nand U10035 (N_10035,N_6412,N_7229);
nand U10036 (N_10036,N_9535,N_5355);
and U10037 (N_10037,N_9182,N_6438);
nand U10038 (N_10038,N_8637,N_5443);
nand U10039 (N_10039,N_9088,N_8288);
nand U10040 (N_10040,N_6181,N_9627);
nand U10041 (N_10041,N_5352,N_5548);
or U10042 (N_10042,N_8014,N_6572);
or U10043 (N_10043,N_8203,N_5071);
and U10044 (N_10044,N_7387,N_5211);
or U10045 (N_10045,N_7865,N_7881);
nand U10046 (N_10046,N_9665,N_7236);
and U10047 (N_10047,N_7058,N_7190);
nor U10048 (N_10048,N_6128,N_6546);
nand U10049 (N_10049,N_6231,N_8510);
and U10050 (N_10050,N_6701,N_9610);
and U10051 (N_10051,N_9845,N_7671);
and U10052 (N_10052,N_5347,N_7146);
or U10053 (N_10053,N_7351,N_8420);
or U10054 (N_10054,N_7450,N_5594);
nor U10055 (N_10055,N_7515,N_7007);
or U10056 (N_10056,N_6050,N_8666);
nor U10057 (N_10057,N_9761,N_9573);
or U10058 (N_10058,N_6133,N_5439);
or U10059 (N_10059,N_7418,N_8170);
nand U10060 (N_10060,N_6769,N_7696);
or U10061 (N_10061,N_9951,N_6669);
and U10062 (N_10062,N_8596,N_6400);
nand U10063 (N_10063,N_7322,N_8214);
nor U10064 (N_10064,N_7323,N_9750);
and U10065 (N_10065,N_6614,N_7402);
or U10066 (N_10066,N_6383,N_7597);
nand U10067 (N_10067,N_7304,N_5907);
and U10068 (N_10068,N_7261,N_6459);
and U10069 (N_10069,N_6313,N_7148);
nor U10070 (N_10070,N_5329,N_6109);
or U10071 (N_10071,N_5479,N_6361);
or U10072 (N_10072,N_5277,N_9460);
nor U10073 (N_10073,N_9205,N_8444);
nor U10074 (N_10074,N_6152,N_5328);
or U10075 (N_10075,N_9221,N_8428);
nand U10076 (N_10076,N_9033,N_6282);
nand U10077 (N_10077,N_8164,N_9608);
nor U10078 (N_10078,N_5399,N_5823);
nand U10079 (N_10079,N_6319,N_5701);
nor U10080 (N_10080,N_9624,N_8879);
nand U10081 (N_10081,N_9904,N_6677);
nand U10082 (N_10082,N_7421,N_6552);
and U10083 (N_10083,N_6086,N_8445);
and U10084 (N_10084,N_8774,N_6148);
nand U10085 (N_10085,N_8163,N_9029);
nor U10086 (N_10086,N_9444,N_9990);
nand U10087 (N_10087,N_7562,N_6999);
and U10088 (N_10088,N_9870,N_5551);
nor U10089 (N_10089,N_8638,N_5540);
nor U10090 (N_10090,N_5693,N_8342);
nor U10091 (N_10091,N_5286,N_6872);
and U10092 (N_10092,N_9612,N_9212);
and U10093 (N_10093,N_6306,N_6463);
and U10094 (N_10094,N_8231,N_7225);
nand U10095 (N_10095,N_8154,N_7006);
and U10096 (N_10096,N_5935,N_6321);
or U10097 (N_10097,N_5408,N_8921);
nor U10098 (N_10098,N_5858,N_6487);
and U10099 (N_10099,N_8837,N_8339);
nand U10100 (N_10100,N_6227,N_5558);
and U10101 (N_10101,N_7014,N_7708);
nor U10102 (N_10102,N_9397,N_5047);
nor U10103 (N_10103,N_6281,N_7847);
nor U10104 (N_10104,N_9325,N_7274);
or U10105 (N_10105,N_5044,N_7937);
nand U10106 (N_10106,N_8625,N_9433);
nor U10107 (N_10107,N_9749,N_6254);
nor U10108 (N_10108,N_6868,N_9216);
nand U10109 (N_10109,N_5856,N_9897);
or U10110 (N_10110,N_9948,N_8304);
nor U10111 (N_10111,N_5948,N_6143);
and U10112 (N_10112,N_9151,N_7518);
or U10113 (N_10113,N_5215,N_9927);
nand U10114 (N_10114,N_5738,N_8605);
nor U10115 (N_10115,N_5792,N_6327);
and U10116 (N_10116,N_5300,N_9137);
nor U10117 (N_10117,N_5975,N_6250);
nor U10118 (N_10118,N_6278,N_5267);
or U10119 (N_10119,N_5798,N_9259);
xnor U10120 (N_10120,N_6234,N_7314);
nand U10121 (N_10121,N_8150,N_8733);
nand U10122 (N_10122,N_9127,N_6731);
and U10123 (N_10123,N_9268,N_5203);
or U10124 (N_10124,N_7997,N_9304);
and U10125 (N_10125,N_8455,N_9168);
nand U10126 (N_10126,N_9368,N_5592);
and U10127 (N_10127,N_9365,N_6906);
nand U10128 (N_10128,N_9344,N_8912);
nor U10129 (N_10129,N_7767,N_7894);
nand U10130 (N_10130,N_6009,N_6055);
nor U10131 (N_10131,N_5430,N_9234);
or U10132 (N_10132,N_6131,N_6146);
or U10133 (N_10133,N_6751,N_7487);
and U10134 (N_10134,N_9655,N_7496);
xnor U10135 (N_10135,N_5445,N_7552);
xor U10136 (N_10136,N_8907,N_5518);
and U10137 (N_10137,N_5569,N_6905);
nor U10138 (N_10138,N_9968,N_7021);
nand U10139 (N_10139,N_7991,N_7919);
nand U10140 (N_10140,N_6388,N_5354);
xor U10141 (N_10141,N_5861,N_9395);
and U10142 (N_10142,N_7337,N_9889);
and U10143 (N_10143,N_9380,N_7590);
nor U10144 (N_10144,N_7163,N_9989);
xnor U10145 (N_10145,N_8616,N_8206);
nand U10146 (N_10146,N_9131,N_5442);
nor U10147 (N_10147,N_6809,N_6532);
nand U10148 (N_10148,N_9780,N_6837);
and U10149 (N_10149,N_7423,N_7295);
and U10150 (N_10150,N_9469,N_9668);
nand U10151 (N_10151,N_8465,N_6026);
nor U10152 (N_10152,N_8081,N_7061);
nor U10153 (N_10153,N_9019,N_8303);
nand U10154 (N_10154,N_5253,N_9426);
nand U10155 (N_10155,N_6293,N_7840);
nor U10156 (N_10156,N_8419,N_5417);
nor U10157 (N_10157,N_7425,N_5593);
nor U10158 (N_10158,N_7916,N_7125);
nor U10159 (N_10159,N_8015,N_5421);
and U10160 (N_10160,N_7710,N_9851);
nor U10161 (N_10161,N_9915,N_8668);
or U10162 (N_10162,N_7167,N_9464);
nor U10163 (N_10163,N_8624,N_6199);
and U10164 (N_10164,N_8253,N_9299);
or U10165 (N_10165,N_9038,N_5862);
and U10166 (N_10166,N_7020,N_7267);
and U10167 (N_10167,N_7876,N_9058);
and U10168 (N_10168,N_6835,N_9917);
and U10169 (N_10169,N_7650,N_6207);
or U10170 (N_10170,N_6822,N_7481);
nand U10171 (N_10171,N_5833,N_7711);
nor U10172 (N_10172,N_5464,N_7660);
or U10173 (N_10173,N_7630,N_8327);
nor U10174 (N_10174,N_6350,N_7041);
or U10175 (N_10175,N_5115,N_7943);
and U10176 (N_10176,N_8710,N_5017);
nor U10177 (N_10177,N_7089,N_5100);
nand U10178 (N_10178,N_7106,N_5212);
nand U10179 (N_10179,N_7294,N_5447);
xnor U10180 (N_10180,N_8427,N_8088);
nor U10181 (N_10181,N_6948,N_7098);
or U10182 (N_10182,N_8134,N_8022);
or U10183 (N_10183,N_8090,N_9626);
or U10184 (N_10184,N_5346,N_9160);
nor U10185 (N_10185,N_5252,N_5634);
or U10186 (N_10186,N_9829,N_6525);
and U10187 (N_10187,N_8116,N_9934);
and U10188 (N_10188,N_6723,N_8277);
and U10189 (N_10189,N_6493,N_8992);
nor U10190 (N_10190,N_5987,N_7349);
nor U10191 (N_10191,N_8513,N_6628);
nand U10192 (N_10192,N_9601,N_7700);
nand U10193 (N_10193,N_7506,N_8740);
and U10194 (N_10194,N_5138,N_5200);
or U10195 (N_10195,N_5670,N_6989);
nor U10196 (N_10196,N_6567,N_8548);
or U10197 (N_10197,N_8798,N_7498);
or U10198 (N_10198,N_6272,N_9370);
or U10199 (N_10199,N_6887,N_8386);
nor U10200 (N_10200,N_7617,N_9119);
or U10201 (N_10201,N_6937,N_7502);
xnor U10202 (N_10202,N_8948,N_8208);
nand U10203 (N_10203,N_5638,N_6395);
or U10204 (N_10204,N_8604,N_5002);
and U10205 (N_10205,N_8323,N_7177);
or U10206 (N_10206,N_7510,N_8533);
xnor U10207 (N_10207,N_8660,N_7382);
nor U10208 (N_10208,N_9276,N_5322);
nor U10209 (N_10209,N_5040,N_6579);
and U10210 (N_10210,N_6640,N_9702);
and U10211 (N_10211,N_7279,N_5112);
and U10212 (N_10212,N_5938,N_5343);
xor U10213 (N_10213,N_7761,N_7026);
and U10214 (N_10214,N_8285,N_7601);
and U10215 (N_10215,N_5461,N_7795);
nand U10216 (N_10216,N_8600,N_9609);
or U10217 (N_10217,N_6680,N_9682);
nand U10218 (N_10218,N_8401,N_9978);
nand U10219 (N_10219,N_6967,N_6985);
and U10220 (N_10220,N_9318,N_5678);
or U10221 (N_10221,N_9252,N_7352);
or U10222 (N_10222,N_9054,N_5029);
nor U10223 (N_10223,N_5660,N_9223);
and U10224 (N_10224,N_6834,N_8443);
nand U10225 (N_10225,N_5591,N_8389);
and U10226 (N_10226,N_6574,N_5315);
and U10227 (N_10227,N_5295,N_9499);
nor U10228 (N_10228,N_7676,N_7582);
or U10229 (N_10229,N_7675,N_5389);
nor U10230 (N_10230,N_9579,N_6670);
and U10231 (N_10231,N_9218,N_5639);
and U10232 (N_10232,N_7479,N_6602);
nand U10233 (N_10233,N_7565,N_9706);
nand U10234 (N_10234,N_6266,N_5018);
and U10235 (N_10235,N_6144,N_7200);
nand U10236 (N_10236,N_8628,N_6716);
and U10237 (N_10237,N_6918,N_6955);
and U10238 (N_10238,N_7830,N_8071);
and U10239 (N_10239,N_7107,N_9675);
and U10240 (N_10240,N_9109,N_5304);
nor U10241 (N_10241,N_6084,N_7988);
and U10242 (N_10242,N_7374,N_5799);
nand U10243 (N_10243,N_8030,N_6924);
and U10244 (N_10244,N_8937,N_8158);
nor U10245 (N_10245,N_7204,N_9312);
or U10246 (N_10246,N_5719,N_6735);
and U10247 (N_10247,N_7420,N_6775);
nand U10248 (N_10248,N_8129,N_8571);
and U10249 (N_10249,N_6829,N_5788);
and U10250 (N_10250,N_9742,N_7731);
or U10251 (N_10251,N_6894,N_6288);
or U10252 (N_10252,N_7090,N_6208);
nand U10253 (N_10253,N_8518,N_5013);
and U10254 (N_10254,N_6428,N_6023);
and U10255 (N_10255,N_8464,N_9028);
or U10256 (N_10256,N_5407,N_7180);
nand U10257 (N_10257,N_8562,N_9485);
or U10258 (N_10258,N_6218,N_5760);
nand U10259 (N_10259,N_8369,N_8563);
nor U10260 (N_10260,N_5469,N_6619);
or U10261 (N_10261,N_7931,N_9906);
and U10262 (N_10262,N_8366,N_9497);
xnor U10263 (N_10263,N_7029,N_5073);
nand U10264 (N_10264,N_5208,N_8019);
and U10265 (N_10265,N_5883,N_6569);
nand U10266 (N_10266,N_9023,N_8822);
nand U10267 (N_10267,N_5288,N_5960);
nor U10268 (N_10268,N_8475,N_6486);
and U10269 (N_10269,N_8058,N_7380);
nand U10270 (N_10270,N_9577,N_7371);
nor U10271 (N_10271,N_6859,N_9139);
nor U10272 (N_10272,N_6936,N_8067);
nand U10273 (N_10273,N_8699,N_8582);
or U10274 (N_10274,N_9465,N_5618);
or U10275 (N_10275,N_5801,N_8402);
nand U10276 (N_10276,N_8580,N_5713);
xor U10277 (N_10277,N_7717,N_7213);
nor U10278 (N_10278,N_9885,N_8639);
or U10279 (N_10279,N_6307,N_6334);
and U10280 (N_10280,N_5381,N_5658);
or U10281 (N_10281,N_5214,N_7614);
or U10282 (N_10282,N_6824,N_7212);
nor U10283 (N_10283,N_6064,N_5980);
nand U10284 (N_10284,N_7867,N_7832);
or U10285 (N_10285,N_5985,N_5366);
and U10286 (N_10286,N_6401,N_9301);
and U10287 (N_10287,N_7193,N_7333);
or U10288 (N_10288,N_5285,N_5458);
nor U10289 (N_10289,N_6638,N_9138);
and U10290 (N_10290,N_8099,N_6591);
nor U10291 (N_10291,N_9207,N_5494);
and U10292 (N_10292,N_7612,N_6944);
xnor U10293 (N_10293,N_9687,N_9129);
nor U10294 (N_10294,N_7680,N_8190);
or U10295 (N_10295,N_7205,N_8051);
and U10296 (N_10296,N_6729,N_7470);
nand U10297 (N_10297,N_5722,N_9393);
and U10298 (N_10298,N_8577,N_6509);
and U10299 (N_10299,N_9891,N_5613);
nor U10300 (N_10300,N_6817,N_9521);
nand U10301 (N_10301,N_7191,N_7608);
nor U10302 (N_10302,N_9701,N_9183);
and U10303 (N_10303,N_6903,N_6177);
nand U10304 (N_10304,N_9554,N_7490);
and U10305 (N_10305,N_9560,N_9993);
nand U10306 (N_10306,N_8499,N_6041);
and U10307 (N_10307,N_6149,N_8784);
nor U10308 (N_10308,N_5140,N_7604);
nand U10309 (N_10309,N_7035,N_9507);
and U10310 (N_10310,N_9970,N_8125);
or U10311 (N_10311,N_7571,N_8260);
nor U10312 (N_10312,N_8523,N_6326);
or U10313 (N_10313,N_9636,N_8529);
or U10314 (N_10314,N_9495,N_6523);
nand U10315 (N_10315,N_9941,N_5635);
nor U10316 (N_10316,N_6566,N_9518);
or U10317 (N_10317,N_8292,N_6507);
and U10318 (N_10318,N_5522,N_7275);
or U10319 (N_10319,N_6928,N_5683);
nand U10320 (N_10320,N_5153,N_9728);
nand U10321 (N_10321,N_8996,N_5934);
nor U10322 (N_10322,N_5394,N_5106);
and U10323 (N_10323,N_9913,N_8632);
nor U10324 (N_10324,N_8576,N_6245);
nor U10325 (N_10325,N_5500,N_5096);
or U10326 (N_10326,N_5945,N_9716);
and U10327 (N_10327,N_6380,N_5240);
nor U10328 (N_10328,N_8805,N_7281);
nor U10329 (N_10329,N_7122,N_5832);
nor U10330 (N_10330,N_5180,N_9901);
nand U10331 (N_10331,N_9826,N_7049);
or U10332 (N_10332,N_6382,N_7299);
nand U10333 (N_10333,N_7248,N_7367);
or U10334 (N_10334,N_8298,N_5213);
and U10335 (N_10335,N_5537,N_5852);
or U10336 (N_10336,N_7398,N_7097);
and U10337 (N_10337,N_8944,N_8631);
nand U10338 (N_10338,N_6742,N_5275);
nor U10339 (N_10339,N_7960,N_7720);
nand U10340 (N_10340,N_7341,N_9621);
nand U10341 (N_10341,N_7264,N_5675);
nor U10342 (N_10342,N_9606,N_9463);
nand U10343 (N_10343,N_5111,N_5667);
nor U10344 (N_10344,N_8209,N_8815);
nor U10345 (N_10345,N_6727,N_9104);
and U10346 (N_10346,N_8459,N_7113);
nand U10347 (N_10347,N_7395,N_6930);
nor U10348 (N_10348,N_8578,N_8845);
nand U10349 (N_10349,N_8957,N_7230);
and U10350 (N_10350,N_8955,N_6404);
and U10351 (N_10351,N_6171,N_6103);
nand U10352 (N_10352,N_9817,N_9721);
nand U10353 (N_10353,N_5911,N_5444);
nor U10354 (N_10354,N_8685,N_9201);
nor U10355 (N_10355,N_6940,N_7554);
and U10356 (N_10356,N_9258,N_6981);
and U10357 (N_10357,N_7912,N_9653);
and U10358 (N_10358,N_5955,N_7160);
or U10359 (N_10359,N_8642,N_9337);
and U10360 (N_10360,N_9413,N_7348);
or U10361 (N_10361,N_7385,N_5089);
nand U10362 (N_10362,N_9288,N_9146);
nor U10363 (N_10363,N_5769,N_8640);
or U10364 (N_10364,N_7640,N_7593);
nor U10365 (N_10365,N_7201,N_5098);
and U10366 (N_10366,N_5113,N_8535);
nor U10367 (N_10367,N_6949,N_5508);
and U10368 (N_10368,N_7189,N_7632);
nand U10369 (N_10369,N_7269,N_5341);
nor U10370 (N_10370,N_5133,N_5094);
nor U10371 (N_10371,N_8110,N_6469);
xnor U10372 (N_10372,N_7768,N_5405);
nor U10373 (N_10373,N_6004,N_6352);
or U10374 (N_10374,N_9354,N_7084);
and U10375 (N_10375,N_8738,N_9166);
and U10376 (N_10376,N_8602,N_8078);
or U10377 (N_10377,N_8020,N_5129);
nor U10378 (N_10378,N_6213,N_6860);
nand U10379 (N_10379,N_6778,N_6538);
nand U10380 (N_10380,N_5564,N_8036);
or U10381 (N_10381,N_9068,N_9583);
or U10382 (N_10382,N_6202,N_5117);
nand U10383 (N_10383,N_9032,N_6205);
or U10384 (N_10384,N_6375,N_6984);
or U10385 (N_10385,N_9747,N_7667);
and U10386 (N_10386,N_6494,N_8528);
and U10387 (N_10387,N_6974,N_9000);
or U10388 (N_10388,N_8794,N_9003);
or U10389 (N_10389,N_6687,N_5142);
nand U10390 (N_10390,N_8112,N_8320);
and U10391 (N_10391,N_7968,N_5109);
and U10392 (N_10392,N_5107,N_5541);
and U10393 (N_10393,N_7219,N_7484);
and U10394 (N_10394,N_9740,N_8601);
or U10395 (N_10395,N_9593,N_6719);
or U10396 (N_10396,N_8612,N_9625);
nor U10397 (N_10397,N_6060,N_7482);
or U10398 (N_10398,N_8573,N_8313);
nand U10399 (N_10399,N_6908,N_7625);
or U10400 (N_10400,N_9331,N_8831);
or U10401 (N_10401,N_6754,N_8338);
and U10402 (N_10402,N_6795,N_7953);
or U10403 (N_10403,N_9273,N_7272);
or U10404 (N_10404,N_7643,N_9417);
nor U10405 (N_10405,N_8848,N_6374);
and U10406 (N_10406,N_9734,N_7331);
nand U10407 (N_10407,N_7540,N_6006);
nand U10408 (N_10408,N_5470,N_7393);
and U10409 (N_10409,N_8057,N_9001);
and U10410 (N_10410,N_6798,N_8745);
nor U10411 (N_10411,N_5642,N_5779);
nand U10412 (N_10412,N_7024,N_7779);
or U10413 (N_10413,N_8187,N_6066);
nor U10414 (N_10414,N_8244,N_7679);
nand U10415 (N_10415,N_9434,N_7312);
nor U10416 (N_10416,N_9095,N_6875);
or U10417 (N_10417,N_6444,N_7973);
nor U10418 (N_10418,N_8804,N_7172);
nor U10419 (N_10419,N_9775,N_6479);
nor U10420 (N_10420,N_6563,N_7971);
or U10421 (N_10421,N_5493,N_5104);
or U10422 (N_10422,N_9456,N_5229);
nand U10423 (N_10423,N_8031,N_7055);
and U10424 (N_10424,N_6709,N_8176);
nand U10425 (N_10425,N_6449,N_6675);
and U10426 (N_10426,N_7358,N_8314);
nor U10427 (N_10427,N_7882,N_6115);
nor U10428 (N_10428,N_5726,N_6200);
xor U10429 (N_10429,N_9284,N_6190);
and U10430 (N_10430,N_7899,N_8149);
nor U10431 (N_10431,N_5489,N_8603);
and U10432 (N_10432,N_9523,N_5482);
nor U10433 (N_10433,N_6220,N_7197);
and U10434 (N_10434,N_9963,N_6134);
or U10435 (N_10435,N_7032,N_5590);
or U10436 (N_10436,N_8273,N_7568);
and U10437 (N_10437,N_5636,N_6414);
nor U10438 (N_10438,N_5772,N_7414);
nor U10439 (N_10439,N_7884,N_8991);
nor U10440 (N_10440,N_9087,N_9987);
nand U10441 (N_10441,N_7462,N_8073);
and U10442 (N_10442,N_6216,N_7709);
or U10443 (N_10443,N_9164,N_9149);
nand U10444 (N_10444,N_6242,N_8915);
nor U10445 (N_10445,N_7362,N_7137);
and U10446 (N_10446,N_5531,N_8761);
and U10447 (N_10447,N_5156,N_9388);
nand U10448 (N_10448,N_7086,N_8156);
nor U10449 (N_10449,N_9106,N_7819);
and U10450 (N_10450,N_6472,N_7366);
nor U10451 (N_10451,N_7871,N_6789);
nand U10452 (N_10452,N_7218,N_5588);
and U10453 (N_10453,N_8440,N_8439);
nand U10454 (N_10454,N_9219,N_9004);
or U10455 (N_10455,N_7737,N_6214);
or U10456 (N_10456,N_5307,N_5246);
nor U10457 (N_10457,N_5785,N_9458);
or U10458 (N_10458,N_9524,N_7474);
or U10459 (N_10459,N_8230,N_8433);
nor U10460 (N_10460,N_5308,N_6298);
or U10461 (N_10461,N_7436,N_7639);
and U10462 (N_10462,N_7196,N_5720);
nor U10463 (N_10463,N_6416,N_6237);
nand U10464 (N_10464,N_7188,N_5155);
nand U10465 (N_10465,N_9454,N_5737);
nor U10466 (N_10466,N_9931,N_7375);
nor U10467 (N_10467,N_8343,N_5969);
nor U10468 (N_10468,N_9572,N_7182);
or U10469 (N_10469,N_9392,N_7658);
nor U10470 (N_10470,N_8516,N_6154);
and U10471 (N_10471,N_6738,N_7079);
nor U10472 (N_10472,N_5392,N_7745);
and U10473 (N_10473,N_6273,N_5375);
nor U10474 (N_10474,N_8372,N_5640);
nand U10475 (N_10475,N_9666,N_9905);
nor U10476 (N_10476,N_7430,N_8109);
and U10477 (N_10477,N_8388,N_7751);
and U10478 (N_10478,N_8537,N_9296);
nor U10479 (N_10479,N_9421,N_9988);
or U10480 (N_10480,N_9966,N_6431);
nand U10481 (N_10481,N_9056,N_8196);
and U10482 (N_10482,N_9387,N_9759);
nand U10483 (N_10483,N_5222,N_9663);
and U10484 (N_10484,N_5780,N_9616);
nand U10485 (N_10485,N_9541,N_6612);
or U10486 (N_10486,N_6490,N_5169);
and U10487 (N_10487,N_8453,N_9103);
nor U10488 (N_10488,N_6842,N_5269);
nor U10489 (N_10489,N_6774,N_8038);
or U10490 (N_10490,N_7980,N_9812);
and U10491 (N_10491,N_7434,N_8215);
nand U10492 (N_10492,N_7642,N_7101);
and U10493 (N_10493,N_5601,N_8311);
nand U10494 (N_10494,N_7047,N_8938);
and U10495 (N_10495,N_6087,N_6169);
nand U10496 (N_10496,N_6106,N_8717);
and U10497 (N_10497,N_7929,N_5822);
nor U10498 (N_10498,N_9008,N_9016);
or U10499 (N_10499,N_6166,N_6407);
and U10500 (N_10500,N_8467,N_9170);
nand U10501 (N_10501,N_7918,N_9562);
and U10502 (N_10502,N_9765,N_7306);
or U10503 (N_10503,N_9980,N_7016);
nand U10504 (N_10504,N_9739,N_7154);
nand U10505 (N_10505,N_6083,N_5595);
and U10506 (N_10506,N_6547,N_8542);
or U10507 (N_10507,N_9522,N_5451);
or U10508 (N_10508,N_8649,N_7415);
nor U10509 (N_10509,N_9834,N_8574);
nor U10510 (N_10510,N_9591,N_5645);
nor U10511 (N_10511,N_5365,N_5066);
or U10512 (N_10512,N_5998,N_9459);
nor U10513 (N_10513,N_5686,N_9178);
and U10514 (N_10514,N_5922,N_7005);
nand U10515 (N_10515,N_5284,N_8168);
nor U10516 (N_10516,N_5255,N_7111);
nand U10517 (N_10517,N_6419,N_7845);
and U10518 (N_10518,N_9515,N_5152);
nor U10519 (N_10519,N_9064,N_6011);
nand U10520 (N_10520,N_9237,N_5901);
or U10521 (N_10521,N_7290,N_6938);
and U10522 (N_10522,N_6355,N_8689);
nor U10523 (N_10523,N_6108,N_5249);
nand U10524 (N_10524,N_5299,N_8694);
nor U10525 (N_10525,N_5904,N_5092);
and U10526 (N_10526,N_6965,N_9848);
or U10527 (N_10527,N_7906,N_8583);
nor U10528 (N_10528,N_6926,N_5748);
nand U10529 (N_10529,N_6519,N_9559);
nor U10530 (N_10530,N_8979,N_9872);
and U10531 (N_10531,N_5570,N_5149);
and U10532 (N_10532,N_5816,N_8536);
and U10533 (N_10533,N_6228,N_6855);
nand U10534 (N_10534,N_6505,N_9225);
nor U10535 (N_10535,N_7879,N_9180);
nor U10536 (N_10536,N_5199,N_7599);
and U10537 (N_10537,N_7417,N_9967);
and U10538 (N_10538,N_7042,N_9389);
nand U10539 (N_10539,N_9360,N_7541);
nand U10540 (N_10540,N_6454,N_7805);
or U10541 (N_10541,N_5610,N_8515);
or U10542 (N_10542,N_7456,N_9143);
nand U10543 (N_10543,N_9586,N_9698);
nor U10544 (N_10544,N_5765,N_7378);
nor U10545 (N_10545,N_8796,N_9719);
or U10546 (N_10546,N_7011,N_7195);
and U10547 (N_10547,N_9245,N_7232);
or U10548 (N_10548,N_6644,N_9316);
or U10549 (N_10549,N_7332,N_5396);
and U10550 (N_10550,N_8850,N_6063);
nor U10551 (N_10551,N_9821,N_5431);
nand U10552 (N_10552,N_5994,N_5778);
nor U10553 (N_10553,N_7930,N_9236);
nand U10554 (N_10554,N_5317,N_5878);
nor U10555 (N_10555,N_5506,N_5692);
xor U10556 (N_10556,N_5139,N_8834);
or U10557 (N_10557,N_9254,N_5586);
or U10558 (N_10558,N_8539,N_7764);
and U10559 (N_10559,N_9140,N_5181);
nor U10560 (N_10560,N_7802,N_9802);
nor U10561 (N_10561,N_9753,N_8123);
nor U10562 (N_10562,N_7572,N_9881);
and U10563 (N_10563,N_5710,N_9264);
or U10564 (N_10564,N_8335,N_6561);
and U10565 (N_10565,N_9918,N_7575);
nor U10566 (N_10566,N_5051,N_8788);
or U10567 (N_10567,N_5560,N_9141);
or U10568 (N_10568,N_5859,N_6943);
or U10569 (N_10569,N_7780,N_7466);
xor U10570 (N_10570,N_9673,N_6482);
nand U10571 (N_10571,N_5929,N_5599);
or U10572 (N_10572,N_7648,N_5078);
and U10573 (N_10573,N_8731,N_8584);
and U10574 (N_10574,N_8653,N_5952);
nor U10575 (N_10575,N_9346,N_7311);
and U10576 (N_10576,N_5236,N_9472);
or U10577 (N_10577,N_6074,N_6102);
nor U10578 (N_10578,N_9022,N_9133);
nor U10579 (N_10579,N_6840,N_8290);
nand U10580 (N_10580,N_7485,N_8025);
xor U10581 (N_10581,N_8037,N_7716);
nor U10582 (N_10582,N_9925,N_7600);
nand U10583 (N_10583,N_6168,N_7260);
or U10584 (N_10584,N_9692,N_6617);
nor U10585 (N_10585,N_9811,N_5190);
nand U10586 (N_10586,N_6057,N_9145);
and U10587 (N_10587,N_9911,N_9007);
xnor U10588 (N_10588,N_8177,N_5184);
nor U10589 (N_10589,N_5465,N_9002);
nor U10590 (N_10590,N_7908,N_9091);
and U10591 (N_10591,N_6892,N_8534);
nand U10592 (N_10592,N_9961,N_9374);
xor U10593 (N_10593,N_7532,N_9537);
nor U10594 (N_10594,N_9824,N_7411);
nand U10595 (N_10595,N_8050,N_5819);
and U10596 (N_10596,N_9050,N_8945);
and U10597 (N_10597,N_8316,N_5781);
nor U10598 (N_10598,N_9363,N_7784);
or U10599 (N_10599,N_6553,N_5523);
nor U10600 (N_10600,N_9115,N_5943);
and U10601 (N_10601,N_9340,N_5024);
nand U10602 (N_10602,N_6722,N_5371);
or U10603 (N_10603,N_8896,N_7488);
nand U10604 (N_10604,N_8243,N_5360);
or U10605 (N_10605,N_9820,N_6065);
nand U10606 (N_10606,N_9754,N_7659);
nor U10607 (N_10607,N_8477,N_7270);
nand U10608 (N_10608,N_7838,N_6252);
xnor U10609 (N_10609,N_7834,N_5986);
and U10610 (N_10610,N_5696,N_6730);
or U10611 (N_10611,N_9806,N_8886);
nand U10612 (N_10612,N_9694,N_5336);
nor U10613 (N_10613,N_6934,N_9938);
nand U10614 (N_10614,N_9726,N_5028);
nand U10615 (N_10615,N_7437,N_7883);
or U10616 (N_10616,N_8613,N_8264);
and U10617 (N_10617,N_6013,N_9267);
or U10618 (N_10618,N_8854,N_9595);
and U10619 (N_10619,N_7507,N_7889);
or U10620 (N_10620,N_7956,N_6781);
nand U10621 (N_10621,N_5807,N_8590);
and U10622 (N_10622,N_8119,N_6788);
nand U10623 (N_10623,N_7610,N_9158);
nor U10624 (N_10624,N_7896,N_8132);
or U10625 (N_10625,N_7303,N_7268);
nor U10626 (N_10626,N_6770,N_9695);
xor U10627 (N_10627,N_7944,N_7256);
nor U10628 (N_10628,N_7873,N_5700);
and U10629 (N_10629,N_7844,N_9017);
and U10630 (N_10630,N_6800,N_9882);
nand U10631 (N_10631,N_6997,N_8310);
and U10632 (N_10632,N_8709,N_5292);
nand U10633 (N_10633,N_6299,N_9313);
nor U10634 (N_10634,N_8210,N_8222);
xnor U10635 (N_10635,N_9204,N_5455);
and U10636 (N_10636,N_7150,N_9262);
and U10637 (N_10637,N_7846,N_6461);
and U10638 (N_10638,N_6554,N_9399);
nor U10639 (N_10639,N_6568,N_7609);
and U10640 (N_10640,N_9489,N_8540);
nor U10641 (N_10641,N_6570,N_5991);
or U10642 (N_10642,N_6192,N_8005);
and U10643 (N_10643,N_8856,N_7583);
or U10644 (N_10644,N_6806,N_7945);
or U10645 (N_10645,N_6297,N_5080);
nand U10646 (N_10646,N_7903,N_5749);
or U10647 (N_10647,N_5305,N_8267);
nand U10648 (N_10648,N_8704,N_9442);
nor U10649 (N_10649,N_7854,N_6263);
and U10650 (N_10650,N_6070,N_5176);
and U10651 (N_10651,N_6305,N_9420);
nand U10652 (N_10652,N_5831,N_8949);
nand U10653 (N_10653,N_5187,N_6264);
or U10654 (N_10654,N_5641,N_9154);
nand U10655 (N_10655,N_8393,N_6145);
and U10656 (N_10656,N_9132,N_8570);
nand U10657 (N_10657,N_7072,N_8454);
nor U10658 (N_10658,N_6746,N_5794);
nand U10659 (N_10659,N_8851,N_9390);
nor U10660 (N_10660,N_7928,N_7773);
or U10661 (N_10661,N_7979,N_8897);
nor U10662 (N_10662,N_6785,N_9618);
or U10663 (N_10663,N_9998,N_7463);
nand U10664 (N_10664,N_6964,N_7292);
nand U10665 (N_10665,N_6448,N_7723);
nor U10666 (N_10666,N_5653,N_9377);
nand U10667 (N_10667,N_5084,N_9874);
nand U10668 (N_10668,N_7060,N_9298);
nand U10669 (N_10669,N_9315,N_9884);
nand U10670 (N_10670,N_6067,N_7948);
nand U10671 (N_10671,N_9150,N_6111);
and U10672 (N_10672,N_8270,N_5606);
nor U10673 (N_10673,N_5755,N_6947);
nand U10674 (N_10674,N_8361,N_6092);
or U10675 (N_10675,N_5244,N_5646);
nor U10676 (N_10676,N_8852,N_6194);
nand U10677 (N_10677,N_9770,N_9764);
nand U10678 (N_10678,N_8678,N_7116);
nor U10679 (N_10679,N_9321,N_9112);
or U10680 (N_10680,N_6239,N_6161);
nand U10681 (N_10681,N_5499,N_6748);
nor U10682 (N_10682,N_6900,N_5565);
or U10683 (N_10683,N_9453,N_6226);
and U10684 (N_10684,N_8873,N_6632);
or U10685 (N_10685,N_9379,N_7054);
or U10686 (N_10686,N_6173,N_5918);
or U10687 (N_10687,N_5023,N_7752);
nor U10688 (N_10688,N_7584,N_9813);
nor U10689 (N_10689,N_8186,N_8595);
nor U10690 (N_10690,N_6585,N_8076);
nand U10691 (N_10691,N_6631,N_8994);
and U10692 (N_10692,N_7941,N_9660);
xor U10693 (N_10693,N_7741,N_7949);
nor U10694 (N_10694,N_8211,N_6162);
and U10695 (N_10695,N_5507,N_5763);
or U10696 (N_10696,N_7112,N_9659);
and U10697 (N_10697,N_6188,N_7198);
nor U10698 (N_10698,N_5178,N_8966);
and U10699 (N_10699,N_9707,N_7258);
nand U10700 (N_10700,N_5034,N_9047);
nand U10701 (N_10701,N_6127,N_6587);
or U10702 (N_10702,N_5903,N_8843);
xor U10703 (N_10703,N_7678,N_8964);
and U10704 (N_10704,N_7793,N_7068);
and U10705 (N_10705,N_7749,N_8087);
and U10706 (N_10706,N_6346,N_7424);
or U10707 (N_10707,N_9441,N_5457);
or U10708 (N_10708,N_6405,N_5566);
or U10709 (N_10709,N_9053,N_9949);
nand U10710 (N_10710,N_5734,N_8718);
and U10711 (N_10711,N_9386,N_9857);
and U10712 (N_10712,N_6816,N_6725);
nand U10713 (N_10713,N_6694,N_8737);
nor U10714 (N_10714,N_8497,N_5312);
or U10715 (N_10715,N_8456,N_9720);
nor U10716 (N_10716,N_7344,N_9944);
nand U10717 (N_10717,N_7376,N_5243);
and U10718 (N_10718,N_7277,N_7446);
or U10719 (N_10719,N_6752,N_5910);
nand U10720 (N_10720,N_7729,N_6432);
and U10721 (N_10721,N_8754,N_9815);
nand U10722 (N_10722,N_8449,N_8842);
and U10723 (N_10723,N_6849,N_7656);
nor U10724 (N_10724,N_6659,N_9974);
nand U10725 (N_10725,N_7057,N_5131);
nand U10726 (N_10726,N_9873,N_9614);
or U10727 (N_10727,N_6693,N_6185);
and U10728 (N_10728,N_7581,N_5691);
and U10729 (N_10729,N_5492,N_5517);
and U10730 (N_10730,N_5966,N_9403);
nor U10731 (N_10731,N_8375,N_6804);
or U10732 (N_10732,N_7579,N_6864);
nand U10733 (N_10733,N_6373,N_7921);
nand U10734 (N_10734,N_8870,N_8925);
nor U10735 (N_10735,N_9994,N_8572);
or U10736 (N_10736,N_8166,N_5395);
and U10737 (N_10737,N_6686,N_5698);
or U10738 (N_10738,N_7080,N_8350);
nand U10739 (N_10739,N_9903,N_5825);
or U10740 (N_10740,N_5533,N_7370);
and U10741 (N_10741,N_8162,N_7251);
nor U10742 (N_10742,N_8478,N_5218);
or U10743 (N_10743,N_5627,N_6700);
and U10744 (N_10744,N_8491,N_6582);
nand U10745 (N_10745,N_5689,N_9320);
and U10746 (N_10746,N_7501,N_8976);
nand U10747 (N_10747,N_8713,N_8876);
and U10748 (N_10748,N_9427,N_8880);
and U10749 (N_10749,N_8262,N_7544);
and U10750 (N_10750,N_6029,N_6531);
and U10751 (N_10751,N_7339,N_5192);
or U10752 (N_10752,N_7210,N_7243);
nand U10753 (N_10753,N_7155,N_7620);
or U10754 (N_10754,N_7273,N_6425);
nor U10755 (N_10755,N_8780,N_5123);
nand U10756 (N_10756,N_8760,N_5563);
and U10757 (N_10757,N_8823,N_7747);
nand U10758 (N_10758,N_9040,N_8307);
or U10759 (N_10759,N_7066,N_8145);
and U10760 (N_10760,N_8508,N_9490);
or U10761 (N_10761,N_8008,N_9511);
nand U10762 (N_10762,N_9831,N_9287);
and U10763 (N_10763,N_6717,N_5477);
nor U10764 (N_10764,N_8160,N_5870);
and U10765 (N_10765,N_5154,N_7069);
or U10766 (N_10766,N_6916,N_5743);
or U10767 (N_10767,N_5707,N_5727);
nand U10768 (N_10768,N_9783,N_5614);
xnor U10769 (N_10769,N_7162,N_7853);
or U10770 (N_10770,N_7158,N_8192);
nor U10771 (N_10771,N_5682,N_9677);
nand U10772 (N_10772,N_8460,N_9639);
and U10773 (N_10773,N_5397,N_7136);
or U10774 (N_10774,N_9529,N_9335);
nand U10775 (N_10775,N_6262,N_8652);
or U10776 (N_10776,N_6805,N_6684);
and U10777 (N_10777,N_8355,N_5311);
and U10778 (N_10778,N_5136,N_7603);
and U10779 (N_10779,N_5804,N_7563);
nor U10780 (N_10780,N_9876,N_8202);
or U10781 (N_10781,N_8868,N_9730);
or U10782 (N_10782,N_5924,N_6290);
nand U10783 (N_10783,N_6624,N_9167);
nand U10784 (N_10784,N_6034,N_7015);
or U10785 (N_10785,N_6890,N_8706);
or U10786 (N_10786,N_5281,N_8909);
or U10787 (N_10787,N_7216,N_7519);
nand U10788 (N_10788,N_6539,N_5932);
nand U10789 (N_10789,N_8667,N_6003);
and U10790 (N_10790,N_9637,N_6508);
nor U10791 (N_10791,N_9048,N_6812);
and U10792 (N_10792,N_7967,N_8234);
and U10793 (N_10793,N_9202,N_7173);
or U10794 (N_10794,N_5348,N_5326);
or U10795 (N_10795,N_9587,N_5103);
or U10796 (N_10796,N_5402,N_5543);
and U10797 (N_10797,N_7984,N_8349);
and U10798 (N_10798,N_6457,N_9186);
nor U10799 (N_10799,N_6015,N_7255);
or U10800 (N_10800,N_7556,N_6773);
nand U10801 (N_10801,N_7665,N_7859);
or U10802 (N_10802,N_9638,N_9916);
or U10803 (N_10803,N_7619,N_5297);
and U10804 (N_10804,N_5363,N_6271);
or U10805 (N_10805,N_7688,N_7489);
nand U10806 (N_10806,N_6100,N_7451);
nor U10807 (N_10807,N_5278,N_8191);
nand U10808 (N_10808,N_5045,N_5694);
or U10809 (N_10809,N_5515,N_6980);
nor U10810 (N_10810,N_5379,N_5753);
or U10811 (N_10811,N_7338,N_6595);
nand U10812 (N_10812,N_6711,N_8217);
nor U10813 (N_10813,N_9709,N_6747);
nor U10814 (N_10814,N_5899,N_5981);
or U10815 (N_10815,N_8013,N_7818);
or U10816 (N_10816,N_5331,N_5597);
and U10817 (N_10817,N_9628,N_6973);
nand U10818 (N_10818,N_7577,N_8636);
or U10819 (N_10819,N_8011,N_6886);
nand U10820 (N_10820,N_5920,N_7901);
or U10821 (N_10821,N_5248,N_8178);
nand U10822 (N_10822,N_7970,N_5386);
nor U10823 (N_10823,N_7091,N_8630);
and U10824 (N_10824,N_5438,N_6466);
nor U10825 (N_10825,N_8034,N_7791);
or U10826 (N_10826,N_7383,N_6368);
nor U10827 (N_10827,N_6615,N_6082);
nand U10828 (N_10828,N_7467,N_6000);
xor U10829 (N_10829,N_5179,N_8860);
nor U10830 (N_10830,N_5195,N_7207);
or U10831 (N_10831,N_8684,N_8471);
and U10832 (N_10832,N_9110,N_6782);
nor U10833 (N_10833,N_6261,N_5951);
and U10834 (N_10834,N_8027,N_6238);
nand U10835 (N_10835,N_5126,N_8026);
nand U10836 (N_10836,N_9997,N_5061);
and U10837 (N_10837,N_5893,N_8184);
or U10838 (N_10838,N_5607,N_7159);
nand U10839 (N_10839,N_7756,N_8839);
nor U10840 (N_10840,N_9500,N_8965);
nand U10841 (N_10841,N_5775,N_7397);
or U10842 (N_10842,N_6033,N_5052);
and U10843 (N_10843,N_6961,N_6225);
or U10844 (N_10844,N_7759,N_9036);
nand U10845 (N_10845,N_9307,N_9187);
nor U10846 (N_10846,N_7396,N_6224);
nor U10847 (N_10847,N_6592,N_6933);
and U10848 (N_10848,N_5097,N_5879);
or U10849 (N_10849,N_5673,N_9382);
or U10850 (N_10850,N_8783,N_6215);
or U10851 (N_10851,N_8238,N_7635);
nand U10852 (N_10852,N_8939,N_6663);
and U10853 (N_10853,N_6378,N_7799);
and U10854 (N_10854,N_6163,N_7513);
or U10855 (N_10855,N_7736,N_7529);
nor U10856 (N_10856,N_8223,N_8266);
or U10857 (N_10857,N_9708,N_5947);
and U10858 (N_10858,N_5340,N_8670);
nor U10859 (N_10859,N_9120,N_8579);
nand U10860 (N_10860,N_5046,N_9394);
nor U10861 (N_10861,N_7786,N_5849);
nor U10862 (N_10862,N_8414,N_7654);
and U10863 (N_10863,N_5385,N_9836);
or U10864 (N_10864,N_7491,N_5373);
and U10865 (N_10865,N_8835,N_6843);
nand U10866 (N_10866,N_8898,N_9455);
nand U10867 (N_10867,N_5198,N_8521);
nand U10868 (N_10868,N_5811,N_9658);
or U10869 (N_10869,N_6891,N_6206);
or U10870 (N_10870,N_6362,N_8664);
nand U10871 (N_10871,N_9714,N_6878);
xor U10872 (N_10872,N_6674,N_8336);
nand U10873 (N_10873,N_5806,N_6367);
nor U10874 (N_10874,N_5090,N_6662);
nor U10875 (N_10875,N_9517,N_9005);
and U10876 (N_10876,N_8418,N_8483);
and U10877 (N_10877,N_6360,N_5074);
and U10878 (N_10878,N_7986,N_6104);
and U10879 (N_10879,N_9156,N_9396);
nand U10880 (N_10880,N_8035,N_6756);
nor U10881 (N_10881,N_5839,N_5235);
or U10882 (N_10882,N_6402,N_8494);
nand U10883 (N_10883,N_9062,N_9011);
nand U10884 (N_10884,N_9108,N_8826);
and U10885 (N_10885,N_9311,N_6174);
or U10886 (N_10886,N_7038,N_7757);
nor U10887 (N_10887,N_5056,N_8807);
nor U10888 (N_10888,N_9226,N_5488);
and U10889 (N_10889,N_5463,N_5260);
and U10890 (N_10890,N_5349,N_8606);
or U10891 (N_10891,N_9633,N_5130);
nor U10892 (N_10892,N_6734,N_9135);
or U10893 (N_10893,N_5841,N_8920);
and U10894 (N_10894,N_9272,N_9482);
nand U10895 (N_10895,N_5196,N_8072);
nor U10896 (N_10896,N_7346,N_6323);
nor U10897 (N_10897,N_7169,N_6436);
xor U10898 (N_10898,N_9886,N_6826);
nor U10899 (N_10899,N_6516,N_8565);
or U10900 (N_10900,N_7143,N_8874);
nand U10901 (N_10901,N_9835,N_5632);
and U10902 (N_10902,N_8940,N_9952);
nand U10903 (N_10903,N_5838,N_6338);
nor U10904 (N_10904,N_9398,N_9705);
or U10905 (N_10905,N_7758,N_5654);
and U10906 (N_10906,N_9034,N_9842);
nor U10907 (N_10907,N_8289,N_7618);
nand U10908 (N_10908,N_6498,N_5940);
nor U10909 (N_10909,N_7849,N_6007);
xor U10910 (N_10910,N_7063,N_6863);
and U10911 (N_10911,N_8148,N_7202);
nand U10912 (N_10912,N_5448,N_7616);
nand U10913 (N_10913,N_6504,N_5339);
nand U10914 (N_10914,N_7335,N_9240);
nand U10915 (N_10915,N_8877,N_9727);
and U10916 (N_10916,N_5369,N_5193);
nand U10917 (N_10917,N_8543,N_8597);
or U10918 (N_10918,N_5383,N_8318);
and U10919 (N_10919,N_5612,N_7735);
and U10920 (N_10920,N_9285,N_5364);
nand U10921 (N_10921,N_9457,N_9067);
or U10922 (N_10922,N_6618,N_5521);
xor U10923 (N_10923,N_6576,N_8069);
nor U10924 (N_10924,N_8904,N_5014);
or U10925 (N_10925,N_5121,N_7018);
nor U10926 (N_10926,N_9045,N_7316);
or U10927 (N_10927,N_7807,N_6841);
xor U10928 (N_10928,N_8657,N_5995);
nor U10929 (N_10929,N_9194,N_9114);
nand U10930 (N_10930,N_5917,N_6784);
and U10931 (N_10931,N_8988,N_6324);
and U10932 (N_10932,N_5848,N_5576);
or U10933 (N_10933,N_9935,N_6715);
nor U10934 (N_10934,N_8549,N_6014);
or U10935 (N_10935,N_7525,N_7558);
nand U10936 (N_10936,N_5826,N_9641);
and U10937 (N_10937,N_7445,N_7013);
or U10938 (N_10938,N_8358,N_9798);
nand U10939 (N_10939,N_8053,N_8319);
or U10940 (N_10940,N_5228,N_7989);
nand U10941 (N_10941,N_9169,N_5912);
nor U10942 (N_10942,N_8009,N_6430);
nand U10943 (N_10943,N_7870,N_5988);
nand U10944 (N_10944,N_6991,N_9230);
nor U10945 (N_10945,N_9116,N_8102);
nor U10946 (N_10946,N_7923,N_9546);
or U10947 (N_10947,N_6089,N_9757);
or U10948 (N_10948,N_7099,N_6643);
or U10949 (N_10949,N_7081,N_8167);
xnor U10950 (N_10950,N_7495,N_7442);
and U10951 (N_10951,N_9896,N_7356);
and U10952 (N_10952,N_9973,N_5323);
nor U10953 (N_10953,N_7932,N_6019);
or U10954 (N_10954,N_6337,N_9118);
nand U10955 (N_10955,N_5063,N_7776);
nand U10956 (N_10956,N_6394,N_7598);
nor U10957 (N_10957,N_9875,N_6253);
or U10958 (N_10958,N_6599,N_8193);
and U10959 (N_10959,N_7982,N_7117);
or U10960 (N_10960,N_9082,N_7611);
or U10961 (N_10961,N_7969,N_7301);
nor U10962 (N_10962,N_5587,N_5462);
nor U10963 (N_10963,N_8075,N_6529);
and U10964 (N_10964,N_9549,N_6446);
and U10965 (N_10965,N_6335,N_6331);
nor U10966 (N_10966,N_9792,N_7669);
nor U10967 (N_10967,N_5608,N_8055);
and U10968 (N_10968,N_8864,N_8012);
nand U10969 (N_10969,N_9250,N_5172);
or U10970 (N_10970,N_9662,N_6986);
and U10971 (N_10971,N_5851,N_9926);
or U10972 (N_10972,N_5008,N_9712);
or U10973 (N_10973,N_8271,N_9909);
nand U10974 (N_10974,N_5409,N_8520);
or U10975 (N_10975,N_7589,N_8545);
and U10976 (N_10976,N_8430,N_9629);
nor U10977 (N_10977,N_6823,N_9093);
or U10978 (N_10978,N_5401,N_8095);
xor U10979 (N_10979,N_9776,N_8984);
or U10980 (N_10980,N_6625,N_7500);
or U10981 (N_10981,N_7149,N_8396);
nand U10982 (N_10982,N_5680,N_9134);
and U10983 (N_10983,N_8492,N_8139);
nand U10984 (N_10984,N_6777,N_7860);
nor U10985 (N_10985,N_6118,N_5937);
nand U10986 (N_10986,N_9477,N_7156);
nand U10987 (N_10987,N_8263,N_8284);
nor U10988 (N_10988,N_7740,N_5147);
or U10989 (N_10989,N_6032,N_6295);
nor U10990 (N_10990,N_6291,N_5256);
or U10991 (N_10991,N_6197,N_6037);
nand U10992 (N_10992,N_8806,N_8914);
nor U10993 (N_10993,N_5035,N_6935);
or U10994 (N_10994,N_9704,N_6819);
and U10995 (N_10995,N_9255,N_7992);
nor U10996 (N_10996,N_9084,N_7523);
nor U10997 (N_10997,N_9488,N_9171);
nor U10998 (N_10998,N_9407,N_6153);
nor U10999 (N_10999,N_8764,N_6349);
or U11000 (N_11000,N_8383,N_9009);
or U11001 (N_11001,N_6844,N_6705);
nand U11002 (N_11002,N_9405,N_6626);
nor U11003 (N_11003,N_9355,N_7891);
and U11004 (N_11004,N_8524,N_6672);
xnor U11005 (N_11005,N_6381,N_6536);
or U11006 (N_11006,N_6212,N_5580);
and U11007 (N_11007,N_8751,N_6714);
and U11008 (N_11008,N_5182,N_6069);
nor U11009 (N_11009,N_6803,N_5062);
nand U11010 (N_11010,N_6620,N_5992);
and U11011 (N_11011,N_7083,N_7718);
nor U11012 (N_11012,N_5863,N_9246);
and U11013 (N_11013,N_7977,N_8086);
nand U11014 (N_11014,N_5997,N_7145);
and U11015 (N_11015,N_7278,N_8397);
nor U11016 (N_11016,N_6939,N_6332);
and U11017 (N_11017,N_8098,N_7074);
and U11018 (N_11018,N_8171,N_5502);
or U11019 (N_11019,N_7226,N_5472);
nor U11020 (N_11020,N_5688,N_6603);
and U11021 (N_11021,N_7836,N_6357);
xnor U11022 (N_11022,N_6358,N_6796);
nand U11023 (N_11023,N_8911,N_8567);
nor U11024 (N_11024,N_8802,N_8546);
nor U11025 (N_11025,N_7924,N_6303);
nand U11026 (N_11026,N_9890,N_9483);
or U11027 (N_11027,N_6707,N_5846);
nor U11028 (N_11028,N_5424,N_8743);
nand U11029 (N_11029,N_7293,N_8849);
or U11030 (N_11030,N_9085,N_7936);
and U11031 (N_11031,N_7320,N_6126);
nand U11032 (N_11032,N_9092,N_5527);
nand U11033 (N_11033,N_9676,N_5735);
and U11034 (N_11034,N_9852,N_5999);
nand U11035 (N_11035,N_5530,N_8133);
nand U11036 (N_11036,N_5664,N_6753);
nand U11037 (N_11037,N_5723,N_5075);
nand U11038 (N_11038,N_6330,N_5895);
or U11039 (N_11039,N_8778,N_8321);
nand U11040 (N_11040,N_9767,N_7045);
or U11041 (N_11041,N_7567,N_6911);
nand U11042 (N_11042,N_7453,N_9270);
nor U11043 (N_11043,N_6656,N_8131);
nor U11044 (N_11044,N_6158,N_8782);
nand U11045 (N_11045,N_6101,N_7677);
or U11046 (N_11046,N_5175,N_8247);
or U11047 (N_11047,N_8544,N_8447);
nand U11048 (N_11048,N_8960,N_5231);
nand U11049 (N_11049,N_5668,N_9424);
or U11050 (N_11050,N_5483,N_8931);
or U11051 (N_11051,N_5643,N_9858);
nor U11052 (N_11052,N_8197,N_7464);
and U11053 (N_11053,N_6175,N_6904);
nand U11054 (N_11054,N_5695,N_5372);
nor U11055 (N_11055,N_8328,N_9070);
nor U11056 (N_11056,N_5320,N_6597);
nand U11057 (N_11057,N_7206,N_6580);
and U11058 (N_11058,N_6956,N_9208);
xnor U11059 (N_11059,N_8658,N_6135);
xor U11060 (N_11060,N_5733,N_8564);
nor U11061 (N_11061,N_7161,N_6838);
nor U11062 (N_11062,N_6410,N_8043);
or U11063 (N_11063,N_8884,N_9342);
xnor U11064 (N_11064,N_8276,N_9383);
nor U11065 (N_11065,N_9548,N_8504);
nand U11066 (N_11066,N_9274,N_9605);
nor U11067 (N_11067,N_5079,N_8525);
and U11068 (N_11068,N_7053,N_9525);
or U11069 (N_11069,N_9619,N_9580);
or U11070 (N_11070,N_9286,N_6571);
nor U11071 (N_11071,N_7806,N_8114);
nand U11072 (N_11072,N_9176,N_6873);
and U11073 (N_11073,N_5572,N_8041);
nand U11074 (N_11074,N_5321,N_7093);
xnor U11075 (N_11075,N_8265,N_7363);
nand U11076 (N_11076,N_6049,N_6613);
and U11077 (N_11077,N_7034,N_8220);
and U11078 (N_11078,N_8021,N_7622);
nor U11079 (N_11079,N_5037,N_5820);
and U11080 (N_11080,N_8240,N_5791);
and U11081 (N_11081,N_9756,N_5221);
nand U11082 (N_11082,N_8555,N_7324);
nand U11083 (N_11083,N_8331,N_7211);
or U11084 (N_11084,N_6794,N_6879);
nand U11085 (N_11085,N_7864,N_8479);
or U11086 (N_11086,N_9197,N_5514);
nor U11087 (N_11087,N_7353,N_9615);
xnor U11088 (N_11088,N_8091,N_6370);
and U11089 (N_11089,N_9418,N_9228);
or U11090 (N_11090,N_9868,N_7077);
nand U11091 (N_11091,N_7874,N_9348);
and U11092 (N_11092,N_8274,N_7940);
nor U11093 (N_11093,N_5342,N_9039);
or U11094 (N_11094,N_8074,N_6017);
nand U11095 (N_11095,N_8643,N_9649);
nor U11096 (N_11096,N_8334,N_9799);
nand U11097 (N_11097,N_8983,N_8146);
and U11098 (N_11098,N_5547,N_6914);
or U11099 (N_11099,N_8930,N_7902);
nand U11100 (N_11100,N_6302,N_9324);
and U11101 (N_11101,N_8626,N_9671);
xnor U11102 (N_11102,N_5413,N_6257);
nor U11103 (N_11103,N_8859,N_6095);
and U11104 (N_11104,N_5611,N_9865);
or U11105 (N_11105,N_6056,N_7682);
and U11106 (N_11106,N_7861,N_9281);
and U11107 (N_11107,N_6098,N_8827);
or U11108 (N_11108,N_8236,N_8627);
nor U11109 (N_11109,N_5128,N_5205);
and U11110 (N_11110,N_7259,N_8248);
nor U11111 (N_11111,N_7379,N_8297);
nand U11112 (N_11112,N_8872,N_5021);
nor U11113 (N_11113,N_9516,N_6530);
nand U11114 (N_11114,N_8681,N_7580);
nand U11115 (N_11115,N_7790,N_6121);
and U11116 (N_11116,N_7942,N_6848);
nand U11117 (N_11117,N_5876,N_7743);
and U11118 (N_11118,N_8282,N_7646);
and U11119 (N_11119,N_9947,N_6209);
and U11120 (N_11120,N_5519,N_5065);
or U11121 (N_11121,N_7493,N_6246);
or U11122 (N_11122,N_8517,N_9520);
xor U11123 (N_11123,N_8332,N_9907);
nor U11124 (N_11124,N_8933,N_9553);
nand U11125 (N_11125,N_9795,N_8781);
or U11126 (N_11126,N_7974,N_6421);
or U11127 (N_11127,N_6699,N_5855);
or U11128 (N_11128,N_7694,N_7555);
nor U11129 (N_11129,N_8963,N_7168);
nand U11130 (N_11130,N_5752,N_9510);
nor U11131 (N_11131,N_7297,N_7666);
nor U11132 (N_11132,N_5054,N_6703);
nand U11133 (N_11133,N_5890,N_6204);
nor U11134 (N_11134,N_5812,N_8039);
nand U11135 (N_11135,N_9892,N_6078);
nand U11136 (N_11136,N_7237,N_8405);
and U11137 (N_11137,N_5435,N_7785);
and U11138 (N_11138,N_6452,N_5866);
nor U11139 (N_11139,N_9031,N_8669);
and U11140 (N_11140,N_5202,N_7983);
nor U11141 (N_11141,N_6183,N_7405);
nor U11142 (N_11142,N_5793,N_8341);
and U11143 (N_11143,N_6502,N_7534);
nor U11144 (N_11144,N_8085,N_8906);
xor U11145 (N_11145,N_6451,N_8448);
xor U11146 (N_11146,N_5624,N_7958);
nand U11147 (N_11147,N_7176,N_7153);
and U11148 (N_11148,N_9381,N_5429);
xnor U11149 (N_11149,N_8324,N_7308);
nor U11150 (N_11150,N_5944,N_9430);
nor U11151 (N_11151,N_7981,N_6365);
and U11152 (N_11152,N_7321,N_7056);
nor U11153 (N_11153,N_8018,N_6895);
or U11154 (N_11154,N_5813,N_8296);
nor U11155 (N_11155,N_6422,N_8675);
or U11156 (N_11156,N_6396,N_8503);
nand U11157 (N_11157,N_5974,N_6506);
and U11158 (N_11158,N_9065,N_6959);
nor U11159 (N_11159,N_6755,N_6920);
and U11160 (N_11160,N_5344,N_6341);
or U11161 (N_11161,N_8729,N_8474);
nor U11162 (N_11162,N_5795,N_5459);
nand U11163 (N_11163,N_5758,N_6424);
nand U11164 (N_11164,N_8422,N_7472);
xnor U11165 (N_11165,N_5581,N_5495);
or U11166 (N_11166,N_5163,N_9428);
nand U11167 (N_11167,N_8825,N_8084);
nor U11168 (N_11168,N_8588,N_7300);
or U11169 (N_11169,N_9526,N_9772);
nor U11170 (N_11170,N_6315,N_7685);
nand U11171 (N_11171,N_7448,N_7126);
nand U11172 (N_11172,N_5247,N_7223);
and U11173 (N_11173,N_6623,N_8560);
or U11174 (N_11174,N_6186,N_8958);
nor U11175 (N_11175,N_6847,N_5486);
nand U11176 (N_11176,N_8978,N_8708);
nand U11177 (N_11177,N_9603,N_9599);
or U11178 (N_11178,N_6995,N_5629);
nand U11179 (N_11179,N_6386,N_6882);
and U11180 (N_11180,N_9263,N_8741);
nand U11181 (N_11181,N_6423,N_6690);
nand U11182 (N_11182,N_5690,N_9416);
nand U11183 (N_11183,N_9943,N_7391);
or U11184 (N_11184,N_9854,N_5291);
and U11185 (N_11185,N_6052,N_6909);
nor U11186 (N_11186,N_5625,N_8382);
and U11187 (N_11187,N_5889,N_5845);
nand U11188 (N_11188,N_9958,N_9651);
nand U11189 (N_11189,N_5022,N_9481);
or U11190 (N_11190,N_6309,N_9153);
or U11191 (N_11191,N_5783,N_8725);
nor U11192 (N_11192,N_5233,N_7291);
nand U11193 (N_11193,N_5434,N_7851);
nor U11194 (N_11194,N_8552,N_8721);
or U11195 (N_11195,N_5873,N_9762);
nor U11196 (N_11196,N_8093,N_9247);
nor U11197 (N_11197,N_9479,N_6312);
nor U11198 (N_11198,N_9536,N_9664);
nand U11199 (N_11199,N_7334,N_8905);
and U11200 (N_11200,N_5864,N_9075);
or U11201 (N_11201,N_8189,N_7439);
and U11202 (N_11202,N_8614,N_7208);
nand U11203 (N_11203,N_6702,N_8946);
and U11204 (N_11204,N_6353,N_5330);
nand U11205 (N_11205,N_6713,N_9098);
or U11206 (N_11206,N_9558,N_9013);
and U11207 (N_11207,N_5913,N_6897);
and U11208 (N_11208,N_7328,N_6793);
and U11209 (N_11209,N_9744,N_9414);
nand U11210 (N_11210,N_8608,N_7432);
or U11211 (N_11211,N_6649,N_7138);
nand U11212 (N_11212,N_6776,N_6071);
nand U11213 (N_11213,N_7661,N_9986);
nand U11214 (N_11214,N_7224,N_5473);
and U11215 (N_11215,N_9841,N_8291);
nand U11216 (N_11216,N_9763,N_7287);
nand U11217 (N_11217,N_9117,N_8246);
and U11218 (N_11218,N_6391,N_7863);
nor U11219 (N_11219,N_5358,N_8758);
nor U11220 (N_11220,N_6189,N_8813);
and U11221 (N_11221,N_6792,N_6247);
nand U11222 (N_11222,N_5549,N_8329);
or U11223 (N_11223,N_8990,N_5433);
nor U11224 (N_11224,N_6634,N_5239);
nand U11225 (N_11225,N_9243,N_5105);
or U11226 (N_11226,N_8734,N_8348);
and U11227 (N_11227,N_5705,N_5584);
and U11228 (N_11228,N_7626,N_7911);
nor U11229 (N_11229,N_6222,N_5842);
and U11230 (N_11230,N_7246,N_9788);
nand U11231 (N_11231,N_7135,N_8867);
and U11232 (N_11232,N_5471,N_7388);
nor U11233 (N_11233,N_5077,N_6219);
or U11234 (N_11234,N_8399,N_8352);
or U11235 (N_11235,N_9853,N_5258);
nor U11236 (N_11236,N_7996,N_8130);
nand U11237 (N_11237,N_8426,N_9411);
nor U11238 (N_11238,N_5257,N_7826);
nand U11239 (N_11239,N_9338,N_7127);
and U11240 (N_11240,N_5579,N_9329);
and U11241 (N_11241,N_8619,N_5091);
or U11242 (N_11242,N_6002,N_5058);
nand U11243 (N_11243,N_9094,N_6411);
or U11244 (N_11244,N_6081,N_8901);
xnor U11245 (N_11245,N_8028,N_7179);
and U11246 (N_11246,N_5030,N_9491);
xor U11247 (N_11247,N_6594,N_5837);
or U11248 (N_11248,N_6047,N_6172);
nand U11249 (N_11249,N_7797,N_9645);
or U11250 (N_11250,N_8682,N_8249);
nand U11251 (N_11251,N_8793,N_8862);
and U11252 (N_11252,N_7721,N_5025);
and U11253 (N_11253,N_7927,N_8429);
or U11254 (N_11254,N_9235,N_5990);
nand U11255 (N_11255,N_9366,N_9785);
and U11256 (N_11256,N_7115,N_5972);
or U11257 (N_11257,N_7594,N_9900);
or U11258 (N_11258,N_8007,N_8228);
nand U11259 (N_11259,N_7964,N_9165);
nand U11260 (N_11260,N_6827,N_7872);
or U11261 (N_11261,N_8720,N_5989);
and U11262 (N_11262,N_8003,N_9611);
and U11263 (N_11263,N_8216,N_9644);
nor U11264 (N_11264,N_5501,N_9060);
and U11265 (N_11265,N_5412,N_6460);
nand U11266 (N_11266,N_9352,N_8121);
xnor U11267 (N_11267,N_6280,N_8462);
or U11268 (N_11268,N_7538,N_9043);
or U11269 (N_11269,N_9732,N_5388);
or U11270 (N_11270,N_5009,N_8810);
nor U11271 (N_11271,N_9796,N_7390);
nor U11272 (N_11272,N_9044,N_5232);
nand U11273 (N_11273,N_7181,N_7071);
nor U11274 (N_11274,N_9330,N_8951);
nand U11275 (N_11275,N_7010,N_6975);
or U11276 (N_11276,N_6712,N_5450);
and U11277 (N_11277,N_8047,N_9581);
or U11278 (N_11278,N_8739,N_5005);
or U11279 (N_11279,N_9055,N_9373);
nor U11280 (N_11280,N_9550,N_8033);
or U11281 (N_11281,N_6954,N_8714);
and U11282 (N_11282,N_7003,N_5926);
and U11283 (N_11283,N_5333,N_7559);
or U11284 (N_11284,N_9996,N_9242);
nand U11285 (N_11285,N_5148,N_9960);
or U11286 (N_11286,N_5750,N_8308);
or U11287 (N_11287,N_6871,N_6921);
or U11288 (N_11288,N_8269,N_5534);
and U11289 (N_11289,N_9402,N_8024);
and U11290 (N_11290,N_6198,N_8194);
or U11291 (N_11291,N_8359,N_6275);
and U11292 (N_11292,N_7095,N_8861);
nor U11293 (N_11293,N_5032,N_9310);
nor U11294 (N_11294,N_7228,N_8671);
nand U11295 (N_11295,N_9670,N_9534);
or U11296 (N_11296,N_9895,N_8410);
and U11297 (N_11297,N_8812,N_6971);
nand U11298 (N_11298,N_8354,N_9327);
nand U11299 (N_11299,N_9295,N_8531);
and U11300 (N_11300,N_8693,N_9474);
nor U11301 (N_11301,N_6447,N_8482);
nor U11302 (N_11302,N_9552,N_9302);
or U11303 (N_11303,N_6376,N_7046);
nor U11304 (N_11304,N_5119,N_9932);
nor U11305 (N_11305,N_6359,N_8701);
and U11306 (N_11306,N_8942,N_7247);
nor U11307 (N_11307,N_6304,N_7227);
nand U11308 (N_11308,N_5016,N_8432);
nor U11309 (N_11309,N_5964,N_5982);
nand U11310 (N_11310,N_6345,N_5206);
and U11311 (N_11311,N_9078,N_8108);
nand U11312 (N_11312,N_7392,N_9322);
nor U11313 (N_11313,N_9494,N_9575);
nor U11314 (N_11314,N_6035,N_9122);
or U11315 (N_11315,N_8340,N_8113);
and U11316 (N_11316,N_5238,N_9174);
or U11317 (N_11317,N_6736,N_7009);
xor U11318 (N_11318,N_8486,N_7342);
and U11319 (N_11319,N_5745,N_9096);
nand U11320 (N_11320,N_5854,N_7913);
and U11321 (N_11321,N_5325,N_5491);
and U11322 (N_11322,N_8680,N_5279);
nand U11323 (N_11323,N_7244,N_5270);
and U11324 (N_11324,N_8065,N_9063);
and U11325 (N_11325,N_8157,N_7587);
and U11326 (N_11326,N_6682,N_8926);
nand U11327 (N_11327,N_6385,N_7178);
or U11328 (N_11328,N_9969,N_8629);
or U11329 (N_11329,N_8501,N_6828);
nor U11330 (N_11330,N_5425,N_5134);
and U11331 (N_11331,N_8690,N_5853);
or U11332 (N_11332,N_6025,N_7103);
and U11333 (N_11333,N_7438,N_6073);
nand U11334 (N_11334,N_9607,N_8235);
or U11335 (N_11335,N_6726,N_8705);
or U11336 (N_11336,N_9012,N_8875);
nor U11337 (N_11337,N_5484,N_7576);
or U11338 (N_11338,N_5880,N_5335);
nand U11339 (N_11339,N_5057,N_7885);
or U11340 (N_11340,N_6076,N_8237);
nor U11341 (N_11341,N_8688,N_8814);
nor U11342 (N_11342,N_8547,N_7774);
and U11343 (N_11343,N_8413,N_6697);
nor U11344 (N_11344,N_6988,N_9807);
nor U11345 (N_11345,N_9077,N_8586);
and U11346 (N_11346,N_6718,N_5894);
nor U11347 (N_11347,N_7664,N_6556);
nor U11348 (N_11348,N_9215,N_5338);
nor U11349 (N_11349,N_5081,N_9199);
nor U11350 (N_11350,N_6720,N_7771);
or U11351 (N_11351,N_6658,N_7280);
and U11352 (N_11352,N_6260,N_5356);
and U11353 (N_11353,N_6586,N_7715);
nor U11354 (N_11354,N_5357,N_8659);
nor U11355 (N_11355,N_8645,N_9722);
nor U11356 (N_11356,N_9823,N_5950);
nor U11357 (N_11357,N_6577,N_6044);
and U11358 (N_11358,N_7769,N_9415);
nor U11359 (N_11359,N_5318,N_7985);
nor U11360 (N_11360,N_9856,N_6998);
xnor U11361 (N_11361,N_6593,N_9191);
nor U11362 (N_11362,N_9404,N_7276);
nor U11363 (N_11363,N_5432,N_5665);
nand U11364 (N_11364,N_7763,N_8785);
nand U11365 (N_11365,N_8079,N_9261);
or U11366 (N_11366,N_9480,N_8554);
xor U11367 (N_11367,N_7183,N_7551);
and U11368 (N_11368,N_5146,N_6403);
nor U11369 (N_11369,N_6917,N_8700);
or U11370 (N_11370,N_9336,N_8779);
nand U11371 (N_11371,N_5504,N_8212);
nor U11372 (N_11372,N_7728,N_9241);
or U11373 (N_11373,N_9445,N_5452);
or U11374 (N_11374,N_7050,N_7025);
nor U11375 (N_11375,N_6130,N_8438);
or U11376 (N_11376,N_5230,N_5886);
and U11377 (N_11377,N_8672,N_5137);
nor U11378 (N_11378,N_8771,N_8278);
nor U11379 (N_11379,N_7033,N_9547);
xnor U11380 (N_11380,N_7073,N_8919);
and U11381 (N_11381,N_7655,N_9190);
nand U11382 (N_11382,N_5767,N_7707);
nand U11383 (N_11383,N_6555,N_5273);
nor U11384 (N_11384,N_8617,N_9871);
nand U11385 (N_11385,N_8665,N_9565);
and U11386 (N_11386,N_7355,N_7962);
nand U11387 (N_11387,N_6342,N_6548);
or U11388 (N_11388,N_7878,N_8803);
and U11389 (N_11389,N_8280,N_9206);
and U11390 (N_11390,N_6772,N_8281);
nand U11391 (N_11391,N_6167,N_9431);
or U11392 (N_11392,N_6627,N_7954);
or U11393 (N_11393,N_9684,N_9793);
or U11394 (N_11394,N_9685,N_7004);
nor U11395 (N_11395,N_6808,N_9590);
and U11396 (N_11396,N_9214,N_8924);
and U11397 (N_11397,N_5302,N_8373);
or U11398 (N_11398,N_9564,N_7811);
and U11399 (N_11399,N_9343,N_7543);
nand U11400 (N_11400,N_5721,N_6267);
nand U11401 (N_11401,N_7336,N_7469);
nand U11402 (N_11402,N_7965,N_9125);
nor U11403 (N_11403,N_6983,N_8756);
or U11404 (N_11404,N_5404,N_5183);
or U11405 (N_11405,N_8923,N_7546);
nor U11406 (N_11406,N_6589,N_5512);
nand U11407 (N_11407,N_9364,N_8890);
or U11408 (N_11408,N_5403,N_7027);
and U11409 (N_11409,N_5087,N_8514);
and U11410 (N_11410,N_7561,N_8469);
and U11411 (N_11411,N_8811,N_6813);
or U11412 (N_11412,N_7788,N_5662);
nor U11413 (N_11413,N_8830,N_8838);
nor U11414 (N_11414,N_7787,N_5909);
nand U11415 (N_11415,N_8275,N_5101);
nand U11416 (N_11416,N_9162,N_5637);
nor U11417 (N_11417,N_5511,N_9152);
and U11418 (N_11418,N_6259,N_5072);
nand U11419 (N_11419,N_5480,N_8558);
nand U11420 (N_11420,N_7535,N_9213);
or U11421 (N_11421,N_9406,N_8633);
and U11422 (N_11422,N_7809,N_5387);
or U11423 (N_11423,N_8551,N_6406);
and U11424 (N_11424,N_6336,N_5568);
or U11425 (N_11425,N_8962,N_9102);
nand U11426 (N_11426,N_5936,N_6542);
nand U11427 (N_11427,N_5102,N_9717);
nor U11428 (N_11428,N_5818,N_8061);
or U11429 (N_11429,N_9693,N_7134);
nor U11430 (N_11430,N_7732,N_7813);
nor U11431 (N_11431,N_5217,N_8161);
nor U11432 (N_11432,N_6646,N_8376);
or U11433 (N_11433,N_7030,N_5027);
or U11434 (N_11434,N_8412,N_7239);
nand U11435 (N_11435,N_8968,N_6500);
nor U11436 (N_11436,N_5774,N_7088);
and U11437 (N_11437,N_6314,N_7995);
and U11438 (N_11438,N_7426,N_6235);
nand U11439 (N_11439,N_9361,N_6018);
and U11440 (N_11440,N_6802,N_7804);
nand U11441 (N_11441,N_8362,N_5857);
nor U11442 (N_11442,N_5110,N_9375);
nand U11443 (N_11443,N_7697,N_9667);
or U11444 (N_11444,N_7043,N_7214);
nand U11445 (N_11445,N_5416,N_8357);
nand U11446 (N_11446,N_6578,N_6630);
or U11447 (N_11447,N_8591,N_9462);
and U11448 (N_11448,N_7139,N_9506);
or U11449 (N_11449,N_8155,N_7739);
nand U11450 (N_11450,N_5082,N_8251);
or U11451 (N_11451,N_9277,N_8124);
or U11452 (N_11452,N_9347,N_9787);
nor U11453 (N_11453,N_5191,N_7284);
and U11454 (N_11454,N_5562,N_7298);
nor U11455 (N_11455,N_7875,N_5261);
nor U11456 (N_11456,N_5914,N_6865);
or U11457 (N_11457,N_6907,N_5882);
nor U11458 (N_11458,N_7151,N_6870);
and U11459 (N_11459,N_7895,N_6866);
nand U11460 (N_11460,N_8142,N_6957);
nand U11461 (N_11461,N_6691,N_7926);
xor U11462 (N_11462,N_5031,N_8695);
nor U11463 (N_11463,N_6042,N_6850);
and U11464 (N_11464,N_8466,N_6503);
or U11465 (N_11465,N_5210,N_8561);
and U11466 (N_11466,N_9172,N_7880);
nor U11467 (N_11467,N_9929,N_7429);
and U11468 (N_11468,N_9080,N_5805);
and U11469 (N_11469,N_5604,N_9076);
nand U11470 (N_11470,N_8651,N_5868);
or U11471 (N_11471,N_6596,N_7633);
nand U11472 (N_11472,N_5623,N_7503);
and U11473 (N_11473,N_5535,N_7569);
nor U11474 (N_11474,N_6836,N_5185);
nor U11475 (N_11475,N_9648,N_6607);
or U11476 (N_11476,N_5298,N_9026);
or U11477 (N_11477,N_6852,N_8305);
nor U11478 (N_11478,N_6068,N_6480);
or U11479 (N_11479,N_7062,N_9613);
nand U11480 (N_11480,N_7843,N_7877);
and U11481 (N_11481,N_7692,N_9126);
and U11482 (N_11482,N_8755,N_6137);
or U11483 (N_11483,N_6048,N_9643);
nand U11484 (N_11484,N_5353,N_6369);
and U11485 (N_11485,N_5931,N_9345);
nand U11486 (N_11486,N_6993,N_5746);
and U11487 (N_11487,N_5209,N_8299);
or U11488 (N_11488,N_9185,N_9530);
nor U11489 (N_11489,N_8406,N_8749);
and U11490 (N_11490,N_9278,N_9193);
nand U11491 (N_11491,N_6740,N_7394);
or U11492 (N_11492,N_7730,N_6739);
or U11493 (N_11493,N_5897,N_6196);
or U11494 (N_11494,N_8772,N_9773);
or U11495 (N_11495,N_8556,N_7221);
nor U11496 (N_11496,N_9544,N_8106);
and U11497 (N_11497,N_5747,N_6832);
nand U11498 (N_11498,N_7386,N_6815);
nand U11499 (N_11499,N_5770,N_6758);
nor U11500 (N_11500,N_5728,N_5316);
or U11501 (N_11501,N_5790,N_6453);
and U11502 (N_11502,N_7354,N_7823);
nor U11503 (N_11503,N_5241,N_7288);
nor U11504 (N_11504,N_8644,N_5885);
nand U11505 (N_11505,N_6797,N_7691);
nor U11506 (N_11506,N_9257,N_8097);
nand U11507 (N_11507,N_9735,N_8676);
or U11508 (N_11508,N_5374,N_9314);
or U11509 (N_11509,N_6676,N_6598);
or U11510 (N_11510,N_9328,N_7422);
and U11511 (N_11511,N_7748,N_6340);
nor U11512 (N_11512,N_9503,N_5161);
nand U11513 (N_11513,N_5265,N_5546);
or U11514 (N_11514,N_5797,N_6704);
nand U11515 (N_11515,N_9492,N_8715);
and U11516 (N_11516,N_7357,N_8434);
or U11517 (N_11517,N_8488,N_8816);
or U11518 (N_11518,N_8421,N_7078);
and U11519 (N_11519,N_6654,N_7184);
and U11520 (N_11520,N_9585,N_5577);
nand U11521 (N_11521,N_5603,N_9372);
xnor U11522 (N_11522,N_7781,N_5532);
and U11523 (N_11523,N_6535,N_6666);
nor U11524 (N_11524,N_6526,N_9159);
or U11525 (N_11525,N_5946,N_9238);
or U11526 (N_11526,N_9439,N_6061);
or U11527 (N_11527,N_6440,N_7400);
or U11528 (N_11528,N_8165,N_8137);
and U11529 (N_11529,N_6528,N_8956);
or U11530 (N_11530,N_6005,N_7634);
nand U11531 (N_11531,N_5059,N_9863);
nor U11532 (N_11532,N_5226,N_7241);
or U11533 (N_11533,N_5706,N_6901);
and U11534 (N_11534,N_9451,N_7536);
and U11535 (N_11535,N_7031,N_8961);
or U11536 (N_11536,N_5605,N_8615);
or U11537 (N_11537,N_7454,N_8143);
nand U11538 (N_11538,N_5170,N_6471);
and U11539 (N_11539,N_5699,N_5382);
and U11540 (N_11540,N_9425,N_9729);
or U11541 (N_11541,N_9249,N_9177);
and U11542 (N_11542,N_8415,N_5539);
and U11543 (N_11543,N_6673,N_5262);
and U11544 (N_11544,N_6389,N_9450);
nor U11545 (N_11545,N_5725,N_9220);
nor U11546 (N_11546,N_7531,N_5542);
nor U11547 (N_11547,N_5135,N_6329);
xnor U11548 (N_11548,N_9731,N_5896);
nand U11549 (N_11549,N_8029,N_5303);
or U11550 (N_11550,N_7952,N_7578);
and U11551 (N_11551,N_6051,N_7142);
and U11552 (N_11552,N_6351,N_7452);
and U11553 (N_11553,N_6476,N_6562);
nor U11554 (N_11554,N_8424,N_6645);
nand U11555 (N_11555,N_7408,N_9024);
nor U11556 (N_11556,N_9010,N_9940);
and U11557 (N_11557,N_7317,N_5671);
xor U11558 (N_11558,N_6899,N_7085);
nor U11559 (N_11559,N_9568,N_5835);
nand U11560 (N_11560,N_8201,N_9317);
and U11561 (N_11561,N_5513,N_5900);
nor U11562 (N_11562,N_5245,N_9349);
or U11563 (N_11563,N_6112,N_9760);
or U11564 (N_11564,N_5916,N_7157);
nand U11565 (N_11565,N_5124,N_8337);
or U11566 (N_11566,N_9408,N_7186);
or U11567 (N_11567,N_7778,N_5167);
xnor U11568 (N_11568,N_8918,N_5718);
or U11569 (N_11569,N_8752,N_8832);
or U11570 (N_11570,N_9051,N_5224);
nand U11571 (N_11571,N_5093,N_8620);
and U11572 (N_11572,N_6371,N_7458);
and U11573 (N_11573,N_7573,N_9540);
nand U11574 (N_11574,N_5796,N_9576);
xnor U11575 (N_11575,N_9914,N_5223);
or U11576 (N_11576,N_8437,N_8364);
nand U11577 (N_11577,N_9470,N_8115);
and U11578 (N_11578,N_7670,N_5422);
and U11579 (N_11579,N_9357,N_6165);
nand U11580 (N_11580,N_8472,N_7419);
or U11581 (N_11581,N_5143,N_5709);
and U11582 (N_11582,N_6176,N_9280);
or U11583 (N_11583,N_9046,N_9822);
xor U11584 (N_11584,N_5616,N_7441);
and U11585 (N_11585,N_6105,N_5157);
and U11586 (N_11586,N_7435,N_7808);
nor U11587 (N_11587,N_7798,N_7087);
and U11588 (N_11588,N_9819,N_5784);
xnor U11589 (N_11589,N_7530,N_9020);
or U11590 (N_11590,N_6952,N_8049);
nand U11591 (N_11591,N_7461,N_6296);
or U11592 (N_11592,N_5337,N_9229);
nor U11593 (N_11593,N_9883,N_7407);
nand U11594 (N_11594,N_9306,N_5053);
nand U11595 (N_11595,N_9493,N_5617);
nand U11596 (N_11596,N_7512,N_8484);
or U11597 (N_11597,N_7777,N_6779);
xnor U11598 (N_11598,N_7898,N_6780);
nor U11599 (N_11599,N_7124,N_5583);
or U11600 (N_11600,N_7123,N_5661);
and U11601 (N_11601,N_6125,N_7064);
or U11602 (N_11602,N_6664,N_5327);
nand U11603 (N_11603,N_5836,N_6001);
xor U11604 (N_11604,N_6274,N_7065);
nand U11605 (N_11605,N_8726,N_6771);
nand U11606 (N_11606,N_5971,N_9300);
nor U11607 (N_11607,N_6867,N_6560);
and U11608 (N_11608,N_8023,N_6636);
and U11609 (N_11609,N_6898,N_8819);
nand U11610 (N_11610,N_7307,N_7067);
and U11611 (N_11611,N_5669,N_8847);
or U11612 (N_11612,N_8384,N_7947);
nand U11613 (N_11613,N_8724,N_6661);
nand U11614 (N_11614,N_8351,N_9556);
nand U11615 (N_11615,N_6728,N_9188);
and U11616 (N_11616,N_6564,N_6441);
nor U11617 (N_11617,N_9566,N_7444);
nor U11618 (N_11618,N_7262,N_6384);
or U11619 (N_11619,N_5875,N_5419);
nand U11620 (N_11620,N_8450,N_5380);
nor U11621 (N_11621,N_6606,N_9266);
nor U11622 (N_11622,N_6635,N_9097);
or U11623 (N_11623,N_7994,N_5487);
or U11624 (N_11624,N_6426,N_7282);
nand U11625 (N_11625,N_9542,N_5050);
and U11626 (N_11626,N_6534,N_9072);
and U11627 (N_11627,N_9089,N_5108);
or U11628 (N_11628,N_7428,N_8322);
nand U11629 (N_11629,N_9452,N_8006);
nor U11630 (N_11630,N_8301,N_6982);
or U11631 (N_11631,N_9681,N_9898);
nand U11632 (N_11632,N_7465,N_9332);
nand U11633 (N_11633,N_6581,N_9592);
nor U11634 (N_11634,N_7564,N_6244);
nand U11635 (N_11635,N_5843,N_7812);
nor U11636 (N_11636,N_6485,N_6488);
or U11637 (N_11637,N_7835,N_6880);
or U11638 (N_11638,N_5731,N_8789);
nor U11639 (N_11639,N_8808,N_7990);
nand U11640 (N_11640,N_8105,N_5824);
or U11641 (N_11641,N_9101,N_5559);
nand U11642 (N_11642,N_7939,N_5234);
and U11643 (N_11643,N_9839,N_6668);
and U11644 (N_11644,N_6854,N_5908);
and U11645 (N_11645,N_8490,N_8980);
nor U11646 (N_11646,N_5015,N_8128);
or U11647 (N_11647,N_6953,N_5378);
or U11648 (N_11648,N_8922,N_5554);
nor U11649 (N_11649,N_8763,N_6915);
and U11650 (N_11650,N_7403,N_6122);
nor U11651 (N_11651,N_9690,N_7526);
and U11652 (N_11652,N_8817,N_5766);
nor U11653 (N_11653,N_5978,N_5280);
and U11654 (N_11654,N_5803,N_6399);
or U11655 (N_11655,N_7909,N_7978);
nand U11656 (N_11656,N_7699,N_9888);
nor U11657 (N_11657,N_8175,N_8046);
nand U11658 (N_11658,N_9184,N_6513);
or U11659 (N_11659,N_9083,N_7684);
nand U11660 (N_11660,N_6170,N_7511);
or U11661 (N_11661,N_8742,N_7613);
nor U11662 (N_11662,N_7494,N_8054);
nand U11663 (N_11663,N_9496,N_9860);
and U11664 (N_11664,N_8801,N_9423);
nand U11665 (N_11665,N_9545,N_9059);
nand U11666 (N_11666,N_7250,N_9400);
or U11667 (N_11667,N_5194,N_5925);
and U11668 (N_11668,N_8844,N_8592);
nand U11669 (N_11669,N_9869,N_5400);
nor U11670 (N_11670,N_9899,N_8900);
nand U11671 (N_11671,N_9661,N_7668);
and U11672 (N_11672,N_9049,N_6851);
xor U11673 (N_11673,N_7109,N_8986);
nand U11674 (N_11674,N_6565,N_7627);
and U11675 (N_11675,N_8089,N_9269);
or U11676 (N_11676,N_7369,N_7174);
nor U11677 (N_11677,N_5652,N_9291);
or U11678 (N_11678,N_5324,N_6474);
and U11679 (N_11679,N_9596,N_6858);
or U11680 (N_11680,N_5001,N_9680);
xnor U11681 (N_11681,N_6527,N_8522);
and U11682 (N_11682,N_7831,N_8395);
or U11683 (N_11683,N_7856,N_9473);
or U11684 (N_11684,N_6710,N_9743);
and U11685 (N_11685,N_9789,N_8126);
or U11686 (N_11686,N_5306,N_5621);
nand U11687 (N_11687,N_9121,N_5525);
nor U11688 (N_11688,N_9843,N_5038);
or U11689 (N_11689,N_7549,N_9147);
nand U11690 (N_11690,N_6203,N_5589);
xnor U11691 (N_11691,N_9136,N_8229);
or U11692 (N_11692,N_6757,N_9210);
and U11693 (N_11693,N_9844,N_6012);
nand U11694 (N_11694,N_8792,N_5165);
nand U11695 (N_11695,N_8408,N_5717);
and U11696 (N_11696,N_5345,N_8952);
nand U11697 (N_11697,N_7606,N_5963);
nand U11698 (N_11698,N_5834,N_8441);
or U11699 (N_11699,N_8887,N_6966);
and U11700 (N_11700,N_6839,N_9954);
nand U11701 (N_11701,N_6045,N_6515);
and U11702 (N_11702,N_8082,N_6230);
or U11703 (N_11703,N_8446,N_5984);
nor U11704 (N_11704,N_6077,N_7520);
and U11705 (N_11705,N_7762,N_6951);
or U11706 (N_11706,N_5600,N_7814);
or U11707 (N_11707,N_8245,N_5840);
nor U11708 (N_11708,N_7527,N_7792);
nand U11709 (N_11709,N_5150,N_9519);
xor U11710 (N_11710,N_5441,N_6093);
and U11711 (N_11711,N_7959,N_6030);
and U11712 (N_11712,N_6695,N_5919);
nand U11713 (N_11713,N_5575,N_9939);
or U11714 (N_11714,N_9982,N_6020);
or U11715 (N_11715,N_8776,N_5977);
nand U11716 (N_11716,N_8279,N_9933);
and U11717 (N_11717,N_6058,N_8435);
and U11718 (N_11718,N_9623,N_6521);
or U11719 (N_11719,N_7917,N_9200);
nor U11720 (N_11720,N_7165,N_6611);
or U11721 (N_11721,N_8293,N_6931);
or U11722 (N_11722,N_5703,N_6922);
and U11723 (N_11723,N_8252,N_9803);
or U11724 (N_11724,N_9983,N_8587);
or U11725 (N_11725,N_6279,N_7999);
or U11726 (N_11726,N_8423,N_7215);
or U11727 (N_11727,N_8716,N_6119);
or U11728 (N_11728,N_5739,N_6099);
nor U11729 (N_11729,N_9021,N_9674);
and U11730 (N_11730,N_6008,N_9689);
nor U11731 (N_11731,N_7770,N_6927);
nand U11732 (N_11732,N_8509,N_6495);
or U11733 (N_11733,N_9723,N_5757);
and U11734 (N_11734,N_5715,N_5287);
xor U11735 (N_11735,N_9725,N_5891);
or U11736 (N_11736,N_9598,N_7130);
nor U11737 (N_11737,N_7602,N_8107);
and U11738 (N_11738,N_7686,N_9105);
nor U11739 (N_11739,N_9378,N_7641);
nand U11740 (N_11740,N_8913,N_5756);
and U11741 (N_11741,N_8404,N_9175);
nand U11742 (N_11742,N_6945,N_8111);
nand U11743 (N_11743,N_9265,N_5367);
nor U11744 (N_11744,N_8295,N_7585);
nand U11745 (N_11745,N_8205,N_5276);
and U11746 (N_11746,N_7966,N_9879);
and U11747 (N_11747,N_8728,N_8762);
or U11748 (N_11748,N_9196,N_9350);
or U11749 (N_11749,N_6996,N_9256);
or U11750 (N_11750,N_9924,N_8768);
nand U11751 (N_11751,N_7028,N_7373);
or U11752 (N_11752,N_5293,N_6629);
nor U11753 (N_11753,N_6642,N_6657);
and U11754 (N_11754,N_9654,N_6437);
and U11755 (N_11755,N_6088,N_9189);
nor U11756 (N_11756,N_8254,N_5888);
or U11757 (N_11757,N_7242,N_8092);
or U11758 (N_11758,N_8846,N_6833);
nor U11759 (N_11759,N_9923,N_7972);
nand U11760 (N_11760,N_9449,N_5332);
nand U11761 (N_11761,N_8863,N_7629);
and U11762 (N_11762,N_8356,N_7217);
nor U11763 (N_11763,N_7783,N_6195);
or U11764 (N_11764,N_5552,N_6150);
nand U11765 (N_11765,N_9297,N_8016);
or U11766 (N_11766,N_5188,N_9791);
and U11767 (N_11767,N_6217,N_6987);
and U11768 (N_11768,N_6786,N_5553);
or U11769 (N_11769,N_9308,N_5505);
or U11770 (N_11770,N_8101,N_9710);
or U11771 (N_11771,N_6464,N_7108);
or U11772 (N_11772,N_6877,N_5933);
and U11773 (N_11773,N_8791,N_6766);
and U11774 (N_11774,N_5742,N_6142);
nor U11775 (N_11775,N_7289,N_9198);
or U11776 (N_11776,N_5789,N_8881);
nor U11777 (N_11777,N_7492,N_8489);
nand U11778 (N_11778,N_7542,N_9713);
or U11779 (N_11779,N_8417,N_9752);
and U11780 (N_11780,N_9155,N_6588);
nor U11781 (N_11781,N_8511,N_8077);
nand U11782 (N_11782,N_9992,N_6992);
nor U11783 (N_11783,N_6418,N_5160);
nand U11784 (N_11784,N_9319,N_7129);
or U11785 (N_11785,N_8302,N_8294);
nand U11786 (N_11786,N_9751,N_9232);
nor U11787 (N_11787,N_7987,N_9902);
nor U11788 (N_11788,N_9440,N_5207);
nand U11789 (N_11789,N_5423,N_6046);
and U11790 (N_11790,N_8345,N_6807);
xor U11791 (N_11791,N_9688,N_8621);
and U11792 (N_11792,N_7816,N_7703);
nand U11793 (N_11793,N_6499,N_7855);
nor U11794 (N_11794,N_5679,N_6990);
nand U11795 (N_11795,N_7096,N_5036);
nand U11796 (N_11796,N_5993,N_7283);
nor U11797 (N_11797,N_5171,N_7829);
nor U11798 (N_11798,N_7310,N_6767);
nand U11799 (N_11799,N_8757,N_7372);
nor U11800 (N_11800,N_9025,N_5006);
nand U11801 (N_11801,N_5983,N_5225);
xor U11802 (N_11802,N_8344,N_7922);
and U11803 (N_11803,N_8927,N_9672);
or U11804 (N_11804,N_9248,N_9631);
and U11805 (N_11805,N_8442,N_8506);
or U11806 (N_11806,N_9640,N_6053);
and U11807 (N_11807,N_9282,N_8306);
or U11808 (N_11808,N_9512,N_5961);
nand U11809 (N_11809,N_6294,N_6540);
nand U11810 (N_11810,N_5266,N_8853);
nor U11811 (N_11811,N_6465,N_9894);
xnor U11812 (N_11812,N_5510,N_5956);
and U11813 (N_11813,N_7475,N_9642);
nand U11814 (N_11814,N_9253,N_9142);
nand U11815 (N_11815,N_9786,N_7822);
nand U11816 (N_11816,N_6031,N_6608);
nor U11817 (N_11817,N_8325,N_5771);
nor U11818 (N_11818,N_7023,N_5649);
nand U11819 (N_11819,N_6141,N_8368);
or U11820 (N_11820,N_6489,N_5454);
or U11821 (N_11821,N_6641,N_8635);
nor U11822 (N_11822,N_5466,N_5351);
or U11823 (N_11823,N_6533,N_8179);
and U11824 (N_11824,N_7713,N_7017);
nand U11825 (N_11825,N_8218,N_5498);
and U11826 (N_11826,N_9964,N_8987);
and U11827 (N_11827,N_5440,N_7360);
nand U11828 (N_11828,N_7886,N_6333);
nor U11829 (N_11829,N_5159,N_6912);
nor U11830 (N_11830,N_9797,N_8646);
and U11831 (N_11831,N_5007,N_5561);
nand U11832 (N_11832,N_8970,N_5368);
and U11833 (N_11833,N_9755,N_8893);
and U11834 (N_11834,N_5777,N_7621);
nor U11835 (N_11835,N_5996,N_5314);
or U11836 (N_11836,N_7404,N_6477);
nor U11837 (N_11837,N_7907,N_6885);
and U11838 (N_11838,N_7296,N_8917);
nor U11839 (N_11839,N_6387,N_7810);
or U11840 (N_11840,N_5953,N_5099);
nor U11841 (N_11841,N_6210,N_8268);
nor U11842 (N_11842,N_5418,N_7008);
and U11843 (N_11843,N_8622,N_8759);
or U11844 (N_11844,N_7588,N_5536);
nor U11845 (N_11845,N_5122,N_8103);
nand U11846 (N_11846,N_6559,N_7828);
nor U11847 (N_11847,N_8180,N_9061);
or U11848 (N_11848,N_6846,N_6409);
and U11849 (N_11849,N_9173,N_8932);
nor U11850 (N_11850,N_9859,N_9691);
or U11851 (N_11851,N_9391,N_8894);
nand U11852 (N_11852,N_9771,N_7663);
nor U11853 (N_11853,N_5309,N_8068);
nor U11854 (N_11854,N_6027,N_9777);
or U11855 (N_11855,N_5083,N_6761);
or U11856 (N_11856,N_7570,N_6651);
nor U11857 (N_11857,N_9699,N_8140);
nor U11858 (N_11858,N_5898,N_6110);
or U11859 (N_11859,N_8242,N_7413);
or U11860 (N_11860,N_5467,N_7933);
nand U11861 (N_11861,N_8959,N_7803);
and U11862 (N_11862,N_7092,N_6688);
nand U11863 (N_11863,N_9561,N_7302);
nand U11864 (N_11864,N_9991,N_8809);
and U11865 (N_11865,N_7591,N_8436);
and U11866 (N_11866,N_6653,N_9401);
or U11867 (N_11867,N_9484,N_7233);
and U11868 (N_11868,N_6443,N_6814);
or U11869 (N_11869,N_7133,N_9919);
xnor U11870 (N_11870,N_9588,N_5716);
nor U11871 (N_11871,N_6968,N_9498);
or U11872 (N_11872,N_5659,N_5712);
and U11873 (N_11873,N_7480,N_5954);
xnor U11874 (N_11874,N_8883,N_8457);
or U11875 (N_11875,N_8594,N_5250);
and U11876 (N_11876,N_8744,N_8787);
and U11877 (N_11877,N_6232,N_5456);
nand U11878 (N_11878,N_8032,N_6178);
and U11879 (N_11879,N_7102,N_6667);
or U11880 (N_11880,N_8892,N_6622);
nand U11881 (N_11881,N_7645,N_8727);
and U11882 (N_11882,N_5867,N_8403);
or U11883 (N_11883,N_7628,N_8730);
or U11884 (N_11884,N_8409,N_6919);
and U11885 (N_11885,N_8697,N_5436);
nor U11886 (N_11886,N_9509,N_7837);
nand U11887 (N_11887,N_5930,N_6241);
and U11888 (N_11888,N_6180,N_6036);
and U11889 (N_11889,N_9828,N_6665);
or U11890 (N_11890,N_7059,N_8833);
and U11891 (N_11891,N_5043,N_7416);
xor U11892 (N_11892,N_5319,N_6655);
or U11893 (N_11893,N_6028,N_5829);
nand U11894 (N_11894,N_5496,N_8972);
and U11895 (N_11895,N_8080,N_7187);
nand U11896 (N_11896,N_5509,N_7638);
and U11897 (N_11897,N_8250,N_9211);
or U11898 (N_11898,N_8541,N_8502);
nand U11899 (N_11899,N_9830,N_5114);
nand U11900 (N_11900,N_9700,N_5393);
nand U11901 (N_11901,N_7690,N_5874);
nand U11902 (N_11902,N_5545,N_7234);
or U11903 (N_11903,N_7869,N_9810);
and U11904 (N_11904,N_9292,N_7384);
nor U11905 (N_11905,N_8159,N_9950);
xnor U11906 (N_11906,N_6300,N_5164);
or U11907 (N_11907,N_7457,N_6648);
nand U11908 (N_11908,N_9971,N_8648);
and U11909 (N_11909,N_7993,N_8641);
or U11910 (N_11910,N_6483,N_6609);
or U11911 (N_11911,N_8367,N_9475);
and U11912 (N_11912,N_9501,N_6601);
or U11913 (N_11913,N_9686,N_6325);
or U11914 (N_11914,N_7796,N_6268);
nand U11915 (N_11915,N_7746,N_7381);
nand U11916 (N_11916,N_8233,N_9724);
nor U11917 (N_11917,N_6080,N_8451);
nand U11918 (N_11918,N_9569,N_6151);
nor U11919 (N_11919,N_8696,N_8387);
nor U11920 (N_11920,N_8775,N_7036);
or U11921 (N_11921,N_7076,N_6318);
nand U11922 (N_11922,N_7514,N_6442);
xnor U11923 (N_11923,N_5630,N_6745);
nor U11924 (N_11924,N_6277,N_8371);
or U11925 (N_11925,N_9646,N_7624);
or U11926 (N_11926,N_7318,N_9748);
nor U11927 (N_11927,N_7887,N_9081);
nand U11928 (N_11928,N_6397,N_7935);
or U11929 (N_11929,N_9371,N_8550);
or U11930 (N_11930,N_8507,N_9782);
or U11931 (N_11931,N_6978,N_7755);
and U11932 (N_11932,N_5626,N_8589);
and U11933 (N_11933,N_8662,N_6896);
nor U11934 (N_11934,N_8686,N_6962);
or U11935 (N_11935,N_5860,N_9955);
nand U11936 (N_11936,N_9594,N_6129);
nor U11937 (N_11937,N_5227,N_9209);
or U11938 (N_11938,N_6310,N_7235);
nor U11939 (N_11939,N_6191,N_5158);
and U11940 (N_11940,N_7001,N_6706);
or U11941 (N_11941,N_6140,N_8004);
and U11942 (N_11942,N_9912,N_9069);
and U11943 (N_11943,N_6760,N_6462);
nor U11944 (N_11944,N_8064,N_5620);
nor U11945 (N_11945,N_8379,N_7245);
nor U11946 (N_11946,N_7852,N_5808);
nor U11947 (N_11947,N_9578,N_7459);
nor U11948 (N_11948,N_7505,N_6286);
or U11949 (N_11949,N_6201,N_6136);
and U11950 (N_11950,N_8773,N_8213);
xnor U11951 (N_11951,N_5497,N_9015);
nor U11952 (N_11952,N_7473,N_6255);
nor U11953 (N_11953,N_5468,N_6040);
and U11954 (N_11954,N_8981,N_5237);
and U11955 (N_11955,N_6258,N_8977);
nand U11956 (N_11956,N_9244,N_5782);
or U11957 (N_11957,N_9715,N_7185);
and U11958 (N_11958,N_7104,N_7257);
nor U11959 (N_11959,N_9582,N_7249);
and U11960 (N_11960,N_5359,N_8200);
xor U11961 (N_11961,N_9600,N_9294);
and U11962 (N_11962,N_7147,N_9231);
nand U11963 (N_11963,N_8999,N_6708);
nor U11964 (N_11964,N_5453,N_5741);
nor U11965 (N_11965,N_5251,N_6236);
nor U11966 (N_11966,N_5538,N_8882);
and U11967 (N_11967,N_5173,N_8127);
nand U11968 (N_11968,N_7719,N_6075);
or U11969 (N_11969,N_9679,N_8452);
and U11970 (N_11970,N_8747,N_7253);
nor U11971 (N_11971,N_9574,N_6138);
nor U11972 (N_11972,N_8607,N_6434);
nand U11973 (N_11973,N_6265,N_7596);
and U11974 (N_11974,N_9362,N_8647);
nor U11975 (N_11975,N_7477,N_5672);
xnor U11976 (N_11976,N_7132,N_9504);
or U11977 (N_11977,N_7175,N_6132);
nand U11978 (N_11978,N_6977,N_9571);
and U11979 (N_11979,N_6159,N_5516);
or U11980 (N_11980,N_5026,N_8871);
nor U11981 (N_11981,N_7938,N_6941);
and U11982 (N_11982,N_8895,N_8407);
nor U11983 (N_11983,N_9827,N_8750);
or U11984 (N_11984,N_7765,N_7075);
and U11985 (N_11985,N_8232,N_8378);
nand U11986 (N_11986,N_9809,N_8498);
and U11987 (N_11987,N_9505,N_8120);
and U11988 (N_11988,N_5674,N_9233);
or U11989 (N_11989,N_7265,N_7858);
nand U11990 (N_11990,N_9289,N_6354);
and U11991 (N_11991,N_8663,N_6456);
nor U11992 (N_11992,N_7842,N_9862);
and U11993 (N_11993,N_5003,N_6484);
nor U11994 (N_11994,N_8568,N_5151);
nand U11995 (N_11995,N_9309,N_6470);
and U11996 (N_11996,N_7605,N_6317);
nor U11997 (N_11997,N_9195,N_7313);
nor U11998 (N_11998,N_7760,N_5220);
or U11999 (N_11999,N_6696,N_9910);
nand U12000 (N_12000,N_7012,N_6590);
or U12001 (N_12001,N_5012,N_9161);
nand U12002 (N_12002,N_6249,N_8118);
nand U12003 (N_12003,N_8173,N_9847);
and U12004 (N_12004,N_6610,N_9376);
nor U12005 (N_12005,N_7998,N_8777);
or U12006 (N_12006,N_8040,N_7976);
nand U12007 (N_12007,N_7509,N_6379);
xor U12008 (N_12008,N_7961,N_9014);
nand U12009 (N_12009,N_6759,N_9358);
nand U12010 (N_12010,N_8655,N_5474);
and U12011 (N_12011,N_8790,N_9733);
or U12012 (N_12012,N_8692,N_5095);
and U12013 (N_12013,N_7315,N_6689);
nand U12014 (N_12014,N_6522,N_9584);
xor U12015 (N_12015,N_8941,N_9533);
nand U12016 (N_12016,N_9461,N_6289);
and U12017 (N_12017,N_7330,N_9634);
nor U12018 (N_12018,N_9042,N_6856);
or U12019 (N_12019,N_6435,N_5906);
nor U12020 (N_12020,N_6541,N_9604);
nand U12021 (N_12021,N_7574,N_8711);
nand U12022 (N_12022,N_8735,N_5406);
nand U12023 (N_12023,N_7254,N_6517);
and U12024 (N_12024,N_7772,N_5631);
and U12025 (N_12025,N_7553,N_5362);
nor U12026 (N_12026,N_6639,N_6652);
nor U12027 (N_12027,N_5939,N_9946);
and U12028 (N_12028,N_5524,N_6557);
nor U12029 (N_12029,N_7476,N_5578);
and U12030 (N_12030,N_8869,N_8654);
or U12031 (N_12031,N_5923,N_9435);
or U12032 (N_12032,N_8723,N_8569);
or U12033 (N_12033,N_8889,N_9678);
and U12034 (N_12034,N_6799,N_5446);
and U12035 (N_12035,N_6883,N_8315);
or U12036 (N_12036,N_8916,N_5704);
nor U12037 (N_12037,N_5020,N_6790);
nand U12038 (N_12038,N_8888,N_8153);
and U12039 (N_12039,N_6059,N_7738);
nand U12040 (N_12040,N_5350,N_7521);
nand U12041 (N_12041,N_8100,N_6763);
or U12042 (N_12042,N_7662,N_6750);
or U12043 (N_12043,N_7704,N_7841);
nor U12044 (N_12044,N_9385,N_6116);
or U12045 (N_12045,N_6491,N_8557);
nor U12046 (N_12046,N_6284,N_9100);
or U12047 (N_12047,N_5810,N_7557);
and U12048 (N_12048,N_9437,N_5732);
nand U12049 (N_12049,N_5676,N_5391);
or U12050 (N_12050,N_6363,N_7427);
or U12051 (N_12051,N_9528,N_5773);
and U12052 (N_12052,N_7449,N_6478);
nand U12053 (N_12053,N_7389,N_6889);
nor U12054 (N_12054,N_7340,N_8828);
nor U12055 (N_12055,N_7409,N_6417);
nor U12056 (N_12056,N_7533,N_5573);
nand U12057 (N_12057,N_6155,N_9683);
nand U12058 (N_12058,N_9833,N_8673);
nand U12059 (N_12059,N_6724,N_8935);
and U12060 (N_12060,N_7040,N_8480);
or U12061 (N_12061,N_7673,N_5915);
or U12062 (N_12062,N_9432,N_9936);
xnor U12063 (N_12063,N_5927,N_8059);
nor U12064 (N_12064,N_8891,N_7963);
nor U12065 (N_12065,N_8748,N_9741);
and U12066 (N_12066,N_6316,N_5724);
nand U12067 (N_12067,N_8286,N_6743);
nand U12068 (N_12068,N_7693,N_8707);
nand U12069 (N_12069,N_9953,N_8753);
nand U12070 (N_12070,N_9419,N_7052);
or U12071 (N_12071,N_7305,N_6179);
or U12072 (N_12072,N_5174,N_5427);
nand U12073 (N_12073,N_5529,N_7695);
or U12074 (N_12074,N_7406,N_8104);
and U12075 (N_12075,N_5000,N_9866);
or U12076 (N_12076,N_6791,N_6021);
or U12077 (N_12077,N_6514,N_9555);
nor U12078 (N_12078,N_8634,N_6550);
and U12079 (N_12079,N_8947,N_9620);
or U12080 (N_12080,N_5216,N_5428);
nor U12081 (N_12081,N_5254,N_5478);
and U12082 (N_12082,N_6415,N_7271);
nor U12083 (N_12083,N_5264,N_9323);
and U12084 (N_12084,N_5574,N_9861);
nor U12085 (N_12085,N_6450,N_6520);
nand U12086 (N_12086,N_6496,N_5787);
and U12087 (N_12087,N_9339,N_7286);
or U12088 (N_12088,N_8538,N_8687);
or U12089 (N_12089,N_7110,N_7754);
or U12090 (N_12090,N_6248,N_9832);
or U12091 (N_12091,N_8857,N_5628);
or U12092 (N_12092,N_7934,N_9849);
nor U12093 (N_12093,N_6923,N_7550);
or U12094 (N_12094,N_9995,N_9224);
nor U12095 (N_12095,N_5602,N_9622);
nand U12096 (N_12096,N_5039,N_8493);
and U12097 (N_12097,N_6811,N_5301);
or U12098 (N_12098,N_8207,N_6583);
or U12099 (N_12099,N_7131,N_5033);
nand U12100 (N_12100,N_9937,N_9563);
nand U12101 (N_12101,N_9502,N_5294);
nand U12102 (N_12102,N_7702,N_7345);
or U12103 (N_12103,N_8818,N_7652);
nand U12104 (N_12104,N_6256,N_9351);
nand U12105 (N_12105,N_8062,N_9341);
xor U12106 (N_12106,N_7827,N_5064);
nand U12107 (N_12107,N_5544,N_8936);
and U12108 (N_12108,N_9367,N_7801);
nor U12109 (N_12109,N_5881,N_6276);
and U12110 (N_12110,N_9570,N_9567);
or U12111 (N_12111,N_9538,N_6372);
or U12112 (N_12112,N_6685,N_8829);
nand U12113 (N_12113,N_6475,N_5555);
nor U12114 (N_12114,N_5666,N_8346);
or U12115 (N_12115,N_7789,N_7955);
and U12116 (N_12116,N_9239,N_8141);
nor U12117 (N_12117,N_5821,N_8765);
nand U12118 (N_12118,N_5420,N_6733);
nand U12119 (N_12119,N_9981,N_6678);
nand U12120 (N_12120,N_5125,N_5877);
or U12121 (N_12121,N_7508,N_6801);
and U12122 (N_12122,N_8770,N_8183);
nor U12123 (N_12123,N_9466,N_9703);
or U12124 (N_12124,N_6072,N_6113);
nor U12125 (N_12125,N_8195,N_7522);
or U12126 (N_12126,N_8144,N_7100);
nand U12127 (N_12127,N_7350,N_7504);
nor U12128 (N_12128,N_8182,N_6857);
nand U12129 (N_12129,N_9774,N_8797);
and U12130 (N_12130,N_5708,N_5283);
or U12131 (N_12131,N_9192,N_5361);
or U12132 (N_12132,N_5271,N_9867);
or U12133 (N_12133,N_8000,N_5296);
nand U12134 (N_12134,N_6328,N_5144);
nand U12135 (N_12135,N_7171,N_7377);
nand U12136 (N_12136,N_8224,N_8365);
or U12137 (N_12137,N_9959,N_8989);
nand U12138 (N_12138,N_9356,N_8618);
and U12139 (N_12139,N_7051,N_8855);
or U12140 (N_12140,N_5965,N_6929);
nor U12141 (N_12141,N_8017,N_5219);
or U12142 (N_12142,N_8722,N_6744);
and U12143 (N_12143,N_6096,N_7238);
nor U12144 (N_12144,N_5850,N_6193);
nor U12145 (N_12145,N_5681,N_8953);
nor U12146 (N_12146,N_5949,N_7566);
nor U12147 (N_12147,N_9041,N_5655);
xnor U12148 (N_12148,N_7825,N_9422);
or U12149 (N_12149,N_9908,N_5761);
nand U12150 (N_12150,N_6737,N_5828);
nor U12151 (N_12151,N_9921,N_8661);
xor U12152 (N_12152,N_7002,N_7683);
nand U12153 (N_12153,N_6147,N_5800);
and U12154 (N_12154,N_5485,N_6085);
nand U12155 (N_12155,N_6413,N_8950);
and U12156 (N_12156,N_5596,N_9290);
and U12157 (N_12157,N_6043,N_8392);
and U12158 (N_12158,N_8002,N_6016);
nand U12159 (N_12159,N_9409,N_5697);
and U12160 (N_12160,N_8010,N_9669);
nand U12161 (N_12161,N_9283,N_7866);
and U12162 (N_12162,N_8820,N_9630);
or U12163 (N_12163,N_7140,N_6932);
and U12164 (N_12164,N_5088,N_8599);
nand U12165 (N_12165,N_8221,N_9217);
nand U12166 (N_12166,N_5426,N_8188);
xor U12167 (N_12167,N_6398,N_9090);
and U12168 (N_12168,N_5556,N_7329);
and U12169 (N_12169,N_5503,N_6039);
and U12170 (N_12170,N_5526,N_6783);
nand U12171 (N_12171,N_8993,N_7724);
and U12172 (N_12172,N_9333,N_8928);
and U12173 (N_12173,N_6647,N_8585);
nand U12174 (N_12174,N_6960,N_9838);
and U12175 (N_12175,N_6845,N_8610);
and U12176 (N_12176,N_8060,N_8063);
nor U12177 (N_12177,N_8096,N_8732);
nor U12178 (N_12178,N_5520,N_8702);
nand U12179 (N_12179,N_8799,N_6420);
nor U12180 (N_12180,N_8746,N_6408);
or U12181 (N_12181,N_5370,N_8902);
nor U12182 (N_12182,N_8593,N_8070);
nor U12183 (N_12183,N_7545,N_9486);
nor U12184 (N_12184,N_7800,N_5714);
nand U12185 (N_12185,N_8309,N_8257);
or U12186 (N_12186,N_5865,N_6184);
nand U12187 (N_12187,N_5189,N_6497);
and U12188 (N_12188,N_8398,N_5145);
nor U12189 (N_12189,N_8824,N_5197);
or U12190 (N_12190,N_5048,N_5242);
or U12191 (N_12191,N_6473,N_7689);
and U12192 (N_12192,N_7775,N_8370);
or U12193 (N_12193,N_7222,N_9508);
nand U12194 (N_12194,N_5460,N_8650);
or U12195 (N_12195,N_8934,N_9930);
nand U12196 (N_12196,N_5475,N_5585);
and U12197 (N_12197,N_8530,N_7483);
nor U12198 (N_12198,N_8865,N_6356);
and U12199 (N_12199,N_8169,N_6976);
nor U12200 (N_12200,N_7347,N_8800);
or U12201 (N_12201,N_5764,N_9878);
and U12202 (N_12202,N_8975,N_9157);
and U12203 (N_12203,N_5086,N_6320);
nand U12204 (N_12204,N_5830,N_6633);
nand U12205 (N_12205,N_5815,N_6283);
and U12206 (N_12206,N_9111,N_7651);
or U12207 (N_12207,N_9531,N_9303);
nand U12208 (N_12208,N_9825,N_8609);
and U12209 (N_12209,N_9030,N_8866);
and U12210 (N_12210,N_5204,N_5390);
and U12211 (N_12211,N_9800,N_6433);
and U12212 (N_12212,N_8677,N_9446);
and U12213 (N_12213,N_8623,N_8598);
nand U12214 (N_12214,N_7537,N_7019);
and U12215 (N_12215,N_5740,N_6524);
nor U12216 (N_12216,N_9478,N_8929);
nand U12217 (N_12217,N_8056,N_5582);
and U12218 (N_12218,N_6558,N_7742);
and U12219 (N_12219,N_7850,N_9027);
or U12220 (N_12220,N_8394,N_7120);
and U12221 (N_12221,N_6160,N_6621);
nor U12222 (N_12222,N_9052,N_7044);
nand U12223 (N_12223,N_7649,N_9738);
or U12224 (N_12224,N_8899,N_7361);
or U12225 (N_12225,N_5962,N_7343);
or U12226 (N_12226,N_6573,N_9957);
or U12227 (N_12227,N_7528,N_7499);
and U12228 (N_12228,N_9071,N_5070);
and U12229 (N_12229,N_8858,N_9976);
or U12230 (N_12230,N_8500,N_9922);
nand U12231 (N_12231,N_7734,N_8431);
and U12232 (N_12232,N_7722,N_8353);
or U12233 (N_12233,N_9086,N_6511);
nor U12234 (N_12234,N_6679,N_6090);
nand U12235 (N_12235,N_9840,N_9718);
nor U12236 (N_12236,N_7705,N_7325);
or U12237 (N_12237,N_9635,N_6512);
nand U12238 (N_12238,N_7725,N_5410);
nand U12239 (N_12239,N_8198,N_7900);
nand U12240 (N_12240,N_6874,N_5768);
and U12241 (N_12241,N_6862,N_5055);
or U12242 (N_12242,N_7144,N_7359);
xor U12243 (N_12243,N_5869,N_6117);
and U12244 (N_12244,N_9543,N_8679);
or U12245 (N_12245,N_7194,N_8766);
and U12246 (N_12246,N_7631,N_7119);
nand U12247 (N_12247,N_7623,N_8841);
nand U12248 (N_12248,N_7946,N_7128);
nand U12249 (N_12249,N_7170,N_8066);
and U12250 (N_12250,N_6348,N_8411);
and U12251 (N_12251,N_5905,N_7263);
or U12252 (N_12252,N_9758,N_8691);
or U12253 (N_12253,N_6820,N_6950);
nand U12254 (N_12254,N_8312,N_5622);
xnor U12255 (N_12255,N_7750,N_8227);
nor U12256 (N_12256,N_8151,N_8767);
or U12257 (N_12257,N_9476,N_9251);
nand U12258 (N_12258,N_9271,N_7455);
nor U12259 (N_12259,N_6492,N_6650);
nor U12260 (N_12260,N_9711,N_9222);
nor U12261 (N_12261,N_8481,N_9203);
and U12262 (N_12262,N_8581,N_7890);
nand U12263 (N_12263,N_9279,N_9006);
nand U12264 (N_12264,N_8532,N_8174);
and U12265 (N_12265,N_7517,N_8425);
and U12266 (N_12266,N_9438,N_5398);
nand U12267 (N_12267,N_7220,N_6902);
nand U12268 (N_12268,N_5268,N_5377);
nand U12269 (N_12269,N_7326,N_7857);
and U12270 (N_12270,N_5069,N_7105);
and U12271 (N_12271,N_8967,N_7560);
or U12272 (N_12272,N_9513,N_9818);
and U12273 (N_12273,N_6211,N_5847);
nor U12274 (N_12274,N_7950,N_6223);
or U12275 (N_12275,N_5633,N_6054);
and U12276 (N_12276,N_7368,N_8152);
and U12277 (N_12277,N_8736,N_5663);
nor U12278 (N_12278,N_8380,N_8526);
nor U12279 (N_12279,N_8470,N_6551);
nor U12280 (N_12280,N_5872,N_8001);
nand U12281 (N_12281,N_5384,N_5647);
nand U12282 (N_12282,N_8135,N_9965);
nor U12283 (N_12283,N_8712,N_6768);
nor U12284 (N_12284,N_5166,N_7839);
nand U12285 (N_12285,N_6468,N_6364);
nor U12286 (N_12286,N_9179,N_9985);
or U12287 (N_12287,N_9850,N_9736);
or U12288 (N_12288,N_9487,N_7782);
or U12289 (N_12289,N_8381,N_5786);
nand U12290 (N_12290,N_9804,N_7152);
and U12291 (N_12291,N_5557,N_6942);
nor U12292 (N_12292,N_5817,N_8400);
or U12293 (N_12293,N_9972,N_9816);
and U12294 (N_12294,N_6124,N_5141);
or U12295 (N_12295,N_5942,N_8971);
nand U12296 (N_12296,N_7672,N_8283);
or U12297 (N_12297,N_7636,N_9778);
or U12298 (N_12298,N_8258,N_6024);
and U12299 (N_12299,N_5759,N_7586);
or U12300 (N_12300,N_6925,N_8703);
nand U12301 (N_12301,N_7951,N_7712);
or U12302 (N_12302,N_8683,N_5968);
xnor U12303 (N_12303,N_5776,N_6311);
nor U12304 (N_12304,N_7431,N_5313);
nand U12305 (N_12305,N_9602,N_7766);
or U12306 (N_12306,N_5177,N_7868);
nor U12307 (N_12307,N_9632,N_5677);
nor U12308 (N_12308,N_9057,N_7266);
nand U12309 (N_12309,N_8485,N_9326);
nand U12310 (N_12310,N_5619,N_5744);
nor U12311 (N_12311,N_8138,N_5814);
and U12312 (N_12312,N_9527,N_7443);
nand U12313 (N_12313,N_6946,N_5827);
or U12314 (N_12314,N_8512,N_9260);
nor U12315 (N_12315,N_8969,N_8566);
and U12316 (N_12316,N_7412,N_7440);
or U12317 (N_12317,N_8241,N_7460);
or U12318 (N_12318,N_8476,N_8094);
nor U12319 (N_12319,N_5201,N_9551);
or U12320 (N_12320,N_7920,N_6584);
or U12321 (N_12321,N_8117,N_7252);
or U12322 (N_12322,N_5892,N_7048);
xnor U12323 (N_12323,N_9079,N_5887);
nor U12324 (N_12324,N_6698,N_7824);
and U12325 (N_12325,N_9107,N_6038);
nand U12326 (N_12326,N_6831,N_7815);
and U12327 (N_12327,N_6888,N_5118);
or U12328 (N_12328,N_7486,N_9880);
nand U12329 (N_12329,N_6157,N_5019);
nor U12330 (N_12330,N_9037,N_8719);
or U12331 (N_12331,N_6979,N_6853);
xor U12332 (N_12332,N_8147,N_9181);
nor U12333 (N_12333,N_6810,N_8908);
nor U12334 (N_12334,N_9148,N_9074);
nand U12335 (N_12335,N_9410,N_6229);
and U12336 (N_12336,N_5957,N_9656);
nor U12337 (N_12337,N_6269,N_5259);
nor U12338 (N_12338,N_6097,N_8496);
nand U12339 (N_12339,N_5042,N_9130);
and U12340 (N_12340,N_5762,N_9766);
nor U12341 (N_12341,N_7114,N_8044);
or U12342 (N_12342,N_5609,N_8122);
or U12343 (N_12343,N_8998,N_7199);
or U12344 (N_12344,N_9532,N_9293);
nand U12345 (N_12345,N_5060,N_6884);
nor U12346 (N_12346,N_6339,N_8083);
or U12347 (N_12347,N_6458,N_5970);
and U12348 (N_12348,N_9227,N_9737);
or U12349 (N_12349,N_5334,N_7094);
and U12350 (N_12350,N_7862,N_5289);
and U12351 (N_12351,N_9768,N_7915);
nand U12352 (N_12352,N_6762,N_8903);
nand U12353 (N_12353,N_8943,N_8611);
nor U12354 (N_12354,N_6660,N_8495);
nand U12355 (N_12355,N_8974,N_9369);
and U12356 (N_12356,N_5976,N_5844);
nand U12357 (N_12357,N_6347,N_6062);
nand U12358 (N_12358,N_7637,N_7365);
nand U12359 (N_12359,N_8390,N_5730);
nand U12360 (N_12360,N_7727,N_5274);
nand U12361 (N_12361,N_9877,N_6022);
nor U12362 (N_12362,N_5644,N_7039);
nor U12363 (N_12363,N_9790,N_9746);
or U12364 (N_12364,N_9066,N_5490);
nand U12365 (N_12365,N_7698,N_7118);
nand U12366 (N_12366,N_7975,N_6322);
nor U12367 (N_12367,N_8487,N_9467);
nand U12368 (N_12368,N_9864,N_7821);
nor U12369 (N_12369,N_5711,N_7595);
nand U12370 (N_12370,N_9128,N_8199);
nand U12371 (N_12371,N_9779,N_6366);
nand U12372 (N_12372,N_7925,N_8261);
nand U12373 (N_12373,N_8786,N_7905);
or U12374 (N_12374,N_9928,N_9956);
nor U12375 (N_12375,N_8048,N_7674);
nand U12376 (N_12376,N_6721,N_7647);
or U12377 (N_12377,N_8226,N_8239);
or U12378 (N_12378,N_6445,N_6187);
xor U12379 (N_12379,N_9769,N_6869);
and U12380 (N_12380,N_6549,N_9745);
nand U12381 (N_12381,N_9412,N_6390);
and U12382 (N_12382,N_9275,N_7681);
or U12383 (N_12383,N_9429,N_9144);
or U12384 (N_12384,N_7524,N_5376);
and U12385 (N_12385,N_7726,N_5684);
nand U12386 (N_12386,N_9443,N_7733);
nand U12387 (N_12387,N_6545,N_9447);
nand U12388 (N_12388,N_7364,N_5615);
nor U12389 (N_12389,N_6732,N_5871);
nor U12390 (N_12390,N_6544,N_5120);
or U12391 (N_12391,N_6972,N_6518);
and U12392 (N_12392,N_5476,N_8391);
nand U12393 (N_12393,N_6994,N_8674);
and U12394 (N_12394,N_6221,N_5979);
nor U12395 (N_12395,N_9448,N_6683);
nor U12396 (N_12396,N_5068,N_8656);
nand U12397 (N_12397,N_8287,N_8416);
and U12398 (N_12398,N_8468,N_9979);
or U12399 (N_12399,N_5263,N_5598);
xor U12400 (N_12400,N_6094,N_5959);
and U12401 (N_12401,N_6681,N_9334);
nand U12402 (N_12402,N_7539,N_8272);
nand U12403 (N_12403,N_6787,N_5011);
and U12404 (N_12404,N_8982,N_5941);
nor U12405 (N_12405,N_8840,N_7121);
nand U12406 (N_12406,N_6343,N_6344);
and U12407 (N_12407,N_9468,N_8553);
nor U12408 (N_12408,N_6120,N_5973);
or U12409 (N_12409,N_5567,N_6251);
or U12410 (N_12410,N_7820,N_5168);
nor U12411 (N_12411,N_8185,N_7744);
xor U12412 (N_12412,N_9887,N_6233);
and U12413 (N_12413,N_7701,N_6765);
and U12414 (N_12414,N_9962,N_8374);
nand U12415 (N_12415,N_7070,N_9099);
nor U12416 (N_12416,N_9814,N_5004);
and U12417 (N_12417,N_5415,N_9942);
or U12418 (N_12418,N_9471,N_7401);
nor U12419 (N_12419,N_7447,N_6818);
nor U12420 (N_12420,N_8136,N_7037);
nand U12421 (N_12421,N_8042,N_6091);
or U12422 (N_12422,N_8045,N_6393);
nor U12423 (N_12423,N_6156,N_6107);
and U12424 (N_12424,N_9163,N_5729);
or U12425 (N_12425,N_7848,N_8505);
and U12426 (N_12426,N_8519,N_5282);
and U12427 (N_12427,N_5132,N_9124);
nand U12428 (N_12428,N_8885,N_9801);
and U12429 (N_12429,N_7817,N_7468);
and U12430 (N_12430,N_6692,N_9984);
nor U12431 (N_12431,N_6287,N_7231);
and U12432 (N_12432,N_5650,N_6182);
nor U12433 (N_12433,N_5736,N_9697);
and U12434 (N_12434,N_5967,N_5648);
and U12435 (N_12435,N_8219,N_7615);
nor U12436 (N_12436,N_7319,N_6467);
or U12437 (N_12437,N_5802,N_8360);
and U12438 (N_12438,N_5076,N_6963);
and U12439 (N_12439,N_5085,N_6377);
nor U12440 (N_12440,N_6876,N_6270);
nand U12441 (N_12441,N_8225,N_6575);
nor U12442 (N_12442,N_8347,N_6893);
nor U12443 (N_12443,N_8559,N_6913);
or U12444 (N_12444,N_9557,N_9647);
nand U12445 (N_12445,N_6825,N_6958);
nor U12446 (N_12446,N_5884,N_8698);
nor U12447 (N_12447,N_5049,N_7209);
nand U12448 (N_12448,N_9696,N_9855);
and U12449 (N_12449,N_5414,N_6821);
or U12450 (N_12450,N_8995,N_6861);
and U12451 (N_12451,N_7888,N_9977);
nor U12452 (N_12452,N_9617,N_8473);
or U12453 (N_12453,N_5186,N_9018);
or U12454 (N_12454,N_8463,N_8385);
and U12455 (N_12455,N_9999,N_9589);
and U12456 (N_12456,N_7399,N_9113);
or U12457 (N_12457,N_6123,N_9597);
nor U12458 (N_12458,N_5902,N_5550);
nor U12459 (N_12459,N_9945,N_5449);
nand U12460 (N_12460,N_7914,N_9035);
and U12461 (N_12461,N_9652,N_6637);
nor U12462 (N_12462,N_5754,N_5437);
xor U12463 (N_12463,N_7904,N_8575);
nand U12464 (N_12464,N_9893,N_9657);
nand U12465 (N_12465,N_9359,N_5411);
or U12466 (N_12466,N_8821,N_9837);
nor U12467 (N_12467,N_9781,N_6292);
or U12468 (N_12468,N_9305,N_7607);
or U12469 (N_12469,N_8300,N_7657);
and U12470 (N_12470,N_6501,N_8836);
nor U12471 (N_12471,N_9384,N_8878);
nor U12472 (N_12472,N_5571,N_8973);
nor U12473 (N_12473,N_6392,N_7497);
nor U12474 (N_12474,N_8769,N_6455);
xor U12475 (N_12475,N_7433,N_9436);
or U12476 (N_12476,N_7714,N_8910);
nor U12477 (N_12477,N_6079,N_5809);
nand U12478 (N_12478,N_8256,N_5528);
nand U12479 (N_12479,N_7910,N_7706);
and U12480 (N_12480,N_8954,N_9975);
nand U12481 (N_12481,N_6285,N_6439);
and U12482 (N_12482,N_9539,N_6749);
nor U12483 (N_12483,N_7892,N_7410);
and U12484 (N_12484,N_7141,N_8204);
nor U12485 (N_12485,N_7592,N_5067);
nand U12486 (N_12486,N_7687,N_5010);
nand U12487 (N_12487,N_6139,N_7478);
and U12488 (N_12488,N_5162,N_9794);
and U12489 (N_12489,N_8333,N_9808);
xor U12490 (N_12490,N_5656,N_7082);
nand U12491 (N_12491,N_5702,N_5116);
xnor U12492 (N_12492,N_8997,N_6600);
nand U12493 (N_12493,N_7653,N_8795);
nor U12494 (N_12494,N_7240,N_5921);
nand U12495 (N_12495,N_7516,N_7957);
nor U12496 (N_12496,N_5687,N_7192);
and U12497 (N_12497,N_7471,N_6010);
nand U12498 (N_12498,N_6671,N_8461);
and U12499 (N_12499,N_8259,N_6969);
or U12500 (N_12500,N_9953,N_9157);
or U12501 (N_12501,N_8230,N_6816);
or U12502 (N_12502,N_9565,N_6780);
or U12503 (N_12503,N_6162,N_8139);
nor U12504 (N_12504,N_9811,N_7796);
nand U12505 (N_12505,N_6324,N_6034);
or U12506 (N_12506,N_5422,N_9464);
nand U12507 (N_12507,N_6092,N_5490);
nand U12508 (N_12508,N_9563,N_7505);
or U12509 (N_12509,N_5030,N_8470);
or U12510 (N_12510,N_8077,N_5255);
nand U12511 (N_12511,N_8327,N_9207);
or U12512 (N_12512,N_8037,N_9733);
nor U12513 (N_12513,N_6913,N_8223);
and U12514 (N_12514,N_9660,N_6102);
and U12515 (N_12515,N_8182,N_6839);
and U12516 (N_12516,N_7663,N_7947);
nand U12517 (N_12517,N_6853,N_7925);
nand U12518 (N_12518,N_5237,N_9745);
and U12519 (N_12519,N_6601,N_8264);
or U12520 (N_12520,N_8799,N_6223);
nor U12521 (N_12521,N_7755,N_9811);
nor U12522 (N_12522,N_9157,N_6686);
and U12523 (N_12523,N_8678,N_9680);
and U12524 (N_12524,N_5079,N_6068);
nand U12525 (N_12525,N_7113,N_8762);
and U12526 (N_12526,N_5512,N_6926);
nor U12527 (N_12527,N_9227,N_9109);
nor U12528 (N_12528,N_5684,N_8612);
nor U12529 (N_12529,N_5621,N_5159);
and U12530 (N_12530,N_8988,N_7012);
nor U12531 (N_12531,N_7726,N_8362);
nand U12532 (N_12532,N_5212,N_5817);
and U12533 (N_12533,N_7732,N_6754);
or U12534 (N_12534,N_5133,N_5488);
and U12535 (N_12535,N_6999,N_6573);
or U12536 (N_12536,N_6813,N_6607);
nor U12537 (N_12537,N_5647,N_7801);
and U12538 (N_12538,N_9739,N_9787);
or U12539 (N_12539,N_8129,N_5993);
nor U12540 (N_12540,N_5538,N_9102);
xnor U12541 (N_12541,N_7450,N_5268);
and U12542 (N_12542,N_5150,N_6613);
nand U12543 (N_12543,N_9907,N_9172);
and U12544 (N_12544,N_9429,N_8742);
or U12545 (N_12545,N_8293,N_6344);
and U12546 (N_12546,N_9955,N_8236);
nand U12547 (N_12547,N_7795,N_6709);
or U12548 (N_12548,N_7748,N_9929);
nand U12549 (N_12549,N_8870,N_7041);
nand U12550 (N_12550,N_7811,N_9756);
xor U12551 (N_12551,N_6427,N_7781);
nor U12552 (N_12552,N_7043,N_8826);
nor U12553 (N_12553,N_6251,N_6795);
or U12554 (N_12554,N_6722,N_9307);
and U12555 (N_12555,N_7264,N_5771);
and U12556 (N_12556,N_9585,N_5031);
and U12557 (N_12557,N_5666,N_6380);
xor U12558 (N_12558,N_7024,N_9148);
nand U12559 (N_12559,N_9070,N_7025);
and U12560 (N_12560,N_8283,N_8891);
and U12561 (N_12561,N_8644,N_8847);
and U12562 (N_12562,N_6722,N_7763);
nor U12563 (N_12563,N_7925,N_6226);
or U12564 (N_12564,N_8642,N_6090);
and U12565 (N_12565,N_8707,N_7276);
or U12566 (N_12566,N_5551,N_9563);
nor U12567 (N_12567,N_8053,N_6951);
nor U12568 (N_12568,N_8730,N_9250);
and U12569 (N_12569,N_7588,N_6800);
nor U12570 (N_12570,N_7722,N_7473);
and U12571 (N_12571,N_8654,N_6225);
or U12572 (N_12572,N_6153,N_6426);
nand U12573 (N_12573,N_5603,N_7423);
nand U12574 (N_12574,N_7642,N_6367);
nand U12575 (N_12575,N_8250,N_9010);
nor U12576 (N_12576,N_7873,N_8833);
or U12577 (N_12577,N_9972,N_7356);
and U12578 (N_12578,N_6760,N_9094);
nor U12579 (N_12579,N_5851,N_8554);
nor U12580 (N_12580,N_7255,N_9709);
nand U12581 (N_12581,N_8289,N_5571);
nand U12582 (N_12582,N_7995,N_8487);
and U12583 (N_12583,N_9520,N_6880);
and U12584 (N_12584,N_9138,N_7673);
nor U12585 (N_12585,N_5546,N_5060);
or U12586 (N_12586,N_8577,N_5958);
or U12587 (N_12587,N_8898,N_6055);
or U12588 (N_12588,N_9422,N_7831);
nor U12589 (N_12589,N_5885,N_9055);
or U12590 (N_12590,N_6699,N_6528);
or U12591 (N_12591,N_9248,N_9645);
and U12592 (N_12592,N_5285,N_9327);
and U12593 (N_12593,N_5206,N_6761);
and U12594 (N_12594,N_7021,N_9563);
nand U12595 (N_12595,N_8286,N_9014);
and U12596 (N_12596,N_8606,N_8365);
nand U12597 (N_12597,N_9954,N_9234);
or U12598 (N_12598,N_9873,N_8731);
and U12599 (N_12599,N_6721,N_9149);
and U12600 (N_12600,N_8508,N_9106);
and U12601 (N_12601,N_9503,N_8993);
xor U12602 (N_12602,N_5500,N_9833);
or U12603 (N_12603,N_5736,N_8052);
and U12604 (N_12604,N_6121,N_5713);
nor U12605 (N_12605,N_5024,N_8502);
nor U12606 (N_12606,N_9808,N_5400);
and U12607 (N_12607,N_6484,N_6126);
or U12608 (N_12608,N_6462,N_5321);
nor U12609 (N_12609,N_7628,N_8535);
and U12610 (N_12610,N_9976,N_6905);
nor U12611 (N_12611,N_6074,N_5768);
nand U12612 (N_12612,N_7146,N_7384);
or U12613 (N_12613,N_9387,N_5156);
and U12614 (N_12614,N_9120,N_8162);
and U12615 (N_12615,N_7051,N_7995);
nor U12616 (N_12616,N_5619,N_5314);
or U12617 (N_12617,N_6903,N_5086);
nor U12618 (N_12618,N_9706,N_9633);
and U12619 (N_12619,N_5010,N_5120);
and U12620 (N_12620,N_7599,N_7898);
or U12621 (N_12621,N_5376,N_9340);
nand U12622 (N_12622,N_5500,N_7124);
nor U12623 (N_12623,N_5933,N_7614);
and U12624 (N_12624,N_6397,N_5451);
nand U12625 (N_12625,N_9002,N_9622);
nor U12626 (N_12626,N_7630,N_9319);
nand U12627 (N_12627,N_5584,N_6125);
and U12628 (N_12628,N_7695,N_6670);
nor U12629 (N_12629,N_6592,N_9052);
or U12630 (N_12630,N_6742,N_9292);
nand U12631 (N_12631,N_5769,N_8048);
xor U12632 (N_12632,N_6656,N_9762);
or U12633 (N_12633,N_7783,N_6125);
nor U12634 (N_12634,N_6606,N_5308);
nor U12635 (N_12635,N_6476,N_9240);
or U12636 (N_12636,N_6893,N_5913);
nand U12637 (N_12637,N_5489,N_8567);
and U12638 (N_12638,N_7133,N_8655);
or U12639 (N_12639,N_9828,N_9439);
nor U12640 (N_12640,N_8615,N_7215);
or U12641 (N_12641,N_9830,N_5596);
or U12642 (N_12642,N_8172,N_5065);
nor U12643 (N_12643,N_8147,N_7048);
or U12644 (N_12644,N_5457,N_6152);
and U12645 (N_12645,N_7953,N_8998);
nand U12646 (N_12646,N_9863,N_8875);
nor U12647 (N_12647,N_6887,N_7278);
and U12648 (N_12648,N_7921,N_9336);
xor U12649 (N_12649,N_8478,N_8516);
nor U12650 (N_12650,N_6261,N_6992);
and U12651 (N_12651,N_8876,N_9102);
and U12652 (N_12652,N_7383,N_7147);
or U12653 (N_12653,N_8376,N_7400);
nor U12654 (N_12654,N_7795,N_8582);
or U12655 (N_12655,N_5984,N_9927);
and U12656 (N_12656,N_5201,N_7780);
xnor U12657 (N_12657,N_5889,N_9191);
nor U12658 (N_12658,N_8250,N_6605);
or U12659 (N_12659,N_8805,N_6604);
or U12660 (N_12660,N_8772,N_8698);
xnor U12661 (N_12661,N_7372,N_8415);
or U12662 (N_12662,N_7895,N_8398);
nor U12663 (N_12663,N_5563,N_9453);
and U12664 (N_12664,N_9212,N_8470);
nor U12665 (N_12665,N_6552,N_6925);
or U12666 (N_12666,N_8764,N_7199);
and U12667 (N_12667,N_6478,N_6121);
nand U12668 (N_12668,N_9867,N_7349);
or U12669 (N_12669,N_9247,N_8664);
and U12670 (N_12670,N_9423,N_8967);
and U12671 (N_12671,N_7865,N_7022);
or U12672 (N_12672,N_5368,N_9577);
nor U12673 (N_12673,N_7899,N_9144);
nor U12674 (N_12674,N_8366,N_7454);
or U12675 (N_12675,N_6767,N_5628);
nor U12676 (N_12676,N_8887,N_5663);
nand U12677 (N_12677,N_6094,N_5048);
and U12678 (N_12678,N_6541,N_6812);
and U12679 (N_12679,N_5689,N_9997);
nor U12680 (N_12680,N_9258,N_6710);
nand U12681 (N_12681,N_5139,N_6625);
or U12682 (N_12682,N_8620,N_6631);
nor U12683 (N_12683,N_5091,N_9366);
or U12684 (N_12684,N_9747,N_5468);
and U12685 (N_12685,N_7816,N_7111);
nand U12686 (N_12686,N_8718,N_9006);
or U12687 (N_12687,N_9879,N_7466);
nor U12688 (N_12688,N_5186,N_5371);
or U12689 (N_12689,N_9060,N_6316);
and U12690 (N_12690,N_6138,N_5906);
nand U12691 (N_12691,N_6960,N_9752);
or U12692 (N_12692,N_5836,N_5783);
nor U12693 (N_12693,N_6524,N_9275);
or U12694 (N_12694,N_6502,N_5342);
or U12695 (N_12695,N_8570,N_9989);
or U12696 (N_12696,N_7844,N_7172);
and U12697 (N_12697,N_8729,N_8809);
and U12698 (N_12698,N_8411,N_9369);
xor U12699 (N_12699,N_8924,N_5739);
and U12700 (N_12700,N_6062,N_8378);
nor U12701 (N_12701,N_9705,N_8235);
xnor U12702 (N_12702,N_9896,N_6005);
nand U12703 (N_12703,N_7899,N_6859);
nand U12704 (N_12704,N_6272,N_7863);
nand U12705 (N_12705,N_9889,N_7704);
or U12706 (N_12706,N_5467,N_5292);
or U12707 (N_12707,N_7019,N_6517);
nor U12708 (N_12708,N_5084,N_7155);
nand U12709 (N_12709,N_7027,N_5095);
or U12710 (N_12710,N_5714,N_9277);
nand U12711 (N_12711,N_5559,N_6516);
or U12712 (N_12712,N_7944,N_7788);
nand U12713 (N_12713,N_5014,N_6921);
or U12714 (N_12714,N_8332,N_6108);
nand U12715 (N_12715,N_9590,N_7381);
and U12716 (N_12716,N_7758,N_8288);
nor U12717 (N_12717,N_7261,N_7445);
or U12718 (N_12718,N_6021,N_9116);
nor U12719 (N_12719,N_7207,N_7691);
or U12720 (N_12720,N_6770,N_8211);
or U12721 (N_12721,N_7961,N_8270);
and U12722 (N_12722,N_7481,N_8125);
nor U12723 (N_12723,N_7775,N_8835);
and U12724 (N_12724,N_7948,N_8849);
nand U12725 (N_12725,N_9131,N_8399);
or U12726 (N_12726,N_9258,N_5361);
or U12727 (N_12727,N_8578,N_8307);
nor U12728 (N_12728,N_5748,N_8520);
or U12729 (N_12729,N_5547,N_7451);
nor U12730 (N_12730,N_6585,N_7479);
nand U12731 (N_12731,N_8406,N_7131);
nand U12732 (N_12732,N_9935,N_5502);
and U12733 (N_12733,N_6410,N_7325);
or U12734 (N_12734,N_8367,N_6173);
and U12735 (N_12735,N_9381,N_6928);
nand U12736 (N_12736,N_7952,N_8647);
nor U12737 (N_12737,N_8778,N_9201);
nand U12738 (N_12738,N_5697,N_7837);
nand U12739 (N_12739,N_7880,N_7507);
xnor U12740 (N_12740,N_6007,N_5223);
or U12741 (N_12741,N_8405,N_5522);
nand U12742 (N_12742,N_7618,N_6989);
nand U12743 (N_12743,N_5473,N_6784);
nor U12744 (N_12744,N_6541,N_6302);
or U12745 (N_12745,N_8856,N_7451);
or U12746 (N_12746,N_6754,N_6514);
or U12747 (N_12747,N_6608,N_7428);
nand U12748 (N_12748,N_6030,N_9787);
and U12749 (N_12749,N_5801,N_9663);
nor U12750 (N_12750,N_9118,N_9835);
nor U12751 (N_12751,N_9692,N_9255);
or U12752 (N_12752,N_7866,N_9072);
nand U12753 (N_12753,N_8487,N_5707);
nor U12754 (N_12754,N_6401,N_9748);
or U12755 (N_12755,N_7634,N_7657);
nor U12756 (N_12756,N_8443,N_6780);
and U12757 (N_12757,N_9427,N_6839);
nand U12758 (N_12758,N_6402,N_8754);
or U12759 (N_12759,N_9355,N_7007);
nand U12760 (N_12760,N_8431,N_8968);
and U12761 (N_12761,N_5446,N_6300);
nand U12762 (N_12762,N_9943,N_5626);
and U12763 (N_12763,N_8173,N_9050);
and U12764 (N_12764,N_6126,N_6062);
or U12765 (N_12765,N_6292,N_8412);
nor U12766 (N_12766,N_8942,N_7325);
xnor U12767 (N_12767,N_7830,N_6245);
and U12768 (N_12768,N_5013,N_5517);
nor U12769 (N_12769,N_8175,N_9828);
and U12770 (N_12770,N_8394,N_9677);
nor U12771 (N_12771,N_9777,N_7617);
nor U12772 (N_12772,N_7531,N_7053);
nor U12773 (N_12773,N_5605,N_6109);
and U12774 (N_12774,N_7831,N_7727);
nand U12775 (N_12775,N_5552,N_6250);
nand U12776 (N_12776,N_8081,N_6958);
and U12777 (N_12777,N_8432,N_8651);
nand U12778 (N_12778,N_7173,N_9339);
and U12779 (N_12779,N_7370,N_9262);
or U12780 (N_12780,N_7317,N_5927);
or U12781 (N_12781,N_6308,N_7485);
nand U12782 (N_12782,N_6581,N_7359);
nand U12783 (N_12783,N_5472,N_5639);
nand U12784 (N_12784,N_9509,N_7720);
nor U12785 (N_12785,N_7210,N_9263);
nand U12786 (N_12786,N_9795,N_5367);
nor U12787 (N_12787,N_6337,N_6327);
nor U12788 (N_12788,N_8254,N_7217);
or U12789 (N_12789,N_7481,N_5674);
and U12790 (N_12790,N_9509,N_6168);
nor U12791 (N_12791,N_5788,N_5970);
and U12792 (N_12792,N_5144,N_8026);
or U12793 (N_12793,N_5200,N_9100);
or U12794 (N_12794,N_8401,N_9353);
nor U12795 (N_12795,N_7387,N_5683);
and U12796 (N_12796,N_9343,N_7119);
nor U12797 (N_12797,N_8358,N_9198);
and U12798 (N_12798,N_7486,N_8861);
and U12799 (N_12799,N_8368,N_5377);
or U12800 (N_12800,N_5404,N_9702);
nand U12801 (N_12801,N_8751,N_8305);
nand U12802 (N_12802,N_9428,N_8758);
nor U12803 (N_12803,N_8235,N_8478);
and U12804 (N_12804,N_9930,N_5852);
nand U12805 (N_12805,N_5981,N_7977);
and U12806 (N_12806,N_5570,N_9351);
nor U12807 (N_12807,N_5537,N_6249);
nor U12808 (N_12808,N_6581,N_7592);
and U12809 (N_12809,N_9161,N_9687);
or U12810 (N_12810,N_7575,N_6696);
or U12811 (N_12811,N_9403,N_9378);
or U12812 (N_12812,N_6009,N_8768);
nor U12813 (N_12813,N_7151,N_9934);
nand U12814 (N_12814,N_8506,N_8832);
and U12815 (N_12815,N_7284,N_8753);
or U12816 (N_12816,N_8780,N_8694);
and U12817 (N_12817,N_9351,N_8639);
and U12818 (N_12818,N_9982,N_6423);
or U12819 (N_12819,N_7947,N_8886);
and U12820 (N_12820,N_6352,N_5084);
nand U12821 (N_12821,N_9215,N_5993);
or U12822 (N_12822,N_5649,N_7166);
and U12823 (N_12823,N_8288,N_5155);
xnor U12824 (N_12824,N_6617,N_7297);
nand U12825 (N_12825,N_8329,N_5689);
or U12826 (N_12826,N_8329,N_8651);
nor U12827 (N_12827,N_7300,N_6655);
nor U12828 (N_12828,N_9240,N_6157);
or U12829 (N_12829,N_6561,N_7784);
nor U12830 (N_12830,N_6011,N_8629);
or U12831 (N_12831,N_6531,N_5550);
nor U12832 (N_12832,N_6625,N_5044);
nor U12833 (N_12833,N_8016,N_6724);
or U12834 (N_12834,N_5005,N_6483);
and U12835 (N_12835,N_9500,N_6726);
xnor U12836 (N_12836,N_7788,N_8839);
and U12837 (N_12837,N_6039,N_6371);
and U12838 (N_12838,N_8297,N_8520);
nor U12839 (N_12839,N_5472,N_9579);
and U12840 (N_12840,N_7776,N_7161);
and U12841 (N_12841,N_8105,N_6905);
nand U12842 (N_12842,N_9036,N_9201);
nor U12843 (N_12843,N_9068,N_7826);
and U12844 (N_12844,N_6101,N_7689);
and U12845 (N_12845,N_8894,N_8151);
or U12846 (N_12846,N_8058,N_8945);
or U12847 (N_12847,N_6357,N_6436);
and U12848 (N_12848,N_8765,N_6385);
nor U12849 (N_12849,N_6415,N_9123);
and U12850 (N_12850,N_7538,N_7641);
xnor U12851 (N_12851,N_7242,N_5366);
nor U12852 (N_12852,N_8454,N_7167);
and U12853 (N_12853,N_7513,N_6269);
and U12854 (N_12854,N_5339,N_8366);
and U12855 (N_12855,N_9833,N_6809);
or U12856 (N_12856,N_5002,N_9384);
nand U12857 (N_12857,N_7861,N_8188);
and U12858 (N_12858,N_5244,N_5537);
nand U12859 (N_12859,N_5758,N_8258);
and U12860 (N_12860,N_8174,N_9174);
or U12861 (N_12861,N_9600,N_5975);
and U12862 (N_12862,N_8832,N_9815);
or U12863 (N_12863,N_8208,N_7583);
or U12864 (N_12864,N_9046,N_9065);
nor U12865 (N_12865,N_9401,N_9271);
nor U12866 (N_12866,N_9822,N_9696);
or U12867 (N_12867,N_9933,N_9694);
nand U12868 (N_12868,N_5285,N_7732);
or U12869 (N_12869,N_9789,N_9878);
xor U12870 (N_12870,N_5465,N_8389);
and U12871 (N_12871,N_7542,N_5751);
nand U12872 (N_12872,N_6295,N_8682);
or U12873 (N_12873,N_9439,N_9536);
nand U12874 (N_12874,N_5523,N_7595);
or U12875 (N_12875,N_5243,N_5268);
nand U12876 (N_12876,N_7467,N_5605);
and U12877 (N_12877,N_8576,N_6273);
xor U12878 (N_12878,N_5369,N_8279);
or U12879 (N_12879,N_5348,N_9163);
nand U12880 (N_12880,N_7972,N_7864);
or U12881 (N_12881,N_5040,N_8649);
nand U12882 (N_12882,N_7497,N_6003);
and U12883 (N_12883,N_5007,N_8466);
or U12884 (N_12884,N_7771,N_8356);
nand U12885 (N_12885,N_8738,N_8000);
nand U12886 (N_12886,N_7173,N_7972);
nor U12887 (N_12887,N_6954,N_5663);
or U12888 (N_12888,N_7200,N_6493);
nand U12889 (N_12889,N_9929,N_9859);
or U12890 (N_12890,N_6227,N_7292);
and U12891 (N_12891,N_8173,N_9662);
or U12892 (N_12892,N_9847,N_6830);
nor U12893 (N_12893,N_6149,N_8348);
and U12894 (N_12894,N_7950,N_5961);
and U12895 (N_12895,N_8557,N_8035);
nand U12896 (N_12896,N_8916,N_5917);
and U12897 (N_12897,N_9644,N_8864);
nand U12898 (N_12898,N_8174,N_9718);
nand U12899 (N_12899,N_9589,N_5719);
nand U12900 (N_12900,N_7324,N_5725);
nand U12901 (N_12901,N_6669,N_6954);
or U12902 (N_12902,N_6215,N_8088);
nor U12903 (N_12903,N_6743,N_8629);
nand U12904 (N_12904,N_8402,N_8241);
nor U12905 (N_12905,N_8149,N_7681);
nor U12906 (N_12906,N_8729,N_9862);
or U12907 (N_12907,N_6844,N_7807);
nand U12908 (N_12908,N_5106,N_7417);
and U12909 (N_12909,N_9281,N_7329);
nand U12910 (N_12910,N_9286,N_6737);
nand U12911 (N_12911,N_7235,N_7555);
or U12912 (N_12912,N_6254,N_9349);
nand U12913 (N_12913,N_9063,N_9265);
or U12914 (N_12914,N_9844,N_6185);
nand U12915 (N_12915,N_7456,N_6922);
nand U12916 (N_12916,N_6792,N_9131);
nor U12917 (N_12917,N_8063,N_6085);
or U12918 (N_12918,N_9234,N_8139);
xor U12919 (N_12919,N_7432,N_8559);
nand U12920 (N_12920,N_8548,N_5792);
or U12921 (N_12921,N_9571,N_6704);
nor U12922 (N_12922,N_5575,N_5886);
nor U12923 (N_12923,N_6881,N_5444);
or U12924 (N_12924,N_6466,N_9227);
nor U12925 (N_12925,N_9347,N_6995);
nor U12926 (N_12926,N_9537,N_6589);
and U12927 (N_12927,N_8563,N_9962);
or U12928 (N_12928,N_6430,N_7975);
or U12929 (N_12929,N_5817,N_7199);
or U12930 (N_12930,N_7165,N_8315);
and U12931 (N_12931,N_5681,N_5100);
or U12932 (N_12932,N_5414,N_8887);
nand U12933 (N_12933,N_8638,N_6990);
and U12934 (N_12934,N_9126,N_8956);
and U12935 (N_12935,N_6552,N_6170);
xnor U12936 (N_12936,N_5346,N_9473);
nor U12937 (N_12937,N_6229,N_7550);
and U12938 (N_12938,N_6309,N_8770);
nand U12939 (N_12939,N_9436,N_9281);
or U12940 (N_12940,N_5555,N_6923);
or U12941 (N_12941,N_6882,N_8297);
or U12942 (N_12942,N_9452,N_7276);
nand U12943 (N_12943,N_9889,N_9891);
and U12944 (N_12944,N_9816,N_9294);
or U12945 (N_12945,N_7240,N_6727);
and U12946 (N_12946,N_5201,N_6824);
nor U12947 (N_12947,N_6921,N_5200);
and U12948 (N_12948,N_6516,N_9749);
nand U12949 (N_12949,N_7458,N_5423);
and U12950 (N_12950,N_6464,N_7849);
nor U12951 (N_12951,N_6117,N_9465);
nor U12952 (N_12952,N_6266,N_9150);
and U12953 (N_12953,N_7658,N_8426);
or U12954 (N_12954,N_7238,N_6453);
nor U12955 (N_12955,N_5288,N_7980);
nor U12956 (N_12956,N_6941,N_5907);
or U12957 (N_12957,N_9219,N_7084);
nor U12958 (N_12958,N_9466,N_6419);
or U12959 (N_12959,N_9561,N_7094);
and U12960 (N_12960,N_6564,N_7349);
or U12961 (N_12961,N_5898,N_6389);
or U12962 (N_12962,N_5448,N_7433);
nand U12963 (N_12963,N_7191,N_7541);
nand U12964 (N_12964,N_9511,N_6773);
and U12965 (N_12965,N_7244,N_7695);
or U12966 (N_12966,N_9415,N_8578);
or U12967 (N_12967,N_5480,N_9545);
xor U12968 (N_12968,N_6333,N_8053);
nand U12969 (N_12969,N_8146,N_8177);
nor U12970 (N_12970,N_9663,N_8324);
nand U12971 (N_12971,N_8149,N_5966);
nand U12972 (N_12972,N_8865,N_9606);
nor U12973 (N_12973,N_5706,N_7037);
nand U12974 (N_12974,N_8834,N_7676);
or U12975 (N_12975,N_5642,N_7639);
and U12976 (N_12976,N_8264,N_9301);
and U12977 (N_12977,N_6288,N_5416);
and U12978 (N_12978,N_6113,N_7742);
and U12979 (N_12979,N_8962,N_9865);
nand U12980 (N_12980,N_5853,N_6887);
or U12981 (N_12981,N_5150,N_8411);
or U12982 (N_12982,N_7127,N_7573);
and U12983 (N_12983,N_7614,N_9069);
and U12984 (N_12984,N_8139,N_7288);
or U12985 (N_12985,N_7006,N_6036);
nor U12986 (N_12986,N_9105,N_7135);
nor U12987 (N_12987,N_7964,N_8557);
nand U12988 (N_12988,N_6302,N_5837);
nand U12989 (N_12989,N_8113,N_5993);
nor U12990 (N_12990,N_8333,N_5774);
or U12991 (N_12991,N_5165,N_7161);
and U12992 (N_12992,N_7421,N_9324);
and U12993 (N_12993,N_7554,N_7610);
or U12994 (N_12994,N_9554,N_9016);
nand U12995 (N_12995,N_9013,N_9884);
or U12996 (N_12996,N_7212,N_9582);
nand U12997 (N_12997,N_6395,N_6980);
nand U12998 (N_12998,N_5176,N_8559);
or U12999 (N_12999,N_7949,N_6020);
and U13000 (N_13000,N_7310,N_9861);
nand U13001 (N_13001,N_9737,N_8213);
and U13002 (N_13002,N_7335,N_6961);
or U13003 (N_13003,N_7922,N_9154);
nor U13004 (N_13004,N_6515,N_6353);
nand U13005 (N_13005,N_6817,N_9015);
xor U13006 (N_13006,N_9911,N_7272);
or U13007 (N_13007,N_7498,N_8885);
nand U13008 (N_13008,N_6890,N_8859);
and U13009 (N_13009,N_5094,N_7961);
nand U13010 (N_13010,N_9489,N_6514);
nor U13011 (N_13011,N_8377,N_5631);
or U13012 (N_13012,N_6273,N_5527);
or U13013 (N_13013,N_6577,N_7064);
and U13014 (N_13014,N_9891,N_5331);
nand U13015 (N_13015,N_7375,N_7869);
or U13016 (N_13016,N_6566,N_8121);
nand U13017 (N_13017,N_7273,N_8811);
or U13018 (N_13018,N_6096,N_6826);
nor U13019 (N_13019,N_9980,N_6654);
or U13020 (N_13020,N_6856,N_8217);
nor U13021 (N_13021,N_8377,N_7323);
nand U13022 (N_13022,N_9762,N_8743);
nand U13023 (N_13023,N_5182,N_6575);
nor U13024 (N_13024,N_7249,N_7498);
or U13025 (N_13025,N_6192,N_9359);
nor U13026 (N_13026,N_6009,N_6774);
nand U13027 (N_13027,N_8885,N_7250);
or U13028 (N_13028,N_8190,N_6292);
nand U13029 (N_13029,N_5521,N_6532);
nand U13030 (N_13030,N_9598,N_5050);
or U13031 (N_13031,N_9607,N_6538);
and U13032 (N_13032,N_7838,N_7955);
or U13033 (N_13033,N_7511,N_7292);
or U13034 (N_13034,N_8032,N_6494);
and U13035 (N_13035,N_7525,N_9945);
nand U13036 (N_13036,N_9430,N_5951);
and U13037 (N_13037,N_8070,N_8196);
nor U13038 (N_13038,N_7394,N_6201);
and U13039 (N_13039,N_8864,N_6854);
nor U13040 (N_13040,N_6763,N_8597);
and U13041 (N_13041,N_5933,N_7393);
nor U13042 (N_13042,N_5930,N_8349);
and U13043 (N_13043,N_8798,N_6165);
or U13044 (N_13044,N_5756,N_8618);
and U13045 (N_13045,N_6511,N_7777);
nor U13046 (N_13046,N_7798,N_5462);
and U13047 (N_13047,N_7647,N_6365);
and U13048 (N_13048,N_5653,N_5960);
nand U13049 (N_13049,N_8744,N_7845);
nand U13050 (N_13050,N_5716,N_6773);
and U13051 (N_13051,N_6305,N_7208);
and U13052 (N_13052,N_6006,N_7453);
xnor U13053 (N_13053,N_7379,N_7367);
nand U13054 (N_13054,N_5689,N_8950);
or U13055 (N_13055,N_5196,N_6325);
nand U13056 (N_13056,N_5980,N_6025);
and U13057 (N_13057,N_5520,N_6148);
and U13058 (N_13058,N_7340,N_8289);
or U13059 (N_13059,N_7917,N_5389);
or U13060 (N_13060,N_9279,N_9886);
nor U13061 (N_13061,N_6532,N_5234);
nor U13062 (N_13062,N_5350,N_7405);
nand U13063 (N_13063,N_6587,N_9027);
nand U13064 (N_13064,N_8563,N_7565);
and U13065 (N_13065,N_7200,N_9863);
nand U13066 (N_13066,N_8571,N_7384);
or U13067 (N_13067,N_7932,N_7891);
and U13068 (N_13068,N_8456,N_7817);
and U13069 (N_13069,N_8358,N_7729);
and U13070 (N_13070,N_5647,N_8731);
nand U13071 (N_13071,N_9526,N_7049);
nor U13072 (N_13072,N_7752,N_9412);
or U13073 (N_13073,N_8990,N_6572);
xnor U13074 (N_13074,N_8641,N_5913);
and U13075 (N_13075,N_7143,N_9827);
nor U13076 (N_13076,N_6654,N_5823);
nor U13077 (N_13077,N_7536,N_5355);
and U13078 (N_13078,N_7365,N_6714);
and U13079 (N_13079,N_9423,N_6911);
and U13080 (N_13080,N_6913,N_5608);
nand U13081 (N_13081,N_5077,N_5203);
xnor U13082 (N_13082,N_7153,N_7884);
nor U13083 (N_13083,N_9432,N_9929);
nand U13084 (N_13084,N_5588,N_5239);
nand U13085 (N_13085,N_7827,N_8496);
nand U13086 (N_13086,N_6052,N_8860);
nor U13087 (N_13087,N_5735,N_9020);
nand U13088 (N_13088,N_5809,N_5190);
nor U13089 (N_13089,N_8976,N_7676);
or U13090 (N_13090,N_7632,N_6874);
nor U13091 (N_13091,N_7005,N_8615);
or U13092 (N_13092,N_9516,N_7080);
xor U13093 (N_13093,N_6262,N_9488);
xor U13094 (N_13094,N_6123,N_5879);
or U13095 (N_13095,N_6490,N_7154);
or U13096 (N_13096,N_5732,N_7567);
nand U13097 (N_13097,N_7914,N_9839);
or U13098 (N_13098,N_5772,N_5227);
nand U13099 (N_13099,N_5115,N_8641);
or U13100 (N_13100,N_6881,N_8912);
xor U13101 (N_13101,N_5198,N_9819);
nand U13102 (N_13102,N_7431,N_7755);
nand U13103 (N_13103,N_7742,N_5070);
nor U13104 (N_13104,N_5250,N_6496);
nor U13105 (N_13105,N_6499,N_7902);
and U13106 (N_13106,N_7936,N_9421);
nand U13107 (N_13107,N_6172,N_9424);
nor U13108 (N_13108,N_6902,N_7956);
and U13109 (N_13109,N_9928,N_6741);
nand U13110 (N_13110,N_6239,N_6997);
and U13111 (N_13111,N_6682,N_7952);
nor U13112 (N_13112,N_9639,N_7952);
nand U13113 (N_13113,N_8441,N_9050);
nor U13114 (N_13114,N_8912,N_8565);
or U13115 (N_13115,N_9316,N_8973);
nor U13116 (N_13116,N_5948,N_5610);
and U13117 (N_13117,N_5772,N_9396);
nor U13118 (N_13118,N_7858,N_5361);
nand U13119 (N_13119,N_5672,N_6694);
nor U13120 (N_13120,N_9213,N_8503);
and U13121 (N_13121,N_6684,N_9955);
nand U13122 (N_13122,N_8599,N_7394);
nor U13123 (N_13123,N_9381,N_8199);
nor U13124 (N_13124,N_5077,N_7779);
nor U13125 (N_13125,N_6473,N_5077);
and U13126 (N_13126,N_8585,N_7540);
nor U13127 (N_13127,N_6271,N_5978);
nor U13128 (N_13128,N_8558,N_6121);
or U13129 (N_13129,N_9036,N_5383);
and U13130 (N_13130,N_6874,N_9049);
nor U13131 (N_13131,N_5950,N_5453);
nor U13132 (N_13132,N_6997,N_7015);
nor U13133 (N_13133,N_8181,N_7416);
and U13134 (N_13134,N_7073,N_9442);
nor U13135 (N_13135,N_9563,N_7496);
nor U13136 (N_13136,N_8259,N_6487);
nand U13137 (N_13137,N_5363,N_5781);
nand U13138 (N_13138,N_7337,N_5173);
and U13139 (N_13139,N_9829,N_6243);
nand U13140 (N_13140,N_5227,N_5630);
nand U13141 (N_13141,N_7090,N_6875);
nand U13142 (N_13142,N_6411,N_8470);
nand U13143 (N_13143,N_5359,N_6916);
nor U13144 (N_13144,N_5520,N_6654);
nand U13145 (N_13145,N_7422,N_5137);
or U13146 (N_13146,N_7548,N_8414);
and U13147 (N_13147,N_7337,N_8677);
nand U13148 (N_13148,N_6014,N_5261);
or U13149 (N_13149,N_9825,N_8331);
and U13150 (N_13150,N_7959,N_9119);
nand U13151 (N_13151,N_7193,N_8941);
nor U13152 (N_13152,N_7640,N_6177);
and U13153 (N_13153,N_7324,N_6701);
or U13154 (N_13154,N_7594,N_5527);
or U13155 (N_13155,N_8593,N_8563);
nand U13156 (N_13156,N_9741,N_9479);
nand U13157 (N_13157,N_9579,N_7349);
and U13158 (N_13158,N_8562,N_8800);
nand U13159 (N_13159,N_5853,N_6424);
or U13160 (N_13160,N_5180,N_9815);
nand U13161 (N_13161,N_8589,N_6910);
nor U13162 (N_13162,N_5721,N_8818);
and U13163 (N_13163,N_5397,N_9103);
or U13164 (N_13164,N_7476,N_6756);
and U13165 (N_13165,N_5816,N_8100);
nand U13166 (N_13166,N_9562,N_7607);
nand U13167 (N_13167,N_7357,N_9299);
nand U13168 (N_13168,N_9688,N_6336);
or U13169 (N_13169,N_8925,N_7018);
and U13170 (N_13170,N_7512,N_7515);
or U13171 (N_13171,N_6716,N_9831);
and U13172 (N_13172,N_9105,N_5264);
or U13173 (N_13173,N_9035,N_7380);
nand U13174 (N_13174,N_7279,N_5765);
or U13175 (N_13175,N_5001,N_5847);
nor U13176 (N_13176,N_9008,N_6485);
nor U13177 (N_13177,N_7344,N_7110);
nand U13178 (N_13178,N_6813,N_8032);
and U13179 (N_13179,N_5844,N_8849);
nor U13180 (N_13180,N_7777,N_5303);
nor U13181 (N_13181,N_6998,N_9927);
or U13182 (N_13182,N_6104,N_5514);
nand U13183 (N_13183,N_5899,N_9910);
or U13184 (N_13184,N_5231,N_6367);
and U13185 (N_13185,N_9962,N_6169);
nor U13186 (N_13186,N_6690,N_9168);
nand U13187 (N_13187,N_9082,N_6827);
nor U13188 (N_13188,N_9453,N_8175);
nor U13189 (N_13189,N_7627,N_5178);
nand U13190 (N_13190,N_8249,N_7923);
nand U13191 (N_13191,N_6240,N_9276);
or U13192 (N_13192,N_6361,N_7356);
nor U13193 (N_13193,N_8550,N_6750);
nor U13194 (N_13194,N_9505,N_8069);
nand U13195 (N_13195,N_5034,N_9543);
nor U13196 (N_13196,N_7094,N_7962);
or U13197 (N_13197,N_5542,N_9648);
nand U13198 (N_13198,N_8719,N_6362);
and U13199 (N_13199,N_9968,N_8568);
nor U13200 (N_13200,N_7036,N_5414);
nand U13201 (N_13201,N_5837,N_7497);
nor U13202 (N_13202,N_7554,N_5092);
nor U13203 (N_13203,N_5961,N_8175);
and U13204 (N_13204,N_9953,N_5435);
nand U13205 (N_13205,N_7751,N_5461);
and U13206 (N_13206,N_8206,N_7333);
nand U13207 (N_13207,N_9761,N_5595);
nand U13208 (N_13208,N_9118,N_6228);
nand U13209 (N_13209,N_5425,N_5524);
or U13210 (N_13210,N_6597,N_6877);
or U13211 (N_13211,N_5047,N_7580);
nand U13212 (N_13212,N_9999,N_7806);
or U13213 (N_13213,N_6807,N_5417);
nor U13214 (N_13214,N_7924,N_7960);
nand U13215 (N_13215,N_8938,N_9762);
nor U13216 (N_13216,N_8176,N_8811);
and U13217 (N_13217,N_5918,N_6935);
nor U13218 (N_13218,N_7968,N_6666);
nand U13219 (N_13219,N_6819,N_9297);
and U13220 (N_13220,N_9943,N_6805);
or U13221 (N_13221,N_5932,N_5010);
nor U13222 (N_13222,N_8643,N_5402);
nand U13223 (N_13223,N_6101,N_5201);
nor U13224 (N_13224,N_6927,N_6513);
or U13225 (N_13225,N_7928,N_5287);
or U13226 (N_13226,N_9513,N_9802);
and U13227 (N_13227,N_5560,N_9370);
nor U13228 (N_13228,N_6650,N_8301);
nor U13229 (N_13229,N_8837,N_9678);
nand U13230 (N_13230,N_6527,N_9665);
and U13231 (N_13231,N_5828,N_5868);
or U13232 (N_13232,N_9528,N_9976);
or U13233 (N_13233,N_9113,N_5001);
nand U13234 (N_13234,N_9657,N_9555);
or U13235 (N_13235,N_8226,N_8732);
nand U13236 (N_13236,N_7927,N_9338);
or U13237 (N_13237,N_5521,N_6257);
and U13238 (N_13238,N_6085,N_7594);
and U13239 (N_13239,N_7905,N_9152);
or U13240 (N_13240,N_7279,N_9298);
nand U13241 (N_13241,N_8759,N_9723);
xnor U13242 (N_13242,N_7001,N_7699);
and U13243 (N_13243,N_7980,N_5628);
and U13244 (N_13244,N_6691,N_9371);
or U13245 (N_13245,N_6539,N_9199);
or U13246 (N_13246,N_8246,N_9579);
nor U13247 (N_13247,N_5946,N_8821);
or U13248 (N_13248,N_9426,N_9505);
nand U13249 (N_13249,N_5109,N_6590);
or U13250 (N_13250,N_9718,N_8388);
and U13251 (N_13251,N_9113,N_7123);
nor U13252 (N_13252,N_5812,N_6726);
or U13253 (N_13253,N_8716,N_6880);
or U13254 (N_13254,N_7824,N_9773);
and U13255 (N_13255,N_7454,N_7029);
and U13256 (N_13256,N_7063,N_7321);
nor U13257 (N_13257,N_6353,N_7846);
nor U13258 (N_13258,N_5545,N_5349);
or U13259 (N_13259,N_8135,N_8420);
or U13260 (N_13260,N_8444,N_9792);
and U13261 (N_13261,N_7090,N_6108);
nand U13262 (N_13262,N_9404,N_7169);
nand U13263 (N_13263,N_9759,N_7768);
nor U13264 (N_13264,N_8608,N_8492);
nor U13265 (N_13265,N_7932,N_8958);
nor U13266 (N_13266,N_9403,N_6043);
nand U13267 (N_13267,N_9117,N_8674);
nand U13268 (N_13268,N_9850,N_8096);
or U13269 (N_13269,N_8405,N_6683);
nand U13270 (N_13270,N_9444,N_9646);
nand U13271 (N_13271,N_5575,N_8319);
nand U13272 (N_13272,N_8579,N_6686);
xor U13273 (N_13273,N_9322,N_6486);
nor U13274 (N_13274,N_9904,N_9367);
or U13275 (N_13275,N_6579,N_9902);
nor U13276 (N_13276,N_8726,N_9982);
nor U13277 (N_13277,N_6996,N_8267);
nor U13278 (N_13278,N_5400,N_8296);
nor U13279 (N_13279,N_9285,N_8516);
or U13280 (N_13280,N_9730,N_8008);
nor U13281 (N_13281,N_8682,N_6898);
and U13282 (N_13282,N_6416,N_8707);
nor U13283 (N_13283,N_5873,N_5576);
or U13284 (N_13284,N_9328,N_6797);
or U13285 (N_13285,N_7097,N_9426);
nand U13286 (N_13286,N_8876,N_5419);
nand U13287 (N_13287,N_8687,N_8353);
and U13288 (N_13288,N_8468,N_7892);
or U13289 (N_13289,N_5555,N_9339);
nand U13290 (N_13290,N_9277,N_9942);
nor U13291 (N_13291,N_5909,N_9117);
nor U13292 (N_13292,N_7458,N_5146);
or U13293 (N_13293,N_8116,N_5205);
nand U13294 (N_13294,N_5103,N_9106);
or U13295 (N_13295,N_7776,N_9950);
nor U13296 (N_13296,N_7264,N_5302);
and U13297 (N_13297,N_6025,N_5233);
and U13298 (N_13298,N_9386,N_5481);
nor U13299 (N_13299,N_8860,N_7157);
and U13300 (N_13300,N_9208,N_6958);
nor U13301 (N_13301,N_6526,N_8205);
and U13302 (N_13302,N_7937,N_7750);
nand U13303 (N_13303,N_7184,N_9210);
and U13304 (N_13304,N_6932,N_5627);
and U13305 (N_13305,N_6045,N_6259);
nor U13306 (N_13306,N_6445,N_8772);
nor U13307 (N_13307,N_7102,N_9848);
nor U13308 (N_13308,N_7558,N_5797);
nor U13309 (N_13309,N_6032,N_8583);
or U13310 (N_13310,N_8235,N_7264);
and U13311 (N_13311,N_7383,N_6054);
nor U13312 (N_13312,N_5762,N_7920);
and U13313 (N_13313,N_9682,N_6947);
nor U13314 (N_13314,N_8853,N_7412);
and U13315 (N_13315,N_9275,N_6862);
nand U13316 (N_13316,N_6814,N_5422);
nor U13317 (N_13317,N_6288,N_6430);
xor U13318 (N_13318,N_5913,N_8806);
nor U13319 (N_13319,N_7680,N_8912);
nor U13320 (N_13320,N_9885,N_7364);
nand U13321 (N_13321,N_8958,N_9491);
nand U13322 (N_13322,N_8175,N_6007);
nor U13323 (N_13323,N_6544,N_5718);
or U13324 (N_13324,N_7941,N_8030);
or U13325 (N_13325,N_9724,N_6059);
and U13326 (N_13326,N_8627,N_5005);
nand U13327 (N_13327,N_9848,N_7550);
or U13328 (N_13328,N_8980,N_5952);
nand U13329 (N_13329,N_9086,N_8443);
nand U13330 (N_13330,N_7603,N_9521);
nand U13331 (N_13331,N_6411,N_5753);
or U13332 (N_13332,N_6215,N_9702);
or U13333 (N_13333,N_7052,N_6271);
nor U13334 (N_13334,N_8739,N_5460);
nor U13335 (N_13335,N_9119,N_8584);
nor U13336 (N_13336,N_8382,N_6665);
and U13337 (N_13337,N_8818,N_9445);
or U13338 (N_13338,N_8476,N_9108);
nand U13339 (N_13339,N_6121,N_7567);
nand U13340 (N_13340,N_5598,N_5088);
or U13341 (N_13341,N_6844,N_6373);
nor U13342 (N_13342,N_8118,N_9242);
and U13343 (N_13343,N_5498,N_7365);
nand U13344 (N_13344,N_9649,N_5850);
and U13345 (N_13345,N_7481,N_5775);
or U13346 (N_13346,N_8860,N_8755);
or U13347 (N_13347,N_8288,N_8342);
or U13348 (N_13348,N_8607,N_5575);
and U13349 (N_13349,N_5373,N_7550);
nand U13350 (N_13350,N_5183,N_5851);
nor U13351 (N_13351,N_9687,N_5951);
nand U13352 (N_13352,N_8891,N_8539);
nor U13353 (N_13353,N_9030,N_9625);
or U13354 (N_13354,N_5450,N_9495);
nor U13355 (N_13355,N_8538,N_6572);
or U13356 (N_13356,N_7857,N_5882);
or U13357 (N_13357,N_7270,N_6415);
nor U13358 (N_13358,N_7867,N_7539);
or U13359 (N_13359,N_7699,N_7718);
nand U13360 (N_13360,N_8921,N_6369);
nand U13361 (N_13361,N_6778,N_7776);
xor U13362 (N_13362,N_7800,N_8142);
and U13363 (N_13363,N_5063,N_7423);
nand U13364 (N_13364,N_9408,N_9687);
nand U13365 (N_13365,N_9598,N_8054);
or U13366 (N_13366,N_5135,N_6731);
nor U13367 (N_13367,N_9692,N_5752);
and U13368 (N_13368,N_6482,N_6755);
xnor U13369 (N_13369,N_6283,N_8821);
and U13370 (N_13370,N_9896,N_7273);
nand U13371 (N_13371,N_9038,N_9970);
nor U13372 (N_13372,N_6470,N_7276);
nand U13373 (N_13373,N_5244,N_7296);
or U13374 (N_13374,N_8338,N_9467);
nor U13375 (N_13375,N_5837,N_7679);
nor U13376 (N_13376,N_7405,N_7780);
nor U13377 (N_13377,N_6416,N_7310);
nand U13378 (N_13378,N_6058,N_9644);
or U13379 (N_13379,N_6998,N_7270);
and U13380 (N_13380,N_9999,N_7711);
nand U13381 (N_13381,N_8572,N_5608);
or U13382 (N_13382,N_9087,N_9941);
and U13383 (N_13383,N_5651,N_6080);
and U13384 (N_13384,N_9362,N_9068);
nand U13385 (N_13385,N_6904,N_8759);
or U13386 (N_13386,N_6943,N_6549);
nor U13387 (N_13387,N_7383,N_9795);
and U13388 (N_13388,N_5943,N_9644);
nand U13389 (N_13389,N_9677,N_9305);
and U13390 (N_13390,N_7590,N_6500);
and U13391 (N_13391,N_5944,N_5025);
and U13392 (N_13392,N_7235,N_5386);
and U13393 (N_13393,N_9114,N_8529);
and U13394 (N_13394,N_5949,N_9108);
nand U13395 (N_13395,N_7164,N_7614);
nand U13396 (N_13396,N_7511,N_7443);
and U13397 (N_13397,N_5792,N_8830);
and U13398 (N_13398,N_8788,N_8765);
nand U13399 (N_13399,N_7247,N_9392);
nand U13400 (N_13400,N_8921,N_7991);
and U13401 (N_13401,N_6382,N_5810);
and U13402 (N_13402,N_7289,N_8282);
nand U13403 (N_13403,N_7956,N_6624);
and U13404 (N_13404,N_8551,N_7188);
and U13405 (N_13405,N_6468,N_9404);
nor U13406 (N_13406,N_9021,N_5982);
or U13407 (N_13407,N_9383,N_8591);
and U13408 (N_13408,N_7800,N_5948);
nand U13409 (N_13409,N_5031,N_8664);
or U13410 (N_13410,N_9330,N_5820);
or U13411 (N_13411,N_5116,N_7832);
or U13412 (N_13412,N_5677,N_8765);
or U13413 (N_13413,N_5370,N_6889);
nor U13414 (N_13414,N_5600,N_8593);
or U13415 (N_13415,N_9567,N_6682);
or U13416 (N_13416,N_8343,N_6985);
nand U13417 (N_13417,N_6544,N_5921);
or U13418 (N_13418,N_8745,N_7861);
or U13419 (N_13419,N_9049,N_8201);
and U13420 (N_13420,N_6336,N_9079);
and U13421 (N_13421,N_7745,N_7417);
and U13422 (N_13422,N_8733,N_7426);
nor U13423 (N_13423,N_6760,N_5353);
nor U13424 (N_13424,N_9002,N_8043);
nor U13425 (N_13425,N_5155,N_6999);
or U13426 (N_13426,N_7774,N_7964);
or U13427 (N_13427,N_9774,N_5387);
or U13428 (N_13428,N_7929,N_7022);
and U13429 (N_13429,N_8697,N_8170);
and U13430 (N_13430,N_9040,N_9889);
nand U13431 (N_13431,N_6937,N_5672);
or U13432 (N_13432,N_6516,N_6491);
nor U13433 (N_13433,N_7172,N_6355);
or U13434 (N_13434,N_8499,N_9262);
or U13435 (N_13435,N_7787,N_8490);
nor U13436 (N_13436,N_7909,N_7407);
or U13437 (N_13437,N_6387,N_6196);
and U13438 (N_13438,N_7550,N_5213);
and U13439 (N_13439,N_6965,N_5252);
nor U13440 (N_13440,N_8573,N_9276);
nor U13441 (N_13441,N_9302,N_6713);
and U13442 (N_13442,N_5604,N_5546);
and U13443 (N_13443,N_7047,N_6933);
or U13444 (N_13444,N_9673,N_6621);
and U13445 (N_13445,N_5483,N_8033);
or U13446 (N_13446,N_7524,N_7954);
nand U13447 (N_13447,N_6983,N_8573);
nand U13448 (N_13448,N_8916,N_8341);
nor U13449 (N_13449,N_8020,N_9986);
nor U13450 (N_13450,N_7440,N_6310);
nor U13451 (N_13451,N_6702,N_7052);
nand U13452 (N_13452,N_7789,N_6682);
nor U13453 (N_13453,N_6558,N_8935);
nand U13454 (N_13454,N_6976,N_7531);
or U13455 (N_13455,N_8012,N_8403);
and U13456 (N_13456,N_7818,N_6326);
and U13457 (N_13457,N_6085,N_6276);
and U13458 (N_13458,N_5723,N_9785);
and U13459 (N_13459,N_5396,N_7690);
xnor U13460 (N_13460,N_9121,N_9420);
nor U13461 (N_13461,N_8579,N_8179);
xnor U13462 (N_13462,N_9429,N_7798);
nand U13463 (N_13463,N_9856,N_6286);
and U13464 (N_13464,N_8084,N_6206);
nor U13465 (N_13465,N_8588,N_6316);
nor U13466 (N_13466,N_7701,N_8010);
nor U13467 (N_13467,N_7960,N_9994);
nand U13468 (N_13468,N_5554,N_9219);
or U13469 (N_13469,N_9215,N_9367);
and U13470 (N_13470,N_5459,N_7938);
and U13471 (N_13471,N_7508,N_6123);
nor U13472 (N_13472,N_7907,N_8846);
or U13473 (N_13473,N_8554,N_6641);
or U13474 (N_13474,N_6971,N_8442);
or U13475 (N_13475,N_6668,N_7909);
and U13476 (N_13476,N_5968,N_7783);
or U13477 (N_13477,N_5514,N_5270);
or U13478 (N_13478,N_8479,N_7164);
nand U13479 (N_13479,N_5620,N_6363);
or U13480 (N_13480,N_5383,N_5435);
or U13481 (N_13481,N_5394,N_5850);
nor U13482 (N_13482,N_7581,N_7401);
or U13483 (N_13483,N_8442,N_6825);
nand U13484 (N_13484,N_9955,N_7374);
xnor U13485 (N_13485,N_8857,N_9712);
nor U13486 (N_13486,N_7922,N_8493);
nor U13487 (N_13487,N_8077,N_7544);
and U13488 (N_13488,N_5712,N_6006);
and U13489 (N_13489,N_7168,N_7395);
and U13490 (N_13490,N_8166,N_7734);
nand U13491 (N_13491,N_6579,N_7632);
nor U13492 (N_13492,N_9871,N_9395);
xor U13493 (N_13493,N_6576,N_6707);
or U13494 (N_13494,N_8161,N_5532);
nor U13495 (N_13495,N_8670,N_8486);
and U13496 (N_13496,N_6928,N_8945);
xnor U13497 (N_13497,N_8021,N_5323);
or U13498 (N_13498,N_6628,N_6707);
nand U13499 (N_13499,N_7287,N_7968);
nand U13500 (N_13500,N_7504,N_8168);
and U13501 (N_13501,N_8482,N_6719);
nand U13502 (N_13502,N_9172,N_6953);
nand U13503 (N_13503,N_7980,N_9443);
or U13504 (N_13504,N_6214,N_5563);
or U13505 (N_13505,N_7794,N_6456);
or U13506 (N_13506,N_9541,N_8019);
nor U13507 (N_13507,N_9073,N_8589);
nand U13508 (N_13508,N_5001,N_9190);
nor U13509 (N_13509,N_7566,N_8297);
nor U13510 (N_13510,N_9446,N_5337);
and U13511 (N_13511,N_8212,N_6645);
and U13512 (N_13512,N_7375,N_9812);
nor U13513 (N_13513,N_7436,N_8659);
nand U13514 (N_13514,N_9573,N_9186);
and U13515 (N_13515,N_9807,N_8952);
or U13516 (N_13516,N_9291,N_5804);
nor U13517 (N_13517,N_5246,N_7048);
nor U13518 (N_13518,N_7412,N_9732);
and U13519 (N_13519,N_8066,N_8143);
and U13520 (N_13520,N_7606,N_9915);
and U13521 (N_13521,N_8729,N_9573);
nor U13522 (N_13522,N_6946,N_8261);
or U13523 (N_13523,N_8004,N_5319);
or U13524 (N_13524,N_6150,N_9200);
or U13525 (N_13525,N_5738,N_7046);
nor U13526 (N_13526,N_6171,N_5463);
or U13527 (N_13527,N_8893,N_6240);
and U13528 (N_13528,N_7810,N_8369);
or U13529 (N_13529,N_6827,N_7920);
or U13530 (N_13530,N_6367,N_5099);
and U13531 (N_13531,N_9592,N_7525);
nand U13532 (N_13532,N_7036,N_9260);
nor U13533 (N_13533,N_8447,N_6494);
nand U13534 (N_13534,N_6363,N_8939);
nor U13535 (N_13535,N_5014,N_6958);
nand U13536 (N_13536,N_5320,N_9034);
nor U13537 (N_13537,N_9467,N_5182);
or U13538 (N_13538,N_7021,N_9314);
or U13539 (N_13539,N_7780,N_6068);
xnor U13540 (N_13540,N_6031,N_9400);
or U13541 (N_13541,N_7876,N_7966);
nor U13542 (N_13542,N_9113,N_9177);
nor U13543 (N_13543,N_9730,N_6814);
nand U13544 (N_13544,N_9819,N_8493);
nand U13545 (N_13545,N_7393,N_9138);
and U13546 (N_13546,N_7267,N_9745);
and U13547 (N_13547,N_7889,N_7191);
xnor U13548 (N_13548,N_5106,N_9490);
nor U13549 (N_13549,N_5097,N_9695);
or U13550 (N_13550,N_7009,N_6875);
nand U13551 (N_13551,N_9757,N_5871);
nand U13552 (N_13552,N_6286,N_5895);
nor U13553 (N_13553,N_8169,N_8615);
nor U13554 (N_13554,N_9172,N_8723);
and U13555 (N_13555,N_6498,N_8434);
nand U13556 (N_13556,N_9626,N_8087);
nand U13557 (N_13557,N_9019,N_9301);
nor U13558 (N_13558,N_6745,N_5115);
nor U13559 (N_13559,N_9581,N_6556);
xor U13560 (N_13560,N_5622,N_8137);
nand U13561 (N_13561,N_8020,N_8452);
nor U13562 (N_13562,N_9919,N_6368);
nor U13563 (N_13563,N_7028,N_6085);
nor U13564 (N_13564,N_7419,N_5589);
and U13565 (N_13565,N_7164,N_7772);
or U13566 (N_13566,N_9826,N_7177);
or U13567 (N_13567,N_6965,N_8902);
xor U13568 (N_13568,N_7801,N_9245);
or U13569 (N_13569,N_6888,N_9455);
nor U13570 (N_13570,N_9613,N_9399);
nor U13571 (N_13571,N_6717,N_5343);
nand U13572 (N_13572,N_9253,N_6826);
or U13573 (N_13573,N_8446,N_6202);
nor U13574 (N_13574,N_7813,N_6915);
xor U13575 (N_13575,N_8264,N_6096);
or U13576 (N_13576,N_5917,N_9561);
nor U13577 (N_13577,N_5172,N_6279);
nand U13578 (N_13578,N_9865,N_9887);
nand U13579 (N_13579,N_7442,N_7219);
and U13580 (N_13580,N_9701,N_7019);
nor U13581 (N_13581,N_8596,N_8422);
and U13582 (N_13582,N_5625,N_6463);
nor U13583 (N_13583,N_7068,N_8911);
or U13584 (N_13584,N_7156,N_5420);
and U13585 (N_13585,N_5001,N_5877);
nand U13586 (N_13586,N_9238,N_8653);
and U13587 (N_13587,N_6593,N_6169);
nor U13588 (N_13588,N_9287,N_7868);
or U13589 (N_13589,N_6156,N_9272);
nand U13590 (N_13590,N_9116,N_5090);
and U13591 (N_13591,N_7998,N_5698);
nand U13592 (N_13592,N_8370,N_8034);
and U13593 (N_13593,N_9430,N_8342);
nor U13594 (N_13594,N_7948,N_9131);
nand U13595 (N_13595,N_9635,N_9730);
and U13596 (N_13596,N_7939,N_9562);
or U13597 (N_13597,N_6960,N_7174);
nand U13598 (N_13598,N_8364,N_5874);
or U13599 (N_13599,N_7614,N_8792);
nor U13600 (N_13600,N_7311,N_5396);
and U13601 (N_13601,N_8272,N_8221);
nor U13602 (N_13602,N_9615,N_9402);
and U13603 (N_13603,N_5789,N_8734);
and U13604 (N_13604,N_5320,N_5386);
or U13605 (N_13605,N_8388,N_7749);
or U13606 (N_13606,N_6324,N_5828);
or U13607 (N_13607,N_7949,N_5618);
nor U13608 (N_13608,N_5932,N_8677);
or U13609 (N_13609,N_8339,N_8701);
nand U13610 (N_13610,N_7678,N_6544);
nand U13611 (N_13611,N_8670,N_5792);
nor U13612 (N_13612,N_5845,N_9678);
nor U13613 (N_13613,N_7497,N_6130);
and U13614 (N_13614,N_9943,N_8677);
and U13615 (N_13615,N_6238,N_6234);
or U13616 (N_13616,N_5207,N_5254);
nand U13617 (N_13617,N_7871,N_7681);
nand U13618 (N_13618,N_7177,N_6146);
or U13619 (N_13619,N_9876,N_9801);
nand U13620 (N_13620,N_9908,N_8690);
nand U13621 (N_13621,N_6618,N_6446);
nor U13622 (N_13622,N_5816,N_7016);
nand U13623 (N_13623,N_7178,N_9231);
nand U13624 (N_13624,N_7812,N_9623);
nand U13625 (N_13625,N_8294,N_6562);
or U13626 (N_13626,N_8689,N_6374);
or U13627 (N_13627,N_9560,N_7102);
nand U13628 (N_13628,N_7648,N_5725);
and U13629 (N_13629,N_8753,N_7342);
or U13630 (N_13630,N_6403,N_8589);
nor U13631 (N_13631,N_6253,N_6442);
or U13632 (N_13632,N_8996,N_9026);
nor U13633 (N_13633,N_5339,N_5962);
nor U13634 (N_13634,N_9592,N_5614);
nor U13635 (N_13635,N_8772,N_9097);
and U13636 (N_13636,N_7533,N_6446);
and U13637 (N_13637,N_8046,N_5725);
nand U13638 (N_13638,N_6264,N_9236);
or U13639 (N_13639,N_7502,N_6668);
nor U13640 (N_13640,N_6805,N_5971);
or U13641 (N_13641,N_6180,N_5884);
or U13642 (N_13642,N_9756,N_7853);
and U13643 (N_13643,N_8493,N_8084);
nor U13644 (N_13644,N_6035,N_8144);
nand U13645 (N_13645,N_5548,N_9660);
and U13646 (N_13646,N_8957,N_9015);
and U13647 (N_13647,N_5129,N_6120);
and U13648 (N_13648,N_6607,N_7833);
nor U13649 (N_13649,N_7624,N_8578);
nand U13650 (N_13650,N_5680,N_8365);
nand U13651 (N_13651,N_8562,N_7550);
or U13652 (N_13652,N_9348,N_7554);
or U13653 (N_13653,N_6301,N_9270);
and U13654 (N_13654,N_7233,N_7972);
nor U13655 (N_13655,N_7571,N_9440);
nor U13656 (N_13656,N_9391,N_8013);
or U13657 (N_13657,N_5098,N_6324);
nor U13658 (N_13658,N_5048,N_7418);
or U13659 (N_13659,N_8827,N_9739);
nor U13660 (N_13660,N_8627,N_9988);
or U13661 (N_13661,N_8638,N_6955);
or U13662 (N_13662,N_5685,N_9063);
xnor U13663 (N_13663,N_7508,N_8480);
nand U13664 (N_13664,N_6741,N_6743);
and U13665 (N_13665,N_5486,N_6616);
nor U13666 (N_13666,N_5294,N_5176);
or U13667 (N_13667,N_8201,N_6992);
and U13668 (N_13668,N_5177,N_5109);
xor U13669 (N_13669,N_7900,N_9022);
nand U13670 (N_13670,N_7305,N_5634);
xor U13671 (N_13671,N_7921,N_8926);
or U13672 (N_13672,N_5741,N_8301);
or U13673 (N_13673,N_9514,N_6249);
nor U13674 (N_13674,N_8020,N_9920);
or U13675 (N_13675,N_6836,N_5355);
or U13676 (N_13676,N_5993,N_8202);
nand U13677 (N_13677,N_8231,N_6496);
nor U13678 (N_13678,N_8580,N_6812);
and U13679 (N_13679,N_6320,N_7774);
nor U13680 (N_13680,N_5115,N_7700);
and U13681 (N_13681,N_8203,N_7316);
nor U13682 (N_13682,N_9767,N_9536);
nor U13683 (N_13683,N_7331,N_9914);
nand U13684 (N_13684,N_8978,N_9421);
nand U13685 (N_13685,N_5236,N_9235);
or U13686 (N_13686,N_6260,N_7931);
or U13687 (N_13687,N_5765,N_9847);
nand U13688 (N_13688,N_5297,N_6977);
and U13689 (N_13689,N_8669,N_8909);
nand U13690 (N_13690,N_9763,N_8708);
nand U13691 (N_13691,N_6922,N_7185);
or U13692 (N_13692,N_6516,N_7955);
nor U13693 (N_13693,N_7445,N_8928);
and U13694 (N_13694,N_9459,N_8632);
nand U13695 (N_13695,N_5136,N_5388);
nand U13696 (N_13696,N_6366,N_6764);
or U13697 (N_13697,N_9023,N_7190);
nor U13698 (N_13698,N_8760,N_9199);
or U13699 (N_13699,N_7961,N_9889);
or U13700 (N_13700,N_6544,N_5421);
nand U13701 (N_13701,N_7106,N_9071);
nand U13702 (N_13702,N_8412,N_8425);
and U13703 (N_13703,N_7624,N_7023);
or U13704 (N_13704,N_8215,N_5062);
and U13705 (N_13705,N_5976,N_9829);
or U13706 (N_13706,N_8083,N_7290);
and U13707 (N_13707,N_6450,N_7681);
nand U13708 (N_13708,N_8205,N_7999);
nor U13709 (N_13709,N_7703,N_5983);
or U13710 (N_13710,N_8046,N_8125);
nand U13711 (N_13711,N_7159,N_6310);
nor U13712 (N_13712,N_5571,N_5278);
nor U13713 (N_13713,N_5128,N_7108);
nand U13714 (N_13714,N_7570,N_9078);
or U13715 (N_13715,N_8814,N_5139);
and U13716 (N_13716,N_9217,N_7948);
or U13717 (N_13717,N_8130,N_8605);
and U13718 (N_13718,N_7412,N_9181);
nor U13719 (N_13719,N_9298,N_8572);
nand U13720 (N_13720,N_7785,N_9318);
and U13721 (N_13721,N_9316,N_8055);
nand U13722 (N_13722,N_5972,N_5665);
nand U13723 (N_13723,N_8183,N_6239);
nand U13724 (N_13724,N_6643,N_5714);
nor U13725 (N_13725,N_5126,N_6402);
nand U13726 (N_13726,N_9148,N_6323);
nor U13727 (N_13727,N_6140,N_6800);
and U13728 (N_13728,N_7212,N_7679);
xnor U13729 (N_13729,N_8928,N_8240);
or U13730 (N_13730,N_8611,N_7769);
nand U13731 (N_13731,N_7019,N_9183);
or U13732 (N_13732,N_7549,N_8982);
nor U13733 (N_13733,N_9514,N_8850);
nand U13734 (N_13734,N_5633,N_5135);
and U13735 (N_13735,N_7193,N_6874);
or U13736 (N_13736,N_5791,N_7170);
or U13737 (N_13737,N_7984,N_7029);
nand U13738 (N_13738,N_7811,N_9847);
or U13739 (N_13739,N_7932,N_7282);
or U13740 (N_13740,N_5170,N_9222);
nand U13741 (N_13741,N_9540,N_7011);
or U13742 (N_13742,N_7577,N_7102);
and U13743 (N_13743,N_5509,N_8379);
and U13744 (N_13744,N_5664,N_7880);
nand U13745 (N_13745,N_7891,N_6705);
xor U13746 (N_13746,N_7785,N_5313);
or U13747 (N_13747,N_8657,N_8586);
nor U13748 (N_13748,N_7446,N_6879);
nand U13749 (N_13749,N_6051,N_7210);
or U13750 (N_13750,N_9159,N_9481);
or U13751 (N_13751,N_8169,N_9288);
nand U13752 (N_13752,N_8842,N_6310);
and U13753 (N_13753,N_5560,N_5924);
nor U13754 (N_13754,N_9083,N_6238);
or U13755 (N_13755,N_9013,N_9016);
and U13756 (N_13756,N_7034,N_7968);
nor U13757 (N_13757,N_6748,N_8627);
or U13758 (N_13758,N_8631,N_9957);
or U13759 (N_13759,N_8764,N_6049);
and U13760 (N_13760,N_6870,N_9618);
and U13761 (N_13761,N_5812,N_7669);
nor U13762 (N_13762,N_6533,N_7850);
nor U13763 (N_13763,N_7091,N_9317);
or U13764 (N_13764,N_6084,N_5127);
and U13765 (N_13765,N_9464,N_6762);
and U13766 (N_13766,N_9112,N_6600);
nand U13767 (N_13767,N_5897,N_5823);
or U13768 (N_13768,N_8212,N_8832);
nor U13769 (N_13769,N_7138,N_9448);
or U13770 (N_13770,N_7234,N_7104);
or U13771 (N_13771,N_6550,N_7161);
or U13772 (N_13772,N_9203,N_7486);
xnor U13773 (N_13773,N_7122,N_9601);
nand U13774 (N_13774,N_6349,N_9173);
or U13775 (N_13775,N_7619,N_6564);
nor U13776 (N_13776,N_8454,N_6181);
nand U13777 (N_13777,N_7092,N_8364);
or U13778 (N_13778,N_8671,N_5220);
and U13779 (N_13779,N_5538,N_5488);
and U13780 (N_13780,N_9748,N_7794);
nand U13781 (N_13781,N_5587,N_7976);
or U13782 (N_13782,N_9213,N_6019);
nand U13783 (N_13783,N_9723,N_8954);
nand U13784 (N_13784,N_8536,N_8541);
and U13785 (N_13785,N_9975,N_9557);
or U13786 (N_13786,N_8850,N_6429);
nor U13787 (N_13787,N_6701,N_8138);
nand U13788 (N_13788,N_7533,N_5537);
nor U13789 (N_13789,N_7970,N_7921);
nand U13790 (N_13790,N_5747,N_6196);
nand U13791 (N_13791,N_6224,N_5886);
nor U13792 (N_13792,N_7446,N_6490);
nand U13793 (N_13793,N_8310,N_5192);
nand U13794 (N_13794,N_8168,N_8064);
and U13795 (N_13795,N_6863,N_7037);
or U13796 (N_13796,N_8981,N_7122);
and U13797 (N_13797,N_6046,N_8540);
nand U13798 (N_13798,N_6449,N_6954);
and U13799 (N_13799,N_5145,N_7783);
nor U13800 (N_13800,N_5047,N_6260);
and U13801 (N_13801,N_8969,N_6149);
and U13802 (N_13802,N_9824,N_9063);
nand U13803 (N_13803,N_8156,N_5173);
or U13804 (N_13804,N_8094,N_5523);
or U13805 (N_13805,N_8148,N_6520);
nand U13806 (N_13806,N_8011,N_9607);
and U13807 (N_13807,N_9497,N_6744);
nor U13808 (N_13808,N_8488,N_6431);
and U13809 (N_13809,N_6847,N_7435);
nor U13810 (N_13810,N_6704,N_5185);
or U13811 (N_13811,N_7524,N_9672);
nor U13812 (N_13812,N_8282,N_6270);
nand U13813 (N_13813,N_8033,N_7811);
nand U13814 (N_13814,N_6039,N_6283);
nand U13815 (N_13815,N_6559,N_9738);
and U13816 (N_13816,N_7678,N_8837);
and U13817 (N_13817,N_6556,N_9373);
xor U13818 (N_13818,N_7194,N_9225);
or U13819 (N_13819,N_5916,N_8577);
or U13820 (N_13820,N_7217,N_5550);
or U13821 (N_13821,N_8535,N_7222);
nand U13822 (N_13822,N_5415,N_6069);
nand U13823 (N_13823,N_5976,N_8769);
or U13824 (N_13824,N_5369,N_7795);
nand U13825 (N_13825,N_8567,N_7377);
or U13826 (N_13826,N_7737,N_5340);
and U13827 (N_13827,N_6609,N_6111);
and U13828 (N_13828,N_6359,N_6606);
nand U13829 (N_13829,N_9600,N_8511);
nor U13830 (N_13830,N_7366,N_9640);
nor U13831 (N_13831,N_9498,N_6268);
nand U13832 (N_13832,N_9013,N_9105);
or U13833 (N_13833,N_7153,N_9920);
nor U13834 (N_13834,N_6383,N_7733);
nor U13835 (N_13835,N_5089,N_7180);
nor U13836 (N_13836,N_8075,N_7868);
or U13837 (N_13837,N_8294,N_8298);
nor U13838 (N_13838,N_6576,N_6552);
nor U13839 (N_13839,N_8720,N_6255);
nor U13840 (N_13840,N_9919,N_7013);
nor U13841 (N_13841,N_6641,N_6929);
nand U13842 (N_13842,N_8357,N_7596);
or U13843 (N_13843,N_5129,N_6764);
nor U13844 (N_13844,N_9495,N_8091);
nand U13845 (N_13845,N_5798,N_8036);
or U13846 (N_13846,N_5540,N_6653);
or U13847 (N_13847,N_7075,N_7611);
nand U13848 (N_13848,N_9711,N_5446);
or U13849 (N_13849,N_5118,N_5022);
nor U13850 (N_13850,N_7215,N_6203);
or U13851 (N_13851,N_6876,N_8597);
and U13852 (N_13852,N_7609,N_8826);
nor U13853 (N_13853,N_6051,N_8678);
nand U13854 (N_13854,N_5449,N_9701);
or U13855 (N_13855,N_9406,N_8990);
nand U13856 (N_13856,N_9849,N_8362);
nor U13857 (N_13857,N_8394,N_6014);
nor U13858 (N_13858,N_9517,N_9962);
and U13859 (N_13859,N_8128,N_6270);
nand U13860 (N_13860,N_7054,N_9074);
and U13861 (N_13861,N_5878,N_5457);
or U13862 (N_13862,N_7284,N_7229);
nand U13863 (N_13863,N_9295,N_9871);
nand U13864 (N_13864,N_7753,N_5946);
nor U13865 (N_13865,N_8035,N_5734);
or U13866 (N_13866,N_6486,N_9610);
or U13867 (N_13867,N_5562,N_6582);
nand U13868 (N_13868,N_9843,N_6501);
and U13869 (N_13869,N_5623,N_5876);
or U13870 (N_13870,N_9272,N_6739);
xor U13871 (N_13871,N_9160,N_8164);
or U13872 (N_13872,N_8224,N_8687);
and U13873 (N_13873,N_6077,N_6549);
or U13874 (N_13874,N_6248,N_6446);
nand U13875 (N_13875,N_7048,N_9945);
nand U13876 (N_13876,N_6253,N_8321);
or U13877 (N_13877,N_8611,N_9103);
nand U13878 (N_13878,N_7059,N_7568);
and U13879 (N_13879,N_8651,N_8760);
or U13880 (N_13880,N_8207,N_9265);
or U13881 (N_13881,N_8892,N_6601);
nand U13882 (N_13882,N_7017,N_8453);
or U13883 (N_13883,N_6776,N_5943);
or U13884 (N_13884,N_5733,N_5686);
nor U13885 (N_13885,N_7952,N_5183);
nand U13886 (N_13886,N_8585,N_7017);
nor U13887 (N_13887,N_5195,N_7997);
and U13888 (N_13888,N_8093,N_8564);
and U13889 (N_13889,N_5918,N_5615);
or U13890 (N_13890,N_5924,N_5007);
or U13891 (N_13891,N_8720,N_7190);
xor U13892 (N_13892,N_5976,N_7137);
nand U13893 (N_13893,N_5376,N_6587);
nor U13894 (N_13894,N_8102,N_7218);
nand U13895 (N_13895,N_5361,N_8720);
nor U13896 (N_13896,N_8641,N_6179);
xor U13897 (N_13897,N_5390,N_6224);
nor U13898 (N_13898,N_6586,N_7333);
nor U13899 (N_13899,N_8674,N_7795);
and U13900 (N_13900,N_6420,N_5135);
nand U13901 (N_13901,N_8765,N_9236);
and U13902 (N_13902,N_5881,N_9333);
nand U13903 (N_13903,N_6043,N_7772);
and U13904 (N_13904,N_8222,N_9212);
or U13905 (N_13905,N_6747,N_5462);
xor U13906 (N_13906,N_7408,N_8706);
nor U13907 (N_13907,N_9966,N_6209);
or U13908 (N_13908,N_7315,N_8499);
and U13909 (N_13909,N_5709,N_9581);
nor U13910 (N_13910,N_8238,N_8384);
or U13911 (N_13911,N_7845,N_8411);
or U13912 (N_13912,N_8673,N_5682);
or U13913 (N_13913,N_6432,N_7530);
or U13914 (N_13914,N_8979,N_8994);
nor U13915 (N_13915,N_8764,N_7959);
or U13916 (N_13916,N_6004,N_9754);
nand U13917 (N_13917,N_8173,N_9860);
or U13918 (N_13918,N_7706,N_9243);
nand U13919 (N_13919,N_8617,N_8209);
and U13920 (N_13920,N_6699,N_8745);
and U13921 (N_13921,N_5835,N_7235);
or U13922 (N_13922,N_8677,N_6020);
nor U13923 (N_13923,N_7024,N_7643);
nor U13924 (N_13924,N_7734,N_6048);
nand U13925 (N_13925,N_9580,N_6771);
nand U13926 (N_13926,N_8798,N_5099);
or U13927 (N_13927,N_9914,N_5089);
xnor U13928 (N_13928,N_8408,N_9652);
or U13929 (N_13929,N_5837,N_9869);
and U13930 (N_13930,N_8749,N_5824);
or U13931 (N_13931,N_7503,N_7765);
and U13932 (N_13932,N_6133,N_7283);
nor U13933 (N_13933,N_9994,N_8028);
nand U13934 (N_13934,N_5207,N_9753);
or U13935 (N_13935,N_5411,N_6112);
nand U13936 (N_13936,N_7161,N_7049);
and U13937 (N_13937,N_9474,N_6343);
or U13938 (N_13938,N_6196,N_8165);
nand U13939 (N_13939,N_8601,N_9004);
and U13940 (N_13940,N_9660,N_8959);
nand U13941 (N_13941,N_8765,N_9531);
and U13942 (N_13942,N_9345,N_8394);
xor U13943 (N_13943,N_5357,N_9463);
and U13944 (N_13944,N_7391,N_7320);
and U13945 (N_13945,N_5925,N_7213);
or U13946 (N_13946,N_9437,N_6701);
nand U13947 (N_13947,N_8524,N_5966);
nand U13948 (N_13948,N_6597,N_9113);
or U13949 (N_13949,N_8128,N_9008);
nand U13950 (N_13950,N_9500,N_5426);
nand U13951 (N_13951,N_9625,N_8635);
nand U13952 (N_13952,N_6429,N_8199);
or U13953 (N_13953,N_7053,N_7061);
and U13954 (N_13954,N_9560,N_8475);
nor U13955 (N_13955,N_5595,N_7210);
or U13956 (N_13956,N_5755,N_5792);
nand U13957 (N_13957,N_9683,N_8705);
and U13958 (N_13958,N_5695,N_7894);
and U13959 (N_13959,N_6116,N_8741);
nor U13960 (N_13960,N_6946,N_6751);
nand U13961 (N_13961,N_7629,N_6395);
or U13962 (N_13962,N_9557,N_5392);
or U13963 (N_13963,N_8354,N_8559);
and U13964 (N_13964,N_9746,N_6066);
nor U13965 (N_13965,N_7640,N_8159);
or U13966 (N_13966,N_8545,N_6610);
nor U13967 (N_13967,N_6819,N_5535);
xor U13968 (N_13968,N_5540,N_9508);
nand U13969 (N_13969,N_5219,N_8395);
and U13970 (N_13970,N_6857,N_8320);
and U13971 (N_13971,N_5405,N_7793);
or U13972 (N_13972,N_7393,N_8280);
or U13973 (N_13973,N_6311,N_9780);
and U13974 (N_13974,N_6056,N_6212);
nor U13975 (N_13975,N_8616,N_8442);
nand U13976 (N_13976,N_6398,N_5420);
and U13977 (N_13977,N_6056,N_5330);
nand U13978 (N_13978,N_5443,N_7927);
and U13979 (N_13979,N_5042,N_6990);
nand U13980 (N_13980,N_7353,N_6112);
or U13981 (N_13981,N_9550,N_8472);
or U13982 (N_13982,N_5753,N_5626);
nor U13983 (N_13983,N_5916,N_9577);
and U13984 (N_13984,N_8025,N_7518);
or U13985 (N_13985,N_6155,N_9095);
and U13986 (N_13986,N_6781,N_9405);
or U13987 (N_13987,N_9223,N_8175);
nor U13988 (N_13988,N_9129,N_9038);
nor U13989 (N_13989,N_8155,N_8174);
nor U13990 (N_13990,N_6332,N_6833);
nand U13991 (N_13991,N_5893,N_6490);
nand U13992 (N_13992,N_6699,N_7885);
or U13993 (N_13993,N_6861,N_9378);
nor U13994 (N_13994,N_5774,N_7648);
nand U13995 (N_13995,N_9674,N_8719);
and U13996 (N_13996,N_6366,N_9463);
or U13997 (N_13997,N_8012,N_9567);
nand U13998 (N_13998,N_7718,N_9349);
nand U13999 (N_13999,N_8831,N_7742);
and U14000 (N_14000,N_6303,N_6377);
or U14001 (N_14001,N_9994,N_7667);
nor U14002 (N_14002,N_9605,N_9039);
nor U14003 (N_14003,N_8406,N_9437);
nand U14004 (N_14004,N_7244,N_7419);
or U14005 (N_14005,N_7935,N_7963);
or U14006 (N_14006,N_7899,N_9855);
and U14007 (N_14007,N_6380,N_5774);
nand U14008 (N_14008,N_5537,N_9987);
nand U14009 (N_14009,N_8945,N_9896);
and U14010 (N_14010,N_6777,N_5215);
nor U14011 (N_14011,N_8518,N_5457);
or U14012 (N_14012,N_5844,N_5226);
nor U14013 (N_14013,N_9242,N_6788);
nand U14014 (N_14014,N_5421,N_5401);
and U14015 (N_14015,N_5240,N_6178);
and U14016 (N_14016,N_5255,N_7132);
nor U14017 (N_14017,N_6186,N_7371);
and U14018 (N_14018,N_9334,N_5842);
nand U14019 (N_14019,N_7818,N_8409);
nor U14020 (N_14020,N_9083,N_6383);
or U14021 (N_14021,N_6505,N_9227);
nor U14022 (N_14022,N_7927,N_6294);
nand U14023 (N_14023,N_5205,N_9293);
nor U14024 (N_14024,N_7888,N_8358);
or U14025 (N_14025,N_8956,N_9063);
nor U14026 (N_14026,N_9548,N_7171);
nor U14027 (N_14027,N_8362,N_6630);
nand U14028 (N_14028,N_8580,N_6641);
or U14029 (N_14029,N_7741,N_7147);
and U14030 (N_14030,N_6267,N_8745);
and U14031 (N_14031,N_9730,N_8584);
or U14032 (N_14032,N_5493,N_5859);
and U14033 (N_14033,N_7548,N_5544);
nor U14034 (N_14034,N_7317,N_8110);
nand U14035 (N_14035,N_9027,N_6258);
nor U14036 (N_14036,N_6385,N_8804);
or U14037 (N_14037,N_7671,N_7953);
and U14038 (N_14038,N_9603,N_6432);
nor U14039 (N_14039,N_7811,N_5381);
nand U14040 (N_14040,N_8774,N_9193);
or U14041 (N_14041,N_8823,N_8629);
nor U14042 (N_14042,N_9235,N_9690);
nor U14043 (N_14043,N_5902,N_6849);
nand U14044 (N_14044,N_6830,N_9511);
nand U14045 (N_14045,N_5945,N_8031);
nand U14046 (N_14046,N_8542,N_8150);
nand U14047 (N_14047,N_7763,N_9663);
nor U14048 (N_14048,N_6285,N_8343);
nor U14049 (N_14049,N_7983,N_6273);
nor U14050 (N_14050,N_6448,N_9861);
and U14051 (N_14051,N_7474,N_7862);
nor U14052 (N_14052,N_5816,N_6860);
or U14053 (N_14053,N_7782,N_5021);
or U14054 (N_14054,N_6238,N_8394);
or U14055 (N_14055,N_9155,N_9801);
and U14056 (N_14056,N_6647,N_5930);
or U14057 (N_14057,N_6564,N_8479);
nor U14058 (N_14058,N_9653,N_9789);
nor U14059 (N_14059,N_6379,N_7876);
nor U14060 (N_14060,N_7054,N_7513);
nand U14061 (N_14061,N_6183,N_6757);
or U14062 (N_14062,N_6277,N_8286);
or U14063 (N_14063,N_9410,N_7640);
or U14064 (N_14064,N_9017,N_7191);
nand U14065 (N_14065,N_7300,N_5529);
nor U14066 (N_14066,N_9400,N_6344);
or U14067 (N_14067,N_6797,N_5012);
nor U14068 (N_14068,N_5155,N_6048);
nand U14069 (N_14069,N_7543,N_9310);
and U14070 (N_14070,N_8524,N_8513);
nor U14071 (N_14071,N_9348,N_6535);
nor U14072 (N_14072,N_7601,N_7025);
nand U14073 (N_14073,N_6558,N_8595);
nor U14074 (N_14074,N_8461,N_8158);
and U14075 (N_14075,N_7059,N_7948);
nor U14076 (N_14076,N_9983,N_9002);
and U14077 (N_14077,N_5927,N_7022);
nand U14078 (N_14078,N_8183,N_6035);
or U14079 (N_14079,N_9255,N_8234);
and U14080 (N_14080,N_7537,N_7575);
and U14081 (N_14081,N_8373,N_6968);
or U14082 (N_14082,N_8377,N_5146);
or U14083 (N_14083,N_5991,N_5947);
nor U14084 (N_14084,N_6330,N_6003);
nor U14085 (N_14085,N_9969,N_8672);
nand U14086 (N_14086,N_7560,N_7259);
and U14087 (N_14087,N_6439,N_8530);
nand U14088 (N_14088,N_9386,N_7200);
nor U14089 (N_14089,N_5932,N_8401);
or U14090 (N_14090,N_9262,N_9847);
or U14091 (N_14091,N_8676,N_5817);
or U14092 (N_14092,N_6331,N_8501);
or U14093 (N_14093,N_8598,N_7563);
nor U14094 (N_14094,N_9670,N_8956);
nor U14095 (N_14095,N_5354,N_7949);
nand U14096 (N_14096,N_6523,N_8403);
and U14097 (N_14097,N_7543,N_8047);
or U14098 (N_14098,N_9523,N_8421);
nand U14099 (N_14099,N_8157,N_7994);
and U14100 (N_14100,N_5512,N_7864);
or U14101 (N_14101,N_6341,N_6388);
or U14102 (N_14102,N_6878,N_8800);
nand U14103 (N_14103,N_7684,N_8860);
and U14104 (N_14104,N_6462,N_7815);
nand U14105 (N_14105,N_9011,N_6861);
and U14106 (N_14106,N_5894,N_7640);
nor U14107 (N_14107,N_9461,N_9522);
and U14108 (N_14108,N_5127,N_5555);
nand U14109 (N_14109,N_7400,N_8868);
nand U14110 (N_14110,N_5186,N_6515);
xnor U14111 (N_14111,N_5151,N_9637);
and U14112 (N_14112,N_5930,N_7313);
or U14113 (N_14113,N_7372,N_6567);
or U14114 (N_14114,N_9881,N_5025);
or U14115 (N_14115,N_6183,N_7049);
nor U14116 (N_14116,N_7175,N_7016);
nand U14117 (N_14117,N_5811,N_6117);
nor U14118 (N_14118,N_5285,N_7349);
or U14119 (N_14119,N_9619,N_9724);
or U14120 (N_14120,N_5025,N_8183);
and U14121 (N_14121,N_5047,N_6305);
nand U14122 (N_14122,N_8732,N_7103);
nand U14123 (N_14123,N_7429,N_9187);
and U14124 (N_14124,N_5751,N_6587);
or U14125 (N_14125,N_9347,N_7716);
or U14126 (N_14126,N_6466,N_8742);
and U14127 (N_14127,N_8041,N_7300);
nor U14128 (N_14128,N_5761,N_6392);
and U14129 (N_14129,N_8422,N_8158);
nand U14130 (N_14130,N_8122,N_5256);
and U14131 (N_14131,N_7482,N_9003);
and U14132 (N_14132,N_9557,N_8766);
nor U14133 (N_14133,N_7301,N_7631);
nor U14134 (N_14134,N_5044,N_9534);
and U14135 (N_14135,N_6618,N_5695);
nor U14136 (N_14136,N_9193,N_6842);
nand U14137 (N_14137,N_7513,N_6372);
nor U14138 (N_14138,N_9987,N_7699);
and U14139 (N_14139,N_6917,N_6285);
nand U14140 (N_14140,N_5853,N_8584);
nor U14141 (N_14141,N_6791,N_9896);
nor U14142 (N_14142,N_8318,N_9640);
nand U14143 (N_14143,N_6068,N_9855);
and U14144 (N_14144,N_7984,N_5664);
or U14145 (N_14145,N_6751,N_8330);
and U14146 (N_14146,N_9722,N_9513);
nand U14147 (N_14147,N_9552,N_9160);
nand U14148 (N_14148,N_6011,N_6669);
nand U14149 (N_14149,N_5447,N_6358);
or U14150 (N_14150,N_7925,N_5809);
nor U14151 (N_14151,N_9750,N_6137);
nand U14152 (N_14152,N_8170,N_5036);
nand U14153 (N_14153,N_6906,N_5546);
xnor U14154 (N_14154,N_8470,N_7647);
and U14155 (N_14155,N_8356,N_7453);
nand U14156 (N_14156,N_5129,N_8662);
or U14157 (N_14157,N_7055,N_5548);
or U14158 (N_14158,N_5787,N_9413);
and U14159 (N_14159,N_5069,N_8261);
and U14160 (N_14160,N_6545,N_6538);
and U14161 (N_14161,N_9120,N_8287);
and U14162 (N_14162,N_6932,N_7701);
nand U14163 (N_14163,N_6459,N_7778);
and U14164 (N_14164,N_9097,N_7172);
nor U14165 (N_14165,N_5902,N_5458);
nand U14166 (N_14166,N_8845,N_5884);
or U14167 (N_14167,N_6037,N_6877);
nand U14168 (N_14168,N_6150,N_5887);
and U14169 (N_14169,N_7937,N_9655);
or U14170 (N_14170,N_7178,N_9283);
and U14171 (N_14171,N_9753,N_9912);
and U14172 (N_14172,N_8599,N_7128);
nand U14173 (N_14173,N_5934,N_9060);
or U14174 (N_14174,N_8074,N_5625);
or U14175 (N_14175,N_8277,N_7164);
or U14176 (N_14176,N_5584,N_6549);
nand U14177 (N_14177,N_5047,N_8126);
or U14178 (N_14178,N_7317,N_9308);
or U14179 (N_14179,N_6776,N_8488);
nand U14180 (N_14180,N_8856,N_7338);
or U14181 (N_14181,N_6143,N_9280);
nor U14182 (N_14182,N_8191,N_9893);
nand U14183 (N_14183,N_9832,N_9013);
or U14184 (N_14184,N_9953,N_6486);
nor U14185 (N_14185,N_9449,N_6091);
nand U14186 (N_14186,N_9271,N_6486);
nand U14187 (N_14187,N_8463,N_6443);
nor U14188 (N_14188,N_9596,N_9363);
or U14189 (N_14189,N_7887,N_7494);
and U14190 (N_14190,N_5946,N_7261);
or U14191 (N_14191,N_5689,N_5615);
or U14192 (N_14192,N_7799,N_5889);
nand U14193 (N_14193,N_9765,N_7111);
nand U14194 (N_14194,N_8561,N_9810);
nand U14195 (N_14195,N_8108,N_6689);
and U14196 (N_14196,N_6194,N_8254);
and U14197 (N_14197,N_7057,N_6868);
nand U14198 (N_14198,N_9766,N_7864);
and U14199 (N_14199,N_8660,N_5680);
nor U14200 (N_14200,N_7185,N_6601);
nor U14201 (N_14201,N_8169,N_6707);
nor U14202 (N_14202,N_6049,N_5965);
nor U14203 (N_14203,N_6364,N_8120);
and U14204 (N_14204,N_7106,N_7210);
or U14205 (N_14205,N_7069,N_7586);
or U14206 (N_14206,N_5411,N_9753);
or U14207 (N_14207,N_7149,N_5710);
nand U14208 (N_14208,N_6650,N_6249);
or U14209 (N_14209,N_8648,N_8489);
nand U14210 (N_14210,N_8736,N_5767);
xor U14211 (N_14211,N_5620,N_6662);
and U14212 (N_14212,N_8933,N_5810);
nand U14213 (N_14213,N_8349,N_8091);
nand U14214 (N_14214,N_5612,N_6628);
or U14215 (N_14215,N_7926,N_9784);
nand U14216 (N_14216,N_5338,N_7469);
nor U14217 (N_14217,N_5800,N_9357);
nand U14218 (N_14218,N_6073,N_5883);
and U14219 (N_14219,N_7389,N_8595);
or U14220 (N_14220,N_5619,N_8109);
or U14221 (N_14221,N_7998,N_9317);
nand U14222 (N_14222,N_7157,N_8117);
nor U14223 (N_14223,N_6139,N_8993);
nor U14224 (N_14224,N_5634,N_7728);
nand U14225 (N_14225,N_6556,N_9420);
and U14226 (N_14226,N_9380,N_7735);
and U14227 (N_14227,N_8319,N_5095);
and U14228 (N_14228,N_6606,N_5414);
nor U14229 (N_14229,N_5698,N_5437);
nor U14230 (N_14230,N_5415,N_8260);
nor U14231 (N_14231,N_9213,N_9480);
xor U14232 (N_14232,N_6951,N_7529);
nor U14233 (N_14233,N_5692,N_8398);
and U14234 (N_14234,N_9479,N_9141);
and U14235 (N_14235,N_8743,N_7463);
nand U14236 (N_14236,N_5984,N_6798);
and U14237 (N_14237,N_7089,N_6344);
and U14238 (N_14238,N_5425,N_6066);
nand U14239 (N_14239,N_5177,N_7872);
or U14240 (N_14240,N_7392,N_6436);
or U14241 (N_14241,N_9040,N_5804);
nand U14242 (N_14242,N_7023,N_5492);
nor U14243 (N_14243,N_6841,N_7167);
nor U14244 (N_14244,N_5054,N_6414);
xnor U14245 (N_14245,N_8062,N_5509);
and U14246 (N_14246,N_7016,N_8083);
and U14247 (N_14247,N_8671,N_9995);
nand U14248 (N_14248,N_9156,N_6145);
nand U14249 (N_14249,N_5101,N_7653);
and U14250 (N_14250,N_9556,N_5189);
and U14251 (N_14251,N_7252,N_7133);
and U14252 (N_14252,N_6771,N_9980);
nor U14253 (N_14253,N_5858,N_9989);
and U14254 (N_14254,N_6010,N_6437);
nand U14255 (N_14255,N_6696,N_6301);
nor U14256 (N_14256,N_9915,N_6195);
nand U14257 (N_14257,N_9587,N_9992);
nor U14258 (N_14258,N_7619,N_6168);
nor U14259 (N_14259,N_7665,N_5347);
and U14260 (N_14260,N_7943,N_8812);
nand U14261 (N_14261,N_9399,N_6873);
nor U14262 (N_14262,N_9169,N_9474);
nand U14263 (N_14263,N_7126,N_5494);
nand U14264 (N_14264,N_8616,N_5294);
nor U14265 (N_14265,N_5840,N_8311);
or U14266 (N_14266,N_7435,N_9755);
nand U14267 (N_14267,N_6351,N_5696);
and U14268 (N_14268,N_9457,N_5581);
and U14269 (N_14269,N_6222,N_9823);
and U14270 (N_14270,N_6261,N_7749);
and U14271 (N_14271,N_8299,N_7607);
nor U14272 (N_14272,N_9661,N_7832);
or U14273 (N_14273,N_6010,N_7492);
nand U14274 (N_14274,N_7599,N_7980);
nor U14275 (N_14275,N_7000,N_6927);
nor U14276 (N_14276,N_9234,N_7509);
nand U14277 (N_14277,N_6717,N_7052);
or U14278 (N_14278,N_8007,N_7821);
or U14279 (N_14279,N_6179,N_7608);
or U14280 (N_14280,N_5449,N_7155);
nand U14281 (N_14281,N_9355,N_7819);
nand U14282 (N_14282,N_5597,N_8322);
or U14283 (N_14283,N_7064,N_5849);
nor U14284 (N_14284,N_7486,N_9377);
nor U14285 (N_14285,N_5995,N_9320);
or U14286 (N_14286,N_8880,N_9990);
and U14287 (N_14287,N_8213,N_9521);
or U14288 (N_14288,N_6427,N_9114);
or U14289 (N_14289,N_6830,N_8567);
nor U14290 (N_14290,N_5366,N_7648);
or U14291 (N_14291,N_8184,N_5146);
or U14292 (N_14292,N_6464,N_7493);
xnor U14293 (N_14293,N_5609,N_7539);
or U14294 (N_14294,N_9424,N_9783);
nor U14295 (N_14295,N_6520,N_9197);
and U14296 (N_14296,N_7165,N_9594);
or U14297 (N_14297,N_7074,N_8240);
nor U14298 (N_14298,N_8677,N_5155);
nand U14299 (N_14299,N_7951,N_8710);
or U14300 (N_14300,N_6055,N_5299);
nor U14301 (N_14301,N_6687,N_8170);
nand U14302 (N_14302,N_5134,N_8324);
nand U14303 (N_14303,N_5664,N_8473);
or U14304 (N_14304,N_9320,N_5022);
or U14305 (N_14305,N_7996,N_7196);
and U14306 (N_14306,N_9836,N_6454);
nor U14307 (N_14307,N_7831,N_5933);
or U14308 (N_14308,N_7480,N_6514);
nor U14309 (N_14309,N_5954,N_8077);
nor U14310 (N_14310,N_8808,N_9537);
nor U14311 (N_14311,N_6666,N_5556);
nand U14312 (N_14312,N_9433,N_7782);
and U14313 (N_14313,N_7848,N_8319);
nor U14314 (N_14314,N_7191,N_5126);
and U14315 (N_14315,N_8754,N_6739);
and U14316 (N_14316,N_9579,N_6130);
or U14317 (N_14317,N_5478,N_6875);
nand U14318 (N_14318,N_9939,N_5137);
nand U14319 (N_14319,N_7538,N_6927);
and U14320 (N_14320,N_8599,N_7371);
and U14321 (N_14321,N_9162,N_9857);
nor U14322 (N_14322,N_5698,N_8196);
and U14323 (N_14323,N_6044,N_7341);
or U14324 (N_14324,N_8269,N_7183);
and U14325 (N_14325,N_9902,N_9304);
nor U14326 (N_14326,N_6778,N_8944);
nor U14327 (N_14327,N_8167,N_7326);
or U14328 (N_14328,N_8731,N_6510);
and U14329 (N_14329,N_6269,N_6669);
nand U14330 (N_14330,N_8567,N_5334);
and U14331 (N_14331,N_8641,N_6118);
or U14332 (N_14332,N_5982,N_7159);
nand U14333 (N_14333,N_9992,N_9525);
and U14334 (N_14334,N_6570,N_6761);
and U14335 (N_14335,N_5791,N_8150);
or U14336 (N_14336,N_5996,N_6682);
and U14337 (N_14337,N_6827,N_6518);
nor U14338 (N_14338,N_8601,N_6489);
nor U14339 (N_14339,N_9292,N_9391);
nor U14340 (N_14340,N_6805,N_6139);
or U14341 (N_14341,N_8894,N_5291);
nor U14342 (N_14342,N_5049,N_9875);
nor U14343 (N_14343,N_7395,N_9996);
nand U14344 (N_14344,N_6324,N_6886);
or U14345 (N_14345,N_6095,N_5104);
and U14346 (N_14346,N_6157,N_8648);
nor U14347 (N_14347,N_6230,N_7889);
nor U14348 (N_14348,N_8683,N_5773);
xnor U14349 (N_14349,N_5974,N_5273);
or U14350 (N_14350,N_7487,N_9633);
or U14351 (N_14351,N_7841,N_8407);
and U14352 (N_14352,N_7058,N_6500);
or U14353 (N_14353,N_5428,N_5760);
or U14354 (N_14354,N_8350,N_8882);
nand U14355 (N_14355,N_7392,N_5161);
or U14356 (N_14356,N_6395,N_6451);
and U14357 (N_14357,N_8813,N_5771);
nand U14358 (N_14358,N_5905,N_9509);
xnor U14359 (N_14359,N_5862,N_6375);
nand U14360 (N_14360,N_8867,N_6872);
nand U14361 (N_14361,N_5968,N_6655);
or U14362 (N_14362,N_5112,N_6101);
nand U14363 (N_14363,N_6715,N_9187);
nor U14364 (N_14364,N_5337,N_8982);
nor U14365 (N_14365,N_5751,N_5215);
xor U14366 (N_14366,N_8437,N_7458);
nand U14367 (N_14367,N_7041,N_8740);
and U14368 (N_14368,N_5101,N_6078);
or U14369 (N_14369,N_6179,N_8366);
or U14370 (N_14370,N_7211,N_9811);
and U14371 (N_14371,N_6562,N_9718);
nor U14372 (N_14372,N_7469,N_8987);
or U14373 (N_14373,N_9167,N_7216);
nand U14374 (N_14374,N_8651,N_6201);
or U14375 (N_14375,N_5990,N_5512);
or U14376 (N_14376,N_9402,N_9825);
nor U14377 (N_14377,N_5716,N_6697);
nor U14378 (N_14378,N_7898,N_7701);
nand U14379 (N_14379,N_9235,N_9655);
nand U14380 (N_14380,N_9853,N_5026);
nand U14381 (N_14381,N_6190,N_7509);
nand U14382 (N_14382,N_5246,N_7122);
and U14383 (N_14383,N_6068,N_6637);
and U14384 (N_14384,N_6057,N_8379);
nor U14385 (N_14385,N_6628,N_7767);
nor U14386 (N_14386,N_5869,N_7730);
and U14387 (N_14387,N_7094,N_7389);
nor U14388 (N_14388,N_7581,N_6731);
nand U14389 (N_14389,N_7054,N_5770);
or U14390 (N_14390,N_9299,N_9761);
nor U14391 (N_14391,N_7112,N_7660);
nand U14392 (N_14392,N_8507,N_8696);
or U14393 (N_14393,N_9652,N_8598);
nand U14394 (N_14394,N_6085,N_7692);
nor U14395 (N_14395,N_9842,N_5614);
nand U14396 (N_14396,N_6671,N_5705);
nor U14397 (N_14397,N_6819,N_7251);
nor U14398 (N_14398,N_9594,N_8381);
and U14399 (N_14399,N_7004,N_8195);
nand U14400 (N_14400,N_9342,N_6760);
nand U14401 (N_14401,N_9247,N_8552);
nand U14402 (N_14402,N_7524,N_6736);
nor U14403 (N_14403,N_6123,N_7748);
or U14404 (N_14404,N_7415,N_7449);
or U14405 (N_14405,N_5417,N_7048);
nor U14406 (N_14406,N_7988,N_8848);
nor U14407 (N_14407,N_6050,N_5772);
nand U14408 (N_14408,N_8492,N_6018);
and U14409 (N_14409,N_7677,N_9834);
and U14410 (N_14410,N_6490,N_8691);
nor U14411 (N_14411,N_7591,N_7469);
and U14412 (N_14412,N_6652,N_6581);
or U14413 (N_14413,N_5621,N_7297);
and U14414 (N_14414,N_7190,N_7818);
nand U14415 (N_14415,N_9361,N_7737);
or U14416 (N_14416,N_7930,N_7384);
or U14417 (N_14417,N_6039,N_7713);
and U14418 (N_14418,N_9237,N_8816);
and U14419 (N_14419,N_8831,N_6705);
and U14420 (N_14420,N_5323,N_7325);
and U14421 (N_14421,N_9317,N_8691);
nor U14422 (N_14422,N_8754,N_9859);
nor U14423 (N_14423,N_9023,N_8044);
nor U14424 (N_14424,N_7139,N_6241);
or U14425 (N_14425,N_8736,N_9235);
or U14426 (N_14426,N_5829,N_8215);
and U14427 (N_14427,N_9714,N_7607);
nor U14428 (N_14428,N_7937,N_5047);
nor U14429 (N_14429,N_8355,N_5594);
or U14430 (N_14430,N_9095,N_8250);
and U14431 (N_14431,N_9355,N_9031);
nor U14432 (N_14432,N_8386,N_5465);
or U14433 (N_14433,N_7725,N_9598);
and U14434 (N_14434,N_8104,N_7023);
xnor U14435 (N_14435,N_5374,N_6024);
nor U14436 (N_14436,N_9448,N_6091);
nand U14437 (N_14437,N_7438,N_5095);
or U14438 (N_14438,N_7431,N_7988);
or U14439 (N_14439,N_6840,N_6920);
or U14440 (N_14440,N_9909,N_9500);
nand U14441 (N_14441,N_5046,N_5217);
and U14442 (N_14442,N_5974,N_7110);
or U14443 (N_14443,N_5065,N_8546);
nor U14444 (N_14444,N_6557,N_7210);
or U14445 (N_14445,N_9150,N_7055);
and U14446 (N_14446,N_7243,N_5106);
xor U14447 (N_14447,N_8822,N_9679);
and U14448 (N_14448,N_5143,N_6126);
nor U14449 (N_14449,N_5696,N_9396);
nand U14450 (N_14450,N_9352,N_6383);
nand U14451 (N_14451,N_8225,N_5383);
nand U14452 (N_14452,N_8673,N_8645);
xor U14453 (N_14453,N_9049,N_9120);
and U14454 (N_14454,N_7418,N_7946);
or U14455 (N_14455,N_5339,N_8085);
nor U14456 (N_14456,N_6785,N_5436);
and U14457 (N_14457,N_6876,N_8295);
nor U14458 (N_14458,N_9264,N_5852);
nor U14459 (N_14459,N_5792,N_7137);
or U14460 (N_14460,N_9963,N_7189);
nand U14461 (N_14461,N_6398,N_5783);
and U14462 (N_14462,N_7014,N_9161);
and U14463 (N_14463,N_6692,N_9064);
xnor U14464 (N_14464,N_6599,N_8322);
and U14465 (N_14465,N_8547,N_9421);
and U14466 (N_14466,N_7862,N_7808);
and U14467 (N_14467,N_6551,N_5609);
nor U14468 (N_14468,N_9725,N_7537);
and U14469 (N_14469,N_8585,N_9182);
or U14470 (N_14470,N_9843,N_9768);
and U14471 (N_14471,N_6163,N_7355);
nor U14472 (N_14472,N_7050,N_7078);
nor U14473 (N_14473,N_6213,N_8841);
nand U14474 (N_14474,N_6721,N_7612);
xor U14475 (N_14475,N_9416,N_8393);
nand U14476 (N_14476,N_5506,N_9385);
nand U14477 (N_14477,N_7928,N_7547);
nor U14478 (N_14478,N_6185,N_5967);
or U14479 (N_14479,N_5384,N_5239);
nand U14480 (N_14480,N_8817,N_9412);
or U14481 (N_14481,N_9237,N_7324);
nand U14482 (N_14482,N_6932,N_5713);
nand U14483 (N_14483,N_8517,N_5374);
or U14484 (N_14484,N_8225,N_7119);
nor U14485 (N_14485,N_7102,N_6546);
and U14486 (N_14486,N_6862,N_8663);
nor U14487 (N_14487,N_9829,N_9138);
or U14488 (N_14488,N_7631,N_5879);
nand U14489 (N_14489,N_8762,N_8864);
and U14490 (N_14490,N_5320,N_8368);
and U14491 (N_14491,N_5959,N_6219);
nor U14492 (N_14492,N_5229,N_5538);
or U14493 (N_14493,N_7971,N_5768);
or U14494 (N_14494,N_7862,N_8773);
or U14495 (N_14495,N_8956,N_6551);
nor U14496 (N_14496,N_9431,N_8235);
or U14497 (N_14497,N_6098,N_8346);
and U14498 (N_14498,N_5938,N_8646);
or U14499 (N_14499,N_8102,N_6447);
and U14500 (N_14500,N_7614,N_9212);
nor U14501 (N_14501,N_5574,N_7742);
nor U14502 (N_14502,N_9605,N_7044);
nand U14503 (N_14503,N_9152,N_5947);
nor U14504 (N_14504,N_8931,N_9485);
and U14505 (N_14505,N_9789,N_9615);
or U14506 (N_14506,N_9922,N_8762);
and U14507 (N_14507,N_5894,N_8245);
nand U14508 (N_14508,N_6167,N_9494);
nor U14509 (N_14509,N_6077,N_7404);
nor U14510 (N_14510,N_9236,N_6122);
nand U14511 (N_14511,N_7800,N_9822);
nor U14512 (N_14512,N_9748,N_5405);
and U14513 (N_14513,N_7237,N_6101);
and U14514 (N_14514,N_8094,N_8259);
or U14515 (N_14515,N_8671,N_7682);
nor U14516 (N_14516,N_8809,N_6193);
or U14517 (N_14517,N_6158,N_7862);
and U14518 (N_14518,N_8339,N_9709);
nor U14519 (N_14519,N_9166,N_5729);
and U14520 (N_14520,N_9995,N_5727);
nor U14521 (N_14521,N_8926,N_8228);
or U14522 (N_14522,N_8172,N_9540);
nor U14523 (N_14523,N_7353,N_7675);
nand U14524 (N_14524,N_8285,N_9718);
and U14525 (N_14525,N_7727,N_6755);
xor U14526 (N_14526,N_8127,N_9067);
and U14527 (N_14527,N_8181,N_8617);
nand U14528 (N_14528,N_9740,N_6218);
and U14529 (N_14529,N_9465,N_8185);
nor U14530 (N_14530,N_8961,N_6602);
nand U14531 (N_14531,N_8536,N_9032);
nor U14532 (N_14532,N_9380,N_9148);
or U14533 (N_14533,N_5368,N_7948);
xnor U14534 (N_14534,N_7701,N_9635);
nand U14535 (N_14535,N_9213,N_8608);
nand U14536 (N_14536,N_9388,N_7658);
or U14537 (N_14537,N_6317,N_7195);
and U14538 (N_14538,N_8663,N_9489);
or U14539 (N_14539,N_7049,N_9632);
nor U14540 (N_14540,N_6684,N_9852);
and U14541 (N_14541,N_6684,N_8274);
nand U14542 (N_14542,N_5391,N_8609);
or U14543 (N_14543,N_5478,N_8991);
nor U14544 (N_14544,N_8135,N_7871);
nand U14545 (N_14545,N_6385,N_6658);
nor U14546 (N_14546,N_5840,N_5187);
or U14547 (N_14547,N_9541,N_9988);
nand U14548 (N_14548,N_5491,N_5116);
nor U14549 (N_14549,N_6374,N_8664);
or U14550 (N_14550,N_7909,N_5599);
nor U14551 (N_14551,N_7927,N_6577);
and U14552 (N_14552,N_6150,N_6320);
and U14553 (N_14553,N_9529,N_9282);
nand U14554 (N_14554,N_6994,N_9183);
and U14555 (N_14555,N_8896,N_5284);
and U14556 (N_14556,N_8406,N_6021);
nor U14557 (N_14557,N_5925,N_9289);
nor U14558 (N_14558,N_9761,N_8988);
and U14559 (N_14559,N_6775,N_8035);
nand U14560 (N_14560,N_7257,N_5596);
and U14561 (N_14561,N_5711,N_5309);
or U14562 (N_14562,N_9494,N_5593);
and U14563 (N_14563,N_7930,N_5654);
or U14564 (N_14564,N_8649,N_6656);
or U14565 (N_14565,N_5031,N_8367);
nand U14566 (N_14566,N_7666,N_8186);
nand U14567 (N_14567,N_5155,N_6259);
nor U14568 (N_14568,N_6005,N_8908);
and U14569 (N_14569,N_7919,N_5247);
xnor U14570 (N_14570,N_5268,N_8418);
nor U14571 (N_14571,N_9938,N_5721);
or U14572 (N_14572,N_5365,N_7660);
nand U14573 (N_14573,N_9971,N_5023);
or U14574 (N_14574,N_9773,N_5120);
or U14575 (N_14575,N_7152,N_9716);
nand U14576 (N_14576,N_6777,N_5474);
or U14577 (N_14577,N_6663,N_9837);
nor U14578 (N_14578,N_9944,N_7150);
or U14579 (N_14579,N_7419,N_7473);
nand U14580 (N_14580,N_8982,N_5207);
nand U14581 (N_14581,N_7718,N_8908);
nor U14582 (N_14582,N_7247,N_8572);
nor U14583 (N_14583,N_9499,N_6386);
or U14584 (N_14584,N_5979,N_7810);
nand U14585 (N_14585,N_6998,N_5332);
nor U14586 (N_14586,N_9294,N_9820);
and U14587 (N_14587,N_7411,N_9838);
nand U14588 (N_14588,N_6718,N_9867);
or U14589 (N_14589,N_8464,N_7289);
or U14590 (N_14590,N_8341,N_7710);
and U14591 (N_14591,N_9342,N_8220);
nor U14592 (N_14592,N_9980,N_5656);
nor U14593 (N_14593,N_8128,N_9523);
and U14594 (N_14594,N_8432,N_5086);
and U14595 (N_14595,N_5445,N_6607);
nand U14596 (N_14596,N_5970,N_7944);
nor U14597 (N_14597,N_9687,N_7217);
nand U14598 (N_14598,N_5628,N_8410);
xor U14599 (N_14599,N_7248,N_7886);
nor U14600 (N_14600,N_9843,N_7331);
or U14601 (N_14601,N_9132,N_6400);
nand U14602 (N_14602,N_8886,N_5954);
nand U14603 (N_14603,N_6652,N_8557);
xor U14604 (N_14604,N_5768,N_6657);
nor U14605 (N_14605,N_5341,N_6004);
nand U14606 (N_14606,N_5805,N_6778);
or U14607 (N_14607,N_7313,N_6334);
nand U14608 (N_14608,N_7087,N_5631);
nor U14609 (N_14609,N_6015,N_7786);
and U14610 (N_14610,N_6556,N_5429);
nand U14611 (N_14611,N_7178,N_8855);
nand U14612 (N_14612,N_7380,N_9082);
nor U14613 (N_14613,N_7779,N_8700);
nand U14614 (N_14614,N_5434,N_5539);
nor U14615 (N_14615,N_8602,N_5851);
nor U14616 (N_14616,N_6712,N_6563);
nor U14617 (N_14617,N_8184,N_8217);
nand U14618 (N_14618,N_7585,N_6296);
nand U14619 (N_14619,N_9312,N_5461);
and U14620 (N_14620,N_7387,N_7799);
or U14621 (N_14621,N_7869,N_8150);
and U14622 (N_14622,N_9697,N_6690);
nand U14623 (N_14623,N_5604,N_5994);
and U14624 (N_14624,N_7409,N_7526);
nand U14625 (N_14625,N_9275,N_7961);
or U14626 (N_14626,N_9914,N_5383);
nor U14627 (N_14627,N_7737,N_6022);
or U14628 (N_14628,N_7525,N_8410);
nor U14629 (N_14629,N_5011,N_6317);
or U14630 (N_14630,N_6510,N_6299);
or U14631 (N_14631,N_9415,N_7594);
nor U14632 (N_14632,N_9076,N_6000);
or U14633 (N_14633,N_9126,N_7649);
or U14634 (N_14634,N_9916,N_9337);
or U14635 (N_14635,N_8244,N_6280);
and U14636 (N_14636,N_8835,N_7953);
nand U14637 (N_14637,N_9433,N_7145);
nor U14638 (N_14638,N_9103,N_7692);
nor U14639 (N_14639,N_5898,N_9548);
xor U14640 (N_14640,N_7537,N_9441);
or U14641 (N_14641,N_5776,N_8305);
nor U14642 (N_14642,N_9784,N_8353);
nand U14643 (N_14643,N_6692,N_8644);
xnor U14644 (N_14644,N_8108,N_5259);
nand U14645 (N_14645,N_6944,N_7716);
or U14646 (N_14646,N_8274,N_7210);
nand U14647 (N_14647,N_7372,N_9213);
nand U14648 (N_14648,N_8567,N_8333);
or U14649 (N_14649,N_6982,N_6940);
nor U14650 (N_14650,N_9761,N_8396);
nor U14651 (N_14651,N_9651,N_9388);
nor U14652 (N_14652,N_9710,N_5183);
and U14653 (N_14653,N_6839,N_9596);
nor U14654 (N_14654,N_9083,N_7528);
or U14655 (N_14655,N_8042,N_5578);
nor U14656 (N_14656,N_8774,N_8336);
and U14657 (N_14657,N_7463,N_5053);
nor U14658 (N_14658,N_5060,N_6900);
nand U14659 (N_14659,N_6709,N_7624);
or U14660 (N_14660,N_5453,N_6655);
nor U14661 (N_14661,N_9322,N_9227);
or U14662 (N_14662,N_7130,N_9694);
nor U14663 (N_14663,N_9359,N_8225);
nand U14664 (N_14664,N_8669,N_7295);
nor U14665 (N_14665,N_7728,N_8953);
nor U14666 (N_14666,N_8124,N_5927);
or U14667 (N_14667,N_8228,N_7225);
and U14668 (N_14668,N_7444,N_5609);
xnor U14669 (N_14669,N_8209,N_5388);
and U14670 (N_14670,N_5694,N_6862);
nor U14671 (N_14671,N_5087,N_7375);
or U14672 (N_14672,N_7985,N_6786);
or U14673 (N_14673,N_7957,N_7643);
or U14674 (N_14674,N_6874,N_8075);
nor U14675 (N_14675,N_7745,N_7262);
nor U14676 (N_14676,N_9823,N_9239);
or U14677 (N_14677,N_7748,N_9813);
or U14678 (N_14678,N_9116,N_7406);
or U14679 (N_14679,N_6929,N_7151);
or U14680 (N_14680,N_9433,N_7876);
nand U14681 (N_14681,N_9196,N_6113);
nor U14682 (N_14682,N_9723,N_6293);
and U14683 (N_14683,N_5994,N_6218);
and U14684 (N_14684,N_6315,N_6483);
nand U14685 (N_14685,N_9556,N_7930);
or U14686 (N_14686,N_9183,N_6107);
or U14687 (N_14687,N_5141,N_5948);
and U14688 (N_14688,N_7368,N_9621);
and U14689 (N_14689,N_5116,N_8133);
nor U14690 (N_14690,N_8517,N_6127);
nand U14691 (N_14691,N_9950,N_8080);
and U14692 (N_14692,N_5841,N_5659);
and U14693 (N_14693,N_8500,N_9607);
nor U14694 (N_14694,N_7079,N_5124);
nor U14695 (N_14695,N_7387,N_8444);
nand U14696 (N_14696,N_8278,N_7927);
nor U14697 (N_14697,N_6335,N_6167);
nor U14698 (N_14698,N_7141,N_9128);
or U14699 (N_14699,N_5494,N_5544);
nand U14700 (N_14700,N_5059,N_9312);
nor U14701 (N_14701,N_6625,N_5557);
and U14702 (N_14702,N_7739,N_5886);
and U14703 (N_14703,N_5075,N_8611);
or U14704 (N_14704,N_8140,N_5663);
and U14705 (N_14705,N_6625,N_9734);
or U14706 (N_14706,N_5427,N_6072);
or U14707 (N_14707,N_8112,N_6195);
nor U14708 (N_14708,N_9165,N_5392);
nor U14709 (N_14709,N_6748,N_7106);
nand U14710 (N_14710,N_8805,N_5794);
xnor U14711 (N_14711,N_6920,N_9468);
or U14712 (N_14712,N_9655,N_6046);
or U14713 (N_14713,N_9738,N_7664);
and U14714 (N_14714,N_7696,N_5708);
and U14715 (N_14715,N_9363,N_9865);
and U14716 (N_14716,N_6166,N_9261);
nor U14717 (N_14717,N_6005,N_5520);
nor U14718 (N_14718,N_8842,N_7870);
and U14719 (N_14719,N_8644,N_8488);
or U14720 (N_14720,N_7794,N_7613);
nand U14721 (N_14721,N_7069,N_5927);
or U14722 (N_14722,N_6852,N_9468);
or U14723 (N_14723,N_7859,N_7460);
and U14724 (N_14724,N_6055,N_8037);
and U14725 (N_14725,N_7790,N_5578);
nand U14726 (N_14726,N_6859,N_8481);
xnor U14727 (N_14727,N_5856,N_7744);
nor U14728 (N_14728,N_8593,N_7901);
and U14729 (N_14729,N_9620,N_9855);
and U14730 (N_14730,N_7487,N_6250);
nor U14731 (N_14731,N_7351,N_9632);
nor U14732 (N_14732,N_7932,N_6558);
nand U14733 (N_14733,N_5862,N_7275);
nor U14734 (N_14734,N_9814,N_5102);
nand U14735 (N_14735,N_7849,N_5872);
nor U14736 (N_14736,N_9178,N_9002);
nor U14737 (N_14737,N_5833,N_8641);
nand U14738 (N_14738,N_9860,N_9470);
and U14739 (N_14739,N_9165,N_7716);
or U14740 (N_14740,N_5796,N_7423);
and U14741 (N_14741,N_7189,N_8999);
or U14742 (N_14742,N_5355,N_6896);
or U14743 (N_14743,N_6755,N_5874);
or U14744 (N_14744,N_5357,N_8837);
and U14745 (N_14745,N_6270,N_6922);
or U14746 (N_14746,N_8201,N_8162);
nand U14747 (N_14747,N_8967,N_5896);
nor U14748 (N_14748,N_7941,N_9869);
or U14749 (N_14749,N_7595,N_5263);
or U14750 (N_14750,N_6546,N_9862);
or U14751 (N_14751,N_5089,N_8243);
and U14752 (N_14752,N_9168,N_7081);
nor U14753 (N_14753,N_6871,N_5102);
nand U14754 (N_14754,N_5615,N_8968);
or U14755 (N_14755,N_5416,N_5978);
xor U14756 (N_14756,N_8613,N_8544);
and U14757 (N_14757,N_8602,N_6752);
nor U14758 (N_14758,N_8613,N_9098);
nor U14759 (N_14759,N_8254,N_9732);
nand U14760 (N_14760,N_5771,N_9205);
or U14761 (N_14761,N_6161,N_6893);
or U14762 (N_14762,N_9528,N_9306);
nor U14763 (N_14763,N_6780,N_6368);
nand U14764 (N_14764,N_7106,N_8392);
nor U14765 (N_14765,N_8213,N_8556);
nand U14766 (N_14766,N_7028,N_9483);
and U14767 (N_14767,N_6517,N_7703);
nand U14768 (N_14768,N_8980,N_6109);
and U14769 (N_14769,N_7496,N_8573);
nor U14770 (N_14770,N_9228,N_9124);
xor U14771 (N_14771,N_5568,N_9832);
nand U14772 (N_14772,N_7364,N_7717);
or U14773 (N_14773,N_5800,N_7109);
and U14774 (N_14774,N_7629,N_5009);
and U14775 (N_14775,N_6781,N_9407);
and U14776 (N_14776,N_9482,N_6838);
nor U14777 (N_14777,N_9580,N_7709);
xnor U14778 (N_14778,N_5383,N_6103);
nand U14779 (N_14779,N_9567,N_6101);
nand U14780 (N_14780,N_9981,N_9914);
or U14781 (N_14781,N_9689,N_6971);
or U14782 (N_14782,N_5288,N_8142);
and U14783 (N_14783,N_7777,N_9924);
nor U14784 (N_14784,N_8775,N_7084);
and U14785 (N_14785,N_8002,N_7027);
nor U14786 (N_14786,N_5693,N_6668);
and U14787 (N_14787,N_7965,N_8331);
or U14788 (N_14788,N_6564,N_7918);
and U14789 (N_14789,N_5593,N_7208);
nor U14790 (N_14790,N_8646,N_8723);
or U14791 (N_14791,N_8999,N_5694);
or U14792 (N_14792,N_9563,N_7295);
or U14793 (N_14793,N_7451,N_9056);
and U14794 (N_14794,N_5668,N_5880);
nor U14795 (N_14795,N_8862,N_5614);
and U14796 (N_14796,N_6230,N_7494);
and U14797 (N_14797,N_7796,N_5641);
or U14798 (N_14798,N_6259,N_6246);
nand U14799 (N_14799,N_5359,N_7875);
and U14800 (N_14800,N_6252,N_6204);
or U14801 (N_14801,N_5222,N_6904);
xnor U14802 (N_14802,N_9692,N_6830);
nand U14803 (N_14803,N_9964,N_7640);
nand U14804 (N_14804,N_8605,N_5245);
nor U14805 (N_14805,N_6211,N_7503);
nand U14806 (N_14806,N_8752,N_6044);
or U14807 (N_14807,N_9670,N_5510);
nand U14808 (N_14808,N_9823,N_7396);
and U14809 (N_14809,N_6292,N_5914);
nand U14810 (N_14810,N_7274,N_6631);
nor U14811 (N_14811,N_6674,N_7478);
and U14812 (N_14812,N_6944,N_7129);
nand U14813 (N_14813,N_9821,N_5656);
nor U14814 (N_14814,N_5289,N_8451);
nor U14815 (N_14815,N_8172,N_8568);
nor U14816 (N_14816,N_9120,N_9299);
and U14817 (N_14817,N_9561,N_6684);
and U14818 (N_14818,N_9391,N_9842);
and U14819 (N_14819,N_9144,N_5035);
nand U14820 (N_14820,N_7158,N_6255);
and U14821 (N_14821,N_9353,N_8670);
nor U14822 (N_14822,N_6823,N_7587);
or U14823 (N_14823,N_7747,N_7866);
nand U14824 (N_14824,N_7149,N_9830);
nand U14825 (N_14825,N_7063,N_7472);
xor U14826 (N_14826,N_6645,N_7164);
nand U14827 (N_14827,N_7902,N_8886);
nor U14828 (N_14828,N_5526,N_5002);
xnor U14829 (N_14829,N_7135,N_9408);
or U14830 (N_14830,N_7465,N_6257);
nand U14831 (N_14831,N_7544,N_5647);
nor U14832 (N_14832,N_6554,N_7429);
and U14833 (N_14833,N_7009,N_5736);
nand U14834 (N_14834,N_9395,N_7641);
nand U14835 (N_14835,N_6764,N_5429);
xnor U14836 (N_14836,N_9234,N_5066);
nand U14837 (N_14837,N_8682,N_6140);
or U14838 (N_14838,N_7296,N_9485);
or U14839 (N_14839,N_9950,N_9287);
and U14840 (N_14840,N_6276,N_6849);
or U14841 (N_14841,N_5233,N_8167);
or U14842 (N_14842,N_5680,N_9304);
or U14843 (N_14843,N_8126,N_7674);
or U14844 (N_14844,N_7660,N_9839);
and U14845 (N_14845,N_6850,N_7851);
nor U14846 (N_14846,N_8454,N_8549);
nand U14847 (N_14847,N_7835,N_8717);
or U14848 (N_14848,N_9409,N_9728);
and U14849 (N_14849,N_6805,N_7583);
nor U14850 (N_14850,N_8412,N_7650);
xnor U14851 (N_14851,N_5119,N_5057);
nand U14852 (N_14852,N_9915,N_7186);
and U14853 (N_14853,N_8938,N_9164);
and U14854 (N_14854,N_6078,N_5588);
or U14855 (N_14855,N_5339,N_7105);
and U14856 (N_14856,N_6206,N_8846);
nor U14857 (N_14857,N_7850,N_7657);
nand U14858 (N_14858,N_9309,N_9566);
or U14859 (N_14859,N_8225,N_7475);
nor U14860 (N_14860,N_7785,N_8921);
or U14861 (N_14861,N_5984,N_5164);
or U14862 (N_14862,N_8678,N_6965);
nor U14863 (N_14863,N_6987,N_5635);
and U14864 (N_14864,N_8241,N_7837);
nand U14865 (N_14865,N_7701,N_8261);
nor U14866 (N_14866,N_7796,N_5847);
nand U14867 (N_14867,N_7545,N_8553);
and U14868 (N_14868,N_6123,N_5110);
nand U14869 (N_14869,N_5159,N_8887);
nor U14870 (N_14870,N_6793,N_8808);
and U14871 (N_14871,N_6776,N_7707);
nor U14872 (N_14872,N_8576,N_5199);
and U14873 (N_14873,N_6975,N_5412);
or U14874 (N_14874,N_9697,N_9756);
or U14875 (N_14875,N_8785,N_8932);
nand U14876 (N_14876,N_6346,N_6184);
nor U14877 (N_14877,N_8012,N_9461);
or U14878 (N_14878,N_8169,N_5875);
and U14879 (N_14879,N_5107,N_6004);
nor U14880 (N_14880,N_8869,N_8326);
and U14881 (N_14881,N_5363,N_6012);
and U14882 (N_14882,N_9678,N_6391);
and U14883 (N_14883,N_6224,N_8692);
and U14884 (N_14884,N_9985,N_6155);
nor U14885 (N_14885,N_9729,N_9431);
and U14886 (N_14886,N_7247,N_8305);
nand U14887 (N_14887,N_7793,N_9756);
and U14888 (N_14888,N_5374,N_5762);
or U14889 (N_14889,N_9159,N_7941);
and U14890 (N_14890,N_9370,N_9562);
nand U14891 (N_14891,N_6986,N_6009);
and U14892 (N_14892,N_6367,N_8666);
or U14893 (N_14893,N_7060,N_7433);
nand U14894 (N_14894,N_7693,N_7964);
xor U14895 (N_14895,N_7631,N_8394);
and U14896 (N_14896,N_7037,N_7682);
nor U14897 (N_14897,N_6560,N_6753);
nand U14898 (N_14898,N_5371,N_7565);
nor U14899 (N_14899,N_5916,N_6324);
nor U14900 (N_14900,N_9451,N_6196);
nor U14901 (N_14901,N_9465,N_5464);
nand U14902 (N_14902,N_8752,N_9474);
nand U14903 (N_14903,N_8451,N_8288);
nor U14904 (N_14904,N_8687,N_5010);
or U14905 (N_14905,N_6416,N_8923);
and U14906 (N_14906,N_8295,N_5356);
nor U14907 (N_14907,N_5017,N_9572);
nand U14908 (N_14908,N_5396,N_9813);
and U14909 (N_14909,N_8512,N_8089);
and U14910 (N_14910,N_9040,N_6301);
nand U14911 (N_14911,N_9685,N_8656);
nor U14912 (N_14912,N_5688,N_6609);
and U14913 (N_14913,N_7388,N_8180);
or U14914 (N_14914,N_5425,N_5901);
or U14915 (N_14915,N_9732,N_6463);
and U14916 (N_14916,N_8199,N_8366);
nand U14917 (N_14917,N_5738,N_8512);
or U14918 (N_14918,N_7352,N_6250);
nor U14919 (N_14919,N_8203,N_5279);
nand U14920 (N_14920,N_7873,N_7188);
nand U14921 (N_14921,N_8330,N_8132);
nand U14922 (N_14922,N_8993,N_8509);
or U14923 (N_14923,N_8934,N_9891);
and U14924 (N_14924,N_5821,N_7371);
nand U14925 (N_14925,N_7740,N_7026);
nand U14926 (N_14926,N_8743,N_7132);
or U14927 (N_14927,N_7460,N_8755);
or U14928 (N_14928,N_5587,N_7136);
or U14929 (N_14929,N_9509,N_7669);
nand U14930 (N_14930,N_5720,N_5297);
nand U14931 (N_14931,N_5493,N_5876);
nand U14932 (N_14932,N_7548,N_9925);
or U14933 (N_14933,N_7731,N_6140);
nand U14934 (N_14934,N_6471,N_7666);
nor U14935 (N_14935,N_8876,N_9969);
or U14936 (N_14936,N_6625,N_8604);
or U14937 (N_14937,N_6694,N_6444);
or U14938 (N_14938,N_5037,N_8367);
nor U14939 (N_14939,N_8108,N_8879);
nand U14940 (N_14940,N_7630,N_7284);
nand U14941 (N_14941,N_9153,N_9001);
nand U14942 (N_14942,N_6737,N_7749);
nand U14943 (N_14943,N_5456,N_7174);
nor U14944 (N_14944,N_9802,N_9780);
or U14945 (N_14945,N_9205,N_8126);
nand U14946 (N_14946,N_5937,N_7883);
and U14947 (N_14947,N_9358,N_8286);
and U14948 (N_14948,N_8133,N_8255);
xnor U14949 (N_14949,N_7627,N_8655);
or U14950 (N_14950,N_8147,N_9851);
nand U14951 (N_14951,N_9352,N_7802);
and U14952 (N_14952,N_5815,N_7471);
nor U14953 (N_14953,N_6994,N_5031);
and U14954 (N_14954,N_8514,N_5834);
and U14955 (N_14955,N_6045,N_6603);
nand U14956 (N_14956,N_6214,N_6731);
or U14957 (N_14957,N_6688,N_6041);
nand U14958 (N_14958,N_9336,N_7875);
xor U14959 (N_14959,N_6766,N_8369);
or U14960 (N_14960,N_7982,N_9679);
xor U14961 (N_14961,N_7781,N_9824);
or U14962 (N_14962,N_5463,N_8880);
nor U14963 (N_14963,N_6362,N_5501);
nor U14964 (N_14964,N_5589,N_7300);
nand U14965 (N_14965,N_7435,N_6717);
nor U14966 (N_14966,N_5317,N_8091);
nor U14967 (N_14967,N_5289,N_5166);
nor U14968 (N_14968,N_7327,N_7342);
nand U14969 (N_14969,N_8516,N_9900);
or U14970 (N_14970,N_6410,N_5655);
or U14971 (N_14971,N_8921,N_9442);
or U14972 (N_14972,N_6005,N_8644);
or U14973 (N_14973,N_7059,N_8652);
and U14974 (N_14974,N_9897,N_7882);
nand U14975 (N_14975,N_8257,N_5419);
and U14976 (N_14976,N_8478,N_8852);
nor U14977 (N_14977,N_5851,N_6465);
and U14978 (N_14978,N_8180,N_5162);
nand U14979 (N_14979,N_8829,N_5323);
nand U14980 (N_14980,N_5354,N_9766);
nand U14981 (N_14981,N_8134,N_9712);
nor U14982 (N_14982,N_9194,N_6347);
nor U14983 (N_14983,N_6889,N_8720);
nand U14984 (N_14984,N_9827,N_7057);
xnor U14985 (N_14985,N_9250,N_5859);
nor U14986 (N_14986,N_6060,N_6244);
nand U14987 (N_14987,N_6848,N_8741);
and U14988 (N_14988,N_5381,N_5499);
and U14989 (N_14989,N_5675,N_5554);
or U14990 (N_14990,N_8562,N_6378);
and U14991 (N_14991,N_7673,N_7679);
xor U14992 (N_14992,N_9372,N_8736);
nor U14993 (N_14993,N_9043,N_5269);
nand U14994 (N_14994,N_7404,N_6260);
nand U14995 (N_14995,N_5499,N_7180);
and U14996 (N_14996,N_6441,N_7238);
xnor U14997 (N_14997,N_9772,N_7661);
nand U14998 (N_14998,N_6572,N_8527);
or U14999 (N_14999,N_5558,N_8372);
nor U15000 (N_15000,N_13456,N_14029);
nor U15001 (N_15001,N_12888,N_10094);
or U15002 (N_15002,N_14371,N_14142);
and U15003 (N_15003,N_12873,N_11416);
nor U15004 (N_15004,N_14426,N_14849);
nor U15005 (N_15005,N_11759,N_10228);
and U15006 (N_15006,N_13058,N_12774);
or U15007 (N_15007,N_10136,N_14380);
nor U15008 (N_15008,N_14360,N_14051);
or U15009 (N_15009,N_14798,N_14054);
nand U15010 (N_15010,N_11527,N_11976);
and U15011 (N_15011,N_13093,N_10360);
nand U15012 (N_15012,N_13949,N_13143);
or U15013 (N_15013,N_14555,N_14318);
xor U15014 (N_15014,N_12977,N_14195);
or U15015 (N_15015,N_13596,N_10982);
or U15016 (N_15016,N_13752,N_11870);
and U15017 (N_15017,N_13854,N_14329);
and U15018 (N_15018,N_13794,N_11529);
or U15019 (N_15019,N_10948,N_12872);
xnor U15020 (N_15020,N_13101,N_14908);
nor U15021 (N_15021,N_14560,N_11448);
nor U15022 (N_15022,N_11760,N_10011);
nand U15023 (N_15023,N_13476,N_13386);
nor U15024 (N_15024,N_10915,N_13430);
or U15025 (N_15025,N_12428,N_14885);
and U15026 (N_15026,N_10677,N_14132);
nand U15027 (N_15027,N_10161,N_12999);
or U15028 (N_15028,N_12060,N_12418);
nand U15029 (N_15029,N_14053,N_12221);
xnor U15030 (N_15030,N_12799,N_11902);
and U15031 (N_15031,N_14178,N_13076);
or U15032 (N_15032,N_14827,N_12827);
nand U15033 (N_15033,N_13303,N_14149);
nor U15034 (N_15034,N_11302,N_14543);
nor U15035 (N_15035,N_13384,N_14331);
or U15036 (N_15036,N_11815,N_12082);
and U15037 (N_15037,N_10582,N_12532);
and U15038 (N_15038,N_12416,N_12589);
nand U15039 (N_15039,N_10122,N_14642);
nor U15040 (N_15040,N_11653,N_10601);
nor U15041 (N_15041,N_13610,N_13904);
nor U15042 (N_15042,N_12562,N_13340);
nand U15043 (N_15043,N_11192,N_13919);
and U15044 (N_15044,N_11425,N_10519);
and U15045 (N_15045,N_14205,N_11659);
and U15046 (N_15046,N_11323,N_11668);
and U15047 (N_15047,N_11547,N_11304);
and U15048 (N_15048,N_12363,N_13804);
nor U15049 (N_15049,N_12519,N_14410);
nor U15050 (N_15050,N_13588,N_10637);
and U15051 (N_15051,N_12851,N_12796);
nand U15052 (N_15052,N_13069,N_11288);
and U15053 (N_15053,N_13531,N_13522);
nor U15054 (N_15054,N_10056,N_11827);
or U15055 (N_15055,N_10114,N_13265);
nand U15056 (N_15056,N_11432,N_10185);
nor U15057 (N_15057,N_11266,N_12741);
or U15058 (N_15058,N_11402,N_11142);
and U15059 (N_15059,N_13328,N_10607);
nor U15060 (N_15060,N_11545,N_10709);
or U15061 (N_15061,N_13879,N_14871);
nor U15062 (N_15062,N_10631,N_11755);
or U15063 (N_15063,N_11574,N_12693);
or U15064 (N_15064,N_14981,N_12928);
nand U15065 (N_15065,N_11280,N_13662);
or U15066 (N_15066,N_10788,N_10033);
nor U15067 (N_15067,N_14875,N_11630);
nor U15068 (N_15068,N_13591,N_10400);
or U15069 (N_15069,N_10373,N_10936);
and U15070 (N_15070,N_14946,N_10097);
nand U15071 (N_15071,N_13418,N_12305);
or U15072 (N_15072,N_13862,N_12780);
nor U15073 (N_15073,N_11214,N_14203);
or U15074 (N_15074,N_11235,N_14491);
nand U15075 (N_15075,N_11991,N_13033);
nor U15076 (N_15076,N_10079,N_11049);
or U15077 (N_15077,N_13860,N_12235);
nand U15078 (N_15078,N_14997,N_12571);
and U15079 (N_15079,N_12219,N_11374);
nor U15080 (N_15080,N_14341,N_11460);
nand U15081 (N_15081,N_10213,N_11982);
nand U15082 (N_15082,N_12987,N_14892);
nor U15083 (N_15083,N_12047,N_13491);
or U15084 (N_15084,N_13471,N_10063);
nand U15085 (N_15085,N_10450,N_12370);
and U15086 (N_15086,N_12195,N_12243);
or U15087 (N_15087,N_10370,N_10385);
nand U15088 (N_15088,N_14193,N_12156);
and U15089 (N_15089,N_14277,N_12016);
nand U15090 (N_15090,N_14930,N_14565);
nor U15091 (N_15091,N_11946,N_14514);
and U15092 (N_15092,N_10473,N_10554);
and U15093 (N_15093,N_11826,N_11305);
and U15094 (N_15094,N_12988,N_13912);
or U15095 (N_15095,N_12205,N_11556);
nand U15096 (N_15096,N_13635,N_12509);
nand U15097 (N_15097,N_12770,N_14769);
nor U15098 (N_15098,N_13541,N_13281);
nor U15099 (N_15099,N_13646,N_11297);
and U15100 (N_15100,N_13440,N_14264);
and U15101 (N_15101,N_14084,N_13605);
and U15102 (N_15102,N_10696,N_14335);
and U15103 (N_15103,N_14614,N_13836);
nor U15104 (N_15104,N_11030,N_12289);
nor U15105 (N_15105,N_14472,N_14839);
or U15106 (N_15106,N_14759,N_13562);
or U15107 (N_15107,N_13323,N_10210);
nor U15108 (N_15108,N_13931,N_12450);
or U15109 (N_15109,N_11604,N_14206);
nor U15110 (N_15110,N_12884,N_13208);
or U15111 (N_15111,N_11121,N_11157);
and U15112 (N_15112,N_14237,N_13165);
or U15113 (N_15113,N_12180,N_13917);
nand U15114 (N_15114,N_13630,N_13015);
or U15115 (N_15115,N_10091,N_13393);
nand U15116 (N_15116,N_13296,N_13321);
or U15117 (N_15117,N_10433,N_12762);
nand U15118 (N_15118,N_11639,N_10626);
xnor U15119 (N_15119,N_13047,N_11295);
or U15120 (N_15120,N_10920,N_13534);
or U15121 (N_15121,N_12536,N_11600);
and U15122 (N_15122,N_14461,N_13700);
nor U15123 (N_15123,N_13148,N_13188);
and U15124 (N_15124,N_13008,N_14876);
nor U15125 (N_15125,N_11593,N_14435);
nand U15126 (N_15126,N_14310,N_11511);
or U15127 (N_15127,N_10479,N_11125);
nand U15128 (N_15128,N_13654,N_10883);
nand U15129 (N_15129,N_12169,N_12747);
nor U15130 (N_15130,N_13790,N_10415);
and U15131 (N_15131,N_12614,N_10892);
nor U15132 (N_15132,N_11781,N_12790);
or U15133 (N_15133,N_11013,N_14397);
or U15134 (N_15134,N_11798,N_10065);
nand U15135 (N_15135,N_10076,N_13767);
nand U15136 (N_15136,N_14504,N_13470);
or U15137 (N_15137,N_12506,N_12283);
nor U15138 (N_15138,N_10711,N_14372);
and U15139 (N_15139,N_10869,N_11405);
and U15140 (N_15140,N_12329,N_11139);
nand U15141 (N_15141,N_11627,N_12225);
and U15142 (N_15142,N_11043,N_11813);
or U15143 (N_15143,N_10113,N_11865);
or U15144 (N_15144,N_11223,N_14370);
or U15145 (N_15145,N_11356,N_11825);
or U15146 (N_15146,N_13315,N_10060);
and U15147 (N_15147,N_11528,N_11501);
nor U15148 (N_15148,N_11033,N_11227);
nand U15149 (N_15149,N_10808,N_13335);
and U15150 (N_15150,N_13739,N_11398);
nand U15151 (N_15151,N_14966,N_11892);
or U15152 (N_15152,N_12037,N_10831);
and U15153 (N_15153,N_11924,N_11059);
and U15154 (N_15154,N_14076,N_11829);
nand U15155 (N_15155,N_11099,N_13308);
nand U15156 (N_15156,N_14421,N_12782);
nor U15157 (N_15157,N_10770,N_11480);
and U15158 (N_15158,N_14546,N_14399);
or U15159 (N_15159,N_11393,N_12475);
or U15160 (N_15160,N_11997,N_14141);
nand U15161 (N_15161,N_12193,N_13560);
nor U15162 (N_15162,N_14704,N_10684);
and U15163 (N_15163,N_12278,N_13016);
or U15164 (N_15164,N_12044,N_11419);
or U15165 (N_15165,N_12981,N_13975);
or U15166 (N_15166,N_14446,N_11281);
or U15167 (N_15167,N_10735,N_11621);
or U15168 (N_15168,N_13811,N_10591);
nand U15169 (N_15169,N_12633,N_10769);
and U15170 (N_15170,N_12396,N_12526);
nor U15171 (N_15171,N_11379,N_11625);
or U15172 (N_15172,N_14459,N_10071);
or U15173 (N_15173,N_13273,N_13564);
or U15174 (N_15174,N_13390,N_10988);
nor U15175 (N_15175,N_11298,N_14760);
nor U15176 (N_15176,N_12568,N_11261);
nor U15177 (N_15177,N_11313,N_11736);
or U15178 (N_15178,N_12802,N_14409);
and U15179 (N_15179,N_14602,N_12678);
nor U15180 (N_15180,N_10886,N_12594);
or U15181 (N_15181,N_11417,N_10275);
and U15182 (N_15182,N_12058,N_11819);
and U15183 (N_15183,N_13784,N_10764);
or U15184 (N_15184,N_11749,N_12191);
or U15185 (N_15185,N_11536,N_12876);
or U15186 (N_15186,N_11514,N_12266);
nor U15187 (N_15187,N_10043,N_10317);
nor U15188 (N_15188,N_11381,N_12912);
or U15189 (N_15189,N_11190,N_11628);
nand U15190 (N_15190,N_12212,N_14398);
nor U15191 (N_15191,N_12488,N_12330);
or U15192 (N_15192,N_11583,N_10682);
and U15193 (N_15193,N_10296,N_12164);
and U15194 (N_15194,N_13114,N_12875);
or U15195 (N_15195,N_13758,N_13641);
or U15196 (N_15196,N_13859,N_14775);
nand U15197 (N_15197,N_13771,N_11470);
and U15198 (N_15198,N_12901,N_11029);
nand U15199 (N_15199,N_10146,N_14146);
nor U15200 (N_15200,N_14953,N_13307);
and U15201 (N_15201,N_12449,N_14732);
and U15202 (N_15202,N_12182,N_14117);
nor U15203 (N_15203,N_14327,N_13352);
nand U15204 (N_15204,N_14844,N_11719);
or U15205 (N_15205,N_13978,N_11040);
nand U15206 (N_15206,N_11582,N_11775);
nand U15207 (N_15207,N_11147,N_14973);
nand U15208 (N_15208,N_13104,N_10702);
or U15209 (N_15209,N_11045,N_11879);
and U15210 (N_15210,N_10045,N_12625);
nor U15211 (N_15211,N_13801,N_11727);
nand U15212 (N_15212,N_11874,N_13736);
or U15213 (N_15213,N_12096,N_13772);
or U15214 (N_15214,N_13452,N_12220);
nand U15215 (N_15215,N_13251,N_12099);
nor U15216 (N_15216,N_14626,N_11351);
xnor U15217 (N_15217,N_13220,N_14354);
or U15218 (N_15218,N_12832,N_12391);
nor U15219 (N_15219,N_12337,N_12621);
nand U15220 (N_15220,N_11433,N_12640);
nand U15221 (N_15221,N_10112,N_13398);
or U15222 (N_15222,N_11129,N_14214);
or U15223 (N_15223,N_12176,N_11680);
nor U15224 (N_15224,N_12319,N_13294);
or U15225 (N_15225,N_14692,N_10880);
nand U15226 (N_15226,N_13462,N_11041);
nand U15227 (N_15227,N_14806,N_13995);
and U15228 (N_15228,N_12006,N_12447);
xor U15229 (N_15229,N_12309,N_11489);
nor U15230 (N_15230,N_10145,N_12436);
nand U15231 (N_15231,N_11085,N_11757);
nor U15232 (N_15232,N_14893,N_10566);
nor U15233 (N_15233,N_14709,N_13791);
or U15234 (N_15234,N_14537,N_11786);
xnor U15235 (N_15235,N_13774,N_10881);
nor U15236 (N_15236,N_11250,N_12853);
and U15237 (N_15237,N_11575,N_14025);
nand U15238 (N_15238,N_10587,N_14058);
and U15239 (N_15239,N_13117,N_11932);
nand U15240 (N_15240,N_14328,N_10124);
or U15241 (N_15241,N_13505,N_14506);
and U15242 (N_15242,N_14616,N_13234);
nand U15243 (N_15243,N_13619,N_12073);
or U15244 (N_15244,N_12024,N_14306);
nor U15245 (N_15245,N_12247,N_12575);
nand U15246 (N_15246,N_12124,N_11439);
nor U15247 (N_15247,N_14617,N_12493);
nand U15248 (N_15248,N_12179,N_10812);
or U15249 (N_15249,N_14005,N_10675);
and U15250 (N_15250,N_14168,N_10331);
nor U15251 (N_15251,N_10730,N_13886);
and U15252 (N_15252,N_11221,N_12954);
xnor U15253 (N_15253,N_11360,N_11174);
and U15254 (N_15254,N_12281,N_11116);
or U15255 (N_15255,N_13049,N_12929);
and U15256 (N_15256,N_12542,N_14382);
or U15257 (N_15257,N_13142,N_14803);
and U15258 (N_15258,N_10194,N_14088);
nor U15259 (N_15259,N_13345,N_11361);
or U15260 (N_15260,N_14137,N_10149);
nor U15261 (N_15261,N_13814,N_14119);
nand U15262 (N_15262,N_13403,N_12445);
or U15263 (N_15263,N_10939,N_13996);
or U15264 (N_15264,N_12472,N_12087);
and U15265 (N_15265,N_14162,N_12838);
or U15266 (N_15266,N_12223,N_12806);
and U15267 (N_15267,N_13818,N_12812);
nand U15268 (N_15268,N_14972,N_13834);
or U15269 (N_15269,N_10050,N_13215);
nor U15270 (N_15270,N_10392,N_13973);
or U15271 (N_15271,N_12246,N_11654);
nand U15272 (N_15272,N_10249,N_14585);
and U15273 (N_15273,N_10902,N_11770);
or U15274 (N_15274,N_10109,N_12367);
and U15275 (N_15275,N_14431,N_12053);
nor U15276 (N_15276,N_13622,N_14089);
nor U15277 (N_15277,N_12540,N_11560);
or U15278 (N_15278,N_12725,N_13918);
or U15279 (N_15279,N_12000,N_11367);
and U15280 (N_15280,N_10263,N_12376);
and U15281 (N_15281,N_11595,N_14391);
or U15282 (N_15282,N_11761,N_11546);
nor U15283 (N_15283,N_13813,N_14407);
or U15284 (N_15284,N_10285,N_12446);
or U15285 (N_15285,N_10268,N_11820);
nand U15286 (N_15286,N_14439,N_13029);
or U15287 (N_15287,N_13399,N_12297);
or U15288 (N_15288,N_11024,N_11065);
nand U15289 (N_15289,N_11685,N_11996);
nor U15290 (N_15290,N_10553,N_13846);
xor U15291 (N_15291,N_10064,N_13540);
nand U15292 (N_15292,N_10190,N_11123);
nor U15293 (N_15293,N_13233,N_14877);
nor U15294 (N_15294,N_12545,N_10260);
nor U15295 (N_15295,N_10672,N_11310);
nor U15296 (N_15296,N_10822,N_10496);
nand U15297 (N_15297,N_12383,N_13124);
or U15298 (N_15298,N_10362,N_13503);
nand U15299 (N_15299,N_12649,N_10652);
nand U15300 (N_15300,N_14252,N_11063);
and U15301 (N_15301,N_10817,N_13863);
nor U15302 (N_15302,N_12819,N_10261);
nand U15303 (N_15303,N_11636,N_11275);
and U15304 (N_15304,N_13036,N_11390);
nand U15305 (N_15305,N_10242,N_13937);
nand U15306 (N_15306,N_11316,N_14448);
nand U15307 (N_15307,N_10854,N_11434);
and U15308 (N_15308,N_14753,N_10075);
nand U15309 (N_15309,N_12951,N_13751);
nand U15310 (N_15310,N_14023,N_11741);
or U15311 (N_15311,N_13777,N_13329);
nand U15312 (N_15312,N_10782,N_12910);
and U15313 (N_15313,N_12668,N_14405);
and U15314 (N_15314,N_12117,N_13643);
nand U15315 (N_15315,N_13785,N_13547);
or U15316 (N_15316,N_13759,N_13364);
and U15317 (N_15317,N_10353,N_12320);
and U15318 (N_15318,N_14477,N_12626);
nand U15319 (N_15319,N_13686,N_12325);
nand U15320 (N_15320,N_11590,N_10429);
nand U15321 (N_15321,N_12611,N_10120);
nor U15322 (N_15322,N_12586,N_10690);
nand U15323 (N_15323,N_14682,N_11591);
and U15324 (N_15324,N_13999,N_14796);
nand U15325 (N_15325,N_14569,N_14045);
and U15326 (N_15326,N_14180,N_12345);
or U15327 (N_15327,N_11633,N_14699);
xor U15328 (N_15328,N_11959,N_10164);
xor U15329 (N_15329,N_13874,N_14333);
or U15330 (N_15330,N_12068,N_13652);
and U15331 (N_15331,N_13181,N_10171);
or U15332 (N_15332,N_11472,N_14151);
nor U15333 (N_15333,N_14826,N_13821);
and U15334 (N_15334,N_12271,N_11696);
nand U15335 (N_15335,N_13237,N_13439);
and U15336 (N_15336,N_11388,N_10621);
and U15337 (N_15337,N_10107,N_13623);
or U15338 (N_15338,N_13506,N_14007);
and U15339 (N_15339,N_12482,N_13467);
nor U15340 (N_15340,N_12997,N_11420);
nand U15341 (N_15341,N_11004,N_13783);
and U15342 (N_15342,N_10633,N_13800);
nand U15343 (N_15343,N_10384,N_11601);
or U15344 (N_15344,N_13437,N_12946);
nor U15345 (N_15345,N_14475,N_11913);
and U15346 (N_15346,N_14152,N_10907);
or U15347 (N_15347,N_13896,N_11457);
or U15348 (N_15348,N_11651,N_11073);
nand U15349 (N_15349,N_11833,N_13450);
nand U15350 (N_15350,N_12761,N_13232);
and U15351 (N_15351,N_13461,N_11118);
nand U15352 (N_15352,N_14046,N_12467);
or U15353 (N_15353,N_14735,N_13589);
nor U15354 (N_15354,N_14624,N_14761);
xor U15355 (N_15355,N_10443,N_10932);
and U15356 (N_15356,N_14884,N_12142);
and U15357 (N_15357,N_13548,N_10643);
and U15358 (N_15358,N_11688,N_11692);
and U15359 (N_15359,N_14198,N_10444);
nor U15360 (N_15360,N_12713,N_12809);
nor U15361 (N_15361,N_10090,N_14590);
and U15362 (N_15362,N_12566,N_13414);
and U15363 (N_15363,N_10102,N_12279);
nand U15364 (N_15364,N_10603,N_12676);
and U15365 (N_15365,N_10466,N_10044);
and U15366 (N_15366,N_13536,N_13483);
and U15367 (N_15367,N_10337,N_12046);
or U15368 (N_15368,N_12109,N_13981);
nor U15369 (N_15369,N_12530,N_13446);
and U15370 (N_15370,N_12431,N_14188);
nor U15371 (N_15371,N_10695,N_13826);
or U15372 (N_15372,N_10645,N_12804);
and U15373 (N_15373,N_10398,N_12145);
nor U15374 (N_15374,N_10378,N_11875);
or U15375 (N_15375,N_14797,N_13077);
or U15376 (N_15376,N_13014,N_14041);
or U15377 (N_15377,N_13695,N_13109);
and U15378 (N_15378,N_11691,N_11215);
xnor U15379 (N_15379,N_10078,N_14528);
or U15380 (N_15380,N_11132,N_13799);
nand U15381 (N_15381,N_12338,N_11515);
or U15382 (N_15382,N_13929,N_14618);
nand U15383 (N_15383,N_13655,N_11505);
or U15384 (N_15384,N_10697,N_14358);
and U15385 (N_15385,N_11817,N_13445);
or U15386 (N_15386,N_14395,N_10722);
nor U15387 (N_15387,N_12027,N_12026);
and U15388 (N_15388,N_12161,N_14462);
nor U15389 (N_15389,N_10334,N_11928);
nand U15390 (N_15390,N_13950,N_11914);
or U15391 (N_15391,N_14519,N_14052);
or U15392 (N_15392,N_12089,N_14135);
and U15393 (N_15393,N_12902,N_13797);
and U15394 (N_15394,N_10900,N_14165);
and U15395 (N_15395,N_13163,N_14259);
or U15396 (N_15396,N_10077,N_13162);
and U15397 (N_15397,N_12015,N_12346);
or U15398 (N_15398,N_11573,N_13489);
or U15399 (N_15399,N_13698,N_10501);
nand U15400 (N_15400,N_14492,N_13944);
and U15401 (N_15401,N_10480,N_10423);
and U15402 (N_15402,N_11504,N_14207);
nor U15403 (N_15403,N_12811,N_11780);
xnor U15404 (N_15404,N_11883,N_14578);
nor U15405 (N_15405,N_14281,N_14924);
nand U15406 (N_15406,N_13339,N_10821);
or U15407 (N_15407,N_11734,N_13423);
or U15408 (N_15408,N_12531,N_11869);
and U15409 (N_15409,N_11809,N_11155);
nor U15410 (N_15410,N_11921,N_12425);
nor U15411 (N_15411,N_13824,N_14594);
or U15412 (N_15412,N_12127,N_10184);
nor U15413 (N_15413,N_14595,N_14609);
nor U15414 (N_15414,N_10236,N_10110);
and U15415 (N_15415,N_10917,N_14344);
and U15416 (N_15416,N_14941,N_14452);
and U15417 (N_15417,N_13743,N_11803);
or U15418 (N_15418,N_11710,N_11086);
nor U15419 (N_15419,N_13609,N_11585);
and U15420 (N_15420,N_12742,N_11114);
and U15421 (N_15421,N_13236,N_14963);
nand U15422 (N_15422,N_14218,N_10938);
or U15423 (N_15423,N_12011,N_12410);
and U15424 (N_15424,N_13515,N_13566);
or U15425 (N_15425,N_11876,N_14743);
nor U15426 (N_15426,N_14780,N_14834);
and U15427 (N_15427,N_11689,N_14133);
nor U15428 (N_15428,N_12847,N_11716);
nand U15429 (N_15429,N_11767,N_14542);
nor U15430 (N_15430,N_11683,N_11640);
xor U15431 (N_15431,N_12653,N_10791);
or U15432 (N_15432,N_13575,N_14014);
or U15433 (N_15433,N_12677,N_11701);
nand U15434 (N_15434,N_11626,N_12336);
and U15435 (N_15435,N_14355,N_11602);
or U15436 (N_15436,N_10750,N_11623);
nor U15437 (N_15437,N_12457,N_13554);
nand U15438 (N_15438,N_11906,N_10410);
and U15439 (N_15439,N_13939,N_12599);
or U15440 (N_15440,N_14332,N_13518);
nand U15441 (N_15441,N_10865,N_13718);
and U15442 (N_15442,N_13638,N_12125);
nand U15443 (N_15443,N_12463,N_10540);
or U15444 (N_15444,N_11598,N_14196);
nand U15445 (N_15445,N_12192,N_10338);
nor U15446 (N_15446,N_14664,N_13282);
or U15447 (N_15447,N_10673,N_12318);
and U15448 (N_15448,N_13120,N_14894);
or U15449 (N_15449,N_10320,N_13620);
or U15450 (N_15450,N_14808,N_10118);
nor U15451 (N_15451,N_12317,N_11990);
or U15452 (N_15452,N_10262,N_14778);
or U15453 (N_15453,N_11708,N_14319);
and U15454 (N_15454,N_13568,N_11338);
and U15455 (N_15455,N_14577,N_13795);
or U15456 (N_15456,N_11549,N_14150);
nor U15457 (N_15457,N_13422,N_11347);
nor U15458 (N_15458,N_11110,N_12759);
or U15459 (N_15459,N_10144,N_11507);
nor U15460 (N_15460,N_10374,N_14456);
or U15461 (N_15461,N_14393,N_11103);
or U15462 (N_15462,N_10926,N_11980);
or U15463 (N_15463,N_13664,N_11056);
and U15464 (N_15464,N_13375,N_10840);
and U15465 (N_15465,N_10627,N_10969);
nor U15466 (N_15466,N_12356,N_11438);
nor U15467 (N_15467,N_11199,N_14107);
and U15468 (N_15468,N_11957,N_10350);
or U15469 (N_15469,N_14637,N_11934);
nand U15470 (N_15470,N_12112,N_12100);
and U15471 (N_15471,N_14176,N_12922);
or U15472 (N_15472,N_13984,N_10644);
nand U15473 (N_15473,N_14032,N_14350);
and U15474 (N_15474,N_12308,N_13595);
nor U15475 (N_15475,N_10343,N_10027);
nand U15476 (N_15476,N_13866,N_13288);
or U15477 (N_15477,N_11537,N_10556);
and U15478 (N_15478,N_11181,N_12736);
or U15479 (N_15479,N_14631,N_10083);
nor U15480 (N_15480,N_13388,N_13475);
and U15481 (N_15481,N_13486,N_10314);
and U15482 (N_15482,N_14366,N_11704);
and U15483 (N_15483,N_10613,N_13226);
and U15484 (N_15484,N_10594,N_10584);
nand U15485 (N_15485,N_12576,N_10347);
nor U15486 (N_15486,N_12462,N_12810);
nor U15487 (N_15487,N_14476,N_11909);
or U15488 (N_15488,N_11372,N_13840);
and U15489 (N_15489,N_11948,N_10758);
or U15490 (N_15490,N_10510,N_13644);
and U15491 (N_15491,N_13853,N_12840);
or U15492 (N_15492,N_13395,N_11131);
and U15493 (N_15493,N_13059,N_12645);
nand U15494 (N_15494,N_11559,N_12879);
nor U15495 (N_15495,N_12365,N_10838);
or U15496 (N_15496,N_14028,N_12434);
nand U15497 (N_15497,N_11104,N_14751);
and U15498 (N_15498,N_10402,N_10564);
nand U15499 (N_15499,N_14912,N_11588);
or U15500 (N_15500,N_14776,N_13286);
xnor U15501 (N_15501,N_13733,N_13103);
nor U15502 (N_15502,N_13882,N_13549);
or U15503 (N_15503,N_11748,N_14655);
nand U15504 (N_15504,N_14900,N_14385);
nor U15505 (N_15505,N_14848,N_14437);
nor U15506 (N_15506,N_14254,N_10891);
nor U15507 (N_15507,N_14250,N_13485);
xor U15508 (N_15508,N_13765,N_11618);
nor U15509 (N_15509,N_12858,N_12248);
or U15510 (N_15510,N_12086,N_11860);
nor U15511 (N_15511,N_10342,N_13502);
or U15512 (N_15512,N_14791,N_10871);
nand U15513 (N_15513,N_12581,N_11898);
nand U15514 (N_15514,N_13542,N_14423);
nor U15515 (N_15515,N_10736,N_11321);
nor U15516 (N_15516,N_10291,N_11753);
and U15517 (N_15517,N_10062,N_10619);
and U15518 (N_15518,N_14347,N_13890);
nand U15519 (N_15519,N_14878,N_14861);
nand U15520 (N_15520,N_12299,N_12723);
and U15521 (N_15521,N_13651,N_14605);
nor U15522 (N_15522,N_11482,N_14060);
nand U15523 (N_15523,N_14340,N_10080);
nor U15524 (N_15524,N_11077,N_11415);
nand U15525 (N_15525,N_12122,N_10641);
or U15526 (N_15526,N_13173,N_10328);
and U15527 (N_15527,N_11028,N_14002);
and U15528 (N_15528,N_13574,N_12630);
nand U15529 (N_15529,N_14919,N_11523);
and U15530 (N_15530,N_14719,N_11269);
and U15531 (N_15531,N_10068,N_12049);
or U15532 (N_15532,N_13699,N_12994);
and U15533 (N_15533,N_12515,N_11905);
or U15534 (N_15534,N_13350,N_14762);
and U15535 (N_15535,N_10230,N_12794);
or U15536 (N_15536,N_10803,N_12012);
or U15537 (N_15537,N_12174,N_11805);
nor U15538 (N_15538,N_13827,N_12313);
and U15539 (N_15539,N_11839,N_10719);
nand U15540 (N_15540,N_11768,N_14233);
nor U15541 (N_15541,N_10226,N_11290);
nor U15542 (N_15542,N_10346,N_10639);
nand U15543 (N_15543,N_13108,N_12119);
nand U15544 (N_15544,N_10839,N_14470);
nor U15545 (N_15545,N_14986,N_13078);
or U15546 (N_15546,N_13573,N_13815);
nand U15547 (N_15547,N_10088,N_11988);
or U15548 (N_15548,N_12798,N_14104);
xor U15549 (N_15549,N_13803,N_14050);
or U15550 (N_15550,N_12904,N_11459);
nor U15551 (N_15551,N_14228,N_11154);
nor U15552 (N_15552,N_11057,N_10856);
nor U15553 (N_15553,N_14200,N_10174);
nand U15554 (N_15554,N_12572,N_14563);
or U15555 (N_15555,N_12623,N_12708);
nor U15556 (N_15556,N_10008,N_12148);
or U15557 (N_15557,N_14914,N_13748);
and U15558 (N_15558,N_14703,N_14112);
and U15559 (N_15559,N_10676,N_14374);
or U15560 (N_15560,N_10825,N_13180);
or U15561 (N_15561,N_11072,N_12584);
and U15562 (N_15562,N_14236,N_14515);
or U15563 (N_15563,N_11901,N_10058);
and U15564 (N_15564,N_10596,N_12595);
or U15565 (N_15565,N_12631,N_12837);
or U15566 (N_15566,N_10935,N_11311);
nand U15567 (N_15567,N_11677,N_12939);
and U15568 (N_15568,N_11923,N_14480);
and U15569 (N_15569,N_10588,N_13828);
nand U15570 (N_15570,N_10470,N_14603);
nand U15571 (N_15571,N_12250,N_14708);
or U15572 (N_15572,N_13248,N_12781);
nor U15573 (N_15573,N_12822,N_13262);
nor U15574 (N_15574,N_14469,N_11463);
or U15575 (N_15575,N_11951,N_14387);
and U15576 (N_15576,N_12628,N_10961);
or U15577 (N_15577,N_14969,N_11208);
nand U15578 (N_15578,N_13994,N_13154);
and U15579 (N_15579,N_10586,N_10792);
and U15580 (N_15580,N_10524,N_14521);
and U15581 (N_15581,N_10987,N_11700);
xor U15582 (N_15582,N_10635,N_12883);
nor U15583 (N_15583,N_10267,N_13175);
nand U15584 (N_15584,N_13597,N_14430);
nand U15585 (N_15585,N_12080,N_12083);
or U15586 (N_15586,N_13744,N_14636);
nor U15587 (N_15587,N_14895,N_10014);
or U15588 (N_15588,N_13053,N_14006);
and U15589 (N_15589,N_11418,N_14551);
nand U15590 (N_15590,N_14294,N_12404);
or U15591 (N_15591,N_12056,N_10910);
nor U15592 (N_15592,N_10904,N_14359);
nand U15593 (N_15593,N_10237,N_14771);
nand U15594 (N_15594,N_14865,N_14169);
nand U15595 (N_15595,N_14835,N_12413);
or U15596 (N_15596,N_14592,N_10187);
nor U15597 (N_15597,N_13354,N_10364);
or U15598 (N_15598,N_10772,N_12268);
or U15599 (N_15599,N_14604,N_11384);
and U15600 (N_15600,N_14418,N_13833);
or U15601 (N_15601,N_13192,N_11836);
nand U15602 (N_15602,N_14428,N_14483);
nor U15603 (N_15603,N_11764,N_14113);
nand U15604 (N_15604,N_14702,N_11603);
or U15605 (N_15605,N_13908,N_11245);
nor U15606 (N_15606,N_10680,N_14091);
nand U15607 (N_15607,N_10138,N_12423);
nor U15608 (N_15608,N_13905,N_11872);
and U15609 (N_15609,N_14802,N_10503);
nand U15610 (N_15610,N_10181,N_10495);
nand U15611 (N_15611,N_11107,N_12539);
nand U15612 (N_15612,N_10994,N_13844);
and U15613 (N_15613,N_14773,N_10667);
or U15614 (N_15614,N_11000,N_12441);
or U15615 (N_15615,N_11797,N_12121);
and U15616 (N_15616,N_11152,N_11074);
and U15617 (N_15617,N_14499,N_11191);
and U15618 (N_15618,N_13032,N_11143);
or U15619 (N_15619,N_12619,N_12524);
or U15620 (N_15620,N_10567,N_13145);
nand U15621 (N_15621,N_12971,N_11271);
nand U15622 (N_15622,N_12224,N_10289);
or U15623 (N_15623,N_12787,N_12603);
and U15624 (N_15624,N_13716,N_10927);
or U15625 (N_15625,N_11941,N_12553);
and U15626 (N_15626,N_11133,N_11724);
or U15627 (N_15627,N_10571,N_12375);
and U15628 (N_15628,N_11166,N_12399);
or U15629 (N_15629,N_14217,N_11031);
and U15630 (N_15630,N_13730,N_11728);
or U15631 (N_15631,N_10163,N_12165);
or U15632 (N_15632,N_14381,N_10653);
nand U15633 (N_15633,N_13740,N_13207);
nor U15634 (N_15634,N_13348,N_14921);
nor U15635 (N_15635,N_13734,N_12836);
and U15636 (N_15636,N_13416,N_10276);
or U15637 (N_15637,N_11830,N_11851);
or U15638 (N_15638,N_14275,N_12867);
or U15639 (N_15639,N_11642,N_11744);
xor U15640 (N_15640,N_11476,N_11657);
or U15641 (N_15641,N_11495,N_12214);
or U15642 (N_15642,N_14717,N_11410);
and U15643 (N_15643,N_12153,N_10247);
and U15644 (N_15644,N_13322,N_14942);
nand U15645 (N_15645,N_12055,N_13168);
nor U15646 (N_15646,N_13683,N_13520);
nor U15647 (N_15647,N_10955,N_10401);
and U15648 (N_15648,N_14386,N_13760);
nand U15649 (N_15649,N_11182,N_10894);
nor U15650 (N_15650,N_12953,N_12791);
and U15651 (N_15651,N_10753,N_14211);
and U15652 (N_15652,N_13111,N_13669);
nor U15653 (N_15653,N_11637,N_12372);
or U15654 (N_15654,N_13046,N_14553);
and U15655 (N_15655,N_12906,N_10972);
nor U15656 (N_15656,N_10545,N_14417);
or U15657 (N_15657,N_11319,N_10356);
nand U15658 (N_15658,N_14260,N_12962);
and U15659 (N_15659,N_11524,N_14511);
nor U15660 (N_15660,N_10998,N_14568);
nand U15661 (N_15661,N_14361,N_10021);
or U15662 (N_15662,N_14612,N_10220);
and U15663 (N_15663,N_11960,N_10205);
nand U15664 (N_15664,N_13247,N_13612);
or U15665 (N_15665,N_13965,N_14191);
and U15666 (N_15666,N_13137,N_12014);
nand U15667 (N_15667,N_14994,N_10446);
nor U15668 (N_15668,N_12382,N_12226);
nand U15669 (N_15669,N_14392,N_12216);
nand U15670 (N_15670,N_12609,N_14266);
or U15671 (N_15671,N_10271,N_10906);
nand U15672 (N_15672,N_10660,N_12829);
or U15673 (N_15673,N_11473,N_12892);
and U15674 (N_15674,N_13146,N_12183);
nor U15675 (N_15675,N_12557,N_10156);
and U15676 (N_15676,N_10723,N_12918);
and U15677 (N_15677,N_12147,N_12197);
or U15678 (N_15678,N_14342,N_13593);
or U15679 (N_15679,N_12439,N_14937);
nor U15680 (N_15680,N_10143,N_11984);
nor U15681 (N_15681,N_10622,N_11233);
nand U15682 (N_15682,N_12010,N_10546);
nand U15683 (N_15683,N_13270,N_14201);
nor U15684 (N_15684,N_12944,N_14035);
nor U15685 (N_15685,N_10578,N_14027);
nand U15686 (N_15686,N_12970,N_11855);
or U15687 (N_15687,N_11513,N_11609);
and U15688 (N_15688,N_10028,N_11093);
nor U15689 (N_15689,N_11160,N_14313);
or U15690 (N_15690,N_14125,N_10535);
nor U15691 (N_15691,N_12280,N_11517);
nor U15692 (N_15692,N_10413,N_13510);
or U15693 (N_15693,N_14582,N_10046);
and U15694 (N_15694,N_13711,N_10295);
and U15695 (N_15695,N_11801,N_10489);
nand U15696 (N_15696,N_10379,N_10665);
nor U15697 (N_15697,N_13556,N_13852);
nor U15698 (N_15698,N_14532,N_13501);
or U15699 (N_15699,N_12233,N_13383);
nor U15700 (N_15700,N_10453,N_11571);
nand U15701 (N_15701,N_12800,N_13507);
nor U15702 (N_15702,N_14042,N_12866);
or U15703 (N_15703,N_14038,N_12685);
and U15704 (N_15704,N_13110,N_13203);
xor U15705 (N_15705,N_14182,N_11264);
nand U15706 (N_15706,N_10211,N_14016);
xor U15707 (N_15707,N_11674,N_13687);
or U15708 (N_15708,N_13449,N_12078);
xor U15709 (N_15709,N_13151,N_12417);
nand U15710 (N_15710,N_13285,N_12437);
and U15711 (N_15711,N_13932,N_12485);
nor U15712 (N_15712,N_12737,N_14574);
or U15713 (N_15713,N_11562,N_10203);
or U15714 (N_15714,N_11249,N_14497);
nand U15715 (N_15715,N_12734,N_11493);
nand U15716 (N_15716,N_11841,N_11548);
nand U15717 (N_15717,N_11081,N_14257);
nor U15718 (N_15718,N_10189,N_10529);
nand U15719 (N_15719,N_14993,N_10824);
or U15720 (N_15720,N_10843,N_14887);
nor U15721 (N_15721,N_13953,N_13062);
and U15722 (N_15722,N_14882,N_13199);
xnor U15723 (N_15723,N_13377,N_12465);
nor U15724 (N_15724,N_10387,N_10620);
or U15725 (N_15725,N_13017,N_10048);
and U15726 (N_15726,N_11854,N_11947);
nand U15727 (N_15727,N_14047,N_10377);
or U15728 (N_15728,N_10282,N_10278);
nor U15729 (N_15729,N_13894,N_11406);
or U15730 (N_15730,N_10573,N_13693);
nor U15731 (N_15731,N_13941,N_14600);
nor U15732 (N_15732,N_13068,N_10781);
and U15733 (N_15733,N_10971,N_12260);
or U15734 (N_15734,N_11619,N_12293);
and U15735 (N_15735,N_10497,N_12409);
nand U15736 (N_15736,N_14296,N_13764);
nor U15737 (N_15737,N_11146,N_11006);
and U15738 (N_15738,N_10207,N_14283);
nand U15739 (N_15739,N_10254,N_14615);
nor U15740 (N_15740,N_10921,N_12543);
nor U15741 (N_15741,N_14413,N_11766);
nand U15742 (N_15742,N_10455,N_13424);
nor U15743 (N_15743,N_10092,N_14429);
and U15744 (N_15744,N_10430,N_14864);
or U15745 (N_15745,N_10188,N_11195);
or U15746 (N_15746,N_14096,N_12605);
nand U15747 (N_15747,N_11039,N_14086);
nand U15748 (N_15748,N_13080,N_12777);
or U15749 (N_15749,N_14909,N_14970);
nand U15750 (N_15750,N_12458,N_12138);
nor U15751 (N_15751,N_13697,N_13267);
nor U15752 (N_15752,N_10864,N_11823);
nor U15753 (N_15753,N_13737,N_13583);
xnor U15754 (N_15754,N_13394,N_11397);
xor U15755 (N_15755,N_11762,N_12919);
nor U15756 (N_15756,N_10162,N_14646);
or U15757 (N_15757,N_13235,N_14632);
xor U15758 (N_15758,N_12520,N_10576);
nor U15759 (N_15759,N_12091,N_12384);
nand U15760 (N_15760,N_10416,N_13224);
and U15761 (N_15761,N_13681,N_11520);
or U15762 (N_15762,N_10035,N_13172);
nand U15763 (N_15763,N_12230,N_10965);
or U15764 (N_15764,N_13147,N_12249);
or U15765 (N_15765,N_12881,N_14763);
nor U15766 (N_15766,N_12980,N_13921);
or U15767 (N_15767,N_14870,N_10176);
and U15768 (N_15768,N_13793,N_12664);
nand U15769 (N_15769,N_14723,N_10117);
and U15770 (N_15770,N_10294,N_12222);
nor U15771 (N_15771,N_10333,N_10040);
and U15772 (N_15772,N_12622,N_10600);
nor U15773 (N_15773,N_13391,N_11730);
nor U15774 (N_15774,N_14121,N_12304);
nor U15775 (N_15775,N_11769,N_14010);
or U15776 (N_15776,N_13269,N_12852);
and U15777 (N_15777,N_12263,N_13159);
and U15778 (N_15778,N_12287,N_11130);
and U15779 (N_15779,N_10308,N_12269);
nor U15780 (N_15780,N_12886,N_10125);
nor U15781 (N_15781,N_10966,N_11178);
xnor U15782 (N_15782,N_12130,N_13128);
or U15783 (N_15783,N_11198,N_13297);
xor U15784 (N_15784,N_11064,N_14836);
and U15785 (N_15785,N_10219,N_14000);
nand U15786 (N_15786,N_13088,N_11794);
or U15787 (N_15787,N_10777,N_14714);
nor U15788 (N_15788,N_14030,N_13899);
and U15789 (N_15789,N_13786,N_10448);
nor U15790 (N_15790,N_13634,N_10905);
or U15791 (N_15791,N_14700,N_12422);
or U15792 (N_15792,N_13841,N_11904);
or U15793 (N_15793,N_11979,N_12255);
nand U15794 (N_15794,N_11614,N_11758);
nand U15795 (N_15795,N_10984,N_14216);
nand U15796 (N_15796,N_13382,N_14628);
nor U15797 (N_15797,N_11201,N_13968);
nand U15798 (N_15798,N_11422,N_11232);
nor U15799 (N_15799,N_10302,N_13371);
and U15800 (N_15800,N_12917,N_11586);
nand U15801 (N_15801,N_14977,N_14948);
or U15802 (N_15802,N_12757,N_12783);
nor U15803 (N_15803,N_13243,N_10095);
nor U15804 (N_15804,N_11453,N_11320);
or U15805 (N_15805,N_11705,N_10922);
nor U15806 (N_15806,N_10543,N_13249);
or U15807 (N_15807,N_14815,N_12120);
nor U15808 (N_15808,N_11236,N_14187);
or U15809 (N_15809,N_13749,N_13961);
and U15810 (N_15810,N_14545,N_10467);
nor U15811 (N_15811,N_11027,N_14644);
or U15812 (N_15812,N_11334,N_10826);
nor U15813 (N_15813,N_11485,N_10201);
nor U15814 (N_15814,N_13525,N_14031);
nand U15815 (N_15815,N_11051,N_12374);
nand U15816 (N_15816,N_12393,N_10030);
nor U15817 (N_15817,N_11228,N_14811);
nor U15818 (N_15818,N_11352,N_12899);
nand U15819 (N_15819,N_10708,N_13004);
nor U15820 (N_15820,N_11658,N_10845);
nor U15821 (N_15821,N_13526,N_11779);
nor U15822 (N_15822,N_10299,N_11862);
and U15823 (N_15823,N_13972,N_11880);
nand U15824 (N_15824,N_13552,N_14896);
nor U15825 (N_15825,N_11725,N_11277);
nor U15826 (N_15826,N_11394,N_14066);
nand U15827 (N_15827,N_13205,N_12476);
xor U15828 (N_15828,N_11392,N_13346);
and U15829 (N_15829,N_12185,N_12814);
and U15830 (N_15830,N_11638,N_14320);
nor U15831 (N_15831,N_13411,N_12072);
and U15832 (N_15832,N_10394,N_12552);
or U15833 (N_15833,N_14627,N_10281);
and U15834 (N_15834,N_12460,N_14481);
or U15835 (N_15835,N_14713,N_12956);
nor U15836 (N_15836,N_11484,N_10623);
or U15837 (N_15837,N_12172,N_12009);
nor U15838 (N_15838,N_11522,N_12556);
nor U15839 (N_15839,N_11240,N_14807);
or U15840 (N_15840,N_12135,N_11634);
or U15841 (N_15841,N_14853,N_13843);
or U15842 (N_15842,N_12217,N_12265);
xnor U15843 (N_15843,N_12839,N_13812);
nor U15844 (N_15844,N_14087,N_14130);
nand U15845 (N_15845,N_13466,N_11936);
nand U15846 (N_15846,N_11629,N_10547);
or U15847 (N_15847,N_14675,N_12339);
or U15848 (N_15848,N_13060,N_13768);
and U15849 (N_15849,N_14173,N_11365);
nand U15850 (N_15850,N_10956,N_10973);
and U15851 (N_15851,N_11993,N_14990);
and U15852 (N_15852,N_13035,N_10899);
or U15853 (N_15853,N_14422,N_14580);
nand U15854 (N_15854,N_11225,N_12596);
nor U15855 (N_15855,N_12528,N_10813);
and U15856 (N_15856,N_12636,N_13468);
nor U15857 (N_15857,N_12935,N_10057);
nand U15858 (N_15858,N_13327,N_11816);
nor U15859 (N_15859,N_11832,N_12272);
nor U15860 (N_15860,N_10098,N_13245);
or U15861 (N_15861,N_14548,N_11920);
or U15862 (N_15862,N_10851,N_13185);
nor U15863 (N_15863,N_11238,N_10517);
nand U15864 (N_15864,N_13780,N_12411);
or U15865 (N_15865,N_13091,N_13521);
nand U15866 (N_15866,N_14705,N_12202);
xnor U15867 (N_15867,N_10787,N_12518);
and U15868 (N_15868,N_14596,N_14071);
nand U15869 (N_15869,N_11572,N_13126);
or U15870 (N_15870,N_10642,N_13306);
and U15871 (N_15871,N_13727,N_11519);
and U15872 (N_15872,N_11733,N_11676);
nand U15873 (N_15873,N_10698,N_12491);
xnor U15874 (N_15874,N_13598,N_11969);
nor U15875 (N_15875,N_12704,N_11635);
and U15876 (N_15876,N_10989,N_11447);
or U15877 (N_15877,N_10762,N_12395);
nor U15878 (N_15878,N_13330,N_11699);
or U15879 (N_15879,N_10160,N_14454);
and U15880 (N_15880,N_12252,N_12137);
and U15881 (N_15881,N_13956,N_10233);
or U15882 (N_15882,N_13316,N_13258);
nand U15883 (N_15883,N_10801,N_11009);
nand U15884 (N_15884,N_11690,N_12976);
or U15885 (N_15885,N_12908,N_12701);
nor U15886 (N_15886,N_11193,N_11679);
or U15887 (N_15887,N_12663,N_14728);
nor U15888 (N_15888,N_13970,N_13934);
or U15889 (N_15889,N_10449,N_14274);
or U15890 (N_15890,N_11697,N_11136);
nor U15891 (N_15891,N_13719,N_12288);
nand U15892 (N_15892,N_14265,N_10549);
and U15893 (N_15893,N_14754,N_11443);
and U15894 (N_15894,N_10669,N_10923);
and U15895 (N_15895,N_10321,N_10312);
nand U15896 (N_15896,N_12570,N_10404);
and U15897 (N_15897,N_12824,N_13639);
nand U15898 (N_15898,N_14189,N_11095);
nor U15899 (N_15899,N_13775,N_12464);
nor U15900 (N_15900,N_11983,N_14144);
or U15901 (N_15901,N_10784,N_13149);
or U15902 (N_15902,N_10844,N_12646);
and U15903 (N_15903,N_12473,N_13469);
or U15904 (N_15904,N_12211,N_12076);
nand U15905 (N_15905,N_10970,N_12949);
or U15906 (N_15906,N_14825,N_11437);
nor U15907 (N_15907,N_14273,N_11992);
nand U15908 (N_15908,N_13911,N_13792);
nand U15909 (N_15909,N_11852,N_11012);
nor U15910 (N_15910,N_12635,N_14901);
nor U15911 (N_15911,N_10131,N_11270);
nand U15912 (N_15912,N_13945,N_14379);
and U15913 (N_15913,N_10804,N_14918);
or U15914 (N_15914,N_10816,N_10332);
nand U15915 (N_15915,N_14287,N_11080);
nor U15916 (N_15916,N_11660,N_11021);
or U15917 (N_15917,N_12891,N_10552);
or U15918 (N_15918,N_11655,N_10688);
nor U15919 (N_15919,N_13488,N_12930);
nand U15920 (N_15920,N_12166,N_12102);
nand U15921 (N_15921,N_12534,N_10898);
and U15922 (N_15922,N_12845,N_12237);
or U15923 (N_15923,N_13626,N_12731);
nor U15924 (N_15924,N_11294,N_12732);
and U15925 (N_15925,N_10018,N_13209);
xnor U15926 (N_15926,N_11366,N_12295);
nand U15927 (N_15927,N_11120,N_12392);
nand U15928 (N_15928,N_12565,N_14750);
or U15929 (N_15929,N_13041,N_11508);
and U15930 (N_15930,N_10096,N_12651);
xnor U15931 (N_15931,N_14258,N_10569);
nand U15932 (N_15932,N_13239,N_11255);
nor U15933 (N_15933,N_10548,N_10488);
nand U15934 (N_15934,N_12673,N_14725);
and U15935 (N_15935,N_13946,N_12484);
nor U15936 (N_15936,N_10629,N_12767);
nand U15937 (N_15937,N_13089,N_11149);
nand U15938 (N_15938,N_13504,N_11032);
nor U15939 (N_15939,N_14862,N_12979);
and U15940 (N_15940,N_14999,N_14952);
and U15941 (N_15941,N_13543,N_13266);
nor U15942 (N_15942,N_10855,N_13720);
nor U15943 (N_15943,N_12041,N_12998);
nand U15944 (N_15944,N_14640,N_12752);
and U15945 (N_15945,N_14067,N_14830);
and U15946 (N_15946,N_12090,N_11681);
or U15947 (N_15947,N_12361,N_13951);
or U15948 (N_15948,N_11075,N_11822);
nor U15949 (N_15949,N_10595,N_14523);
nand U15950 (N_15950,N_13897,N_11567);
nand U15951 (N_15951,N_11721,N_10175);
or U15952 (N_15952,N_11260,N_14522);
and U15953 (N_15953,N_11910,N_13332);
or U15954 (N_15954,N_14786,N_13559);
nor U15955 (N_15955,N_14661,N_12347);
nor U15956 (N_15956,N_10744,N_13808);
or U15957 (N_15957,N_14916,N_14153);
or U15958 (N_15958,N_11838,N_11342);
nor U15959 (N_15959,N_13201,N_14989);
and U15960 (N_15960,N_12857,N_14650);
nand U15961 (N_15961,N_10786,N_14813);
nor U15962 (N_15962,N_10919,N_12267);
nor U15963 (N_15963,N_14752,N_14024);
nand U15964 (N_15964,N_14822,N_14938);
or U15965 (N_15965,N_11632,N_14816);
or U15966 (N_15966,N_11848,N_11185);
or U15967 (N_15967,N_11204,N_10053);
nand U15968 (N_15968,N_11005,N_14285);
nor U15969 (N_15969,N_11525,N_12496);
nor U15970 (N_15970,N_12986,N_12788);
nor U15971 (N_15971,N_13809,N_11917);
and U15972 (N_15972,N_11060,N_10403);
nor U15973 (N_15973,N_10605,N_10243);
nand U15974 (N_15974,N_11183,N_11395);
or U15975 (N_15975,N_10002,N_13958);
or U15976 (N_15976,N_13420,N_10944);
and U15977 (N_15977,N_10106,N_12612);
nand U15978 (N_15978,N_12494,N_14443);
and U15979 (N_15979,N_13721,N_12403);
nand U15980 (N_15980,N_14688,N_12025);
nand U15981 (N_15981,N_10022,N_14240);
nor U15982 (N_15982,N_14263,N_13428);
nor U15983 (N_15983,N_14774,N_12801);
or U15984 (N_15984,N_10790,N_14727);
and U15985 (N_15985,N_14249,N_11036);
nor U15986 (N_15986,N_12111,N_14742);
or U15987 (N_15987,N_14855,N_11345);
and U15988 (N_15988,N_11799,N_13892);
or U15989 (N_15989,N_14524,N_12746);
nor U15990 (N_15990,N_13701,N_14787);
and U15991 (N_15991,N_10531,N_14685);
nor U15992 (N_15992,N_13869,N_14906);
or U15993 (N_15993,N_10611,N_10693);
or U15994 (N_15994,N_13616,N_10760);
nand U15995 (N_15995,N_14070,N_10913);
nor U15996 (N_15996,N_14943,N_10756);
nor U15997 (N_15997,N_14767,N_13123);
nand U15998 (N_15998,N_12985,N_14102);
nor U15999 (N_15999,N_12597,N_14526);
nor U16000 (N_16000,N_12818,N_13202);
nand U16001 (N_16001,N_14684,N_11020);
nor U16002 (N_16002,N_11386,N_10924);
or U16003 (N_16003,N_10269,N_12975);
and U16004 (N_16004,N_10086,N_10127);
and U16005 (N_16005,N_14037,N_13691);
nand U16006 (N_16006,N_14389,N_13997);
and U16007 (N_16007,N_13031,N_13670);
nor U16008 (N_16008,N_12616,N_12032);
or U16009 (N_16009,N_14926,N_10390);
or U16010 (N_16010,N_13954,N_13084);
nand U16011 (N_16011,N_13947,N_12036);
nand U16012 (N_16012,N_11899,N_14394);
nand U16013 (N_16013,N_12349,N_13653);
or U16014 (N_16014,N_14648,N_14338);
nand U16015 (N_16015,N_12696,N_11968);
nor U16016 (N_16016,N_10953,N_10134);
and U16017 (N_16017,N_12163,N_12706);
xnor U16018 (N_16018,N_13102,N_10266);
or U16019 (N_16019,N_14368,N_12957);
nor U16020 (N_16020,N_12844,N_10209);
nand U16021 (N_16021,N_13006,N_14814);
and U16022 (N_16022,N_14686,N_13105);
nand U16023 (N_16023,N_11038,N_13113);
nor U16024 (N_16024,N_14414,N_12469);
and U16025 (N_16025,N_11723,N_11084);
or U16026 (N_16026,N_12194,N_14980);
and U16027 (N_16027,N_13964,N_12378);
nor U16028 (N_16028,N_13417,N_10583);
nand U16029 (N_16029,N_10560,N_13925);
or U16030 (N_16030,N_11726,N_10878);
nor U16031 (N_16031,N_12198,N_13660);
or U16032 (N_16032,N_14820,N_14055);
nand U16033 (N_16033,N_14772,N_13259);
and U16034 (N_16034,N_10604,N_12546);
nand U16035 (N_16035,N_14897,N_13825);
nand U16036 (N_16036,N_14243,N_14556);
and U16037 (N_16037,N_14450,N_12535);
nand U16038 (N_16038,N_14181,N_11371);
or U16039 (N_16039,N_12510,N_14369);
or U16040 (N_16040,N_12062,N_11307);
and U16041 (N_16041,N_13454,N_12023);
and U16042 (N_16042,N_14880,N_13550);
and U16043 (N_16043,N_13930,N_10204);
or U16044 (N_16044,N_11844,N_12066);
nand U16045 (N_16045,N_11412,N_10432);
nand U16046 (N_16046,N_11709,N_12499);
xnor U16047 (N_16047,N_10523,N_13642);
nand U16048 (N_16048,N_10749,N_11878);
nor U16049 (N_16049,N_11170,N_12808);
xor U16050 (N_16050,N_13229,N_14487);
and U16051 (N_16051,N_12178,N_12244);
or U16052 (N_16052,N_10768,N_10383);
nor U16053 (N_16053,N_14082,N_14136);
and U16054 (N_16054,N_13051,N_11584);
nand U16055 (N_16055,N_13025,N_13334);
and U16056 (N_16056,N_14406,N_14325);
or U16057 (N_16057,N_14920,N_13986);
nand U16058 (N_16058,N_12816,N_14619);
or U16059 (N_16059,N_13907,N_10229);
nand U16060 (N_16060,N_14376,N_11943);
nand U16061 (N_16061,N_13499,N_14509);
nand U16062 (N_16062,N_11886,N_14518);
and U16063 (N_16063,N_14120,N_12657);
xnor U16064 (N_16064,N_11868,N_11694);
or U16065 (N_16065,N_12554,N_11407);
and U16066 (N_16066,N_13769,N_13959);
and U16067 (N_16067,N_10853,N_14534);
nand U16068 (N_16068,N_10304,N_14681);
nand U16069 (N_16069,N_14740,N_10706);
or U16070 (N_16070,N_12549,N_11134);
and U16071 (N_16071,N_11002,N_13884);
nand U16072 (N_16072,N_11995,N_12561);
and U16073 (N_16073,N_11224,N_11617);
nand U16074 (N_16074,N_10165,N_14415);
and U16075 (N_16075,N_11915,N_13379);
or U16076 (N_16076,N_12059,N_10985);
xnor U16077 (N_16077,N_12606,N_10382);
nand U16078 (N_16078,N_14800,N_10036);
or U16079 (N_16079,N_14512,N_14833);
xor U16080 (N_16080,N_12503,N_10457);
or U16081 (N_16081,N_10662,N_14575);
nand U16082 (N_16082,N_14147,N_12948);
and U16083 (N_16083,N_14701,N_10420);
and U16084 (N_16084,N_14745,N_11669);
and U16085 (N_16085,N_12123,N_11806);
or U16086 (N_16086,N_13529,N_12160);
or U16087 (N_16087,N_13661,N_10658);
and U16088 (N_16088,N_11579,N_14852);
nand U16089 (N_16089,N_11754,N_12719);
and U16090 (N_16090,N_12920,N_13242);
or U16091 (N_16091,N_12903,N_12815);
nor U16092 (N_16092,N_11141,N_12415);
nand U16093 (N_16093,N_12914,N_10481);
and U16094 (N_16094,N_11597,N_14890);
and U16095 (N_16095,N_12007,N_12547);
nor U16096 (N_16096,N_13358,N_11346);
nand U16097 (N_16097,N_13135,N_12916);
nand U16098 (N_16098,N_11348,N_11285);
or U16099 (N_16099,N_12144,N_12306);
and U16100 (N_16100,N_14584,N_11970);
and U16101 (N_16101,N_10714,N_11790);
and U16102 (N_16102,N_12559,N_14625);
or U16103 (N_16103,N_13865,N_13650);
or U16104 (N_16104,N_11089,N_10728);
and U16105 (N_16105,N_12335,N_12715);
nand U16106 (N_16106,N_13153,N_13561);
nand U16107 (N_16107,N_14424,N_13158);
nand U16108 (N_16108,N_14867,N_10395);
xor U16109 (N_16109,N_12699,N_10912);
nor U16110 (N_16110,N_11772,N_11431);
or U16111 (N_16111,N_14613,N_13366);
and U16112 (N_16112,N_10942,N_13712);
and U16113 (N_16113,N_12511,N_12608);
and U16114 (N_16114,N_14507,N_14465);
nand U16115 (N_16115,N_13184,N_14017);
nor U16116 (N_16116,N_14110,N_13513);
nand U16117 (N_16117,N_11314,N_13915);
or U16118 (N_16118,N_12959,N_12691);
and U16119 (N_16119,N_14241,N_11911);
or U16120 (N_16120,N_14339,N_12414);
and U16121 (N_16121,N_14527,N_13442);
and U16122 (N_16122,N_11661,N_14645);
nand U16123 (N_16123,N_13458,N_14768);
nor U16124 (N_16124,N_12889,N_10661);
or U16125 (N_16125,N_13880,N_12648);
nand U16126 (N_16126,N_12843,N_10355);
and U16127 (N_16127,N_11292,N_11399);
nor U16128 (N_16128,N_12894,N_12107);
or U16129 (N_16129,N_13497,N_11521);
nand U16130 (N_16130,N_10947,N_10361);
nor U16131 (N_16131,N_10732,N_10150);
or U16132 (N_16132,N_13913,N_12592);
or U16133 (N_16133,N_14166,N_11187);
nor U16134 (N_16134,N_12604,N_11087);
xnor U16135 (N_16135,N_14077,N_11358);
nor U16136 (N_16136,N_13309,N_12655);
or U16137 (N_16137,N_14711,N_11648);
nand U16138 (N_16138,N_13351,N_14433);
nor U16139 (N_16139,N_10003,N_11135);
or U16140 (N_16140,N_10155,N_11807);
nor U16141 (N_16141,N_12300,N_11773);
and U16142 (N_16142,N_10431,N_12514);
nand U16143 (N_16143,N_14588,N_11022);
and U16144 (N_16144,N_11344,N_14788);
xor U16145 (N_16145,N_10232,N_13280);
or U16146 (N_16146,N_14638,N_13271);
or U16147 (N_16147,N_13039,N_11859);
and U16148 (N_16148,N_10710,N_10013);
and U16149 (N_16149,N_12184,N_12538);
and U16150 (N_16150,N_11211,N_12133);
nand U16151 (N_16151,N_14134,N_12459);
nor U16152 (N_16152,N_13116,N_14039);
xnor U16153 (N_16153,N_10515,N_13304);
and U16154 (N_16154,N_13432,N_10054);
and U16155 (N_16155,N_13373,N_10041);
nor U16156 (N_16156,N_12885,N_13298);
and U16157 (N_16157,N_10411,N_11127);
nor U16158 (N_16158,N_11795,N_11739);
xnor U16159 (N_16159,N_13938,N_10527);
or U16160 (N_16160,N_10111,N_11818);
nor U16161 (N_16161,N_13530,N_14985);
nor U16162 (N_16162,N_12213,N_13579);
nand U16163 (N_16163,N_12097,N_10103);
nand U16164 (N_16164,N_12721,N_11308);
and U16165 (N_16165,N_14957,N_13633);
or U16166 (N_16166,N_12116,N_10137);
or U16167 (N_16167,N_14204,N_14292);
and U16168 (N_16168,N_10557,N_12573);
nor U16169 (N_16169,N_13849,N_12835);
nand U16170 (N_16170,N_10570,N_11461);
and U16171 (N_16171,N_11684,N_11097);
nand U16172 (N_16172,N_13762,N_10129);
nor U16173 (N_16173,N_10796,N_14229);
nand U16174 (N_16174,N_11404,N_11656);
or U16175 (N_16175,N_12358,N_14573);
or U16176 (N_16176,N_10638,N_14956);
or U16177 (N_16177,N_14951,N_10976);
nand U16178 (N_16178,N_12897,N_14840);
nor U16179 (N_16179,N_13820,N_13527);
nand U16180 (N_16180,N_13584,N_12674);
nand U16181 (N_16181,N_13873,N_13902);
or U16182 (N_16182,N_11752,N_10001);
xnor U16183 (N_16183,N_10752,N_12745);
nand U16184 (N_16184,N_10860,N_13565);
nand U16185 (N_16185,N_12820,N_10367);
nor U16186 (N_16186,N_14540,N_11164);
or U16187 (N_16187,N_10368,N_11391);
and U16188 (N_16188,N_10051,N_13713);
or U16189 (N_16189,N_12115,N_11563);
and U16190 (N_16190,N_13013,N_12298);
and U16191 (N_16191,N_11312,N_10949);
or U16192 (N_16192,N_10579,N_14720);
nor U16193 (N_16193,N_14167,N_14799);
or U16194 (N_16194,N_12421,N_11881);
xnor U16195 (N_16195,N_12683,N_13640);
nor U16196 (N_16196,N_11354,N_12785);
or U16197 (N_16197,N_14208,N_12113);
nand U16198 (N_16198,N_10273,N_13276);
nand U16199 (N_16199,N_14804,N_12825);
and U16200 (N_16200,N_11082,N_10157);
and U16201 (N_16201,N_11368,N_13349);
nand U16202 (N_16202,N_12228,N_13129);
nand U16203 (N_16203,N_10369,N_13611);
nand U16204 (N_16204,N_11610,N_12487);
nor U16205 (N_16205,N_10805,N_10525);
nand U16206 (N_16206,N_10793,N_10928);
nor U16207 (N_16207,N_11179,N_14823);
xnor U16208 (N_16208,N_13160,N_13680);
nor U16209 (N_16209,N_14253,N_10126);
or U16210 (N_16210,N_11666,N_13064);
nor U16211 (N_16211,N_11035,N_13508);
nand U16212 (N_16212,N_11671,N_14533);
nor U16213 (N_16213,N_12632,N_14463);
and U16214 (N_16214,N_13342,N_10958);
or U16215 (N_16215,N_11026,N_10039);
and U16216 (N_16216,N_13991,N_14434);
and U16217 (N_16217,N_14722,N_13278);
nor U16218 (N_16218,N_13672,N_12522);
nand U16219 (N_16219,N_12451,N_10025);
or U16220 (N_16220,N_11226,N_14539);
and U16221 (N_16221,N_11333,N_12817);
or U16222 (N_16222,N_12749,N_14079);
and U16223 (N_16223,N_12315,N_13889);
and U16224 (N_16224,N_10819,N_12286);
or U16225 (N_16225,N_12150,N_14513);
nand U16226 (N_16226,N_12050,N_10252);
or U16227 (N_16227,N_13447,N_14171);
and U16228 (N_16228,N_14479,N_13500);
or U16229 (N_16229,N_10344,N_11477);
and U16230 (N_16230,N_14917,N_11070);
nor U16231 (N_16231,N_10789,N_14384);
nand U16232 (N_16232,N_12709,N_13021);
nor U16233 (N_16233,N_14267,N_12913);
nor U16234 (N_16234,N_11490,N_11607);
nand U16235 (N_16235,N_12162,N_14669);
nand U16236 (N_16236,N_14866,N_13480);
xor U16237 (N_16237,N_11329,N_12665);
and U16238 (N_16238,N_12982,N_11244);
or U16239 (N_16239,N_10023,N_11124);
and U16240 (N_16240,N_13336,N_10857);
and U16241 (N_16241,N_13176,N_14194);
and U16242 (N_16242,N_11161,N_10914);
or U16243 (N_16243,N_12188,N_13157);
and U16244 (N_16244,N_11243,N_10967);
nand U16245 (N_16245,N_13341,N_14346);
nand U16246 (N_16246,N_12312,N_10376);
nand U16247 (N_16247,N_12960,N_11444);
or U16248 (N_16248,N_14965,N_11455);
and U16249 (N_16249,N_11487,N_10406);
or U16250 (N_16250,N_13090,N_11745);
and U16251 (N_16251,N_10297,N_11267);
or U16252 (N_16252,N_14623,N_13910);
nor U16253 (N_16253,N_10716,N_13674);
or U16254 (N_16254,N_11427,N_13608);
nor U16255 (N_16255,N_13150,N_13839);
nor U16256 (N_16256,N_13295,N_14706);
nor U16257 (N_16257,N_14843,N_13789);
nor U16258 (N_16258,N_11737,N_10351);
or U16259 (N_16259,N_14114,N_13857);
nor U16260 (N_16260,N_10522,N_14230);
and U16261 (N_16261,N_12501,N_14962);
nand U16262 (N_16262,N_13637,N_12638);
or U16263 (N_16263,N_12593,N_13628);
nand U16264 (N_16264,N_10508,N_11357);
nand U16265 (N_16265,N_11594,N_12588);
nand U16266 (N_16266,N_11023,N_14971);
and U16267 (N_16267,N_11967,N_10452);
or U16268 (N_16268,N_12132,N_12950);
and U16269 (N_16269,N_13134,N_13659);
xor U16270 (N_16270,N_14647,N_14736);
nand U16271 (N_16271,N_13360,N_14074);
nand U16272 (N_16272,N_13532,N_11554);
nand U16273 (N_16273,N_10963,N_14680);
nor U16274 (N_16274,N_14868,N_13152);
and U16275 (N_16275,N_14907,N_11649);
nor U16276 (N_16276,N_13065,N_11930);
nand U16277 (N_16277,N_14464,N_10283);
nand U16278 (N_16278,N_12735,N_12694);
xnor U16279 (N_16279,N_14651,N_13370);
nand U16280 (N_16280,N_14160,N_10511);
nor U16281 (N_16281,N_13189,N_10319);
nor U16282 (N_16282,N_10227,N_12435);
nor U16283 (N_16283,N_10274,N_11387);
nand U16284 (N_16284,N_10575,N_10775);
nor U16285 (N_16285,N_14390,N_13055);
nand U16286 (N_16286,N_10445,N_14508);
or U16287 (N_16287,N_10375,N_12004);
xnor U16288 (N_16288,N_12637,N_11015);
and U16289 (N_16289,N_11207,N_10168);
and U16290 (N_16290,N_13572,N_14352);
or U16291 (N_16291,N_12314,N_14824);
nor U16292 (N_16292,N_11450,N_12955);
nand U16293 (N_16293,N_10418,N_13392);
nor U16294 (N_16294,N_13197,N_14068);
and U16295 (N_16295,N_11885,N_14891);
nand U16296 (N_16296,N_10363,N_14192);
nor U16297 (N_16297,N_11893,N_14812);
or U16298 (N_16298,N_12035,N_14530);
nor U16299 (N_16299,N_12585,N_14251);
or U16300 (N_16300,N_13856,N_14936);
and U16301 (N_16301,N_10492,N_12369);
and U16302 (N_16302,N_11707,N_10151);
nor U16303 (N_16303,N_11242,N_10837);
nor U16304 (N_16304,N_14408,N_10765);
or U16305 (N_16305,N_10354,N_14922);
nor U16306 (N_16306,N_11409,N_14438);
and U16307 (N_16307,N_13823,N_11793);
nor U16308 (N_16308,N_11282,N_11650);
nand U16309 (N_16309,N_12389,N_14108);
and U16310 (N_16310,N_13971,N_12438);
and U16311 (N_16311,N_11938,N_13829);
nand U16312 (N_16312,N_10776,N_12729);
nand U16313 (N_16313,N_11641,N_12720);
xor U16314 (N_16314,N_11592,N_11978);
or U16315 (N_16315,N_11189,N_12697);
or U16316 (N_16316,N_11608,N_11322);
nand U16317 (N_16317,N_11800,N_11128);
and U16318 (N_16318,N_12972,N_12841);
or U16319 (N_16319,N_10284,N_14739);
and U16320 (N_16320,N_10287,N_11882);
nand U16321 (N_16321,N_13167,N_13287);
or U16322 (N_16322,N_13891,N_10000);
nand U16323 (N_16323,N_10323,N_13260);
nand U16324 (N_16324,N_14630,N_14607);
or U16325 (N_16325,N_14440,N_12931);
nor U16326 (N_16326,N_13097,N_12236);
and U16327 (N_16327,N_14693,N_12862);
and U16328 (N_16328,N_13092,N_12718);
and U16329 (N_16329,N_14299,N_13404);
or U16330 (N_16330,N_13179,N_10132);
xor U16331 (N_16331,N_13679,N_10270);
or U16332 (N_16332,N_14598,N_14026);
nor U16333 (N_16333,N_14093,N_13118);
nor U16334 (N_16334,N_10223,N_12498);
and U16335 (N_16335,N_14856,N_11944);
nor U16336 (N_16336,N_11858,N_10251);
nor U16337 (N_16337,N_14581,N_13174);
or U16338 (N_16338,N_14022,N_11663);
or U16339 (N_16339,N_11949,N_12610);
or U16340 (N_16340,N_14232,N_10718);
nor U16341 (N_16341,N_11341,N_14012);
nor U16342 (N_16342,N_14234,N_13096);
nand U16343 (N_16343,N_13374,N_14656);
nand U16344 (N_16344,N_14457,N_14587);
nor U16345 (N_16345,N_14069,N_11383);
nand U16346 (N_16346,N_12270,N_10610);
nand U16347 (N_16347,N_13263,N_13707);
nor U16348 (N_16348,N_10951,N_14531);
or U16349 (N_16349,N_13050,N_12381);
nand U16350 (N_16350,N_11645,N_10133);
or U16351 (N_16351,N_10422,N_10200);
or U16352 (N_16352,N_14482,N_13604);
and U16353 (N_16353,N_10959,N_10931);
and U16354 (N_16354,N_12768,N_11258);
nand U16355 (N_16355,N_11763,N_11543);
and U16356 (N_16356,N_14073,N_12943);
nand U16357 (N_16357,N_11401,N_12672);
nor U16358 (N_16358,N_10288,N_12118);
nor U16359 (N_16359,N_12344,N_11974);
nor U16360 (N_16360,N_10272,N_12786);
or U16361 (N_16361,N_14478,N_12505);
or U16362 (N_16362,N_12813,N_13460);
nor U16363 (N_16363,N_13731,N_11274);
or U16364 (N_16364,N_14671,N_11647);
or U16365 (N_16365,N_14520,N_12478);
nor U16366 (N_16366,N_13131,N_10020);
or U16367 (N_16367,N_13747,N_11925);
nor U16368 (N_16368,N_10179,N_13223);
and U16369 (N_16369,N_12316,N_14271);
or U16370 (N_16370,N_14131,N_10311);
nor U16371 (N_16371,N_13005,N_14529);
nand U16372 (N_16372,N_13735,N_12527);
nor U16373 (N_16373,N_13776,N_13722);
nor U16374 (N_16374,N_10868,N_13990);
and U16375 (N_16375,N_10526,N_12865);
or U16376 (N_16376,N_11965,N_11945);
nor U16377 (N_16377,N_11272,N_10472);
nor U16378 (N_16378,N_11382,N_14793);
and U16379 (N_16379,N_13367,N_11186);
or U16380 (N_16380,N_10879,N_14085);
nand U16381 (N_16381,N_11778,N_10903);
and U16382 (N_16382,N_11540,N_10780);
nor U16383 (N_16383,N_14621,N_13761);
or U16384 (N_16384,N_12974,N_14209);
and U16385 (N_16385,N_10465,N_12397);
nand U16386 (N_16386,N_12863,N_12042);
nor U16387 (N_16387,N_13415,N_13413);
and U16388 (N_16388,N_14111,N_11424);
nor U16389 (N_16389,N_14078,N_11643);
nand U16390 (N_16390,N_13045,N_12196);
and U16391 (N_16391,N_11804,N_12175);
nand U16392 (N_16392,N_13024,N_11435);
and U16393 (N_16393,N_10315,N_10520);
and U16394 (N_16394,N_14282,N_14961);
nor U16395 (N_16395,N_10108,N_14817);
nor U16396 (N_16396,N_10147,N_12470);
or U16397 (N_16397,N_11248,N_11498);
nor U16398 (N_16398,N_10349,N_14660);
nor U16399 (N_16399,N_10705,N_11861);
and U16400 (N_16400,N_14090,N_14291);
nor U16401 (N_16401,N_13802,N_11462);
and U16402 (N_16402,N_10121,N_12065);
or U16403 (N_16403,N_12262,N_12870);
or U16404 (N_16404,N_14724,N_10217);
or U16405 (N_16405,N_13694,N_11008);
nor U16406 (N_16406,N_12098,N_13900);
nand U16407 (N_16407,N_14473,N_10606);
and U16408 (N_16408,N_12710,N_11808);
or U16409 (N_16409,N_11299,N_13363);
and U16410 (N_16410,N_10049,N_10740);
or U16411 (N_16411,N_11939,N_12106);
nor U16412 (N_16412,N_10119,N_12905);
nor U16413 (N_16413,N_14140,N_12753);
nand U16414 (N_16414,N_10073,N_13557);
nor U16415 (N_16415,N_14905,N_11840);
or U16416 (N_16416,N_13022,N_12323);
and U16417 (N_16417,N_13645,N_11776);
nor U16418 (N_16418,N_11516,N_10877);
nor U16419 (N_16419,N_13169,N_14343);
and U16420 (N_16420,N_11046,N_12550);
or U16421 (N_16421,N_10981,N_14979);
or U16422 (N_16422,N_10487,N_13544);
or U16423 (N_16423,N_12173,N_12159);
and U16424 (N_16424,N_10485,N_12424);
or U16425 (N_16425,N_14227,N_12480);
nand U16426 (N_16426,N_11596,N_10774);
or U16427 (N_16427,N_14795,N_10408);
nor U16428 (N_16428,N_11644,N_11673);
and U16429 (N_16429,N_14279,N_13509);
and U16430 (N_16430,N_10424,N_12941);
or U16431 (N_16431,N_11977,N_14072);
nor U16432 (N_16432,N_11145,N_11071);
nand U16433 (N_16433,N_14819,N_11474);
or U16434 (N_16434,N_13888,N_12712);
and U16435 (N_16435,N_14653,N_13983);
and U16436 (N_16436,N_13478,N_14013);
nand U16437 (N_16437,N_11589,N_14860);
nand U16438 (N_16438,N_12310,N_10441);
or U16439 (N_16439,N_14889,N_12933);
nand U16440 (N_16440,N_10442,N_12018);
nor U16441 (N_16441,N_13979,N_11509);
nand U16442 (N_16442,N_10463,N_14500);
nor U16443 (N_16443,N_11646,N_12887);
and U16444 (N_16444,N_14284,N_13183);
nand U16445 (N_16445,N_13875,N_12695);
nand U16446 (N_16446,N_13250,N_13044);
or U16447 (N_16447,N_14486,N_12351);
nand U16448 (N_16448,N_10717,N_13381);
nand U16449 (N_16449,N_10085,N_11117);
nand U16450 (N_16450,N_12652,N_13940);
or U16451 (N_16451,N_11686,N_10577);
or U16452 (N_16452,N_12828,N_11083);
nand U16453 (N_16453,N_11532,N_11268);
nor U16454 (N_16454,N_14738,N_13106);
and U16455 (N_16455,N_14239,N_11445);
or U16456 (N_16456,N_13204,N_12210);
nand U16457 (N_16457,N_13311,N_13448);
xnor U16458 (N_16458,N_11953,N_14818);
and U16459 (N_16459,N_10396,N_12601);
or U16460 (N_16460,N_13300,N_11254);
and U16461 (N_16461,N_10703,N_13816);
or U16462 (N_16462,N_12716,N_10335);
nand U16463 (N_16463,N_12085,N_13704);
nand U16464 (N_16464,N_10482,N_11672);
or U16465 (N_16465,N_14334,N_11253);
xor U16466 (N_16466,N_12748,N_13268);
nor U16467 (N_16467,N_13533,N_13256);
or U16468 (N_16468,N_10867,N_12907);
and U16469 (N_16469,N_12229,N_13459);
xnor U16470 (N_16470,N_10628,N_14597);
nand U16471 (N_16471,N_14324,N_12328);
or U16472 (N_16472,N_12231,N_10182);
and U16473 (N_16473,N_11526,N_10427);
or U16474 (N_16474,N_12541,N_10952);
or U16475 (N_16475,N_14541,N_13861);
nor U16476 (N_16476,N_12245,N_14485);
nand U16477 (N_16477,N_11113,N_13331);
and U16478 (N_16478,N_12548,N_10142);
nor U16479 (N_16479,N_13293,N_12206);
xor U16480 (N_16480,N_10494,N_11981);
and U16481 (N_16481,N_11017,N_12624);
nor U16482 (N_16482,N_11711,N_14170);
nor U16483 (N_16483,N_11168,N_14210);
xnor U16484 (N_16484,N_10169,N_10687);
nor U16485 (N_16485,N_11955,N_10767);
and U16486 (N_16486,N_11230,N_11442);
and U16487 (N_16487,N_12940,N_11481);
and U16488 (N_16488,N_12598,N_10292);
nor U16489 (N_16489,N_12290,N_12357);
nand U16490 (N_16490,N_13472,N_11539);
nand U16491 (N_16491,N_11336,N_14923);
and U16492 (N_16492,N_10874,N_14305);
or U16493 (N_16493,N_11961,N_12681);
nand U16494 (N_16494,N_10099,N_13161);
nor U16495 (N_16495,N_13835,N_14419);
xor U16496 (N_16496,N_12432,N_10436);
nor U16497 (N_16497,N_13898,N_10778);
or U16498 (N_16498,N_13112,N_10042);
and U16499 (N_16499,N_12644,N_13607);
nand U16500 (N_16500,N_11385,N_13496);
and U16501 (N_16501,N_14765,N_10380);
nand U16502 (N_16502,N_11309,N_13806);
and U16503 (N_16503,N_13558,N_11289);
or U16504 (N_16504,N_11587,N_11239);
nand U16505 (N_16505,N_10167,N_11891);
nor U16506 (N_16506,N_12158,N_10848);
nor U16507 (N_16507,N_14792,N_12969);
nand U16508 (N_16508,N_14322,N_10725);
or U16509 (N_16509,N_14779,N_13708);
nor U16510 (N_16510,N_11188,N_14996);
and U16511 (N_16511,N_13380,N_12095);
nor U16512 (N_16512,N_14262,N_11843);
or U16513 (N_16513,N_11263,N_14758);
or U16514 (N_16514,N_10191,N_11203);
nor U16515 (N_16515,N_10602,N_12965);
nand U16516 (N_16516,N_11229,N_10925);
nand U16517 (N_16517,N_11940,N_14444);
nand U16518 (N_16518,N_14098,N_10434);
or U16519 (N_16519,N_12038,N_11069);
and U16520 (N_16520,N_13773,N_14959);
nand U16521 (N_16521,N_14094,N_12925);
xnor U16522 (N_16522,N_14021,N_13009);
xnor U16523 (N_16523,N_13274,N_13253);
nand U16524 (N_16524,N_10739,N_12151);
xor U16525 (N_16525,N_11565,N_11942);
xnor U16526 (N_16526,N_12932,N_11576);
nand U16527 (N_16527,N_13155,N_11698);
nand U16528 (N_16528,N_13570,N_13535);
or U16529 (N_16529,N_12394,N_10806);
and U16530 (N_16530,N_11903,N_14304);
or U16531 (N_16531,N_12307,N_13419);
and U16532 (N_16532,N_10836,N_14353);
nor U16533 (N_16533,N_11303,N_10464);
and U16534 (N_16534,N_12525,N_10491);
nand U16535 (N_16535,N_10538,N_14716);
nand U16536 (N_16536,N_12995,N_14662);
and U16537 (N_16537,N_12523,N_13170);
nor U16538 (N_16538,N_11025,N_10783);
nand U16539 (N_16539,N_13528,N_13127);
nand U16540 (N_16540,N_11912,N_12187);
nand U16541 (N_16541,N_10474,N_14593);
nor U16542 (N_16542,N_14411,N_13632);
and U16543 (N_16543,N_13714,N_11888);
nand U16544 (N_16544,N_14570,N_13592);
or U16545 (N_16545,N_12155,N_13724);
or U16546 (N_16546,N_13763,N_10950);
and U16547 (N_16547,N_13649,N_10212);
or U16548 (N_16548,N_11151,N_11018);
and U16549 (N_16549,N_10290,N_10794);
nand U16550 (N_16550,N_13742,N_10847);
nor U16551 (N_16551,N_10562,N_14124);
or U16552 (N_16552,N_14784,N_10704);
nand U16553 (N_16553,N_11897,N_14741);
nand U16554 (N_16554,N_14988,N_10279);
or U16555 (N_16555,N_12555,N_12052);
nor U16556 (N_16556,N_10192,N_14336);
and U16557 (N_16557,N_13222,N_11355);
and U16558 (N_16558,N_10798,N_13955);
nand U16559 (N_16559,N_13732,N_12360);
nor U16560 (N_16560,N_13629,N_12408);
and U16561 (N_16561,N_13914,N_13957);
nand U16562 (N_16562,N_11612,N_13085);
and U16563 (N_16563,N_14903,N_12966);
nor U16564 (N_16564,N_13138,N_14036);
nor U16565 (N_16565,N_11300,N_10258);
xor U16566 (N_16566,N_12849,N_11544);
or U16567 (N_16567,N_13182,N_14455);
xor U16568 (N_16568,N_10830,N_13436);
and U16569 (N_16569,N_14746,N_12311);
nand U16570 (N_16570,N_12805,N_11530);
and U16571 (N_16571,N_13689,N_10974);
and U16572 (N_16572,N_11871,N_11061);
nor U16573 (N_16573,N_13206,N_10978);
or U16574 (N_16574,N_14869,N_14242);
and U16575 (N_16575,N_12973,N_14730);
nor U16576 (N_16576,N_13977,N_11483);
or U16577 (N_16577,N_12821,N_12688);
nand U16578 (N_16578,N_11887,N_10544);
or U16579 (N_16579,N_13438,N_14288);
or U16580 (N_16580,N_14092,N_13627);
and U16581 (N_16581,N_10469,N_12963);
and U16582 (N_16582,N_13493,N_11916);
or U16583 (N_16583,N_11349,N_11935);
or U16584 (N_16584,N_12453,N_11845);
xor U16585 (N_16585,N_12700,N_12433);
or U16586 (N_16586,N_13738,N_14075);
or U16587 (N_16587,N_14019,N_11273);
nand U16588 (N_16588,N_11210,N_12739);
nand U16589 (N_16589,N_11828,N_14425);
nand U16590 (N_16590,N_14842,N_12094);
or U16591 (N_16591,N_13387,N_13317);
nor U16592 (N_16592,N_11931,N_10241);
and U16593 (N_16593,N_10608,N_13673);
and U16594 (N_16594,N_12040,N_14367);
nand U16595 (N_16595,N_11112,N_14163);
nand U16596 (N_16596,N_13969,N_11966);
and U16597 (N_16597,N_12021,N_12855);
nand U16598 (N_16598,N_10024,N_10326);
nor U16599 (N_16599,N_12141,N_11814);
nor U16600 (N_16600,N_10743,N_13948);
or U16601 (N_16601,N_12743,N_13291);
nand U16602 (N_16602,N_10139,N_12707);
xnor U16603 (N_16603,N_13916,N_11706);
or U16604 (N_16604,N_10990,N_10516);
or U16605 (N_16605,N_11702,N_13903);
and U16606 (N_16606,N_14122,N_14756);
nand U16607 (N_16607,N_11510,N_13284);
nand U16608 (N_16608,N_12517,N_12513);
or U16609 (N_16609,N_11213,N_12942);
nand U16610 (N_16610,N_12650,N_12239);
nor U16611 (N_16611,N_12234,N_14215);
nand U16612 (N_16612,N_13431,N_12291);
and U16613 (N_16613,N_10829,N_13817);
and U16614 (N_16614,N_12756,N_10834);
and U16615 (N_16615,N_10823,N_14226);
nor U16616 (N_16616,N_12789,N_13400);
nor U16617 (N_16617,N_11533,N_10745);
and U16618 (N_16618,N_14268,N_10216);
or U16619 (N_16619,N_10324,N_10761);
nor U16620 (N_16620,N_11922,N_10893);
and U16621 (N_16621,N_10264,N_14222);
and U16622 (N_16622,N_13034,N_10980);
or U16623 (N_16623,N_14810,N_14984);
or U16624 (N_16624,N_10618,N_11359);
nor U16625 (N_16625,N_10530,N_13514);
and U16626 (N_16626,N_11262,N_11205);
nand U16627 (N_16627,N_11989,N_12277);
nand U16628 (N_16628,N_14049,N_11496);
nand U16629 (N_16629,N_14040,N_12583);
nor U16630 (N_16630,N_11497,N_12945);
nor U16631 (N_16631,N_13974,N_12803);
nand U16632 (N_16632,N_13098,N_10130);
nor U16633 (N_16633,N_11985,N_12516);
and U16634 (N_16634,N_14453,N_14115);
nor U16635 (N_16635,N_12352,N_12924);
or U16636 (N_16636,N_13001,N_12241);
nor U16637 (N_16637,N_12507,N_13901);
or U16638 (N_16638,N_14003,N_13171);
or U16639 (N_16639,N_13926,N_11172);
and U16640 (N_16640,N_14831,N_13193);
nor U16641 (N_16641,N_14782,N_12170);
nor U16642 (N_16642,N_12512,N_13217);
nor U16643 (N_16643,N_10010,N_11202);
xnor U16644 (N_16644,N_10399,N_12577);
and U16645 (N_16645,N_14471,N_12689);
nand U16646 (N_16646,N_11108,N_12292);
nand U16647 (N_16647,N_11324,N_14301);
and U16648 (N_16648,N_10609,N_14427);
or U16649 (N_16649,N_10327,N_10318);
xor U16650 (N_16650,N_12154,N_10499);
nor U16651 (N_16651,N_13474,N_10559);
or U16652 (N_16652,N_13241,N_12426);
xor U16653 (N_16653,N_13487,N_14484);
and U16654 (N_16654,N_11122,N_12993);
and U16655 (N_16655,N_10671,N_14516);
xor U16656 (N_16656,N_11929,N_14967);
nand U16657 (N_16657,N_10565,N_12567);
or U16658 (N_16658,N_10504,N_14449);
and U16659 (N_16659,N_13590,N_12332);
nand U16660 (N_16660,N_14549,N_14498);
or U16661 (N_16661,N_12227,N_10322);
and U16662 (N_16662,N_14983,N_11789);
nand U16663 (N_16663,N_12760,N_11693);
nand U16664 (N_16664,N_12744,N_12643);
or U16665 (N_16665,N_12104,N_12698);
and U16666 (N_16666,N_13822,N_12831);
and U16667 (N_16667,N_10084,N_14535);
nor U16668 (N_16668,N_13402,N_14043);
and U16669 (N_16669,N_11158,N_14927);
or U16670 (N_16670,N_11153,N_12354);
nand U16671 (N_16671,N_14670,N_12143);
and U16672 (N_16672,N_10986,N_14718);
and U16673 (N_16673,N_10968,N_10859);
nor U16674 (N_16674,N_11340,N_10128);
and U16675 (N_16675,N_13376,N_14858);
and U16676 (N_16676,N_13477,N_10498);
nor U16677 (N_16677,N_12666,N_11079);
xor U16678 (N_16678,N_14737,N_14128);
nand U16679 (N_16679,N_14365,N_14280);
and U16680 (N_16680,N_14674,N_13130);
nor U16681 (N_16681,N_14123,N_14290);
and U16682 (N_16682,N_11315,N_10507);
and U16683 (N_16683,N_11777,N_11712);
and U16684 (N_16684,N_10186,N_11380);
nor U16685 (N_16685,N_14960,N_10009);
nand U16686 (N_16686,N_14663,N_13988);
nor U16687 (N_16687,N_13618,N_11430);
nor U16688 (N_16688,N_11561,N_13040);
nor U16689 (N_16689,N_11339,N_13441);
or U16690 (N_16690,N_13405,N_10159);
or U16691 (N_16691,N_14348,N_12682);
or U16692 (N_16692,N_14412,N_11287);
nand U16693 (N_16693,N_11937,N_13056);
nand U16694 (N_16694,N_11849,N_11219);
or U16695 (N_16695,N_11171,N_10617);
nand U16696 (N_16696,N_11014,N_12427);
or U16697 (N_16697,N_14161,N_11884);
or U16698 (N_16698,N_13872,N_11278);
nand U16699 (N_16699,N_14351,N_14764);
nor U16700 (N_16700,N_14995,N_10231);
nor U16701 (N_16701,N_13261,N_13966);
nor U16702 (N_16702,N_13368,N_14945);
nor U16703 (N_16703,N_10909,N_12769);
and U16704 (N_16704,N_14309,N_13195);
nor U16705 (N_16705,N_12784,N_10019);
or U16706 (N_16706,N_10458,N_11958);
or U16707 (N_16707,N_11606,N_10012);
or U16708 (N_16708,N_14445,N_10882);
and U16709 (N_16709,N_14841,N_11664);
nand U16710 (N_16710,N_11337,N_12081);
and U16711 (N_16711,N_13481,N_13353);
xor U16712 (N_16712,N_10329,N_14859);
or U16713 (N_16713,N_10235,N_10647);
or U16714 (N_16714,N_14105,N_12703);
and U16715 (N_16715,N_10832,N_10810);
nor U16716 (N_16716,N_13933,N_13473);
nor U16717 (N_16717,N_12077,N_10239);
nor U16718 (N_16718,N_13571,N_13079);
xor U16719 (N_16719,N_12952,N_11283);
nor U16720 (N_16720,N_12466,N_11771);
and U16721 (N_16721,N_14976,N_10685);
or U16722 (N_16722,N_10996,N_12733);
nor U16723 (N_16723,N_10460,N_13427);
or U16724 (N_16724,N_11682,N_10407);
nand U16725 (N_16725,N_13283,N_13924);
or U16726 (N_16726,N_10307,N_14101);
nor U16727 (N_16727,N_12242,N_12020);
nand U16728 (N_16728,N_10861,N_11551);
nand U16729 (N_16729,N_14300,N_10741);
nor U16730 (N_16730,N_11414,N_13344);
and U16731 (N_16731,N_11821,N_10509);
nor U16732 (N_16732,N_12882,N_11326);
or U16733 (N_16733,N_14276,N_11209);
nor U16734 (N_16734,N_10659,N_12569);
or U16735 (N_16735,N_11847,N_10850);
or U16736 (N_16736,N_11491,N_10759);
nand U16737 (N_16737,N_11927,N_14879);
nand U16738 (N_16738,N_12302,N_11197);
nand U16739 (N_16739,N_11908,N_10962);
nor U16740 (N_16740,N_13369,N_11378);
and U16741 (N_16741,N_12373,N_11335);
nor U16742 (N_16742,N_12412,N_10979);
or U16743 (N_16743,N_10238,N_13347);
or U16744 (N_16744,N_10100,N_11616);
and U16745 (N_16745,N_14490,N_14307);
nand U16746 (N_16746,N_12937,N_10359);
and U16747 (N_16747,N_10325,N_11343);
nor U16748 (N_16748,N_10757,N_13314);
nor U16749 (N_16749,N_12468,N_14225);
and U16750 (N_16750,N_12502,N_11926);
and U16751 (N_16751,N_12854,N_12103);
nand U16752 (N_16752,N_14622,N_11101);
or U16753 (N_16753,N_12334,N_11581);
nand U16754 (N_16754,N_10887,N_14873);
xnor U16755 (N_16755,N_13219,N_14501);
nand U16756 (N_16756,N_13624,N_10632);
nand U16757 (N_16757,N_12758,N_13581);
and U16758 (N_16758,N_12968,N_10047);
and U16759 (N_16759,N_13524,N_11169);
or U16760 (N_16760,N_12139,N_14302);
or U16761 (N_16761,N_13603,N_13164);
and U16762 (N_16762,N_14954,N_14377);
and U16763 (N_16763,N_14955,N_12500);
or U16764 (N_16764,N_13246,N_11377);
nor U16765 (N_16765,N_13030,N_13729);
and U16766 (N_16766,N_11156,N_12833);
nand U16767 (N_16767,N_10625,N_14911);
nand U16768 (N_16768,N_14127,N_11542);
xor U16769 (N_16769,N_13457,N_13517);
and U16770 (N_16770,N_11478,N_13987);
and U16771 (N_16771,N_11010,N_10265);
nor U16772 (N_16772,N_12253,N_12034);
nor U16773 (N_16773,N_10502,N_14589);
or U16774 (N_16774,N_13198,N_13788);
or U16775 (N_16775,N_11162,N_12656);
or U16776 (N_16776,N_11237,N_13675);
or U16777 (N_16777,N_14245,N_13923);
or U16778 (N_16778,N_13338,N_10500);
or U16779 (N_16779,N_14383,N_11534);
nand U16780 (N_16780,N_14183,N_12380);
xnor U16781 (N_16781,N_12274,N_11796);
nor U16782 (N_16782,N_14502,N_11180);
and U16783 (N_16783,N_10689,N_10066);
nor U16784 (N_16784,N_14794,N_14396);
and U16785 (N_16785,N_13095,N_13125);
nor U16786 (N_16786,N_13421,N_14635);
or U16787 (N_16787,N_11896,N_14608);
and U16788 (N_16788,N_13277,N_12896);
nor U16789 (N_16789,N_13320,N_11105);
or U16790 (N_16790,N_13196,N_12807);
nand U16791 (N_16791,N_10827,N_13463);
and U16792 (N_16792,N_11252,N_10561);
nor U16793 (N_16793,N_14978,N_14652);
nor U16794 (N_16794,N_13289,N_14416);
nor U16795 (N_16795,N_14337,N_11279);
or U16796 (N_16796,N_14272,N_12048);
nand U16797 (N_16797,N_13429,N_12071);
xnor U16798 (N_16798,N_14466,N_13072);
nand U16799 (N_16799,N_13858,N_14968);
or U16800 (N_16800,N_14247,N_12587);
and U16801 (N_16801,N_11783,N_14729);
nand U16802 (N_16802,N_13037,N_12362);
nand U16803 (N_16803,N_10426,N_13099);
or U16804 (N_16804,N_11566,N_11421);
or U16805 (N_16805,N_10585,N_11148);
nand U16806 (N_16806,N_14676,N_12388);
nand U16807 (N_16807,N_11810,N_14061);
and U16808 (N_16808,N_10257,N_10303);
or U16809 (N_16809,N_13582,N_13682);
nor U16810 (N_16810,N_11564,N_11296);
and U16811 (N_16811,N_10748,N_14364);
nor U16812 (N_16812,N_13696,N_13177);
nor U16813 (N_16813,N_11837,N_10306);
xnor U16814 (N_16814,N_13082,N_12477);
nor U16815 (N_16815,N_13490,N_10339);
or U16816 (N_16816,N_13909,N_10640);
or U16817 (N_16817,N_14998,N_10691);
and U16818 (N_16818,N_12448,N_13187);
nand U16819 (N_16819,N_13567,N_10842);
and U16820 (N_16820,N_14223,N_12110);
or U16821 (N_16821,N_13663,N_13982);
and U16822 (N_16822,N_14388,N_13754);
nand U16823 (N_16823,N_11695,N_12766);
nor U16824 (N_16824,N_11499,N_10435);
nor U16825 (N_16825,N_12326,N_14913);
nor U16826 (N_16826,N_12642,N_11126);
and U16827 (N_16827,N_14174,N_10055);
nor U16828 (N_16828,N_13071,N_14562);
and U16829 (N_16829,N_10082,N_12398);
or U16830 (N_16830,N_12069,N_10713);
and U16831 (N_16831,N_13305,N_12600);
or U16832 (N_16832,N_13166,N_13847);
xnor U16833 (N_16833,N_11362,N_12861);
nand U16834 (N_16834,N_13313,N_14158);
and U16835 (N_16835,N_12795,N_13407);
nand U16836 (N_16836,N_14286,N_14561);
nand U16837 (N_16837,N_13228,N_11306);
nor U16838 (N_16838,N_12075,N_13779);
and U16839 (N_16839,N_10173,N_11894);
nand U16840 (N_16840,N_14185,N_13038);
nor U16841 (N_16841,N_12070,N_10960);
nand U16842 (N_16842,N_10087,N_10026);
nand U16843 (N_16843,N_11552,N_12992);
or U16844 (N_16844,N_10405,N_12348);
nand U16845 (N_16845,N_14330,N_10754);
or U16846 (N_16846,N_10224,N_11364);
and U16847 (N_16847,N_14940,N_11742);
nand U16848 (N_16848,N_12579,N_11098);
or U16849 (N_16849,N_11703,N_10593);
or U16850 (N_16850,N_13710,N_11318);
nand U16851 (N_16851,N_12778,N_11479);
or U16852 (N_16852,N_13444,N_13594);
nand U16853 (N_16853,N_13465,N_13355);
or U16854 (N_16854,N_11092,N_11577);
nor U16855 (N_16855,N_14898,N_13741);
nand U16856 (N_16856,N_14950,N_10818);
or U16857 (N_16857,N_10475,N_12486);
nor U16858 (N_16858,N_10811,N_12692);
or U16859 (N_16859,N_11720,N_14715);
nand U16860 (N_16860,N_14244,N_13389);
nor U16861 (N_16861,N_12705,N_12627);
and U16862 (N_16862,N_11750,N_11176);
and U16863 (N_16863,N_10506,N_14494);
and U16864 (N_16864,N_13019,N_12022);
or U16865 (N_16865,N_13214,N_11488);
or U16866 (N_16866,N_10388,N_11531);
or U16867 (N_16867,N_10890,N_10934);
nand U16868 (N_16868,N_10712,N_14298);
nand U16869 (N_16869,N_12690,N_12647);
nand U16870 (N_16870,N_12521,N_14789);
or U16871 (N_16871,N_14357,N_12537);
or U16872 (N_16872,N_10038,N_14837);
xnor U16873 (N_16873,N_14402,N_11330);
nor U16874 (N_16874,N_10336,N_10572);
nand U16875 (N_16875,N_14255,N_11441);
or U16876 (N_16876,N_13746,N_11740);
nor U16877 (N_16877,N_13578,N_13484);
and U16878 (N_16878,N_14566,N_10615);
nand U16879 (N_16879,N_12670,N_10866);
and U16880 (N_16880,N_10889,N_10081);
xor U16881 (N_16881,N_12497,N_14474);
nand U16882 (N_16882,N_11007,N_14579);
nand U16883 (N_16883,N_13766,N_11265);
or U16884 (N_16884,N_13621,N_11864);
xor U16885 (N_16885,N_14634,N_13967);
nor U16886 (N_16886,N_10248,N_12658);
nand U16887 (N_16887,N_12938,N_12533);
and U16888 (N_16888,N_13778,N_14488);
nor U16889 (N_16889,N_10872,N_11096);
nand U16890 (N_16890,N_11458,N_10666);
and U16891 (N_16891,N_10372,N_13133);
and U16892 (N_16892,N_12490,N_12771);
or U16893 (N_16893,N_11048,N_10152);
nand U16894 (N_16894,N_10699,N_10462);
or U16895 (N_16895,N_12846,N_11467);
nor U16896 (N_16896,N_11173,N_14363);
nand U16897 (N_16897,N_11003,N_14212);
or U16898 (N_16898,N_10412,N_12667);
or U16899 (N_16899,N_14734,N_10841);
nand U16900 (N_16900,N_11396,N_10957);
nand U16901 (N_16901,N_11954,N_14059);
nand U16902 (N_16902,N_11500,N_12190);
or U16903 (N_16903,N_10835,N_10172);
or U16904 (N_16904,N_11873,N_10206);
nor U16905 (N_16905,N_13212,N_14845);
and U16906 (N_16906,N_14863,N_12454);
nor U16907 (N_16907,N_10414,N_12343);
nand U16908 (N_16908,N_13781,N_14564);
or U16909 (N_16909,N_13406,N_13326);
and U16910 (N_16910,N_10493,N_14018);
xor U16911 (N_16911,N_14558,N_11257);
and U16912 (N_16912,N_11568,N_13980);
or U16913 (N_16913,N_11403,N_10447);
nand U16914 (N_16914,N_10214,N_12859);
and U16915 (N_16915,N_13871,N_14156);
or U16916 (N_16916,N_12508,N_14081);
nor U16917 (N_16917,N_14801,N_14677);
or U16918 (N_16918,N_14790,N_11088);
and U16919 (N_16919,N_10417,N_10366);
or U16920 (N_16920,N_14116,N_13073);
nor U16921 (N_16921,N_12471,N_11785);
and U16922 (N_16922,N_14496,N_11102);
nand U16923 (N_16923,N_13665,N_13057);
nor U16924 (N_16924,N_12869,N_11068);
and U16925 (N_16925,N_14505,N_12996);
and U16926 (N_16926,N_14015,N_11220);
or U16927 (N_16927,N_11094,N_12669);
nand U16928 (N_16928,N_14606,N_14832);
and U16929 (N_16929,N_13359,N_12301);
nor U16930 (N_16930,N_10486,N_12238);
or U16931 (N_16931,N_13855,N_10029);
or U16932 (N_16932,N_13671,N_10715);
or U16933 (N_16933,N_10700,N_12779);
or U16934 (N_16934,N_10005,N_12321);
and U16935 (N_16935,N_13238,N_14345);
xnor U16936 (N_16936,N_10727,N_11665);
nand U16937 (N_16937,N_14902,N_12898);
and U16938 (N_16938,N_11428,N_14199);
and U16939 (N_16939,N_11177,N_12639);
nand U16940 (N_16940,N_14145,N_10852);
and U16941 (N_16941,N_12921,N_11423);
and U16942 (N_16942,N_12067,N_12331);
nor U16943 (N_16943,N_10253,N_11774);
nor U16944 (N_16944,N_12105,N_12967);
or U16945 (N_16945,N_14851,N_14947);
nor U16946 (N_16946,N_12340,N_13115);
or U16947 (N_16947,N_12294,N_13186);
nand U16948 (N_16948,N_10828,N_13385);
and U16949 (N_16949,N_13868,N_13870);
or U16950 (N_16950,N_11856,N_11327);
or U16951 (N_16951,N_12259,N_10701);
and U16952 (N_16952,N_14155,N_10648);
nand U16953 (N_16953,N_13495,N_10742);
nand U16954 (N_16954,N_12842,N_11370);
or U16955 (N_16955,N_14935,N_13928);
nand U16956 (N_16956,N_10707,N_12282);
nand U16957 (N_16957,N_12675,N_14554);
or U16958 (N_16958,N_11454,N_13563);
or U16959 (N_16959,N_10807,N_10747);
xnor U16960 (N_16960,N_12860,N_11538);
or U16961 (N_16961,N_13257,N_11284);
or U16962 (N_16962,N_10541,N_10300);
nand U16963 (N_16963,N_13231,N_11570);
or U16964 (N_16964,N_14202,N_11256);
and U16965 (N_16965,N_14312,N_13225);
and U16966 (N_16966,N_14404,N_12961);
and U16967 (N_16967,N_14721,N_10437);
nand U16968 (N_16968,N_10148,N_14915);
and U16969 (N_16969,N_11212,N_13003);
nor U16970 (N_16970,N_11622,N_11835);
nor U16971 (N_16971,N_13837,N_10365);
nand U16972 (N_16972,N_14083,N_10007);
nand U16973 (N_16973,N_14733,N_11109);
or U16974 (N_16974,N_13061,N_11824);
nand U16975 (N_16975,N_12629,N_13706);
or U16976 (N_16976,N_12740,N_14610);
nand U16977 (N_16977,N_11436,N_12714);
nor U16978 (N_16978,N_12203,N_11580);
xnor U16979 (N_16979,N_11464,N_14106);
or U16980 (N_16980,N_10779,N_10246);
nor U16981 (N_16981,N_11599,N_12620);
or U16982 (N_16982,N_13798,N_11194);
nand U16983 (N_16983,N_10069,N_13325);
xor U16984 (N_16984,N_11678,N_13831);
nand U16985 (N_16985,N_10551,N_12149);
or U16986 (N_16986,N_14289,N_10512);
nor U16987 (N_16987,N_10478,N_10170);
and U16988 (N_16988,N_12864,N_11291);
nand U16989 (N_16989,N_14757,N_12848);
and U16990 (N_16990,N_13745,N_11055);
nand U16991 (N_16991,N_10539,N_13144);
and U16992 (N_16992,N_11578,N_12686);
or U16993 (N_16993,N_10624,N_10590);
nor U16994 (N_16994,N_14821,N_14992);
nand U16995 (N_16995,N_13272,N_12990);
and U16996 (N_16996,N_10198,N_13602);
or U16997 (N_16997,N_14256,N_13883);
nor U16998 (N_16998,N_11078,N_10105);
and U16999 (N_16999,N_14672,N_12591);
or U17000 (N_17000,N_11802,N_13020);
or U17001 (N_17001,N_11100,N_13782);
nand U17002 (N_17002,N_11747,N_13753);
or U17003 (N_17003,N_12926,N_12495);
nand U17004 (N_17004,N_10031,N_10451);
or U17005 (N_17005,N_13052,N_12379);
nor U17006 (N_17006,N_13023,N_12479);
and U17007 (N_17007,N_14949,N_12558);
and U17008 (N_17008,N_12936,N_10059);
nand U17009 (N_17009,N_14696,N_11301);
and U17010 (N_17010,N_12684,N_11506);
or U17011 (N_17011,N_14278,N_14659);
or U17012 (N_17012,N_13585,N_10946);
nand U17013 (N_17013,N_14525,N_11866);
and U17014 (N_17014,N_13464,N_12419);
nor U17015 (N_17015,N_13717,N_13410);
nand U17016 (N_17016,N_13087,N_13324);
and U17017 (N_17017,N_10135,N_14020);
or U17018 (N_17018,N_11535,N_12726);
nand U17019 (N_17019,N_10177,N_13299);
and U17020 (N_17020,N_14783,N_11834);
and U17021 (N_17021,N_13494,N_12209);
nor U17022 (N_17022,N_10250,N_14375);
nand U17023 (N_17023,N_11218,N_12140);
nand U17024 (N_17024,N_14401,N_11042);
nand U17025 (N_17025,N_14538,N_11667);
or U17026 (N_17026,N_10664,N_10895);
or U17027 (N_17027,N_14308,N_13845);
nor U17028 (N_17028,N_12492,N_14080);
and U17029 (N_17029,N_10720,N_11376);
xnor U17030 (N_17030,N_13885,N_12031);
and U17031 (N_17031,N_14489,N_12134);
nor U17032 (N_17032,N_14643,N_13893);
and U17033 (N_17033,N_14378,N_13876);
nor U17034 (N_17034,N_13010,N_12871);
and U17035 (N_17035,N_14707,N_14436);
and U17036 (N_17036,N_13577,N_11842);
or U17037 (N_17037,N_10202,N_10513);
nand U17038 (N_17038,N_13586,N_14231);
nand U17039 (N_17039,N_14689,N_10795);
and U17040 (N_17040,N_10954,N_10140);
nand U17041 (N_17041,N_14103,N_11115);
and U17042 (N_17042,N_11746,N_14184);
or U17043 (N_17043,N_11389,N_12146);
nand U17044 (N_17044,N_10916,N_11900);
nor U17045 (N_17045,N_12407,N_10678);
nor U17046 (N_17046,N_14235,N_11167);
nor U17047 (N_17047,N_14095,N_12823);
nor U17048 (N_17048,N_14744,N_10940);
and U17049 (N_17049,N_12189,N_12750);
nor U17050 (N_17050,N_14248,N_12461);
xnor U17051 (N_17051,N_11975,N_13580);
nand U17052 (N_17052,N_11137,N_14224);
and U17053 (N_17053,N_13703,N_11973);
nor U17054 (N_17054,N_14544,N_14100);
nor U17055 (N_17055,N_14881,N_10897);
nor U17056 (N_17056,N_14899,N_13453);
nor U17057 (N_17057,N_12181,N_14649);
nand U17058 (N_17058,N_12208,N_11611);
and U17059 (N_17059,N_13613,N_10896);
and U17060 (N_17060,N_11165,N_10537);
or U17061 (N_17061,N_13048,N_13887);
nand U17062 (N_17062,N_13498,N_14982);
nand U17063 (N_17063,N_11373,N_13043);
or U17064 (N_17064,N_12171,N_12017);
or U17065 (N_17065,N_11729,N_11877);
nand U17066 (N_17066,N_10670,N_11987);
or U17067 (N_17067,N_12680,N_11812);
and U17068 (N_17068,N_12429,N_13107);
nand U17069 (N_17069,N_13985,N_14157);
or U17070 (N_17070,N_14695,N_12613);
or U17071 (N_17071,N_14805,N_13920);
nand U17072 (N_17072,N_11053,N_10574);
nand U17073 (N_17073,N_14766,N_10208);
nor U17074 (N_17074,N_11363,N_14118);
and U17075 (N_17075,N_14886,N_12660);
and U17076 (N_17076,N_10158,N_11999);
xor U17077 (N_17077,N_11163,N_14591);
nand U17078 (N_17078,N_14850,N_10199);
and U17079 (N_17079,N_14639,N_11466);
nand U17080 (N_17080,N_12793,N_14888);
nand U17081 (N_17081,N_12895,N_10650);
or U17082 (N_17082,N_13692,N_12978);
or U17083 (N_17083,N_11469,N_14238);
nor U17084 (N_17084,N_11241,N_13636);
or U17085 (N_17085,N_11722,N_11613);
and U17086 (N_17086,N_12775,N_11411);
nand U17087 (N_17087,N_11325,N_14559);
xor U17088 (N_17088,N_13027,N_10995);
or U17089 (N_17089,N_13805,N_14362);
and U17090 (N_17090,N_14190,N_11159);
and U17091 (N_17091,N_10389,N_12003);
and U17092 (N_17092,N_12442,N_10345);
and U17093 (N_17093,N_14063,N_10301);
or U17094 (N_17094,N_13668,N_11353);
nor U17095 (N_17095,N_13906,N_10589);
or U17096 (N_17096,N_12560,N_13867);
nand U17097 (N_17097,N_12772,N_12390);
or U17098 (N_17098,N_14432,N_14698);
nand U17099 (N_17099,N_10052,N_12030);
nand U17100 (N_17100,N_10930,N_14629);
nor U17101 (N_17101,N_11662,N_13993);
nor U17102 (N_17102,N_10006,N_14987);
nand U17103 (N_17103,N_14599,N_12126);
or U17104 (N_17104,N_13943,N_11718);
and U17105 (N_17105,N_14326,N_12368);
nor U17106 (N_17106,N_13264,N_13935);
xor U17107 (N_17107,N_14510,N_12868);
and U17108 (N_17108,N_10800,N_14373);
and U17109 (N_17109,N_14749,N_14552);
and U17110 (N_17110,N_13252,N_10975);
or U17111 (N_17111,N_13927,N_11011);
nand U17112 (N_17112,N_14928,N_10067);
and U17113 (N_17113,N_12008,N_10649);
nor U17114 (N_17114,N_13796,N_13218);
and U17115 (N_17115,N_13210,N_12327);
or U17116 (N_17116,N_12880,N_10340);
and U17117 (N_17117,N_12830,N_13357);
and U17118 (N_17118,N_14697,N_13658);
xor U17119 (N_17119,N_11512,N_11440);
nand U17120 (N_17120,N_14349,N_13807);
or U17121 (N_17121,N_14710,N_12443);
nor U17122 (N_17122,N_10514,N_14148);
or U17123 (N_17123,N_14691,N_14547);
nand U17124 (N_17124,N_12002,N_11247);
nor U17125 (N_17125,N_13301,N_10310);
and U17126 (N_17126,N_14874,N_13337);
nor U17127 (N_17127,N_11475,N_14317);
nand U17128 (N_17128,N_11919,N_13067);
and U17129 (N_17129,N_13362,N_12341);
or U17130 (N_17130,N_14931,N_12618);
nor U17131 (N_17131,N_10933,N_14785);
and U17132 (N_17132,N_14004,N_10218);
and U17133 (N_17133,N_13086,N_10034);
xnor U17134 (N_17134,N_10799,N_14099);
nand U17135 (N_17135,N_13425,N_10534);
or U17136 (N_17136,N_13832,N_10352);
nor U17137 (N_17137,N_14829,N_13451);
nor U17138 (N_17138,N_11317,N_10256);
nor U17139 (N_17139,N_12856,N_10215);
nand U17140 (N_17140,N_13310,N_10476);
nor U17141 (N_17141,N_10654,N_12923);
nand U17142 (N_17142,N_13666,N_10766);
and U17143 (N_17143,N_11620,N_11206);
or U17144 (N_17144,N_10724,N_13244);
or U17145 (N_17145,N_12005,N_10901);
nand U17146 (N_17146,N_13255,N_12582);
nand U17147 (N_17147,N_11907,N_12722);
nand U17148 (N_17148,N_10490,N_10421);
nand U17149 (N_17149,N_11276,N_13275);
nand U17150 (N_17150,N_13012,N_13551);
nand U17151 (N_17151,N_12679,N_10558);
or U17152 (N_17152,N_13850,N_11465);
nand U17153 (N_17153,N_14468,N_14164);
nor U17154 (N_17154,N_12797,N_10419);
nor U17155 (N_17155,N_12400,N_12074);
or U17156 (N_17156,N_10316,N_12350);
nand U17157 (N_17157,N_11831,N_10885);
and U17158 (N_17158,N_10862,N_12284);
xnor U17159 (N_17159,N_11037,N_11553);
and U17160 (N_17160,N_14665,N_12108);
or U17161 (N_17161,N_13690,N_10773);
and U17162 (N_17162,N_10833,N_14964);
or U17163 (N_17163,N_13960,N_12129);
nand U17164 (N_17164,N_14550,N_10298);
and U17165 (N_17165,N_10532,N_12019);
nor U17166 (N_17166,N_10884,N_11076);
nand U17167 (N_17167,N_10630,N_11890);
and U17168 (N_17168,N_10197,N_12578);
and U17169 (N_17169,N_12481,N_12131);
nand U17170 (N_17170,N_12013,N_14694);
or U17171 (N_17171,N_10004,N_10104);
and U17172 (N_17172,N_12402,N_11541);
and U17173 (N_17173,N_12927,N_14991);
nor U17174 (N_17174,N_10568,N_13372);
nor U17175 (N_17175,N_13848,N_12079);
and U17176 (N_17176,N_11792,N_14726);
and U17177 (N_17177,N_14297,N_14314);
and U17178 (N_17178,N_14932,N_13864);
and U17179 (N_17179,N_10357,N_10870);
or U17180 (N_17180,N_13667,N_13290);
nor U17181 (N_17181,N_10738,N_14186);
nand U17182 (N_17182,N_13976,N_14781);
and U17183 (N_17183,N_13750,N_10809);
and U17184 (N_17184,N_13952,N_12440);
or U17185 (N_17185,N_11150,N_12529);
or U17186 (N_17186,N_11144,N_14712);
and U17187 (N_17187,N_12964,N_14154);
or U17188 (N_17188,N_10875,N_13963);
and U17189 (N_17189,N_10428,N_12167);
or U17190 (N_17190,N_12850,N_12386);
or U17191 (N_17191,N_13227,N_13895);
nand U17192 (N_17192,N_11782,N_12420);
nand U17193 (N_17193,N_13191,N_10180);
nand U17194 (N_17194,N_11615,N_11429);
or U17195 (N_17195,N_12232,N_12947);
nand U17196 (N_17196,N_14583,N_11569);
or U17197 (N_17197,N_10873,N_13007);
and U17198 (N_17198,N_14586,N_14011);
and U17199 (N_17199,N_13312,N_14403);
nand U17200 (N_17200,N_11331,N_14056);
and U17201 (N_17201,N_11050,N_14838);
and U17202 (N_17202,N_12989,N_10763);
or U17203 (N_17203,N_10734,N_12342);
or U17204 (N_17204,N_10259,N_10755);
nor U17205 (N_17205,N_12322,N_11350);
nand U17206 (N_17206,N_14654,N_13728);
nand U17207 (N_17207,N_10937,N_13546);
and U17208 (N_17208,N_11451,N_10166);
and U17209 (N_17209,N_14177,N_14458);
or U17210 (N_17210,N_14503,N_12353);
and U17211 (N_17211,N_13553,N_10196);
nand U17212 (N_17212,N_13989,N_14934);
nand U17213 (N_17213,N_11986,N_13555);
nand U17214 (N_17214,N_11452,N_13396);
and U17215 (N_17215,N_14567,N_12717);
and U17216 (N_17216,N_11555,N_12763);
nand U17217 (N_17217,N_10983,N_13482);
nand U17218 (N_17218,N_12983,N_13881);
nor U17219 (N_17219,N_14315,N_14009);
nand U17220 (N_17220,N_13100,N_10911);
and U17221 (N_17221,N_12455,N_12702);
nand U17222 (N_17222,N_14495,N_13726);
or U17223 (N_17223,N_14748,N_11216);
or U17224 (N_17224,N_10244,N_10348);
nor U17225 (N_17225,N_13569,N_10123);
nand U17226 (N_17226,N_12890,N_11106);
or U17227 (N_17227,N_13443,N_11850);
or U17228 (N_17228,N_11550,N_10456);
nor U17229 (N_17229,N_13537,N_13240);
and U17230 (N_17230,N_11052,N_11738);
and U17231 (N_17231,N_12877,N_14572);
or U17232 (N_17232,N_12590,N_13066);
or U17233 (N_17233,N_10358,N_13318);
nand U17234 (N_17234,N_13676,N_11918);
or U17235 (N_17235,N_10646,N_11963);
xnor U17236 (N_17236,N_13715,N_13615);
or U17237 (N_17237,N_11962,N_11034);
nor U17238 (N_17238,N_12039,N_12385);
nor U17239 (N_17239,N_11413,N_13194);
and U17240 (N_17240,N_14657,N_10992);
nor U17241 (N_17241,N_14731,N_10115);
or U17242 (N_17242,N_10668,N_13702);
nand U17243 (N_17243,N_14034,N_13523);
nor U17244 (N_17244,N_13756,N_10240);
and U17245 (N_17245,N_13877,N_13998);
or U17246 (N_17246,N_11714,N_13412);
and U17247 (N_17247,N_12303,N_12911);
or U17248 (N_17248,N_11735,N_10141);
or U17249 (N_17249,N_14872,N_11286);
nor U17250 (N_17250,N_12186,N_13221);
or U17251 (N_17251,N_13614,N_10943);
nor U17252 (N_17252,N_14601,N_10309);
nand U17253 (N_17253,N_11687,N_11119);
or U17254 (N_17254,N_13709,N_11138);
xnor U17255 (N_17255,N_10222,N_12617);
or U17256 (N_17256,N_14620,N_13333);
nand U17257 (N_17257,N_12544,N_11044);
or U17258 (N_17258,N_12444,N_12893);
nand U17259 (N_17259,N_10731,N_11111);
nand U17260 (N_17260,N_13141,N_13011);
or U17261 (N_17261,N_10305,N_14683);
nand U17262 (N_17262,N_12687,N_11446);
nor U17263 (N_17263,N_10183,N_11140);
or U17264 (N_17264,N_13657,N_12662);
nand U17265 (N_17265,N_12276,N_12387);
or U17266 (N_17266,N_10280,N_10397);
and U17267 (N_17267,N_13757,N_10679);
nand U17268 (N_17268,N_13942,N_13434);
nand U17269 (N_17269,N_12755,N_13408);
nor U17270 (N_17270,N_13190,N_14958);
nor U17271 (N_17271,N_10330,N_11889);
or U17272 (N_17272,N_14777,N_11047);
nand U17273 (N_17273,N_11558,N_12751);
or U17274 (N_17274,N_13302,N_14197);
and U17275 (N_17275,N_13684,N_11062);
or U17276 (N_17276,N_14447,N_10663);
and U17277 (N_17277,N_10195,N_14219);
xnor U17278 (N_17278,N_10694,N_12054);
and U17279 (N_17279,N_10964,N_10393);
and U17280 (N_17280,N_12909,N_13230);
nand U17281 (N_17281,N_13545,N_12738);
and U17282 (N_17282,N_13878,N_14311);
xor U17283 (N_17283,N_11784,N_12377);
and U17284 (N_17284,N_10721,N_12063);
and U17285 (N_17285,N_14097,N_11791);
nor U17286 (N_17286,N_10820,N_12093);
nor U17287 (N_17287,N_12984,N_13000);
or U17288 (N_17288,N_13409,N_10733);
nand U17289 (N_17289,N_12258,N_14270);
or U17290 (N_17290,N_10815,N_10797);
or U17291 (N_17291,N_12728,N_13516);
nor U17292 (N_17292,N_12878,N_13178);
nor U17293 (N_17293,N_13647,N_14668);
and U17294 (N_17294,N_10858,N_13992);
and U17295 (N_17295,N_14057,N_11998);
nor U17296 (N_17296,N_14139,N_14673);
or U17297 (N_17297,N_13139,N_11251);
or U17298 (N_17298,N_13538,N_10908);
nand U17299 (N_17299,N_10771,N_13319);
nand U17300 (N_17300,N_10746,N_10941);
nand U17301 (N_17301,N_14658,N_12001);
nand U17302 (N_17302,N_13083,N_11054);
nor U17303 (N_17303,N_10597,N_10846);
and U17304 (N_17304,N_13936,N_10997);
or U17305 (N_17305,N_13599,N_14172);
nor U17306 (N_17306,N_13063,N_12092);
nor U17307 (N_17307,N_10849,N_10015);
and U17308 (N_17308,N_11328,N_10313);
and U17309 (N_17309,N_12792,N_13094);
nand U17310 (N_17310,N_10074,N_10683);
or U17311 (N_17311,N_10521,N_11857);
nor U17312 (N_17312,N_12776,N_12764);
nor U17313 (N_17313,N_11717,N_10802);
or U17314 (N_17314,N_14460,N_12452);
nand U17315 (N_17315,N_11950,N_14667);
nor U17316 (N_17316,N_12551,N_11972);
nand U17317 (N_17317,N_10193,N_14611);
nand U17318 (N_17318,N_14321,N_14269);
nor U17319 (N_17319,N_13511,N_11196);
nand U17320 (N_17320,N_10070,N_12602);
nor U17321 (N_17321,N_11090,N_10751);
nor U17322 (N_17322,N_10863,N_11731);
nand U17323 (N_17323,N_13819,N_14847);
and U17324 (N_17324,N_13688,N_14770);
and U17325 (N_17325,N_12045,N_13018);
nand U17326 (N_17326,N_14441,N_14939);
nor U17327 (N_17327,N_11067,N_14536);
or U17328 (N_17328,N_14295,N_10178);
and U17329 (N_17329,N_12607,N_12064);
nand U17330 (N_17330,N_11293,N_12504);
or U17331 (N_17331,N_14678,N_13725);
nand U17332 (N_17332,N_11867,N_12580);
or U17333 (N_17333,N_10409,N_13279);
nand U17334 (N_17334,N_12366,N_12215);
nand U17335 (N_17335,N_14356,N_11016);
or U17336 (N_17336,N_11964,N_14293);
nand U17337 (N_17337,N_10371,N_10634);
and U17338 (N_17338,N_11471,N_12256);
and U17339 (N_17339,N_11019,N_14451);
nand U17340 (N_17340,N_13587,N_12765);
and U17341 (N_17341,N_11631,N_11811);
nand U17342 (N_17342,N_12401,N_12051);
nor U17343 (N_17343,N_11369,N_13119);
or U17344 (N_17344,N_12641,N_12730);
nor U17345 (N_17345,N_14138,N_12201);
and U17346 (N_17346,N_10991,N_10505);
nand U17347 (N_17347,N_11449,N_13922);
nor U17348 (N_17348,N_14143,N_12028);
and U17349 (N_17349,N_10101,N_14883);
and U17350 (N_17350,N_11994,N_10037);
and U17351 (N_17351,N_11624,N_11231);
or U17352 (N_17352,N_13705,N_13479);
nor U17353 (N_17353,N_10674,N_14846);
and U17354 (N_17354,N_13356,N_14641);
and U17355 (N_17355,N_12152,N_12483);
and U17356 (N_17356,N_14854,N_11456);
or U17357 (N_17357,N_13213,N_12430);
nor U17358 (N_17358,N_11853,N_10072);
nor U17359 (N_17359,N_13755,N_13600);
nor U17360 (N_17360,N_14975,N_14857);
and U17361 (N_17361,N_10555,N_13074);
or U17362 (N_17362,N_11066,N_10542);
nand U17363 (N_17363,N_14065,N_10729);
nor U17364 (N_17364,N_12474,N_12874);
nor U17365 (N_17365,N_12364,N_11217);
or U17366 (N_17366,N_11001,N_14008);
nand U17367 (N_17367,N_12285,N_13962);
and U17368 (N_17368,N_10616,N_10737);
and U17369 (N_17369,N_14828,N_10599);
or U17370 (N_17370,N_14904,N_10093);
and U17371 (N_17371,N_10225,N_10439);
and U17372 (N_17372,N_13512,N_12355);
nand U17373 (N_17373,N_10154,N_14221);
nand U17374 (N_17374,N_11732,N_13606);
or U17375 (N_17375,N_11557,N_11670);
or U17376 (N_17376,N_10454,N_13200);
nor U17377 (N_17377,N_10440,N_13492);
nor U17378 (N_17378,N_12257,N_12826);
xnor U17379 (N_17379,N_13361,N_10655);
xnor U17380 (N_17380,N_13140,N_13625);
and U17381 (N_17381,N_14679,N_13216);
nor U17382 (N_17382,N_13435,N_13122);
nor U17383 (N_17383,N_14246,N_11605);
and U17384 (N_17384,N_14910,N_13677);
nor U17385 (N_17385,N_10686,N_11751);
nand U17386 (N_17386,N_12200,N_11259);
nand U17387 (N_17387,N_13397,N_13054);
nand U17388 (N_17388,N_14261,N_10386);
and U17389 (N_17389,N_14044,N_11468);
nor U17390 (N_17390,N_14571,N_10483);
or U17391 (N_17391,N_11426,N_12727);
nand U17392 (N_17392,N_13539,N_12934);
or U17393 (N_17393,N_10017,N_10550);
or U17394 (N_17394,N_11652,N_13830);
and U17395 (N_17395,N_13838,N_10286);
nand U17396 (N_17396,N_12273,N_14687);
nand U17397 (N_17397,N_10918,N_13656);
or U17398 (N_17398,N_11058,N_10221);
and U17399 (N_17399,N_12057,N_14033);
nor U17400 (N_17400,N_12958,N_12900);
nor U17401 (N_17401,N_11863,N_10692);
nand U17402 (N_17402,N_10032,N_12177);
nand U17403 (N_17403,N_12834,N_12333);
nor U17404 (N_17404,N_10536,N_13292);
or U17405 (N_17405,N_12043,N_13365);
and U17406 (N_17406,N_12563,N_12634);
and U17407 (N_17407,N_12991,N_10391);
or U17408 (N_17408,N_10277,N_10234);
and U17409 (N_17409,N_10681,N_11518);
nor U17410 (N_17410,N_14316,N_12218);
or U17411 (N_17411,N_10528,N_14493);
nor U17412 (N_17412,N_11952,N_14576);
xnor U17413 (N_17413,N_11494,N_14933);
or U17414 (N_17414,N_10381,N_14633);
nor U17415 (N_17415,N_13026,N_13685);
or U17416 (N_17416,N_11675,N_10563);
nor U17417 (N_17417,N_11895,N_13121);
nor U17418 (N_17418,N_10876,N_13136);
nand U17419 (N_17419,N_12296,N_14809);
and U17420 (N_17420,N_14666,N_13156);
nor U17421 (N_17421,N_14126,N_10785);
nand U17422 (N_17422,N_10999,N_12240);
or U17423 (N_17423,N_12574,N_10255);
nand U17424 (N_17424,N_11787,N_10153);
and U17425 (N_17425,N_13519,N_12264);
nor U17426 (N_17426,N_10656,N_13028);
or U17427 (N_17427,N_12128,N_13723);
nand U17428 (N_17428,N_12564,N_13842);
or U17429 (N_17429,N_10016,N_11743);
or U17430 (N_17430,N_10468,N_11846);
and U17431 (N_17431,N_10533,N_14944);
and U17432 (N_17432,N_14179,N_11715);
nor U17433 (N_17433,N_12661,N_14064);
or U17434 (N_17434,N_11956,N_10888);
nand U17435 (N_17435,N_12136,N_11503);
nand U17436 (N_17436,N_13378,N_13426);
nand U17437 (N_17437,N_11200,N_13810);
nand U17438 (N_17438,N_13617,N_12406);
or U17439 (N_17439,N_11222,N_10461);
nand U17440 (N_17440,N_11486,N_14213);
and U17441 (N_17441,N_10614,N_10580);
and U17442 (N_17442,N_12659,N_12261);
or U17443 (N_17443,N_12915,N_10518);
and U17444 (N_17444,N_12204,N_10341);
nand U17445 (N_17445,N_12101,N_11175);
and U17446 (N_17446,N_12207,N_12254);
nor U17447 (N_17447,N_13648,N_10477);
nand U17448 (N_17448,N_10592,N_13455);
nand U17449 (N_17449,N_12114,N_14048);
nor U17450 (N_17450,N_13132,N_13401);
nand U17451 (N_17451,N_12275,N_13433);
nor U17452 (N_17452,N_13081,N_12456);
nor U17453 (N_17453,N_14175,N_13576);
and U17454 (N_17454,N_14925,N_10484);
nand U17455 (N_17455,N_14517,N_12724);
and U17456 (N_17456,N_11400,N_10636);
or U17457 (N_17457,N_10061,N_13042);
nand U17458 (N_17458,N_14400,N_10977);
nand U17459 (N_17459,N_13851,N_11246);
nand U17460 (N_17460,N_10657,N_11933);
nand U17461 (N_17461,N_12033,N_10651);
and U17462 (N_17462,N_14747,N_10598);
nand U17463 (N_17463,N_14062,N_12711);
and U17464 (N_17464,N_12251,N_14929);
nand U17465 (N_17465,N_12773,N_14303);
nand U17466 (N_17466,N_12084,N_11332);
xor U17467 (N_17467,N_14420,N_14557);
or U17468 (N_17468,N_10293,N_10612);
nor U17469 (N_17469,N_11971,N_14467);
nor U17470 (N_17470,N_11713,N_10425);
nand U17471 (N_17471,N_13070,N_13075);
or U17472 (N_17472,N_13211,N_12615);
nand U17473 (N_17473,N_10116,N_13787);
nor U17474 (N_17474,N_12324,N_11502);
nor U17475 (N_17475,N_13254,N_14220);
or U17476 (N_17476,N_11184,N_12061);
nor U17477 (N_17477,N_14159,N_12157);
or U17478 (N_17478,N_11375,N_14109);
and U17479 (N_17479,N_14690,N_10814);
or U17480 (N_17480,N_13343,N_10471);
and U17481 (N_17481,N_12088,N_10945);
or U17482 (N_17482,N_12754,N_10993);
nor U17483 (N_17483,N_10438,N_14442);
and U17484 (N_17484,N_11091,N_13002);
nor U17485 (N_17485,N_11234,N_10459);
nor U17486 (N_17486,N_13678,N_11756);
nor U17487 (N_17487,N_12359,N_12371);
nor U17488 (N_17488,N_11408,N_14129);
nor U17489 (N_17489,N_10726,N_12405);
or U17490 (N_17490,N_14755,N_12654);
and U17491 (N_17491,N_10929,N_12489);
or U17492 (N_17492,N_12168,N_14323);
nor U17493 (N_17493,N_10245,N_10089);
and U17494 (N_17494,N_13601,N_12671);
and U17495 (N_17495,N_11492,N_11765);
nand U17496 (N_17496,N_12029,N_14974);
or U17497 (N_17497,N_10581,N_11788);
and U17498 (N_17498,N_12199,N_13631);
nor U17499 (N_17499,N_13770,N_14001);
and U17500 (N_17500,N_10200,N_12086);
nor U17501 (N_17501,N_14940,N_14600);
xor U17502 (N_17502,N_13205,N_14473);
nor U17503 (N_17503,N_13325,N_10886);
nand U17504 (N_17504,N_13861,N_13743);
nor U17505 (N_17505,N_11175,N_11915);
nor U17506 (N_17506,N_12982,N_12637);
or U17507 (N_17507,N_13915,N_11391);
nor U17508 (N_17508,N_13921,N_10264);
nor U17509 (N_17509,N_13550,N_10847);
and U17510 (N_17510,N_11094,N_12554);
nand U17511 (N_17511,N_11405,N_12474);
or U17512 (N_17512,N_11838,N_13577);
nand U17513 (N_17513,N_12739,N_10772);
nor U17514 (N_17514,N_14004,N_10188);
nand U17515 (N_17515,N_14406,N_14640);
and U17516 (N_17516,N_11521,N_11656);
or U17517 (N_17517,N_14449,N_11407);
and U17518 (N_17518,N_11453,N_10562);
nor U17519 (N_17519,N_11412,N_12726);
nand U17520 (N_17520,N_13251,N_11431);
nor U17521 (N_17521,N_14900,N_12231);
and U17522 (N_17522,N_14239,N_12622);
and U17523 (N_17523,N_12809,N_13869);
nor U17524 (N_17524,N_14790,N_14036);
or U17525 (N_17525,N_14893,N_14191);
or U17526 (N_17526,N_11090,N_10285);
xor U17527 (N_17527,N_13731,N_12274);
nor U17528 (N_17528,N_10281,N_10792);
nand U17529 (N_17529,N_14196,N_10573);
and U17530 (N_17530,N_13962,N_13888);
xor U17531 (N_17531,N_10114,N_13119);
and U17532 (N_17532,N_14178,N_11480);
nand U17533 (N_17533,N_13483,N_12598);
and U17534 (N_17534,N_10248,N_12892);
nor U17535 (N_17535,N_12418,N_13012);
nor U17536 (N_17536,N_12059,N_13276);
nand U17537 (N_17537,N_13742,N_10903);
nand U17538 (N_17538,N_14427,N_10167);
and U17539 (N_17539,N_11906,N_12161);
nor U17540 (N_17540,N_13579,N_13529);
and U17541 (N_17541,N_10744,N_13252);
nand U17542 (N_17542,N_13849,N_10522);
nand U17543 (N_17543,N_10569,N_14022);
and U17544 (N_17544,N_11868,N_12840);
nor U17545 (N_17545,N_14566,N_11399);
and U17546 (N_17546,N_12712,N_12139);
or U17547 (N_17547,N_12763,N_12537);
and U17548 (N_17548,N_12623,N_12397);
nor U17549 (N_17549,N_14010,N_14474);
and U17550 (N_17550,N_13825,N_14343);
nor U17551 (N_17551,N_10202,N_11630);
and U17552 (N_17552,N_13199,N_11536);
or U17553 (N_17553,N_13646,N_12586);
nor U17554 (N_17554,N_11234,N_14963);
and U17555 (N_17555,N_13370,N_14772);
xnor U17556 (N_17556,N_11597,N_13911);
and U17557 (N_17557,N_12323,N_10716);
and U17558 (N_17558,N_12471,N_12523);
and U17559 (N_17559,N_13285,N_14339);
nor U17560 (N_17560,N_10484,N_13750);
nor U17561 (N_17561,N_12240,N_11327);
and U17562 (N_17562,N_10264,N_12357);
and U17563 (N_17563,N_13766,N_13466);
nor U17564 (N_17564,N_13732,N_10814);
nor U17565 (N_17565,N_12365,N_11786);
nor U17566 (N_17566,N_11286,N_14623);
nor U17567 (N_17567,N_12482,N_13754);
nor U17568 (N_17568,N_12132,N_14570);
or U17569 (N_17569,N_13874,N_13493);
or U17570 (N_17570,N_13422,N_13078);
nor U17571 (N_17571,N_14767,N_14864);
nor U17572 (N_17572,N_13093,N_10440);
nand U17573 (N_17573,N_11565,N_10803);
nor U17574 (N_17574,N_12384,N_10896);
and U17575 (N_17575,N_12976,N_11503);
or U17576 (N_17576,N_10319,N_14187);
nor U17577 (N_17577,N_13502,N_13973);
nand U17578 (N_17578,N_13380,N_11781);
or U17579 (N_17579,N_14387,N_13085);
nand U17580 (N_17580,N_12105,N_10342);
nand U17581 (N_17581,N_10116,N_11743);
and U17582 (N_17582,N_13687,N_14097);
nand U17583 (N_17583,N_12042,N_12603);
or U17584 (N_17584,N_13910,N_13196);
nand U17585 (N_17585,N_14454,N_11012);
or U17586 (N_17586,N_11672,N_11730);
xnor U17587 (N_17587,N_12549,N_14147);
or U17588 (N_17588,N_13663,N_13320);
nand U17589 (N_17589,N_10922,N_11231);
and U17590 (N_17590,N_13459,N_10772);
or U17591 (N_17591,N_13641,N_10973);
and U17592 (N_17592,N_10292,N_11622);
or U17593 (N_17593,N_11200,N_11744);
nor U17594 (N_17594,N_14163,N_10968);
or U17595 (N_17595,N_13969,N_14758);
nand U17596 (N_17596,N_10797,N_14315);
nand U17597 (N_17597,N_12052,N_13522);
nor U17598 (N_17598,N_12141,N_10336);
nor U17599 (N_17599,N_14622,N_14861);
nor U17600 (N_17600,N_10014,N_10668);
nor U17601 (N_17601,N_12782,N_11935);
or U17602 (N_17602,N_10834,N_13482);
and U17603 (N_17603,N_12380,N_13272);
or U17604 (N_17604,N_12148,N_12674);
nor U17605 (N_17605,N_13570,N_10435);
nor U17606 (N_17606,N_14806,N_14195);
nand U17607 (N_17607,N_14596,N_10653);
or U17608 (N_17608,N_10201,N_10965);
or U17609 (N_17609,N_11344,N_12495);
nand U17610 (N_17610,N_12959,N_13296);
or U17611 (N_17611,N_13634,N_11435);
xor U17612 (N_17612,N_12612,N_12124);
nor U17613 (N_17613,N_11762,N_14631);
nand U17614 (N_17614,N_13348,N_14016);
nand U17615 (N_17615,N_10444,N_13143);
nand U17616 (N_17616,N_10733,N_11734);
or U17617 (N_17617,N_13579,N_11207);
and U17618 (N_17618,N_14767,N_14634);
nor U17619 (N_17619,N_12757,N_12237);
or U17620 (N_17620,N_12054,N_10986);
and U17621 (N_17621,N_14289,N_10506);
nor U17622 (N_17622,N_12588,N_13942);
nand U17623 (N_17623,N_12395,N_10706);
and U17624 (N_17624,N_14072,N_13333);
nor U17625 (N_17625,N_14550,N_14410);
and U17626 (N_17626,N_13191,N_12391);
nand U17627 (N_17627,N_12380,N_13970);
nand U17628 (N_17628,N_11847,N_11461);
nor U17629 (N_17629,N_11417,N_13340);
and U17630 (N_17630,N_12161,N_11839);
nor U17631 (N_17631,N_10124,N_10239);
and U17632 (N_17632,N_14494,N_10072);
xor U17633 (N_17633,N_13239,N_10595);
nand U17634 (N_17634,N_11948,N_10741);
nor U17635 (N_17635,N_10006,N_14862);
nand U17636 (N_17636,N_12887,N_14519);
nand U17637 (N_17637,N_12803,N_10712);
nor U17638 (N_17638,N_10800,N_14950);
nor U17639 (N_17639,N_12227,N_11946);
and U17640 (N_17640,N_10113,N_13796);
or U17641 (N_17641,N_10625,N_10482);
nand U17642 (N_17642,N_14633,N_14112);
nand U17643 (N_17643,N_12572,N_14684);
nor U17644 (N_17644,N_13516,N_12566);
or U17645 (N_17645,N_10371,N_11197);
nor U17646 (N_17646,N_11636,N_12809);
and U17647 (N_17647,N_13599,N_10225);
nor U17648 (N_17648,N_11030,N_10180);
and U17649 (N_17649,N_12171,N_12270);
or U17650 (N_17650,N_10015,N_14441);
or U17651 (N_17651,N_11589,N_10528);
and U17652 (N_17652,N_10602,N_10999);
nor U17653 (N_17653,N_14035,N_14911);
or U17654 (N_17654,N_14849,N_13290);
xor U17655 (N_17655,N_12058,N_10864);
nand U17656 (N_17656,N_14907,N_11415);
nor U17657 (N_17657,N_14135,N_14646);
nand U17658 (N_17658,N_10432,N_13936);
nor U17659 (N_17659,N_11624,N_13737);
and U17660 (N_17660,N_10602,N_10356);
nand U17661 (N_17661,N_11116,N_10607);
or U17662 (N_17662,N_10775,N_11332);
or U17663 (N_17663,N_10902,N_10918);
and U17664 (N_17664,N_12542,N_10768);
nand U17665 (N_17665,N_13834,N_13987);
and U17666 (N_17666,N_10111,N_14120);
and U17667 (N_17667,N_14065,N_13206);
nor U17668 (N_17668,N_10319,N_10370);
nand U17669 (N_17669,N_11978,N_12828);
nor U17670 (N_17670,N_12987,N_14141);
nand U17671 (N_17671,N_11469,N_13487);
nand U17672 (N_17672,N_14214,N_13859);
or U17673 (N_17673,N_14448,N_14166);
xor U17674 (N_17674,N_13647,N_10187);
and U17675 (N_17675,N_10804,N_10211);
nand U17676 (N_17676,N_14160,N_12039);
or U17677 (N_17677,N_14598,N_14030);
or U17678 (N_17678,N_10335,N_13125);
or U17679 (N_17679,N_11597,N_10459);
and U17680 (N_17680,N_13057,N_10216);
nor U17681 (N_17681,N_13224,N_12444);
nor U17682 (N_17682,N_11835,N_11686);
nand U17683 (N_17683,N_12306,N_10862);
or U17684 (N_17684,N_11425,N_14604);
nand U17685 (N_17685,N_12388,N_13314);
nand U17686 (N_17686,N_12204,N_14657);
nor U17687 (N_17687,N_14124,N_12573);
nand U17688 (N_17688,N_13943,N_11294);
nor U17689 (N_17689,N_11347,N_13126);
nor U17690 (N_17690,N_13269,N_13065);
nand U17691 (N_17691,N_14018,N_12241);
and U17692 (N_17692,N_12953,N_10850);
or U17693 (N_17693,N_10185,N_12307);
or U17694 (N_17694,N_11013,N_13004);
nand U17695 (N_17695,N_12022,N_11486);
and U17696 (N_17696,N_13769,N_11863);
or U17697 (N_17697,N_12523,N_13980);
nor U17698 (N_17698,N_12414,N_13397);
nand U17699 (N_17699,N_14108,N_12091);
nor U17700 (N_17700,N_10660,N_14825);
nand U17701 (N_17701,N_11442,N_12973);
nor U17702 (N_17702,N_13251,N_11747);
nand U17703 (N_17703,N_13483,N_11698);
nand U17704 (N_17704,N_11420,N_13124);
or U17705 (N_17705,N_12532,N_11546);
nor U17706 (N_17706,N_13456,N_10897);
or U17707 (N_17707,N_11934,N_12965);
nand U17708 (N_17708,N_10509,N_13352);
or U17709 (N_17709,N_13786,N_10342);
nor U17710 (N_17710,N_11994,N_10178);
nor U17711 (N_17711,N_10637,N_11528);
and U17712 (N_17712,N_14274,N_11871);
or U17713 (N_17713,N_10008,N_13709);
nand U17714 (N_17714,N_10618,N_10229);
nand U17715 (N_17715,N_13168,N_12368);
nor U17716 (N_17716,N_12773,N_12707);
or U17717 (N_17717,N_12862,N_14450);
and U17718 (N_17718,N_12481,N_13714);
nor U17719 (N_17719,N_13835,N_11174);
nor U17720 (N_17720,N_13258,N_14495);
and U17721 (N_17721,N_12130,N_14427);
or U17722 (N_17722,N_10939,N_11456);
and U17723 (N_17723,N_11120,N_11420);
nand U17724 (N_17724,N_10873,N_14993);
and U17725 (N_17725,N_13700,N_14809);
xnor U17726 (N_17726,N_13916,N_10674);
and U17727 (N_17727,N_10765,N_14859);
nor U17728 (N_17728,N_12619,N_13704);
nor U17729 (N_17729,N_12165,N_13014);
nor U17730 (N_17730,N_11531,N_12038);
or U17731 (N_17731,N_11428,N_14422);
nor U17732 (N_17732,N_14757,N_11043);
nand U17733 (N_17733,N_11672,N_11252);
nor U17734 (N_17734,N_14541,N_14842);
nand U17735 (N_17735,N_11583,N_14983);
nor U17736 (N_17736,N_13764,N_12364);
nor U17737 (N_17737,N_13695,N_11678);
nand U17738 (N_17738,N_11694,N_12597);
and U17739 (N_17739,N_11911,N_14138);
nor U17740 (N_17740,N_11166,N_13614);
nor U17741 (N_17741,N_14777,N_14792);
and U17742 (N_17742,N_14285,N_11656);
or U17743 (N_17743,N_12133,N_14380);
nand U17744 (N_17744,N_10899,N_13360);
nand U17745 (N_17745,N_13870,N_13047);
and U17746 (N_17746,N_10477,N_14266);
nand U17747 (N_17747,N_10415,N_11592);
or U17748 (N_17748,N_14577,N_14485);
nand U17749 (N_17749,N_12554,N_12219);
nor U17750 (N_17750,N_12051,N_13877);
and U17751 (N_17751,N_10117,N_13859);
nand U17752 (N_17752,N_11691,N_13572);
nand U17753 (N_17753,N_14303,N_14434);
nand U17754 (N_17754,N_13066,N_14659);
nand U17755 (N_17755,N_14311,N_10154);
nand U17756 (N_17756,N_13035,N_12119);
nand U17757 (N_17757,N_12187,N_11575);
or U17758 (N_17758,N_12196,N_11908);
or U17759 (N_17759,N_14609,N_14395);
and U17760 (N_17760,N_10236,N_12357);
or U17761 (N_17761,N_14877,N_13589);
nand U17762 (N_17762,N_11518,N_12942);
nand U17763 (N_17763,N_14265,N_14220);
nand U17764 (N_17764,N_14009,N_10462);
nor U17765 (N_17765,N_14877,N_10747);
xor U17766 (N_17766,N_14496,N_12243);
nand U17767 (N_17767,N_14043,N_10994);
nand U17768 (N_17768,N_11035,N_12950);
nand U17769 (N_17769,N_12335,N_12405);
or U17770 (N_17770,N_12955,N_13604);
or U17771 (N_17771,N_14793,N_13989);
nand U17772 (N_17772,N_12847,N_10298);
nand U17773 (N_17773,N_10752,N_12128);
nor U17774 (N_17774,N_13449,N_11229);
nand U17775 (N_17775,N_10248,N_13683);
nand U17776 (N_17776,N_12195,N_14156);
nand U17777 (N_17777,N_11215,N_12980);
and U17778 (N_17778,N_14079,N_12475);
nand U17779 (N_17779,N_11456,N_12084);
or U17780 (N_17780,N_10821,N_13223);
nor U17781 (N_17781,N_11274,N_11990);
or U17782 (N_17782,N_13985,N_11180);
nand U17783 (N_17783,N_12942,N_12554);
or U17784 (N_17784,N_14770,N_11309);
xor U17785 (N_17785,N_12217,N_14479);
nand U17786 (N_17786,N_11801,N_12670);
and U17787 (N_17787,N_12589,N_14663);
nand U17788 (N_17788,N_12051,N_11729);
nand U17789 (N_17789,N_10897,N_14407);
and U17790 (N_17790,N_13731,N_11038);
nor U17791 (N_17791,N_12909,N_13593);
or U17792 (N_17792,N_14626,N_13643);
or U17793 (N_17793,N_13833,N_11440);
nor U17794 (N_17794,N_14011,N_14849);
xnor U17795 (N_17795,N_11873,N_11696);
nand U17796 (N_17796,N_13002,N_11095);
nand U17797 (N_17797,N_14854,N_10066);
or U17798 (N_17798,N_10832,N_12909);
and U17799 (N_17799,N_10115,N_13131);
nand U17800 (N_17800,N_13987,N_12873);
nand U17801 (N_17801,N_14356,N_14527);
or U17802 (N_17802,N_13757,N_10189);
xnor U17803 (N_17803,N_12716,N_10284);
and U17804 (N_17804,N_10870,N_10006);
or U17805 (N_17805,N_12690,N_10474);
nor U17806 (N_17806,N_13708,N_14014);
nor U17807 (N_17807,N_11695,N_11588);
and U17808 (N_17808,N_10902,N_11889);
nand U17809 (N_17809,N_10426,N_10227);
or U17810 (N_17810,N_12914,N_10048);
nand U17811 (N_17811,N_10299,N_12423);
and U17812 (N_17812,N_11601,N_10405);
nor U17813 (N_17813,N_14481,N_14619);
nand U17814 (N_17814,N_11419,N_13556);
nand U17815 (N_17815,N_10549,N_12974);
and U17816 (N_17816,N_13907,N_12822);
nand U17817 (N_17817,N_14216,N_10044);
nor U17818 (N_17818,N_12979,N_14610);
or U17819 (N_17819,N_10509,N_10985);
nor U17820 (N_17820,N_13467,N_12779);
nor U17821 (N_17821,N_14501,N_14386);
or U17822 (N_17822,N_14922,N_14722);
nand U17823 (N_17823,N_10142,N_11500);
and U17824 (N_17824,N_12562,N_12426);
or U17825 (N_17825,N_10511,N_12932);
or U17826 (N_17826,N_13285,N_14469);
xor U17827 (N_17827,N_10266,N_10416);
nor U17828 (N_17828,N_11196,N_10376);
or U17829 (N_17829,N_12289,N_14740);
nand U17830 (N_17830,N_11374,N_10000);
or U17831 (N_17831,N_10627,N_11093);
nand U17832 (N_17832,N_12806,N_13029);
or U17833 (N_17833,N_11412,N_13466);
nand U17834 (N_17834,N_14222,N_10667);
nor U17835 (N_17835,N_10860,N_14281);
and U17836 (N_17836,N_12001,N_12087);
nor U17837 (N_17837,N_13329,N_13526);
nor U17838 (N_17838,N_11088,N_13371);
xor U17839 (N_17839,N_12993,N_10493);
nand U17840 (N_17840,N_11473,N_14839);
nand U17841 (N_17841,N_11281,N_14202);
nor U17842 (N_17842,N_12422,N_13213);
and U17843 (N_17843,N_13579,N_11805);
xor U17844 (N_17844,N_13592,N_14860);
nor U17845 (N_17845,N_13723,N_12475);
and U17846 (N_17846,N_11312,N_12411);
nand U17847 (N_17847,N_14580,N_14577);
and U17848 (N_17848,N_11110,N_14036);
or U17849 (N_17849,N_14697,N_12130);
or U17850 (N_17850,N_11427,N_10377);
or U17851 (N_17851,N_11379,N_13512);
nand U17852 (N_17852,N_13070,N_13670);
nor U17853 (N_17853,N_14452,N_13966);
nand U17854 (N_17854,N_10787,N_13524);
and U17855 (N_17855,N_11187,N_13303);
nor U17856 (N_17856,N_14239,N_13982);
nor U17857 (N_17857,N_10573,N_13586);
xor U17858 (N_17858,N_14065,N_14449);
and U17859 (N_17859,N_12732,N_12461);
and U17860 (N_17860,N_13189,N_14975);
and U17861 (N_17861,N_11628,N_13317);
nor U17862 (N_17862,N_13267,N_13196);
or U17863 (N_17863,N_10308,N_14247);
and U17864 (N_17864,N_10418,N_14683);
nand U17865 (N_17865,N_11428,N_10025);
and U17866 (N_17866,N_13146,N_14168);
nand U17867 (N_17867,N_11042,N_14708);
or U17868 (N_17868,N_10405,N_10320);
nand U17869 (N_17869,N_10510,N_14594);
or U17870 (N_17870,N_13962,N_12435);
nand U17871 (N_17871,N_11812,N_10082);
or U17872 (N_17872,N_12289,N_10114);
or U17873 (N_17873,N_14397,N_11272);
and U17874 (N_17874,N_13178,N_11105);
nand U17875 (N_17875,N_10377,N_10640);
nand U17876 (N_17876,N_11568,N_14374);
and U17877 (N_17877,N_10284,N_10340);
xor U17878 (N_17878,N_10159,N_11860);
nand U17879 (N_17879,N_10779,N_14463);
nor U17880 (N_17880,N_14127,N_13047);
and U17881 (N_17881,N_14814,N_13172);
nand U17882 (N_17882,N_11363,N_10367);
and U17883 (N_17883,N_10558,N_14413);
and U17884 (N_17884,N_12973,N_12716);
nor U17885 (N_17885,N_12989,N_14895);
nor U17886 (N_17886,N_14352,N_12559);
and U17887 (N_17887,N_11992,N_14638);
xor U17888 (N_17888,N_14868,N_14973);
nand U17889 (N_17889,N_12268,N_10995);
or U17890 (N_17890,N_14870,N_13439);
xnor U17891 (N_17891,N_13731,N_14595);
nand U17892 (N_17892,N_11631,N_10082);
and U17893 (N_17893,N_12385,N_10596);
and U17894 (N_17894,N_10189,N_11245);
and U17895 (N_17895,N_14660,N_14881);
and U17896 (N_17896,N_14890,N_13665);
nand U17897 (N_17897,N_13207,N_11266);
and U17898 (N_17898,N_10718,N_14410);
nor U17899 (N_17899,N_13541,N_11874);
or U17900 (N_17900,N_10171,N_14616);
or U17901 (N_17901,N_14059,N_14296);
nor U17902 (N_17902,N_13590,N_12599);
nor U17903 (N_17903,N_14435,N_14744);
nor U17904 (N_17904,N_10356,N_11011);
nor U17905 (N_17905,N_10941,N_11336);
nand U17906 (N_17906,N_13952,N_11202);
nand U17907 (N_17907,N_14260,N_11998);
xor U17908 (N_17908,N_12166,N_12029);
and U17909 (N_17909,N_10427,N_12048);
and U17910 (N_17910,N_10738,N_10533);
or U17911 (N_17911,N_14597,N_13189);
and U17912 (N_17912,N_13498,N_11866);
nand U17913 (N_17913,N_13552,N_11156);
and U17914 (N_17914,N_11044,N_13080);
nor U17915 (N_17915,N_14493,N_11233);
and U17916 (N_17916,N_14175,N_10909);
nor U17917 (N_17917,N_12632,N_13472);
nor U17918 (N_17918,N_10821,N_13838);
nor U17919 (N_17919,N_12505,N_14126);
nand U17920 (N_17920,N_13299,N_12260);
xor U17921 (N_17921,N_14936,N_10085);
or U17922 (N_17922,N_11568,N_14687);
nor U17923 (N_17923,N_12647,N_14772);
and U17924 (N_17924,N_13835,N_13282);
nor U17925 (N_17925,N_13171,N_14234);
or U17926 (N_17926,N_12232,N_12587);
nand U17927 (N_17927,N_10760,N_11097);
nor U17928 (N_17928,N_14942,N_14877);
and U17929 (N_17929,N_13377,N_12216);
nor U17930 (N_17930,N_11202,N_11709);
nand U17931 (N_17931,N_10104,N_12816);
nor U17932 (N_17932,N_12323,N_14282);
and U17933 (N_17933,N_10106,N_13033);
xor U17934 (N_17934,N_13697,N_11061);
nor U17935 (N_17935,N_13894,N_11470);
or U17936 (N_17936,N_12265,N_13250);
nand U17937 (N_17937,N_11374,N_11779);
nand U17938 (N_17938,N_13805,N_12832);
or U17939 (N_17939,N_10524,N_14902);
and U17940 (N_17940,N_12046,N_10520);
or U17941 (N_17941,N_13709,N_11370);
nor U17942 (N_17942,N_13915,N_12178);
or U17943 (N_17943,N_14900,N_12614);
or U17944 (N_17944,N_11279,N_10638);
and U17945 (N_17945,N_12577,N_13464);
and U17946 (N_17946,N_13578,N_14404);
and U17947 (N_17947,N_10537,N_12619);
nand U17948 (N_17948,N_10329,N_14241);
nand U17949 (N_17949,N_13599,N_14217);
nand U17950 (N_17950,N_12740,N_12943);
or U17951 (N_17951,N_14242,N_13059);
or U17952 (N_17952,N_12991,N_11779);
nor U17953 (N_17953,N_11511,N_10870);
nor U17954 (N_17954,N_12411,N_14176);
nor U17955 (N_17955,N_11536,N_10516);
nor U17956 (N_17956,N_14337,N_10056);
or U17957 (N_17957,N_14916,N_13989);
or U17958 (N_17958,N_12283,N_10595);
or U17959 (N_17959,N_10608,N_10523);
and U17960 (N_17960,N_14080,N_14746);
nor U17961 (N_17961,N_10421,N_12972);
and U17962 (N_17962,N_12479,N_11871);
or U17963 (N_17963,N_14958,N_12522);
and U17964 (N_17964,N_13073,N_11812);
or U17965 (N_17965,N_14911,N_11888);
and U17966 (N_17966,N_13734,N_14984);
and U17967 (N_17967,N_10295,N_13035);
nand U17968 (N_17968,N_13291,N_10606);
and U17969 (N_17969,N_11997,N_11069);
nor U17970 (N_17970,N_13650,N_12702);
nor U17971 (N_17971,N_13874,N_12054);
nor U17972 (N_17972,N_13222,N_14579);
nor U17973 (N_17973,N_13059,N_12315);
nor U17974 (N_17974,N_12738,N_12697);
and U17975 (N_17975,N_11851,N_14027);
nand U17976 (N_17976,N_12966,N_12138);
nor U17977 (N_17977,N_12642,N_11505);
and U17978 (N_17978,N_13464,N_13513);
nand U17979 (N_17979,N_13549,N_10636);
nand U17980 (N_17980,N_10631,N_12022);
xnor U17981 (N_17981,N_11566,N_10900);
or U17982 (N_17982,N_12844,N_14295);
nor U17983 (N_17983,N_14844,N_10603);
nand U17984 (N_17984,N_11708,N_12051);
nor U17985 (N_17985,N_13738,N_10213);
nand U17986 (N_17986,N_13748,N_10882);
and U17987 (N_17987,N_11110,N_10682);
nor U17988 (N_17988,N_13901,N_14514);
nor U17989 (N_17989,N_12124,N_11645);
or U17990 (N_17990,N_13411,N_13885);
nor U17991 (N_17991,N_10923,N_13153);
nand U17992 (N_17992,N_12358,N_10921);
or U17993 (N_17993,N_13487,N_12409);
nor U17994 (N_17994,N_14905,N_10507);
nand U17995 (N_17995,N_14416,N_11500);
nand U17996 (N_17996,N_12703,N_10971);
nand U17997 (N_17997,N_11867,N_10448);
nand U17998 (N_17998,N_12926,N_12220);
and U17999 (N_17999,N_13585,N_11700);
nand U18000 (N_18000,N_14732,N_10942);
and U18001 (N_18001,N_13758,N_11552);
or U18002 (N_18002,N_13990,N_12402);
nor U18003 (N_18003,N_12723,N_12244);
and U18004 (N_18004,N_10866,N_14114);
nor U18005 (N_18005,N_12322,N_11571);
nand U18006 (N_18006,N_14050,N_11140);
nor U18007 (N_18007,N_13633,N_10497);
nand U18008 (N_18008,N_12393,N_12437);
or U18009 (N_18009,N_11327,N_12647);
nand U18010 (N_18010,N_10895,N_11785);
nor U18011 (N_18011,N_10717,N_14370);
nor U18012 (N_18012,N_13583,N_11807);
or U18013 (N_18013,N_10452,N_11048);
nor U18014 (N_18014,N_10543,N_14043);
nand U18015 (N_18015,N_14749,N_11750);
nor U18016 (N_18016,N_11123,N_10564);
nor U18017 (N_18017,N_12662,N_13555);
xnor U18018 (N_18018,N_13393,N_14933);
and U18019 (N_18019,N_14906,N_11534);
and U18020 (N_18020,N_10468,N_14932);
or U18021 (N_18021,N_11517,N_10194);
and U18022 (N_18022,N_14271,N_12257);
nor U18023 (N_18023,N_14265,N_10644);
or U18024 (N_18024,N_12408,N_14832);
nor U18025 (N_18025,N_11577,N_14072);
and U18026 (N_18026,N_14539,N_12655);
or U18027 (N_18027,N_12751,N_14122);
and U18028 (N_18028,N_10536,N_14800);
nor U18029 (N_18029,N_14119,N_12865);
nor U18030 (N_18030,N_12105,N_12008);
nand U18031 (N_18031,N_10737,N_13339);
or U18032 (N_18032,N_10431,N_13669);
nor U18033 (N_18033,N_14585,N_13571);
nand U18034 (N_18034,N_11357,N_11018);
nand U18035 (N_18035,N_11570,N_14878);
and U18036 (N_18036,N_10865,N_10228);
and U18037 (N_18037,N_11429,N_12076);
nand U18038 (N_18038,N_14481,N_14273);
and U18039 (N_18039,N_14606,N_14535);
and U18040 (N_18040,N_11377,N_12316);
nand U18041 (N_18041,N_13430,N_13599);
or U18042 (N_18042,N_14137,N_10892);
nand U18043 (N_18043,N_12121,N_11394);
nor U18044 (N_18044,N_13906,N_10468);
nor U18045 (N_18045,N_12892,N_11520);
or U18046 (N_18046,N_14647,N_14895);
or U18047 (N_18047,N_11688,N_11581);
nand U18048 (N_18048,N_12977,N_11927);
nor U18049 (N_18049,N_12518,N_14031);
nor U18050 (N_18050,N_12026,N_13716);
and U18051 (N_18051,N_10714,N_12050);
and U18052 (N_18052,N_10513,N_12948);
nor U18053 (N_18053,N_14866,N_10234);
nor U18054 (N_18054,N_13921,N_14587);
nor U18055 (N_18055,N_13721,N_11652);
or U18056 (N_18056,N_10437,N_12875);
and U18057 (N_18057,N_13193,N_13264);
and U18058 (N_18058,N_11540,N_12173);
nor U18059 (N_18059,N_14139,N_14543);
nor U18060 (N_18060,N_13261,N_10172);
nor U18061 (N_18061,N_11475,N_10829);
nor U18062 (N_18062,N_13922,N_14234);
or U18063 (N_18063,N_13905,N_11037);
or U18064 (N_18064,N_11648,N_12460);
or U18065 (N_18065,N_11279,N_13902);
nor U18066 (N_18066,N_11039,N_12083);
nor U18067 (N_18067,N_12844,N_14257);
nand U18068 (N_18068,N_12713,N_14080);
nand U18069 (N_18069,N_13858,N_11083);
and U18070 (N_18070,N_13923,N_14164);
nand U18071 (N_18071,N_14248,N_14404);
and U18072 (N_18072,N_12536,N_10098);
nor U18073 (N_18073,N_10990,N_10720);
nor U18074 (N_18074,N_12871,N_10648);
or U18075 (N_18075,N_10244,N_13800);
nor U18076 (N_18076,N_10701,N_11915);
nor U18077 (N_18077,N_14675,N_12278);
nand U18078 (N_18078,N_12067,N_11195);
or U18079 (N_18079,N_10187,N_13406);
and U18080 (N_18080,N_13270,N_14797);
nor U18081 (N_18081,N_14987,N_14680);
nor U18082 (N_18082,N_11227,N_13675);
and U18083 (N_18083,N_13856,N_11630);
or U18084 (N_18084,N_12062,N_11322);
and U18085 (N_18085,N_10222,N_10341);
nand U18086 (N_18086,N_11036,N_13268);
and U18087 (N_18087,N_12346,N_12213);
nor U18088 (N_18088,N_10947,N_14310);
and U18089 (N_18089,N_10425,N_14730);
xnor U18090 (N_18090,N_11814,N_11026);
or U18091 (N_18091,N_10845,N_11609);
nor U18092 (N_18092,N_12211,N_14854);
xor U18093 (N_18093,N_14502,N_14398);
nand U18094 (N_18094,N_12841,N_10220);
and U18095 (N_18095,N_11124,N_12085);
nor U18096 (N_18096,N_12788,N_12382);
or U18097 (N_18097,N_13648,N_12843);
or U18098 (N_18098,N_12036,N_12967);
nand U18099 (N_18099,N_11635,N_11347);
or U18100 (N_18100,N_12235,N_13534);
or U18101 (N_18101,N_10250,N_14438);
nand U18102 (N_18102,N_12359,N_14312);
and U18103 (N_18103,N_14262,N_10477);
nand U18104 (N_18104,N_13716,N_11974);
or U18105 (N_18105,N_11347,N_14930);
and U18106 (N_18106,N_10635,N_13817);
and U18107 (N_18107,N_14982,N_10753);
or U18108 (N_18108,N_11605,N_11945);
nand U18109 (N_18109,N_14662,N_11848);
nor U18110 (N_18110,N_10751,N_14138);
or U18111 (N_18111,N_10115,N_11903);
nor U18112 (N_18112,N_10654,N_14917);
and U18113 (N_18113,N_12328,N_10047);
and U18114 (N_18114,N_10885,N_14931);
and U18115 (N_18115,N_11924,N_10622);
xnor U18116 (N_18116,N_14440,N_10499);
or U18117 (N_18117,N_14124,N_11170);
nand U18118 (N_18118,N_11072,N_13365);
nand U18119 (N_18119,N_12598,N_14850);
nor U18120 (N_18120,N_14655,N_12189);
nor U18121 (N_18121,N_13194,N_10141);
nand U18122 (N_18122,N_12807,N_13345);
nor U18123 (N_18123,N_12209,N_12193);
nand U18124 (N_18124,N_10427,N_13788);
nor U18125 (N_18125,N_13133,N_11429);
or U18126 (N_18126,N_14148,N_13537);
nand U18127 (N_18127,N_12677,N_12384);
or U18128 (N_18128,N_10666,N_11828);
or U18129 (N_18129,N_14527,N_11186);
and U18130 (N_18130,N_12088,N_12710);
nand U18131 (N_18131,N_11174,N_13518);
nand U18132 (N_18132,N_14576,N_10476);
or U18133 (N_18133,N_10700,N_11277);
and U18134 (N_18134,N_12763,N_14686);
nor U18135 (N_18135,N_11960,N_14129);
nor U18136 (N_18136,N_10473,N_12569);
nor U18137 (N_18137,N_12495,N_12183);
nand U18138 (N_18138,N_14722,N_13001);
nand U18139 (N_18139,N_12192,N_11969);
nand U18140 (N_18140,N_14774,N_14566);
and U18141 (N_18141,N_10098,N_11557);
nor U18142 (N_18142,N_13574,N_11452);
nor U18143 (N_18143,N_13479,N_12246);
and U18144 (N_18144,N_14400,N_14538);
nand U18145 (N_18145,N_14018,N_14864);
nor U18146 (N_18146,N_12485,N_13496);
and U18147 (N_18147,N_10300,N_14337);
or U18148 (N_18148,N_11604,N_12956);
nor U18149 (N_18149,N_12315,N_13184);
or U18150 (N_18150,N_14563,N_12492);
or U18151 (N_18151,N_13431,N_14587);
or U18152 (N_18152,N_14428,N_10694);
nand U18153 (N_18153,N_11346,N_11881);
nor U18154 (N_18154,N_14400,N_13366);
nor U18155 (N_18155,N_11366,N_12035);
nor U18156 (N_18156,N_13900,N_13381);
and U18157 (N_18157,N_14450,N_13006);
nand U18158 (N_18158,N_14509,N_13317);
nand U18159 (N_18159,N_12764,N_14784);
xnor U18160 (N_18160,N_13303,N_12268);
and U18161 (N_18161,N_13843,N_13457);
nor U18162 (N_18162,N_12531,N_14391);
nor U18163 (N_18163,N_10292,N_13779);
nand U18164 (N_18164,N_13899,N_13431);
and U18165 (N_18165,N_11025,N_13835);
or U18166 (N_18166,N_12726,N_12908);
and U18167 (N_18167,N_12706,N_11197);
nand U18168 (N_18168,N_14110,N_13120);
and U18169 (N_18169,N_10406,N_13514);
xnor U18170 (N_18170,N_10057,N_14077);
or U18171 (N_18171,N_12839,N_14325);
nor U18172 (N_18172,N_11993,N_14009);
or U18173 (N_18173,N_10038,N_11970);
and U18174 (N_18174,N_14944,N_14260);
nor U18175 (N_18175,N_12416,N_10898);
or U18176 (N_18176,N_14148,N_12996);
xnor U18177 (N_18177,N_10423,N_14179);
or U18178 (N_18178,N_11391,N_14030);
and U18179 (N_18179,N_13055,N_13404);
or U18180 (N_18180,N_12180,N_14392);
and U18181 (N_18181,N_12558,N_10090);
and U18182 (N_18182,N_14353,N_13449);
or U18183 (N_18183,N_13834,N_13929);
and U18184 (N_18184,N_13426,N_11365);
nand U18185 (N_18185,N_11941,N_14407);
or U18186 (N_18186,N_13282,N_10261);
nor U18187 (N_18187,N_12635,N_10965);
or U18188 (N_18188,N_13180,N_11134);
or U18189 (N_18189,N_11489,N_14743);
and U18190 (N_18190,N_10126,N_14100);
and U18191 (N_18191,N_11311,N_14727);
nor U18192 (N_18192,N_10989,N_14105);
nor U18193 (N_18193,N_13907,N_12279);
nand U18194 (N_18194,N_14410,N_12915);
nand U18195 (N_18195,N_11072,N_11985);
nor U18196 (N_18196,N_13343,N_10105);
nand U18197 (N_18197,N_11282,N_10982);
nor U18198 (N_18198,N_10212,N_12111);
or U18199 (N_18199,N_14461,N_11299);
xor U18200 (N_18200,N_11885,N_11490);
nand U18201 (N_18201,N_13729,N_10242);
or U18202 (N_18202,N_12683,N_14360);
and U18203 (N_18203,N_12135,N_13123);
or U18204 (N_18204,N_13625,N_14254);
or U18205 (N_18205,N_14461,N_12642);
nand U18206 (N_18206,N_11437,N_11098);
nand U18207 (N_18207,N_10147,N_13034);
nor U18208 (N_18208,N_11587,N_10616);
and U18209 (N_18209,N_12369,N_12917);
or U18210 (N_18210,N_12823,N_12971);
and U18211 (N_18211,N_11185,N_13813);
or U18212 (N_18212,N_14748,N_10935);
xor U18213 (N_18213,N_14854,N_10256);
nor U18214 (N_18214,N_12776,N_11659);
nor U18215 (N_18215,N_14735,N_13841);
nand U18216 (N_18216,N_12985,N_11300);
or U18217 (N_18217,N_12595,N_11098);
nand U18218 (N_18218,N_12515,N_13342);
or U18219 (N_18219,N_12762,N_12144);
nand U18220 (N_18220,N_10838,N_13031);
or U18221 (N_18221,N_13779,N_14684);
nand U18222 (N_18222,N_12860,N_14758);
nand U18223 (N_18223,N_13499,N_14495);
and U18224 (N_18224,N_10374,N_13999);
or U18225 (N_18225,N_14860,N_11607);
nor U18226 (N_18226,N_10763,N_11330);
xor U18227 (N_18227,N_11693,N_12336);
nor U18228 (N_18228,N_10548,N_11351);
or U18229 (N_18229,N_14053,N_12904);
or U18230 (N_18230,N_11899,N_14800);
or U18231 (N_18231,N_11700,N_12759);
or U18232 (N_18232,N_10825,N_12845);
or U18233 (N_18233,N_11050,N_11355);
and U18234 (N_18234,N_14872,N_11552);
nand U18235 (N_18235,N_13700,N_11592);
and U18236 (N_18236,N_10403,N_12696);
nand U18237 (N_18237,N_14692,N_12437);
and U18238 (N_18238,N_12262,N_13256);
and U18239 (N_18239,N_14940,N_14169);
nand U18240 (N_18240,N_12434,N_12570);
nor U18241 (N_18241,N_11841,N_13572);
or U18242 (N_18242,N_12784,N_13716);
and U18243 (N_18243,N_13662,N_12521);
nor U18244 (N_18244,N_12063,N_14261);
nand U18245 (N_18245,N_11493,N_12252);
or U18246 (N_18246,N_14717,N_11256);
and U18247 (N_18247,N_14364,N_11474);
or U18248 (N_18248,N_10183,N_10383);
and U18249 (N_18249,N_12164,N_14990);
xor U18250 (N_18250,N_13495,N_13644);
and U18251 (N_18251,N_14739,N_11856);
or U18252 (N_18252,N_11150,N_14980);
xnor U18253 (N_18253,N_14413,N_10167);
and U18254 (N_18254,N_12092,N_14210);
or U18255 (N_18255,N_10309,N_14721);
and U18256 (N_18256,N_10010,N_10735);
nand U18257 (N_18257,N_12826,N_11751);
nor U18258 (N_18258,N_11755,N_12228);
nor U18259 (N_18259,N_11058,N_13312);
nand U18260 (N_18260,N_10895,N_13533);
nor U18261 (N_18261,N_14929,N_12571);
or U18262 (N_18262,N_11263,N_11255);
or U18263 (N_18263,N_13162,N_11736);
and U18264 (N_18264,N_13243,N_12167);
nor U18265 (N_18265,N_11294,N_11828);
nand U18266 (N_18266,N_13896,N_12708);
nor U18267 (N_18267,N_13594,N_11153);
nor U18268 (N_18268,N_14709,N_12650);
and U18269 (N_18269,N_11331,N_14507);
nand U18270 (N_18270,N_14879,N_10042);
nor U18271 (N_18271,N_11760,N_13112);
and U18272 (N_18272,N_13204,N_14980);
nor U18273 (N_18273,N_11254,N_12507);
and U18274 (N_18274,N_11013,N_11388);
and U18275 (N_18275,N_10187,N_10326);
nand U18276 (N_18276,N_10944,N_10021);
nand U18277 (N_18277,N_14840,N_14112);
and U18278 (N_18278,N_14884,N_11687);
and U18279 (N_18279,N_11127,N_11369);
and U18280 (N_18280,N_11008,N_10761);
or U18281 (N_18281,N_11791,N_14082);
and U18282 (N_18282,N_11991,N_11432);
xnor U18283 (N_18283,N_13118,N_13056);
xor U18284 (N_18284,N_13891,N_10559);
nor U18285 (N_18285,N_13509,N_10238);
and U18286 (N_18286,N_11029,N_10706);
and U18287 (N_18287,N_12199,N_10198);
or U18288 (N_18288,N_10376,N_10657);
and U18289 (N_18289,N_13158,N_12592);
and U18290 (N_18290,N_13928,N_12729);
or U18291 (N_18291,N_11614,N_11090);
nand U18292 (N_18292,N_14446,N_12222);
nor U18293 (N_18293,N_14286,N_13541);
nand U18294 (N_18294,N_10661,N_12369);
or U18295 (N_18295,N_13191,N_13682);
nand U18296 (N_18296,N_12061,N_10527);
and U18297 (N_18297,N_12770,N_13966);
nor U18298 (N_18298,N_12341,N_12285);
xnor U18299 (N_18299,N_14111,N_14555);
nor U18300 (N_18300,N_11871,N_13949);
nand U18301 (N_18301,N_10991,N_11037);
and U18302 (N_18302,N_14308,N_14088);
nor U18303 (N_18303,N_12354,N_10735);
nand U18304 (N_18304,N_12774,N_14659);
or U18305 (N_18305,N_14752,N_11419);
and U18306 (N_18306,N_12272,N_14354);
and U18307 (N_18307,N_14374,N_10802);
and U18308 (N_18308,N_10702,N_11420);
nor U18309 (N_18309,N_13409,N_11352);
and U18310 (N_18310,N_13244,N_11254);
and U18311 (N_18311,N_13312,N_10895);
and U18312 (N_18312,N_13284,N_14620);
or U18313 (N_18313,N_12954,N_11689);
nand U18314 (N_18314,N_13241,N_10788);
and U18315 (N_18315,N_12143,N_13654);
nor U18316 (N_18316,N_12800,N_13655);
nand U18317 (N_18317,N_10069,N_11954);
nand U18318 (N_18318,N_12376,N_12119);
nor U18319 (N_18319,N_12504,N_12430);
and U18320 (N_18320,N_11220,N_11086);
or U18321 (N_18321,N_14323,N_12335);
nand U18322 (N_18322,N_12545,N_14434);
and U18323 (N_18323,N_13589,N_11535);
or U18324 (N_18324,N_11425,N_13469);
or U18325 (N_18325,N_10789,N_14092);
nor U18326 (N_18326,N_10256,N_12417);
nand U18327 (N_18327,N_10412,N_11870);
nand U18328 (N_18328,N_12262,N_12105);
nand U18329 (N_18329,N_13935,N_13754);
nor U18330 (N_18330,N_14333,N_14201);
or U18331 (N_18331,N_13158,N_10688);
and U18332 (N_18332,N_12515,N_13868);
or U18333 (N_18333,N_12016,N_12964);
and U18334 (N_18334,N_10737,N_12939);
and U18335 (N_18335,N_14442,N_14889);
or U18336 (N_18336,N_14167,N_10982);
or U18337 (N_18337,N_10847,N_11987);
nor U18338 (N_18338,N_12550,N_14594);
nor U18339 (N_18339,N_12509,N_10763);
and U18340 (N_18340,N_14548,N_13350);
and U18341 (N_18341,N_12083,N_13497);
nor U18342 (N_18342,N_12913,N_14056);
and U18343 (N_18343,N_14482,N_14965);
or U18344 (N_18344,N_13967,N_12670);
nand U18345 (N_18345,N_13770,N_13551);
nor U18346 (N_18346,N_12373,N_10604);
or U18347 (N_18347,N_11075,N_14346);
nor U18348 (N_18348,N_11449,N_14119);
or U18349 (N_18349,N_13946,N_13658);
nor U18350 (N_18350,N_11122,N_10058);
or U18351 (N_18351,N_14775,N_11543);
or U18352 (N_18352,N_13657,N_10443);
and U18353 (N_18353,N_10657,N_14351);
nor U18354 (N_18354,N_11769,N_12431);
nor U18355 (N_18355,N_10539,N_14921);
and U18356 (N_18356,N_14383,N_13266);
nor U18357 (N_18357,N_10877,N_13557);
or U18358 (N_18358,N_14548,N_12174);
or U18359 (N_18359,N_10173,N_11594);
or U18360 (N_18360,N_10555,N_12957);
and U18361 (N_18361,N_10164,N_14293);
or U18362 (N_18362,N_14233,N_12011);
or U18363 (N_18363,N_14516,N_12824);
nor U18364 (N_18364,N_14872,N_10175);
or U18365 (N_18365,N_14925,N_12005);
nand U18366 (N_18366,N_10267,N_11939);
nand U18367 (N_18367,N_11012,N_10147);
nand U18368 (N_18368,N_10053,N_14518);
nor U18369 (N_18369,N_10188,N_11381);
nand U18370 (N_18370,N_13433,N_14780);
nand U18371 (N_18371,N_13410,N_14042);
or U18372 (N_18372,N_13714,N_10314);
nand U18373 (N_18373,N_12311,N_14082);
nand U18374 (N_18374,N_13292,N_10441);
nand U18375 (N_18375,N_13640,N_13473);
or U18376 (N_18376,N_13332,N_13111);
and U18377 (N_18377,N_11676,N_14873);
nor U18378 (N_18378,N_12308,N_14879);
and U18379 (N_18379,N_12266,N_10270);
or U18380 (N_18380,N_11385,N_11494);
nor U18381 (N_18381,N_14747,N_11325);
nor U18382 (N_18382,N_12619,N_13188);
and U18383 (N_18383,N_10837,N_10875);
nand U18384 (N_18384,N_14363,N_12254);
xor U18385 (N_18385,N_10961,N_14177);
nor U18386 (N_18386,N_12503,N_12712);
and U18387 (N_18387,N_11336,N_12023);
or U18388 (N_18388,N_14448,N_11094);
nor U18389 (N_18389,N_13365,N_13142);
nand U18390 (N_18390,N_10688,N_10141);
and U18391 (N_18391,N_13392,N_10299);
and U18392 (N_18392,N_12430,N_14331);
xnor U18393 (N_18393,N_14030,N_10387);
nor U18394 (N_18394,N_10012,N_11010);
and U18395 (N_18395,N_13878,N_11683);
and U18396 (N_18396,N_13274,N_13999);
or U18397 (N_18397,N_10092,N_13815);
nor U18398 (N_18398,N_12477,N_13085);
xnor U18399 (N_18399,N_12969,N_10812);
nand U18400 (N_18400,N_11814,N_14433);
and U18401 (N_18401,N_13484,N_10602);
nor U18402 (N_18402,N_13316,N_12918);
and U18403 (N_18403,N_13216,N_11155);
nand U18404 (N_18404,N_12886,N_12203);
or U18405 (N_18405,N_13846,N_14320);
nand U18406 (N_18406,N_13598,N_10469);
nand U18407 (N_18407,N_12777,N_12406);
or U18408 (N_18408,N_12343,N_14912);
and U18409 (N_18409,N_13740,N_11066);
or U18410 (N_18410,N_11673,N_10575);
or U18411 (N_18411,N_11941,N_12123);
nor U18412 (N_18412,N_11785,N_11092);
nand U18413 (N_18413,N_14289,N_14146);
nand U18414 (N_18414,N_11855,N_13540);
or U18415 (N_18415,N_12452,N_13621);
or U18416 (N_18416,N_13552,N_13413);
and U18417 (N_18417,N_10274,N_13799);
and U18418 (N_18418,N_14407,N_13397);
and U18419 (N_18419,N_10354,N_14200);
nand U18420 (N_18420,N_12876,N_14095);
nor U18421 (N_18421,N_11985,N_12499);
nand U18422 (N_18422,N_12975,N_11648);
and U18423 (N_18423,N_11363,N_10561);
and U18424 (N_18424,N_10829,N_10675);
nor U18425 (N_18425,N_11803,N_10407);
nand U18426 (N_18426,N_14570,N_14518);
nor U18427 (N_18427,N_11722,N_11575);
and U18428 (N_18428,N_10487,N_12989);
and U18429 (N_18429,N_14593,N_13049);
and U18430 (N_18430,N_14809,N_13263);
nand U18431 (N_18431,N_13284,N_10211);
or U18432 (N_18432,N_14421,N_11757);
or U18433 (N_18433,N_13929,N_11390);
and U18434 (N_18434,N_13841,N_12727);
and U18435 (N_18435,N_11737,N_12670);
or U18436 (N_18436,N_12872,N_10879);
nand U18437 (N_18437,N_11859,N_13030);
or U18438 (N_18438,N_10570,N_13941);
nor U18439 (N_18439,N_14617,N_10871);
and U18440 (N_18440,N_10465,N_13204);
and U18441 (N_18441,N_14641,N_14620);
nor U18442 (N_18442,N_12518,N_11286);
and U18443 (N_18443,N_13159,N_11061);
or U18444 (N_18444,N_12582,N_12541);
nand U18445 (N_18445,N_12121,N_12304);
nor U18446 (N_18446,N_13071,N_13164);
and U18447 (N_18447,N_13208,N_13180);
nor U18448 (N_18448,N_10369,N_14693);
and U18449 (N_18449,N_13086,N_12240);
or U18450 (N_18450,N_13954,N_11799);
and U18451 (N_18451,N_10158,N_10587);
and U18452 (N_18452,N_12053,N_10455);
nand U18453 (N_18453,N_11138,N_12441);
or U18454 (N_18454,N_14764,N_12751);
nand U18455 (N_18455,N_14687,N_10467);
or U18456 (N_18456,N_14530,N_14613);
nor U18457 (N_18457,N_12447,N_14755);
nand U18458 (N_18458,N_13340,N_11992);
and U18459 (N_18459,N_10966,N_13177);
and U18460 (N_18460,N_11130,N_11491);
and U18461 (N_18461,N_11489,N_14641);
or U18462 (N_18462,N_11133,N_14109);
nor U18463 (N_18463,N_10270,N_11868);
nand U18464 (N_18464,N_11799,N_10326);
or U18465 (N_18465,N_10216,N_14590);
nor U18466 (N_18466,N_13130,N_10224);
or U18467 (N_18467,N_12837,N_10182);
or U18468 (N_18468,N_10739,N_12543);
or U18469 (N_18469,N_11399,N_10429);
and U18470 (N_18470,N_10457,N_11511);
nor U18471 (N_18471,N_10761,N_10276);
and U18472 (N_18472,N_14223,N_11850);
or U18473 (N_18473,N_12129,N_10630);
nor U18474 (N_18474,N_12092,N_14449);
and U18475 (N_18475,N_12384,N_11930);
and U18476 (N_18476,N_10192,N_10041);
nor U18477 (N_18477,N_13188,N_10287);
nor U18478 (N_18478,N_11659,N_12265);
nor U18479 (N_18479,N_12014,N_12753);
and U18480 (N_18480,N_13858,N_10391);
and U18481 (N_18481,N_12804,N_13916);
nand U18482 (N_18482,N_13354,N_13096);
nor U18483 (N_18483,N_10625,N_11363);
and U18484 (N_18484,N_10123,N_14620);
or U18485 (N_18485,N_13503,N_11442);
nand U18486 (N_18486,N_14012,N_10807);
or U18487 (N_18487,N_13871,N_12544);
nor U18488 (N_18488,N_10768,N_12238);
or U18489 (N_18489,N_13788,N_11211);
and U18490 (N_18490,N_10140,N_12288);
nand U18491 (N_18491,N_10420,N_11842);
and U18492 (N_18492,N_11167,N_11542);
nand U18493 (N_18493,N_12327,N_10175);
nand U18494 (N_18494,N_10831,N_14786);
or U18495 (N_18495,N_10585,N_13890);
or U18496 (N_18496,N_13179,N_14483);
or U18497 (N_18497,N_13212,N_13666);
and U18498 (N_18498,N_11607,N_11414);
or U18499 (N_18499,N_13365,N_11655);
nand U18500 (N_18500,N_13356,N_13184);
nand U18501 (N_18501,N_11074,N_11919);
nor U18502 (N_18502,N_10096,N_14027);
or U18503 (N_18503,N_14334,N_13298);
and U18504 (N_18504,N_13223,N_12890);
and U18505 (N_18505,N_10074,N_10535);
or U18506 (N_18506,N_13618,N_11261);
nand U18507 (N_18507,N_14303,N_13034);
xnor U18508 (N_18508,N_13297,N_11968);
and U18509 (N_18509,N_13553,N_10776);
and U18510 (N_18510,N_14284,N_11249);
or U18511 (N_18511,N_13456,N_10990);
xor U18512 (N_18512,N_13191,N_14247);
and U18513 (N_18513,N_10024,N_11910);
and U18514 (N_18514,N_12630,N_13134);
or U18515 (N_18515,N_13305,N_14732);
or U18516 (N_18516,N_14908,N_13560);
or U18517 (N_18517,N_13301,N_11832);
or U18518 (N_18518,N_11299,N_12097);
and U18519 (N_18519,N_11141,N_12874);
or U18520 (N_18520,N_11008,N_13037);
or U18521 (N_18521,N_14559,N_12892);
or U18522 (N_18522,N_10628,N_11867);
nand U18523 (N_18523,N_12389,N_11574);
or U18524 (N_18524,N_12088,N_12550);
and U18525 (N_18525,N_10839,N_12690);
nor U18526 (N_18526,N_11539,N_14878);
nor U18527 (N_18527,N_12978,N_10863);
nand U18528 (N_18528,N_10860,N_14230);
nand U18529 (N_18529,N_14803,N_12123);
xor U18530 (N_18530,N_10881,N_13585);
or U18531 (N_18531,N_13044,N_14090);
or U18532 (N_18532,N_12274,N_13222);
nand U18533 (N_18533,N_13092,N_12415);
nor U18534 (N_18534,N_12347,N_11407);
nor U18535 (N_18535,N_13792,N_13238);
or U18536 (N_18536,N_11202,N_12153);
or U18537 (N_18537,N_10199,N_13763);
nand U18538 (N_18538,N_12708,N_13833);
or U18539 (N_18539,N_12415,N_12511);
or U18540 (N_18540,N_12887,N_14131);
and U18541 (N_18541,N_11161,N_11836);
and U18542 (N_18542,N_10660,N_13751);
nand U18543 (N_18543,N_14682,N_12717);
nand U18544 (N_18544,N_10872,N_10730);
or U18545 (N_18545,N_13434,N_12030);
or U18546 (N_18546,N_12486,N_14199);
or U18547 (N_18547,N_14293,N_10884);
nor U18548 (N_18548,N_14028,N_13616);
or U18549 (N_18549,N_11842,N_12225);
nand U18550 (N_18550,N_10260,N_12100);
and U18551 (N_18551,N_13475,N_10923);
xnor U18552 (N_18552,N_13767,N_14721);
or U18553 (N_18553,N_14108,N_14051);
nor U18554 (N_18554,N_10493,N_11440);
nor U18555 (N_18555,N_12367,N_12743);
and U18556 (N_18556,N_10493,N_11661);
and U18557 (N_18557,N_12581,N_14736);
and U18558 (N_18558,N_14223,N_11219);
nor U18559 (N_18559,N_14953,N_10574);
and U18560 (N_18560,N_11655,N_12924);
nor U18561 (N_18561,N_13230,N_14316);
nand U18562 (N_18562,N_10012,N_14635);
nand U18563 (N_18563,N_10594,N_14105);
or U18564 (N_18564,N_12096,N_13340);
nand U18565 (N_18565,N_10771,N_14092);
nand U18566 (N_18566,N_12114,N_10172);
nand U18567 (N_18567,N_11251,N_11623);
nand U18568 (N_18568,N_14450,N_13324);
and U18569 (N_18569,N_13882,N_14013);
nand U18570 (N_18570,N_13369,N_12780);
nor U18571 (N_18571,N_13906,N_10764);
and U18572 (N_18572,N_11629,N_14214);
nand U18573 (N_18573,N_14740,N_11747);
xor U18574 (N_18574,N_13343,N_13287);
nor U18575 (N_18575,N_14253,N_10236);
nand U18576 (N_18576,N_14393,N_10030);
and U18577 (N_18577,N_11760,N_10572);
nor U18578 (N_18578,N_10037,N_12805);
nand U18579 (N_18579,N_13763,N_10953);
or U18580 (N_18580,N_10528,N_10743);
or U18581 (N_18581,N_10968,N_11357);
nand U18582 (N_18582,N_14723,N_12293);
or U18583 (N_18583,N_12079,N_12814);
nor U18584 (N_18584,N_14141,N_14568);
nand U18585 (N_18585,N_11490,N_11636);
nand U18586 (N_18586,N_14106,N_12069);
nand U18587 (N_18587,N_11488,N_10836);
and U18588 (N_18588,N_11179,N_12142);
nor U18589 (N_18589,N_13723,N_13648);
and U18590 (N_18590,N_13816,N_13915);
and U18591 (N_18591,N_14626,N_14684);
nor U18592 (N_18592,N_10384,N_14822);
and U18593 (N_18593,N_14049,N_12538);
nor U18594 (N_18594,N_11744,N_10977);
nor U18595 (N_18595,N_13234,N_13941);
nor U18596 (N_18596,N_14664,N_12688);
nand U18597 (N_18597,N_12714,N_14083);
and U18598 (N_18598,N_10870,N_12254);
nor U18599 (N_18599,N_14542,N_11356);
nand U18600 (N_18600,N_10963,N_11694);
nand U18601 (N_18601,N_11757,N_10251);
nand U18602 (N_18602,N_14336,N_13028);
or U18603 (N_18603,N_12852,N_11085);
or U18604 (N_18604,N_13314,N_10064);
or U18605 (N_18605,N_14376,N_11653);
nor U18606 (N_18606,N_13162,N_14990);
nor U18607 (N_18607,N_11581,N_13664);
nor U18608 (N_18608,N_14548,N_10015);
and U18609 (N_18609,N_12342,N_13631);
or U18610 (N_18610,N_13463,N_11807);
and U18611 (N_18611,N_13902,N_13828);
nor U18612 (N_18612,N_10143,N_13485);
nor U18613 (N_18613,N_11975,N_12679);
nand U18614 (N_18614,N_12111,N_13263);
and U18615 (N_18615,N_10089,N_10356);
nor U18616 (N_18616,N_14053,N_10327);
and U18617 (N_18617,N_13500,N_11845);
or U18618 (N_18618,N_14557,N_14728);
nand U18619 (N_18619,N_11005,N_12172);
nor U18620 (N_18620,N_10668,N_12231);
nor U18621 (N_18621,N_14968,N_10213);
and U18622 (N_18622,N_14778,N_14764);
nand U18623 (N_18623,N_12686,N_12968);
nand U18624 (N_18624,N_14528,N_13268);
nand U18625 (N_18625,N_13291,N_12548);
nor U18626 (N_18626,N_14438,N_10295);
or U18627 (N_18627,N_14140,N_10664);
nor U18628 (N_18628,N_14094,N_11399);
nor U18629 (N_18629,N_14996,N_13284);
nor U18630 (N_18630,N_14041,N_12304);
xnor U18631 (N_18631,N_14713,N_11574);
nor U18632 (N_18632,N_14738,N_12040);
or U18633 (N_18633,N_11649,N_12163);
nand U18634 (N_18634,N_10706,N_13459);
nor U18635 (N_18635,N_14103,N_14381);
or U18636 (N_18636,N_10671,N_10561);
nor U18637 (N_18637,N_13497,N_13345);
nor U18638 (N_18638,N_12113,N_11844);
nor U18639 (N_18639,N_13669,N_13814);
or U18640 (N_18640,N_13312,N_13173);
nand U18641 (N_18641,N_14380,N_11817);
and U18642 (N_18642,N_12019,N_14083);
nand U18643 (N_18643,N_13962,N_10664);
and U18644 (N_18644,N_11184,N_14383);
or U18645 (N_18645,N_10474,N_11543);
and U18646 (N_18646,N_11554,N_14097);
or U18647 (N_18647,N_13397,N_11875);
nor U18648 (N_18648,N_11286,N_12007);
nand U18649 (N_18649,N_10321,N_12069);
or U18650 (N_18650,N_12625,N_10914);
nor U18651 (N_18651,N_12401,N_11316);
and U18652 (N_18652,N_11068,N_14802);
nand U18653 (N_18653,N_13610,N_10663);
or U18654 (N_18654,N_13644,N_13367);
and U18655 (N_18655,N_12864,N_12148);
and U18656 (N_18656,N_13650,N_12830);
nand U18657 (N_18657,N_13191,N_13868);
nor U18658 (N_18658,N_14456,N_14944);
or U18659 (N_18659,N_10185,N_10462);
nor U18660 (N_18660,N_10517,N_11374);
or U18661 (N_18661,N_12731,N_14507);
nand U18662 (N_18662,N_12923,N_11785);
or U18663 (N_18663,N_14159,N_14619);
or U18664 (N_18664,N_14394,N_12881);
or U18665 (N_18665,N_10448,N_13860);
nand U18666 (N_18666,N_10216,N_11381);
and U18667 (N_18667,N_12586,N_13871);
and U18668 (N_18668,N_12614,N_10690);
nor U18669 (N_18669,N_12456,N_14552);
or U18670 (N_18670,N_14365,N_12576);
nor U18671 (N_18671,N_12515,N_12883);
or U18672 (N_18672,N_13385,N_13617);
nor U18673 (N_18673,N_10317,N_10819);
or U18674 (N_18674,N_10699,N_13941);
or U18675 (N_18675,N_14216,N_13429);
and U18676 (N_18676,N_11471,N_13257);
nor U18677 (N_18677,N_13076,N_10599);
nand U18678 (N_18678,N_12929,N_13318);
nand U18679 (N_18679,N_11714,N_11652);
or U18680 (N_18680,N_12428,N_14038);
nand U18681 (N_18681,N_13098,N_14071);
and U18682 (N_18682,N_13155,N_14190);
nand U18683 (N_18683,N_13300,N_10480);
or U18684 (N_18684,N_10810,N_10192);
or U18685 (N_18685,N_14412,N_14257);
and U18686 (N_18686,N_12639,N_11358);
nand U18687 (N_18687,N_10704,N_13197);
and U18688 (N_18688,N_10431,N_10613);
nand U18689 (N_18689,N_12523,N_11107);
and U18690 (N_18690,N_12967,N_10769);
nor U18691 (N_18691,N_14059,N_12262);
or U18692 (N_18692,N_10483,N_13141);
or U18693 (N_18693,N_12940,N_10585);
and U18694 (N_18694,N_10453,N_10341);
nor U18695 (N_18695,N_11221,N_12103);
and U18696 (N_18696,N_11037,N_14494);
or U18697 (N_18697,N_11702,N_14516);
or U18698 (N_18698,N_14398,N_12460);
xor U18699 (N_18699,N_14612,N_10128);
or U18700 (N_18700,N_12130,N_12306);
and U18701 (N_18701,N_13106,N_14099);
nor U18702 (N_18702,N_13723,N_10504);
nor U18703 (N_18703,N_11121,N_14605);
or U18704 (N_18704,N_11452,N_12015);
nor U18705 (N_18705,N_11653,N_10902);
nand U18706 (N_18706,N_12565,N_13653);
and U18707 (N_18707,N_10688,N_14239);
and U18708 (N_18708,N_12583,N_11613);
nand U18709 (N_18709,N_12960,N_12042);
nor U18710 (N_18710,N_10935,N_12334);
or U18711 (N_18711,N_12410,N_12758);
or U18712 (N_18712,N_12943,N_11807);
and U18713 (N_18713,N_10269,N_11978);
nand U18714 (N_18714,N_10996,N_12713);
nand U18715 (N_18715,N_13550,N_10162);
or U18716 (N_18716,N_13295,N_11801);
xor U18717 (N_18717,N_10678,N_11550);
or U18718 (N_18718,N_13649,N_10445);
and U18719 (N_18719,N_12562,N_13457);
nor U18720 (N_18720,N_14798,N_14248);
or U18721 (N_18721,N_13600,N_14423);
nor U18722 (N_18722,N_14909,N_11331);
and U18723 (N_18723,N_13595,N_10365);
nor U18724 (N_18724,N_13412,N_12449);
nor U18725 (N_18725,N_12222,N_13788);
and U18726 (N_18726,N_13152,N_11581);
and U18727 (N_18727,N_14597,N_14251);
and U18728 (N_18728,N_14502,N_12405);
or U18729 (N_18729,N_11209,N_11321);
or U18730 (N_18730,N_10513,N_11128);
nand U18731 (N_18731,N_13210,N_13071);
xnor U18732 (N_18732,N_13406,N_14068);
nand U18733 (N_18733,N_14727,N_11380);
nand U18734 (N_18734,N_11386,N_10370);
nand U18735 (N_18735,N_12213,N_12008);
and U18736 (N_18736,N_10633,N_11839);
and U18737 (N_18737,N_14418,N_14327);
and U18738 (N_18738,N_11768,N_14856);
and U18739 (N_18739,N_13970,N_10402);
nor U18740 (N_18740,N_12444,N_13263);
nor U18741 (N_18741,N_11672,N_13248);
and U18742 (N_18742,N_11206,N_11161);
and U18743 (N_18743,N_12507,N_10017);
and U18744 (N_18744,N_13817,N_14769);
and U18745 (N_18745,N_14048,N_13488);
or U18746 (N_18746,N_13555,N_14752);
or U18747 (N_18747,N_10508,N_10865);
or U18748 (N_18748,N_14008,N_14585);
nand U18749 (N_18749,N_11126,N_12805);
or U18750 (N_18750,N_13303,N_11074);
xnor U18751 (N_18751,N_14741,N_13856);
xnor U18752 (N_18752,N_13703,N_11204);
nand U18753 (N_18753,N_13657,N_14663);
or U18754 (N_18754,N_11322,N_12419);
and U18755 (N_18755,N_11403,N_11911);
and U18756 (N_18756,N_14089,N_12622);
and U18757 (N_18757,N_11840,N_13283);
nand U18758 (N_18758,N_14973,N_10445);
nand U18759 (N_18759,N_13368,N_13169);
and U18760 (N_18760,N_12807,N_11882);
and U18761 (N_18761,N_12289,N_13772);
and U18762 (N_18762,N_12187,N_14391);
and U18763 (N_18763,N_13116,N_10353);
nor U18764 (N_18764,N_13688,N_12488);
and U18765 (N_18765,N_10348,N_14293);
nor U18766 (N_18766,N_12609,N_11460);
or U18767 (N_18767,N_12454,N_14588);
nor U18768 (N_18768,N_14899,N_11502);
and U18769 (N_18769,N_10332,N_11682);
nor U18770 (N_18770,N_11800,N_10495);
or U18771 (N_18771,N_13129,N_14957);
or U18772 (N_18772,N_14333,N_13308);
nand U18773 (N_18773,N_13441,N_11443);
and U18774 (N_18774,N_11862,N_11190);
or U18775 (N_18775,N_12792,N_10613);
and U18776 (N_18776,N_14900,N_12173);
and U18777 (N_18777,N_11154,N_14707);
nand U18778 (N_18778,N_11572,N_14472);
nand U18779 (N_18779,N_10336,N_14830);
and U18780 (N_18780,N_14408,N_10597);
nor U18781 (N_18781,N_14127,N_12921);
nor U18782 (N_18782,N_13812,N_10929);
nand U18783 (N_18783,N_13419,N_13689);
and U18784 (N_18784,N_10509,N_11463);
nand U18785 (N_18785,N_10120,N_14762);
xnor U18786 (N_18786,N_11054,N_14232);
nand U18787 (N_18787,N_10082,N_12195);
and U18788 (N_18788,N_14757,N_14306);
and U18789 (N_18789,N_14862,N_14511);
nor U18790 (N_18790,N_12968,N_11268);
nor U18791 (N_18791,N_14446,N_14443);
nor U18792 (N_18792,N_13556,N_10745);
or U18793 (N_18793,N_11263,N_11128);
and U18794 (N_18794,N_12734,N_14774);
or U18795 (N_18795,N_14873,N_10631);
or U18796 (N_18796,N_14195,N_11037);
and U18797 (N_18797,N_11084,N_10074);
or U18798 (N_18798,N_12786,N_11375);
or U18799 (N_18799,N_11404,N_11243);
or U18800 (N_18800,N_14660,N_11271);
nor U18801 (N_18801,N_14718,N_11450);
nor U18802 (N_18802,N_12494,N_13015);
xor U18803 (N_18803,N_14489,N_10541);
nor U18804 (N_18804,N_12377,N_14747);
nor U18805 (N_18805,N_11596,N_11129);
nand U18806 (N_18806,N_13162,N_12262);
and U18807 (N_18807,N_11574,N_13290);
and U18808 (N_18808,N_13214,N_10202);
nor U18809 (N_18809,N_12009,N_14609);
or U18810 (N_18810,N_13618,N_10366);
and U18811 (N_18811,N_10988,N_13240);
nor U18812 (N_18812,N_11618,N_12620);
or U18813 (N_18813,N_14427,N_10194);
xor U18814 (N_18814,N_13399,N_11708);
or U18815 (N_18815,N_10525,N_12148);
or U18816 (N_18816,N_14289,N_11652);
xor U18817 (N_18817,N_13601,N_12356);
or U18818 (N_18818,N_11280,N_11732);
or U18819 (N_18819,N_10943,N_11035);
nand U18820 (N_18820,N_10195,N_11786);
nand U18821 (N_18821,N_13333,N_12828);
nand U18822 (N_18822,N_11759,N_11173);
nand U18823 (N_18823,N_14317,N_10456);
and U18824 (N_18824,N_12253,N_14686);
nand U18825 (N_18825,N_14945,N_10119);
nor U18826 (N_18826,N_10826,N_13245);
and U18827 (N_18827,N_12121,N_13741);
and U18828 (N_18828,N_13006,N_11615);
nand U18829 (N_18829,N_10946,N_10942);
and U18830 (N_18830,N_14531,N_12718);
nor U18831 (N_18831,N_10739,N_10440);
and U18832 (N_18832,N_10675,N_13757);
and U18833 (N_18833,N_11384,N_13874);
and U18834 (N_18834,N_12795,N_14944);
and U18835 (N_18835,N_14218,N_10169);
or U18836 (N_18836,N_10080,N_10185);
nor U18837 (N_18837,N_10661,N_12687);
nor U18838 (N_18838,N_13816,N_11779);
or U18839 (N_18839,N_12505,N_11553);
nand U18840 (N_18840,N_10473,N_11250);
nor U18841 (N_18841,N_14417,N_14066);
xor U18842 (N_18842,N_12448,N_12214);
nor U18843 (N_18843,N_14788,N_11437);
nor U18844 (N_18844,N_11430,N_10058);
or U18845 (N_18845,N_14700,N_12778);
nor U18846 (N_18846,N_12418,N_11731);
or U18847 (N_18847,N_10160,N_12130);
nor U18848 (N_18848,N_11707,N_11930);
nor U18849 (N_18849,N_13251,N_11204);
xor U18850 (N_18850,N_13278,N_11554);
nand U18851 (N_18851,N_12040,N_11943);
and U18852 (N_18852,N_11212,N_11095);
and U18853 (N_18853,N_11391,N_14025);
and U18854 (N_18854,N_12188,N_10456);
and U18855 (N_18855,N_12877,N_13271);
and U18856 (N_18856,N_13454,N_10137);
and U18857 (N_18857,N_14556,N_11801);
and U18858 (N_18858,N_10421,N_13928);
nor U18859 (N_18859,N_13312,N_14285);
and U18860 (N_18860,N_10522,N_12863);
nand U18861 (N_18861,N_10864,N_11478);
nor U18862 (N_18862,N_11523,N_10955);
nor U18863 (N_18863,N_13730,N_11118);
nor U18864 (N_18864,N_13148,N_14046);
or U18865 (N_18865,N_12276,N_14321);
and U18866 (N_18866,N_14338,N_13821);
xor U18867 (N_18867,N_12714,N_10739);
and U18868 (N_18868,N_10857,N_12603);
nor U18869 (N_18869,N_13299,N_10528);
nor U18870 (N_18870,N_10796,N_10144);
and U18871 (N_18871,N_13372,N_13032);
and U18872 (N_18872,N_10235,N_13933);
and U18873 (N_18873,N_12961,N_13900);
or U18874 (N_18874,N_13457,N_14144);
and U18875 (N_18875,N_14845,N_14069);
or U18876 (N_18876,N_13431,N_12551);
nand U18877 (N_18877,N_12550,N_11162);
nand U18878 (N_18878,N_14484,N_13590);
and U18879 (N_18879,N_10585,N_13192);
nand U18880 (N_18880,N_13031,N_11120);
xor U18881 (N_18881,N_13985,N_11698);
or U18882 (N_18882,N_14711,N_11081);
nor U18883 (N_18883,N_12323,N_10959);
or U18884 (N_18884,N_11115,N_13981);
xnor U18885 (N_18885,N_13338,N_10410);
nand U18886 (N_18886,N_11880,N_12848);
and U18887 (N_18887,N_12116,N_14156);
or U18888 (N_18888,N_11992,N_11815);
or U18889 (N_18889,N_13275,N_10175);
nand U18890 (N_18890,N_13096,N_10948);
and U18891 (N_18891,N_10598,N_11031);
and U18892 (N_18892,N_10158,N_13370);
nand U18893 (N_18893,N_10661,N_12861);
and U18894 (N_18894,N_11630,N_11217);
and U18895 (N_18895,N_11713,N_12951);
nor U18896 (N_18896,N_13066,N_13626);
nand U18897 (N_18897,N_14224,N_10144);
and U18898 (N_18898,N_10435,N_10119);
nand U18899 (N_18899,N_11102,N_14309);
and U18900 (N_18900,N_12301,N_11525);
nand U18901 (N_18901,N_12512,N_10532);
and U18902 (N_18902,N_14732,N_10645);
nor U18903 (N_18903,N_12000,N_14433);
nor U18904 (N_18904,N_13700,N_11436);
nor U18905 (N_18905,N_10799,N_12173);
nor U18906 (N_18906,N_13069,N_12595);
or U18907 (N_18907,N_11969,N_11643);
nand U18908 (N_18908,N_11942,N_14334);
or U18909 (N_18909,N_11870,N_13879);
or U18910 (N_18910,N_14181,N_12768);
nor U18911 (N_18911,N_12222,N_14524);
and U18912 (N_18912,N_14555,N_14128);
nor U18913 (N_18913,N_10864,N_12413);
nor U18914 (N_18914,N_12785,N_11372);
and U18915 (N_18915,N_14712,N_13544);
nand U18916 (N_18916,N_12729,N_13672);
nor U18917 (N_18917,N_10057,N_12587);
nor U18918 (N_18918,N_14943,N_10496);
and U18919 (N_18919,N_11445,N_14210);
or U18920 (N_18920,N_10621,N_14838);
and U18921 (N_18921,N_10200,N_13840);
nand U18922 (N_18922,N_11297,N_13598);
and U18923 (N_18923,N_12669,N_10561);
and U18924 (N_18924,N_13321,N_11367);
nand U18925 (N_18925,N_13422,N_10289);
nor U18926 (N_18926,N_13077,N_13141);
and U18927 (N_18927,N_12155,N_10074);
xor U18928 (N_18928,N_11504,N_14094);
or U18929 (N_18929,N_13792,N_12507);
or U18930 (N_18930,N_14682,N_11185);
and U18931 (N_18931,N_12158,N_10067);
nand U18932 (N_18932,N_13611,N_13413);
or U18933 (N_18933,N_13970,N_12954);
or U18934 (N_18934,N_12941,N_11703);
or U18935 (N_18935,N_14561,N_10949);
xnor U18936 (N_18936,N_14678,N_11112);
nand U18937 (N_18937,N_13266,N_13945);
or U18938 (N_18938,N_11981,N_10005);
nor U18939 (N_18939,N_14618,N_10817);
or U18940 (N_18940,N_12852,N_14158);
nor U18941 (N_18941,N_12709,N_11662);
nor U18942 (N_18942,N_12327,N_10779);
xnor U18943 (N_18943,N_14024,N_13148);
and U18944 (N_18944,N_11879,N_10656);
or U18945 (N_18945,N_14780,N_10274);
and U18946 (N_18946,N_10837,N_10381);
and U18947 (N_18947,N_14955,N_12129);
or U18948 (N_18948,N_13168,N_14436);
or U18949 (N_18949,N_13302,N_12171);
and U18950 (N_18950,N_12178,N_14923);
xnor U18951 (N_18951,N_12935,N_12197);
nor U18952 (N_18952,N_12192,N_11167);
and U18953 (N_18953,N_13573,N_14216);
nand U18954 (N_18954,N_11089,N_13254);
nand U18955 (N_18955,N_14195,N_14134);
nor U18956 (N_18956,N_13310,N_14375);
or U18957 (N_18957,N_11219,N_13954);
xor U18958 (N_18958,N_12551,N_12014);
nor U18959 (N_18959,N_13798,N_12694);
nor U18960 (N_18960,N_13050,N_11696);
or U18961 (N_18961,N_13950,N_11677);
nand U18962 (N_18962,N_14948,N_11019);
and U18963 (N_18963,N_13273,N_11568);
nor U18964 (N_18964,N_12914,N_10397);
or U18965 (N_18965,N_11176,N_13023);
nand U18966 (N_18966,N_11278,N_14321);
nor U18967 (N_18967,N_14038,N_10199);
nand U18968 (N_18968,N_13062,N_12512);
and U18969 (N_18969,N_13949,N_12842);
nand U18970 (N_18970,N_12666,N_11305);
and U18971 (N_18971,N_10913,N_12673);
and U18972 (N_18972,N_10047,N_12452);
nand U18973 (N_18973,N_13017,N_14744);
xnor U18974 (N_18974,N_14159,N_13876);
nand U18975 (N_18975,N_14250,N_10124);
or U18976 (N_18976,N_14091,N_11722);
and U18977 (N_18977,N_10086,N_13574);
or U18978 (N_18978,N_13705,N_14591);
nand U18979 (N_18979,N_12215,N_13721);
and U18980 (N_18980,N_13066,N_11804);
and U18981 (N_18981,N_13048,N_14068);
nand U18982 (N_18982,N_11606,N_10107);
nor U18983 (N_18983,N_12865,N_14756);
and U18984 (N_18984,N_10724,N_10763);
and U18985 (N_18985,N_10527,N_12417);
xor U18986 (N_18986,N_11627,N_11498);
or U18987 (N_18987,N_10469,N_12755);
nor U18988 (N_18988,N_13850,N_14682);
nor U18989 (N_18989,N_14236,N_11835);
nand U18990 (N_18990,N_13806,N_11632);
or U18991 (N_18991,N_13473,N_11142);
and U18992 (N_18992,N_11671,N_13518);
and U18993 (N_18993,N_14212,N_14653);
nand U18994 (N_18994,N_14837,N_14834);
xor U18995 (N_18995,N_14043,N_10152);
nand U18996 (N_18996,N_11394,N_13489);
or U18997 (N_18997,N_13105,N_13485);
nor U18998 (N_18998,N_10642,N_11648);
nand U18999 (N_18999,N_10778,N_10058);
or U19000 (N_19000,N_11346,N_13810);
nor U19001 (N_19001,N_12942,N_13912);
and U19002 (N_19002,N_10168,N_12473);
and U19003 (N_19003,N_14294,N_10298);
nor U19004 (N_19004,N_12996,N_13284);
and U19005 (N_19005,N_10480,N_12377);
nand U19006 (N_19006,N_14317,N_11517);
nand U19007 (N_19007,N_14052,N_10501);
nor U19008 (N_19008,N_14530,N_13183);
nor U19009 (N_19009,N_13375,N_14576);
nor U19010 (N_19010,N_12701,N_13044);
xnor U19011 (N_19011,N_10851,N_14689);
nand U19012 (N_19012,N_11670,N_10859);
and U19013 (N_19013,N_11006,N_12812);
nand U19014 (N_19014,N_14057,N_12143);
nor U19015 (N_19015,N_11225,N_10318);
nand U19016 (N_19016,N_10836,N_12308);
and U19017 (N_19017,N_12876,N_11495);
or U19018 (N_19018,N_12813,N_12337);
or U19019 (N_19019,N_14838,N_12451);
nand U19020 (N_19020,N_13073,N_13498);
or U19021 (N_19021,N_13236,N_13849);
and U19022 (N_19022,N_13660,N_11599);
and U19023 (N_19023,N_12284,N_14954);
or U19024 (N_19024,N_10921,N_10078);
and U19025 (N_19025,N_14784,N_12905);
or U19026 (N_19026,N_13602,N_13989);
nand U19027 (N_19027,N_13955,N_11021);
and U19028 (N_19028,N_14206,N_11560);
and U19029 (N_19029,N_14694,N_10936);
nand U19030 (N_19030,N_13456,N_12978);
or U19031 (N_19031,N_11149,N_14709);
or U19032 (N_19032,N_13483,N_14483);
and U19033 (N_19033,N_10785,N_14842);
nor U19034 (N_19034,N_12655,N_12573);
and U19035 (N_19035,N_12774,N_10001);
xor U19036 (N_19036,N_13254,N_14633);
or U19037 (N_19037,N_11553,N_13443);
or U19038 (N_19038,N_12131,N_13352);
nor U19039 (N_19039,N_11492,N_14385);
nor U19040 (N_19040,N_14325,N_12550);
nand U19041 (N_19041,N_12752,N_12887);
nand U19042 (N_19042,N_10561,N_12892);
nand U19043 (N_19043,N_12969,N_13278);
nor U19044 (N_19044,N_11941,N_13249);
xor U19045 (N_19045,N_12749,N_13081);
nor U19046 (N_19046,N_13987,N_11424);
nand U19047 (N_19047,N_12178,N_13334);
and U19048 (N_19048,N_10930,N_13994);
xnor U19049 (N_19049,N_12808,N_14384);
and U19050 (N_19050,N_13708,N_10563);
nor U19051 (N_19051,N_10838,N_13427);
or U19052 (N_19052,N_12848,N_12868);
or U19053 (N_19053,N_11519,N_12012);
and U19054 (N_19054,N_14614,N_11833);
and U19055 (N_19055,N_14579,N_14708);
or U19056 (N_19056,N_10636,N_10694);
or U19057 (N_19057,N_14513,N_12878);
and U19058 (N_19058,N_11365,N_11355);
nand U19059 (N_19059,N_12238,N_12803);
or U19060 (N_19060,N_14234,N_14081);
or U19061 (N_19061,N_11393,N_14079);
or U19062 (N_19062,N_12270,N_14763);
nor U19063 (N_19063,N_14315,N_12615);
and U19064 (N_19064,N_14639,N_12703);
nor U19065 (N_19065,N_13585,N_10164);
and U19066 (N_19066,N_11493,N_12609);
nor U19067 (N_19067,N_13756,N_11210);
nand U19068 (N_19068,N_12743,N_14591);
and U19069 (N_19069,N_11866,N_12856);
and U19070 (N_19070,N_10672,N_10171);
or U19071 (N_19071,N_12945,N_13321);
and U19072 (N_19072,N_14205,N_10873);
nand U19073 (N_19073,N_12482,N_13470);
nand U19074 (N_19074,N_12458,N_11022);
nor U19075 (N_19075,N_12391,N_12502);
and U19076 (N_19076,N_13633,N_12596);
nor U19077 (N_19077,N_14129,N_10045);
or U19078 (N_19078,N_14161,N_14378);
nand U19079 (N_19079,N_13210,N_10649);
and U19080 (N_19080,N_11386,N_11181);
nor U19081 (N_19081,N_13673,N_13217);
nand U19082 (N_19082,N_14397,N_14988);
nor U19083 (N_19083,N_11836,N_10826);
or U19084 (N_19084,N_10487,N_12963);
or U19085 (N_19085,N_13388,N_14843);
and U19086 (N_19086,N_13498,N_10781);
nor U19087 (N_19087,N_13882,N_12140);
or U19088 (N_19088,N_13956,N_14597);
xor U19089 (N_19089,N_10049,N_14791);
nand U19090 (N_19090,N_12359,N_13657);
or U19091 (N_19091,N_13467,N_14425);
xor U19092 (N_19092,N_10255,N_14138);
and U19093 (N_19093,N_13549,N_14224);
or U19094 (N_19094,N_13659,N_12579);
nand U19095 (N_19095,N_10462,N_11441);
or U19096 (N_19096,N_12529,N_14427);
nand U19097 (N_19097,N_12722,N_10807);
nand U19098 (N_19098,N_10931,N_11694);
nor U19099 (N_19099,N_10960,N_12052);
or U19100 (N_19100,N_11274,N_10858);
nor U19101 (N_19101,N_14765,N_12546);
nand U19102 (N_19102,N_11365,N_10484);
and U19103 (N_19103,N_11218,N_10918);
nand U19104 (N_19104,N_10718,N_10003);
or U19105 (N_19105,N_12199,N_11700);
or U19106 (N_19106,N_14095,N_12131);
nand U19107 (N_19107,N_10994,N_14528);
or U19108 (N_19108,N_13659,N_10175);
nand U19109 (N_19109,N_11717,N_14857);
nand U19110 (N_19110,N_12475,N_14922);
and U19111 (N_19111,N_12579,N_12948);
or U19112 (N_19112,N_11179,N_11963);
nor U19113 (N_19113,N_12302,N_12647);
nor U19114 (N_19114,N_10697,N_14527);
nor U19115 (N_19115,N_13897,N_12115);
or U19116 (N_19116,N_10081,N_14686);
nand U19117 (N_19117,N_14201,N_13489);
or U19118 (N_19118,N_14204,N_12955);
nor U19119 (N_19119,N_13495,N_14114);
and U19120 (N_19120,N_14834,N_14865);
or U19121 (N_19121,N_13328,N_12394);
and U19122 (N_19122,N_13205,N_10181);
nand U19123 (N_19123,N_13313,N_11519);
nand U19124 (N_19124,N_12375,N_12265);
nor U19125 (N_19125,N_11376,N_11413);
nand U19126 (N_19126,N_10635,N_11970);
nand U19127 (N_19127,N_12771,N_12086);
and U19128 (N_19128,N_10947,N_14926);
or U19129 (N_19129,N_11893,N_12753);
nand U19130 (N_19130,N_12580,N_10227);
xnor U19131 (N_19131,N_11447,N_14069);
and U19132 (N_19132,N_14530,N_13065);
nor U19133 (N_19133,N_12621,N_12147);
or U19134 (N_19134,N_10910,N_12137);
nand U19135 (N_19135,N_12260,N_14837);
nor U19136 (N_19136,N_14854,N_14608);
xnor U19137 (N_19137,N_11657,N_14786);
nor U19138 (N_19138,N_10035,N_12307);
nor U19139 (N_19139,N_14097,N_14228);
nor U19140 (N_19140,N_10330,N_13292);
and U19141 (N_19141,N_11975,N_13890);
nand U19142 (N_19142,N_11184,N_14473);
and U19143 (N_19143,N_14459,N_11159);
or U19144 (N_19144,N_13710,N_10728);
or U19145 (N_19145,N_14173,N_14917);
and U19146 (N_19146,N_13305,N_12883);
and U19147 (N_19147,N_13617,N_10409);
nand U19148 (N_19148,N_13110,N_13779);
and U19149 (N_19149,N_11620,N_12376);
nor U19150 (N_19150,N_13237,N_11800);
nand U19151 (N_19151,N_14879,N_14112);
or U19152 (N_19152,N_12323,N_10657);
or U19153 (N_19153,N_10451,N_10571);
and U19154 (N_19154,N_12983,N_14139);
and U19155 (N_19155,N_12528,N_14853);
nor U19156 (N_19156,N_12412,N_10834);
or U19157 (N_19157,N_10351,N_10171);
nand U19158 (N_19158,N_13517,N_11138);
or U19159 (N_19159,N_14539,N_12746);
and U19160 (N_19160,N_10745,N_13139);
and U19161 (N_19161,N_12693,N_10989);
nor U19162 (N_19162,N_14055,N_14073);
or U19163 (N_19163,N_13039,N_11308);
nor U19164 (N_19164,N_14607,N_13907);
and U19165 (N_19165,N_10974,N_10185);
nor U19166 (N_19166,N_11567,N_12125);
nor U19167 (N_19167,N_11212,N_12043);
nand U19168 (N_19168,N_14692,N_12963);
and U19169 (N_19169,N_14313,N_10975);
nor U19170 (N_19170,N_11722,N_12327);
nor U19171 (N_19171,N_12885,N_13375);
and U19172 (N_19172,N_13317,N_11546);
nor U19173 (N_19173,N_11624,N_10567);
nand U19174 (N_19174,N_10022,N_12408);
nor U19175 (N_19175,N_13431,N_14812);
and U19176 (N_19176,N_12863,N_12355);
nor U19177 (N_19177,N_12359,N_11052);
nor U19178 (N_19178,N_13946,N_10555);
nor U19179 (N_19179,N_13903,N_10200);
or U19180 (N_19180,N_11236,N_13329);
nor U19181 (N_19181,N_11529,N_12018);
or U19182 (N_19182,N_14003,N_12547);
or U19183 (N_19183,N_14110,N_14475);
nand U19184 (N_19184,N_13251,N_12446);
nand U19185 (N_19185,N_10758,N_14884);
nand U19186 (N_19186,N_14441,N_11066);
nand U19187 (N_19187,N_11938,N_13097);
and U19188 (N_19188,N_14034,N_14521);
and U19189 (N_19189,N_13646,N_10819);
nand U19190 (N_19190,N_10036,N_12307);
nor U19191 (N_19191,N_13584,N_11586);
nand U19192 (N_19192,N_12183,N_13990);
nand U19193 (N_19193,N_11877,N_10964);
nand U19194 (N_19194,N_11818,N_12237);
nor U19195 (N_19195,N_11158,N_14406);
and U19196 (N_19196,N_13025,N_14670);
or U19197 (N_19197,N_13008,N_11071);
nand U19198 (N_19198,N_11266,N_13070);
nand U19199 (N_19199,N_13896,N_12586);
xnor U19200 (N_19200,N_12697,N_12267);
nand U19201 (N_19201,N_10679,N_13349);
nor U19202 (N_19202,N_11666,N_13205);
and U19203 (N_19203,N_12615,N_13037);
nand U19204 (N_19204,N_11597,N_12808);
or U19205 (N_19205,N_14486,N_11657);
or U19206 (N_19206,N_14814,N_13604);
nand U19207 (N_19207,N_10903,N_12404);
and U19208 (N_19208,N_14542,N_11511);
nor U19209 (N_19209,N_11627,N_12638);
nand U19210 (N_19210,N_10293,N_10745);
or U19211 (N_19211,N_11127,N_10120);
nand U19212 (N_19212,N_10718,N_13365);
nor U19213 (N_19213,N_11112,N_13134);
nand U19214 (N_19214,N_12906,N_13414);
nor U19215 (N_19215,N_12592,N_14549);
nor U19216 (N_19216,N_14584,N_10457);
nor U19217 (N_19217,N_14085,N_11102);
or U19218 (N_19218,N_12415,N_10035);
nand U19219 (N_19219,N_14435,N_13102);
nand U19220 (N_19220,N_11391,N_13466);
or U19221 (N_19221,N_13017,N_10440);
or U19222 (N_19222,N_10996,N_12501);
or U19223 (N_19223,N_12383,N_10721);
or U19224 (N_19224,N_11928,N_12892);
and U19225 (N_19225,N_14267,N_12811);
and U19226 (N_19226,N_12905,N_11211);
and U19227 (N_19227,N_13113,N_13537);
nor U19228 (N_19228,N_10974,N_14627);
and U19229 (N_19229,N_13288,N_11637);
nand U19230 (N_19230,N_10434,N_12108);
and U19231 (N_19231,N_11124,N_11883);
and U19232 (N_19232,N_11155,N_13548);
nor U19233 (N_19233,N_10009,N_11808);
nor U19234 (N_19234,N_14098,N_14971);
nand U19235 (N_19235,N_10541,N_10808);
and U19236 (N_19236,N_11492,N_13070);
nand U19237 (N_19237,N_12037,N_12847);
and U19238 (N_19238,N_11648,N_14589);
nor U19239 (N_19239,N_13421,N_11113);
and U19240 (N_19240,N_14761,N_12100);
nand U19241 (N_19241,N_12871,N_11512);
and U19242 (N_19242,N_13250,N_13244);
and U19243 (N_19243,N_13366,N_10325);
nor U19244 (N_19244,N_13734,N_10080);
and U19245 (N_19245,N_13473,N_14224);
nor U19246 (N_19246,N_11880,N_14274);
or U19247 (N_19247,N_14541,N_14168);
nand U19248 (N_19248,N_10822,N_13904);
or U19249 (N_19249,N_12026,N_13279);
and U19250 (N_19250,N_14106,N_11922);
nor U19251 (N_19251,N_11469,N_13549);
or U19252 (N_19252,N_12376,N_10696);
xnor U19253 (N_19253,N_11042,N_14774);
or U19254 (N_19254,N_14255,N_14861);
nand U19255 (N_19255,N_12613,N_14202);
nand U19256 (N_19256,N_14430,N_14365);
or U19257 (N_19257,N_10720,N_10193);
nor U19258 (N_19258,N_14286,N_11515);
and U19259 (N_19259,N_14234,N_10531);
nor U19260 (N_19260,N_14758,N_10501);
and U19261 (N_19261,N_14975,N_11054);
and U19262 (N_19262,N_11265,N_11971);
nor U19263 (N_19263,N_10556,N_12431);
and U19264 (N_19264,N_12920,N_12968);
and U19265 (N_19265,N_13519,N_14367);
or U19266 (N_19266,N_10225,N_12229);
or U19267 (N_19267,N_12208,N_10860);
nor U19268 (N_19268,N_10546,N_14451);
nand U19269 (N_19269,N_12448,N_14755);
nor U19270 (N_19270,N_10107,N_11451);
nor U19271 (N_19271,N_11927,N_13498);
and U19272 (N_19272,N_13957,N_14709);
nand U19273 (N_19273,N_11988,N_10147);
and U19274 (N_19274,N_11433,N_14800);
or U19275 (N_19275,N_10671,N_11500);
or U19276 (N_19276,N_12859,N_11548);
nand U19277 (N_19277,N_11394,N_11703);
or U19278 (N_19278,N_11022,N_10555);
or U19279 (N_19279,N_14942,N_10805);
or U19280 (N_19280,N_12141,N_13861);
xor U19281 (N_19281,N_14911,N_14552);
nand U19282 (N_19282,N_12129,N_11061);
nor U19283 (N_19283,N_12974,N_13215);
and U19284 (N_19284,N_13423,N_14273);
or U19285 (N_19285,N_12231,N_10897);
or U19286 (N_19286,N_11727,N_13591);
nand U19287 (N_19287,N_12442,N_13198);
and U19288 (N_19288,N_12925,N_13362);
nor U19289 (N_19289,N_14546,N_12007);
and U19290 (N_19290,N_12068,N_12998);
nor U19291 (N_19291,N_11052,N_12701);
and U19292 (N_19292,N_10831,N_13128);
or U19293 (N_19293,N_13686,N_12717);
nand U19294 (N_19294,N_12226,N_12524);
nor U19295 (N_19295,N_10625,N_13156);
nor U19296 (N_19296,N_12830,N_10336);
and U19297 (N_19297,N_13827,N_10921);
or U19298 (N_19298,N_13984,N_10132);
and U19299 (N_19299,N_14143,N_12329);
nand U19300 (N_19300,N_13016,N_12298);
nor U19301 (N_19301,N_10332,N_13040);
nor U19302 (N_19302,N_12624,N_14184);
and U19303 (N_19303,N_11311,N_10473);
and U19304 (N_19304,N_12457,N_10533);
and U19305 (N_19305,N_11648,N_13429);
nand U19306 (N_19306,N_13499,N_13936);
nor U19307 (N_19307,N_12586,N_13255);
nand U19308 (N_19308,N_13058,N_11265);
and U19309 (N_19309,N_13382,N_13514);
or U19310 (N_19310,N_12096,N_14000);
or U19311 (N_19311,N_13222,N_12882);
nor U19312 (N_19312,N_10962,N_12552);
nand U19313 (N_19313,N_10556,N_14772);
nor U19314 (N_19314,N_13562,N_14569);
or U19315 (N_19315,N_13580,N_14997);
nand U19316 (N_19316,N_12759,N_13941);
and U19317 (N_19317,N_13915,N_10555);
nor U19318 (N_19318,N_13101,N_12916);
nor U19319 (N_19319,N_14465,N_11673);
and U19320 (N_19320,N_11696,N_10907);
and U19321 (N_19321,N_10498,N_12224);
and U19322 (N_19322,N_13661,N_11286);
nor U19323 (N_19323,N_10284,N_11019);
nand U19324 (N_19324,N_10486,N_11039);
or U19325 (N_19325,N_11294,N_11607);
nand U19326 (N_19326,N_11317,N_10961);
or U19327 (N_19327,N_14607,N_11766);
nor U19328 (N_19328,N_10237,N_12264);
and U19329 (N_19329,N_14284,N_13097);
or U19330 (N_19330,N_12938,N_12578);
nor U19331 (N_19331,N_13903,N_10155);
and U19332 (N_19332,N_10754,N_10489);
nand U19333 (N_19333,N_14783,N_13098);
nand U19334 (N_19334,N_12580,N_14446);
nor U19335 (N_19335,N_11663,N_10932);
or U19336 (N_19336,N_14420,N_11368);
nor U19337 (N_19337,N_11540,N_10020);
and U19338 (N_19338,N_11456,N_13530);
nor U19339 (N_19339,N_11386,N_12330);
nand U19340 (N_19340,N_10628,N_12147);
nor U19341 (N_19341,N_11205,N_10036);
nor U19342 (N_19342,N_13932,N_11681);
or U19343 (N_19343,N_14879,N_10804);
nor U19344 (N_19344,N_11281,N_11610);
nand U19345 (N_19345,N_12730,N_12508);
and U19346 (N_19346,N_11456,N_10125);
or U19347 (N_19347,N_13363,N_14896);
or U19348 (N_19348,N_12812,N_12862);
nand U19349 (N_19349,N_12166,N_14911);
xnor U19350 (N_19350,N_13618,N_14991);
nor U19351 (N_19351,N_11671,N_11419);
nand U19352 (N_19352,N_12646,N_14908);
and U19353 (N_19353,N_10273,N_12748);
or U19354 (N_19354,N_11568,N_11648);
or U19355 (N_19355,N_11060,N_13396);
nand U19356 (N_19356,N_14555,N_14266);
nand U19357 (N_19357,N_13169,N_14918);
nor U19358 (N_19358,N_11841,N_10456);
nand U19359 (N_19359,N_10120,N_11064);
nand U19360 (N_19360,N_12416,N_10786);
nor U19361 (N_19361,N_11454,N_13590);
and U19362 (N_19362,N_12236,N_14143);
xor U19363 (N_19363,N_13057,N_11597);
xor U19364 (N_19364,N_13346,N_14566);
or U19365 (N_19365,N_11495,N_11393);
nand U19366 (N_19366,N_11972,N_12541);
or U19367 (N_19367,N_12724,N_12857);
and U19368 (N_19368,N_11542,N_13781);
or U19369 (N_19369,N_12229,N_14370);
xnor U19370 (N_19370,N_14563,N_11099);
nand U19371 (N_19371,N_10892,N_13581);
and U19372 (N_19372,N_13290,N_13060);
or U19373 (N_19373,N_11239,N_10679);
and U19374 (N_19374,N_10268,N_12411);
nand U19375 (N_19375,N_14360,N_12890);
nor U19376 (N_19376,N_11955,N_11291);
nor U19377 (N_19377,N_12701,N_11174);
and U19378 (N_19378,N_11153,N_13810);
or U19379 (N_19379,N_14430,N_14978);
or U19380 (N_19380,N_10961,N_12296);
nor U19381 (N_19381,N_14034,N_12254);
nor U19382 (N_19382,N_10105,N_14738);
xnor U19383 (N_19383,N_14487,N_11206);
nand U19384 (N_19384,N_11210,N_14042);
nor U19385 (N_19385,N_11067,N_10885);
or U19386 (N_19386,N_14666,N_12740);
nor U19387 (N_19387,N_10931,N_13309);
or U19388 (N_19388,N_10910,N_10384);
nor U19389 (N_19389,N_11155,N_12401);
or U19390 (N_19390,N_10556,N_12969);
or U19391 (N_19391,N_13894,N_10026);
nor U19392 (N_19392,N_11421,N_11947);
or U19393 (N_19393,N_11218,N_10539);
and U19394 (N_19394,N_13607,N_14367);
or U19395 (N_19395,N_10958,N_14578);
nor U19396 (N_19396,N_13726,N_10551);
or U19397 (N_19397,N_11041,N_13205);
nand U19398 (N_19398,N_12740,N_14720);
nand U19399 (N_19399,N_14388,N_14562);
or U19400 (N_19400,N_14812,N_10377);
nand U19401 (N_19401,N_11627,N_12983);
and U19402 (N_19402,N_13983,N_10892);
nor U19403 (N_19403,N_12824,N_14250);
nand U19404 (N_19404,N_12231,N_11344);
and U19405 (N_19405,N_13665,N_11933);
and U19406 (N_19406,N_13363,N_10759);
nor U19407 (N_19407,N_11896,N_10290);
or U19408 (N_19408,N_12584,N_14177);
or U19409 (N_19409,N_10650,N_13485);
nand U19410 (N_19410,N_10358,N_14158);
nor U19411 (N_19411,N_11360,N_11802);
nor U19412 (N_19412,N_13323,N_12652);
and U19413 (N_19413,N_14010,N_12332);
nand U19414 (N_19414,N_10928,N_13834);
or U19415 (N_19415,N_13581,N_12666);
or U19416 (N_19416,N_10422,N_12522);
nor U19417 (N_19417,N_13138,N_13042);
and U19418 (N_19418,N_11560,N_13069);
or U19419 (N_19419,N_13947,N_13275);
or U19420 (N_19420,N_11452,N_11878);
nor U19421 (N_19421,N_12473,N_12564);
xor U19422 (N_19422,N_12407,N_13685);
or U19423 (N_19423,N_10871,N_14995);
nor U19424 (N_19424,N_14546,N_11222);
and U19425 (N_19425,N_13926,N_11771);
and U19426 (N_19426,N_13235,N_14502);
and U19427 (N_19427,N_12825,N_12521);
nand U19428 (N_19428,N_10534,N_11575);
and U19429 (N_19429,N_10904,N_13259);
and U19430 (N_19430,N_12032,N_14975);
and U19431 (N_19431,N_10725,N_13420);
and U19432 (N_19432,N_12552,N_14765);
nor U19433 (N_19433,N_11169,N_14060);
xnor U19434 (N_19434,N_10366,N_11730);
and U19435 (N_19435,N_14989,N_10601);
nor U19436 (N_19436,N_11595,N_10361);
nor U19437 (N_19437,N_11310,N_10073);
and U19438 (N_19438,N_10762,N_12637);
and U19439 (N_19439,N_13143,N_10693);
or U19440 (N_19440,N_13233,N_14294);
and U19441 (N_19441,N_13543,N_13163);
and U19442 (N_19442,N_14646,N_10746);
nor U19443 (N_19443,N_11235,N_13476);
nand U19444 (N_19444,N_11233,N_14427);
nor U19445 (N_19445,N_12499,N_14655);
and U19446 (N_19446,N_12781,N_13470);
or U19447 (N_19447,N_11135,N_10656);
nand U19448 (N_19448,N_11074,N_10058);
and U19449 (N_19449,N_13957,N_10075);
or U19450 (N_19450,N_10351,N_13273);
and U19451 (N_19451,N_14979,N_12454);
nor U19452 (N_19452,N_14873,N_11675);
and U19453 (N_19453,N_11459,N_14487);
nor U19454 (N_19454,N_12478,N_13996);
nor U19455 (N_19455,N_14739,N_11923);
nand U19456 (N_19456,N_12337,N_11744);
or U19457 (N_19457,N_12160,N_10880);
nand U19458 (N_19458,N_10065,N_11467);
nor U19459 (N_19459,N_11240,N_10633);
nand U19460 (N_19460,N_14375,N_10885);
and U19461 (N_19461,N_13481,N_12219);
nor U19462 (N_19462,N_14529,N_10327);
nor U19463 (N_19463,N_10302,N_13683);
nor U19464 (N_19464,N_14424,N_12742);
nand U19465 (N_19465,N_10154,N_11362);
nor U19466 (N_19466,N_10234,N_10723);
nor U19467 (N_19467,N_13621,N_13516);
and U19468 (N_19468,N_11332,N_14615);
or U19469 (N_19469,N_13868,N_12452);
nand U19470 (N_19470,N_11766,N_13248);
nor U19471 (N_19471,N_10160,N_10130);
and U19472 (N_19472,N_14452,N_12014);
nand U19473 (N_19473,N_11747,N_14485);
nor U19474 (N_19474,N_10077,N_12514);
and U19475 (N_19475,N_13790,N_13101);
nand U19476 (N_19476,N_11154,N_13823);
and U19477 (N_19477,N_14377,N_14835);
or U19478 (N_19478,N_12177,N_10920);
or U19479 (N_19479,N_13026,N_12560);
and U19480 (N_19480,N_14558,N_10549);
nor U19481 (N_19481,N_12904,N_14460);
nand U19482 (N_19482,N_12637,N_12743);
xnor U19483 (N_19483,N_13213,N_14918);
nand U19484 (N_19484,N_10210,N_11838);
nor U19485 (N_19485,N_10459,N_13536);
and U19486 (N_19486,N_13587,N_11313);
nor U19487 (N_19487,N_12803,N_12358);
or U19488 (N_19488,N_13050,N_14814);
nand U19489 (N_19489,N_13038,N_14652);
nor U19490 (N_19490,N_12274,N_13143);
nand U19491 (N_19491,N_11631,N_13256);
xnor U19492 (N_19492,N_12187,N_12591);
nand U19493 (N_19493,N_14667,N_14423);
nand U19494 (N_19494,N_11213,N_14974);
nor U19495 (N_19495,N_13184,N_14076);
nor U19496 (N_19496,N_10674,N_13079);
or U19497 (N_19497,N_12481,N_13098);
nand U19498 (N_19498,N_11413,N_10865);
nand U19499 (N_19499,N_12150,N_11345);
nand U19500 (N_19500,N_13210,N_12367);
and U19501 (N_19501,N_12031,N_10609);
nor U19502 (N_19502,N_10840,N_12382);
nand U19503 (N_19503,N_11619,N_10537);
xor U19504 (N_19504,N_13906,N_11998);
or U19505 (N_19505,N_12029,N_12972);
and U19506 (N_19506,N_11563,N_14443);
or U19507 (N_19507,N_13084,N_14665);
or U19508 (N_19508,N_12039,N_12206);
nor U19509 (N_19509,N_14542,N_10288);
and U19510 (N_19510,N_13290,N_11344);
and U19511 (N_19511,N_11257,N_12151);
nand U19512 (N_19512,N_13386,N_10856);
nand U19513 (N_19513,N_13012,N_14533);
nand U19514 (N_19514,N_13312,N_13961);
and U19515 (N_19515,N_11150,N_14232);
or U19516 (N_19516,N_13831,N_12258);
nor U19517 (N_19517,N_13291,N_12971);
or U19518 (N_19518,N_14206,N_11570);
and U19519 (N_19519,N_14360,N_12526);
or U19520 (N_19520,N_14576,N_13487);
nand U19521 (N_19521,N_13739,N_14849);
or U19522 (N_19522,N_11409,N_14737);
or U19523 (N_19523,N_11906,N_12895);
nor U19524 (N_19524,N_14030,N_12853);
or U19525 (N_19525,N_13432,N_12175);
nand U19526 (N_19526,N_11377,N_13572);
and U19527 (N_19527,N_10932,N_13077);
nor U19528 (N_19528,N_13229,N_12704);
or U19529 (N_19529,N_13164,N_14192);
and U19530 (N_19530,N_10602,N_13465);
and U19531 (N_19531,N_10219,N_13013);
xor U19532 (N_19532,N_14927,N_14430);
nand U19533 (N_19533,N_13714,N_12342);
xor U19534 (N_19534,N_12150,N_12962);
nand U19535 (N_19535,N_11295,N_14891);
or U19536 (N_19536,N_12275,N_11205);
or U19537 (N_19537,N_12643,N_12230);
nor U19538 (N_19538,N_13478,N_13267);
nor U19539 (N_19539,N_11102,N_13599);
or U19540 (N_19540,N_11467,N_10491);
nand U19541 (N_19541,N_14244,N_12764);
nand U19542 (N_19542,N_12288,N_10653);
nand U19543 (N_19543,N_11309,N_11541);
nand U19544 (N_19544,N_13647,N_14832);
nor U19545 (N_19545,N_10251,N_14095);
or U19546 (N_19546,N_10521,N_13128);
or U19547 (N_19547,N_10713,N_10785);
and U19548 (N_19548,N_14240,N_12655);
and U19549 (N_19549,N_10341,N_12948);
nor U19550 (N_19550,N_12601,N_14791);
nand U19551 (N_19551,N_13763,N_11411);
and U19552 (N_19552,N_10601,N_14399);
nor U19553 (N_19553,N_13437,N_12698);
nand U19554 (N_19554,N_13502,N_14324);
nand U19555 (N_19555,N_10123,N_11389);
nor U19556 (N_19556,N_13340,N_11262);
or U19557 (N_19557,N_11502,N_10570);
and U19558 (N_19558,N_14929,N_14353);
or U19559 (N_19559,N_12918,N_14160);
and U19560 (N_19560,N_12038,N_10874);
and U19561 (N_19561,N_14542,N_13111);
nor U19562 (N_19562,N_11739,N_10007);
xnor U19563 (N_19563,N_12559,N_14170);
or U19564 (N_19564,N_13603,N_12735);
or U19565 (N_19565,N_12647,N_11891);
nand U19566 (N_19566,N_12176,N_14652);
nand U19567 (N_19567,N_11050,N_13097);
nor U19568 (N_19568,N_10145,N_14523);
nor U19569 (N_19569,N_11545,N_10361);
nor U19570 (N_19570,N_14901,N_14025);
nand U19571 (N_19571,N_11420,N_13239);
and U19572 (N_19572,N_14466,N_11272);
nor U19573 (N_19573,N_10762,N_11491);
nor U19574 (N_19574,N_10729,N_14919);
nor U19575 (N_19575,N_14220,N_13409);
nand U19576 (N_19576,N_10053,N_13783);
nand U19577 (N_19577,N_13777,N_14111);
or U19578 (N_19578,N_13887,N_13473);
and U19579 (N_19579,N_14411,N_13251);
nand U19580 (N_19580,N_14428,N_11892);
or U19581 (N_19581,N_10035,N_13113);
or U19582 (N_19582,N_10454,N_14269);
and U19583 (N_19583,N_13928,N_13790);
nand U19584 (N_19584,N_10782,N_11768);
or U19585 (N_19585,N_11260,N_10542);
nor U19586 (N_19586,N_11233,N_13401);
or U19587 (N_19587,N_13937,N_13189);
and U19588 (N_19588,N_10849,N_13876);
and U19589 (N_19589,N_11121,N_10569);
or U19590 (N_19590,N_12367,N_14076);
nor U19591 (N_19591,N_12168,N_12056);
and U19592 (N_19592,N_14139,N_13175);
nor U19593 (N_19593,N_12304,N_13608);
nor U19594 (N_19594,N_10648,N_12504);
nor U19595 (N_19595,N_10358,N_13853);
and U19596 (N_19596,N_12158,N_10390);
nor U19597 (N_19597,N_10869,N_14678);
nand U19598 (N_19598,N_11490,N_10810);
and U19599 (N_19599,N_10528,N_11398);
or U19600 (N_19600,N_12527,N_11129);
or U19601 (N_19601,N_13596,N_13312);
and U19602 (N_19602,N_13430,N_10864);
nand U19603 (N_19603,N_10070,N_14603);
and U19604 (N_19604,N_12634,N_10273);
nand U19605 (N_19605,N_13991,N_13291);
and U19606 (N_19606,N_13035,N_14617);
nand U19607 (N_19607,N_11528,N_11564);
and U19608 (N_19608,N_11861,N_11363);
or U19609 (N_19609,N_10064,N_14599);
nand U19610 (N_19610,N_12369,N_10538);
xnor U19611 (N_19611,N_13005,N_11748);
and U19612 (N_19612,N_11751,N_10827);
or U19613 (N_19613,N_14041,N_14823);
or U19614 (N_19614,N_12404,N_12112);
and U19615 (N_19615,N_11057,N_14684);
or U19616 (N_19616,N_14378,N_11720);
nor U19617 (N_19617,N_11897,N_13958);
and U19618 (N_19618,N_14946,N_12829);
nor U19619 (N_19619,N_13924,N_12465);
xnor U19620 (N_19620,N_13610,N_11752);
or U19621 (N_19621,N_12084,N_13804);
nor U19622 (N_19622,N_11242,N_10901);
or U19623 (N_19623,N_13795,N_14952);
nor U19624 (N_19624,N_12912,N_10428);
xor U19625 (N_19625,N_14387,N_10087);
nor U19626 (N_19626,N_12843,N_13608);
and U19627 (N_19627,N_14002,N_10240);
and U19628 (N_19628,N_14365,N_11140);
nand U19629 (N_19629,N_14589,N_12980);
nor U19630 (N_19630,N_10071,N_12917);
nand U19631 (N_19631,N_10647,N_11794);
or U19632 (N_19632,N_14686,N_10125);
nor U19633 (N_19633,N_11158,N_11796);
and U19634 (N_19634,N_12286,N_13703);
nor U19635 (N_19635,N_10457,N_14930);
and U19636 (N_19636,N_14156,N_13340);
and U19637 (N_19637,N_11350,N_10559);
nor U19638 (N_19638,N_14436,N_11310);
nand U19639 (N_19639,N_11555,N_14059);
nand U19640 (N_19640,N_13342,N_14191);
or U19641 (N_19641,N_10810,N_13977);
nand U19642 (N_19642,N_12629,N_12460);
nand U19643 (N_19643,N_10752,N_11463);
or U19644 (N_19644,N_13916,N_14438);
and U19645 (N_19645,N_13233,N_12216);
nor U19646 (N_19646,N_12642,N_10145);
nor U19647 (N_19647,N_14172,N_10555);
or U19648 (N_19648,N_13314,N_10444);
nor U19649 (N_19649,N_13962,N_12222);
nor U19650 (N_19650,N_10610,N_10085);
nand U19651 (N_19651,N_12863,N_10214);
nand U19652 (N_19652,N_12847,N_10731);
and U19653 (N_19653,N_10352,N_11400);
nor U19654 (N_19654,N_12213,N_14028);
or U19655 (N_19655,N_12750,N_14813);
or U19656 (N_19656,N_11904,N_12950);
or U19657 (N_19657,N_13762,N_10628);
nor U19658 (N_19658,N_14967,N_14840);
and U19659 (N_19659,N_10965,N_10250);
nand U19660 (N_19660,N_10172,N_12309);
or U19661 (N_19661,N_11524,N_13003);
or U19662 (N_19662,N_12093,N_11063);
and U19663 (N_19663,N_14602,N_13766);
or U19664 (N_19664,N_14472,N_10533);
nor U19665 (N_19665,N_13428,N_13416);
nand U19666 (N_19666,N_14731,N_12523);
and U19667 (N_19667,N_13741,N_14885);
nand U19668 (N_19668,N_12361,N_12065);
or U19669 (N_19669,N_12456,N_10634);
nor U19670 (N_19670,N_13352,N_10587);
nand U19671 (N_19671,N_13747,N_12864);
and U19672 (N_19672,N_10792,N_10472);
and U19673 (N_19673,N_14294,N_14291);
and U19674 (N_19674,N_14276,N_14460);
nand U19675 (N_19675,N_14319,N_12758);
nand U19676 (N_19676,N_13635,N_10049);
and U19677 (N_19677,N_11088,N_11303);
nor U19678 (N_19678,N_11896,N_14436);
and U19679 (N_19679,N_10985,N_14612);
and U19680 (N_19680,N_10396,N_10707);
and U19681 (N_19681,N_10100,N_10110);
nor U19682 (N_19682,N_13004,N_13046);
nor U19683 (N_19683,N_13614,N_14702);
nor U19684 (N_19684,N_14644,N_10158);
or U19685 (N_19685,N_14438,N_13968);
nor U19686 (N_19686,N_10828,N_11779);
nor U19687 (N_19687,N_11394,N_14456);
and U19688 (N_19688,N_11861,N_14705);
nor U19689 (N_19689,N_13077,N_14518);
nand U19690 (N_19690,N_11243,N_13815);
nor U19691 (N_19691,N_12853,N_12005);
or U19692 (N_19692,N_11162,N_14694);
and U19693 (N_19693,N_11934,N_11707);
or U19694 (N_19694,N_13923,N_13125);
or U19695 (N_19695,N_13565,N_12260);
nand U19696 (N_19696,N_13341,N_11321);
nor U19697 (N_19697,N_13855,N_11017);
and U19698 (N_19698,N_12028,N_11455);
or U19699 (N_19699,N_11648,N_11613);
and U19700 (N_19700,N_13364,N_12727);
nand U19701 (N_19701,N_13907,N_12834);
nor U19702 (N_19702,N_14961,N_10215);
nor U19703 (N_19703,N_11839,N_11321);
or U19704 (N_19704,N_11404,N_12357);
and U19705 (N_19705,N_13647,N_13242);
and U19706 (N_19706,N_10588,N_10423);
nand U19707 (N_19707,N_13095,N_13801);
and U19708 (N_19708,N_13413,N_10839);
nor U19709 (N_19709,N_10170,N_11760);
nor U19710 (N_19710,N_11805,N_10577);
nor U19711 (N_19711,N_11263,N_10094);
nor U19712 (N_19712,N_12114,N_13911);
nand U19713 (N_19713,N_14543,N_11618);
nor U19714 (N_19714,N_10037,N_11436);
nand U19715 (N_19715,N_11503,N_13992);
and U19716 (N_19716,N_10865,N_11365);
or U19717 (N_19717,N_14384,N_14779);
nand U19718 (N_19718,N_13282,N_13442);
nand U19719 (N_19719,N_13774,N_13276);
and U19720 (N_19720,N_14975,N_13451);
or U19721 (N_19721,N_11803,N_10849);
and U19722 (N_19722,N_10651,N_12598);
and U19723 (N_19723,N_12923,N_12253);
or U19724 (N_19724,N_12736,N_13848);
nand U19725 (N_19725,N_13285,N_12060);
nand U19726 (N_19726,N_12089,N_14758);
nor U19727 (N_19727,N_11883,N_13915);
nor U19728 (N_19728,N_13238,N_11413);
nor U19729 (N_19729,N_10134,N_10137);
and U19730 (N_19730,N_13666,N_13349);
or U19731 (N_19731,N_13098,N_11480);
or U19732 (N_19732,N_11974,N_11817);
or U19733 (N_19733,N_10592,N_14297);
nor U19734 (N_19734,N_13255,N_11843);
xor U19735 (N_19735,N_12018,N_14217);
and U19736 (N_19736,N_10239,N_14433);
nor U19737 (N_19737,N_11726,N_14889);
and U19738 (N_19738,N_10155,N_11587);
nor U19739 (N_19739,N_12717,N_12349);
or U19740 (N_19740,N_11682,N_10061);
or U19741 (N_19741,N_13893,N_11559);
and U19742 (N_19742,N_10177,N_11485);
and U19743 (N_19743,N_10668,N_14575);
and U19744 (N_19744,N_13421,N_12912);
or U19745 (N_19745,N_14918,N_13311);
and U19746 (N_19746,N_12772,N_13093);
or U19747 (N_19747,N_12106,N_13929);
or U19748 (N_19748,N_11774,N_14283);
xnor U19749 (N_19749,N_13277,N_14914);
or U19750 (N_19750,N_13428,N_12943);
or U19751 (N_19751,N_10357,N_11189);
nor U19752 (N_19752,N_14017,N_11840);
xnor U19753 (N_19753,N_13621,N_12888);
and U19754 (N_19754,N_13801,N_11811);
and U19755 (N_19755,N_12440,N_12199);
xor U19756 (N_19756,N_13348,N_14349);
or U19757 (N_19757,N_11907,N_10850);
or U19758 (N_19758,N_14122,N_11914);
nand U19759 (N_19759,N_14398,N_13298);
or U19760 (N_19760,N_11911,N_12699);
nand U19761 (N_19761,N_10064,N_14967);
nand U19762 (N_19762,N_12806,N_11341);
and U19763 (N_19763,N_11913,N_11430);
nand U19764 (N_19764,N_12238,N_10832);
nand U19765 (N_19765,N_11823,N_11571);
nand U19766 (N_19766,N_12739,N_13160);
or U19767 (N_19767,N_12035,N_10015);
and U19768 (N_19768,N_13510,N_10924);
or U19769 (N_19769,N_10430,N_12868);
or U19770 (N_19770,N_11368,N_14474);
nor U19771 (N_19771,N_10867,N_13483);
or U19772 (N_19772,N_14615,N_12601);
or U19773 (N_19773,N_11202,N_12570);
and U19774 (N_19774,N_13271,N_10094);
nand U19775 (N_19775,N_14930,N_12227);
or U19776 (N_19776,N_12374,N_14057);
nor U19777 (N_19777,N_10799,N_14598);
nand U19778 (N_19778,N_13904,N_11115);
or U19779 (N_19779,N_12838,N_10358);
nand U19780 (N_19780,N_14276,N_13934);
xor U19781 (N_19781,N_10141,N_10946);
nor U19782 (N_19782,N_14137,N_14267);
or U19783 (N_19783,N_14781,N_13983);
or U19784 (N_19784,N_10530,N_14815);
or U19785 (N_19785,N_12098,N_12101);
or U19786 (N_19786,N_10398,N_13989);
or U19787 (N_19787,N_12465,N_11262);
or U19788 (N_19788,N_13235,N_13031);
nor U19789 (N_19789,N_12488,N_10199);
nor U19790 (N_19790,N_12506,N_12854);
or U19791 (N_19791,N_10913,N_11319);
and U19792 (N_19792,N_10452,N_11630);
nand U19793 (N_19793,N_12944,N_10769);
and U19794 (N_19794,N_14178,N_11058);
nor U19795 (N_19795,N_10687,N_13472);
nand U19796 (N_19796,N_12442,N_12490);
and U19797 (N_19797,N_11907,N_14006);
or U19798 (N_19798,N_13520,N_14021);
and U19799 (N_19799,N_12137,N_10932);
nor U19800 (N_19800,N_11690,N_12345);
or U19801 (N_19801,N_10767,N_11100);
or U19802 (N_19802,N_13231,N_11891);
nand U19803 (N_19803,N_13607,N_10152);
and U19804 (N_19804,N_11080,N_11510);
nor U19805 (N_19805,N_14711,N_13702);
nand U19806 (N_19806,N_11550,N_13635);
or U19807 (N_19807,N_11414,N_10715);
or U19808 (N_19808,N_13932,N_12204);
nor U19809 (N_19809,N_10050,N_10475);
or U19810 (N_19810,N_10375,N_11574);
nor U19811 (N_19811,N_10520,N_13846);
and U19812 (N_19812,N_11541,N_11014);
and U19813 (N_19813,N_10554,N_14763);
or U19814 (N_19814,N_13114,N_11617);
nor U19815 (N_19815,N_13587,N_11824);
or U19816 (N_19816,N_13891,N_12433);
or U19817 (N_19817,N_10413,N_10739);
nor U19818 (N_19818,N_10322,N_11853);
and U19819 (N_19819,N_12471,N_11806);
nor U19820 (N_19820,N_14414,N_13693);
or U19821 (N_19821,N_13484,N_12082);
and U19822 (N_19822,N_12494,N_11926);
and U19823 (N_19823,N_10060,N_10928);
and U19824 (N_19824,N_12407,N_11653);
or U19825 (N_19825,N_12924,N_13771);
nor U19826 (N_19826,N_14173,N_11816);
or U19827 (N_19827,N_11585,N_13621);
or U19828 (N_19828,N_14354,N_12882);
or U19829 (N_19829,N_13606,N_14413);
nor U19830 (N_19830,N_10836,N_13856);
nor U19831 (N_19831,N_12017,N_10621);
or U19832 (N_19832,N_10054,N_14533);
or U19833 (N_19833,N_14200,N_14525);
or U19834 (N_19834,N_13991,N_12548);
or U19835 (N_19835,N_10618,N_12764);
or U19836 (N_19836,N_14456,N_11608);
nor U19837 (N_19837,N_11322,N_14884);
nand U19838 (N_19838,N_11216,N_14127);
xor U19839 (N_19839,N_11906,N_13017);
nand U19840 (N_19840,N_10383,N_13513);
xnor U19841 (N_19841,N_11362,N_10273);
nand U19842 (N_19842,N_13132,N_12101);
and U19843 (N_19843,N_10393,N_14841);
and U19844 (N_19844,N_10549,N_13794);
nand U19845 (N_19845,N_10275,N_11631);
or U19846 (N_19846,N_11155,N_12940);
and U19847 (N_19847,N_14478,N_14874);
nor U19848 (N_19848,N_12441,N_14481);
and U19849 (N_19849,N_10867,N_10837);
or U19850 (N_19850,N_14766,N_13686);
nor U19851 (N_19851,N_11947,N_10923);
nor U19852 (N_19852,N_14727,N_13900);
nor U19853 (N_19853,N_12934,N_10815);
nand U19854 (N_19854,N_14522,N_12255);
nor U19855 (N_19855,N_13419,N_13973);
or U19856 (N_19856,N_12010,N_14789);
nor U19857 (N_19857,N_12574,N_13912);
nor U19858 (N_19858,N_14577,N_12161);
or U19859 (N_19859,N_14414,N_11102);
or U19860 (N_19860,N_12491,N_12566);
or U19861 (N_19861,N_13379,N_13841);
or U19862 (N_19862,N_14011,N_10941);
and U19863 (N_19863,N_14655,N_12061);
nor U19864 (N_19864,N_14572,N_14460);
and U19865 (N_19865,N_14888,N_10722);
nand U19866 (N_19866,N_12243,N_10067);
or U19867 (N_19867,N_12302,N_10849);
and U19868 (N_19868,N_13067,N_10236);
nor U19869 (N_19869,N_11712,N_11808);
or U19870 (N_19870,N_12272,N_12457);
nand U19871 (N_19871,N_11891,N_12487);
nor U19872 (N_19872,N_14498,N_11927);
or U19873 (N_19873,N_10627,N_14706);
and U19874 (N_19874,N_13547,N_14343);
and U19875 (N_19875,N_13939,N_10676);
and U19876 (N_19876,N_11735,N_12348);
nor U19877 (N_19877,N_13115,N_11594);
or U19878 (N_19878,N_10840,N_11023);
or U19879 (N_19879,N_13938,N_14878);
or U19880 (N_19880,N_12722,N_14684);
or U19881 (N_19881,N_10018,N_13557);
nand U19882 (N_19882,N_14820,N_14693);
and U19883 (N_19883,N_10497,N_11967);
and U19884 (N_19884,N_11905,N_12827);
nor U19885 (N_19885,N_12050,N_10648);
nor U19886 (N_19886,N_12245,N_14472);
nor U19887 (N_19887,N_10538,N_12963);
or U19888 (N_19888,N_10918,N_12842);
and U19889 (N_19889,N_11413,N_12292);
nand U19890 (N_19890,N_12939,N_13671);
or U19891 (N_19891,N_11811,N_10690);
nor U19892 (N_19892,N_14193,N_10950);
or U19893 (N_19893,N_14847,N_11309);
and U19894 (N_19894,N_13896,N_10601);
or U19895 (N_19895,N_11328,N_11612);
nor U19896 (N_19896,N_12933,N_10041);
nand U19897 (N_19897,N_12581,N_12667);
and U19898 (N_19898,N_14223,N_13564);
or U19899 (N_19899,N_14984,N_14699);
nand U19900 (N_19900,N_10620,N_11172);
or U19901 (N_19901,N_12184,N_11814);
nand U19902 (N_19902,N_14317,N_11862);
nor U19903 (N_19903,N_14081,N_10803);
nor U19904 (N_19904,N_12816,N_10272);
nor U19905 (N_19905,N_14787,N_14404);
nand U19906 (N_19906,N_11002,N_11742);
nor U19907 (N_19907,N_11747,N_12706);
nor U19908 (N_19908,N_12568,N_12115);
xnor U19909 (N_19909,N_11038,N_14262);
nand U19910 (N_19910,N_12500,N_13518);
and U19911 (N_19911,N_11371,N_11812);
xor U19912 (N_19912,N_11006,N_11982);
nand U19913 (N_19913,N_12857,N_12268);
or U19914 (N_19914,N_14017,N_10004);
or U19915 (N_19915,N_13832,N_14738);
and U19916 (N_19916,N_11566,N_14392);
nor U19917 (N_19917,N_12408,N_14537);
or U19918 (N_19918,N_14982,N_11874);
and U19919 (N_19919,N_10816,N_11583);
nand U19920 (N_19920,N_13858,N_13076);
or U19921 (N_19921,N_14450,N_10109);
and U19922 (N_19922,N_12221,N_11965);
or U19923 (N_19923,N_12792,N_10617);
nand U19924 (N_19924,N_10103,N_11213);
nor U19925 (N_19925,N_11918,N_13582);
xor U19926 (N_19926,N_14402,N_10198);
nor U19927 (N_19927,N_14455,N_12205);
nor U19928 (N_19928,N_10311,N_11937);
or U19929 (N_19929,N_11295,N_14416);
or U19930 (N_19930,N_13104,N_13882);
nor U19931 (N_19931,N_10496,N_10903);
nor U19932 (N_19932,N_10222,N_12424);
nand U19933 (N_19933,N_13319,N_11913);
and U19934 (N_19934,N_11228,N_14925);
nand U19935 (N_19935,N_13379,N_10932);
and U19936 (N_19936,N_10769,N_14677);
nand U19937 (N_19937,N_11349,N_11097);
nand U19938 (N_19938,N_13056,N_11658);
nand U19939 (N_19939,N_13031,N_11986);
and U19940 (N_19940,N_14627,N_10430);
or U19941 (N_19941,N_13000,N_10497);
nor U19942 (N_19942,N_10680,N_13179);
nand U19943 (N_19943,N_11027,N_13275);
nand U19944 (N_19944,N_13520,N_11916);
and U19945 (N_19945,N_10393,N_12034);
nand U19946 (N_19946,N_13505,N_11249);
and U19947 (N_19947,N_10145,N_10154);
and U19948 (N_19948,N_10844,N_13416);
and U19949 (N_19949,N_13013,N_14323);
and U19950 (N_19950,N_10094,N_11148);
nor U19951 (N_19951,N_11573,N_13218);
or U19952 (N_19952,N_13761,N_13114);
nand U19953 (N_19953,N_12965,N_13376);
nor U19954 (N_19954,N_10818,N_14922);
nand U19955 (N_19955,N_11553,N_14529);
nor U19956 (N_19956,N_11162,N_11871);
or U19957 (N_19957,N_12164,N_12231);
nor U19958 (N_19958,N_12210,N_13287);
nand U19959 (N_19959,N_13222,N_13603);
nor U19960 (N_19960,N_14040,N_12507);
nor U19961 (N_19961,N_13234,N_11980);
and U19962 (N_19962,N_12077,N_14188);
nor U19963 (N_19963,N_12733,N_13235);
nand U19964 (N_19964,N_11743,N_12137);
nand U19965 (N_19965,N_12851,N_11243);
nor U19966 (N_19966,N_13689,N_12882);
or U19967 (N_19967,N_13700,N_11338);
and U19968 (N_19968,N_10404,N_14775);
xnor U19969 (N_19969,N_14650,N_14379);
and U19970 (N_19970,N_13009,N_10754);
nor U19971 (N_19971,N_14179,N_11812);
nor U19972 (N_19972,N_14458,N_13154);
and U19973 (N_19973,N_10073,N_14114);
or U19974 (N_19974,N_10685,N_11915);
xnor U19975 (N_19975,N_13125,N_13041);
nand U19976 (N_19976,N_10710,N_11006);
nand U19977 (N_19977,N_12509,N_12814);
or U19978 (N_19978,N_13313,N_10415);
or U19979 (N_19979,N_14837,N_11979);
nand U19980 (N_19980,N_13403,N_12821);
or U19981 (N_19981,N_14898,N_10890);
and U19982 (N_19982,N_14941,N_10304);
or U19983 (N_19983,N_12135,N_14165);
and U19984 (N_19984,N_13514,N_13158);
nor U19985 (N_19985,N_11621,N_12912);
nor U19986 (N_19986,N_12385,N_10256);
or U19987 (N_19987,N_13534,N_11036);
nor U19988 (N_19988,N_10264,N_14460);
nand U19989 (N_19989,N_11060,N_10000);
or U19990 (N_19990,N_14697,N_10494);
or U19991 (N_19991,N_10980,N_14194);
or U19992 (N_19992,N_12286,N_14912);
and U19993 (N_19993,N_10976,N_11661);
nor U19994 (N_19994,N_10078,N_13784);
nor U19995 (N_19995,N_13033,N_10912);
nor U19996 (N_19996,N_12614,N_11238);
nor U19997 (N_19997,N_11281,N_12772);
or U19998 (N_19998,N_11884,N_10075);
and U19999 (N_19999,N_10182,N_14779);
or U20000 (N_20000,N_18018,N_15157);
nor U20001 (N_20001,N_18953,N_19201);
or U20002 (N_20002,N_16400,N_19188);
nor U20003 (N_20003,N_15300,N_16051);
nand U20004 (N_20004,N_15115,N_19828);
nand U20005 (N_20005,N_15452,N_19434);
nand U20006 (N_20006,N_15713,N_16218);
nor U20007 (N_20007,N_15118,N_16197);
or U20008 (N_20008,N_19449,N_15168);
and U20009 (N_20009,N_18071,N_17498);
and U20010 (N_20010,N_19132,N_19672);
or U20011 (N_20011,N_15373,N_18745);
nor U20012 (N_20012,N_19680,N_18184);
nor U20013 (N_20013,N_19870,N_15725);
and U20014 (N_20014,N_17445,N_15439);
and U20015 (N_20015,N_15034,N_17816);
xor U20016 (N_20016,N_18771,N_18848);
or U20017 (N_20017,N_18143,N_16925);
nand U20018 (N_20018,N_18947,N_16377);
nor U20019 (N_20019,N_15987,N_17468);
nand U20020 (N_20020,N_15128,N_17318);
nor U20021 (N_20021,N_17725,N_16978);
and U20022 (N_20022,N_19322,N_16044);
nand U20023 (N_20023,N_19992,N_17769);
or U20024 (N_20024,N_15990,N_15763);
nand U20025 (N_20025,N_17357,N_15038);
and U20026 (N_20026,N_16015,N_17044);
nand U20027 (N_20027,N_19304,N_19288);
or U20028 (N_20028,N_19377,N_18639);
nand U20029 (N_20029,N_18204,N_15814);
or U20030 (N_20030,N_16237,N_17108);
and U20031 (N_20031,N_18797,N_15818);
or U20032 (N_20032,N_16369,N_15614);
or U20033 (N_20033,N_17767,N_16178);
xnor U20034 (N_20034,N_16785,N_18139);
and U20035 (N_20035,N_17989,N_19323);
or U20036 (N_20036,N_15766,N_18834);
and U20037 (N_20037,N_18701,N_18826);
nor U20038 (N_20038,N_16936,N_17556);
or U20039 (N_20039,N_19348,N_15385);
nand U20040 (N_20040,N_19755,N_18839);
nor U20041 (N_20041,N_15687,N_16652);
or U20042 (N_20042,N_16518,N_16048);
or U20043 (N_20043,N_17724,N_19292);
and U20044 (N_20044,N_17535,N_15060);
nor U20045 (N_20045,N_19813,N_16143);
or U20046 (N_20046,N_16150,N_15553);
and U20047 (N_20047,N_18296,N_15602);
nor U20048 (N_20048,N_18636,N_18115);
and U20049 (N_20049,N_15556,N_16277);
nor U20050 (N_20050,N_17890,N_15925);
and U20051 (N_20051,N_19553,N_17995);
nand U20052 (N_20052,N_18183,N_17040);
and U20053 (N_20053,N_18161,N_15457);
or U20054 (N_20054,N_18149,N_15174);
or U20055 (N_20055,N_18337,N_19613);
and U20056 (N_20056,N_16406,N_19668);
nand U20057 (N_20057,N_17781,N_16991);
nor U20058 (N_20058,N_18147,N_16522);
and U20059 (N_20059,N_17833,N_18578);
nor U20060 (N_20060,N_19407,N_15285);
nand U20061 (N_20061,N_16901,N_16834);
nand U20062 (N_20062,N_17695,N_19231);
or U20063 (N_20063,N_17519,N_19906);
nand U20064 (N_20064,N_19543,N_16697);
or U20065 (N_20065,N_17934,N_19776);
nor U20066 (N_20066,N_18682,N_15829);
or U20067 (N_20067,N_18440,N_18882);
nand U20068 (N_20068,N_16288,N_16055);
or U20069 (N_20069,N_17828,N_16095);
and U20070 (N_20070,N_17495,N_16350);
nand U20071 (N_20071,N_19485,N_19661);
and U20072 (N_20072,N_18508,N_19749);
nand U20073 (N_20073,N_17999,N_18692);
and U20074 (N_20074,N_19036,N_19071);
nor U20075 (N_20075,N_18698,N_17602);
nor U20076 (N_20076,N_19152,N_17452);
nand U20077 (N_20077,N_17238,N_16361);
nor U20078 (N_20078,N_19197,N_15479);
or U20079 (N_20079,N_19226,N_16425);
nand U20080 (N_20080,N_17815,N_19985);
nor U20081 (N_20081,N_17218,N_18408);
nand U20082 (N_20082,N_18786,N_18145);
and U20083 (N_20083,N_15578,N_15121);
nor U20084 (N_20084,N_16411,N_19527);
or U20085 (N_20085,N_17497,N_18423);
nor U20086 (N_20086,N_19843,N_17196);
nand U20087 (N_20087,N_19957,N_16018);
or U20088 (N_20088,N_15098,N_15521);
or U20089 (N_20089,N_16307,N_17773);
and U20090 (N_20090,N_17149,N_15887);
or U20091 (N_20091,N_19691,N_18643);
and U20092 (N_20092,N_16152,N_15377);
or U20093 (N_20093,N_17782,N_18413);
nor U20094 (N_20094,N_16465,N_15771);
nor U20095 (N_20095,N_15628,N_18274);
or U20096 (N_20096,N_17908,N_17041);
and U20097 (N_20097,N_17619,N_17387);
nor U20098 (N_20098,N_19903,N_18481);
nor U20099 (N_20099,N_16679,N_17487);
nor U20100 (N_20100,N_15367,N_19161);
and U20101 (N_20101,N_16003,N_18835);
nor U20102 (N_20102,N_18124,N_18637);
or U20103 (N_20103,N_15085,N_16342);
and U20104 (N_20104,N_15131,N_17838);
and U20105 (N_20105,N_18689,N_16185);
nor U20106 (N_20106,N_19917,N_17391);
nand U20107 (N_20107,N_18671,N_18005);
or U20108 (N_20108,N_18220,N_18444);
nor U20109 (N_20109,N_15580,N_18592);
and U20110 (N_20110,N_18031,N_18503);
or U20111 (N_20111,N_18978,N_15716);
nand U20112 (N_20112,N_16035,N_17346);
and U20113 (N_20113,N_19009,N_18244);
and U20114 (N_20114,N_16610,N_19682);
and U20115 (N_20115,N_16247,N_16891);
xnor U20116 (N_20116,N_16759,N_18970);
nor U20117 (N_20117,N_19673,N_16407);
nor U20118 (N_20118,N_18109,N_19390);
nor U20119 (N_20119,N_16558,N_15234);
or U20120 (N_20120,N_15254,N_16402);
nand U20121 (N_20121,N_18350,N_16319);
or U20122 (N_20122,N_17875,N_15317);
or U20123 (N_20123,N_15133,N_15808);
nor U20124 (N_20124,N_18465,N_18590);
or U20125 (N_20125,N_19967,N_15338);
nand U20126 (N_20126,N_18787,N_16111);
nand U20127 (N_20127,N_18420,N_19825);
and U20128 (N_20128,N_19632,N_17668);
or U20129 (N_20129,N_18895,N_18487);
nand U20130 (N_20130,N_17775,N_18063);
nand U20131 (N_20131,N_16793,N_15828);
or U20132 (N_20132,N_16364,N_16000);
or U20133 (N_20133,N_16501,N_18373);
and U20134 (N_20134,N_15957,N_16204);
and U20135 (N_20135,N_15113,N_15981);
or U20136 (N_20136,N_18176,N_18218);
and U20137 (N_20137,N_19573,N_17779);
and U20138 (N_20138,N_19261,N_19314);
and U20139 (N_20139,N_17499,N_16931);
or U20140 (N_20140,N_17020,N_17605);
or U20141 (N_20141,N_16630,N_19548);
nand U20142 (N_20142,N_15383,N_17263);
nor U20143 (N_20143,N_17871,N_18309);
nor U20144 (N_20144,N_18362,N_15093);
nand U20145 (N_20145,N_17190,N_19147);
nor U20146 (N_20146,N_15599,N_17293);
or U20147 (N_20147,N_19236,N_16794);
nor U20148 (N_20148,N_19832,N_15052);
and U20149 (N_20149,N_19091,N_18751);
and U20150 (N_20150,N_18633,N_15185);
or U20151 (N_20151,N_18261,N_15425);
xnor U20152 (N_20152,N_16948,N_18320);
or U20153 (N_20153,N_16061,N_19834);
nor U20154 (N_20154,N_18602,N_16315);
nand U20155 (N_20155,N_19396,N_17693);
nor U20156 (N_20156,N_15799,N_18422);
or U20157 (N_20157,N_16126,N_18984);
or U20158 (N_20158,N_16201,N_17913);
or U20159 (N_20159,N_18484,N_17262);
or U20160 (N_20160,N_15688,N_19025);
xnor U20161 (N_20161,N_16603,N_16725);
nand U20162 (N_20162,N_15076,N_18428);
nor U20163 (N_20163,N_16956,N_18126);
nand U20164 (N_20164,N_19972,N_16193);
and U20165 (N_20165,N_17208,N_19833);
nor U20166 (N_20166,N_17155,N_16967);
or U20167 (N_20167,N_18432,N_15105);
and U20168 (N_20168,N_19073,N_18347);
and U20169 (N_20169,N_17427,N_16109);
nand U20170 (N_20170,N_18608,N_18506);
nand U20171 (N_20171,N_15645,N_18459);
nor U20172 (N_20172,N_17527,N_17162);
and U20173 (N_20173,N_18644,N_15576);
and U20174 (N_20174,N_19773,N_16284);
nand U20175 (N_20175,N_16225,N_19808);
nand U20176 (N_20176,N_19165,N_19339);
nor U20177 (N_20177,N_18686,N_16796);
and U20178 (N_20178,N_17233,N_17652);
or U20179 (N_20179,N_17579,N_15730);
or U20180 (N_20180,N_15621,N_18498);
and U20181 (N_20181,N_17603,N_18431);
nor U20182 (N_20182,N_19928,N_18036);
or U20183 (N_20183,N_19757,N_16324);
and U20184 (N_20184,N_16092,N_18348);
nand U20185 (N_20185,N_19409,N_16259);
or U20186 (N_20186,N_15414,N_19358);
nand U20187 (N_20187,N_15805,N_17270);
nand U20188 (N_20188,N_17277,N_18868);
or U20189 (N_20189,N_19079,N_17545);
and U20190 (N_20190,N_16134,N_15978);
and U20191 (N_20191,N_18884,N_15833);
or U20192 (N_20192,N_17011,N_18023);
nand U20193 (N_20193,N_18368,N_19370);
and U20194 (N_20194,N_18222,N_16024);
nand U20195 (N_20195,N_15236,N_15964);
or U20196 (N_20196,N_19248,N_15288);
or U20197 (N_20197,N_19417,N_17068);
and U20198 (N_20198,N_18930,N_15907);
nand U20199 (N_20199,N_19877,N_16171);
nand U20200 (N_20200,N_19986,N_15301);
and U20201 (N_20201,N_17549,N_16886);
nor U20202 (N_20202,N_17830,N_17470);
nor U20203 (N_20203,N_15468,N_15665);
nor U20204 (N_20204,N_15485,N_15582);
or U20205 (N_20205,N_16168,N_15411);
or U20206 (N_20206,N_17111,N_15913);
or U20207 (N_20207,N_15988,N_18951);
and U20208 (N_20208,N_18116,N_18666);
xor U20209 (N_20209,N_18790,N_18726);
nor U20210 (N_20210,N_15504,N_19500);
nor U20211 (N_20211,N_18769,N_18680);
nand U20212 (N_20212,N_15033,N_15870);
nor U20213 (N_20213,N_19621,N_18938);
nand U20214 (N_20214,N_19999,N_16699);
xor U20215 (N_20215,N_18704,N_18825);
and U20216 (N_20216,N_17244,N_15140);
nor U20217 (N_20217,N_15705,N_18104);
nor U20218 (N_20218,N_19931,N_17230);
nor U20219 (N_20219,N_17751,N_15287);
or U20220 (N_20220,N_17415,N_17146);
nor U20221 (N_20221,N_15448,N_18395);
and U20222 (N_20222,N_15011,N_19206);
nand U20223 (N_20223,N_17007,N_19253);
or U20224 (N_20224,N_15890,N_19331);
nand U20225 (N_20225,N_15107,N_18525);
nand U20226 (N_20226,N_18768,N_19614);
or U20227 (N_20227,N_19402,N_18775);
nand U20228 (N_20228,N_17479,N_19320);
nor U20229 (N_20229,N_19752,N_16352);
and U20230 (N_20230,N_17307,N_18851);
nand U20231 (N_20231,N_17932,N_18630);
or U20232 (N_20232,N_19422,N_17043);
xnor U20233 (N_20233,N_15190,N_15183);
nand U20234 (N_20234,N_19041,N_15908);
or U20235 (N_20235,N_17223,N_18194);
nand U20236 (N_20236,N_15119,N_17584);
nand U20237 (N_20237,N_18609,N_16008);
nor U20238 (N_20238,N_16657,N_18522);
nand U20239 (N_20239,N_15002,N_19096);
nor U20240 (N_20240,N_15765,N_18449);
nand U20241 (N_20241,N_18561,N_16912);
nand U20242 (N_20242,N_16928,N_17551);
or U20243 (N_20243,N_18312,N_15712);
nand U20244 (N_20244,N_17435,N_15658);
nand U20245 (N_20245,N_16619,N_17430);
nand U20246 (N_20246,N_17685,N_16641);
and U20247 (N_20247,N_18017,N_18324);
and U20248 (N_20248,N_15848,N_18131);
xnor U20249 (N_20249,N_17600,N_19866);
nor U20250 (N_20250,N_16158,N_19347);
and U20251 (N_20251,N_19381,N_15611);
and U20252 (N_20252,N_18100,N_18725);
nand U20253 (N_20253,N_15530,N_15864);
or U20254 (N_20254,N_19905,N_15594);
or U20255 (N_20255,N_18586,N_17206);
nand U20256 (N_20256,N_15027,N_18392);
nor U20257 (N_20257,N_15144,N_19232);
nor U20258 (N_20258,N_17016,N_19809);
nand U20259 (N_20259,N_17951,N_19030);
and U20260 (N_20260,N_18537,N_19975);
nor U20261 (N_20261,N_17836,N_16039);
or U20262 (N_20262,N_18495,N_17275);
nor U20263 (N_20263,N_19305,N_15895);
nor U20264 (N_20264,N_19419,N_15363);
nand U20265 (N_20265,N_19574,N_17219);
or U20266 (N_20266,N_15559,N_19272);
nand U20267 (N_20267,N_15492,N_18605);
xor U20268 (N_20268,N_19094,N_18654);
nor U20269 (N_20269,N_17532,N_16676);
nand U20270 (N_20270,N_16066,N_17115);
nor U20271 (N_20271,N_15415,N_17911);
nor U20272 (N_20272,N_18518,N_17753);
nand U20273 (N_20273,N_19430,N_15336);
nand U20274 (N_20274,N_16496,N_17594);
and U20275 (N_20275,N_17159,N_16394);
nor U20276 (N_20276,N_18103,N_19919);
and U20277 (N_20277,N_15748,N_18824);
and U20278 (N_20278,N_17083,N_15695);
nand U20279 (N_20279,N_19850,N_19101);
nand U20280 (N_20280,N_18833,N_18599);
nor U20281 (N_20281,N_16615,N_15255);
nor U20282 (N_20282,N_15539,N_16416);
xnor U20283 (N_20283,N_18809,N_15785);
nand U20284 (N_20284,N_18723,N_19782);
nor U20285 (N_20285,N_19117,N_18200);
nor U20286 (N_20286,N_16002,N_17849);
or U20287 (N_20287,N_17744,N_17252);
nand U20288 (N_20288,N_17312,N_17475);
nand U20289 (N_20289,N_17938,N_19839);
and U20290 (N_20290,N_16596,N_17260);
nand U20291 (N_20291,N_19436,N_17258);
and U20292 (N_20292,N_15718,N_18946);
or U20293 (N_20293,N_18750,N_19530);
and U20294 (N_20294,N_18285,N_18094);
or U20295 (N_20295,N_19921,N_15616);
nor U20296 (N_20296,N_19733,N_15560);
or U20297 (N_20297,N_16175,N_18539);
and U20298 (N_20298,N_17009,N_17082);
or U20299 (N_20299,N_19788,N_16401);
and U20300 (N_20300,N_15866,N_19863);
nand U20301 (N_20301,N_16627,N_17033);
or U20302 (N_20302,N_18155,N_16285);
and U20303 (N_20303,N_16223,N_18494);
nor U20304 (N_20304,N_15752,N_19851);
nand U20305 (N_20305,N_17364,N_15470);
or U20306 (N_20306,N_17133,N_15063);
nor U20307 (N_20307,N_16161,N_17559);
or U20308 (N_20308,N_18904,N_19059);
nand U20309 (N_20309,N_18684,N_19031);
nand U20310 (N_20310,N_16575,N_15181);
and U20311 (N_20311,N_17440,N_18893);
and U20312 (N_20312,N_16778,N_15788);
nand U20313 (N_20313,N_18897,N_18173);
nor U20314 (N_20314,N_18697,N_16238);
and U20315 (N_20315,N_19431,N_15004);
and U20316 (N_20316,N_18016,N_17735);
or U20317 (N_20317,N_17237,N_16494);
and U20318 (N_20318,N_18687,N_15565);
nor U20319 (N_20319,N_16325,N_17311);
and U20320 (N_20320,N_19544,N_17862);
nor U20321 (N_20321,N_15428,N_17176);
and U20322 (N_20322,N_19926,N_15784);
and U20323 (N_20323,N_17654,N_15329);
or U20324 (N_20324,N_17558,N_19357);
nand U20325 (N_20325,N_16846,N_18044);
nand U20326 (N_20326,N_17937,N_15700);
nand U20327 (N_20327,N_17847,N_16074);
nor U20328 (N_20328,N_16644,N_18264);
or U20329 (N_20329,N_19476,N_16792);
or U20330 (N_20330,N_17632,N_17842);
and U20331 (N_20331,N_17548,N_16638);
or U20332 (N_20332,N_19074,N_17462);
nand U20333 (N_20333,N_16137,N_15178);
and U20334 (N_20334,N_19250,N_19647);
or U20335 (N_20335,N_15787,N_18932);
nand U20336 (N_20336,N_16128,N_16437);
or U20337 (N_20337,N_16892,N_15648);
or U20338 (N_20338,N_15996,N_16952);
xor U20339 (N_20339,N_16403,N_17340);
or U20340 (N_20340,N_15324,N_15495);
xor U20341 (N_20341,N_18646,N_15571);
or U20342 (N_20342,N_15677,N_19715);
or U20343 (N_20343,N_18998,N_16296);
nand U20344 (N_20344,N_17129,N_17099);
and U20345 (N_20345,N_18479,N_17178);
and U20346 (N_20346,N_17413,N_19504);
and U20347 (N_20347,N_19064,N_17513);
xor U20348 (N_20348,N_17997,N_18955);
nor U20349 (N_20349,N_17521,N_17682);
and U20350 (N_20350,N_19066,N_16538);
nand U20351 (N_20351,N_15047,N_16224);
and U20352 (N_20352,N_19051,N_16981);
xnor U20353 (N_20353,N_15424,N_17097);
nor U20354 (N_20354,N_18042,N_17386);
nand U20355 (N_20355,N_18836,N_15949);
and U20356 (N_20356,N_15597,N_19075);
nand U20357 (N_20357,N_15213,N_15170);
nor U20358 (N_20358,N_19677,N_19435);
nor U20359 (N_20359,N_17402,N_16413);
nor U20360 (N_20360,N_15362,N_17666);
nand U20361 (N_20361,N_16739,N_17571);
nor U20362 (N_20362,N_19191,N_15447);
and U20363 (N_20363,N_15745,N_17780);
nand U20364 (N_20364,N_18782,N_19328);
nor U20365 (N_20365,N_18731,N_15500);
nand U20366 (N_20366,N_18753,N_18593);
and U20367 (N_20367,N_19960,N_17360);
nor U20368 (N_20368,N_19103,N_16426);
and U20369 (N_20369,N_15820,N_19125);
nand U20370 (N_20370,N_15333,N_18365);
and U20371 (N_20371,N_15880,N_19675);
nor U20372 (N_20372,N_15477,N_19093);
nor U20373 (N_20373,N_16862,N_17590);
nor U20374 (N_20374,N_17810,N_15159);
or U20375 (N_20375,N_16379,N_16316);
nand U20376 (N_20376,N_18253,N_18118);
nand U20377 (N_20377,N_17761,N_18177);
and U20378 (N_20378,N_17931,N_17800);
or U20379 (N_20379,N_16970,N_16208);
and U20380 (N_20380,N_17152,N_19607);
nor U20381 (N_20381,N_15782,N_18729);
or U20382 (N_20382,N_15789,N_19455);
nor U20383 (N_20383,N_16682,N_19873);
or U20384 (N_20384,N_18794,N_19216);
and U20385 (N_20385,N_17737,N_18454);
or U20386 (N_20386,N_17803,N_18781);
and U20387 (N_20387,N_19172,N_18263);
nand U20388 (N_20388,N_19349,N_15844);
and U20389 (N_20389,N_16810,N_19134);
nor U20390 (N_20390,N_15619,N_18394);
and U20391 (N_20391,N_18961,N_16607);
and U20392 (N_20392,N_15767,N_18547);
nor U20393 (N_20393,N_18798,N_16056);
nor U20394 (N_20394,N_17128,N_18976);
nor U20395 (N_20395,N_15821,N_16669);
nor U20396 (N_20396,N_15845,N_15497);
nor U20397 (N_20397,N_19518,N_18265);
and U20398 (N_20398,N_18128,N_16539);
or U20399 (N_20399,N_18409,N_16083);
or U20400 (N_20400,N_17713,N_18744);
and U20401 (N_20401,N_18795,N_15846);
nand U20402 (N_20402,N_18702,N_19107);
and U20403 (N_20403,N_15146,N_19441);
nand U20404 (N_20404,N_19592,N_16144);
nand U20405 (N_20405,N_15867,N_15192);
or U20406 (N_20406,N_16821,N_16177);
nand U20407 (N_20407,N_16578,N_18854);
and U20408 (N_20408,N_17031,N_15370);
nor U20409 (N_20409,N_16833,N_15145);
nor U20410 (N_20410,N_17329,N_15360);
nand U20411 (N_20411,N_16436,N_16703);
and U20412 (N_20412,N_18617,N_19380);
nor U20413 (N_20413,N_15777,N_18530);
nor U20414 (N_20414,N_16852,N_19619);
and U20415 (N_20415,N_17483,N_15350);
or U20416 (N_20416,N_19575,N_16447);
and U20417 (N_20417,N_19277,N_19516);
nor U20418 (N_20418,N_19800,N_19251);
and U20419 (N_20419,N_19506,N_15888);
and U20420 (N_20420,N_18910,N_18496);
nand U20421 (N_20421,N_16365,N_15282);
and U20422 (N_20422,N_18127,N_16303);
or U20423 (N_20423,N_16561,N_15847);
nand U20424 (N_20424,N_18532,N_19252);
nand U20425 (N_20425,N_19481,N_18690);
nor U20426 (N_20426,N_19589,N_17586);
or U20427 (N_20427,N_19984,N_17118);
nand U20428 (N_20428,N_19037,N_15815);
nand U20429 (N_20429,N_15358,N_19141);
and U20430 (N_20430,N_15876,N_17096);
nor U20431 (N_20431,N_17471,N_15618);
nand U20432 (N_20432,N_17887,N_18972);
or U20433 (N_20433,N_17198,N_19652);
nor U20434 (N_20434,N_17689,N_18371);
or U20435 (N_20435,N_15983,N_18401);
nand U20436 (N_20436,N_19955,N_16357);
and U20437 (N_20437,N_16019,N_16849);
or U20438 (N_20438,N_16060,N_16478);
nor U20439 (N_20439,N_18950,N_18258);
nor U20440 (N_20440,N_15603,N_18317);
or U20441 (N_20441,N_18847,N_16932);
or U20442 (N_20442,N_18962,N_18006);
nor U20443 (N_20443,N_19149,N_18445);
nand U20444 (N_20444,N_17211,N_16301);
nor U20445 (N_20445,N_17382,N_15882);
and U20446 (N_20446,N_15778,N_18247);
and U20447 (N_20447,N_19080,N_15155);
and U20448 (N_20448,N_15064,N_17651);
or U20449 (N_20449,N_18516,N_15268);
nor U20450 (N_20450,N_19403,N_15933);
and U20451 (N_20451,N_19519,N_16546);
or U20452 (N_20452,N_15281,N_18448);
or U20453 (N_20453,N_17840,N_16995);
nand U20454 (N_20454,N_15496,N_18675);
nand U20455 (N_20455,N_15904,N_15195);
and U20456 (N_20456,N_17848,N_19317);
nor U20457 (N_20457,N_16755,N_19943);
and U20458 (N_20458,N_16283,N_17540);
and U20459 (N_20459,N_18164,N_16151);
and U20460 (N_20460,N_15094,N_16495);
nor U20461 (N_20461,N_19827,N_17640);
nor U20462 (N_20462,N_18133,N_17557);
and U20463 (N_20463,N_19491,N_16651);
nand U20464 (N_20464,N_17952,N_17730);
or U20465 (N_20465,N_17524,N_17375);
xor U20466 (N_20466,N_18733,N_15466);
nand U20467 (N_20467,N_19872,N_16840);
or U20468 (N_20468,N_18476,N_16441);
nand U20469 (N_20469,N_17877,N_18566);
and U20470 (N_20470,N_15364,N_19653);
and U20471 (N_20471,N_19745,N_16408);
nand U20472 (N_20472,N_15985,N_17696);
nor U20473 (N_20473,N_18385,N_19439);
and U20474 (N_20474,N_18575,N_15852);
nor U20475 (N_20475,N_19609,N_18649);
nor U20476 (N_20476,N_16213,N_16349);
and U20477 (N_20477,N_16409,N_16842);
and U20478 (N_20478,N_19517,N_15441);
and U20479 (N_20479,N_16587,N_15859);
and U20480 (N_20480,N_16242,N_16639);
nand U20481 (N_20481,N_17804,N_19535);
xnor U20482 (N_20482,N_15652,N_18523);
nand U20483 (N_20483,N_16454,N_15494);
nor U20484 (N_20484,N_18340,N_15642);
nand U20485 (N_20485,N_18555,N_17570);
or U20486 (N_20486,N_17676,N_16383);
nor U20487 (N_20487,N_18252,N_18902);
nor U20488 (N_20488,N_19166,N_16022);
or U20489 (N_20489,N_17589,N_18764);
nor U20490 (N_20490,N_16076,N_16067);
and U20491 (N_20491,N_16873,N_19708);
and U20492 (N_20492,N_18082,N_19704);
nand U20493 (N_20493,N_19362,N_17817);
nand U20494 (N_20494,N_18339,N_16690);
and U20495 (N_20495,N_17073,N_15206);
nor U20496 (N_20496,N_18217,N_17726);
nor U20497 (N_20497,N_15111,N_17698);
and U20498 (N_20498,N_16354,N_18308);
nor U20499 (N_20499,N_18918,N_16512);
and U20500 (N_20500,N_18820,N_17740);
and U20501 (N_20501,N_16551,N_15982);
or U20502 (N_20502,N_17745,N_19204);
and U20503 (N_20503,N_18914,N_15309);
and U20504 (N_20504,N_18249,N_19842);
and U20505 (N_20505,N_18681,N_17691);
or U20506 (N_20506,N_16773,N_18211);
and U20507 (N_20507,N_18327,N_19977);
nor U20508 (N_20508,N_16255,N_19119);
nor U20509 (N_20509,N_16841,N_19330);
nor U20510 (N_20510,N_16986,N_18858);
or U20511 (N_20511,N_18841,N_19656);
and U20512 (N_20512,N_15433,N_16291);
nand U20513 (N_20513,N_18160,N_17986);
nor U20514 (N_20514,N_15232,N_15082);
and U20515 (N_20515,N_19214,N_19560);
nand U20516 (N_20516,N_18658,N_15334);
or U20517 (N_20517,N_19319,N_18192);
nand U20518 (N_20518,N_16199,N_19908);
xnor U20519 (N_20519,N_15632,N_18638);
nor U20520 (N_20520,N_19948,N_19978);
xnor U20521 (N_20521,N_15555,N_17322);
and U20522 (N_20522,N_15493,N_16065);
xnor U20523 (N_20523,N_17212,N_18270);
xnor U20524 (N_20524,N_17976,N_16129);
or U20525 (N_20525,N_18528,N_18332);
or U20526 (N_20526,N_18812,N_16906);
nor U20527 (N_20527,N_19286,N_15971);
and U20528 (N_20528,N_19545,N_15629);
or U20529 (N_20529,N_16813,N_18936);
nand U20530 (N_20530,N_16599,N_18840);
nor U20531 (N_20531,N_19720,N_15813);
or U20532 (N_20532,N_15838,N_18310);
nor U20533 (N_20533,N_19791,N_16336);
nor U20534 (N_20534,N_17087,N_18709);
or U20535 (N_20535,N_18367,N_15921);
or U20536 (N_20536,N_19572,N_19238);
nand U20537 (N_20537,N_19712,N_15233);
and U20538 (N_20538,N_16311,N_17958);
or U20539 (N_20539,N_17410,N_17002);
nor U20540 (N_20540,N_18534,N_18334);
nand U20541 (N_20541,N_18306,N_15676);
and U20542 (N_20542,N_16358,N_16613);
and U20543 (N_20543,N_19684,N_15250);
nor U20544 (N_20544,N_15352,N_17981);
and U20545 (N_20545,N_17088,N_16875);
and U20546 (N_20546,N_17880,N_18655);
nor U20547 (N_20547,N_19930,N_19775);
nor U20548 (N_20548,N_19650,N_18239);
nand U20549 (N_20549,N_17010,N_17175);
nand U20550 (N_20550,N_17720,N_16474);
and U20551 (N_20551,N_19706,N_17143);
and U20552 (N_20552,N_17463,N_16040);
nor U20553 (N_20553,N_18114,N_16655);
or U20554 (N_20554,N_17345,N_17843);
or U20555 (N_20555,N_17091,N_15179);
nand U20556 (N_20556,N_16477,N_19634);
or U20557 (N_20557,N_19212,N_17778);
nor U20558 (N_20558,N_18182,N_16781);
nand U20559 (N_20559,N_15823,N_16355);
or U20560 (N_20560,N_17655,N_15562);
or U20561 (N_20561,N_19528,N_15357);
and U20562 (N_20562,N_15152,N_19584);
or U20563 (N_20563,N_17331,N_17940);
and U20564 (N_20564,N_15343,N_16902);
nor U20565 (N_20565,N_15786,N_16733);
and U20566 (N_20566,N_17358,N_16890);
and U20567 (N_20567,N_16112,N_18915);
nor U20568 (N_20568,N_15734,N_17625);
and U20569 (N_20569,N_18908,N_15110);
and U20570 (N_20570,N_17205,N_16788);
or U20571 (N_20571,N_15995,N_19750);
nand U20572 (N_20572,N_16216,N_18468);
nor U20573 (N_20573,N_17736,N_19418);
nor U20574 (N_20574,N_15227,N_18527);
or U20575 (N_20575,N_15217,N_15694);
and U20576 (N_20576,N_16735,N_15761);
nor U20577 (N_20577,N_18033,N_18075);
nand U20578 (N_20578,N_19954,N_19624);
and U20579 (N_20579,N_17975,N_19269);
or U20580 (N_20580,N_19658,N_16410);
or U20581 (N_20581,N_17451,N_19356);
or U20582 (N_20582,N_18906,N_17458);
nand U20583 (N_20583,N_19932,N_17859);
nor U20584 (N_20584,N_19089,N_17138);
xnor U20585 (N_20585,N_18907,N_15526);
nor U20586 (N_20586,N_16632,N_15164);
or U20587 (N_20587,N_18529,N_17588);
or U20588 (N_20588,N_15125,N_17624);
nor U20589 (N_20589,N_19335,N_17119);
or U20590 (N_20590,N_19070,N_17174);
and U20591 (N_20591,N_18271,N_17147);
nor U20592 (N_20592,N_18142,N_19388);
nand U20593 (N_20593,N_17642,N_18355);
nor U20594 (N_20594,N_18819,N_16321);
nor U20595 (N_20595,N_19368,N_19293);
nor U20596 (N_20596,N_17661,N_15691);
nand U20597 (N_20597,N_19770,N_18469);
and U20598 (N_20598,N_19427,N_15382);
nand U20599 (N_20599,N_17376,N_19502);
xnor U20600 (N_20600,N_17139,N_15266);
nor U20601 (N_20601,N_18916,N_16190);
or U20602 (N_20602,N_18966,N_15592);
nand U20603 (N_20603,N_17144,N_16674);
nor U20604 (N_20604,N_19379,N_16577);
and U20605 (N_20605,N_18284,N_15931);
and U20606 (N_20606,N_16855,N_17669);
nand U20607 (N_20607,N_18038,N_17921);
and U20608 (N_20608,N_18703,N_16455);
nand U20609 (N_20609,N_18993,N_19265);
or U20610 (N_20610,N_17494,N_16562);
nor U20611 (N_20611,N_15215,N_16582);
nor U20612 (N_20612,N_19284,N_19296);
nor U20613 (N_20613,N_19525,N_18969);
nor U20614 (N_20614,N_16172,N_18635);
and U20615 (N_20615,N_16068,N_18607);
or U20616 (N_20616,N_16337,N_18937);
and U20617 (N_20617,N_16547,N_19979);
or U20618 (N_20618,N_17290,N_18721);
and U20619 (N_20619,N_15605,N_19270);
and U20620 (N_20620,N_19638,N_15454);
and U20621 (N_20621,N_16380,N_15003);
or U20622 (N_20622,N_18093,N_19857);
nand U20623 (N_20623,N_16320,N_15482);
nand U20624 (N_20624,N_15096,N_18716);
nand U20625 (N_20625,N_18980,N_18159);
and U20626 (N_20626,N_18977,N_17615);
nor U20627 (N_20627,N_16675,N_16822);
or U20628 (N_20628,N_17629,N_18480);
nor U20629 (N_20629,N_18521,N_15760);
nand U20630 (N_20630,N_17702,N_15806);
and U20631 (N_20631,N_19641,N_18774);
and U20632 (N_20632,N_15337,N_17591);
nand U20633 (N_20633,N_17085,N_19018);
or U20634 (N_20634,N_18991,N_19886);
nand U20635 (N_20635,N_15561,N_16930);
xor U20636 (N_20636,N_17802,N_18975);
nand U20637 (N_20637,N_17384,N_18535);
or U20638 (N_20638,N_16326,N_15442);
nand U20639 (N_20639,N_18927,N_16159);
xor U20640 (N_20640,N_15136,N_15418);
nor U20641 (N_20641,N_18992,N_16244);
or U20642 (N_20642,N_17900,N_18673);
nand U20643 (N_20643,N_16527,N_17127);
and U20644 (N_20644,N_15451,N_18313);
and U20645 (N_20645,N_16101,N_15631);
or U20646 (N_20646,N_16047,N_17034);
or U20647 (N_20647,N_16427,N_17675);
or U20648 (N_20648,N_18879,N_18443);
nand U20649 (N_20649,N_16449,N_15764);
nor U20650 (N_20650,N_16287,N_17006);
nor U20651 (N_20651,N_17770,N_16836);
or U20652 (N_20652,N_15942,N_18780);
and U20653 (N_20653,N_17330,N_19365);
nor U20654 (N_20654,N_16504,N_16064);
or U20655 (N_20655,N_16241,N_18273);
nor U20656 (N_20656,N_15049,N_18552);
and U20657 (N_20657,N_16233,N_18559);
nand U20658 (N_20658,N_15245,N_18434);
nand U20659 (N_20659,N_19239,N_17049);
nand U20660 (N_20660,N_17953,N_17069);
and U20661 (N_20661,N_19484,N_16537);
and U20662 (N_20662,N_16963,N_19190);
xor U20663 (N_20663,N_15335,N_15261);
or U20664 (N_20664,N_19375,N_15673);
nand U20665 (N_20665,N_16323,N_19939);
nand U20666 (N_20666,N_15017,N_18453);
or U20667 (N_20667,N_16868,N_15381);
or U20668 (N_20668,N_16209,N_18758);
or U20669 (N_20669,N_18342,N_18054);
nand U20670 (N_20670,N_19000,N_19736);
or U20671 (N_20671,N_18749,N_18570);
nor U20672 (N_20672,N_17261,N_18933);
nand U20673 (N_20673,N_17438,N_15130);
or U20674 (N_20674,N_19333,N_16798);
nor U20675 (N_20675,N_15948,N_15068);
nor U20676 (N_20676,N_17581,N_16282);
nand U20677 (N_20677,N_18471,N_18412);
nand U20678 (N_20678,N_19373,N_15579);
nand U20679 (N_20679,N_15708,N_18762);
or U20680 (N_20680,N_16686,N_19185);
nor U20681 (N_20681,N_16322,N_17705);
and U20682 (N_20682,N_19689,N_17776);
nand U20683 (N_20683,N_18994,N_15307);
nor U20684 (N_20684,N_16919,N_17946);
nor U20685 (N_20685,N_18297,N_19763);
nand U20686 (N_20686,N_15219,N_17457);
nor U20687 (N_20687,N_16202,N_18954);
nand U20688 (N_20688,N_15963,N_17421);
or U20689 (N_20689,N_15540,N_19086);
nand U20690 (N_20690,N_18359,N_17919);
nor U20691 (N_20691,N_19499,N_18549);
nand U20692 (N_20692,N_15023,N_15550);
nor U20693 (N_20693,N_19741,N_17759);
nand U20694 (N_20694,N_19976,N_18035);
xnor U20695 (N_20695,N_18818,N_15318);
xor U20696 (N_20696,N_17878,N_17061);
nor U20697 (N_20697,N_15375,N_19164);
nor U20698 (N_20698,N_17657,N_17439);
and U20699 (N_20699,N_18718,N_15811);
and U20700 (N_20700,N_18203,N_17222);
nand U20701 (N_20701,N_18280,N_15757);
and U20702 (N_20702,N_18421,N_15544);
nand U20703 (N_20703,N_17081,N_15678);
nor U20704 (N_20704,N_16913,N_18442);
nor U20705 (N_20705,N_19895,N_15163);
or U20706 (N_20706,N_16646,N_18490);
and U20707 (N_20707,N_16173,N_15061);
nor U20708 (N_20708,N_16492,N_19142);
nor U20709 (N_20709,N_16780,N_16450);
or U20710 (N_20710,N_15109,N_15406);
nand U20711 (N_20711,N_18956,N_19234);
and U20712 (N_20712,N_18079,N_16490);
and U20713 (N_20713,N_17077,N_16876);
or U20714 (N_20714,N_19210,N_15384);
nor U20715 (N_20715,N_18514,N_16863);
nand U20716 (N_20716,N_18742,N_19996);
and U20717 (N_20717,N_16753,N_16100);
and U20718 (N_20718,N_19266,N_15488);
nand U20719 (N_20719,N_15161,N_17648);
or U20720 (N_20720,N_17825,N_19274);
nand U20721 (N_20721,N_19868,N_17449);
nor U20722 (N_20722,N_16934,N_19826);
nor U20723 (N_20723,N_17269,N_19336);
and U20724 (N_20724,N_17325,N_15795);
and U20725 (N_20725,N_17103,N_17249);
and U20726 (N_20726,N_18197,N_17893);
and U20727 (N_20727,N_15259,N_17604);
or U20728 (N_20728,N_18830,N_17708);
or U20729 (N_20729,N_16343,N_15744);
nand U20730 (N_20730,N_15203,N_15458);
and U20731 (N_20731,N_18949,N_19970);
nor U20732 (N_20732,N_19754,N_17716);
and U20733 (N_20733,N_18941,N_19579);
nor U20734 (N_20734,N_19840,N_19110);
and U20735 (N_20735,N_17281,N_16629);
nor U20736 (N_20736,N_16222,N_18553);
nor U20737 (N_20737,N_19629,N_15886);
nor U20738 (N_20738,N_15698,N_16300);
or U20739 (N_20739,N_18857,N_17255);
nor U20740 (N_20740,N_16014,N_17392);
and U20741 (N_20741,N_15970,N_18504);
xor U20742 (N_20742,N_19307,N_16069);
and U20743 (N_20743,N_19471,N_17378);
or U20744 (N_20744,N_17057,N_18485);
nand U20745 (N_20745,N_15810,N_16853);
nand U20746 (N_20746,N_18267,N_15936);
nor U20747 (N_20747,N_19456,N_17419);
nor U20748 (N_20748,N_17105,N_18241);
xor U20749 (N_20749,N_19475,N_17285);
nand U20750 (N_20750,N_17954,N_16503);
and U20751 (N_20751,N_18488,N_15284);
or U20752 (N_20752,N_15427,N_16797);
and U20753 (N_20753,N_19801,N_17231);
and U20754 (N_20754,N_17158,N_19262);
nor U20755 (N_20755,N_17630,N_19256);
and U20756 (N_20756,N_17188,N_16262);
xor U20757 (N_20757,N_15857,N_15932);
and U20758 (N_20758,N_19264,N_18232);
and U20759 (N_20759,N_17416,N_18162);
nor U20760 (N_20760,N_15551,N_18662);
nor U20761 (N_20761,N_18905,N_17465);
and U20762 (N_20762,N_18292,N_19923);
nor U20763 (N_20763,N_17100,N_16977);
nor U20764 (N_20764,N_18172,N_17641);
nor U20765 (N_20765,N_17210,N_19523);
and U20766 (N_20766,N_17426,N_17172);
and U20767 (N_20767,N_17925,N_19151);
nor U20768 (N_20768,N_15069,N_16649);
xnor U20769 (N_20769,N_18855,N_15420);
nand U20770 (N_20770,N_18773,N_15891);
or U20771 (N_20771,N_19235,N_16857);
nor U20772 (N_20772,N_17537,N_15575);
nor U20773 (N_20773,N_15395,N_16428);
nor U20774 (N_20774,N_16530,N_18759);
and U20775 (N_20775,N_18064,N_18437);
nand U20776 (N_20776,N_19795,N_17437);
nand U20777 (N_20777,N_17114,N_18333);
or U20778 (N_20778,N_19705,N_15345);
nand U20779 (N_20779,N_19470,N_15371);
nand U20780 (N_20780,N_18403,N_17649);
nand U20781 (N_20781,N_16110,N_18406);
and U20782 (N_20782,N_18791,N_15967);
and U20783 (N_20783,N_18619,N_15581);
nand U20784 (N_20784,N_15390,N_18713);
and U20785 (N_20785,N_16989,N_15952);
nor U20786 (N_20786,N_19805,N_19971);
or U20787 (N_20787,N_15651,N_16414);
nand U20788 (N_20788,N_16502,N_19291);
or U20789 (N_20789,N_19707,N_15510);
nand U20790 (N_20790,N_17259,N_17955);
nand U20791 (N_20791,N_18509,N_16270);
and U20792 (N_20792,N_18580,N_16643);
or U20793 (N_20793,N_17005,N_17755);
nand U20794 (N_20794,N_19578,N_17171);
and U20795 (N_20795,N_19940,N_19891);
nor U20796 (N_20796,N_18356,N_17722);
or U20797 (N_20797,N_16894,N_19880);
nor U20798 (N_20798,N_19411,N_16289);
or U20799 (N_20799,N_17282,N_16707);
or U20800 (N_20800,N_18226,N_19894);
or U20801 (N_20801,N_16373,N_15535);
nand U20802 (N_20802,N_17420,N_15137);
xnor U20803 (N_20803,N_19721,N_16747);
nor U20804 (N_20804,N_19681,N_15732);
nor U20805 (N_20805,N_15640,N_17530);
nor U20806 (N_20806,N_16543,N_18743);
and U20807 (N_20807,N_17117,N_19211);
and U20808 (N_20808,N_17502,N_17343);
or U20809 (N_20809,N_19016,N_17864);
nor U20810 (N_20810,N_17942,N_15456);
nor U20811 (N_20811,N_15230,N_18279);
nor U20812 (N_20812,N_17974,N_16823);
nor U20813 (N_20813,N_18411,N_18384);
and U20814 (N_20814,N_15926,N_19751);
nand U20815 (N_20815,N_17949,N_16695);
and U20816 (N_20816,N_18243,N_15991);
nor U20817 (N_20817,N_19925,N_18971);
and U20818 (N_20818,N_16818,N_16265);
or U20819 (N_20819,N_16872,N_19224);
nand U20820 (N_20820,N_18587,N_18659);
nor U20821 (N_20821,N_19084,N_15714);
and U20822 (N_20822,N_16104,N_17731);
nor U20823 (N_20823,N_16580,N_16293);
or U20824 (N_20824,N_19282,N_16461);
or U20825 (N_20825,N_17036,N_18772);
and U20826 (N_20826,N_16859,N_18084);
and U20827 (N_20827,N_19524,N_16604);
nand U20828 (N_20828,N_15262,N_19155);
nand U20829 (N_20829,N_17317,N_15707);
and U20830 (N_20830,N_18298,N_16529);
and U20831 (N_20831,N_18816,N_19138);
and U20832 (N_20832,N_19562,N_15412);
nand U20833 (N_20833,N_17371,N_19316);
xor U20834 (N_20834,N_16524,N_18935);
and U20835 (N_20835,N_19920,N_18180);
nand U20836 (N_20836,N_16910,N_16572);
nor U20837 (N_20837,N_15862,N_19822);
nor U20838 (N_20838,N_15552,N_19810);
xor U20839 (N_20839,N_16335,N_19318);
and U20840 (N_20840,N_17610,N_16738);
nand U20841 (N_20841,N_16102,N_16290);
nor U20842 (N_20842,N_16467,N_16054);
or U20843 (N_20843,N_16664,N_17789);
and U20844 (N_20844,N_16672,N_15951);
and U20845 (N_20845,N_16049,N_18806);
nor U20846 (N_20846,N_15517,N_15874);
or U20847 (N_20847,N_18067,N_15054);
nor U20848 (N_20848,N_15878,N_19399);
nor U20849 (N_20849,N_15689,N_15546);
nor U20850 (N_20850,N_16256,N_15409);
or U20851 (N_20851,N_18925,N_15431);
nand U20852 (N_20852,N_18810,N_17101);
xnor U20853 (N_20853,N_16133,N_17351);
and U20854 (N_20854,N_18294,N_17894);
and U20855 (N_20855,N_15666,N_15095);
nand U20856 (N_20856,N_17522,N_15976);
and U20857 (N_20857,N_17607,N_18860);
xnor U20858 (N_20858,N_19604,N_16684);
nor U20859 (N_20859,N_15308,N_17353);
nor U20860 (N_20860,N_18011,N_17704);
nor U20861 (N_20861,N_15208,N_18601);
or U20862 (N_20862,N_17749,N_18456);
nand U20863 (N_20863,N_16677,N_15116);
and U20864 (N_20864,N_18543,N_16353);
or U20865 (N_20865,N_18502,N_19010);
or U20866 (N_20866,N_17297,N_16642);
nand U20867 (N_20867,N_18641,N_15310);
nor U20868 (N_20868,N_16508,N_19642);
nand U20869 (N_20869,N_15953,N_18515);
nand U20870 (N_20870,N_18873,N_19443);
and U20871 (N_20871,N_18551,N_15816);
nor U20872 (N_20872,N_17023,N_19616);
nand U20873 (N_20873,N_16505,N_16789);
and U20874 (N_20874,N_15762,N_18366);
and U20875 (N_20875,N_18717,N_17186);
and U20876 (N_20876,N_16103,N_19167);
nand U20877 (N_20877,N_19596,N_15875);
nor U20878 (N_20878,N_19122,N_17276);
or U20879 (N_20879,N_19676,N_19196);
xor U20880 (N_20880,N_19764,N_16117);
and U20881 (N_20881,N_16927,N_16837);
or U20882 (N_20882,N_18817,N_18558);
nand U20883 (N_20883,N_16271,N_19130);
nor U20884 (N_20884,N_19065,N_15251);
nor U20885 (N_20885,N_18122,N_16581);
nor U20886 (N_20886,N_18407,N_18014);
or U20887 (N_20887,N_19163,N_15800);
nor U20888 (N_20888,N_17928,N_18301);
nand U20889 (N_20889,N_17790,N_19654);
nand U20890 (N_20890,N_15021,N_16273);
and U20891 (N_20891,N_16549,N_19962);
or U20892 (N_20892,N_15104,N_16760);
nor U20893 (N_20893,N_19221,N_18588);
and U20894 (N_20894,N_15453,N_18231);
nor U20895 (N_20895,N_16783,N_17839);
nand U20896 (N_20896,N_17857,N_16924);
or U20897 (N_20897,N_19012,N_19035);
and U20898 (N_20898,N_15832,N_17466);
and U20899 (N_20899,N_15912,N_19598);
nor U20900 (N_20900,N_19267,N_15662);
and U20901 (N_20901,N_16958,N_15303);
nand U20902 (N_20902,N_19637,N_17807);
nor U20903 (N_20903,N_19796,N_16182);
nor U20904 (N_20904,N_18026,N_15241);
or U20905 (N_20905,N_19774,N_18170);
xnor U20906 (N_20906,N_17443,N_19783);
or U20907 (N_20907,N_18959,N_17701);
and U20908 (N_20908,N_19469,N_19882);
and U20909 (N_20909,N_19734,N_19448);
or U20910 (N_20910,N_16705,N_19406);
or U20911 (N_20911,N_15661,N_18389);
or U20912 (N_20912,N_19577,N_17080);
nor U20913 (N_20913,N_16525,N_17076);
and U20914 (N_20914,N_17544,N_15503);
or U20915 (N_20915,N_19309,N_19424);
or U20916 (N_20916,N_15740,N_17968);
nor U20917 (N_20917,N_15660,N_16591);
nand U20918 (N_20918,N_18417,N_15809);
or U20919 (N_20919,N_17688,N_19968);
or U20920 (N_20920,N_18123,N_19473);
nand U20921 (N_20921,N_18705,N_17777);
nand U20922 (N_20922,N_17021,N_18567);
nand U20923 (N_20923,N_15413,N_15917);
nand U20924 (N_20924,N_16540,N_18737);
or U20925 (N_20925,N_15754,N_17039);
nor U20926 (N_20926,N_19350,N_16548);
or U20927 (N_20927,N_16253,N_16935);
and U20928 (N_20928,N_18196,N_16696);
nor U20929 (N_20929,N_19935,N_19085);
and U20930 (N_20930,N_17822,N_16023);
or U20931 (N_20931,N_15135,N_17450);
nand U20932 (N_20932,N_15958,N_15944);
and U20933 (N_20933,N_18399,N_19104);
and U20934 (N_20934,N_16660,N_16617);
or U20935 (N_20935,N_15000,N_18141);
nand U20936 (N_20936,N_17837,N_17289);
xnor U20937 (N_20937,N_16228,N_17961);
or U20938 (N_20938,N_19490,N_17093);
nand U20939 (N_20939,N_18130,N_15798);
or U20940 (N_20940,N_16563,N_18544);
nand U20941 (N_20941,N_16557,N_15176);
and U20942 (N_20942,N_18099,N_16345);
and U20943 (N_20943,N_15781,N_17234);
nor U20944 (N_20944,N_18576,N_15702);
nor U20945 (N_20945,N_16926,N_18120);
nor U20946 (N_20946,N_19732,N_17089);
nand U20947 (N_20947,N_17215,N_15372);
nand U20948 (N_20948,N_15044,N_16971);
nor U20949 (N_20949,N_16210,N_15885);
nor U20950 (N_20950,N_17302,N_18021);
nor U20951 (N_20951,N_18875,N_18486);
nor U20952 (N_20952,N_15590,N_19344);
nor U20953 (N_20953,N_17515,N_15294);
nor U20954 (N_20954,N_15750,N_17983);
nand U20955 (N_20955,N_16232,N_16715);
nor U20956 (N_20956,N_16712,N_19413);
nor U20957 (N_20957,N_19205,N_16980);
nand U20958 (N_20958,N_15824,N_17969);
and U20959 (N_20959,N_19114,N_19203);
nand U20960 (N_20960,N_19218,N_18233);
or U20961 (N_20961,N_15074,N_16688);
nand U20962 (N_20962,N_16059,N_18837);
nand U20963 (N_20963,N_15220,N_19557);
nand U20964 (N_20964,N_18564,N_16305);
nor U20965 (N_20965,N_18996,N_16294);
nand U20966 (N_20966,N_15934,N_17873);
nand U20967 (N_20967,N_19043,N_19392);
nand U20968 (N_20968,N_17300,N_18880);
and U20969 (N_20969,N_19222,N_18917);
nand U20970 (N_20970,N_15898,N_15649);
or U20971 (N_20971,N_15389,N_16328);
nor U20972 (N_20972,N_18785,N_17038);
nor U20973 (N_20973,N_16559,N_17063);
nor U20974 (N_20974,N_17113,N_17869);
nor U20975 (N_20975,N_19566,N_18107);
and U20976 (N_20976,N_18765,N_15256);
or U20977 (N_20977,N_17899,N_18685);
or U20978 (N_20978,N_17403,N_16396);
and U20979 (N_20979,N_15572,N_19599);
nand U20980 (N_20980,N_17578,N_18931);
nor U20981 (N_20981,N_15747,N_17247);
nand U20982 (N_20982,N_19283,N_15518);
nor U20983 (N_20983,N_18277,N_17339);
nand U20984 (N_20984,N_16471,N_16240);
and U20985 (N_20985,N_19966,N_15704);
or U20986 (N_20986,N_16463,N_15679);
or U20987 (N_20987,N_16473,N_15315);
or U20988 (N_20988,N_19078,N_15739);
and U20989 (N_20989,N_16972,N_15984);
nor U20990 (N_20990,N_15994,N_17891);
and U20991 (N_20991,N_15899,N_18376);
nor U20992 (N_20992,N_16153,N_16805);
nand U20993 (N_20993,N_19213,N_15316);
xnor U20994 (N_20994,N_17943,N_18229);
and U20995 (N_20995,N_16803,N_16476);
or U20996 (N_20996,N_18302,N_17496);
and U20997 (N_20997,N_19464,N_18028);
nand U20998 (N_20998,N_19639,N_17441);
and U20999 (N_20999,N_16754,N_15960);
xnor U21000 (N_21000,N_16114,N_17609);
nor U21001 (N_21001,N_16653,N_16565);
nand U21002 (N_21002,N_18378,N_15922);
nor U21003 (N_21003,N_19915,N_17052);
nand U21004 (N_21004,N_17332,N_17298);
and U21005 (N_21005,N_19714,N_15751);
nand U21006 (N_21006,N_17047,N_19173);
and U21007 (N_21007,N_16802,N_19457);
nand U21008 (N_21008,N_19664,N_18622);
nor U21009 (N_21009,N_17528,N_15228);
and U21010 (N_21010,N_16230,N_16309);
and U21011 (N_21011,N_16614,N_19511);
nand U21012 (N_21012,N_19761,N_15332);
nand U21013 (N_21013,N_16544,N_19993);
nand U21014 (N_21014,N_17611,N_18185);
nand U21015 (N_21015,N_17835,N_16356);
or U21016 (N_21016,N_18074,N_15077);
nand U21017 (N_21017,N_16949,N_17831);
nand U21018 (N_21018,N_18240,N_16090);
xnor U21019 (N_21019,N_16272,N_19184);
xor U21020 (N_21020,N_16568,N_19459);
nand U21021 (N_21021,N_19640,N_16742);
nor U21022 (N_21022,N_16236,N_18154);
and U21023 (N_21023,N_17752,N_17315);
nor U21024 (N_21024,N_16861,N_18080);
nand U21025 (N_21025,N_19332,N_18727);
nand U21026 (N_21026,N_19997,N_17214);
nand U21027 (N_21027,N_16499,N_16941);
and U21028 (N_21028,N_19697,N_18066);
and U21029 (N_21029,N_15445,N_16816);
nor U21030 (N_21030,N_15040,N_15770);
and U21031 (N_21031,N_17990,N_15013);
nor U21032 (N_21032,N_16534,N_19744);
or U21033 (N_21033,N_17663,N_16028);
nor U21034 (N_21034,N_16718,N_19933);
and U21035 (N_21035,N_17858,N_17341);
and U21036 (N_21036,N_16274,N_16645);
nand U21037 (N_21037,N_15664,N_17762);
nor U21038 (N_21038,N_19229,N_19586);
or U21039 (N_21039,N_18354,N_16207);
or U21040 (N_21040,N_17447,N_15659);
and U21041 (N_21041,N_15326,N_17795);
xnor U21042 (N_21042,N_19433,N_17408);
nor U21043 (N_21043,N_18049,N_16929);
nor U21044 (N_21044,N_17792,N_16955);
nand U21045 (N_21045,N_18004,N_19227);
and U21046 (N_21046,N_15090,N_18426);
xnor U21047 (N_21047,N_16609,N_16487);
xnor U21048 (N_21048,N_19472,N_19837);
and U21049 (N_21049,N_18757,N_17184);
or U21050 (N_21050,N_19606,N_15378);
nand U21051 (N_21051,N_15346,N_17401);
and U21052 (N_21052,N_16466,N_16851);
or U21053 (N_21053,N_18472,N_19951);
and U21054 (N_21054,N_19342,N_15577);
or U21055 (N_21055,N_16900,N_16418);
and U21056 (N_21056,N_18072,N_15522);
or U21057 (N_21057,N_16765,N_17235);
or U21058 (N_21058,N_17772,N_18866);
and U21059 (N_21059,N_15240,N_15892);
nand U21060 (N_21060,N_17783,N_16231);
or U21061 (N_21061,N_18266,N_15475);
and U21062 (N_21062,N_19374,N_18435);
or U21063 (N_21063,N_19559,N_15753);
or U21064 (N_21064,N_16458,N_18171);
or U21065 (N_21065,N_15796,N_18181);
nand U21066 (N_21066,N_17645,N_17381);
and U21067 (N_21067,N_17303,N_15434);
nor U21068 (N_21068,N_19703,N_19400);
nor U21069 (N_21069,N_15663,N_17070);
and U21070 (N_21070,N_16895,N_17508);
nand U21071 (N_21071,N_16191,N_19028);
and U21072 (N_21072,N_17352,N_17721);
and U21073 (N_21073,N_17189,N_16826);
nor U21074 (N_21074,N_18455,N_17852);
xnor U21075 (N_21075,N_15855,N_15610);
and U21076 (N_21076,N_17316,N_15306);
nor U21077 (N_21077,N_17484,N_16734);
nand U21078 (N_21078,N_18752,N_15391);
nor U21079 (N_21079,N_18645,N_15035);
nor U21080 (N_21080,N_19295,N_15009);
nor U21081 (N_21081,N_16983,N_17424);
nand U21082 (N_21082,N_15743,N_18397);
nand U21083 (N_21083,N_18328,N_17058);
and U21084 (N_21084,N_15969,N_19973);
nor U21085 (N_21085,N_15022,N_17182);
nand U21086 (N_21086,N_17490,N_17929);
nor U21087 (N_21087,N_18070,N_15432);
or U21088 (N_21088,N_18584,N_16937);
xnor U21089 (N_21089,N_15103,N_16251);
or U21090 (N_21090,N_15290,N_17327);
or U21091 (N_21091,N_18065,N_19969);
and U21092 (N_21092,N_19299,N_17246);
and U21093 (N_21093,N_16279,N_18616);
or U21094 (N_21094,N_19852,N_19911);
or U21095 (N_21095,N_18871,N_15302);
or U21096 (N_21096,N_17664,N_17506);
or U21097 (N_21097,N_18043,N_15243);
nand U21098 (N_21098,N_19458,N_16154);
and U21099 (N_21099,N_18799,N_19040);
and U21100 (N_21100,N_15900,N_19618);
and U21101 (N_21101,N_19936,N_16457);
or U21102 (N_21102,N_15975,N_19879);
nor U21103 (N_21103,N_17608,N_16113);
or U21104 (N_21104,N_18542,N_16012);
nor U21105 (N_21105,N_15177,N_18429);
or U21106 (N_21106,N_18278,N_18651);
or U21107 (N_21107,N_16390,N_19311);
or U21108 (N_21108,N_17950,N_17396);
nand U21109 (N_21109,N_18225,N_19001);
and U21110 (N_21110,N_18734,N_16959);
and U21111 (N_21111,N_19869,N_18573);
or U21112 (N_21112,N_17094,N_15901);
nor U21113 (N_21113,N_19462,N_19526);
and U21114 (N_21114,N_19804,N_18620);
and U21115 (N_21115,N_18919,N_17690);
nand U21116 (N_21116,N_18493,N_16743);
and U21117 (N_21117,N_17715,N_17801);
or U21118 (N_21118,N_15929,N_16331);
nand U21119 (N_21119,N_19127,N_16887);
nor U21120 (N_21120,N_15298,N_19378);
and U21121 (N_21121,N_17639,N_19902);
or U21122 (N_21122,N_15935,N_16254);
and U21123 (N_21123,N_15410,N_16532);
nor U21124 (N_21124,N_15169,N_15609);
and U21125 (N_21125,N_15993,N_15499);
or U21126 (N_21126,N_17213,N_16858);
nand U21127 (N_21127,N_16605,N_16034);
nor U21128 (N_21128,N_17075,N_17733);
nor U21129 (N_21129,N_18052,N_17897);
nor U21130 (N_21130,N_18338,N_18450);
and U21131 (N_21131,N_19076,N_15102);
nor U21132 (N_21132,N_19884,N_18940);
and U21133 (N_21133,N_17574,N_18224);
and U21134 (N_21134,N_16701,N_16037);
or U21135 (N_21135,N_18778,N_19489);
xor U21136 (N_21136,N_16121,N_15042);
and U21137 (N_21137,N_15675,N_17904);
nor U21138 (N_21138,N_18227,N_18097);
or U21139 (N_21139,N_18219,N_18653);
nor U21140 (N_21140,N_19521,N_17092);
nor U21141 (N_21141,N_15016,N_18051);
and U21142 (N_21142,N_18585,N_18600);
nor U21143 (N_21143,N_15742,N_18827);
nor U21144 (N_21144,N_19135,N_19892);
or U21145 (N_21145,N_19083,N_18150);
and U21146 (N_21146,N_16880,N_17273);
nor U21147 (N_21147,N_15484,N_19108);
nor U21148 (N_21148,N_15041,N_16870);
and U21149 (N_21149,N_19990,N_17941);
or U21150 (N_21150,N_16800,N_19785);
nand U21151 (N_21151,N_19507,N_18881);
and U21152 (N_21152,N_19829,N_17994);
nand U21153 (N_21153,N_16500,N_17692);
and U21154 (N_21154,N_19003,N_19696);
or U21155 (N_21155,N_15127,N_19113);
or U21156 (N_21156,N_18269,N_17678);
and U21157 (N_21157,N_15062,N_18574);
or U21158 (N_21158,N_16085,N_15078);
nor U21159 (N_21159,N_15624,N_19769);
nand U21160 (N_21160,N_17248,N_16790);
or U21161 (N_21161,N_17892,N_15291);
nor U21162 (N_21162,N_19595,N_19198);
and U21163 (N_21163,N_18179,N_19099);
nand U21164 (N_21164,N_16091,N_16378);
nand U21165 (N_21165,N_19050,N_19174);
and U21166 (N_21166,N_16722,N_15706);
nand U21167 (N_21167,N_17525,N_15968);
or U21168 (N_21168,N_16269,N_17395);
nor U21169 (N_21169,N_16893,N_16127);
or U21170 (N_21170,N_18874,N_19963);
nand U21171 (N_21171,N_18129,N_15106);
nor U21172 (N_21172,N_17226,N_17793);
nor U21173 (N_21173,N_17201,N_17193);
or U21174 (N_21174,N_17697,N_15670);
nand U21175 (N_21175,N_19501,N_19087);
nand U21176 (N_21176,N_15180,N_16220);
or U21177 (N_21177,N_19766,N_19896);
nor U21178 (N_21178,N_17930,N_18482);
nor U21179 (N_21179,N_18125,N_18466);
or U21180 (N_21180,N_16681,N_17035);
nor U21181 (N_21181,N_16731,N_19546);
or U21182 (N_21182,N_18865,N_19709);
and U21183 (N_21183,N_15211,N_18981);
nor U21184 (N_21184,N_18008,N_16554);
nand U21185 (N_21185,N_17670,N_17635);
nand U21186 (N_21186,N_15138,N_17425);
or U21187 (N_21187,N_18524,N_18119);
xor U21188 (N_21188,N_17204,N_18793);
or U21189 (N_21189,N_15489,N_16693);
nand U21190 (N_21190,N_15008,N_19739);
nor U21191 (N_21191,N_18661,N_16268);
nand U21192 (N_21192,N_19981,N_18541);
nand U21193 (N_21193,N_18805,N_16583);
and U21194 (N_21194,N_17914,N_17996);
and U21195 (N_21195,N_17160,N_15480);
nand U21196 (N_21196,N_15450,N_18803);
and U21197 (N_21197,N_18859,N_16176);
nand U21198 (N_21198,N_15741,N_15914);
nand U21199 (N_21199,N_17592,N_15910);
and U21200 (N_21200,N_15481,N_15657);
or U21201 (N_21201,N_17136,N_17656);
or U21202 (N_21202,N_16045,N_18730);
nor U21203 (N_21203,N_16423,N_19479);
or U21204 (N_21204,N_17399,N_19207);
nand U21205 (N_21205,N_18167,N_16879);
and U21206 (N_21206,N_19032,N_16536);
nand U21207 (N_21207,N_18110,N_19247);
nand U21208 (N_21208,N_18582,N_19713);
or U21209 (N_21209,N_15668,N_15873);
and U21210 (N_21210,N_17760,N_15237);
and U21211 (N_21211,N_17257,N_16756);
nor U21212 (N_21212,N_15772,N_16985);
nor U21213 (N_21213,N_15906,N_15126);
nand U21214 (N_21214,N_17493,N_18862);
and U21215 (N_21215,N_17662,N_16809);
or U21216 (N_21216,N_18614,N_15902);
or U21217 (N_21217,N_19129,N_18492);
nor U21218 (N_21218,N_17320,N_15099);
nor U21219 (N_21219,N_16430,N_16786);
nand U21220 (N_21220,N_17723,N_17161);
nand U21221 (N_21221,N_17998,N_17896);
or U21222 (N_21222,N_19498,N_19643);
nand U21223 (N_21223,N_19539,N_15583);
nand U21224 (N_21224,N_17157,N_16634);
nand U21225 (N_21225,N_18688,N_15568);
nor U21226 (N_21226,N_16119,N_16346);
nand U21227 (N_21227,N_16626,N_17916);
nand U21228 (N_21228,N_16493,N_16556);
and U21229 (N_21229,N_16806,N_15045);
or U21230 (N_21230,N_16914,N_17291);
or U21231 (N_21231,N_18300,N_16922);
xor U21232 (N_21232,N_16481,N_19193);
and U21233 (N_21233,N_15685,N_17785);
nand U21234 (N_21234,N_18475,N_16689);
or U21235 (N_21235,N_15071,N_19395);
or U21236 (N_21236,N_16118,N_16513);
nand U21237 (N_21237,N_19088,N_19260);
nand U21238 (N_21238,N_18986,N_19635);
or U21239 (N_21239,N_16616,N_18577);
and U21240 (N_21240,N_18728,N_15030);
nor U21241 (N_21241,N_18069,N_19118);
nand U21242 (N_21242,N_15918,N_16446);
and U21243 (N_21243,N_17254,N_17388);
or U21244 (N_21244,N_18861,N_19728);
nand U21245 (N_21245,N_16898,N_17333);
or U21246 (N_21246,N_15353,N_16752);
nor U21247 (N_21247,N_15965,N_18507);
nand U21248 (N_21248,N_16939,N_18223);
or U21249 (N_21249,N_17053,N_16597);
xnor U21250 (N_21250,N_16825,N_19182);
nor U21251 (N_21251,N_16763,N_17531);
or U21252 (N_21252,N_19440,N_18712);
and U21253 (N_21253,N_18900,N_19090);
and U21254 (N_21254,N_16180,N_18583);
or U21255 (N_21255,N_19959,N_16399);
nor U21256 (N_21256,N_18377,N_15347);
nor U21257 (N_21257,N_17709,N_15257);
nand U21258 (N_21258,N_18168,N_15915);
nor U21259 (N_21259,N_19723,N_19364);
nor U21260 (N_21260,N_19802,N_17874);
and U21261 (N_21261,N_17582,N_19463);
nand U21262 (N_21262,N_19771,N_19608);
nand U21263 (N_21263,N_19394,N_19428);
and U21264 (N_21264,N_16043,N_15114);
nor U21265 (N_21265,N_16661,N_16904);
nor U21266 (N_21266,N_18315,N_18548);
or U21267 (N_21267,N_17566,N_16659);
and U21268 (N_21268,N_17568,N_19558);
and U21269 (N_21269,N_15401,N_16033);
nand U21270 (N_21270,N_15723,N_17389);
nor U21271 (N_21271,N_15506,N_17130);
and U21272 (N_21272,N_17126,N_17397);
and U21273 (N_21273,N_15674,N_17918);
nand U21274 (N_21274,N_17819,N_17295);
and U21275 (N_21275,N_17220,N_19063);
nor U21276 (N_21276,N_18776,N_19263);
and U21277 (N_21277,N_15212,N_16969);
and U21278 (N_21278,N_16156,N_19856);
and U21279 (N_21279,N_18390,N_19995);
nor U21280 (N_21280,N_19157,N_17805);
or U21281 (N_21281,N_18281,N_15856);
or U21282 (N_21282,N_17434,N_17717);
or U21283 (N_21283,N_17000,N_18958);
nor U21284 (N_21284,N_15826,N_18767);
nand U21285 (N_21285,N_17987,N_17347);
and U21286 (N_21286,N_16123,N_15903);
or U21287 (N_21287,N_16376,N_16775);
nor U21288 (N_21288,N_17711,N_18844);
nand U21289 (N_21289,N_15422,N_19432);
or U21290 (N_21290,N_17718,N_18461);
or U21291 (N_21291,N_17583,N_17356);
and U21292 (N_21292,N_17550,N_16951);
or U21293 (N_21293,N_18230,N_19657);
nor U21294 (N_21294,N_16030,N_16576);
xnor U21295 (N_21295,N_18314,N_16946);
nor U21296 (N_21296,N_17626,N_17120);
or U21297 (N_21297,N_18922,N_16593);
or U21298 (N_21298,N_18921,N_15031);
and U21299 (N_21299,N_19371,N_18000);
and U21300 (N_21300,N_19494,N_19176);
xor U21301 (N_21301,N_17121,N_19743);
or U21302 (N_21302,N_15825,N_17939);
or U21303 (N_21303,N_15289,N_19753);
nor U21304 (N_21304,N_16257,N_18656);
nand U21305 (N_21305,N_17194,N_17879);
and U21306 (N_21306,N_18789,N_16214);
nand U21307 (N_21307,N_19628,N_15046);
or U21308 (N_21308,N_15331,N_16389);
or U21309 (N_21309,N_16650,N_16938);
and U21310 (N_21310,N_15015,N_15467);
xnor U21311 (N_21311,N_19735,N_17765);
nor U21312 (N_21312,N_16566,N_18477);
and U21313 (N_21313,N_18208,N_16098);
nand U21314 (N_21314,N_17017,N_15726);
or U21315 (N_21315,N_15617,N_16234);
and U21316 (N_21316,N_16830,N_16770);
xnor U21317 (N_21317,N_19171,N_17367);
nor U21318 (N_21318,N_15293,N_16570);
nand U21319 (N_21319,N_15435,N_16444);
or U21320 (N_21320,N_17242,N_15837);
and U21321 (N_21321,N_15955,N_19958);
xnor U21322 (N_21322,N_17125,N_16434);
nand U21323 (N_21323,N_16306,N_15292);
nor U21324 (N_21324,N_15641,N_16395);
nor U21325 (N_21325,N_16384,N_19513);
nor U21326 (N_21326,N_17923,N_17511);
nor U21327 (N_21327,N_15339,N_17409);
nand U21328 (N_21328,N_16052,N_16031);
nand U21329 (N_21329,N_16854,N_16187);
nand U21330 (N_21330,N_19482,N_15513);
nand U21331 (N_21331,N_18870,N_18942);
nor U21332 (N_21332,N_15311,N_18030);
nand U21333 (N_21333,N_16749,N_16071);
and U21334 (N_21334,N_16990,N_15314);
nand U21335 (N_21335,N_18117,N_16470);
xnor U21336 (N_21336,N_15498,N_16072);
xnor U21337 (N_21337,N_15928,N_16086);
nor U21338 (N_21338,N_16700,N_17456);
nor U21339 (N_21339,N_15710,N_19854);
or U21340 (N_21340,N_15817,N_15055);
or U21341 (N_21341,N_19622,N_19393);
xnor U21342 (N_21342,N_15697,N_19495);
nand U21343 (N_21343,N_17267,N_16122);
nor U21344 (N_21344,N_15014,N_19636);
and U21345 (N_21345,N_19465,N_15635);
nand U21346 (N_21346,N_18670,N_19778);
nor U21347 (N_21347,N_19047,N_15026);
nor U21348 (N_21348,N_19814,N_16004);
or U21349 (N_21349,N_15142,N_18596);
nand U21350 (N_21350,N_18415,N_19354);
nand U21351 (N_21351,N_16709,N_18957);
nor U21352 (N_21352,N_15515,N_15554);
nor U21353 (N_21353,N_19678,N_19860);
or U21354 (N_21354,N_15534,N_19821);
nor U21355 (N_21355,N_17132,N_17055);
or U21356 (N_21356,N_16497,N_19340);
nand U21357 (N_21357,N_18113,N_18370);
or U21358 (N_21358,N_17813,N_16832);
or U21359 (N_21359,N_19550,N_19631);
nand U21360 (N_21360,N_17072,N_16339);
nand U21361 (N_21361,N_19561,N_15407);
nor U21362 (N_21362,N_16845,N_19765);
or U21363 (N_21363,N_16865,N_16736);
nand U21364 (N_21364,N_15399,N_17617);
nand U21365 (N_21365,N_18513,N_15134);
or U21366 (N_21366,N_15446,N_18111);
or U21367 (N_21367,N_15511,N_18624);
or U21368 (N_21368,N_19055,N_19593);
nand U21369 (N_21369,N_18358,N_18489);
and U21370 (N_21370,N_15637,N_17562);
nor U21371 (N_21371,N_16456,N_16828);
or U21372 (N_21372,N_17203,N_16469);
and U21373 (N_21373,N_15123,N_17025);
or U21374 (N_21374,N_16885,N_17823);
and U21375 (N_21375,N_18715,N_19790);
nor U21376 (N_21376,N_17595,N_17472);
nor U21377 (N_21377,N_19798,N_18706);
nand U21378 (N_21378,N_19924,N_17365);
nor U21379 (N_21379,N_17719,N_17278);
nand U21380 (N_21380,N_16586,N_15221);
xor U21381 (N_21381,N_15323,N_18611);
nor U21382 (N_21382,N_19451,N_15210);
nor U21383 (N_21383,N_18305,N_16075);
nor U21384 (N_21384,N_17944,N_17305);
nand U21385 (N_21385,N_19509,N_15089);
nand U21386 (N_21386,N_16439,N_18201);
nor U21387 (N_21387,N_18571,N_17001);
nor U21388 (N_21388,N_18010,N_18568);
or U21389 (N_21389,N_19359,N_18388);
or U21390 (N_21390,N_18188,N_15440);
nand U21391 (N_21391,N_19777,N_16347);
nor U21392 (N_21392,N_16200,N_19571);
or U21393 (N_21393,N_17454,N_16648);
nand U21394 (N_21394,N_17766,N_18291);
nor U21395 (N_21395,N_15394,N_17543);
nor U21396 (N_21396,N_16438,N_17841);
nand U21397 (N_21397,N_15731,N_18032);
nor U21398 (N_21398,N_16338,N_17173);
or U21399 (N_21399,N_19865,N_15091);
or U21400 (N_21400,N_19549,N_17593);
or U21401 (N_21401,N_16923,N_18345);
or U21402 (N_21402,N_16909,N_16658);
and U21403 (N_21403,N_15531,N_19789);
nand U21404 (N_21404,N_16982,N_15669);
and U21405 (N_21405,N_17576,N_18391);
or U21406 (N_21406,N_18707,N_15989);
or U21407 (N_21407,N_18536,N_16281);
nand U21408 (N_21408,N_18760,N_18187);
nor U21409 (N_21409,N_16814,N_19831);
nor U21410 (N_21410,N_17653,N_18892);
nand U21411 (N_21411,N_17786,N_17606);
and U21412 (N_21412,N_19162,N_17195);
nor U21413 (N_21413,N_19942,N_16966);
and U21414 (N_21414,N_19410,N_19153);
or U21415 (N_21415,N_17948,N_15182);
nand U21416 (N_21416,N_18452,N_17268);
nor U21417 (N_21417,N_19615,N_18629);
or U21418 (N_21418,N_17684,N_15269);
nor U21419 (N_21419,N_18650,N_19505);
or U21420 (N_21420,N_17224,N_16724);
nor U21421 (N_21421,N_17850,N_16138);
nand U21422 (N_21422,N_17013,N_16723);
nand U21423 (N_21423,N_18901,N_15735);
nor U21424 (N_21424,N_16370,N_16226);
or U21425 (N_21425,N_15361,N_15278);
nor U21426 (N_21426,N_16592,N_17738);
nor U21427 (N_21427,N_17861,N_18349);
nand U21428 (N_21428,N_19115,N_17907);
nand U21429 (N_21429,N_15613,N_18148);
nand U21430 (N_21430,N_15053,N_18083);
and U21431 (N_21431,N_17411,N_18418);
nor U21432 (N_21432,N_16089,N_19404);
nand U21433 (N_21433,N_16878,N_18098);
nor U21434 (N_21434,N_18676,N_18669);
or U21435 (N_21435,N_19686,N_19659);
or U21436 (N_21436,N_17433,N_19057);
or U21437 (N_21437,N_17032,N_18322);
or U21438 (N_21438,N_19382,N_16264);
nor U21439 (N_21439,N_15505,N_19019);
nor U21440 (N_21440,N_18491,N_17507);
nand U21441 (N_21441,N_15853,N_18679);
nor U21442 (N_21442,N_18813,N_17323);
and U21443 (N_21443,N_19569,N_19327);
and U21444 (N_21444,N_17856,N_15827);
nor U21445 (N_21445,N_15636,N_16482);
or U21446 (N_21446,N_19603,N_17398);
nor U21447 (N_21447,N_16673,N_17250);
or U21448 (N_21448,N_15919,N_17045);
and U21449 (N_21449,N_17993,N_17650);
nand U21450 (N_21450,N_19772,N_15769);
or U21451 (N_21451,N_15455,N_18076);
or U21452 (N_21452,N_18446,N_19724);
or U21453 (N_21453,N_19974,N_16386);
xor U21454 (N_21454,N_15473,N_18623);
nand U21455 (N_21455,N_17972,N_19054);
nor U21456 (N_21456,N_17102,N_16011);
and U21457 (N_21457,N_16680,N_17181);
nor U21458 (N_21458,N_16327,N_17885);
nor U21459 (N_21459,N_15198,N_18674);
and U21460 (N_21460,N_19688,N_19278);
nand U21461 (N_21461,N_16954,N_16671);
nor U21462 (N_21462,N_18714,N_19120);
and U21463 (N_21463,N_19133,N_17027);
or U21464 (N_21464,N_15355,N_18924);
or U21465 (N_21465,N_15153,N_16514);
nand U21466 (N_21466,N_15525,N_17555);
or U21467 (N_21467,N_17933,N_17199);
or U21468 (N_21468,N_19623,N_17019);
nand U21469 (N_21469,N_15075,N_17672);
and U21470 (N_21470,N_17977,N_15148);
and U21471 (N_21471,N_15029,N_19666);
nand U21472 (N_21472,N_18250,N_18973);
nor U21473 (N_21473,N_15950,N_16489);
nand U21474 (N_21474,N_18510,N_19453);
and U21475 (N_21475,N_17787,N_19477);
or U21476 (N_21476,N_17442,N_19890);
nand U21477 (N_21477,N_15962,N_15327);
and U21478 (N_21478,N_17633,N_15005);
and U21479 (N_21479,N_15946,N_17980);
and U21480 (N_21480,N_17066,N_15775);
and U21481 (N_21481,N_19956,N_16625);
nor U21482 (N_21482,N_16729,N_16917);
and U21483 (N_21483,N_18741,N_18207);
and U21484 (N_21484,N_15235,N_16333);
and U21485 (N_21485,N_19315,N_18997);
nand U21486 (N_21486,N_15073,N_18288);
nand U21487 (N_21487,N_18101,N_19722);
and U21488 (N_21488,N_18381,N_16124);
nor U21489 (N_21489,N_18952,N_17978);
and U21490 (N_21490,N_15680,N_17636);
nor U21491 (N_21491,N_18606,N_18346);
xor U21492 (N_21492,N_18968,N_18105);
nand U21493 (N_21493,N_19111,N_15643);
and U21494 (N_21494,N_18740,N_18321);
nor U21495 (N_21495,N_18242,N_18724);
nand U21496 (N_21496,N_18678,N_17910);
nand U21497 (N_21497,N_19450,N_16258);
nor U21498 (N_21498,N_17227,N_15387);
nand U21499 (N_21499,N_17957,N_18387);
and U21500 (N_21500,N_16611,N_17794);
nand U21501 (N_21501,N_19244,N_16163);
or U21502 (N_21502,N_17504,N_17665);
and U21503 (N_21503,N_16009,N_19024);
nor U21504 (N_21504,N_17286,N_15402);
and U21505 (N_21505,N_16330,N_19137);
and U21506 (N_21506,N_18202,N_18003);
xor U21507 (N_21507,N_16491,N_16297);
nand U21508 (N_21508,N_19610,N_16608);
and U21509 (N_21509,N_18887,N_16768);
or U21510 (N_21510,N_15258,N_17882);
or U21511 (N_21511,N_15028,N_19026);
nor U21512 (N_21512,N_19109,N_18628);
nor U21513 (N_21513,N_18078,N_16571);
nor U21514 (N_21514,N_17644,N_15541);
and U21515 (N_21515,N_19178,N_17481);
nand U21516 (N_21516,N_15320,N_19862);
and U21517 (N_21517,N_18002,N_15408);
nand U21518 (N_21518,N_18379,N_19366);
nand U21519 (N_21519,N_16062,N_19242);
nand U21520 (N_21520,N_15426,N_16730);
or U21521 (N_21521,N_15330,N_15249);
nor U21522 (N_21522,N_16141,N_17336);
nand U21523 (N_21523,N_17148,N_17292);
nand U21524 (N_21524,N_17851,N_16907);
nor U21525 (N_21525,N_18068,N_19536);
nor U21526 (N_21526,N_16636,N_17876);
nor U21527 (N_21527,N_17750,N_18474);
nor U21528 (N_21528,N_19300,N_18057);
nand U21529 (N_21529,N_16656,N_19853);
and U21530 (N_21530,N_19583,N_18665);
and U21531 (N_21531,N_17104,N_17962);
or U21532 (N_21532,N_17573,N_17432);
or U21533 (N_21533,N_16612,N_17563);
and U21534 (N_21534,N_17500,N_16542);
and U21535 (N_21535,N_15299,N_15270);
and U21536 (N_21536,N_15340,N_15587);
nand U21537 (N_21537,N_15861,N_17970);
nand U21538 (N_21538,N_15139,N_18526);
nor U21539 (N_21539,N_17004,N_15462);
nand U21540 (N_21540,N_15253,N_18040);
and U21541 (N_21541,N_17319,N_19885);
nor U21542 (N_21542,N_16164,N_15398);
nand U21543 (N_21543,N_15465,N_16769);
and U21544 (N_21544,N_19929,N_15973);
nor U21545 (N_21545,N_15889,N_16079);
and U21546 (N_21546,N_17310,N_19492);
or U21547 (N_21547,N_15274,N_18458);
nand U21548 (N_21548,N_16211,N_15593);
or U21549 (N_21549,N_15151,N_19325);
or U21550 (N_21550,N_15397,N_15514);
and U21551 (N_21551,N_16569,N_17756);
or U21552 (N_21552,N_19662,N_17712);
and U21553 (N_21553,N_17078,N_17414);
or U21554 (N_21554,N_15601,N_17960);
or U21555 (N_21555,N_18304,N_15585);
or U21556 (N_21556,N_17359,N_18037);
and U21557 (N_21557,N_16998,N_17601);
nand U21558 (N_21558,N_17628,N_15079);
xnor U21559 (N_21559,N_16710,N_19310);
or U21560 (N_21560,N_17844,N_19759);
and U21561 (N_21561,N_15404,N_16727);
xor U21562 (N_21562,N_16808,N_15600);
nand U21563 (N_21563,N_16235,N_15272);
xnor U21564 (N_21564,N_19062,N_17757);
and U21565 (N_21565,N_16920,N_15066);
or U21566 (N_21566,N_18579,N_18886);
nand U21567 (N_21567,N_16404,N_19799);
xnor U21568 (N_21568,N_16239,N_18779);
or U21569 (N_21569,N_18934,N_19437);
or U21570 (N_21570,N_17460,N_17284);
nor U21571 (N_21571,N_15868,N_16771);
and U21572 (N_21572,N_18877,N_18519);
nand U21573 (N_21573,N_15252,N_18007);
and U21574 (N_21574,N_17084,N_19867);
nand U21575 (N_21575,N_16149,N_17855);
nand U21576 (N_21576,N_15992,N_19158);
and U21577 (N_21577,N_17200,N_18691);
or U21578 (N_21578,N_15369,N_15276);
or U21579 (N_21579,N_17660,N_19648);
nor U21580 (N_21580,N_17631,N_17870);
nand U21581 (N_21581,N_18165,N_17547);
or U21582 (N_21582,N_15464,N_15630);
nor U21583 (N_21583,N_16026,N_17992);
or U21584 (N_21584,N_18554,N_16622);
or U21585 (N_21585,N_19048,N_19245);
nand U21586 (N_21586,N_16882,N_19937);
nand U21587 (N_21587,N_16475,N_15267);
or U21588 (N_21588,N_17826,N_17453);
nand U21589 (N_21589,N_15851,N_16510);
nor U21590 (N_21590,N_19082,N_17534);
nand U21591 (N_21591,N_15101,N_18766);
nor U21592 (N_21592,N_16670,N_15849);
nand U21593 (N_21593,N_16624,N_16961);
nand U21594 (N_21594,N_15998,N_16286);
nor U21595 (N_21595,N_19989,N_19423);
nor U21596 (N_21596,N_17122,N_16382);
nor U21597 (N_21597,N_15790,N_16843);
nor U21598 (N_21598,N_17095,N_19991);
and U21599 (N_21599,N_17565,N_16987);
and U21600 (N_21600,N_17860,N_15502);
or U21601 (N_21601,N_18929,N_18894);
and U21602 (N_21602,N_18238,N_18963);
nand U21603 (N_21603,N_19876,N_16623);
nand U21604 (N_21604,N_15263,N_18344);
nor U21605 (N_21605,N_17012,N_16804);
nand U21606 (N_21606,N_17637,N_15625);
and U21607 (N_21607,N_15943,N_19625);
and U21608 (N_21608,N_15871,N_18262);
and U21609 (N_21609,N_19081,N_18174);
or U21610 (N_21610,N_19097,N_15122);
or U21611 (N_21611,N_18089,N_19600);
or U21612 (N_21612,N_17647,N_17074);
or U21613 (N_21613,N_17846,N_19522);
nand U21614 (N_21614,N_15961,N_17232);
or U21615 (N_21615,N_15570,N_18777);
or U21616 (N_21616,N_17667,N_15449);
nor U21617 (N_21617,N_16600,N_17552);
nor U21618 (N_21618,N_19397,N_15319);
and U21619 (N_21619,N_15469,N_15086);
nor U21620 (N_21620,N_18293,N_18060);
and U21621 (N_21621,N_15717,N_18563);
nor U21622 (N_21622,N_15937,N_19425);
nor U21623 (N_21623,N_16053,N_19701);
or U21624 (N_21624,N_15877,N_15443);
nor U21625 (N_21625,N_16745,N_18988);
nor U21626 (N_21626,N_16766,N_16162);
nand U21627 (N_21627,N_19762,N_18199);
nand U21628 (N_21628,N_15158,N_17191);
or U21629 (N_21629,N_15374,N_15598);
and U21630 (N_21630,N_17338,N_18944);
or U21631 (N_21631,N_19871,N_15797);
or U21632 (N_21632,N_19312,N_19611);
nor U21633 (N_21633,N_16993,N_18783);
or U21634 (N_21634,N_17832,N_16762);
nor U21635 (N_21635,N_18193,N_16728);
and U21636 (N_21636,N_19255,N_17686);
and U21637 (N_21637,N_15172,N_16740);
or U21638 (N_21638,N_15072,N_15156);
and U21639 (N_21639,N_17488,N_17820);
and U21640 (N_21640,N_15839,N_17390);
nand U21641 (N_21641,N_19461,N_18677);
and U21642 (N_21642,N_16125,N_19670);
or U21643 (N_21643,N_15112,N_15549);
and U21644 (N_21644,N_16484,N_16081);
nor U21645 (N_21645,N_19058,N_19156);
nor U21646 (N_21646,N_16106,N_15523);
or U21647 (N_21647,N_18276,N_18531);
nor U21648 (N_21648,N_18694,N_15209);
nand U21649 (N_21649,N_19859,N_15558);
or U21650 (N_21650,N_19532,N_17187);
nor U21651 (N_21651,N_15897,N_17597);
or U21652 (N_21652,N_15474,N_17431);
nand U21653 (N_21653,N_15692,N_16585);
and U21654 (N_21654,N_17369,N_17596);
xor U21655 (N_21655,N_17217,N_17394);
nand U21656 (N_21656,N_15006,N_19591);
or U21657 (N_21657,N_16988,N_19225);
nand U21658 (N_21658,N_18318,N_16602);
nand U21659 (N_21659,N_17404,N_18255);
nand U21660 (N_21660,N_18360,N_19913);
or U21661 (N_21661,N_16381,N_15124);
and U21662 (N_21662,N_18696,N_16713);
nand U21663 (N_21663,N_17829,N_17107);
nand U21664 (N_21664,N_16856,N_17124);
nand U21665 (N_21665,N_15056,N_17177);
nand U21666 (N_21666,N_19786,N_19486);
nor U21667 (N_21667,N_19044,N_19692);
or U21668 (N_21668,N_19343,N_19824);
and U21669 (N_21669,N_19938,N_16807);
nand U21670 (N_21670,N_15966,N_15348);
nand U21671 (N_21671,N_16429,N_17763);
nand U21672 (N_21672,N_19233,N_17621);
nor U21673 (N_21673,N_19160,N_17746);
or U21674 (N_21674,N_16280,N_16391);
nand U21675 (N_21675,N_15644,N_19334);
xnor U21676 (N_21676,N_19398,N_18889);
nor U21677 (N_21677,N_17153,N_15132);
or U21678 (N_21678,N_19324,N_15801);
or U21679 (N_21679,N_19602,N_15001);
nand U21680 (N_21680,N_15945,N_16157);
nand U21681 (N_21681,N_16217,N_15623);
nor U21682 (N_21682,N_17868,N_17446);
and U21683 (N_21683,N_17140,N_17505);
and U21684 (N_21684,N_18195,N_18846);
or U21685 (N_21685,N_16940,N_19699);
nand U21686 (N_21686,N_18869,N_17473);
nand U21687 (N_21687,N_19052,N_19590);
or U21688 (N_21688,N_19053,N_15638);
nor U21689 (N_21689,N_19408,N_17797);
and U21690 (N_21690,N_17304,N_19588);
nor U21691 (N_21691,N_17098,N_19819);
nand U21692 (N_21692,N_17612,N_19386);
and U21693 (N_21693,N_17623,N_15622);
nand U21694 (N_21694,N_19580,N_18025);
or U21695 (N_21695,N_15696,N_18353);
and U21696 (N_21696,N_18621,N_19415);
and U21697 (N_21697,N_16420,N_18053);
xor U21698 (N_21698,N_19228,N_15150);
nand U21699 (N_21699,N_15207,N_19241);
or U21700 (N_21700,N_15205,N_17884);
or U21701 (N_21701,N_16195,N_16662);
or U21702 (N_21702,N_15612,N_16229);
and U21703 (N_21703,N_17564,N_16295);
or U21704 (N_21704,N_18210,N_15911);
nand U21705 (N_21705,N_18275,N_17216);
and U21706 (N_21706,N_17774,N_16278);
or U21707 (N_21707,N_16663,N_16640);
and U21708 (N_21708,N_17294,N_19980);
and U21709 (N_21709,N_17988,N_17110);
xor U21710 (N_21710,N_15672,N_15296);
and U21711 (N_21711,N_15699,N_15567);
nor U21712 (N_21712,N_15893,N_19748);
nor U21713 (N_21713,N_17374,N_15650);
or U21714 (N_21714,N_18831,N_16573);
nand U21715 (N_21715,N_15160,N_15633);
or U21716 (N_21716,N_19387,N_19405);
nor U21717 (N_21717,N_15802,N_18538);
or U21718 (N_21718,N_16422,N_17732);
and U21719 (N_21719,N_17142,N_17889);
or U21720 (N_21720,N_18911,N_17170);
and U21721 (N_21721,N_15542,N_19964);
nor U21722 (N_21722,N_17865,N_16189);
or U21723 (N_21723,N_18398,N_19646);
or U21724 (N_21724,N_17956,N_15065);
nand U21725 (N_21725,N_16721,N_15608);
nor U21726 (N_21726,N_16942,N_18987);
nor U21727 (N_21727,N_17706,N_19626);
and U21728 (N_21728,N_19195,N_18626);
nor U21729 (N_21729,N_17510,N_16545);
and U21730 (N_21730,N_17845,N_16359);
nor U21731 (N_21731,N_18157,N_19899);
and U21732 (N_21732,N_15313,N_18299);
or U21733 (N_21733,N_18059,N_15831);
nor U21734 (N_21734,N_15905,N_19746);
and U21735 (N_21735,N_15429,N_16944);
and U21736 (N_21736,N_18186,N_15386);
nor U21737 (N_21737,N_18335,N_18137);
nand U21738 (N_21738,N_18121,N_16348);
nand U21739 (N_21739,N_18132,N_18085);
and U21740 (N_21740,N_17030,N_15349);
and U21741 (N_21741,N_17123,N_16896);
or U21742 (N_21742,N_15634,N_18086);
and U21743 (N_21743,N_18228,N_19067);
and U21744 (N_21744,N_16943,N_18091);
and U21745 (N_21745,N_16375,N_19478);
or U21746 (N_21746,N_17577,N_16332);
or U21747 (N_21747,N_17241,N_19864);
nand U21748 (N_21748,N_15032,N_16819);
xor U21749 (N_21749,N_15167,N_19694);
or U21750 (N_21750,N_15459,N_16933);
nand U21751 (N_21751,N_16021,N_19014);
and U21752 (N_21752,N_19693,N_19426);
nand U21753 (N_21753,N_17936,N_18045);
nand U21754 (N_21754,N_19140,N_19006);
nand U21755 (N_21755,N_16215,N_16267);
or U21756 (N_21756,N_15656,N_16523);
nand U21757 (N_21757,N_17523,N_16667);
nor U21758 (N_21758,N_17971,N_18589);
nor U21759 (N_21759,N_17963,N_19338);
or U21760 (N_21760,N_19797,N_16442);
or U21761 (N_21761,N_16567,N_16317);
nand U21762 (N_21762,N_19846,N_16777);
nor U21763 (N_21763,N_17818,N_15080);
nand U21764 (N_21764,N_19922,N_15709);
and U21765 (N_21765,N_17455,N_16628);
or U21766 (N_21766,N_16589,N_18995);
nand U21767 (N_21767,N_17796,N_17056);
xor U21768 (N_21768,N_18090,N_15392);
nand U21769 (N_21769,N_17065,N_19148);
or U21770 (N_21770,N_18478,N_18152);
nor U21771 (N_21771,N_17966,N_15147);
nor U21772 (N_21772,N_19355,N_17265);
nor U21773 (N_21773,N_16550,N_19570);
or U21774 (N_21774,N_17553,N_15909);
nor U21775 (N_21775,N_17197,N_17710);
nand U21776 (N_21776,N_19257,N_16483);
and U21777 (N_21777,N_19289,N_17927);
or U21778 (N_21778,N_16351,N_16094);
or U21779 (N_21779,N_16452,N_18283);
nand U21780 (N_21780,N_19002,N_19794);
nor U21781 (N_21781,N_16405,N_16552);
xnor U21782 (N_21782,N_16691,N_19944);
and U21783 (N_21783,N_17180,N_15703);
or U21784 (N_21784,N_18888,N_17228);
xnor U21785 (N_21785,N_16132,N_15997);
and U21786 (N_21786,N_15977,N_15566);
nor U21787 (N_21787,N_15792,N_19154);
and U21788 (N_21788,N_17572,N_16179);
nor U21789 (N_21789,N_17898,N_15746);
nor U21790 (N_21790,N_15461,N_15736);
or U21791 (N_21791,N_15244,N_16073);
or U21792 (N_21792,N_19807,N_15779);
nand U21793 (N_21793,N_19180,N_19934);
nor U21794 (N_21794,N_16136,N_15863);
or U21795 (N_21795,N_18829,N_15584);
nand U21796 (N_21796,N_18899,N_17673);
nor U21797 (N_21797,N_19179,N_18603);
nor U21798 (N_21798,N_15460,N_19987);
and U21799 (N_21799,N_16005,N_19186);
and U21800 (N_21800,N_18326,N_16751);
xnor U21801 (N_21801,N_17380,N_19230);
nor U21802 (N_21802,N_16767,N_15547);
and U21803 (N_21803,N_16464,N_16654);
and U21804 (N_21804,N_15280,N_18414);
and U21805 (N_21805,N_16784,N_15843);
nor U21806 (N_21806,N_18735,N_19468);
or U21807 (N_21807,N_16692,N_16116);
nand U21808 (N_21808,N_19376,N_17334);
nor U21809 (N_21809,N_18845,N_17151);
nor U21810 (N_21810,N_15667,N_19541);
and U21811 (N_21811,N_16155,N_15328);
nor U21812 (N_21812,N_19015,N_19901);
nand U21813 (N_21813,N_18683,N_18290);
nand U21814 (N_21814,N_15165,N_17271);
nor U21815 (N_21815,N_16275,N_16719);
nor U21816 (N_21816,N_18463,N_15533);
nand U21817 (N_21817,N_18891,N_19169);
nand U21818 (N_21818,N_15202,N_19844);
nor U21819 (N_21819,N_16276,N_17658);
and U21820 (N_21820,N_16479,N_19369);
and U21821 (N_21821,N_19102,N_18386);
and U21822 (N_21822,N_16957,N_19551);
nor U21823 (N_21823,N_19803,N_19202);
and U21824 (N_21824,N_19533,N_16899);
or U21825 (N_21825,N_15794,N_18102);
nor U21826 (N_21826,N_15653,N_19881);
and U21827 (N_21827,N_17444,N_19716);
or U21828 (N_21828,N_18364,N_17618);
nor U21829 (N_21829,N_16292,N_19861);
or U21830 (N_21830,N_17616,N_15312);
nor U21831 (N_21831,N_18864,N_19563);
or U21832 (N_21832,N_18746,N_16774);
nor U21833 (N_21833,N_18804,N_16260);
nor U21834 (N_21834,N_19046,N_19898);
xor U21835 (N_21835,N_16714,N_19189);
or U21836 (N_21836,N_17370,N_17788);
or U21837 (N_21837,N_16298,N_17054);
nor U21838 (N_21838,N_19904,N_18216);
nor U21839 (N_21839,N_17366,N_18983);
nor U21840 (N_21840,N_15841,N_19219);
or U21841 (N_21841,N_16016,N_17901);
or U21842 (N_21842,N_17137,N_18591);
and U21843 (N_21843,N_19540,N_19056);
nand U21844 (N_21844,N_16779,N_15242);
or U21845 (N_21845,N_17799,N_18470);
or U21846 (N_21846,N_16245,N_18190);
nor U21847 (N_21847,N_16633,N_19912);
nor U21848 (N_21848,N_19758,N_15478);
or U21849 (N_21849,N_16334,N_17363);
and U21850 (N_21850,N_17221,N_17806);
nand U21851 (N_21851,N_16903,N_15524);
and U21852 (N_21852,N_18943,N_18770);
nand U21853 (N_21853,N_16574,N_16312);
and U21854 (N_21854,N_18416,N_17680);
nand U21855 (N_21855,N_19946,N_19565);
nor U21856 (N_21856,N_16708,N_15351);
or U21857 (N_21857,N_19487,N_19192);
nor U21858 (N_21858,N_15100,N_15606);
or U21859 (N_21859,N_18863,N_16105);
nand U21860 (N_21860,N_19756,N_17883);
nor U21861 (N_21861,N_17854,N_15463);
nor U21862 (N_21862,N_17881,N_18505);
nand U21863 (N_21863,N_18382,N_16815);
nand U21864 (N_21864,N_16341,N_18191);
xnor U21865 (N_21865,N_17062,N_15812);
nor U21866 (N_21866,N_17245,N_15604);
and U21867 (N_21867,N_19695,N_17784);
nor U21868 (N_21868,N_16448,N_19564);
nor U21869 (N_21869,N_16884,N_15200);
and U21870 (N_21870,N_15405,N_18156);
nand U21871 (N_21871,N_19360,N_15020);
nand U21872 (N_21872,N_19816,N_19737);
and U21873 (N_21873,N_19784,N_19718);
nor U21874 (N_21874,N_16535,N_17022);
or U21875 (N_21875,N_19633,N_17748);
nand U21876 (N_21876,N_15199,N_15025);
nor U21877 (N_21877,N_16620,N_18634);
and U21878 (N_21878,N_16367,N_15189);
nor U21879 (N_21879,N_19128,N_16799);
nand U21880 (N_21880,N_17681,N_17349);
and U21881 (N_21881,N_16871,N_19298);
nor U21882 (N_21882,N_17707,N_16146);
or U21883 (N_21883,N_18557,N_15627);
or U21884 (N_21884,N_19587,N_18562);
and U21885 (N_21885,N_18473,N_15048);
and U21886 (N_21886,N_15171,N_15247);
nand U21887 (N_21887,N_16560,N_17428);
and U21888 (N_21888,N_17741,N_17747);
and U21889 (N_21889,N_18711,N_18520);
nor U21890 (N_21890,N_15117,N_16698);
nand U21891 (N_21891,N_19285,N_18720);
and U21892 (N_21892,N_15527,N_19220);
nor U21893 (N_21893,N_15365,N_19849);
nor U21894 (N_21894,N_18153,N_16647);
or U21895 (N_21895,N_19045,N_15421);
nor U21896 (N_21896,N_16025,N_15277);
nor U21897 (N_21897,N_18251,N_18572);
nand U21898 (N_21898,N_16631,N_19674);
nand U21899 (N_21899,N_18828,N_17554);
nand U21900 (N_21900,N_17926,N_18361);
xor U21901 (N_21901,N_19663,N_17324);
nand U21902 (N_21902,N_15930,N_16372);
and U21903 (N_21903,N_17383,N_18738);
and U21904 (N_21904,N_17742,N_16480);
nor U21905 (N_21905,N_17253,N_15701);
or U21906 (N_21906,N_19768,N_15684);
or U21907 (N_21907,N_15472,N_19594);
and U21908 (N_21908,N_15804,N_18784);
or U21909 (N_21909,N_15538,N_18425);
nor U21910 (N_21910,N_18029,N_18756);
and U21911 (N_21911,N_18647,N_19170);
nand U21912 (N_21912,N_16299,N_15018);
nor U21913 (N_21913,N_17895,N_18260);
or U21914 (N_21914,N_18427,N_15865);
nand U21915 (N_21915,N_19143,N_19249);
and U21916 (N_21916,N_15491,N_19568);
or U21917 (N_21917,N_15512,N_17350);
or U21918 (N_21918,N_15058,N_15980);
nor U21919 (N_21919,N_16058,N_16526);
or U21920 (N_21920,N_15733,N_19644);
and U21921 (N_21921,N_16992,N_18560);
and U21922 (N_21922,N_18311,N_16761);
and U21923 (N_21923,N_17348,N_17979);
nor U21924 (N_21924,N_16440,N_18999);
nand U21925 (N_21925,N_15218,N_17037);
and U21926 (N_21926,N_16170,N_19841);
or U21927 (N_21927,N_18990,N_19276);
nand U21928 (N_21928,N_18979,N_17526);
or U21929 (N_21929,N_17406,N_17812);
nand U21930 (N_21930,N_19072,N_16183);
or U21931 (N_21931,N_19008,N_17964);
nor U21932 (N_21932,N_19994,N_15595);
and U21933 (N_21933,N_18383,N_16460);
and U21934 (N_21934,N_16041,N_17798);
nand U21935 (N_21935,N_15295,N_15438);
xnor U21936 (N_21936,N_15647,N_18982);
nor U21937 (N_21937,N_18323,N_18945);
nand U21938 (N_21938,N_15081,N_17163);
nand U21939 (N_21939,N_16261,N_19175);
and U21940 (N_21940,N_16598,N_18178);
nand U21941 (N_21941,N_17167,N_17264);
and U21942 (N_21942,N_16387,N_19363);
nand U21943 (N_21943,N_18221,N_15260);
and U21944 (N_21944,N_16050,N_16078);
nand U21945 (N_21945,N_19534,N_15279);
nand U21946 (N_21946,N_15501,N_15376);
or U21947 (N_21947,N_17905,N_16431);
or U21948 (N_21948,N_18898,N_19645);
nand U21949 (N_21949,N_19021,N_16385);
nand U21950 (N_21950,N_16517,N_15724);
and U21951 (N_21951,N_16145,N_15520);
nand U21952 (N_21952,N_17354,N_18436);
and U21953 (N_21953,N_19061,N_18815);
or U21954 (N_21954,N_17202,N_16997);
or U21955 (N_21955,N_18640,N_19243);
nor U21956 (N_21956,N_16847,N_17529);
nand U21957 (N_21957,N_16443,N_18928);
nor U21958 (N_21958,N_17326,N_17135);
or U21959 (N_21959,N_18457,N_15711);
and U21960 (N_21960,N_17164,N_17536);
nor U21961 (N_21961,N_19106,N_15239);
nand U21962 (N_21962,N_16194,N_16533);
nand U21963 (N_21963,N_17546,N_17622);
and U21964 (N_21964,N_18055,N_18974);
nor U21965 (N_21965,N_18796,N_17886);
nor U21966 (N_21966,N_16077,N_17314);
and U21967 (N_21967,N_18546,N_15940);
nand U21968 (N_21968,N_16181,N_15275);
or U21969 (N_21969,N_15191,N_16388);
nor U21970 (N_21970,N_17060,N_18048);
and U21971 (N_21971,N_19793,N_17464);
nor U21972 (N_21972,N_16205,N_18369);
and U21973 (N_21973,N_16839,N_15050);
or U21974 (N_21974,N_18719,N_15403);
or U21975 (N_21975,N_19421,N_19683);
and U21976 (N_21976,N_18319,N_19830);
and U21977 (N_21977,N_19060,N_16046);
nor U21978 (N_21978,N_15204,N_17309);
or U21979 (N_21979,N_15487,N_19215);
nor U21980 (N_21980,N_19098,N_16010);
nand U21981 (N_21981,N_15654,N_16088);
or U21982 (N_21982,N_19496,N_16188);
nand U21983 (N_21983,N_18087,N_17342);
nor U21984 (N_21984,N_19836,N_19011);
or U21985 (N_21985,N_15214,N_18693);
and U21986 (N_21986,N_17272,N_17924);
nor U21987 (N_21987,N_19665,N_18248);
nand U21988 (N_21988,N_19815,N_16424);
nand U21989 (N_21989,N_19887,N_16057);
and U21990 (N_21990,N_17599,N_19273);
and U21991 (N_21991,N_16911,N_19855);
or U21992 (N_21992,N_19217,N_16772);
nand U21993 (N_21993,N_18013,N_16006);
or U21994 (N_21994,N_18878,N_18331);
nor U21995 (N_21995,N_15545,N_16313);
and U21996 (N_21996,N_16246,N_17301);
or U21997 (N_21997,N_17866,N_15591);
and U21998 (N_21998,N_19223,N_19918);
nor U21999 (N_21999,N_16965,N_18960);
nand U22000 (N_22000,N_17627,N_17824);
nor U22001 (N_22001,N_16947,N_15872);
or U22002 (N_22002,N_17821,N_17296);
nand U22003 (N_22003,N_16820,N_19352);
or U22004 (N_22004,N_15759,N_17679);
nor U22005 (N_22005,N_18343,N_16860);
and U22006 (N_22006,N_18801,N_15043);
nor U22007 (N_22007,N_15986,N_18852);
and U22008 (N_22008,N_18850,N_17809);
nand U22009 (N_22009,N_18138,N_19412);
nor U22010 (N_22010,N_18710,N_16964);
and U22011 (N_22011,N_15776,N_17683);
nand U22012 (N_22012,N_18144,N_17814);
nor U22013 (N_22013,N_17417,N_16945);
nor U22014 (N_22014,N_19187,N_17308);
and U22015 (N_22015,N_16844,N_19116);
and U22016 (N_22016,N_17372,N_17287);
xnor U22017 (N_22017,N_16897,N_17026);
or U22018 (N_22018,N_17520,N_17492);
nor U22019 (N_22019,N_18512,N_15881);
xor U22020 (N_22020,N_19965,N_16318);
nor U22021 (N_22021,N_19268,N_17412);
nand U22022 (N_22022,N_17008,N_17236);
or U22023 (N_22023,N_16717,N_15620);
nor U22024 (N_22024,N_15197,N_17888);
and U22025 (N_22025,N_19687,N_18396);
or U22026 (N_22026,N_17459,N_19679);
nand U22027 (N_22027,N_15120,N_17423);
xor U22028 (N_22028,N_16433,N_16702);
or U22029 (N_22029,N_19069,N_17368);
nor U22030 (N_22030,N_18287,N_16310);
and U22031 (N_22031,N_15860,N_18307);
and U22032 (N_22032,N_17965,N_18282);
and U22033 (N_22033,N_19700,N_15596);
or U22034 (N_22034,N_19467,N_19177);
nor U22035 (N_22035,N_17109,N_15615);
nor U22036 (N_22036,N_18140,N_18792);
nor U22037 (N_22037,N_16732,N_18295);
xnor U22038 (N_22038,N_16186,N_16737);
nand U22039 (N_22039,N_17185,N_16212);
nand U22040 (N_22040,N_16115,N_17405);
xnor U22041 (N_22041,N_19445,N_17274);
nand U22042 (N_22042,N_15729,N_17018);
and U22043 (N_22043,N_18664,N_17156);
or U22044 (N_22044,N_18872,N_16515);
nand U22045 (N_22045,N_16097,N_19542);
nor U22046 (N_22046,N_17283,N_15012);
nand U22047 (N_22047,N_17728,N_18965);
nor U22048 (N_22048,N_18811,N_17067);
xnor U22049 (N_22049,N_17945,N_19341);
nand U22050 (N_22050,N_18236,N_15690);
nor U22051 (N_22051,N_17086,N_19848);
or U22052 (N_22052,N_15939,N_15342);
nor U22053 (N_22053,N_17485,N_19297);
or U22054 (N_22054,N_16511,N_19013);
nand U22055 (N_22055,N_19383,N_16848);
or U22056 (N_22056,N_19983,N_16507);
xor U22057 (N_22057,N_16417,N_18460);
nand U22058 (N_22058,N_19909,N_17385);
nand U22059 (N_22059,N_19690,N_15671);
nand U22060 (N_22060,N_16908,N_18374);
nand U22061 (N_22061,N_15223,N_18012);
nor U22062 (N_22062,N_15780,N_18732);
or U22063 (N_22063,N_15286,N_15537);
and U22064 (N_22064,N_19685,N_19531);
nand U22065 (N_22065,N_15143,N_18214);
and U22066 (N_22066,N_19698,N_15693);
nand U22067 (N_22067,N_16084,N_16344);
or U22068 (N_22068,N_18722,N_16968);
and U22069 (N_22069,N_19159,N_19438);
xor U22070 (N_22070,N_19947,N_15341);
nand U22071 (N_22071,N_18009,N_18352);
nor U22072 (N_22072,N_16973,N_16070);
nor U22073 (N_22073,N_16107,N_15858);
nor U22074 (N_22074,N_16838,N_19660);
nor U22075 (N_22075,N_17991,N_15528);
and U22076 (N_22076,N_16668,N_18081);
or U22077 (N_22077,N_17912,N_18788);
nand U22078 (N_22078,N_15084,N_15569);
and U22079 (N_22079,N_16203,N_18330);
or U22080 (N_22080,N_19907,N_17739);
or U22081 (N_22081,N_15507,N_18034);
nand U22082 (N_22082,N_15356,N_17183);
or U22083 (N_22083,N_17048,N_17902);
or U22084 (N_22084,N_16921,N_16165);
or U22085 (N_22085,N_15166,N_15444);
nand U22086 (N_22086,N_15626,N_19710);
and U22087 (N_22087,N_15224,N_19027);
nand U22088 (N_22088,N_15573,N_17561);
nand U22089 (N_22089,N_17489,N_15783);
or U22090 (N_22090,N_17059,N_19095);
nand U22091 (N_22091,N_18163,N_19820);
nand U22092 (N_22092,N_15683,N_18433);
nand U22093 (N_22093,N_18325,N_19655);
or U22094 (N_22094,N_16791,N_16371);
nand U22095 (N_22095,N_19279,N_19240);
nor U22096 (N_22096,N_17154,N_17743);
or U22097 (N_22097,N_16415,N_16881);
nor U22098 (N_22098,N_18989,N_19488);
nor U22099 (N_22099,N_19004,N_16635);
nand U22100 (N_22100,N_15248,N_18823);
or U22101 (N_22101,N_16363,N_15024);
nor U22102 (N_22102,N_15321,N_19897);
nor U22103 (N_22103,N_17585,N_18909);
xnor U22104 (N_22104,N_18213,N_17192);
or U22105 (N_22105,N_19302,N_15380);
and U22106 (N_22106,N_16131,N_15490);
or U22107 (N_22107,N_15822,N_15536);
nor U22108 (N_22108,N_16252,N_15720);
nor U22109 (N_22109,N_16867,N_18695);
and U22110 (N_22110,N_15379,N_19567);
nor U22111 (N_22111,N_15755,N_15194);
nor U22112 (N_22112,N_16139,N_15529);
or U22113 (N_22113,N_16606,N_15092);
and U22114 (N_22114,N_17567,N_18134);
nor U22115 (N_22115,N_19792,N_15979);
nand U22116 (N_22116,N_18410,N_19597);
and U22117 (N_22117,N_18363,N_15229);
nor U22118 (N_22118,N_15070,N_19183);
and U22119 (N_22119,N_16711,N_19555);
or U22120 (N_22120,N_16678,N_16243);
or U22121 (N_22121,N_17051,N_18058);
nand U22122 (N_22122,N_15721,N_18198);
or U22123 (N_22123,N_18912,N_18375);
nor U22124 (N_22124,N_19326,N_15793);
nor U22125 (N_22125,N_18739,N_17229);
nand U22126 (N_22126,N_18631,N_17461);
nor U22127 (N_22127,N_16001,N_19878);
and U22128 (N_22128,N_15173,N_18964);
or U22129 (N_22129,N_16130,N_15393);
and U22130 (N_22130,N_17024,N_16994);
nor U22131 (N_22131,N_18175,N_17476);
nand U22132 (N_22132,N_15359,N_19005);
or U22133 (N_22133,N_19237,N_16419);
nand U22134 (N_22134,N_15396,N_16704);
and U22135 (N_22135,N_17947,N_17243);
nand U22136 (N_22136,N_18146,N_17306);
nor U22137 (N_22137,N_15273,N_18511);
and U22138 (N_22138,N_16462,N_19515);
and U22139 (N_22139,N_19998,N_17225);
nand U22140 (N_22140,N_17580,N_16519);
and U22141 (N_22141,N_17984,N_15175);
and U22142 (N_22142,N_18598,N_16362);
nor U22143 (N_22143,N_17643,N_17811);
and U22144 (N_22144,N_15959,N_16042);
and U22145 (N_22145,N_19280,N_19982);
nor U22146 (N_22146,N_19007,N_15476);
and U22147 (N_22147,N_18404,N_15927);
or U22148 (N_22148,N_17491,N_18372);
or U22149 (N_22149,N_17071,N_19529);
or U22150 (N_22150,N_19835,N_18920);
and U22151 (N_22151,N_17422,N_19208);
nor U22152 (N_22152,N_15059,N_17906);
xnor U22153 (N_22153,N_19508,N_16017);
nor U22154 (N_22154,N_19630,N_17361);
and U22155 (N_22155,N_17560,N_18497);
and U22156 (N_22156,N_19585,N_15201);
and U22157 (N_22157,N_19910,N_17699);
xnor U22158 (N_22158,N_19145,N_15423);
or U22159 (N_22159,N_17808,N_17209);
nand U22160 (N_22160,N_17791,N_18540);
and U22161 (N_22161,N_17542,N_19514);
nand U22162 (N_22162,N_18316,N_17015);
nor U22163 (N_22163,N_19100,N_17429);
nand U22164 (N_22164,N_19401,N_19460);
and U22165 (N_22165,N_15924,N_15574);
or U22166 (N_22166,N_18020,N_18500);
nand U22167 (N_22167,N_17407,N_17516);
and U22168 (N_22168,N_17079,N_18748);
nand U22169 (N_22169,N_19294,N_18166);
or U22170 (N_22170,N_15036,N_16250);
nor U22171 (N_22171,N_17313,N_19346);
nor U22172 (N_22172,N_18569,N_16521);
and U22173 (N_22173,N_16412,N_19466);
and U22174 (N_22174,N_18245,N_16850);
nor U22175 (N_22175,N_18657,N_16468);
and U22176 (N_22176,N_16036,N_17915);
xnor U22177 (N_22177,N_16974,N_15956);
and U22178 (N_22178,N_18019,N_15231);
nor U22179 (N_22179,N_15088,N_16960);
or U22180 (N_22180,N_17501,N_15322);
nor U22181 (N_22181,N_17362,N_17754);
nand U22182 (N_22182,N_18108,N_19303);
nor U22183 (N_22183,N_18761,N_19649);
nand U22184 (N_22184,N_19914,N_16221);
nand U22185 (N_22185,N_17335,N_15543);
or U22186 (N_22186,N_17131,N_18357);
or U22187 (N_22187,N_16716,N_18821);
xnor U22188 (N_22188,N_18736,N_16782);
and U22189 (N_22189,N_15010,N_19126);
or U22190 (N_22190,N_18073,N_18672);
nand U22191 (N_22191,N_15129,N_15719);
nor U22192 (N_22192,N_15563,N_18212);
or U22193 (N_22193,N_15999,N_17150);
nor U22194 (N_22194,N_19949,N_18545);
nor U22195 (N_22195,N_15325,N_15516);
and U22196 (N_22196,N_16588,N_16950);
nor U22197 (N_22197,N_15686,N_18441);
nand U22198 (N_22198,N_19725,N_18808);
and U22199 (N_22199,N_15588,N_18842);
nand U22200 (N_22200,N_18268,N_19038);
nor U22201 (N_22201,N_18610,N_15749);
and U22202 (N_22202,N_18215,N_19581);
or U22203 (N_22203,N_17266,N_15483);
nor U22204 (N_22204,N_16746,N_18209);
nand U22205 (N_22205,N_19875,N_19194);
or U22206 (N_22206,N_19760,N_15057);
or U22207 (N_22207,N_17050,N_15835);
and U22208 (N_22208,N_18660,N_19200);
nor U22209 (N_22209,N_15039,N_18430);
nand U22210 (N_22210,N_19806,N_18708);
and U22211 (N_22211,N_18896,N_18106);
nand U22212 (N_22212,N_19306,N_16665);
nand U22213 (N_22213,N_15557,N_17116);
or U22214 (N_22214,N_16329,N_18652);
nor U22215 (N_22215,N_15646,N_19446);
or U22216 (N_22216,N_16776,N_18041);
nor U22217 (N_22217,N_16795,N_19077);
nor U22218 (N_22218,N_15854,N_16888);
nand U22219 (N_22219,N_16541,N_18062);
nand U22220 (N_22220,N_19576,N_18464);
and U22221 (N_22221,N_15354,N_16590);
and U22222 (N_22222,N_19372,N_19416);
nand U22223 (N_22223,N_16169,N_18056);
or U22224 (N_22224,N_17355,N_18259);
xor U22225 (N_22225,N_18151,N_17575);
nor U22226 (N_22226,N_17714,N_19811);
or U22227 (N_22227,N_15819,N_17251);
nor U22228 (N_22228,N_15850,N_19367);
nand U22229 (N_22229,N_16984,N_19361);
nand U22230 (N_22230,N_16485,N_18189);
and U22231 (N_22231,N_18642,N_17758);
or U22232 (N_22232,N_17377,N_16108);
or U22233 (N_22233,N_15972,N_16831);
and U22234 (N_22234,N_17003,N_19787);
and U22235 (N_22235,N_17166,N_19181);
or U22236 (N_22236,N_17379,N_16509);
or U22237 (N_22237,N_17863,N_18272);
and U22238 (N_22238,N_16013,N_16801);
or U22239 (N_22239,N_15607,N_19199);
or U22240 (N_22240,N_19121,N_16198);
nand U22241 (N_22241,N_17687,N_17014);
nor U22242 (N_22242,N_16393,N_15344);
nand U22243 (N_22243,N_17659,N_18254);
and U22244 (N_22244,N_17853,N_16835);
and U22245 (N_22245,N_17517,N_19838);
or U22246 (N_22246,N_15548,N_16877);
or U22247 (N_22247,N_18047,N_18755);
nand U22248 (N_22248,N_15067,N_15366);
and U22249 (N_22249,N_17337,N_17917);
and U22250 (N_22250,N_19961,N_16392);
or U22251 (N_22251,N_18700,N_17598);
nand U22252 (N_22252,N_16748,N_19246);
and U22253 (N_22253,N_19105,N_18061);
nor U22254 (N_22254,N_16916,N_17042);
nor U22255 (N_22255,N_15225,N_18565);
nor U22256 (N_22256,N_19414,N_19729);
nand U22257 (N_22257,N_16263,N_17344);
or U22258 (N_22258,N_17169,N_19480);
and U22259 (N_22259,N_17539,N_18867);
nand U22260 (N_22260,N_16869,N_17256);
nand U22261 (N_22261,N_15019,N_15894);
or U22262 (N_22262,N_19927,N_18256);
or U22263 (N_22263,N_19321,N_15974);
and U22264 (N_22264,N_16366,N_16685);
and U22265 (N_22265,N_15681,N_16637);
xor U22266 (N_22266,N_19112,N_18581);
nand U22267 (N_22267,N_19275,N_17764);
xnor U22268 (N_22268,N_16374,N_15368);
and U22269 (N_22269,N_19029,N_18849);
nor U22270 (N_22270,N_19329,N_17165);
or U22271 (N_22271,N_17569,N_19747);
or U22272 (N_22272,N_19612,N_19131);
nand U22273 (N_22273,N_16082,N_16147);
nor U22274 (N_22274,N_19420,N_18625);
or U22275 (N_22275,N_17903,N_16451);
nand U22276 (N_22276,N_17482,N_15187);
nand U22277 (N_22277,N_18754,N_18039);
nand U22278 (N_22278,N_18612,N_17872);
and U22279 (N_22279,N_19042,N_19017);
or U22280 (N_22280,N_16432,N_18329);
nand U22281 (N_22281,N_16741,N_16757);
nand U22282 (N_22282,N_16555,N_19702);
nor U22283 (N_22283,N_15941,N_17448);
and U22284 (N_22284,N_16516,N_18135);
and U22285 (N_22285,N_15246,N_18257);
and U22286 (N_22286,N_15807,N_19812);
nand U22287 (N_22287,N_18402,N_19717);
nor U22288 (N_22288,N_15773,N_17834);
nand U22289 (N_22289,N_19454,N_15097);
nand U22290 (N_22290,N_17240,N_15430);
nor U22291 (N_22291,N_17503,N_16962);
nor U22292 (N_22292,N_16979,N_16750);
or U22293 (N_22293,N_17509,N_19780);
or U22294 (N_22294,N_19671,N_17935);
nor U22295 (N_22295,N_16020,N_17827);
nor U22296 (N_22296,N_19150,N_19136);
or U22297 (N_22297,N_15954,N_16618);
or U22298 (N_22298,N_19556,N_17982);
and U22299 (N_22299,N_16726,N_18303);
nor U22300 (N_22300,N_16531,N_17959);
nor U22301 (N_22301,N_15803,N_19537);
xnor U22302 (N_22302,N_17279,N_15923);
or U22303 (N_22303,N_19538,N_17299);
nor U22304 (N_22304,N_15417,N_15222);
or U22305 (N_22305,N_18380,N_18447);
nand U22306 (N_22306,N_18169,N_15682);
and U22307 (N_22307,N_17729,N_17134);
or U22308 (N_22308,N_16687,N_19719);
nand U22309 (N_22309,N_17638,N_17634);
or U22310 (N_22310,N_15193,N_17393);
and U22311 (N_22311,N_18246,N_18885);
nand U22312 (N_22312,N_18814,N_18022);
and U22313 (N_22313,N_15226,N_17674);
nor U22314 (N_22314,N_19168,N_18438);
nor U22315 (N_22315,N_19845,N_19123);
or U22316 (N_22316,N_19823,N_18351);
nand U22317 (N_22317,N_18667,N_19023);
nor U22318 (N_22318,N_16093,N_18618);
nand U22319 (N_22319,N_16435,N_19092);
or U22320 (N_22320,N_15162,N_19889);
and U22321 (N_22321,N_16080,N_17321);
and U22322 (N_22322,N_18136,N_16883);
and U22323 (N_22323,N_18024,N_17207);
or U22324 (N_22324,N_19667,N_18483);
or U22325 (N_22325,N_16976,N_16140);
nand U22326 (N_22326,N_16579,N_18050);
nor U22327 (N_22327,N_17985,N_15738);
or U22328 (N_22328,N_17400,N_15264);
and U22329 (N_22329,N_19950,N_17418);
nand U22330 (N_22330,N_18648,N_16905);
and U22331 (N_22331,N_17145,N_16007);
nor U22332 (N_22332,N_19353,N_15436);
nor U22333 (N_22333,N_15419,N_19883);
nand U22334 (N_22334,N_16553,N_18822);
nor U22335 (N_22335,N_15304,N_15564);
or U22336 (N_22336,N_17141,N_17867);
nand U22337 (N_22337,N_17734,N_16915);
and U22338 (N_22338,N_18604,N_15196);
nor U22339 (N_22339,N_18923,N_19711);
nand U22340 (N_22340,N_19742,N_19474);
nor U22341 (N_22341,N_16360,N_15639);
or U22342 (N_22342,N_17973,N_19738);
nand U22343 (N_22343,N_16249,N_18843);
xnor U22344 (N_22344,N_19779,N_15920);
or U22345 (N_22345,N_19582,N_15589);
nor U22346 (N_22346,N_16184,N_19888);
and U22347 (N_22347,N_18939,N_18286);
nand U22348 (N_22348,N_17469,N_18533);
or U22349 (N_22349,N_19308,N_15471);
nand U22350 (N_22350,N_15768,N_16219);
and U22351 (N_22351,N_19049,N_15938);
nand U22352 (N_22352,N_18913,N_16087);
or U22353 (N_22353,N_17046,N_15655);
and U22354 (N_22354,N_18517,N_19033);
nor U22355 (N_22355,N_16758,N_19493);
nor U22356 (N_22356,N_16308,N_18206);
or U22357 (N_22357,N_19139,N_19627);
nand U22358 (N_22358,N_17538,N_17514);
and U22359 (N_22359,N_17909,N_19520);
or U22360 (N_22360,N_16174,N_18967);
and U22361 (N_22361,N_16584,N_18763);
and U22362 (N_22362,N_16029,N_15840);
nand U22363 (N_22363,N_19020,N_15265);
nand U22364 (N_22364,N_19254,N_18341);
nand U22365 (N_22365,N_18499,N_16486);
or U22366 (N_22366,N_16206,N_18550);
or U22367 (N_22367,N_16506,N_17478);
or U22368 (N_22368,N_16999,N_18800);
nand U22369 (N_22369,N_19893,N_18832);
nand U22370 (N_22370,N_19444,N_17646);
or U22371 (N_22371,N_19945,N_19818);
and U22372 (N_22372,N_15416,N_17768);
or U22373 (N_22373,N_18807,N_19429);
nand U22374 (N_22374,N_19952,N_17920);
or U22375 (N_22375,N_15830,N_19605);
nand U22376 (N_22376,N_19384,N_19452);
nor U22377 (N_22377,N_16621,N_19767);
or U22378 (N_22378,N_19483,N_18890);
and U22379 (N_22379,N_19447,N_16720);
nor U22380 (N_22380,N_17436,N_15774);
and U22381 (N_22381,N_18501,N_18095);
nand U22382 (N_22382,N_17512,N_19022);
nor U22383 (N_22383,N_15271,N_16975);
nor U22384 (N_22384,N_15388,N_18393);
or U22385 (N_22385,N_16824,N_19345);
and U22386 (N_22386,N_18112,N_18088);
nor U22387 (N_22387,N_17613,N_19442);
nor U22388 (N_22388,N_15400,N_18747);
or U22389 (N_22389,N_16488,N_16421);
nand U22390 (N_22390,N_17922,N_17288);
or U22391 (N_22391,N_15756,N_19988);
nand U22392 (N_22392,N_15758,N_16196);
or U22393 (N_22393,N_19617,N_16314);
xor U22394 (N_22394,N_17518,N_18451);
nand U22395 (N_22395,N_19039,N_17477);
nand U22396 (N_22396,N_15728,N_16099);
nor U22397 (N_22397,N_18205,N_19554);
or U22398 (N_22398,N_19281,N_16120);
and U22399 (N_22399,N_19497,N_18926);
nor U22400 (N_22400,N_18883,N_15519);
or U22401 (N_22401,N_16829,N_16744);
and U22402 (N_22402,N_16706,N_17328);
xor U22403 (N_22403,N_18400,N_17474);
nor U22404 (N_22404,N_16397,N_19858);
nor U22405 (N_22405,N_18405,N_19068);
nand U22406 (N_22406,N_19351,N_19337);
nand U22407 (N_22407,N_19669,N_15083);
nand U22408 (N_22408,N_19900,N_16248);
xnor U22409 (N_22409,N_18336,N_19503);
or U22410 (N_22410,N_16683,N_19389);
xor U22411 (N_22411,N_18663,N_17239);
and U22412 (N_22412,N_19124,N_19034);
and U22413 (N_22413,N_16889,N_17090);
nor U22414 (N_22414,N_18046,N_15037);
and U22415 (N_22415,N_16302,N_15188);
nand U22416 (N_22416,N_19385,N_18597);
nor U22417 (N_22417,N_18838,N_16498);
nand U22418 (N_22418,N_19847,N_17700);
or U22419 (N_22419,N_16027,N_19391);
or U22420 (N_22420,N_18802,N_16953);
xor U22421 (N_22421,N_18699,N_16666);
or U22422 (N_22422,N_19512,N_19301);
or U22423 (N_22423,N_15884,N_16787);
nand U22424 (N_22424,N_19730,N_16160);
nor U22425 (N_22425,N_16038,N_15297);
and U22426 (N_22426,N_15509,N_16918);
or U22427 (N_22427,N_18594,N_15883);
nor U22428 (N_22428,N_15896,N_17064);
nor U22429 (N_22429,N_18158,N_16032);
xor U22430 (N_22430,N_18001,N_19731);
and U22431 (N_22431,N_18948,N_17467);
or U22432 (N_22432,N_18613,N_18903);
nand U22433 (N_22433,N_16864,N_19290);
and U22434 (N_22434,N_16304,N_16827);
nor U22435 (N_22435,N_18424,N_16167);
and U22436 (N_22436,N_18462,N_17112);
nor U22437 (N_22437,N_17533,N_19953);
nand U22438 (N_22438,N_18856,N_15216);
nand U22439 (N_22439,N_15836,N_16472);
nor U22440 (N_22440,N_16594,N_16694);
nor U22441 (N_22441,N_15947,N_15108);
or U22442 (N_22442,N_19874,N_18419);
and U22443 (N_22443,N_19601,N_18876);
nor U22444 (N_22444,N_15916,N_19259);
nor U22445 (N_22445,N_17694,N_18668);
nor U22446 (N_22446,N_17106,N_16063);
and U22447 (N_22447,N_17029,N_17967);
nor U22448 (N_22448,N_18027,N_16192);
nand U22449 (N_22449,N_19781,N_16459);
or U22450 (N_22450,N_16764,N_16866);
xnor U22451 (N_22451,N_17671,N_17168);
nor U22452 (N_22452,N_17587,N_18015);
nor U22453 (N_22453,N_15834,N_15141);
or U22454 (N_22454,N_15238,N_19651);
nand U22455 (N_22455,N_16135,N_15586);
nand U22456 (N_22456,N_16445,N_17620);
or U22457 (N_22457,N_16996,N_18077);
nand U22458 (N_22458,N_17727,N_18627);
nand U22459 (N_22459,N_17179,N_18853);
or U22460 (N_22460,N_16398,N_19144);
nor U22461 (N_22461,N_15715,N_17028);
nand U22462 (N_22462,N_18556,N_17771);
nor U22463 (N_22463,N_17373,N_17480);
nor U22464 (N_22464,N_16520,N_19941);
xnor U22465 (N_22465,N_16142,N_18237);
nor U22466 (N_22466,N_19287,N_15869);
and U22467 (N_22467,N_16148,N_15186);
nand U22468 (N_22468,N_16564,N_19727);
or U22469 (N_22469,N_16595,N_18595);
nor U22470 (N_22470,N_16874,N_18615);
nor U22471 (N_22471,N_15737,N_16227);
nand U22472 (N_22472,N_19313,N_19510);
and U22473 (N_22473,N_18439,N_15727);
and U22474 (N_22474,N_15722,N_19209);
nand U22475 (N_22475,N_15791,N_18985);
and U22476 (N_22476,N_16601,N_19726);
or U22477 (N_22477,N_15842,N_17541);
or U22478 (N_22478,N_15087,N_15532);
nand U22479 (N_22479,N_19271,N_18235);
nor U22480 (N_22480,N_19740,N_19547);
nor U22481 (N_22481,N_15879,N_17614);
or U22482 (N_22482,N_18467,N_16266);
nand U22483 (N_22483,N_19620,N_18632);
nor U22484 (N_22484,N_16096,N_16528);
and U22485 (N_22485,N_17280,N_16817);
nor U22486 (N_22486,N_15149,N_16812);
or U22487 (N_22487,N_18096,N_18234);
nor U22488 (N_22488,N_16453,N_18289);
nor U22489 (N_22489,N_15486,N_19258);
nor U22490 (N_22490,N_19817,N_16368);
or U22491 (N_22491,N_15051,N_15305);
nand U22492 (N_22492,N_15154,N_15007);
nand U22493 (N_22493,N_19552,N_17703);
nand U22494 (N_22494,N_15508,N_19146);
or U22495 (N_22495,N_18092,N_17486);
nor U22496 (N_22496,N_19916,N_15283);
nor U22497 (N_22497,N_15437,N_15184);
nand U22498 (N_22498,N_16811,N_17677);
and U22499 (N_22499,N_16340,N_16166);
xnor U22500 (N_22500,N_16949,N_16413);
nor U22501 (N_22501,N_17871,N_16268);
nand U22502 (N_22502,N_19809,N_17453);
and U22503 (N_22503,N_17019,N_17482);
nand U22504 (N_22504,N_15615,N_16762);
nor U22505 (N_22505,N_18615,N_16088);
nor U22506 (N_22506,N_17186,N_16753);
and U22507 (N_22507,N_16697,N_19776);
nor U22508 (N_22508,N_16117,N_16893);
nor U22509 (N_22509,N_17583,N_15657);
nand U22510 (N_22510,N_17588,N_16904);
nor U22511 (N_22511,N_16972,N_15811);
nand U22512 (N_22512,N_16994,N_16127);
and U22513 (N_22513,N_18356,N_18499);
nand U22514 (N_22514,N_19271,N_19671);
nor U22515 (N_22515,N_18736,N_18286);
nor U22516 (N_22516,N_19014,N_19939);
nor U22517 (N_22517,N_15155,N_15660);
nor U22518 (N_22518,N_15776,N_18738);
nor U22519 (N_22519,N_17881,N_19027);
nand U22520 (N_22520,N_17753,N_19768);
and U22521 (N_22521,N_19853,N_19158);
or U22522 (N_22522,N_17502,N_16862);
or U22523 (N_22523,N_19072,N_15208);
nand U22524 (N_22524,N_19468,N_18386);
nor U22525 (N_22525,N_19804,N_15969);
nand U22526 (N_22526,N_19843,N_19736);
or U22527 (N_22527,N_16211,N_19199);
nand U22528 (N_22528,N_17911,N_18867);
xnor U22529 (N_22529,N_17590,N_16060);
nand U22530 (N_22530,N_18222,N_17704);
or U22531 (N_22531,N_17406,N_15614);
nor U22532 (N_22532,N_19723,N_16840);
and U22533 (N_22533,N_16001,N_17362);
and U22534 (N_22534,N_17797,N_18401);
and U22535 (N_22535,N_15975,N_16585);
nor U22536 (N_22536,N_16013,N_16607);
nor U22537 (N_22537,N_16438,N_18559);
nand U22538 (N_22538,N_18460,N_15814);
or U22539 (N_22539,N_17647,N_18167);
nand U22540 (N_22540,N_18945,N_15219);
nor U22541 (N_22541,N_16786,N_17063);
nor U22542 (N_22542,N_19585,N_15816);
nand U22543 (N_22543,N_17154,N_19542);
and U22544 (N_22544,N_18315,N_17205);
nor U22545 (N_22545,N_17438,N_17302);
nand U22546 (N_22546,N_16341,N_18131);
or U22547 (N_22547,N_19351,N_19130);
and U22548 (N_22548,N_15067,N_19003);
nor U22549 (N_22549,N_17461,N_19215);
and U22550 (N_22550,N_18693,N_15211);
nand U22551 (N_22551,N_16613,N_15510);
nand U22552 (N_22552,N_17340,N_15517);
or U22553 (N_22553,N_15368,N_15885);
and U22554 (N_22554,N_15899,N_15572);
nand U22555 (N_22555,N_16010,N_19203);
or U22556 (N_22556,N_16670,N_18578);
and U22557 (N_22557,N_15667,N_19645);
and U22558 (N_22558,N_15432,N_18168);
nand U22559 (N_22559,N_19904,N_17554);
nor U22560 (N_22560,N_18718,N_18520);
xnor U22561 (N_22561,N_19651,N_15321);
nor U22562 (N_22562,N_16814,N_17523);
xor U22563 (N_22563,N_15697,N_15406);
and U22564 (N_22564,N_15582,N_19471);
and U22565 (N_22565,N_18663,N_16550);
or U22566 (N_22566,N_18110,N_17720);
nor U22567 (N_22567,N_17052,N_19405);
or U22568 (N_22568,N_19505,N_16735);
xnor U22569 (N_22569,N_15264,N_16786);
nor U22570 (N_22570,N_16468,N_17138);
nand U22571 (N_22571,N_16313,N_19499);
nor U22572 (N_22572,N_18745,N_19941);
or U22573 (N_22573,N_18567,N_16365);
nor U22574 (N_22574,N_16338,N_17980);
nor U22575 (N_22575,N_16292,N_18118);
nand U22576 (N_22576,N_15594,N_19178);
nand U22577 (N_22577,N_18493,N_19329);
and U22578 (N_22578,N_17168,N_15505);
nor U22579 (N_22579,N_16547,N_19586);
and U22580 (N_22580,N_16610,N_15591);
or U22581 (N_22581,N_15953,N_15764);
or U22582 (N_22582,N_17578,N_16443);
nand U22583 (N_22583,N_19703,N_19385);
or U22584 (N_22584,N_19501,N_15769);
nand U22585 (N_22585,N_19544,N_15688);
xnor U22586 (N_22586,N_19686,N_19228);
or U22587 (N_22587,N_16455,N_18417);
or U22588 (N_22588,N_15255,N_19158);
or U22589 (N_22589,N_17565,N_19399);
or U22590 (N_22590,N_17986,N_16949);
or U22591 (N_22591,N_17441,N_17196);
nand U22592 (N_22592,N_18332,N_17997);
nor U22593 (N_22593,N_18499,N_15194);
nor U22594 (N_22594,N_17709,N_18908);
nand U22595 (N_22595,N_17762,N_18394);
xnor U22596 (N_22596,N_19842,N_18300);
nor U22597 (N_22597,N_16016,N_19119);
nand U22598 (N_22598,N_19727,N_18368);
nand U22599 (N_22599,N_15884,N_15402);
nand U22600 (N_22600,N_17806,N_17414);
or U22601 (N_22601,N_18197,N_17518);
nand U22602 (N_22602,N_18050,N_18273);
nand U22603 (N_22603,N_19847,N_15473);
nand U22604 (N_22604,N_15371,N_17053);
nor U22605 (N_22605,N_17549,N_15841);
nor U22606 (N_22606,N_19196,N_16286);
or U22607 (N_22607,N_19553,N_16343);
nor U22608 (N_22608,N_17108,N_19699);
nand U22609 (N_22609,N_15708,N_16139);
and U22610 (N_22610,N_19769,N_15318);
or U22611 (N_22611,N_19625,N_18441);
nor U22612 (N_22612,N_18950,N_17391);
nor U22613 (N_22613,N_18502,N_15632);
nor U22614 (N_22614,N_18864,N_15311);
nand U22615 (N_22615,N_16762,N_18864);
and U22616 (N_22616,N_15292,N_18129);
nor U22617 (N_22617,N_16776,N_15147);
or U22618 (N_22618,N_18813,N_17075);
and U22619 (N_22619,N_15603,N_18521);
and U22620 (N_22620,N_15544,N_18197);
nand U22621 (N_22621,N_15697,N_17494);
nor U22622 (N_22622,N_15603,N_18720);
and U22623 (N_22623,N_18811,N_17250);
or U22624 (N_22624,N_19747,N_18573);
nor U22625 (N_22625,N_16840,N_18778);
nor U22626 (N_22626,N_15617,N_17167);
nor U22627 (N_22627,N_19352,N_18728);
nand U22628 (N_22628,N_15800,N_17014);
and U22629 (N_22629,N_18400,N_16989);
nor U22630 (N_22630,N_18990,N_16519);
nand U22631 (N_22631,N_18449,N_19351);
nor U22632 (N_22632,N_18188,N_19958);
nand U22633 (N_22633,N_19850,N_17618);
and U22634 (N_22634,N_15410,N_16189);
and U22635 (N_22635,N_19911,N_19776);
nor U22636 (N_22636,N_18899,N_17620);
nor U22637 (N_22637,N_15989,N_18012);
or U22638 (N_22638,N_17932,N_19536);
and U22639 (N_22639,N_18563,N_19249);
and U22640 (N_22640,N_18773,N_16220);
and U22641 (N_22641,N_17746,N_18242);
xnor U22642 (N_22642,N_15024,N_15430);
and U22643 (N_22643,N_16998,N_16423);
or U22644 (N_22644,N_15577,N_19216);
nand U22645 (N_22645,N_16883,N_16009);
and U22646 (N_22646,N_18260,N_18565);
and U22647 (N_22647,N_17703,N_16039);
nand U22648 (N_22648,N_19426,N_19566);
and U22649 (N_22649,N_19616,N_16045);
and U22650 (N_22650,N_16767,N_15051);
and U22651 (N_22651,N_19722,N_16534);
nand U22652 (N_22652,N_17118,N_19011);
or U22653 (N_22653,N_17847,N_18796);
or U22654 (N_22654,N_19885,N_18466);
or U22655 (N_22655,N_15355,N_17413);
and U22656 (N_22656,N_16735,N_18126);
and U22657 (N_22657,N_15173,N_19329);
and U22658 (N_22658,N_17221,N_16950);
nor U22659 (N_22659,N_18018,N_19142);
and U22660 (N_22660,N_18535,N_17281);
nand U22661 (N_22661,N_19038,N_18111);
and U22662 (N_22662,N_16857,N_18746);
or U22663 (N_22663,N_19645,N_19245);
nor U22664 (N_22664,N_17014,N_17676);
nand U22665 (N_22665,N_19942,N_17322);
xor U22666 (N_22666,N_18993,N_15349);
nor U22667 (N_22667,N_15947,N_19079);
nor U22668 (N_22668,N_16601,N_15105);
nand U22669 (N_22669,N_17929,N_15628);
or U22670 (N_22670,N_16887,N_17044);
nor U22671 (N_22671,N_17303,N_17193);
nand U22672 (N_22672,N_19318,N_15846);
or U22673 (N_22673,N_19598,N_18817);
and U22674 (N_22674,N_17842,N_19273);
nor U22675 (N_22675,N_16785,N_16164);
or U22676 (N_22676,N_19951,N_19373);
or U22677 (N_22677,N_19306,N_18032);
nor U22678 (N_22678,N_16776,N_18869);
nor U22679 (N_22679,N_19152,N_18597);
and U22680 (N_22680,N_17072,N_16230);
and U22681 (N_22681,N_15509,N_16765);
and U22682 (N_22682,N_16323,N_17916);
nor U22683 (N_22683,N_15663,N_19122);
nand U22684 (N_22684,N_17971,N_15174);
or U22685 (N_22685,N_18766,N_15746);
nand U22686 (N_22686,N_19089,N_16819);
nor U22687 (N_22687,N_17549,N_19076);
and U22688 (N_22688,N_19247,N_16739);
and U22689 (N_22689,N_19675,N_18501);
nand U22690 (N_22690,N_19619,N_18967);
nand U22691 (N_22691,N_18134,N_16502);
nor U22692 (N_22692,N_18485,N_16918);
nor U22693 (N_22693,N_19636,N_17601);
or U22694 (N_22694,N_15515,N_18561);
and U22695 (N_22695,N_16824,N_18233);
and U22696 (N_22696,N_15162,N_15732);
or U22697 (N_22697,N_16148,N_19318);
nor U22698 (N_22698,N_15182,N_17054);
nand U22699 (N_22699,N_16950,N_18880);
nor U22700 (N_22700,N_17329,N_16499);
nand U22701 (N_22701,N_17816,N_15335);
nor U22702 (N_22702,N_16126,N_18027);
or U22703 (N_22703,N_19401,N_16033);
nor U22704 (N_22704,N_17582,N_17690);
or U22705 (N_22705,N_19610,N_15362);
or U22706 (N_22706,N_15208,N_15626);
nor U22707 (N_22707,N_19330,N_15053);
nor U22708 (N_22708,N_15960,N_15745);
xor U22709 (N_22709,N_18332,N_17301);
nor U22710 (N_22710,N_18334,N_16494);
xor U22711 (N_22711,N_16293,N_16203);
or U22712 (N_22712,N_15903,N_17739);
nor U22713 (N_22713,N_18963,N_17653);
and U22714 (N_22714,N_16504,N_19576);
and U22715 (N_22715,N_19908,N_15798);
or U22716 (N_22716,N_18552,N_19421);
nand U22717 (N_22717,N_17554,N_18402);
and U22718 (N_22718,N_16793,N_18830);
nand U22719 (N_22719,N_16603,N_16919);
and U22720 (N_22720,N_16254,N_16220);
and U22721 (N_22721,N_16749,N_16625);
nor U22722 (N_22722,N_17913,N_17921);
or U22723 (N_22723,N_17581,N_19473);
nor U22724 (N_22724,N_17132,N_17592);
or U22725 (N_22725,N_15989,N_15504);
nand U22726 (N_22726,N_18971,N_19424);
or U22727 (N_22727,N_17670,N_18724);
nand U22728 (N_22728,N_18603,N_19651);
nand U22729 (N_22729,N_17066,N_16216);
xnor U22730 (N_22730,N_16056,N_19481);
or U22731 (N_22731,N_18636,N_17150);
nor U22732 (N_22732,N_16938,N_17483);
nand U22733 (N_22733,N_16732,N_16710);
or U22734 (N_22734,N_19604,N_18419);
and U22735 (N_22735,N_16121,N_17242);
and U22736 (N_22736,N_18255,N_16091);
and U22737 (N_22737,N_15480,N_19690);
nor U22738 (N_22738,N_15829,N_19605);
nor U22739 (N_22739,N_18143,N_15292);
or U22740 (N_22740,N_17499,N_17767);
nor U22741 (N_22741,N_17468,N_15582);
nor U22742 (N_22742,N_17092,N_17984);
nor U22743 (N_22743,N_17261,N_17844);
nand U22744 (N_22744,N_19814,N_16225);
nor U22745 (N_22745,N_16797,N_15124);
or U22746 (N_22746,N_15710,N_16243);
nand U22747 (N_22747,N_16086,N_15332);
or U22748 (N_22748,N_18736,N_17981);
nand U22749 (N_22749,N_16938,N_16398);
or U22750 (N_22750,N_17278,N_16910);
or U22751 (N_22751,N_16033,N_17431);
and U22752 (N_22752,N_17972,N_15336);
and U22753 (N_22753,N_16882,N_17925);
nand U22754 (N_22754,N_19669,N_19347);
or U22755 (N_22755,N_18623,N_15009);
or U22756 (N_22756,N_18963,N_17059);
nand U22757 (N_22757,N_19913,N_17293);
or U22758 (N_22758,N_15423,N_17564);
and U22759 (N_22759,N_18078,N_17410);
nand U22760 (N_22760,N_16697,N_17657);
nand U22761 (N_22761,N_19610,N_17264);
nand U22762 (N_22762,N_19833,N_15972);
nand U22763 (N_22763,N_15469,N_17793);
nor U22764 (N_22764,N_19308,N_15527);
or U22765 (N_22765,N_15723,N_19149);
or U22766 (N_22766,N_18918,N_16362);
or U22767 (N_22767,N_15654,N_16365);
xor U22768 (N_22768,N_18116,N_16650);
xnor U22769 (N_22769,N_19340,N_17424);
nand U22770 (N_22770,N_18999,N_17610);
or U22771 (N_22771,N_17725,N_16290);
xnor U22772 (N_22772,N_19760,N_16571);
nand U22773 (N_22773,N_18182,N_18487);
nor U22774 (N_22774,N_17143,N_16901);
nand U22775 (N_22775,N_19323,N_19931);
or U22776 (N_22776,N_16854,N_18022);
xnor U22777 (N_22777,N_17371,N_19254);
nor U22778 (N_22778,N_18665,N_18861);
nand U22779 (N_22779,N_17858,N_15349);
or U22780 (N_22780,N_16341,N_15311);
or U22781 (N_22781,N_17071,N_18977);
and U22782 (N_22782,N_19055,N_18778);
nand U22783 (N_22783,N_19673,N_19182);
or U22784 (N_22784,N_19426,N_15055);
nor U22785 (N_22785,N_18546,N_19011);
nand U22786 (N_22786,N_17983,N_16028);
nand U22787 (N_22787,N_16086,N_18853);
nand U22788 (N_22788,N_19722,N_15735);
or U22789 (N_22789,N_15818,N_16995);
nand U22790 (N_22790,N_18450,N_15635);
nand U22791 (N_22791,N_19788,N_15169);
nand U22792 (N_22792,N_18171,N_19085);
nand U22793 (N_22793,N_17588,N_18755);
nand U22794 (N_22794,N_18161,N_19614);
and U22795 (N_22795,N_15466,N_18333);
and U22796 (N_22796,N_15404,N_15437);
nand U22797 (N_22797,N_18308,N_17193);
nand U22798 (N_22798,N_16035,N_18508);
nand U22799 (N_22799,N_19269,N_19480);
nor U22800 (N_22800,N_16512,N_19938);
nor U22801 (N_22801,N_19258,N_15887);
nor U22802 (N_22802,N_19674,N_19349);
and U22803 (N_22803,N_18999,N_16595);
or U22804 (N_22804,N_17497,N_15774);
nand U22805 (N_22805,N_19124,N_15454);
nor U22806 (N_22806,N_16357,N_16677);
xnor U22807 (N_22807,N_19106,N_15589);
and U22808 (N_22808,N_15564,N_19050);
nor U22809 (N_22809,N_17893,N_16020);
nor U22810 (N_22810,N_18140,N_16198);
xnor U22811 (N_22811,N_15368,N_17993);
or U22812 (N_22812,N_16467,N_18839);
and U22813 (N_22813,N_17341,N_17764);
nand U22814 (N_22814,N_16796,N_17822);
nor U22815 (N_22815,N_16429,N_17656);
xor U22816 (N_22816,N_17756,N_19929);
nor U22817 (N_22817,N_16269,N_16325);
nand U22818 (N_22818,N_19377,N_15171);
or U22819 (N_22819,N_18779,N_18574);
nand U22820 (N_22820,N_19735,N_16945);
nor U22821 (N_22821,N_18110,N_16112);
nand U22822 (N_22822,N_17013,N_18840);
or U22823 (N_22823,N_15312,N_15689);
and U22824 (N_22824,N_15236,N_17796);
or U22825 (N_22825,N_17206,N_18229);
or U22826 (N_22826,N_15942,N_19256);
and U22827 (N_22827,N_17791,N_17772);
nand U22828 (N_22828,N_18945,N_17113);
nand U22829 (N_22829,N_15649,N_18921);
nor U22830 (N_22830,N_18346,N_16345);
or U22831 (N_22831,N_17862,N_16515);
nand U22832 (N_22832,N_15919,N_17123);
nand U22833 (N_22833,N_18422,N_19815);
nand U22834 (N_22834,N_18911,N_18537);
or U22835 (N_22835,N_15426,N_18800);
nor U22836 (N_22836,N_19825,N_15363);
nor U22837 (N_22837,N_15556,N_18297);
and U22838 (N_22838,N_17465,N_15300);
or U22839 (N_22839,N_19891,N_15686);
and U22840 (N_22840,N_15115,N_15112);
and U22841 (N_22841,N_18725,N_15398);
and U22842 (N_22842,N_16225,N_18437);
or U22843 (N_22843,N_15092,N_19143);
nor U22844 (N_22844,N_19533,N_17520);
nand U22845 (N_22845,N_18862,N_17313);
and U22846 (N_22846,N_16289,N_17155);
nor U22847 (N_22847,N_17285,N_15065);
and U22848 (N_22848,N_15013,N_19296);
nor U22849 (N_22849,N_17357,N_15823);
nand U22850 (N_22850,N_18428,N_15287);
or U22851 (N_22851,N_19843,N_18833);
nor U22852 (N_22852,N_16981,N_15792);
xor U22853 (N_22853,N_17994,N_18011);
nor U22854 (N_22854,N_19100,N_17411);
nand U22855 (N_22855,N_15692,N_16786);
or U22856 (N_22856,N_16111,N_18071);
nand U22857 (N_22857,N_17061,N_16124);
and U22858 (N_22858,N_19086,N_18571);
or U22859 (N_22859,N_15483,N_17520);
or U22860 (N_22860,N_16566,N_16012);
nand U22861 (N_22861,N_19599,N_19500);
and U22862 (N_22862,N_15396,N_19949);
or U22863 (N_22863,N_16856,N_19759);
or U22864 (N_22864,N_15943,N_15278);
and U22865 (N_22865,N_18223,N_15346);
nor U22866 (N_22866,N_18444,N_18014);
or U22867 (N_22867,N_17362,N_19647);
nor U22868 (N_22868,N_17722,N_18067);
nor U22869 (N_22869,N_19832,N_16538);
or U22870 (N_22870,N_19241,N_16209);
or U22871 (N_22871,N_15532,N_15324);
nor U22872 (N_22872,N_18758,N_19590);
nor U22873 (N_22873,N_16271,N_16914);
nand U22874 (N_22874,N_19867,N_19194);
nor U22875 (N_22875,N_15746,N_15355);
nand U22876 (N_22876,N_19974,N_16469);
nand U22877 (N_22877,N_19321,N_18727);
or U22878 (N_22878,N_19964,N_15687);
nand U22879 (N_22879,N_19306,N_16702);
or U22880 (N_22880,N_18467,N_18138);
or U22881 (N_22881,N_16775,N_16617);
and U22882 (N_22882,N_18426,N_15577);
or U22883 (N_22883,N_16031,N_15831);
nor U22884 (N_22884,N_15015,N_16542);
and U22885 (N_22885,N_16587,N_16558);
and U22886 (N_22886,N_19546,N_17647);
nor U22887 (N_22887,N_17813,N_19677);
and U22888 (N_22888,N_19479,N_18636);
or U22889 (N_22889,N_18380,N_17739);
nand U22890 (N_22890,N_18543,N_16167);
nor U22891 (N_22891,N_15844,N_18607);
and U22892 (N_22892,N_18281,N_15669);
and U22893 (N_22893,N_19517,N_19261);
or U22894 (N_22894,N_17463,N_15393);
nor U22895 (N_22895,N_17029,N_16294);
and U22896 (N_22896,N_19589,N_18688);
nand U22897 (N_22897,N_15717,N_19156);
and U22898 (N_22898,N_15138,N_17808);
nand U22899 (N_22899,N_15961,N_19998);
and U22900 (N_22900,N_19114,N_16466);
nor U22901 (N_22901,N_16109,N_18523);
nor U22902 (N_22902,N_19314,N_15022);
and U22903 (N_22903,N_15705,N_17296);
nand U22904 (N_22904,N_16885,N_19509);
nor U22905 (N_22905,N_15870,N_17641);
and U22906 (N_22906,N_17443,N_15844);
and U22907 (N_22907,N_16787,N_18909);
nand U22908 (N_22908,N_15490,N_17032);
nand U22909 (N_22909,N_17407,N_19062);
nor U22910 (N_22910,N_16892,N_16624);
and U22911 (N_22911,N_15482,N_16520);
or U22912 (N_22912,N_19989,N_17766);
xnor U22913 (N_22913,N_17954,N_18611);
nand U22914 (N_22914,N_16860,N_15929);
nor U22915 (N_22915,N_16226,N_15807);
nor U22916 (N_22916,N_17149,N_15726);
or U22917 (N_22917,N_15863,N_17904);
or U22918 (N_22918,N_18075,N_19274);
or U22919 (N_22919,N_19734,N_18948);
or U22920 (N_22920,N_17276,N_17475);
and U22921 (N_22921,N_19708,N_19738);
or U22922 (N_22922,N_17371,N_15265);
or U22923 (N_22923,N_16188,N_16311);
nand U22924 (N_22924,N_15302,N_16514);
nor U22925 (N_22925,N_15398,N_17981);
or U22926 (N_22926,N_17240,N_17177);
and U22927 (N_22927,N_16267,N_19715);
and U22928 (N_22928,N_15508,N_18717);
or U22929 (N_22929,N_18377,N_17723);
and U22930 (N_22930,N_17251,N_16098);
or U22931 (N_22931,N_15295,N_17566);
and U22932 (N_22932,N_19933,N_18428);
and U22933 (N_22933,N_18311,N_19130);
xnor U22934 (N_22934,N_16942,N_19336);
and U22935 (N_22935,N_17543,N_19311);
and U22936 (N_22936,N_17656,N_19136);
or U22937 (N_22937,N_19971,N_15295);
nor U22938 (N_22938,N_18135,N_15593);
nor U22939 (N_22939,N_19288,N_19981);
nor U22940 (N_22940,N_18494,N_19340);
nand U22941 (N_22941,N_16534,N_16024);
nor U22942 (N_22942,N_18067,N_18366);
nor U22943 (N_22943,N_17449,N_16893);
or U22944 (N_22944,N_15360,N_17766);
and U22945 (N_22945,N_19332,N_16685);
or U22946 (N_22946,N_16366,N_18299);
xor U22947 (N_22947,N_15734,N_17742);
or U22948 (N_22948,N_15659,N_19715);
nand U22949 (N_22949,N_18117,N_15519);
nor U22950 (N_22950,N_19918,N_19499);
or U22951 (N_22951,N_15766,N_16517);
nor U22952 (N_22952,N_19158,N_17205);
and U22953 (N_22953,N_16513,N_18319);
and U22954 (N_22954,N_16606,N_16651);
nand U22955 (N_22955,N_17804,N_18601);
nand U22956 (N_22956,N_17202,N_19700);
nand U22957 (N_22957,N_16553,N_19483);
nor U22958 (N_22958,N_19687,N_15574);
nand U22959 (N_22959,N_16799,N_18914);
and U22960 (N_22960,N_19493,N_18851);
nor U22961 (N_22961,N_18833,N_16189);
nand U22962 (N_22962,N_17739,N_16477);
nor U22963 (N_22963,N_19646,N_19448);
or U22964 (N_22964,N_17120,N_19823);
nor U22965 (N_22965,N_16810,N_17438);
nand U22966 (N_22966,N_17065,N_18974);
or U22967 (N_22967,N_15437,N_17926);
and U22968 (N_22968,N_18103,N_19878);
and U22969 (N_22969,N_15871,N_18319);
or U22970 (N_22970,N_19895,N_15637);
and U22971 (N_22971,N_15935,N_18765);
or U22972 (N_22972,N_16830,N_16717);
nor U22973 (N_22973,N_15313,N_19481);
or U22974 (N_22974,N_18762,N_16383);
nor U22975 (N_22975,N_18792,N_16464);
nand U22976 (N_22976,N_18217,N_17909);
or U22977 (N_22977,N_15309,N_15017);
xnor U22978 (N_22978,N_15854,N_16267);
nand U22979 (N_22979,N_15628,N_17843);
nor U22980 (N_22980,N_17699,N_19616);
and U22981 (N_22981,N_18507,N_15649);
or U22982 (N_22982,N_15452,N_16259);
nor U22983 (N_22983,N_17207,N_17502);
or U22984 (N_22984,N_17014,N_19831);
nand U22985 (N_22985,N_18199,N_19587);
and U22986 (N_22986,N_17323,N_17771);
and U22987 (N_22987,N_19576,N_15372);
and U22988 (N_22988,N_15122,N_18233);
nor U22989 (N_22989,N_15845,N_18812);
nor U22990 (N_22990,N_16678,N_15023);
nand U22991 (N_22991,N_19389,N_19254);
and U22992 (N_22992,N_16424,N_18644);
and U22993 (N_22993,N_17789,N_16304);
and U22994 (N_22994,N_16054,N_18494);
and U22995 (N_22995,N_17435,N_15305);
or U22996 (N_22996,N_19185,N_19055);
nand U22997 (N_22997,N_19786,N_16096);
or U22998 (N_22998,N_19865,N_17256);
and U22999 (N_22999,N_17019,N_17875);
nor U23000 (N_23000,N_16366,N_18603);
and U23001 (N_23001,N_19568,N_19054);
nor U23002 (N_23002,N_15181,N_17055);
nor U23003 (N_23003,N_16708,N_18071);
and U23004 (N_23004,N_18674,N_15547);
nand U23005 (N_23005,N_18142,N_15810);
nand U23006 (N_23006,N_18682,N_18687);
and U23007 (N_23007,N_18451,N_19604);
or U23008 (N_23008,N_17196,N_17296);
nor U23009 (N_23009,N_18724,N_15718);
nor U23010 (N_23010,N_18576,N_19160);
nor U23011 (N_23011,N_15015,N_16921);
or U23012 (N_23012,N_19757,N_15636);
nand U23013 (N_23013,N_18568,N_19149);
nor U23014 (N_23014,N_16493,N_15017);
nand U23015 (N_23015,N_15852,N_16551);
and U23016 (N_23016,N_17345,N_15075);
nand U23017 (N_23017,N_17051,N_19083);
and U23018 (N_23018,N_17830,N_17306);
and U23019 (N_23019,N_16356,N_19745);
nor U23020 (N_23020,N_19466,N_15810);
nor U23021 (N_23021,N_19591,N_16887);
and U23022 (N_23022,N_19041,N_17309);
nor U23023 (N_23023,N_17695,N_17115);
and U23024 (N_23024,N_15393,N_17612);
nor U23025 (N_23025,N_16115,N_19162);
nand U23026 (N_23026,N_16280,N_19287);
or U23027 (N_23027,N_15118,N_19148);
and U23028 (N_23028,N_16421,N_16765);
nor U23029 (N_23029,N_19179,N_18749);
nor U23030 (N_23030,N_16536,N_19517);
nor U23031 (N_23031,N_18395,N_18152);
nor U23032 (N_23032,N_19460,N_18474);
nand U23033 (N_23033,N_15623,N_16439);
nand U23034 (N_23034,N_15294,N_16038);
and U23035 (N_23035,N_16926,N_18242);
and U23036 (N_23036,N_18642,N_19530);
nor U23037 (N_23037,N_16544,N_19866);
or U23038 (N_23038,N_18258,N_16904);
and U23039 (N_23039,N_18071,N_18705);
or U23040 (N_23040,N_18721,N_18011);
nor U23041 (N_23041,N_15768,N_19962);
nor U23042 (N_23042,N_19322,N_19003);
or U23043 (N_23043,N_17748,N_19261);
nor U23044 (N_23044,N_15810,N_18000);
nand U23045 (N_23045,N_17652,N_19341);
nand U23046 (N_23046,N_15332,N_19426);
or U23047 (N_23047,N_19260,N_15556);
or U23048 (N_23048,N_17131,N_18350);
and U23049 (N_23049,N_18333,N_18858);
and U23050 (N_23050,N_18960,N_17159);
and U23051 (N_23051,N_18720,N_18414);
and U23052 (N_23052,N_19353,N_16042);
nor U23053 (N_23053,N_15698,N_18116);
nor U23054 (N_23054,N_16244,N_16325);
nand U23055 (N_23055,N_17048,N_17296);
or U23056 (N_23056,N_19835,N_17189);
xnor U23057 (N_23057,N_15579,N_16909);
or U23058 (N_23058,N_15638,N_18603);
nor U23059 (N_23059,N_17271,N_15241);
xnor U23060 (N_23060,N_17267,N_17402);
nand U23061 (N_23061,N_15481,N_16174);
and U23062 (N_23062,N_17168,N_16360);
nor U23063 (N_23063,N_17502,N_19010);
nand U23064 (N_23064,N_15767,N_17737);
and U23065 (N_23065,N_16639,N_18697);
nor U23066 (N_23066,N_16413,N_16350);
and U23067 (N_23067,N_17219,N_17428);
or U23068 (N_23068,N_19870,N_16723);
xor U23069 (N_23069,N_18051,N_19104);
nand U23070 (N_23070,N_17970,N_18185);
and U23071 (N_23071,N_16623,N_19535);
and U23072 (N_23072,N_19699,N_19426);
or U23073 (N_23073,N_17573,N_16254);
nor U23074 (N_23074,N_17862,N_15738);
or U23075 (N_23075,N_17594,N_16247);
nand U23076 (N_23076,N_18980,N_15998);
nor U23077 (N_23077,N_16375,N_17460);
nor U23078 (N_23078,N_17801,N_15062);
xor U23079 (N_23079,N_16008,N_16220);
or U23080 (N_23080,N_17356,N_15614);
or U23081 (N_23081,N_19785,N_15246);
and U23082 (N_23082,N_19014,N_16217);
nand U23083 (N_23083,N_16080,N_17200);
and U23084 (N_23084,N_19201,N_18961);
nor U23085 (N_23085,N_19788,N_18718);
and U23086 (N_23086,N_19888,N_19456);
or U23087 (N_23087,N_16436,N_15769);
nand U23088 (N_23088,N_15375,N_16004);
nand U23089 (N_23089,N_17619,N_16503);
and U23090 (N_23090,N_15503,N_16058);
nor U23091 (N_23091,N_19303,N_18826);
or U23092 (N_23092,N_19192,N_16277);
nor U23093 (N_23093,N_17939,N_19230);
nor U23094 (N_23094,N_16784,N_17581);
or U23095 (N_23095,N_18465,N_15179);
nand U23096 (N_23096,N_18563,N_15973);
nor U23097 (N_23097,N_19530,N_16672);
or U23098 (N_23098,N_19106,N_15677);
nand U23099 (N_23099,N_17034,N_18904);
or U23100 (N_23100,N_15325,N_19061);
and U23101 (N_23101,N_15473,N_15883);
and U23102 (N_23102,N_18550,N_19450);
and U23103 (N_23103,N_16974,N_17709);
nor U23104 (N_23104,N_18699,N_15586);
or U23105 (N_23105,N_17827,N_15067);
xnor U23106 (N_23106,N_17609,N_17593);
and U23107 (N_23107,N_15621,N_15542);
or U23108 (N_23108,N_16375,N_17333);
nand U23109 (N_23109,N_15632,N_16269);
and U23110 (N_23110,N_17622,N_15109);
or U23111 (N_23111,N_15517,N_16759);
nand U23112 (N_23112,N_15399,N_17908);
nor U23113 (N_23113,N_16459,N_15755);
or U23114 (N_23114,N_15356,N_17480);
xnor U23115 (N_23115,N_16532,N_15735);
and U23116 (N_23116,N_19097,N_16007);
nand U23117 (N_23117,N_19592,N_15762);
nor U23118 (N_23118,N_15353,N_18550);
nand U23119 (N_23119,N_19132,N_18227);
or U23120 (N_23120,N_15653,N_15680);
nor U23121 (N_23121,N_19984,N_16853);
and U23122 (N_23122,N_15149,N_19742);
and U23123 (N_23123,N_18930,N_16106);
nand U23124 (N_23124,N_17198,N_16719);
nor U23125 (N_23125,N_15420,N_17587);
nor U23126 (N_23126,N_17161,N_15203);
xnor U23127 (N_23127,N_17356,N_16828);
nor U23128 (N_23128,N_15682,N_18301);
xnor U23129 (N_23129,N_16209,N_18831);
nor U23130 (N_23130,N_19622,N_17909);
nor U23131 (N_23131,N_19514,N_17139);
or U23132 (N_23132,N_15528,N_16886);
xor U23133 (N_23133,N_15571,N_19925);
and U23134 (N_23134,N_15048,N_17322);
nand U23135 (N_23135,N_18986,N_16685);
xor U23136 (N_23136,N_15559,N_16563);
xor U23137 (N_23137,N_16696,N_15877);
or U23138 (N_23138,N_16040,N_15787);
nand U23139 (N_23139,N_15870,N_18128);
or U23140 (N_23140,N_15327,N_16232);
or U23141 (N_23141,N_18312,N_17736);
or U23142 (N_23142,N_15710,N_17621);
and U23143 (N_23143,N_15442,N_17820);
and U23144 (N_23144,N_17788,N_16293);
nand U23145 (N_23145,N_19680,N_18031);
nor U23146 (N_23146,N_17664,N_15063);
and U23147 (N_23147,N_15395,N_18721);
or U23148 (N_23148,N_17290,N_18709);
nand U23149 (N_23149,N_19351,N_15813);
or U23150 (N_23150,N_18020,N_16388);
and U23151 (N_23151,N_18806,N_15721);
nor U23152 (N_23152,N_18424,N_18369);
nor U23153 (N_23153,N_16578,N_16716);
nor U23154 (N_23154,N_19405,N_15835);
or U23155 (N_23155,N_16956,N_16716);
or U23156 (N_23156,N_16921,N_16892);
nor U23157 (N_23157,N_16089,N_18193);
or U23158 (N_23158,N_15487,N_18939);
nor U23159 (N_23159,N_18754,N_19256);
nand U23160 (N_23160,N_16397,N_18701);
and U23161 (N_23161,N_19599,N_19541);
nor U23162 (N_23162,N_16479,N_15512);
nand U23163 (N_23163,N_15711,N_19857);
and U23164 (N_23164,N_17201,N_16401);
and U23165 (N_23165,N_16187,N_17659);
or U23166 (N_23166,N_16294,N_18291);
or U23167 (N_23167,N_18580,N_19988);
and U23168 (N_23168,N_18539,N_18397);
or U23169 (N_23169,N_15217,N_19398);
nand U23170 (N_23170,N_17463,N_15143);
nor U23171 (N_23171,N_17069,N_19606);
nand U23172 (N_23172,N_16464,N_15882);
nor U23173 (N_23173,N_15318,N_16204);
or U23174 (N_23174,N_18759,N_17451);
nor U23175 (N_23175,N_18714,N_16441);
or U23176 (N_23176,N_15452,N_18399);
nor U23177 (N_23177,N_18907,N_18073);
xor U23178 (N_23178,N_18151,N_18531);
and U23179 (N_23179,N_19587,N_19356);
nand U23180 (N_23180,N_18142,N_17027);
and U23181 (N_23181,N_17229,N_17878);
or U23182 (N_23182,N_15565,N_16544);
xor U23183 (N_23183,N_16560,N_17157);
and U23184 (N_23184,N_16140,N_19314);
nand U23185 (N_23185,N_15603,N_18177);
or U23186 (N_23186,N_16894,N_16342);
and U23187 (N_23187,N_16831,N_18388);
nor U23188 (N_23188,N_16075,N_18372);
xor U23189 (N_23189,N_18859,N_15233);
or U23190 (N_23190,N_17648,N_15725);
or U23191 (N_23191,N_19601,N_19489);
and U23192 (N_23192,N_18085,N_15827);
nand U23193 (N_23193,N_17303,N_17903);
nand U23194 (N_23194,N_15849,N_17026);
nor U23195 (N_23195,N_15882,N_19565);
nor U23196 (N_23196,N_16790,N_17900);
or U23197 (N_23197,N_18922,N_16976);
nor U23198 (N_23198,N_15403,N_19907);
or U23199 (N_23199,N_19977,N_17610);
nor U23200 (N_23200,N_16364,N_19755);
and U23201 (N_23201,N_16692,N_17571);
and U23202 (N_23202,N_17474,N_18193);
nand U23203 (N_23203,N_19179,N_16121);
or U23204 (N_23204,N_18923,N_17548);
or U23205 (N_23205,N_15006,N_19280);
nand U23206 (N_23206,N_16338,N_19126);
nor U23207 (N_23207,N_19209,N_17006);
or U23208 (N_23208,N_16837,N_17347);
nor U23209 (N_23209,N_19489,N_17510);
or U23210 (N_23210,N_16920,N_15076);
nor U23211 (N_23211,N_19036,N_17878);
nor U23212 (N_23212,N_16605,N_16220);
nand U23213 (N_23213,N_19523,N_16921);
nand U23214 (N_23214,N_16186,N_15651);
nand U23215 (N_23215,N_19220,N_16334);
and U23216 (N_23216,N_16906,N_18097);
nor U23217 (N_23217,N_17246,N_17983);
nand U23218 (N_23218,N_15848,N_19672);
or U23219 (N_23219,N_18638,N_15825);
nand U23220 (N_23220,N_18524,N_16001);
nand U23221 (N_23221,N_18134,N_15671);
xor U23222 (N_23222,N_18193,N_16922);
and U23223 (N_23223,N_16070,N_17971);
nand U23224 (N_23224,N_15217,N_19271);
or U23225 (N_23225,N_19203,N_18113);
nor U23226 (N_23226,N_19551,N_18441);
nor U23227 (N_23227,N_15636,N_19909);
nand U23228 (N_23228,N_17910,N_19271);
or U23229 (N_23229,N_15372,N_19015);
nand U23230 (N_23230,N_16024,N_15606);
and U23231 (N_23231,N_17795,N_18833);
nor U23232 (N_23232,N_16274,N_18644);
or U23233 (N_23233,N_16130,N_17930);
nand U23234 (N_23234,N_15913,N_15713);
or U23235 (N_23235,N_19259,N_16483);
nand U23236 (N_23236,N_19960,N_18673);
nand U23237 (N_23237,N_18677,N_19487);
nor U23238 (N_23238,N_15824,N_16328);
nand U23239 (N_23239,N_15173,N_15310);
or U23240 (N_23240,N_19100,N_16390);
and U23241 (N_23241,N_15454,N_15683);
and U23242 (N_23242,N_16542,N_16403);
nor U23243 (N_23243,N_18520,N_17895);
and U23244 (N_23244,N_18582,N_15346);
nand U23245 (N_23245,N_16891,N_15636);
and U23246 (N_23246,N_17262,N_15790);
and U23247 (N_23247,N_17194,N_16120);
or U23248 (N_23248,N_17042,N_16684);
nor U23249 (N_23249,N_16169,N_16161);
nor U23250 (N_23250,N_18838,N_17667);
nand U23251 (N_23251,N_16844,N_15302);
nor U23252 (N_23252,N_19658,N_16720);
or U23253 (N_23253,N_17115,N_16917);
or U23254 (N_23254,N_17407,N_16502);
nor U23255 (N_23255,N_18943,N_18233);
nand U23256 (N_23256,N_19740,N_17927);
or U23257 (N_23257,N_15388,N_17768);
and U23258 (N_23258,N_19655,N_16343);
nand U23259 (N_23259,N_19938,N_19082);
nor U23260 (N_23260,N_18558,N_18780);
or U23261 (N_23261,N_16140,N_16770);
and U23262 (N_23262,N_15829,N_15076);
or U23263 (N_23263,N_15668,N_15540);
nand U23264 (N_23264,N_15053,N_16515);
and U23265 (N_23265,N_15027,N_16680);
or U23266 (N_23266,N_17469,N_19977);
or U23267 (N_23267,N_17106,N_17287);
nor U23268 (N_23268,N_18274,N_18107);
xor U23269 (N_23269,N_16150,N_17846);
nor U23270 (N_23270,N_15597,N_15003);
or U23271 (N_23271,N_16345,N_16266);
nor U23272 (N_23272,N_17230,N_18716);
nor U23273 (N_23273,N_18055,N_16107);
or U23274 (N_23274,N_19500,N_19027);
nand U23275 (N_23275,N_19082,N_16851);
nand U23276 (N_23276,N_17974,N_15152);
nor U23277 (N_23277,N_17840,N_19766);
or U23278 (N_23278,N_19078,N_16921);
and U23279 (N_23279,N_18463,N_18156);
nand U23280 (N_23280,N_17888,N_16822);
and U23281 (N_23281,N_19500,N_19810);
and U23282 (N_23282,N_17918,N_16211);
or U23283 (N_23283,N_19164,N_15716);
and U23284 (N_23284,N_16438,N_19522);
nand U23285 (N_23285,N_19060,N_16193);
nand U23286 (N_23286,N_18701,N_15932);
nand U23287 (N_23287,N_19295,N_17760);
nand U23288 (N_23288,N_19733,N_18427);
and U23289 (N_23289,N_17433,N_16573);
or U23290 (N_23290,N_16316,N_16031);
nor U23291 (N_23291,N_19823,N_16322);
or U23292 (N_23292,N_16030,N_19895);
nor U23293 (N_23293,N_18187,N_16110);
and U23294 (N_23294,N_19140,N_15328);
nor U23295 (N_23295,N_18025,N_15124);
or U23296 (N_23296,N_16976,N_19634);
or U23297 (N_23297,N_15864,N_15069);
nand U23298 (N_23298,N_15174,N_19022);
nor U23299 (N_23299,N_16733,N_18726);
nand U23300 (N_23300,N_15512,N_18511);
and U23301 (N_23301,N_16024,N_17505);
nor U23302 (N_23302,N_19159,N_17401);
nand U23303 (N_23303,N_17662,N_18608);
and U23304 (N_23304,N_18428,N_17438);
nor U23305 (N_23305,N_17682,N_17993);
or U23306 (N_23306,N_16317,N_15666);
nand U23307 (N_23307,N_16977,N_15477);
and U23308 (N_23308,N_17507,N_16477);
and U23309 (N_23309,N_17162,N_18221);
and U23310 (N_23310,N_16379,N_15033);
and U23311 (N_23311,N_19251,N_15595);
and U23312 (N_23312,N_17782,N_18608);
nand U23313 (N_23313,N_16330,N_19266);
nor U23314 (N_23314,N_16744,N_15214);
or U23315 (N_23315,N_18346,N_18136);
xor U23316 (N_23316,N_16851,N_16490);
and U23317 (N_23317,N_17226,N_18552);
nor U23318 (N_23318,N_16931,N_19580);
and U23319 (N_23319,N_17023,N_15429);
and U23320 (N_23320,N_16768,N_16457);
nand U23321 (N_23321,N_19855,N_15792);
and U23322 (N_23322,N_19019,N_19510);
nor U23323 (N_23323,N_16064,N_19369);
and U23324 (N_23324,N_19781,N_17549);
nor U23325 (N_23325,N_18400,N_19633);
and U23326 (N_23326,N_18835,N_18756);
nor U23327 (N_23327,N_18143,N_18183);
nor U23328 (N_23328,N_19356,N_19142);
or U23329 (N_23329,N_16707,N_18967);
and U23330 (N_23330,N_15288,N_15039);
nand U23331 (N_23331,N_18367,N_15564);
and U23332 (N_23332,N_16615,N_17901);
nand U23333 (N_23333,N_16520,N_16589);
nand U23334 (N_23334,N_16879,N_16866);
and U23335 (N_23335,N_17719,N_15348);
or U23336 (N_23336,N_19072,N_15347);
or U23337 (N_23337,N_15754,N_17363);
or U23338 (N_23338,N_17812,N_19671);
nor U23339 (N_23339,N_16334,N_17923);
nand U23340 (N_23340,N_17576,N_19570);
or U23341 (N_23341,N_15331,N_18457);
nand U23342 (N_23342,N_15427,N_15428);
and U23343 (N_23343,N_18588,N_16377);
or U23344 (N_23344,N_16091,N_18853);
or U23345 (N_23345,N_15543,N_19861);
nand U23346 (N_23346,N_19899,N_15291);
and U23347 (N_23347,N_19118,N_19710);
nor U23348 (N_23348,N_18281,N_18836);
nor U23349 (N_23349,N_17434,N_19794);
nor U23350 (N_23350,N_19541,N_16233);
nor U23351 (N_23351,N_18208,N_18259);
or U23352 (N_23352,N_18147,N_18751);
and U23353 (N_23353,N_17975,N_19864);
and U23354 (N_23354,N_16542,N_17157);
nand U23355 (N_23355,N_17576,N_17648);
and U23356 (N_23356,N_17185,N_17078);
nand U23357 (N_23357,N_17444,N_15076);
xor U23358 (N_23358,N_15377,N_18861);
nor U23359 (N_23359,N_15109,N_18121);
or U23360 (N_23360,N_18392,N_17597);
nand U23361 (N_23361,N_18257,N_19919);
xor U23362 (N_23362,N_19827,N_17905);
and U23363 (N_23363,N_16027,N_18194);
nand U23364 (N_23364,N_17849,N_18291);
nor U23365 (N_23365,N_17606,N_16541);
nand U23366 (N_23366,N_15844,N_17581);
nand U23367 (N_23367,N_16327,N_19457);
and U23368 (N_23368,N_19095,N_16987);
and U23369 (N_23369,N_19926,N_19249);
nand U23370 (N_23370,N_17202,N_15574);
and U23371 (N_23371,N_18436,N_19541);
nor U23372 (N_23372,N_17483,N_17929);
and U23373 (N_23373,N_19307,N_18606);
nor U23374 (N_23374,N_17935,N_17895);
nor U23375 (N_23375,N_17390,N_16838);
nand U23376 (N_23376,N_18978,N_18507);
or U23377 (N_23377,N_19201,N_16041);
or U23378 (N_23378,N_19040,N_19382);
nor U23379 (N_23379,N_17444,N_17734);
or U23380 (N_23380,N_17182,N_17001);
nor U23381 (N_23381,N_15590,N_19561);
and U23382 (N_23382,N_15648,N_15303);
nand U23383 (N_23383,N_19049,N_15455);
xnor U23384 (N_23384,N_17664,N_15785);
or U23385 (N_23385,N_17810,N_17424);
nand U23386 (N_23386,N_17050,N_18520);
nand U23387 (N_23387,N_16856,N_15082);
nor U23388 (N_23388,N_18606,N_15573);
nor U23389 (N_23389,N_15554,N_19110);
or U23390 (N_23390,N_18314,N_17120);
and U23391 (N_23391,N_19970,N_17083);
or U23392 (N_23392,N_18735,N_16990);
nand U23393 (N_23393,N_17348,N_15172);
and U23394 (N_23394,N_18485,N_17938);
nor U23395 (N_23395,N_17155,N_18067);
nand U23396 (N_23396,N_17543,N_17576);
and U23397 (N_23397,N_18249,N_16183);
and U23398 (N_23398,N_16986,N_18598);
and U23399 (N_23399,N_19296,N_18453);
or U23400 (N_23400,N_17327,N_19024);
and U23401 (N_23401,N_15740,N_19376);
nand U23402 (N_23402,N_15980,N_18750);
or U23403 (N_23403,N_16099,N_16323);
nand U23404 (N_23404,N_17048,N_19028);
nor U23405 (N_23405,N_18921,N_16648);
nor U23406 (N_23406,N_19481,N_19140);
nand U23407 (N_23407,N_16075,N_19152);
xor U23408 (N_23408,N_17694,N_15553);
or U23409 (N_23409,N_17023,N_19553);
nand U23410 (N_23410,N_16883,N_18407);
or U23411 (N_23411,N_19816,N_15259);
nor U23412 (N_23412,N_16065,N_15064);
and U23413 (N_23413,N_18029,N_15251);
or U23414 (N_23414,N_18276,N_16665);
or U23415 (N_23415,N_18016,N_17825);
nand U23416 (N_23416,N_18804,N_18622);
nand U23417 (N_23417,N_18714,N_18394);
and U23418 (N_23418,N_16520,N_16880);
nand U23419 (N_23419,N_18522,N_15352);
and U23420 (N_23420,N_17980,N_18207);
or U23421 (N_23421,N_17482,N_19058);
and U23422 (N_23422,N_18621,N_15123);
or U23423 (N_23423,N_17284,N_17383);
nor U23424 (N_23424,N_16411,N_15143);
nor U23425 (N_23425,N_17538,N_17310);
nand U23426 (N_23426,N_16883,N_16587);
nor U23427 (N_23427,N_15238,N_18843);
nand U23428 (N_23428,N_18542,N_17432);
nor U23429 (N_23429,N_15998,N_15808);
nand U23430 (N_23430,N_16826,N_18180);
nand U23431 (N_23431,N_15413,N_16037);
or U23432 (N_23432,N_15689,N_18298);
nor U23433 (N_23433,N_18490,N_17387);
or U23434 (N_23434,N_19979,N_17253);
or U23435 (N_23435,N_18217,N_19427);
nand U23436 (N_23436,N_17967,N_15602);
or U23437 (N_23437,N_15669,N_17700);
or U23438 (N_23438,N_19322,N_18687);
or U23439 (N_23439,N_16086,N_19058);
nand U23440 (N_23440,N_15048,N_18565);
or U23441 (N_23441,N_18878,N_19382);
nor U23442 (N_23442,N_17353,N_16316);
nor U23443 (N_23443,N_18714,N_16361);
nor U23444 (N_23444,N_19156,N_17931);
and U23445 (N_23445,N_19204,N_16966);
nor U23446 (N_23446,N_19081,N_17812);
nor U23447 (N_23447,N_15978,N_15495);
nand U23448 (N_23448,N_19152,N_16871);
nor U23449 (N_23449,N_15000,N_16533);
or U23450 (N_23450,N_17233,N_18422);
and U23451 (N_23451,N_18763,N_15495);
or U23452 (N_23452,N_16188,N_17668);
nand U23453 (N_23453,N_18172,N_15827);
and U23454 (N_23454,N_15155,N_18827);
or U23455 (N_23455,N_16095,N_15320);
nand U23456 (N_23456,N_15495,N_15290);
and U23457 (N_23457,N_15757,N_15641);
nor U23458 (N_23458,N_16530,N_18732);
nand U23459 (N_23459,N_19964,N_15199);
or U23460 (N_23460,N_18390,N_16083);
and U23461 (N_23461,N_18866,N_19958);
and U23462 (N_23462,N_18036,N_18231);
or U23463 (N_23463,N_15366,N_18159);
and U23464 (N_23464,N_18727,N_16878);
nand U23465 (N_23465,N_18938,N_16053);
or U23466 (N_23466,N_19146,N_16729);
nor U23467 (N_23467,N_19317,N_18564);
or U23468 (N_23468,N_17103,N_19493);
and U23469 (N_23469,N_19272,N_18433);
nand U23470 (N_23470,N_19844,N_17503);
nand U23471 (N_23471,N_18152,N_18793);
nor U23472 (N_23472,N_15342,N_19421);
nor U23473 (N_23473,N_17836,N_18001);
nor U23474 (N_23474,N_17624,N_19929);
or U23475 (N_23475,N_19147,N_17298);
or U23476 (N_23476,N_17675,N_16474);
and U23477 (N_23477,N_16025,N_16241);
and U23478 (N_23478,N_18040,N_18044);
and U23479 (N_23479,N_17802,N_15709);
or U23480 (N_23480,N_18311,N_19251);
nand U23481 (N_23481,N_16185,N_19605);
nor U23482 (N_23482,N_19255,N_16533);
and U23483 (N_23483,N_19348,N_19055);
nor U23484 (N_23484,N_19235,N_19676);
nand U23485 (N_23485,N_19107,N_15503);
nand U23486 (N_23486,N_15269,N_16701);
or U23487 (N_23487,N_15916,N_19657);
or U23488 (N_23488,N_15905,N_17880);
and U23489 (N_23489,N_15050,N_16412);
or U23490 (N_23490,N_16107,N_19880);
nand U23491 (N_23491,N_16549,N_17291);
or U23492 (N_23492,N_17894,N_17684);
nand U23493 (N_23493,N_17382,N_19276);
nor U23494 (N_23494,N_18515,N_18600);
or U23495 (N_23495,N_15053,N_17537);
and U23496 (N_23496,N_18735,N_16532);
xor U23497 (N_23497,N_16469,N_15270);
and U23498 (N_23498,N_19734,N_15809);
nor U23499 (N_23499,N_15767,N_18830);
nand U23500 (N_23500,N_16471,N_16313);
or U23501 (N_23501,N_16273,N_17680);
or U23502 (N_23502,N_17237,N_15652);
and U23503 (N_23503,N_16692,N_19734);
and U23504 (N_23504,N_18513,N_16623);
nand U23505 (N_23505,N_15429,N_19489);
nand U23506 (N_23506,N_19505,N_15382);
nor U23507 (N_23507,N_18258,N_15496);
nor U23508 (N_23508,N_18790,N_19796);
and U23509 (N_23509,N_17069,N_16865);
nand U23510 (N_23510,N_15862,N_18061);
xnor U23511 (N_23511,N_19552,N_18166);
nand U23512 (N_23512,N_16043,N_17124);
nor U23513 (N_23513,N_16607,N_16799);
or U23514 (N_23514,N_19116,N_18649);
nor U23515 (N_23515,N_16195,N_15658);
and U23516 (N_23516,N_17622,N_19460);
nor U23517 (N_23517,N_17622,N_19828);
nor U23518 (N_23518,N_19289,N_17715);
and U23519 (N_23519,N_19793,N_18352);
nor U23520 (N_23520,N_19748,N_16718);
and U23521 (N_23521,N_19095,N_18808);
and U23522 (N_23522,N_18011,N_19534);
nor U23523 (N_23523,N_19649,N_17763);
nand U23524 (N_23524,N_19866,N_16316);
and U23525 (N_23525,N_19419,N_15949);
or U23526 (N_23526,N_18463,N_15162);
nor U23527 (N_23527,N_18582,N_18341);
or U23528 (N_23528,N_18299,N_15468);
or U23529 (N_23529,N_17918,N_15780);
nor U23530 (N_23530,N_18891,N_15893);
nor U23531 (N_23531,N_15272,N_16414);
and U23532 (N_23532,N_17063,N_17237);
and U23533 (N_23533,N_17600,N_18032);
or U23534 (N_23534,N_19432,N_15222);
or U23535 (N_23535,N_15060,N_17459);
or U23536 (N_23536,N_19572,N_19393);
nor U23537 (N_23537,N_15909,N_16595);
nor U23538 (N_23538,N_18865,N_15191);
nor U23539 (N_23539,N_18420,N_15812);
nand U23540 (N_23540,N_17392,N_17239);
nor U23541 (N_23541,N_17242,N_16735);
or U23542 (N_23542,N_17963,N_16811);
or U23543 (N_23543,N_19762,N_18556);
nor U23544 (N_23544,N_18703,N_17712);
and U23545 (N_23545,N_17773,N_18277);
nand U23546 (N_23546,N_19490,N_19998);
and U23547 (N_23547,N_17626,N_16416);
nand U23548 (N_23548,N_17134,N_18033);
or U23549 (N_23549,N_18800,N_17649);
or U23550 (N_23550,N_17532,N_18331);
and U23551 (N_23551,N_18799,N_18562);
and U23552 (N_23552,N_17718,N_18026);
and U23553 (N_23553,N_19690,N_18154);
xor U23554 (N_23554,N_19627,N_19684);
nand U23555 (N_23555,N_18477,N_16444);
or U23556 (N_23556,N_19144,N_17516);
and U23557 (N_23557,N_16144,N_18744);
or U23558 (N_23558,N_17057,N_17073);
xor U23559 (N_23559,N_15610,N_19188);
nor U23560 (N_23560,N_16621,N_17680);
and U23561 (N_23561,N_15389,N_18645);
and U23562 (N_23562,N_16281,N_16401);
nor U23563 (N_23563,N_16131,N_16929);
nand U23564 (N_23564,N_15543,N_16698);
nor U23565 (N_23565,N_18778,N_17839);
nor U23566 (N_23566,N_19446,N_18679);
and U23567 (N_23567,N_18428,N_16183);
or U23568 (N_23568,N_15617,N_18545);
nand U23569 (N_23569,N_17060,N_18673);
nand U23570 (N_23570,N_19907,N_18175);
or U23571 (N_23571,N_16191,N_19151);
and U23572 (N_23572,N_19557,N_15998);
xor U23573 (N_23573,N_19233,N_19193);
nand U23574 (N_23574,N_17180,N_16800);
and U23575 (N_23575,N_18906,N_17186);
nor U23576 (N_23576,N_16297,N_18140);
nor U23577 (N_23577,N_16323,N_16453);
nor U23578 (N_23578,N_19599,N_19458);
or U23579 (N_23579,N_18792,N_16768);
nor U23580 (N_23580,N_16772,N_16196);
nand U23581 (N_23581,N_18629,N_15295);
and U23582 (N_23582,N_19671,N_18177);
or U23583 (N_23583,N_17102,N_18882);
or U23584 (N_23584,N_16356,N_16335);
nand U23585 (N_23585,N_15656,N_17580);
or U23586 (N_23586,N_17918,N_19900);
or U23587 (N_23587,N_17887,N_15610);
nor U23588 (N_23588,N_16898,N_18318);
and U23589 (N_23589,N_18833,N_16336);
nand U23590 (N_23590,N_16314,N_17655);
nor U23591 (N_23591,N_16654,N_17632);
nor U23592 (N_23592,N_17999,N_17117);
or U23593 (N_23593,N_15666,N_16669);
nand U23594 (N_23594,N_16840,N_18804);
nor U23595 (N_23595,N_15919,N_17223);
nor U23596 (N_23596,N_19366,N_15663);
nor U23597 (N_23597,N_16291,N_16998);
nor U23598 (N_23598,N_17066,N_15389);
and U23599 (N_23599,N_15007,N_15368);
and U23600 (N_23600,N_17742,N_16459);
or U23601 (N_23601,N_16028,N_15363);
and U23602 (N_23602,N_17253,N_16807);
nand U23603 (N_23603,N_17144,N_16172);
nand U23604 (N_23604,N_16978,N_17274);
or U23605 (N_23605,N_17932,N_15090);
nand U23606 (N_23606,N_15800,N_15022);
nand U23607 (N_23607,N_18078,N_18056);
and U23608 (N_23608,N_16266,N_15449);
and U23609 (N_23609,N_17484,N_18836);
or U23610 (N_23610,N_19930,N_15765);
nand U23611 (N_23611,N_17936,N_16975);
or U23612 (N_23612,N_16478,N_19637);
nor U23613 (N_23613,N_15776,N_16389);
nor U23614 (N_23614,N_17975,N_19076);
or U23615 (N_23615,N_17096,N_18382);
nor U23616 (N_23616,N_15923,N_18924);
nand U23617 (N_23617,N_16276,N_18691);
xnor U23618 (N_23618,N_18094,N_19759);
nand U23619 (N_23619,N_15265,N_15453);
nand U23620 (N_23620,N_16179,N_16437);
nand U23621 (N_23621,N_18531,N_15594);
and U23622 (N_23622,N_15956,N_16517);
or U23623 (N_23623,N_15227,N_19605);
nor U23624 (N_23624,N_18830,N_15107);
and U23625 (N_23625,N_19499,N_16365);
or U23626 (N_23626,N_16728,N_18496);
and U23627 (N_23627,N_17702,N_18615);
nor U23628 (N_23628,N_15083,N_17819);
nor U23629 (N_23629,N_15693,N_18893);
nand U23630 (N_23630,N_18729,N_17981);
nand U23631 (N_23631,N_16298,N_16836);
nand U23632 (N_23632,N_19081,N_16779);
nand U23633 (N_23633,N_19274,N_19137);
nor U23634 (N_23634,N_19557,N_17333);
and U23635 (N_23635,N_16846,N_16327);
or U23636 (N_23636,N_19549,N_19623);
nor U23637 (N_23637,N_15988,N_17121);
nor U23638 (N_23638,N_15236,N_17586);
or U23639 (N_23639,N_16859,N_18948);
nand U23640 (N_23640,N_16060,N_19133);
or U23641 (N_23641,N_19519,N_19584);
or U23642 (N_23642,N_17161,N_17432);
and U23643 (N_23643,N_18836,N_19833);
or U23644 (N_23644,N_15316,N_15028);
or U23645 (N_23645,N_17828,N_19039);
and U23646 (N_23646,N_18270,N_19416);
or U23647 (N_23647,N_18862,N_16692);
nor U23648 (N_23648,N_18441,N_18353);
and U23649 (N_23649,N_15051,N_15598);
nand U23650 (N_23650,N_19003,N_16301);
nor U23651 (N_23651,N_18078,N_19536);
and U23652 (N_23652,N_15639,N_18251);
nor U23653 (N_23653,N_18505,N_17208);
nor U23654 (N_23654,N_15566,N_17953);
or U23655 (N_23655,N_17490,N_19468);
or U23656 (N_23656,N_15449,N_18222);
nor U23657 (N_23657,N_17217,N_17447);
nand U23658 (N_23658,N_16783,N_16967);
nand U23659 (N_23659,N_18133,N_15264);
nand U23660 (N_23660,N_19571,N_16572);
nand U23661 (N_23661,N_16217,N_17957);
and U23662 (N_23662,N_17449,N_19559);
nor U23663 (N_23663,N_15692,N_15939);
or U23664 (N_23664,N_15204,N_15674);
nor U23665 (N_23665,N_15291,N_15399);
and U23666 (N_23666,N_18281,N_19134);
and U23667 (N_23667,N_16827,N_18843);
xor U23668 (N_23668,N_16020,N_19405);
and U23669 (N_23669,N_18055,N_16481);
or U23670 (N_23670,N_15586,N_15604);
nor U23671 (N_23671,N_18470,N_17078);
and U23672 (N_23672,N_16775,N_19567);
nand U23673 (N_23673,N_15513,N_16157);
nand U23674 (N_23674,N_17091,N_17068);
nand U23675 (N_23675,N_17128,N_15480);
nand U23676 (N_23676,N_16225,N_18593);
or U23677 (N_23677,N_15214,N_18192);
nand U23678 (N_23678,N_19885,N_16275);
or U23679 (N_23679,N_18835,N_17329);
and U23680 (N_23680,N_15280,N_15597);
and U23681 (N_23681,N_16451,N_16163);
or U23682 (N_23682,N_19266,N_19358);
and U23683 (N_23683,N_18081,N_16529);
nor U23684 (N_23684,N_15566,N_16443);
xor U23685 (N_23685,N_19857,N_17574);
and U23686 (N_23686,N_15837,N_18096);
and U23687 (N_23687,N_18439,N_15264);
nor U23688 (N_23688,N_18824,N_17359);
nand U23689 (N_23689,N_18270,N_19947);
or U23690 (N_23690,N_17850,N_16947);
xnor U23691 (N_23691,N_16856,N_19584);
nand U23692 (N_23692,N_18011,N_18617);
or U23693 (N_23693,N_15213,N_19037);
nor U23694 (N_23694,N_17163,N_16918);
and U23695 (N_23695,N_18168,N_18928);
or U23696 (N_23696,N_16216,N_19688);
and U23697 (N_23697,N_15426,N_19323);
and U23698 (N_23698,N_15915,N_18908);
and U23699 (N_23699,N_18914,N_18636);
nand U23700 (N_23700,N_15201,N_17926);
nor U23701 (N_23701,N_15370,N_17743);
nor U23702 (N_23702,N_18518,N_15600);
nand U23703 (N_23703,N_17635,N_15187);
or U23704 (N_23704,N_16803,N_18447);
or U23705 (N_23705,N_19310,N_16155);
or U23706 (N_23706,N_15722,N_17514);
nor U23707 (N_23707,N_15670,N_19020);
nor U23708 (N_23708,N_19834,N_16103);
or U23709 (N_23709,N_15638,N_17663);
nand U23710 (N_23710,N_18043,N_19344);
or U23711 (N_23711,N_18092,N_19856);
nand U23712 (N_23712,N_17856,N_17384);
or U23713 (N_23713,N_18677,N_18719);
nor U23714 (N_23714,N_18213,N_19403);
nor U23715 (N_23715,N_18190,N_16291);
and U23716 (N_23716,N_17433,N_17451);
nor U23717 (N_23717,N_16225,N_15808);
or U23718 (N_23718,N_17070,N_15284);
nand U23719 (N_23719,N_16965,N_15507);
nor U23720 (N_23720,N_18511,N_19893);
nand U23721 (N_23721,N_15352,N_19517);
or U23722 (N_23722,N_15598,N_15416);
nand U23723 (N_23723,N_17058,N_15064);
nor U23724 (N_23724,N_16950,N_19900);
nor U23725 (N_23725,N_19571,N_15865);
nand U23726 (N_23726,N_15874,N_18684);
nand U23727 (N_23727,N_19390,N_15885);
or U23728 (N_23728,N_16747,N_18723);
nand U23729 (N_23729,N_18488,N_19150);
nor U23730 (N_23730,N_15458,N_18713);
or U23731 (N_23731,N_15653,N_15288);
or U23732 (N_23732,N_18743,N_16403);
or U23733 (N_23733,N_19700,N_16544);
or U23734 (N_23734,N_15970,N_17206);
and U23735 (N_23735,N_15046,N_17216);
xor U23736 (N_23736,N_16112,N_16529);
and U23737 (N_23737,N_17499,N_19914);
and U23738 (N_23738,N_15797,N_18565);
or U23739 (N_23739,N_18863,N_19032);
and U23740 (N_23740,N_17066,N_16414);
and U23741 (N_23741,N_17923,N_16454);
nand U23742 (N_23742,N_17438,N_19490);
and U23743 (N_23743,N_17773,N_15832);
nor U23744 (N_23744,N_19281,N_16201);
nor U23745 (N_23745,N_16440,N_17714);
and U23746 (N_23746,N_15436,N_15348);
or U23747 (N_23747,N_16630,N_18142);
and U23748 (N_23748,N_19198,N_17726);
nand U23749 (N_23749,N_18376,N_17343);
or U23750 (N_23750,N_17856,N_18228);
nand U23751 (N_23751,N_15200,N_18277);
nor U23752 (N_23752,N_19240,N_16464);
or U23753 (N_23753,N_15163,N_18628);
and U23754 (N_23754,N_18849,N_16133);
or U23755 (N_23755,N_16764,N_16099);
and U23756 (N_23756,N_17531,N_17999);
and U23757 (N_23757,N_15919,N_17122);
and U23758 (N_23758,N_18971,N_17687);
nand U23759 (N_23759,N_18658,N_15814);
nor U23760 (N_23760,N_15015,N_19137);
nor U23761 (N_23761,N_16353,N_15403);
or U23762 (N_23762,N_16158,N_17296);
or U23763 (N_23763,N_18548,N_17962);
or U23764 (N_23764,N_18713,N_17795);
nand U23765 (N_23765,N_18126,N_18079);
nand U23766 (N_23766,N_19051,N_18429);
nor U23767 (N_23767,N_16844,N_18464);
nand U23768 (N_23768,N_18565,N_19074);
nand U23769 (N_23769,N_18400,N_19013);
or U23770 (N_23770,N_15919,N_19738);
or U23771 (N_23771,N_18248,N_18120);
and U23772 (N_23772,N_16423,N_15742);
or U23773 (N_23773,N_19835,N_19748);
xnor U23774 (N_23774,N_17168,N_19552);
nor U23775 (N_23775,N_15731,N_16316);
nor U23776 (N_23776,N_19628,N_18743);
nor U23777 (N_23777,N_18980,N_19170);
nor U23778 (N_23778,N_16607,N_16223);
nand U23779 (N_23779,N_19131,N_17852);
nand U23780 (N_23780,N_15252,N_16834);
nand U23781 (N_23781,N_18684,N_16459);
or U23782 (N_23782,N_18923,N_16487);
nor U23783 (N_23783,N_15550,N_15155);
and U23784 (N_23784,N_19149,N_19962);
xnor U23785 (N_23785,N_19484,N_19198);
and U23786 (N_23786,N_17396,N_17020);
nand U23787 (N_23787,N_18364,N_19657);
nor U23788 (N_23788,N_18527,N_19484);
or U23789 (N_23789,N_18197,N_19762);
nor U23790 (N_23790,N_18020,N_17979);
and U23791 (N_23791,N_16152,N_19092);
or U23792 (N_23792,N_18113,N_19621);
and U23793 (N_23793,N_17468,N_18315);
nor U23794 (N_23794,N_19387,N_15240);
xnor U23795 (N_23795,N_18012,N_16454);
xor U23796 (N_23796,N_19544,N_17501);
or U23797 (N_23797,N_15954,N_19825);
nand U23798 (N_23798,N_17575,N_16130);
nand U23799 (N_23799,N_18830,N_17365);
or U23800 (N_23800,N_15178,N_16564);
xor U23801 (N_23801,N_15515,N_19433);
or U23802 (N_23802,N_16154,N_16731);
nand U23803 (N_23803,N_15423,N_15031);
nand U23804 (N_23804,N_16706,N_18656);
nand U23805 (N_23805,N_18622,N_15609);
or U23806 (N_23806,N_19164,N_18150);
nor U23807 (N_23807,N_15432,N_17160);
and U23808 (N_23808,N_17762,N_19881);
nor U23809 (N_23809,N_18460,N_17995);
nor U23810 (N_23810,N_15420,N_18826);
and U23811 (N_23811,N_17447,N_16550);
and U23812 (N_23812,N_19807,N_19675);
or U23813 (N_23813,N_16046,N_16050);
or U23814 (N_23814,N_18125,N_19600);
nor U23815 (N_23815,N_15277,N_15532);
nor U23816 (N_23816,N_18556,N_17155);
nand U23817 (N_23817,N_15014,N_16846);
or U23818 (N_23818,N_15811,N_16022);
or U23819 (N_23819,N_15687,N_19142);
nor U23820 (N_23820,N_17164,N_16812);
nor U23821 (N_23821,N_17486,N_19135);
nand U23822 (N_23822,N_18060,N_17461);
nor U23823 (N_23823,N_19556,N_19338);
nor U23824 (N_23824,N_16600,N_17101);
nor U23825 (N_23825,N_19406,N_16408);
nor U23826 (N_23826,N_16804,N_15982);
or U23827 (N_23827,N_15214,N_19419);
nor U23828 (N_23828,N_17423,N_19412);
and U23829 (N_23829,N_16350,N_17957);
nand U23830 (N_23830,N_17771,N_16018);
and U23831 (N_23831,N_18463,N_15002);
nand U23832 (N_23832,N_15254,N_17753);
nor U23833 (N_23833,N_15359,N_15368);
nor U23834 (N_23834,N_16215,N_19859);
nand U23835 (N_23835,N_19332,N_18863);
and U23836 (N_23836,N_17715,N_15489);
nor U23837 (N_23837,N_18082,N_18443);
and U23838 (N_23838,N_19285,N_17834);
or U23839 (N_23839,N_18496,N_19320);
or U23840 (N_23840,N_15419,N_17713);
nor U23841 (N_23841,N_19055,N_17930);
nor U23842 (N_23842,N_18348,N_19125);
nor U23843 (N_23843,N_17865,N_16738);
and U23844 (N_23844,N_17300,N_18564);
nand U23845 (N_23845,N_18029,N_15342);
or U23846 (N_23846,N_15966,N_19081);
nor U23847 (N_23847,N_18716,N_18883);
and U23848 (N_23848,N_16021,N_17447);
or U23849 (N_23849,N_18593,N_19722);
and U23850 (N_23850,N_18803,N_15916);
and U23851 (N_23851,N_17911,N_15733);
or U23852 (N_23852,N_15447,N_17747);
xor U23853 (N_23853,N_15873,N_19314);
and U23854 (N_23854,N_17237,N_19569);
nand U23855 (N_23855,N_18246,N_19799);
or U23856 (N_23856,N_15167,N_16281);
nor U23857 (N_23857,N_19948,N_15356);
nand U23858 (N_23858,N_19227,N_15311);
nor U23859 (N_23859,N_17804,N_19389);
or U23860 (N_23860,N_15860,N_18248);
nor U23861 (N_23861,N_15893,N_16942);
and U23862 (N_23862,N_18345,N_18650);
and U23863 (N_23863,N_15269,N_16458);
nand U23864 (N_23864,N_16483,N_19436);
nor U23865 (N_23865,N_19956,N_16443);
and U23866 (N_23866,N_19337,N_17513);
nor U23867 (N_23867,N_18215,N_18350);
and U23868 (N_23868,N_17690,N_16189);
or U23869 (N_23869,N_19734,N_19903);
nand U23870 (N_23870,N_18274,N_16902);
and U23871 (N_23871,N_17268,N_17802);
nor U23872 (N_23872,N_19052,N_16035);
and U23873 (N_23873,N_15128,N_19962);
and U23874 (N_23874,N_17359,N_18756);
nand U23875 (N_23875,N_16511,N_19489);
nand U23876 (N_23876,N_19862,N_18954);
or U23877 (N_23877,N_19370,N_19242);
or U23878 (N_23878,N_19266,N_17966);
nor U23879 (N_23879,N_16927,N_15198);
nor U23880 (N_23880,N_15274,N_17417);
nor U23881 (N_23881,N_16840,N_18240);
nor U23882 (N_23882,N_17431,N_15551);
or U23883 (N_23883,N_17365,N_19461);
nor U23884 (N_23884,N_15772,N_16802);
or U23885 (N_23885,N_15138,N_15903);
nor U23886 (N_23886,N_15175,N_17642);
and U23887 (N_23887,N_19727,N_18987);
and U23888 (N_23888,N_19470,N_15995);
or U23889 (N_23889,N_16153,N_15572);
nand U23890 (N_23890,N_15445,N_15090);
and U23891 (N_23891,N_15649,N_16638);
nor U23892 (N_23892,N_15216,N_16504);
nand U23893 (N_23893,N_19412,N_17760);
and U23894 (N_23894,N_16226,N_18863);
nor U23895 (N_23895,N_18698,N_16093);
or U23896 (N_23896,N_16332,N_15631);
nor U23897 (N_23897,N_19251,N_17936);
and U23898 (N_23898,N_15099,N_15387);
and U23899 (N_23899,N_18003,N_16104);
nand U23900 (N_23900,N_17448,N_16755);
nand U23901 (N_23901,N_15822,N_17934);
or U23902 (N_23902,N_19726,N_18298);
nor U23903 (N_23903,N_19636,N_15870);
or U23904 (N_23904,N_18862,N_18204);
xnor U23905 (N_23905,N_15449,N_15397);
nand U23906 (N_23906,N_17242,N_15802);
and U23907 (N_23907,N_17814,N_15292);
or U23908 (N_23908,N_17120,N_16650);
and U23909 (N_23909,N_16494,N_18364);
and U23910 (N_23910,N_17126,N_16809);
nand U23911 (N_23911,N_17759,N_19886);
nor U23912 (N_23912,N_19263,N_18130);
nand U23913 (N_23913,N_16539,N_15609);
and U23914 (N_23914,N_17563,N_15657);
or U23915 (N_23915,N_19559,N_17840);
or U23916 (N_23916,N_17475,N_17369);
nor U23917 (N_23917,N_16335,N_18959);
or U23918 (N_23918,N_16530,N_15654);
xor U23919 (N_23919,N_17037,N_19083);
nor U23920 (N_23920,N_15624,N_18439);
nor U23921 (N_23921,N_15003,N_15290);
or U23922 (N_23922,N_19204,N_17218);
or U23923 (N_23923,N_18674,N_17252);
xnor U23924 (N_23924,N_17451,N_18944);
nor U23925 (N_23925,N_15118,N_15098);
nand U23926 (N_23926,N_16576,N_19166);
nor U23927 (N_23927,N_16383,N_17953);
and U23928 (N_23928,N_17478,N_19668);
or U23929 (N_23929,N_18651,N_19452);
nor U23930 (N_23930,N_15461,N_15314);
and U23931 (N_23931,N_18281,N_17913);
and U23932 (N_23932,N_16983,N_19929);
or U23933 (N_23933,N_16982,N_16266);
nor U23934 (N_23934,N_17202,N_16565);
and U23935 (N_23935,N_15624,N_19425);
and U23936 (N_23936,N_16428,N_19842);
or U23937 (N_23937,N_18099,N_19398);
and U23938 (N_23938,N_17981,N_19530);
nand U23939 (N_23939,N_17431,N_17112);
nand U23940 (N_23940,N_17320,N_19020);
nand U23941 (N_23941,N_19768,N_16555);
or U23942 (N_23942,N_15933,N_17499);
and U23943 (N_23943,N_16481,N_16133);
or U23944 (N_23944,N_19211,N_18589);
nand U23945 (N_23945,N_15994,N_18855);
nand U23946 (N_23946,N_15818,N_17718);
and U23947 (N_23947,N_17605,N_19195);
or U23948 (N_23948,N_17485,N_19859);
nand U23949 (N_23949,N_15639,N_16383);
nand U23950 (N_23950,N_16730,N_16459);
or U23951 (N_23951,N_17390,N_19332);
and U23952 (N_23952,N_17783,N_17584);
or U23953 (N_23953,N_17008,N_16845);
nor U23954 (N_23954,N_16918,N_17567);
nor U23955 (N_23955,N_19956,N_15484);
or U23956 (N_23956,N_15363,N_15152);
nand U23957 (N_23957,N_19124,N_18618);
nor U23958 (N_23958,N_19466,N_19531);
nand U23959 (N_23959,N_15260,N_19088);
nand U23960 (N_23960,N_16471,N_17075);
and U23961 (N_23961,N_15308,N_18722);
or U23962 (N_23962,N_17715,N_18148);
and U23963 (N_23963,N_17841,N_15228);
or U23964 (N_23964,N_15957,N_19364);
nand U23965 (N_23965,N_16786,N_17111);
nand U23966 (N_23966,N_19791,N_19169);
or U23967 (N_23967,N_17928,N_16913);
nor U23968 (N_23968,N_17626,N_15320);
and U23969 (N_23969,N_16062,N_16852);
or U23970 (N_23970,N_15963,N_15865);
or U23971 (N_23971,N_17981,N_19643);
and U23972 (N_23972,N_18288,N_17284);
or U23973 (N_23973,N_16377,N_18007);
and U23974 (N_23974,N_17014,N_18731);
and U23975 (N_23975,N_15833,N_18229);
nor U23976 (N_23976,N_19286,N_18040);
nand U23977 (N_23977,N_17025,N_18890);
nor U23978 (N_23978,N_16759,N_16256);
and U23979 (N_23979,N_16504,N_19712);
nor U23980 (N_23980,N_17559,N_19208);
nand U23981 (N_23981,N_15852,N_16935);
and U23982 (N_23982,N_17831,N_16879);
nor U23983 (N_23983,N_16925,N_16867);
nand U23984 (N_23984,N_19469,N_16722);
and U23985 (N_23985,N_18029,N_19103);
nand U23986 (N_23986,N_16613,N_19017);
and U23987 (N_23987,N_17076,N_18218);
nor U23988 (N_23988,N_18327,N_17309);
nand U23989 (N_23989,N_19967,N_17154);
or U23990 (N_23990,N_15170,N_19771);
nor U23991 (N_23991,N_19373,N_16842);
nor U23992 (N_23992,N_19269,N_16869);
and U23993 (N_23993,N_19587,N_17388);
nand U23994 (N_23994,N_17265,N_16184);
nand U23995 (N_23995,N_19390,N_19787);
or U23996 (N_23996,N_17365,N_15795);
nor U23997 (N_23997,N_15436,N_15700);
nand U23998 (N_23998,N_19634,N_18097);
nor U23999 (N_23999,N_15006,N_15042);
and U24000 (N_24000,N_16536,N_16068);
nand U24001 (N_24001,N_15700,N_17823);
nand U24002 (N_24002,N_18053,N_16735);
or U24003 (N_24003,N_19555,N_16165);
or U24004 (N_24004,N_19920,N_19862);
nand U24005 (N_24005,N_19494,N_19336);
nand U24006 (N_24006,N_19795,N_19895);
nand U24007 (N_24007,N_17050,N_19215);
or U24008 (N_24008,N_18347,N_17743);
nand U24009 (N_24009,N_19459,N_17837);
nor U24010 (N_24010,N_15777,N_18342);
and U24011 (N_24011,N_18598,N_17056);
and U24012 (N_24012,N_16356,N_18531);
nand U24013 (N_24013,N_18122,N_19847);
xnor U24014 (N_24014,N_19881,N_18036);
nand U24015 (N_24015,N_16928,N_18221);
and U24016 (N_24016,N_18537,N_15576);
and U24017 (N_24017,N_17519,N_15619);
or U24018 (N_24018,N_16969,N_16398);
and U24019 (N_24019,N_17766,N_15226);
nand U24020 (N_24020,N_15588,N_19233);
or U24021 (N_24021,N_16667,N_15714);
nand U24022 (N_24022,N_17198,N_17766);
or U24023 (N_24023,N_19871,N_18394);
nand U24024 (N_24024,N_16655,N_15765);
nand U24025 (N_24025,N_17719,N_18767);
nand U24026 (N_24026,N_18886,N_18943);
or U24027 (N_24027,N_15304,N_19335);
nor U24028 (N_24028,N_19799,N_18736);
and U24029 (N_24029,N_19127,N_16368);
nor U24030 (N_24030,N_18506,N_18322);
or U24031 (N_24031,N_18646,N_19430);
nand U24032 (N_24032,N_15684,N_16650);
nand U24033 (N_24033,N_17508,N_15452);
nor U24034 (N_24034,N_19840,N_17318);
or U24035 (N_24035,N_17932,N_16128);
or U24036 (N_24036,N_15487,N_15997);
nor U24037 (N_24037,N_15795,N_18215);
and U24038 (N_24038,N_18498,N_17658);
nor U24039 (N_24039,N_19149,N_15474);
nand U24040 (N_24040,N_15372,N_15272);
and U24041 (N_24041,N_18854,N_19069);
or U24042 (N_24042,N_15691,N_19489);
nand U24043 (N_24043,N_19851,N_18153);
and U24044 (N_24044,N_19914,N_18927);
or U24045 (N_24045,N_15961,N_16084);
or U24046 (N_24046,N_17572,N_19336);
xor U24047 (N_24047,N_16286,N_15564);
nand U24048 (N_24048,N_18646,N_18851);
nor U24049 (N_24049,N_17866,N_16565);
or U24050 (N_24050,N_16663,N_17855);
or U24051 (N_24051,N_19946,N_15713);
and U24052 (N_24052,N_15126,N_19634);
or U24053 (N_24053,N_17745,N_17398);
nand U24054 (N_24054,N_16504,N_18680);
nor U24055 (N_24055,N_18607,N_15017);
and U24056 (N_24056,N_17473,N_17885);
nand U24057 (N_24057,N_17215,N_19594);
nor U24058 (N_24058,N_15979,N_15528);
nor U24059 (N_24059,N_18543,N_19503);
xor U24060 (N_24060,N_16427,N_15336);
nand U24061 (N_24061,N_17811,N_16538);
nand U24062 (N_24062,N_18523,N_17503);
or U24063 (N_24063,N_15406,N_16852);
or U24064 (N_24064,N_17299,N_15680);
nor U24065 (N_24065,N_17038,N_16172);
nor U24066 (N_24066,N_18073,N_16477);
nand U24067 (N_24067,N_19263,N_18008);
nand U24068 (N_24068,N_16405,N_16447);
nand U24069 (N_24069,N_16223,N_17131);
nor U24070 (N_24070,N_16583,N_15603);
or U24071 (N_24071,N_18063,N_18717);
nand U24072 (N_24072,N_16678,N_19795);
and U24073 (N_24073,N_15090,N_19764);
nand U24074 (N_24074,N_19918,N_15625);
nor U24075 (N_24075,N_15912,N_18432);
or U24076 (N_24076,N_15232,N_19327);
nor U24077 (N_24077,N_19378,N_16840);
or U24078 (N_24078,N_15608,N_15860);
nand U24079 (N_24079,N_16085,N_18608);
and U24080 (N_24080,N_18144,N_15634);
or U24081 (N_24081,N_18982,N_19051);
or U24082 (N_24082,N_19132,N_18658);
nor U24083 (N_24083,N_19837,N_15441);
or U24084 (N_24084,N_15858,N_15960);
xnor U24085 (N_24085,N_16322,N_18008);
nand U24086 (N_24086,N_17022,N_15268);
nor U24087 (N_24087,N_15446,N_17608);
nand U24088 (N_24088,N_16513,N_18848);
nand U24089 (N_24089,N_17183,N_18099);
and U24090 (N_24090,N_18888,N_15998);
or U24091 (N_24091,N_16686,N_18194);
nor U24092 (N_24092,N_15579,N_16577);
or U24093 (N_24093,N_18140,N_18326);
nor U24094 (N_24094,N_18982,N_15063);
nor U24095 (N_24095,N_19895,N_17963);
or U24096 (N_24096,N_17832,N_18984);
or U24097 (N_24097,N_16614,N_17370);
nand U24098 (N_24098,N_15770,N_19087);
nor U24099 (N_24099,N_19681,N_18262);
nand U24100 (N_24100,N_17700,N_16109);
nor U24101 (N_24101,N_16386,N_17706);
or U24102 (N_24102,N_16979,N_19605);
nor U24103 (N_24103,N_16585,N_15919);
nor U24104 (N_24104,N_15422,N_17477);
nand U24105 (N_24105,N_18556,N_19036);
and U24106 (N_24106,N_18172,N_17859);
or U24107 (N_24107,N_18615,N_15127);
or U24108 (N_24108,N_18532,N_17497);
nand U24109 (N_24109,N_15820,N_16852);
or U24110 (N_24110,N_18392,N_16000);
or U24111 (N_24111,N_19691,N_18231);
or U24112 (N_24112,N_15738,N_16149);
and U24113 (N_24113,N_17751,N_16856);
and U24114 (N_24114,N_16014,N_17760);
and U24115 (N_24115,N_16288,N_17091);
nand U24116 (N_24116,N_17700,N_19189);
nand U24117 (N_24117,N_16955,N_18815);
and U24118 (N_24118,N_15529,N_19552);
nand U24119 (N_24119,N_19051,N_15524);
nor U24120 (N_24120,N_16242,N_15668);
nand U24121 (N_24121,N_18236,N_16192);
and U24122 (N_24122,N_15876,N_15756);
nor U24123 (N_24123,N_17574,N_15020);
and U24124 (N_24124,N_18513,N_17659);
nor U24125 (N_24125,N_17270,N_16730);
nand U24126 (N_24126,N_19260,N_19248);
nand U24127 (N_24127,N_19806,N_17720);
or U24128 (N_24128,N_18271,N_15314);
nand U24129 (N_24129,N_17148,N_16828);
nand U24130 (N_24130,N_19659,N_17724);
or U24131 (N_24131,N_17932,N_18462);
and U24132 (N_24132,N_19431,N_16798);
nand U24133 (N_24133,N_15957,N_17371);
or U24134 (N_24134,N_19135,N_17149);
nor U24135 (N_24135,N_15671,N_15624);
or U24136 (N_24136,N_17908,N_15500);
xnor U24137 (N_24137,N_16328,N_15647);
nand U24138 (N_24138,N_16611,N_17856);
nor U24139 (N_24139,N_15620,N_18767);
nor U24140 (N_24140,N_18072,N_16045);
or U24141 (N_24141,N_18555,N_19669);
or U24142 (N_24142,N_16145,N_16560);
nor U24143 (N_24143,N_19819,N_19116);
and U24144 (N_24144,N_18063,N_17556);
or U24145 (N_24145,N_18524,N_18543);
or U24146 (N_24146,N_16150,N_15093);
and U24147 (N_24147,N_18852,N_15051);
or U24148 (N_24148,N_17933,N_18043);
nor U24149 (N_24149,N_19215,N_17893);
nand U24150 (N_24150,N_18808,N_18855);
or U24151 (N_24151,N_19339,N_19794);
nand U24152 (N_24152,N_15059,N_15898);
nand U24153 (N_24153,N_15511,N_17110);
or U24154 (N_24154,N_19230,N_15370);
nand U24155 (N_24155,N_19551,N_16543);
or U24156 (N_24156,N_17967,N_18367);
nand U24157 (N_24157,N_18444,N_17935);
nor U24158 (N_24158,N_15815,N_15025);
or U24159 (N_24159,N_18070,N_16668);
or U24160 (N_24160,N_18925,N_18834);
or U24161 (N_24161,N_19768,N_18850);
and U24162 (N_24162,N_15269,N_15297);
or U24163 (N_24163,N_15721,N_15511);
nor U24164 (N_24164,N_18139,N_15206);
and U24165 (N_24165,N_16215,N_15485);
nor U24166 (N_24166,N_16489,N_18307);
nor U24167 (N_24167,N_17879,N_18359);
or U24168 (N_24168,N_15317,N_19191);
or U24169 (N_24169,N_15081,N_15054);
or U24170 (N_24170,N_17143,N_18050);
or U24171 (N_24171,N_17405,N_16118);
nand U24172 (N_24172,N_17757,N_18759);
nor U24173 (N_24173,N_15967,N_18015);
nand U24174 (N_24174,N_18564,N_17959);
and U24175 (N_24175,N_18916,N_19042);
and U24176 (N_24176,N_16205,N_18303);
and U24177 (N_24177,N_15848,N_19061);
nand U24178 (N_24178,N_15340,N_18840);
nor U24179 (N_24179,N_17243,N_17858);
nor U24180 (N_24180,N_19291,N_18460);
nand U24181 (N_24181,N_19999,N_19308);
xnor U24182 (N_24182,N_16526,N_18569);
and U24183 (N_24183,N_15440,N_16361);
and U24184 (N_24184,N_18526,N_17802);
and U24185 (N_24185,N_19733,N_16050);
xor U24186 (N_24186,N_18216,N_19025);
and U24187 (N_24187,N_19628,N_15176);
nand U24188 (N_24188,N_17143,N_17093);
nand U24189 (N_24189,N_16210,N_15091);
or U24190 (N_24190,N_16347,N_19563);
or U24191 (N_24191,N_15209,N_16219);
and U24192 (N_24192,N_16207,N_16674);
nand U24193 (N_24193,N_18972,N_16614);
nand U24194 (N_24194,N_15673,N_16968);
nor U24195 (N_24195,N_17939,N_17274);
nor U24196 (N_24196,N_16116,N_16214);
and U24197 (N_24197,N_16997,N_18935);
nor U24198 (N_24198,N_18651,N_18777);
or U24199 (N_24199,N_19245,N_17320);
or U24200 (N_24200,N_17551,N_19343);
nand U24201 (N_24201,N_17563,N_15049);
and U24202 (N_24202,N_19550,N_19245);
or U24203 (N_24203,N_15056,N_15746);
xor U24204 (N_24204,N_19799,N_16200);
and U24205 (N_24205,N_15526,N_15689);
nand U24206 (N_24206,N_15827,N_18289);
nand U24207 (N_24207,N_16398,N_15537);
nor U24208 (N_24208,N_18031,N_19914);
and U24209 (N_24209,N_19205,N_16790);
nand U24210 (N_24210,N_19485,N_17142);
nand U24211 (N_24211,N_19122,N_16483);
nand U24212 (N_24212,N_16704,N_18337);
nor U24213 (N_24213,N_19357,N_16966);
or U24214 (N_24214,N_15042,N_15799);
and U24215 (N_24215,N_19983,N_15030);
and U24216 (N_24216,N_16436,N_16965);
and U24217 (N_24217,N_19667,N_16940);
nor U24218 (N_24218,N_18640,N_19711);
nor U24219 (N_24219,N_16787,N_18738);
xor U24220 (N_24220,N_17554,N_15773);
nor U24221 (N_24221,N_19598,N_15779);
or U24222 (N_24222,N_15257,N_16743);
or U24223 (N_24223,N_19925,N_17947);
or U24224 (N_24224,N_15752,N_16522);
nor U24225 (N_24225,N_19713,N_17558);
and U24226 (N_24226,N_18368,N_16045);
nor U24227 (N_24227,N_15152,N_18654);
nand U24228 (N_24228,N_18517,N_16108);
nand U24229 (N_24229,N_19067,N_19691);
or U24230 (N_24230,N_15069,N_18851);
nand U24231 (N_24231,N_19915,N_15884);
and U24232 (N_24232,N_16199,N_19790);
and U24233 (N_24233,N_16408,N_17549);
nand U24234 (N_24234,N_15376,N_17288);
or U24235 (N_24235,N_16449,N_18582);
and U24236 (N_24236,N_17365,N_19264);
nand U24237 (N_24237,N_17462,N_15800);
nand U24238 (N_24238,N_18977,N_16014);
nor U24239 (N_24239,N_17769,N_15048);
and U24240 (N_24240,N_18818,N_16115);
or U24241 (N_24241,N_19165,N_16826);
and U24242 (N_24242,N_17902,N_19639);
nor U24243 (N_24243,N_16603,N_18636);
and U24244 (N_24244,N_17547,N_16191);
or U24245 (N_24245,N_19725,N_19790);
nand U24246 (N_24246,N_15339,N_19955);
nor U24247 (N_24247,N_17248,N_18473);
xnor U24248 (N_24248,N_16362,N_16208);
and U24249 (N_24249,N_18633,N_16539);
and U24250 (N_24250,N_17273,N_16023);
nand U24251 (N_24251,N_17405,N_16452);
or U24252 (N_24252,N_17179,N_15403);
and U24253 (N_24253,N_16555,N_19467);
and U24254 (N_24254,N_19799,N_17784);
nor U24255 (N_24255,N_16489,N_18873);
nor U24256 (N_24256,N_17763,N_17131);
nand U24257 (N_24257,N_15136,N_19877);
and U24258 (N_24258,N_18205,N_16330);
nor U24259 (N_24259,N_15642,N_19185);
or U24260 (N_24260,N_16147,N_15963);
or U24261 (N_24261,N_16721,N_16369);
xor U24262 (N_24262,N_17617,N_18895);
nor U24263 (N_24263,N_19035,N_16171);
nor U24264 (N_24264,N_17479,N_19243);
and U24265 (N_24265,N_19045,N_15161);
nor U24266 (N_24266,N_18200,N_19671);
or U24267 (N_24267,N_16016,N_15816);
or U24268 (N_24268,N_16970,N_16945);
and U24269 (N_24269,N_18809,N_15672);
and U24270 (N_24270,N_18659,N_18456);
nand U24271 (N_24271,N_18939,N_19256);
and U24272 (N_24272,N_19217,N_19675);
or U24273 (N_24273,N_17969,N_16404);
xnor U24274 (N_24274,N_15512,N_17231);
nor U24275 (N_24275,N_18932,N_18055);
nand U24276 (N_24276,N_19596,N_15605);
and U24277 (N_24277,N_18531,N_17820);
nand U24278 (N_24278,N_16362,N_15432);
nor U24279 (N_24279,N_16853,N_16282);
nand U24280 (N_24280,N_19855,N_15400);
nor U24281 (N_24281,N_16521,N_16064);
and U24282 (N_24282,N_19054,N_16493);
nor U24283 (N_24283,N_16691,N_19831);
nand U24284 (N_24284,N_18550,N_17924);
xnor U24285 (N_24285,N_16073,N_19545);
nand U24286 (N_24286,N_19411,N_18529);
nand U24287 (N_24287,N_18447,N_16436);
nor U24288 (N_24288,N_19480,N_19233);
and U24289 (N_24289,N_16852,N_16589);
nor U24290 (N_24290,N_16851,N_19483);
nand U24291 (N_24291,N_17843,N_15084);
or U24292 (N_24292,N_17133,N_17503);
nor U24293 (N_24293,N_17405,N_17307);
or U24294 (N_24294,N_16819,N_17613);
nor U24295 (N_24295,N_16644,N_16631);
nand U24296 (N_24296,N_16441,N_15310);
or U24297 (N_24297,N_16390,N_16987);
and U24298 (N_24298,N_19422,N_18491);
or U24299 (N_24299,N_16613,N_19195);
nand U24300 (N_24300,N_19556,N_16787);
nand U24301 (N_24301,N_16112,N_15270);
or U24302 (N_24302,N_18059,N_18365);
and U24303 (N_24303,N_15631,N_18680);
nor U24304 (N_24304,N_15673,N_17533);
and U24305 (N_24305,N_19662,N_18145);
and U24306 (N_24306,N_18524,N_17291);
or U24307 (N_24307,N_18558,N_18814);
and U24308 (N_24308,N_15825,N_17463);
or U24309 (N_24309,N_16992,N_15614);
nand U24310 (N_24310,N_17601,N_16936);
nand U24311 (N_24311,N_18213,N_16675);
and U24312 (N_24312,N_19634,N_15282);
or U24313 (N_24313,N_17963,N_17116);
nand U24314 (N_24314,N_16279,N_17879);
or U24315 (N_24315,N_19021,N_19273);
nor U24316 (N_24316,N_19767,N_15114);
and U24317 (N_24317,N_17906,N_16844);
nand U24318 (N_24318,N_15596,N_18534);
nand U24319 (N_24319,N_15699,N_19484);
or U24320 (N_24320,N_15760,N_15295);
and U24321 (N_24321,N_18150,N_19046);
nand U24322 (N_24322,N_16241,N_15731);
nor U24323 (N_24323,N_18372,N_16250);
nor U24324 (N_24324,N_15166,N_16194);
nor U24325 (N_24325,N_19622,N_19343);
nor U24326 (N_24326,N_17978,N_16508);
and U24327 (N_24327,N_15748,N_16165);
and U24328 (N_24328,N_17462,N_19278);
nor U24329 (N_24329,N_17227,N_15064);
nand U24330 (N_24330,N_18563,N_19327);
nor U24331 (N_24331,N_19701,N_17545);
or U24332 (N_24332,N_19546,N_17698);
and U24333 (N_24333,N_18058,N_16901);
xnor U24334 (N_24334,N_18325,N_18370);
nor U24335 (N_24335,N_18042,N_17294);
or U24336 (N_24336,N_17074,N_17788);
nor U24337 (N_24337,N_17292,N_16402);
nand U24338 (N_24338,N_19722,N_16474);
and U24339 (N_24339,N_18327,N_16027);
and U24340 (N_24340,N_16226,N_16839);
nor U24341 (N_24341,N_18772,N_18300);
nor U24342 (N_24342,N_17078,N_19801);
nor U24343 (N_24343,N_15209,N_16577);
and U24344 (N_24344,N_18692,N_15070);
nand U24345 (N_24345,N_15930,N_15330);
nor U24346 (N_24346,N_17303,N_15451);
or U24347 (N_24347,N_19924,N_17556);
and U24348 (N_24348,N_16553,N_18345);
or U24349 (N_24349,N_16108,N_19863);
nand U24350 (N_24350,N_16171,N_15132);
and U24351 (N_24351,N_16838,N_18463);
nor U24352 (N_24352,N_16495,N_18722);
or U24353 (N_24353,N_18576,N_17945);
nand U24354 (N_24354,N_18497,N_17897);
nor U24355 (N_24355,N_17394,N_16864);
nand U24356 (N_24356,N_17239,N_18223);
nand U24357 (N_24357,N_19163,N_18041);
nand U24358 (N_24358,N_15904,N_19557);
nor U24359 (N_24359,N_15482,N_15530);
and U24360 (N_24360,N_16907,N_18902);
and U24361 (N_24361,N_15360,N_15957);
or U24362 (N_24362,N_18459,N_17125);
nor U24363 (N_24363,N_17269,N_18589);
and U24364 (N_24364,N_16898,N_19014);
nor U24365 (N_24365,N_18461,N_17072);
nor U24366 (N_24366,N_17314,N_15219);
and U24367 (N_24367,N_15450,N_19991);
nand U24368 (N_24368,N_15861,N_18962);
and U24369 (N_24369,N_17827,N_19651);
or U24370 (N_24370,N_19687,N_17594);
nand U24371 (N_24371,N_18041,N_18247);
and U24372 (N_24372,N_17686,N_19032);
and U24373 (N_24373,N_15137,N_18572);
or U24374 (N_24374,N_17141,N_15892);
nand U24375 (N_24375,N_15820,N_18631);
and U24376 (N_24376,N_15853,N_18342);
nand U24377 (N_24377,N_15141,N_19077);
or U24378 (N_24378,N_18411,N_17405);
nand U24379 (N_24379,N_19528,N_15963);
and U24380 (N_24380,N_15529,N_19828);
or U24381 (N_24381,N_17530,N_17232);
nand U24382 (N_24382,N_17297,N_15805);
and U24383 (N_24383,N_18820,N_18033);
nor U24384 (N_24384,N_17275,N_17987);
nor U24385 (N_24385,N_15852,N_19704);
nor U24386 (N_24386,N_15036,N_18777);
nor U24387 (N_24387,N_15784,N_17123);
or U24388 (N_24388,N_16114,N_15353);
or U24389 (N_24389,N_16366,N_17255);
and U24390 (N_24390,N_18809,N_15952);
nand U24391 (N_24391,N_16413,N_16700);
nand U24392 (N_24392,N_19396,N_17524);
and U24393 (N_24393,N_15214,N_15144);
nand U24394 (N_24394,N_18681,N_18620);
or U24395 (N_24395,N_19210,N_17092);
and U24396 (N_24396,N_16499,N_17401);
or U24397 (N_24397,N_15348,N_18173);
xor U24398 (N_24398,N_16799,N_19831);
nand U24399 (N_24399,N_15115,N_15087);
nor U24400 (N_24400,N_16322,N_18995);
nand U24401 (N_24401,N_18144,N_19632);
nor U24402 (N_24402,N_19423,N_18892);
and U24403 (N_24403,N_19917,N_19190);
nand U24404 (N_24404,N_15432,N_16112);
nand U24405 (N_24405,N_16452,N_18693);
or U24406 (N_24406,N_17948,N_15382);
nand U24407 (N_24407,N_16207,N_15133);
and U24408 (N_24408,N_15751,N_15312);
and U24409 (N_24409,N_17454,N_19391);
nor U24410 (N_24410,N_18451,N_19872);
and U24411 (N_24411,N_16853,N_18545);
and U24412 (N_24412,N_15908,N_16922);
and U24413 (N_24413,N_18814,N_17193);
nor U24414 (N_24414,N_16944,N_18162);
nor U24415 (N_24415,N_15426,N_19107);
or U24416 (N_24416,N_16922,N_15961);
and U24417 (N_24417,N_17812,N_16183);
nand U24418 (N_24418,N_18275,N_19617);
nor U24419 (N_24419,N_17750,N_15781);
nor U24420 (N_24420,N_15191,N_15820);
nand U24421 (N_24421,N_16276,N_16877);
nor U24422 (N_24422,N_18024,N_16752);
nand U24423 (N_24423,N_19523,N_15380);
and U24424 (N_24424,N_19445,N_17952);
and U24425 (N_24425,N_17499,N_18292);
and U24426 (N_24426,N_17452,N_17213);
and U24427 (N_24427,N_16396,N_16893);
nor U24428 (N_24428,N_15646,N_17177);
nor U24429 (N_24429,N_18411,N_18767);
and U24430 (N_24430,N_15292,N_16486);
nor U24431 (N_24431,N_15900,N_15673);
and U24432 (N_24432,N_15912,N_16305);
nand U24433 (N_24433,N_15061,N_18404);
nor U24434 (N_24434,N_16622,N_18409);
or U24435 (N_24435,N_18890,N_18804);
or U24436 (N_24436,N_15792,N_19936);
nand U24437 (N_24437,N_15821,N_15716);
nor U24438 (N_24438,N_16160,N_17450);
and U24439 (N_24439,N_17701,N_19945);
nor U24440 (N_24440,N_17182,N_17873);
nand U24441 (N_24441,N_17664,N_19718);
or U24442 (N_24442,N_16379,N_15179);
nor U24443 (N_24443,N_15003,N_15014);
nand U24444 (N_24444,N_17217,N_19320);
nand U24445 (N_24445,N_16689,N_18389);
and U24446 (N_24446,N_16277,N_19505);
nor U24447 (N_24447,N_16834,N_19913);
and U24448 (N_24448,N_19941,N_16206);
nand U24449 (N_24449,N_19303,N_16549);
and U24450 (N_24450,N_16096,N_16037);
nor U24451 (N_24451,N_16827,N_17229);
nand U24452 (N_24452,N_19715,N_15100);
nor U24453 (N_24453,N_19793,N_19810);
nor U24454 (N_24454,N_15440,N_18929);
nor U24455 (N_24455,N_15105,N_19734);
and U24456 (N_24456,N_15436,N_16419);
and U24457 (N_24457,N_15416,N_18159);
nand U24458 (N_24458,N_16319,N_19733);
or U24459 (N_24459,N_18777,N_15827);
and U24460 (N_24460,N_19388,N_16060);
and U24461 (N_24461,N_15296,N_15053);
or U24462 (N_24462,N_18601,N_18144);
nor U24463 (N_24463,N_15645,N_15649);
nand U24464 (N_24464,N_15257,N_19955);
nor U24465 (N_24465,N_15227,N_17315);
xor U24466 (N_24466,N_15289,N_15489);
and U24467 (N_24467,N_16177,N_19498);
or U24468 (N_24468,N_19909,N_15476);
or U24469 (N_24469,N_16529,N_18345);
nand U24470 (N_24470,N_16735,N_18812);
or U24471 (N_24471,N_15725,N_17911);
and U24472 (N_24472,N_16512,N_17916);
nor U24473 (N_24473,N_18296,N_16890);
or U24474 (N_24474,N_19168,N_19604);
and U24475 (N_24475,N_17174,N_18252);
or U24476 (N_24476,N_17605,N_15752);
and U24477 (N_24477,N_18132,N_19958);
nor U24478 (N_24478,N_19548,N_17459);
nor U24479 (N_24479,N_15729,N_16487);
or U24480 (N_24480,N_18575,N_15763);
nor U24481 (N_24481,N_17564,N_17900);
or U24482 (N_24482,N_19141,N_15704);
nand U24483 (N_24483,N_16704,N_17125);
and U24484 (N_24484,N_17585,N_15722);
nand U24485 (N_24485,N_15306,N_15330);
and U24486 (N_24486,N_18804,N_16394);
or U24487 (N_24487,N_16752,N_17191);
and U24488 (N_24488,N_16818,N_17857);
and U24489 (N_24489,N_17483,N_16607);
and U24490 (N_24490,N_16981,N_17199);
nand U24491 (N_24491,N_16578,N_16153);
or U24492 (N_24492,N_15816,N_17076);
nand U24493 (N_24493,N_19324,N_18465);
nor U24494 (N_24494,N_16990,N_17821);
or U24495 (N_24495,N_19895,N_17509);
nand U24496 (N_24496,N_15937,N_18872);
or U24497 (N_24497,N_19363,N_15339);
or U24498 (N_24498,N_19458,N_17580);
or U24499 (N_24499,N_16110,N_15883);
nand U24500 (N_24500,N_16838,N_18786);
or U24501 (N_24501,N_17113,N_16980);
nor U24502 (N_24502,N_15837,N_15262);
and U24503 (N_24503,N_18242,N_19334);
and U24504 (N_24504,N_16062,N_18400);
nand U24505 (N_24505,N_19569,N_15052);
nor U24506 (N_24506,N_15679,N_15512);
xor U24507 (N_24507,N_15913,N_19019);
or U24508 (N_24508,N_18682,N_17433);
and U24509 (N_24509,N_17523,N_15859);
nor U24510 (N_24510,N_16052,N_15658);
nand U24511 (N_24511,N_19938,N_15877);
or U24512 (N_24512,N_15193,N_19526);
nor U24513 (N_24513,N_18676,N_19621);
nand U24514 (N_24514,N_16317,N_19480);
or U24515 (N_24515,N_19256,N_17335);
or U24516 (N_24516,N_16723,N_15424);
nand U24517 (N_24517,N_15992,N_17452);
and U24518 (N_24518,N_19098,N_15872);
nand U24519 (N_24519,N_18836,N_19893);
and U24520 (N_24520,N_17298,N_19008);
nor U24521 (N_24521,N_19668,N_16580);
or U24522 (N_24522,N_19366,N_17088);
or U24523 (N_24523,N_19332,N_17076);
nor U24524 (N_24524,N_17523,N_17921);
and U24525 (N_24525,N_18896,N_16056);
or U24526 (N_24526,N_17278,N_17336);
nor U24527 (N_24527,N_19958,N_16697);
nand U24528 (N_24528,N_19324,N_17061);
and U24529 (N_24529,N_15342,N_16481);
and U24530 (N_24530,N_16189,N_16316);
nand U24531 (N_24531,N_15382,N_16792);
and U24532 (N_24532,N_17266,N_18945);
or U24533 (N_24533,N_17445,N_18992);
xor U24534 (N_24534,N_17627,N_16423);
xor U24535 (N_24535,N_19062,N_16310);
nor U24536 (N_24536,N_17292,N_16270);
nor U24537 (N_24537,N_17531,N_19647);
or U24538 (N_24538,N_18672,N_19426);
or U24539 (N_24539,N_15262,N_18316);
and U24540 (N_24540,N_18077,N_18226);
and U24541 (N_24541,N_19887,N_17958);
and U24542 (N_24542,N_16574,N_18210);
or U24543 (N_24543,N_19441,N_18118);
nor U24544 (N_24544,N_18477,N_18179);
or U24545 (N_24545,N_17654,N_17507);
nand U24546 (N_24546,N_17371,N_18162);
and U24547 (N_24547,N_18732,N_18813);
or U24548 (N_24548,N_17766,N_15078);
or U24549 (N_24549,N_19971,N_19216);
nand U24550 (N_24550,N_17402,N_17389);
xnor U24551 (N_24551,N_17211,N_16076);
nand U24552 (N_24552,N_18209,N_17124);
and U24553 (N_24553,N_18684,N_16654);
nor U24554 (N_24554,N_18828,N_16731);
nor U24555 (N_24555,N_15423,N_18806);
nor U24556 (N_24556,N_17514,N_16470);
or U24557 (N_24557,N_18076,N_16262);
or U24558 (N_24558,N_15370,N_18586);
and U24559 (N_24559,N_18770,N_15142);
nor U24560 (N_24560,N_18533,N_16767);
or U24561 (N_24561,N_16952,N_15200);
nor U24562 (N_24562,N_18656,N_17774);
nand U24563 (N_24563,N_17435,N_17758);
or U24564 (N_24564,N_16851,N_19547);
and U24565 (N_24565,N_19396,N_18214);
nand U24566 (N_24566,N_16075,N_18483);
or U24567 (N_24567,N_17872,N_15297);
nand U24568 (N_24568,N_19023,N_16112);
nor U24569 (N_24569,N_16566,N_19632);
or U24570 (N_24570,N_19663,N_17207);
and U24571 (N_24571,N_18555,N_17012);
nand U24572 (N_24572,N_17313,N_15809);
nand U24573 (N_24573,N_15855,N_17575);
or U24574 (N_24574,N_18045,N_16222);
nand U24575 (N_24575,N_18117,N_15669);
nor U24576 (N_24576,N_17615,N_18939);
and U24577 (N_24577,N_17631,N_17639);
and U24578 (N_24578,N_15671,N_16388);
nand U24579 (N_24579,N_17287,N_17055);
or U24580 (N_24580,N_18158,N_15239);
nand U24581 (N_24581,N_16042,N_16778);
nor U24582 (N_24582,N_15861,N_18632);
or U24583 (N_24583,N_17412,N_19632);
nor U24584 (N_24584,N_17917,N_18870);
or U24585 (N_24585,N_18391,N_17809);
nor U24586 (N_24586,N_17458,N_19873);
nor U24587 (N_24587,N_16528,N_16659);
or U24588 (N_24588,N_17460,N_18647);
or U24589 (N_24589,N_16892,N_19301);
nor U24590 (N_24590,N_19575,N_15585);
nand U24591 (N_24591,N_16423,N_19811);
nand U24592 (N_24592,N_15422,N_17533);
nand U24593 (N_24593,N_17254,N_16865);
nand U24594 (N_24594,N_19095,N_19407);
or U24595 (N_24595,N_16822,N_16257);
nand U24596 (N_24596,N_15140,N_16135);
xnor U24597 (N_24597,N_16317,N_16714);
or U24598 (N_24598,N_19500,N_17356);
nor U24599 (N_24599,N_16764,N_18049);
nand U24600 (N_24600,N_16717,N_15253);
nand U24601 (N_24601,N_16234,N_15805);
and U24602 (N_24602,N_16340,N_15222);
or U24603 (N_24603,N_16699,N_16589);
nor U24604 (N_24604,N_15839,N_19164);
xor U24605 (N_24605,N_15182,N_16954);
and U24606 (N_24606,N_17627,N_16400);
xor U24607 (N_24607,N_15005,N_15984);
or U24608 (N_24608,N_15026,N_16824);
or U24609 (N_24609,N_17846,N_15079);
and U24610 (N_24610,N_17557,N_18809);
and U24611 (N_24611,N_18970,N_18386);
nor U24612 (N_24612,N_15834,N_17313);
nand U24613 (N_24613,N_18598,N_17560);
nor U24614 (N_24614,N_16908,N_16038);
nor U24615 (N_24615,N_16203,N_16003);
and U24616 (N_24616,N_18192,N_15083);
or U24617 (N_24617,N_17445,N_16351);
or U24618 (N_24618,N_17822,N_19010);
or U24619 (N_24619,N_17035,N_19566);
and U24620 (N_24620,N_16123,N_15029);
or U24621 (N_24621,N_19638,N_16175);
nand U24622 (N_24622,N_16551,N_18194);
and U24623 (N_24623,N_18525,N_15830);
xnor U24624 (N_24624,N_18079,N_15878);
or U24625 (N_24625,N_16788,N_16238);
and U24626 (N_24626,N_19426,N_17432);
nor U24627 (N_24627,N_19544,N_17770);
and U24628 (N_24628,N_15736,N_16637);
and U24629 (N_24629,N_18833,N_18098);
or U24630 (N_24630,N_17704,N_15840);
or U24631 (N_24631,N_17226,N_16291);
or U24632 (N_24632,N_17598,N_17939);
nand U24633 (N_24633,N_19980,N_19337);
nand U24634 (N_24634,N_15939,N_15158);
xor U24635 (N_24635,N_16328,N_16497);
or U24636 (N_24636,N_16429,N_19757);
or U24637 (N_24637,N_18544,N_19457);
and U24638 (N_24638,N_18725,N_18312);
nand U24639 (N_24639,N_17186,N_15854);
nand U24640 (N_24640,N_15076,N_19854);
nand U24641 (N_24641,N_17950,N_18191);
nand U24642 (N_24642,N_17443,N_16571);
nor U24643 (N_24643,N_15945,N_18026);
nand U24644 (N_24644,N_16143,N_18788);
or U24645 (N_24645,N_17280,N_19344);
nand U24646 (N_24646,N_18688,N_18693);
xor U24647 (N_24647,N_17241,N_18921);
and U24648 (N_24648,N_15920,N_16109);
and U24649 (N_24649,N_19365,N_15849);
nor U24650 (N_24650,N_19807,N_18703);
nand U24651 (N_24651,N_16345,N_16424);
nor U24652 (N_24652,N_15790,N_15644);
nand U24653 (N_24653,N_16038,N_19315);
or U24654 (N_24654,N_19756,N_16347);
nor U24655 (N_24655,N_18516,N_19460);
nand U24656 (N_24656,N_16355,N_16531);
nand U24657 (N_24657,N_19551,N_16114);
or U24658 (N_24658,N_19800,N_15886);
nand U24659 (N_24659,N_17791,N_19599);
nor U24660 (N_24660,N_17836,N_18198);
nor U24661 (N_24661,N_18801,N_15681);
nor U24662 (N_24662,N_16062,N_15614);
or U24663 (N_24663,N_18249,N_17272);
and U24664 (N_24664,N_16545,N_17583);
and U24665 (N_24665,N_16209,N_15317);
nor U24666 (N_24666,N_17737,N_16168);
or U24667 (N_24667,N_15063,N_15218);
and U24668 (N_24668,N_18063,N_16287);
and U24669 (N_24669,N_16059,N_19239);
nand U24670 (N_24670,N_18295,N_17017);
or U24671 (N_24671,N_16456,N_18983);
or U24672 (N_24672,N_16989,N_17256);
nor U24673 (N_24673,N_19637,N_15784);
or U24674 (N_24674,N_16308,N_15948);
or U24675 (N_24675,N_15851,N_18320);
nor U24676 (N_24676,N_18087,N_17914);
and U24677 (N_24677,N_19119,N_18726);
or U24678 (N_24678,N_18816,N_18377);
nor U24679 (N_24679,N_16919,N_17579);
or U24680 (N_24680,N_17077,N_18746);
or U24681 (N_24681,N_19745,N_15203);
or U24682 (N_24682,N_15633,N_17323);
and U24683 (N_24683,N_17850,N_18931);
xnor U24684 (N_24684,N_15005,N_18351);
nand U24685 (N_24685,N_15736,N_15808);
nand U24686 (N_24686,N_19260,N_18110);
or U24687 (N_24687,N_15918,N_15354);
or U24688 (N_24688,N_19883,N_17883);
and U24689 (N_24689,N_17954,N_19140);
and U24690 (N_24690,N_15705,N_19868);
or U24691 (N_24691,N_18889,N_18723);
or U24692 (N_24692,N_16129,N_16662);
nor U24693 (N_24693,N_16098,N_15122);
nor U24694 (N_24694,N_19333,N_18488);
nand U24695 (N_24695,N_16359,N_19435);
or U24696 (N_24696,N_19778,N_16214);
and U24697 (N_24697,N_19452,N_16243);
nor U24698 (N_24698,N_18768,N_15567);
and U24699 (N_24699,N_15360,N_17265);
or U24700 (N_24700,N_15232,N_16756);
nand U24701 (N_24701,N_19889,N_19984);
and U24702 (N_24702,N_16210,N_15689);
nor U24703 (N_24703,N_15938,N_15247);
and U24704 (N_24704,N_18715,N_16669);
nor U24705 (N_24705,N_19661,N_17264);
nor U24706 (N_24706,N_16951,N_16711);
nand U24707 (N_24707,N_18274,N_19605);
nor U24708 (N_24708,N_15153,N_17256);
nand U24709 (N_24709,N_15853,N_15867);
nor U24710 (N_24710,N_19146,N_19002);
and U24711 (N_24711,N_19185,N_18467);
and U24712 (N_24712,N_17247,N_18030);
or U24713 (N_24713,N_18351,N_18072);
or U24714 (N_24714,N_17786,N_16576);
nand U24715 (N_24715,N_19669,N_15318);
nand U24716 (N_24716,N_19428,N_17982);
and U24717 (N_24717,N_17431,N_19874);
and U24718 (N_24718,N_15048,N_16356);
nor U24719 (N_24719,N_16063,N_16403);
or U24720 (N_24720,N_15634,N_17318);
or U24721 (N_24721,N_16962,N_19734);
or U24722 (N_24722,N_18201,N_18740);
nand U24723 (N_24723,N_17350,N_15291);
or U24724 (N_24724,N_15696,N_17242);
or U24725 (N_24725,N_18262,N_17596);
nand U24726 (N_24726,N_18339,N_19672);
nand U24727 (N_24727,N_18642,N_19298);
or U24728 (N_24728,N_17300,N_19118);
nor U24729 (N_24729,N_19759,N_17460);
nand U24730 (N_24730,N_16295,N_17777);
and U24731 (N_24731,N_18835,N_19416);
nor U24732 (N_24732,N_18571,N_17329);
nor U24733 (N_24733,N_18210,N_16777);
xor U24734 (N_24734,N_15684,N_16082);
or U24735 (N_24735,N_15559,N_17181);
nor U24736 (N_24736,N_17167,N_17756);
nand U24737 (N_24737,N_19384,N_19889);
or U24738 (N_24738,N_15114,N_18710);
or U24739 (N_24739,N_15054,N_18619);
and U24740 (N_24740,N_18400,N_16601);
nand U24741 (N_24741,N_16429,N_16990);
or U24742 (N_24742,N_18012,N_19666);
nand U24743 (N_24743,N_16240,N_16780);
or U24744 (N_24744,N_17953,N_19274);
and U24745 (N_24745,N_15763,N_18305);
nand U24746 (N_24746,N_17556,N_16637);
and U24747 (N_24747,N_19377,N_17970);
or U24748 (N_24748,N_15159,N_19256);
and U24749 (N_24749,N_18864,N_18725);
nand U24750 (N_24750,N_16756,N_19922);
and U24751 (N_24751,N_15475,N_19388);
nor U24752 (N_24752,N_16742,N_16338);
and U24753 (N_24753,N_18346,N_19797);
nand U24754 (N_24754,N_15424,N_15638);
xnor U24755 (N_24755,N_17484,N_16651);
or U24756 (N_24756,N_19607,N_16031);
or U24757 (N_24757,N_19270,N_15986);
nand U24758 (N_24758,N_18405,N_18001);
and U24759 (N_24759,N_15485,N_19349);
nand U24760 (N_24760,N_18674,N_19587);
or U24761 (N_24761,N_18280,N_19901);
or U24762 (N_24762,N_18232,N_18246);
and U24763 (N_24763,N_19177,N_17060);
and U24764 (N_24764,N_19709,N_15683);
or U24765 (N_24765,N_15215,N_18777);
and U24766 (N_24766,N_18020,N_17496);
and U24767 (N_24767,N_15197,N_16105);
and U24768 (N_24768,N_18444,N_18435);
and U24769 (N_24769,N_17505,N_19465);
nor U24770 (N_24770,N_18615,N_15510);
and U24771 (N_24771,N_18939,N_17806);
nor U24772 (N_24772,N_16621,N_15243);
nand U24773 (N_24773,N_17111,N_19533);
nor U24774 (N_24774,N_17117,N_19042);
nand U24775 (N_24775,N_17434,N_15413);
or U24776 (N_24776,N_19014,N_19280);
or U24777 (N_24777,N_19399,N_16632);
and U24778 (N_24778,N_18652,N_19559);
or U24779 (N_24779,N_18433,N_19261);
and U24780 (N_24780,N_16964,N_17953);
and U24781 (N_24781,N_19186,N_19605);
or U24782 (N_24782,N_19276,N_17152);
or U24783 (N_24783,N_15685,N_18077);
nand U24784 (N_24784,N_18095,N_16758);
nand U24785 (N_24785,N_17449,N_18237);
nand U24786 (N_24786,N_16659,N_19994);
or U24787 (N_24787,N_15105,N_15690);
nor U24788 (N_24788,N_16511,N_17923);
nand U24789 (N_24789,N_19571,N_18577);
nor U24790 (N_24790,N_15464,N_18927);
nand U24791 (N_24791,N_18616,N_15680);
nor U24792 (N_24792,N_17785,N_17677);
nor U24793 (N_24793,N_15578,N_18516);
or U24794 (N_24794,N_18408,N_18052);
nor U24795 (N_24795,N_16789,N_18790);
and U24796 (N_24796,N_18927,N_16504);
nand U24797 (N_24797,N_17996,N_16847);
nand U24798 (N_24798,N_19684,N_15377);
and U24799 (N_24799,N_19382,N_19210);
or U24800 (N_24800,N_18591,N_16677);
nand U24801 (N_24801,N_15149,N_16798);
nor U24802 (N_24802,N_16974,N_16087);
xor U24803 (N_24803,N_16469,N_15282);
or U24804 (N_24804,N_15214,N_17480);
or U24805 (N_24805,N_17423,N_17928);
or U24806 (N_24806,N_18980,N_19120);
nand U24807 (N_24807,N_15718,N_15608);
nor U24808 (N_24808,N_16592,N_19649);
xnor U24809 (N_24809,N_17580,N_16288);
and U24810 (N_24810,N_15684,N_16375);
nor U24811 (N_24811,N_18012,N_18017);
xnor U24812 (N_24812,N_19189,N_17806);
and U24813 (N_24813,N_18378,N_15144);
and U24814 (N_24814,N_16742,N_16083);
or U24815 (N_24815,N_19800,N_16494);
or U24816 (N_24816,N_19920,N_19118);
or U24817 (N_24817,N_18076,N_19115);
nor U24818 (N_24818,N_18578,N_19832);
nor U24819 (N_24819,N_15235,N_16472);
or U24820 (N_24820,N_19678,N_18515);
and U24821 (N_24821,N_18082,N_17507);
or U24822 (N_24822,N_17991,N_15211);
or U24823 (N_24823,N_19406,N_17033);
or U24824 (N_24824,N_15241,N_17255);
nor U24825 (N_24825,N_18585,N_16888);
and U24826 (N_24826,N_17166,N_15120);
nor U24827 (N_24827,N_18343,N_18922);
nor U24828 (N_24828,N_19057,N_19164);
nor U24829 (N_24829,N_19564,N_16636);
and U24830 (N_24830,N_18131,N_15932);
or U24831 (N_24831,N_16739,N_19487);
and U24832 (N_24832,N_15581,N_15818);
nand U24833 (N_24833,N_19440,N_16235);
xor U24834 (N_24834,N_17127,N_18810);
nand U24835 (N_24835,N_19510,N_15782);
and U24836 (N_24836,N_15173,N_19889);
nand U24837 (N_24837,N_15998,N_19219);
nor U24838 (N_24838,N_15909,N_16371);
and U24839 (N_24839,N_19653,N_19517);
and U24840 (N_24840,N_17284,N_15023);
or U24841 (N_24841,N_16729,N_18141);
nor U24842 (N_24842,N_18185,N_16134);
or U24843 (N_24843,N_19104,N_19269);
nand U24844 (N_24844,N_18846,N_18250);
nand U24845 (N_24845,N_19104,N_16806);
and U24846 (N_24846,N_17752,N_19094);
nor U24847 (N_24847,N_18034,N_18435);
nand U24848 (N_24848,N_17144,N_16147);
and U24849 (N_24849,N_17469,N_19553);
or U24850 (N_24850,N_17935,N_15371);
nand U24851 (N_24851,N_19828,N_18645);
and U24852 (N_24852,N_15158,N_19223);
and U24853 (N_24853,N_16295,N_18254);
or U24854 (N_24854,N_17477,N_17097);
or U24855 (N_24855,N_16197,N_18806);
or U24856 (N_24856,N_15412,N_19982);
and U24857 (N_24857,N_16659,N_18887);
or U24858 (N_24858,N_16224,N_15639);
nand U24859 (N_24859,N_15388,N_18652);
nand U24860 (N_24860,N_16954,N_16339);
and U24861 (N_24861,N_17207,N_17603);
nor U24862 (N_24862,N_17871,N_17538);
nand U24863 (N_24863,N_15489,N_18262);
or U24864 (N_24864,N_17944,N_16920);
xnor U24865 (N_24865,N_17497,N_16987);
nand U24866 (N_24866,N_15747,N_15764);
nor U24867 (N_24867,N_19722,N_18857);
nand U24868 (N_24868,N_16102,N_18646);
nand U24869 (N_24869,N_19055,N_16768);
nand U24870 (N_24870,N_17553,N_19169);
or U24871 (N_24871,N_19700,N_18590);
nand U24872 (N_24872,N_18267,N_18885);
nor U24873 (N_24873,N_18859,N_18424);
and U24874 (N_24874,N_19029,N_16807);
and U24875 (N_24875,N_19653,N_18729);
and U24876 (N_24876,N_16687,N_19125);
or U24877 (N_24877,N_17443,N_18885);
nand U24878 (N_24878,N_16237,N_19265);
nor U24879 (N_24879,N_18053,N_17698);
and U24880 (N_24880,N_19743,N_16001);
or U24881 (N_24881,N_15781,N_18195);
nor U24882 (N_24882,N_17804,N_19137);
or U24883 (N_24883,N_18516,N_16580);
nand U24884 (N_24884,N_19734,N_18284);
or U24885 (N_24885,N_19459,N_15630);
nor U24886 (N_24886,N_19263,N_19427);
and U24887 (N_24887,N_15378,N_17474);
nand U24888 (N_24888,N_18835,N_15321);
nor U24889 (N_24889,N_17327,N_16299);
nand U24890 (N_24890,N_19331,N_19538);
nand U24891 (N_24891,N_18196,N_19840);
or U24892 (N_24892,N_19693,N_19102);
nand U24893 (N_24893,N_19062,N_17813);
or U24894 (N_24894,N_15457,N_19805);
nor U24895 (N_24895,N_18938,N_15809);
nor U24896 (N_24896,N_16444,N_16953);
or U24897 (N_24897,N_17768,N_17224);
nor U24898 (N_24898,N_16169,N_15915);
nand U24899 (N_24899,N_19334,N_16697);
xor U24900 (N_24900,N_18997,N_18076);
nand U24901 (N_24901,N_15153,N_16311);
and U24902 (N_24902,N_18276,N_17158);
and U24903 (N_24903,N_16295,N_17445);
and U24904 (N_24904,N_19079,N_15117);
nor U24905 (N_24905,N_19721,N_19212);
nand U24906 (N_24906,N_15840,N_17847);
or U24907 (N_24907,N_16489,N_19055);
nor U24908 (N_24908,N_15996,N_18968);
and U24909 (N_24909,N_15759,N_17829);
nor U24910 (N_24910,N_18488,N_16165);
nor U24911 (N_24911,N_15540,N_17932);
nor U24912 (N_24912,N_19782,N_16327);
or U24913 (N_24913,N_19928,N_16480);
or U24914 (N_24914,N_15047,N_19984);
nor U24915 (N_24915,N_18903,N_18114);
nor U24916 (N_24916,N_17593,N_17042);
nor U24917 (N_24917,N_18684,N_16673);
or U24918 (N_24918,N_15928,N_19252);
nor U24919 (N_24919,N_17036,N_18539);
or U24920 (N_24920,N_19929,N_15657);
nor U24921 (N_24921,N_15998,N_19264);
nor U24922 (N_24922,N_15751,N_18047);
nand U24923 (N_24923,N_18520,N_19219);
nand U24924 (N_24924,N_16076,N_17105);
nor U24925 (N_24925,N_18089,N_17373);
nor U24926 (N_24926,N_18492,N_17724);
nand U24927 (N_24927,N_18091,N_15457);
nor U24928 (N_24928,N_15543,N_17169);
nor U24929 (N_24929,N_19914,N_16566);
nor U24930 (N_24930,N_18827,N_15017);
and U24931 (N_24931,N_15226,N_15747);
and U24932 (N_24932,N_16808,N_18725);
or U24933 (N_24933,N_17002,N_19593);
nand U24934 (N_24934,N_17764,N_16218);
or U24935 (N_24935,N_15041,N_19190);
nand U24936 (N_24936,N_16878,N_17508);
or U24937 (N_24937,N_18505,N_17613);
nand U24938 (N_24938,N_19366,N_17966);
nor U24939 (N_24939,N_17538,N_15916);
and U24940 (N_24940,N_19106,N_17455);
or U24941 (N_24941,N_16387,N_15143);
or U24942 (N_24942,N_15362,N_15518);
or U24943 (N_24943,N_19305,N_17027);
and U24944 (N_24944,N_18091,N_16432);
or U24945 (N_24945,N_15495,N_18417);
and U24946 (N_24946,N_17129,N_18384);
and U24947 (N_24947,N_19600,N_17474);
or U24948 (N_24948,N_18469,N_15868);
and U24949 (N_24949,N_18132,N_17942);
nor U24950 (N_24950,N_19875,N_17535);
or U24951 (N_24951,N_19831,N_16525);
nand U24952 (N_24952,N_16813,N_16468);
or U24953 (N_24953,N_15598,N_18203);
nand U24954 (N_24954,N_17868,N_15552);
nor U24955 (N_24955,N_18246,N_15959);
or U24956 (N_24956,N_18429,N_16996);
nand U24957 (N_24957,N_17846,N_16846);
and U24958 (N_24958,N_18609,N_18586);
or U24959 (N_24959,N_16290,N_17089);
or U24960 (N_24960,N_18909,N_16538);
or U24961 (N_24961,N_18057,N_15375);
nor U24962 (N_24962,N_15076,N_15479);
or U24963 (N_24963,N_15109,N_18283);
and U24964 (N_24964,N_17395,N_16500);
or U24965 (N_24965,N_17424,N_16328);
nor U24966 (N_24966,N_16317,N_19608);
nor U24967 (N_24967,N_15716,N_17775);
or U24968 (N_24968,N_15239,N_16717);
nor U24969 (N_24969,N_16809,N_19991);
nor U24970 (N_24970,N_15744,N_17427);
or U24971 (N_24971,N_17252,N_15690);
and U24972 (N_24972,N_17235,N_16570);
or U24973 (N_24973,N_15313,N_16033);
nand U24974 (N_24974,N_15167,N_17710);
nand U24975 (N_24975,N_15651,N_16016);
or U24976 (N_24976,N_17562,N_15920);
or U24977 (N_24977,N_15479,N_17978);
and U24978 (N_24978,N_16082,N_19785);
nand U24979 (N_24979,N_17103,N_17034);
nor U24980 (N_24980,N_17915,N_16969);
nor U24981 (N_24981,N_17248,N_15057);
and U24982 (N_24982,N_18231,N_16901);
and U24983 (N_24983,N_16894,N_17455);
nor U24984 (N_24984,N_15689,N_17034);
nand U24985 (N_24985,N_18157,N_16346);
nor U24986 (N_24986,N_18542,N_16755);
nand U24987 (N_24987,N_18977,N_17675);
nor U24988 (N_24988,N_19449,N_18349);
and U24989 (N_24989,N_15815,N_16747);
nand U24990 (N_24990,N_18944,N_18015);
nor U24991 (N_24991,N_16996,N_18976);
or U24992 (N_24992,N_17091,N_19708);
nand U24993 (N_24993,N_16560,N_16594);
or U24994 (N_24994,N_16833,N_17173);
nand U24995 (N_24995,N_15060,N_19891);
nor U24996 (N_24996,N_19522,N_18867);
nand U24997 (N_24997,N_17904,N_16732);
and U24998 (N_24998,N_19637,N_16272);
nor U24999 (N_24999,N_19991,N_17804);
nand UO_0 (O_0,N_20428,N_22901);
and UO_1 (O_1,N_22517,N_23062);
and UO_2 (O_2,N_22242,N_21944);
and UO_3 (O_3,N_24560,N_20505);
or UO_4 (O_4,N_20709,N_24529);
and UO_5 (O_5,N_23886,N_24834);
nand UO_6 (O_6,N_21375,N_24666);
nor UO_7 (O_7,N_21584,N_22940);
and UO_8 (O_8,N_21489,N_21995);
xnor UO_9 (O_9,N_20020,N_23979);
and UO_10 (O_10,N_24286,N_22976);
nor UO_11 (O_11,N_20330,N_20626);
and UO_12 (O_12,N_23554,N_24226);
nand UO_13 (O_13,N_22275,N_20141);
and UO_14 (O_14,N_24931,N_20175);
nor UO_15 (O_15,N_24592,N_21220);
or UO_16 (O_16,N_24315,N_22464);
xor UO_17 (O_17,N_24853,N_20530);
nor UO_18 (O_18,N_20051,N_24102);
nand UO_19 (O_19,N_23177,N_22992);
or UO_20 (O_20,N_23137,N_24332);
or UO_21 (O_21,N_23473,N_22364);
or UO_22 (O_22,N_20804,N_20356);
nor UO_23 (O_23,N_23928,N_21858);
and UO_24 (O_24,N_23503,N_21330);
or UO_25 (O_25,N_20912,N_21819);
and UO_26 (O_26,N_21946,N_24370);
and UO_27 (O_27,N_23216,N_23582);
nand UO_28 (O_28,N_21133,N_22030);
nor UO_29 (O_29,N_21204,N_21026);
nor UO_30 (O_30,N_24464,N_23020);
nand UO_31 (O_31,N_23936,N_24958);
or UO_32 (O_32,N_21561,N_22107);
xor UO_33 (O_33,N_24523,N_21817);
or UO_34 (O_34,N_20904,N_21101);
or UO_35 (O_35,N_22393,N_22466);
nor UO_36 (O_36,N_21765,N_21901);
or UO_37 (O_37,N_20016,N_24389);
or UO_38 (O_38,N_21723,N_24770);
nand UO_39 (O_39,N_23723,N_22936);
and UO_40 (O_40,N_20797,N_22158);
or UO_41 (O_41,N_21215,N_23262);
nor UO_42 (O_42,N_21301,N_24297);
or UO_43 (O_43,N_22877,N_22622);
and UO_44 (O_44,N_22688,N_20542);
and UO_45 (O_45,N_23189,N_23383);
or UO_46 (O_46,N_21080,N_20315);
and UO_47 (O_47,N_21036,N_24108);
nor UO_48 (O_48,N_21320,N_20683);
nand UO_49 (O_49,N_21966,N_23657);
nand UO_50 (O_50,N_22014,N_21720);
or UO_51 (O_51,N_22382,N_24468);
nand UO_52 (O_52,N_24946,N_23700);
nor UO_53 (O_53,N_20533,N_24861);
or UO_54 (O_54,N_24899,N_24790);
nand UO_55 (O_55,N_21905,N_20259);
nand UO_56 (O_56,N_24534,N_21423);
and UO_57 (O_57,N_24282,N_21877);
or UO_58 (O_58,N_20941,N_24661);
nand UO_59 (O_59,N_23399,N_23633);
and UO_60 (O_60,N_23516,N_22343);
nor UO_61 (O_61,N_24624,N_21702);
nor UO_62 (O_62,N_21013,N_24120);
and UO_63 (O_63,N_20999,N_21211);
nand UO_64 (O_64,N_22598,N_23654);
and UO_65 (O_65,N_23249,N_23025);
nand UO_66 (O_66,N_24670,N_23431);
xor UO_67 (O_67,N_23609,N_22731);
or UO_68 (O_68,N_22284,N_21855);
and UO_69 (O_69,N_24222,N_22018);
and UO_70 (O_70,N_22113,N_20959);
or UO_71 (O_71,N_22804,N_22770);
or UO_72 (O_72,N_22852,N_23217);
and UO_73 (O_73,N_20907,N_22300);
and UO_74 (O_74,N_22495,N_23321);
and UO_75 (O_75,N_23069,N_20691);
nor UO_76 (O_76,N_22069,N_22036);
nand UO_77 (O_77,N_20773,N_21650);
or UO_78 (O_78,N_23378,N_24803);
nand UO_79 (O_79,N_21477,N_24347);
nor UO_80 (O_80,N_23222,N_21803);
or UO_81 (O_81,N_23898,N_22982);
or UO_82 (O_82,N_21506,N_20599);
nor UO_83 (O_83,N_23032,N_20837);
nand UO_84 (O_84,N_23983,N_23155);
or UO_85 (O_85,N_20460,N_23231);
or UO_86 (O_86,N_20423,N_21774);
nor UO_87 (O_87,N_22781,N_23679);
xor UO_88 (O_88,N_21100,N_20081);
and UO_89 (O_89,N_23009,N_23371);
nor UO_90 (O_90,N_21799,N_24986);
and UO_91 (O_91,N_21219,N_22060);
nand UO_92 (O_92,N_21106,N_24037);
and UO_93 (O_93,N_22886,N_21422);
and UO_94 (O_94,N_21728,N_21870);
nand UO_95 (O_95,N_22075,N_23507);
and UO_96 (O_96,N_21351,N_20977);
xnor UO_97 (O_97,N_21150,N_24708);
nor UO_98 (O_98,N_24311,N_24463);
nor UO_99 (O_99,N_20426,N_21078);
nor UO_100 (O_100,N_21170,N_23082);
or UO_101 (O_101,N_23299,N_21923);
nand UO_102 (O_102,N_23131,N_21947);
or UO_103 (O_103,N_21383,N_22739);
nor UO_104 (O_104,N_24554,N_20277);
nand UO_105 (O_105,N_21257,N_22779);
and UO_106 (O_106,N_24049,N_22285);
nor UO_107 (O_107,N_20944,N_24836);
nor UO_108 (O_108,N_24442,N_24025);
nor UO_109 (O_109,N_24299,N_22013);
nor UO_110 (O_110,N_24180,N_23454);
and UO_111 (O_111,N_21781,N_21726);
nand UO_112 (O_112,N_20603,N_24824);
or UO_113 (O_113,N_22006,N_23492);
and UO_114 (O_114,N_20240,N_20586);
and UO_115 (O_115,N_20117,N_22857);
xnor UO_116 (O_116,N_21465,N_24075);
or UO_117 (O_117,N_24218,N_20256);
and UO_118 (O_118,N_24187,N_21750);
nand UO_119 (O_119,N_24132,N_22951);
nor UO_120 (O_120,N_20747,N_22818);
nor UO_121 (O_121,N_22921,N_22851);
and UO_122 (O_122,N_24911,N_23790);
and UO_123 (O_123,N_20017,N_20661);
or UO_124 (O_124,N_21867,N_20763);
and UO_125 (O_125,N_20873,N_24065);
or UO_126 (O_126,N_21488,N_23143);
nor UO_127 (O_127,N_23859,N_20920);
and UO_128 (O_128,N_24147,N_24746);
and UO_129 (O_129,N_22706,N_20805);
nor UO_130 (O_130,N_24493,N_24952);
and UO_131 (O_131,N_21428,N_21826);
nand UO_132 (O_132,N_22863,N_23161);
or UO_133 (O_133,N_20278,N_24190);
nor UO_134 (O_134,N_21532,N_24385);
nor UO_135 (O_135,N_21712,N_22288);
and UO_136 (O_136,N_22338,N_22048);
nand UO_137 (O_137,N_24904,N_22766);
or UO_138 (O_138,N_23574,N_24637);
nand UO_139 (O_139,N_21034,N_24266);
and UO_140 (O_140,N_22783,N_20810);
or UO_141 (O_141,N_20276,N_23565);
or UO_142 (O_142,N_21050,N_24436);
nand UO_143 (O_143,N_21929,N_23498);
or UO_144 (O_144,N_21969,N_24967);
or UO_145 (O_145,N_24500,N_24481);
nand UO_146 (O_146,N_21071,N_22083);
nor UO_147 (O_147,N_23505,N_22313);
nand UO_148 (O_148,N_22103,N_24644);
nand UO_149 (O_149,N_20170,N_24123);
nand UO_150 (O_150,N_24677,N_23170);
or UO_151 (O_151,N_20584,N_24325);
and UO_152 (O_152,N_22438,N_23445);
and UO_153 (O_153,N_23400,N_24198);
nor UO_154 (O_154,N_23775,N_23880);
nor UO_155 (O_155,N_20187,N_22718);
nand UO_156 (O_156,N_21910,N_20079);
and UO_157 (O_157,N_22229,N_20689);
nor UO_158 (O_158,N_22442,N_20345);
nand UO_159 (O_159,N_23406,N_21055);
nor UO_160 (O_160,N_23452,N_21533);
xor UO_161 (O_161,N_23786,N_22281);
nor UO_162 (O_162,N_20642,N_21976);
nor UO_163 (O_163,N_22260,N_24652);
nand UO_164 (O_164,N_23858,N_22828);
or UO_165 (O_165,N_23885,N_23640);
nand UO_166 (O_166,N_21403,N_24636);
or UO_167 (O_167,N_23846,N_24989);
nor UO_168 (O_168,N_23667,N_20302);
nor UO_169 (O_169,N_22677,N_21970);
nand UO_170 (O_170,N_22835,N_21876);
nor UO_171 (O_171,N_23261,N_21154);
and UO_172 (O_172,N_20730,N_21567);
or UO_173 (O_173,N_23678,N_21708);
or UO_174 (O_174,N_20605,N_22259);
nand UO_175 (O_175,N_24997,N_22296);
or UO_176 (O_176,N_20712,N_22150);
and UO_177 (O_177,N_20848,N_21493);
xor UO_178 (O_178,N_21560,N_24409);
and UO_179 (O_179,N_21865,N_21511);
nor UO_180 (O_180,N_22925,N_20785);
or UO_181 (O_181,N_20355,N_22055);
or UO_182 (O_182,N_21908,N_24014);
nand UO_183 (O_183,N_20475,N_22891);
nand UO_184 (O_184,N_24879,N_22400);
or UO_185 (O_185,N_20002,N_21044);
and UO_186 (O_186,N_20334,N_23921);
or UO_187 (O_187,N_24762,N_24936);
nor UO_188 (O_188,N_22843,N_21345);
or UO_189 (O_189,N_20693,N_24469);
nor UO_190 (O_190,N_22855,N_20323);
and UO_191 (O_191,N_24489,N_22590);
nand UO_192 (O_192,N_21129,N_22673);
or UO_193 (O_193,N_22511,N_21636);
nand UO_194 (O_194,N_23192,N_21042);
and UO_195 (O_195,N_23479,N_22581);
nor UO_196 (O_196,N_20112,N_24597);
nand UO_197 (O_197,N_24305,N_22720);
or UO_198 (O_198,N_23124,N_20638);
or UO_199 (O_199,N_21789,N_20148);
nor UO_200 (O_200,N_22805,N_22063);
or UO_201 (O_201,N_22865,N_24687);
nor UO_202 (O_202,N_24369,N_24038);
nand UO_203 (O_203,N_24263,N_20369);
and UO_204 (O_204,N_21656,N_20838);
nor UO_205 (O_205,N_21741,N_20125);
nand UO_206 (O_206,N_24012,N_20310);
or UO_207 (O_207,N_23533,N_20764);
or UO_208 (O_208,N_21235,N_23377);
nand UO_209 (O_209,N_20153,N_23897);
and UO_210 (O_210,N_21614,N_24850);
nand UO_211 (O_211,N_24998,N_20890);
or UO_212 (O_212,N_21121,N_22687);
nor UO_213 (O_213,N_24058,N_23677);
or UO_214 (O_214,N_21729,N_22552);
or UO_215 (O_215,N_20410,N_23636);
nor UO_216 (O_216,N_24783,N_22170);
nand UO_217 (O_217,N_23627,N_23462);
and UO_218 (O_218,N_24026,N_24261);
nand UO_219 (O_219,N_21812,N_22587);
or UO_220 (O_220,N_23270,N_23536);
and UO_221 (O_221,N_24425,N_24698);
or UO_222 (O_222,N_23080,N_24070);
or UO_223 (O_223,N_22469,N_21677);
or UO_224 (O_224,N_21372,N_23015);
and UO_225 (O_225,N_23969,N_22800);
or UO_226 (O_226,N_22972,N_24055);
nand UO_227 (O_227,N_20199,N_24507);
nor UO_228 (O_228,N_20090,N_20579);
xor UO_229 (O_229,N_23050,N_20224);
nand UO_230 (O_230,N_20550,N_24735);
and UO_231 (O_231,N_20508,N_22733);
nand UO_232 (O_232,N_20831,N_22912);
nor UO_233 (O_233,N_22074,N_22784);
or UO_234 (O_234,N_23799,N_23468);
nand UO_235 (O_235,N_24030,N_21061);
or UO_236 (O_236,N_21268,N_22858);
or UO_237 (O_237,N_24738,N_24013);
and UO_238 (O_238,N_22475,N_23949);
or UO_239 (O_239,N_20732,N_21875);
and UO_240 (O_240,N_21572,N_24710);
nand UO_241 (O_241,N_23112,N_22850);
and UO_242 (O_242,N_21521,N_21370);
or UO_243 (O_243,N_20970,N_24300);
nor UO_244 (O_244,N_21766,N_20412);
or UO_245 (O_245,N_20482,N_20481);
nor UO_246 (O_246,N_23193,N_23506);
and UO_247 (O_247,N_22369,N_21737);
or UO_248 (O_248,N_21289,N_20085);
or UO_249 (O_249,N_20802,N_22777);
or UO_250 (O_250,N_21742,N_22072);
nand UO_251 (O_251,N_23185,N_23601);
or UO_252 (O_252,N_20167,N_23126);
and UO_253 (O_253,N_20519,N_22267);
nand UO_254 (O_254,N_20602,N_20131);
nor UO_255 (O_255,N_23976,N_22088);
nand UO_256 (O_256,N_21162,N_22151);
or UO_257 (O_257,N_24486,N_24435);
and UO_258 (O_258,N_21335,N_20592);
or UO_259 (O_259,N_23968,N_23488);
nor UO_260 (O_260,N_22966,N_21283);
or UO_261 (O_261,N_23393,N_21594);
nor UO_262 (O_262,N_21977,N_20514);
xnor UO_263 (O_263,N_22210,N_21989);
nor UO_264 (O_264,N_21184,N_20026);
and UO_265 (O_265,N_20048,N_24182);
and UO_266 (O_266,N_24526,N_24260);
and UO_267 (O_267,N_21024,N_22467);
nand UO_268 (O_268,N_22146,N_22832);
nor UO_269 (O_269,N_23174,N_20161);
nand UO_270 (O_270,N_24525,N_22512);
nand UO_271 (O_271,N_24514,N_22389);
nand UO_272 (O_272,N_21463,N_22973);
or UO_273 (O_273,N_24696,N_23986);
nor UO_274 (O_274,N_21412,N_24103);
and UO_275 (O_275,N_23521,N_22007);
nor UO_276 (O_276,N_22776,N_21808);
or UO_277 (O_277,N_20803,N_22700);
nor UO_278 (O_278,N_22033,N_22652);
nand UO_279 (O_279,N_21543,N_20662);
or UO_280 (O_280,N_21593,N_22910);
and UO_281 (O_281,N_22572,N_20585);
or UO_282 (O_282,N_23571,N_23650);
and UO_283 (O_283,N_21279,N_21209);
or UO_284 (O_284,N_20630,N_24917);
or UO_285 (O_285,N_24818,N_22374);
and UO_286 (O_286,N_23045,N_24128);
and UO_287 (O_287,N_20464,N_24787);
nand UO_288 (O_288,N_21721,N_20160);
nand UO_289 (O_289,N_22683,N_21380);
or UO_290 (O_290,N_23524,N_21710);
nor UO_291 (O_291,N_22497,N_20996);
xnor UO_292 (O_292,N_20431,N_23373);
nand UO_293 (O_293,N_24029,N_23548);
and UO_294 (O_294,N_24502,N_23147);
nor UO_295 (O_295,N_23618,N_23680);
and UO_296 (O_296,N_23484,N_21625);
nor UO_297 (O_297,N_22065,N_21888);
nor UO_298 (O_298,N_24791,N_20840);
xnor UO_299 (O_299,N_20451,N_23964);
nand UO_300 (O_300,N_21986,N_22744);
nor UO_301 (O_301,N_24138,N_24495);
nand UO_302 (O_302,N_20484,N_20842);
and UO_303 (O_303,N_22640,N_24296);
nor UO_304 (O_304,N_22282,N_22047);
xor UO_305 (O_305,N_21309,N_24386);
nand UO_306 (O_306,N_24384,N_21274);
and UO_307 (O_307,N_21214,N_23926);
or UO_308 (O_308,N_21575,N_21099);
or UO_309 (O_309,N_22949,N_21548);
and UO_310 (O_310,N_21985,N_21173);
and UO_311 (O_311,N_23766,N_23096);
nand UO_312 (O_312,N_20172,N_22454);
or UO_313 (O_313,N_21948,N_21248);
nand UO_314 (O_314,N_20313,N_21717);
or UO_315 (O_315,N_21290,N_24840);
nor UO_316 (O_316,N_24934,N_22024);
or UO_317 (O_317,N_21052,N_22591);
nor UO_318 (O_318,N_20381,N_21321);
nor UO_319 (O_319,N_21518,N_20976);
or UO_320 (O_320,N_22017,N_20449);
nor UO_321 (O_321,N_23925,N_24561);
nand UO_322 (O_322,N_20042,N_23117);
nor UO_323 (O_323,N_20253,N_21053);
nor UO_324 (O_324,N_20522,N_23872);
or UO_325 (O_325,N_21060,N_22142);
and UO_326 (O_326,N_23074,N_22071);
nand UO_327 (O_327,N_22751,N_20485);
xnor UO_328 (O_328,N_23892,N_22838);
nor UO_329 (O_329,N_20521,N_22370);
or UO_330 (O_330,N_21176,N_22307);
and UO_331 (O_331,N_21212,N_24140);
nand UO_332 (O_332,N_21821,N_22980);
nand UO_333 (O_333,N_23810,N_20304);
nor UO_334 (O_334,N_23087,N_22401);
or UO_335 (O_335,N_22830,N_21897);
nor UO_336 (O_336,N_20748,N_23496);
xor UO_337 (O_337,N_22578,N_21968);
nor UO_338 (O_338,N_24000,N_21634);
nor UO_339 (O_339,N_24220,N_24028);
or UO_340 (O_340,N_23471,N_24144);
or UO_341 (O_341,N_20151,N_22432);
nand UO_342 (O_342,N_24487,N_22373);
or UO_343 (O_343,N_20795,N_23142);
nor UO_344 (O_344,N_22719,N_20779);
or UO_345 (O_345,N_24335,N_23720);
or UO_346 (O_346,N_22273,N_22385);
or UO_347 (O_347,N_21963,N_24412);
and UO_348 (O_348,N_21681,N_22574);
and UO_349 (O_349,N_20956,N_24546);
or UO_350 (O_350,N_20853,N_22125);
nand UO_351 (O_351,N_23502,N_20295);
or UO_352 (O_352,N_21961,N_20798);
nand UO_353 (O_353,N_20677,N_20535);
nor UO_354 (O_354,N_24161,N_23544);
xnor UO_355 (O_355,N_24172,N_24255);
nand UO_356 (O_356,N_22435,N_20248);
nor UO_357 (O_357,N_20616,N_21862);
nor UO_358 (O_358,N_24635,N_22953);
and UO_359 (O_359,N_24195,N_23881);
and UO_360 (O_360,N_23570,N_20083);
and UO_361 (O_361,N_23336,N_22480);
nand UO_362 (O_362,N_21714,N_20546);
and UO_363 (O_363,N_23624,N_22334);
nor UO_364 (O_364,N_22878,N_24681);
and UO_365 (O_365,N_22233,N_20984);
nand UO_366 (O_366,N_20308,N_22787);
nor UO_367 (O_367,N_22601,N_23209);
nor UO_368 (O_368,N_20214,N_21928);
nor UO_369 (O_369,N_24839,N_20441);
nand UO_370 (O_370,N_23984,N_24018);
nor UO_371 (O_371,N_21621,N_20594);
and UO_372 (O_372,N_22397,N_21020);
nor UO_373 (O_373,N_23577,N_21601);
nand UO_374 (O_374,N_22710,N_20498);
or UO_375 (O_375,N_23763,N_23000);
nor UO_376 (O_376,N_23658,N_23651);
nand UO_377 (O_377,N_23834,N_20527);
nand UO_378 (O_378,N_21245,N_20937);
nor UO_379 (O_379,N_22775,N_20006);
nand UO_380 (O_380,N_23129,N_20939);
or UO_381 (O_381,N_24980,N_21032);
and UO_382 (O_382,N_24665,N_24253);
nand UO_383 (O_383,N_22894,N_22821);
and UO_384 (O_384,N_24362,N_21558);
nand UO_385 (O_385,N_23247,N_23344);
and UO_386 (O_386,N_21449,N_22553);
nand UO_387 (O_387,N_23599,N_21652);
nand UO_388 (O_388,N_22960,N_23944);
nor UO_389 (O_389,N_21122,N_23370);
or UO_390 (O_390,N_21478,N_22924);
nor UO_391 (O_391,N_24785,N_20588);
nor UO_392 (O_392,N_23312,N_24683);
or UO_393 (O_393,N_20990,N_24765);
nand UO_394 (O_394,N_22748,N_22354);
nor UO_395 (O_395,N_24274,N_23990);
and UO_396 (O_396,N_20891,N_24549);
nand UO_397 (O_397,N_20560,N_24242);
nand UO_398 (O_398,N_21534,N_23759);
and UO_399 (O_399,N_22793,N_23001);
and UO_400 (O_400,N_23065,N_21520);
or UO_401 (O_401,N_23739,N_22540);
nand UO_402 (O_402,N_23758,N_21408);
nor UO_403 (O_403,N_20821,N_22729);
nand UO_404 (O_404,N_20646,N_23661);
nor UO_405 (O_405,N_20528,N_20783);
and UO_406 (O_406,N_21243,N_20872);
nor UO_407 (O_407,N_22262,N_24975);
or UO_408 (O_408,N_21603,N_20438);
and UO_409 (O_409,N_22061,N_23291);
or UO_410 (O_410,N_20714,N_22130);
nor UO_411 (O_411,N_22736,N_21902);
nor UO_412 (O_412,N_20960,N_22448);
nand UO_413 (O_413,N_21302,N_20432);
nand UO_414 (O_414,N_21453,N_21475);
and UO_415 (O_415,N_22009,N_21748);
or UO_416 (O_416,N_22682,N_24878);
and UO_417 (O_417,N_22445,N_23780);
and UO_418 (O_418,N_22003,N_23596);
nand UO_419 (O_419,N_24465,N_24969);
and UO_420 (O_420,N_21999,N_20622);
nor UO_421 (O_421,N_23798,N_21300);
nand UO_422 (O_422,N_20680,N_21882);
nor UO_423 (O_423,N_21743,N_23670);
nand UO_424 (O_424,N_23433,N_23830);
nor UO_425 (O_425,N_23444,N_22263);
and UO_426 (O_426,N_21589,N_22726);
and UO_427 (O_427,N_20930,N_24454);
nand UO_428 (O_428,N_24241,N_21455);
or UO_429 (O_429,N_22773,N_23663);
nand UO_430 (O_430,N_24520,N_24280);
nor UO_431 (O_431,N_21421,N_21670);
nand UO_432 (O_432,N_24916,N_21992);
nor UO_433 (O_433,N_24115,N_23597);
and UO_434 (O_434,N_24522,N_21230);
and UO_435 (O_435,N_24133,N_20948);
and UO_436 (O_436,N_21758,N_24877);
or UO_437 (O_437,N_21158,N_22087);
and UO_438 (O_438,N_23620,N_24568);
nor UO_439 (O_439,N_22359,N_23254);
or UO_440 (O_440,N_23342,N_24736);
nand UO_441 (O_441,N_24621,N_24690);
nand UO_442 (O_442,N_21649,N_21433);
and UO_443 (O_443,N_23622,N_24050);
and UO_444 (O_444,N_22276,N_22478);
and UO_445 (O_445,N_20270,N_20264);
nand UO_446 (O_446,N_20133,N_22546);
nor UO_447 (O_447,N_22619,N_20014);
nor UO_448 (O_448,N_23180,N_21030);
nand UO_449 (O_449,N_24498,N_24866);
nand UO_450 (O_450,N_24884,N_23769);
xor UO_451 (O_451,N_22613,N_22527);
and UO_452 (O_452,N_21432,N_23243);
nand UO_453 (O_453,N_21136,N_20715);
xor UO_454 (O_454,N_23653,N_20650);
nand UO_455 (O_455,N_21687,N_24148);
nor UO_456 (O_456,N_22235,N_24405);
nor UO_457 (O_457,N_22839,N_23701);
and UO_458 (O_458,N_23485,N_21392);
nand UO_459 (O_459,N_22458,N_24176);
nand UO_460 (O_460,N_24515,N_22437);
nand UO_461 (O_461,N_23499,N_23176);
or UO_462 (O_462,N_21627,N_22705);
nor UO_463 (O_463,N_24426,N_20577);
and UO_464 (O_464,N_22176,N_23333);
and UO_465 (O_465,N_24688,N_21114);
and UO_466 (O_466,N_24852,N_24593);
xor UO_467 (O_467,N_20497,N_24519);
or UO_468 (O_468,N_21429,N_21339);
or UO_469 (O_469,N_24569,N_22386);
xor UO_470 (O_470,N_24214,N_24772);
nand UO_471 (O_471,N_23891,N_21485);
and UO_472 (O_472,N_21772,N_24448);
and UO_473 (O_473,N_23747,N_22419);
nand UO_474 (O_474,N_23289,N_23381);
nor UO_475 (O_475,N_23256,N_21324);
and UO_476 (O_476,N_21098,N_20574);
or UO_477 (O_477,N_20686,N_21418);
and UO_478 (O_478,N_22215,N_22384);
and UO_479 (O_479,N_24733,N_22836);
nor UO_480 (O_480,N_23649,N_20819);
nor UO_481 (O_481,N_22429,N_23530);
nand UO_482 (O_482,N_21979,N_20903);
or UO_483 (O_483,N_23776,N_22814);
or UO_484 (O_484,N_22051,N_22114);
nand UO_485 (O_485,N_20835,N_24430);
or UO_486 (O_486,N_23803,N_21271);
nor UO_487 (O_487,N_21419,N_23284);
and UO_488 (O_488,N_20046,N_24246);
nor UO_489 (O_489,N_24974,N_20983);
nor UO_490 (O_490,N_22444,N_23267);
or UO_491 (O_491,N_21771,N_24779);
and UO_492 (O_492,N_24869,N_24365);
or UO_493 (O_493,N_20877,N_23740);
nor UO_494 (O_494,N_22620,N_22570);
nand UO_495 (O_495,N_20695,N_23002);
nand UO_496 (O_496,N_22646,N_20576);
xor UO_497 (O_497,N_21029,N_24235);
nor UO_498 (O_498,N_22637,N_24163);
and UO_499 (O_499,N_21957,N_21447);
and UO_500 (O_500,N_21574,N_22477);
nand UO_501 (O_501,N_21844,N_24124);
nand UO_502 (O_502,N_22101,N_21801);
nor UO_503 (O_503,N_21892,N_23874);
nand UO_504 (O_504,N_24822,N_20411);
or UO_505 (O_505,N_24414,N_24777);
nand UO_506 (O_506,N_21155,N_23614);
nand UO_507 (O_507,N_21093,N_23750);
or UO_508 (O_508,N_24867,N_20563);
nand UO_509 (O_509,N_24328,N_22641);
or UO_510 (O_510,N_24472,N_21382);
and UO_511 (O_511,N_22911,N_23992);
or UO_512 (O_512,N_24651,N_23313);
or UO_513 (O_513,N_22841,N_23806);
and UO_514 (O_514,N_23347,N_23483);
and UO_515 (O_515,N_20477,N_24859);
or UO_516 (O_516,N_23272,N_24716);
and UO_517 (O_517,N_23509,N_22989);
nor UO_518 (O_518,N_24063,N_21836);
or UO_519 (O_519,N_22185,N_24518);
nor UO_520 (O_520,N_21285,N_23041);
xnor UO_521 (O_521,N_24640,N_22460);
nand UO_522 (O_522,N_21400,N_23549);
or UO_523 (O_523,N_24860,N_21580);
or UO_524 (O_524,N_21805,N_24566);
or UO_525 (O_525,N_21954,N_20367);
nor UO_526 (O_526,N_24932,N_24827);
or UO_527 (O_527,N_24798,N_21756);
nor UO_528 (O_528,N_23063,N_21698);
and UO_529 (O_529,N_20916,N_20841);
nand UO_530 (O_530,N_21747,N_24954);
or UO_531 (O_531,N_21576,N_21536);
and UO_532 (O_532,N_23430,N_24606);
nand UO_533 (O_533,N_21031,N_20039);
nand UO_534 (O_534,N_24289,N_24098);
or UO_535 (O_535,N_20813,N_24434);
or UO_536 (O_536,N_24087,N_21775);
nor UO_537 (O_537,N_20119,N_23054);
or UO_538 (O_538,N_20075,N_23413);
nand UO_539 (O_539,N_21238,N_22250);
or UO_540 (O_540,N_23016,N_21503);
or UO_541 (O_541,N_23240,N_21866);
and UO_542 (O_542,N_22969,N_21581);
and UO_543 (O_543,N_20503,N_21563);
nor UO_544 (O_544,N_20578,N_23674);
or UO_545 (O_545,N_20337,N_20022);
and UO_546 (O_546,N_21385,N_22658);
nor UO_547 (O_547,N_21437,N_22155);
or UO_548 (O_548,N_22872,N_22782);
or UO_549 (O_549,N_21833,N_21779);
or UO_550 (O_550,N_24734,N_20972);
or UO_551 (O_551,N_24473,N_23118);
or UO_552 (O_552,N_23781,N_20037);
nor UO_553 (O_553,N_24737,N_24725);
nand UO_554 (O_554,N_23306,N_24813);
nor UO_555 (O_555,N_24964,N_21688);
nor UO_556 (O_556,N_20459,N_20881);
nor UO_557 (O_557,N_20597,N_21438);
nor UO_558 (O_558,N_21040,N_24684);
nor UO_559 (O_559,N_20092,N_21673);
or UO_560 (O_560,N_21987,N_22667);
xor UO_561 (O_561,N_22554,N_23078);
and UO_562 (O_562,N_22978,N_21174);
nor UO_563 (O_563,N_24956,N_22410);
xnor UO_564 (O_564,N_21840,N_21542);
nor UO_565 (O_565,N_20705,N_22371);
nor UO_566 (O_566,N_22349,N_20049);
nor UO_567 (O_567,N_23440,N_20127);
and UO_568 (O_568,N_24283,N_23975);
nor UO_569 (O_569,N_23387,N_21852);
nor UO_570 (O_570,N_21094,N_24817);
nor UO_571 (O_571,N_24372,N_20180);
or UO_572 (O_572,N_22534,N_23474);
nand UO_573 (O_573,N_21691,N_21010);
nand UO_574 (O_574,N_20722,N_23580);
nand UO_575 (O_575,N_21927,N_23362);
nand UO_576 (O_576,N_24106,N_23865);
nor UO_577 (O_577,N_21674,N_22955);
nand UO_578 (O_578,N_23295,N_21073);
nor UO_579 (O_579,N_22124,N_24764);
nand UO_580 (O_580,N_20390,N_20060);
or UO_581 (O_581,N_23339,N_24271);
or UO_582 (O_582,N_20387,N_21322);
nor UO_583 (O_583,N_21311,N_24368);
nor UO_584 (O_584,N_24021,N_20724);
or UO_585 (O_585,N_21357,N_21680);
nor UO_586 (O_586,N_24950,N_24979);
nor UO_587 (O_587,N_21007,N_21361);
or UO_588 (O_588,N_24994,N_23127);
or UO_589 (O_589,N_20068,N_23139);
or UO_590 (O_590,N_21871,N_22795);
and UO_591 (O_591,N_24951,N_23187);
nand UO_592 (O_592,N_20829,N_20880);
nor UO_593 (O_593,N_23007,N_22817);
or UO_594 (O_594,N_20955,N_20050);
or UO_595 (O_595,N_21917,N_23102);
nand UO_596 (O_596,N_23477,N_21544);
and UO_597 (O_597,N_20868,N_22365);
or UO_598 (O_598,N_21725,N_20241);
or UO_599 (O_599,N_24715,N_22157);
and UO_600 (O_600,N_20033,N_20306);
xnor UO_601 (O_601,N_22219,N_24512);
nand UO_602 (O_602,N_21070,N_24823);
nand UO_603 (O_603,N_21899,N_23899);
nor UO_604 (O_604,N_23030,N_21252);
nor UO_605 (O_605,N_23138,N_22500);
nor UO_606 (O_606,N_20740,N_22630);
nand UO_607 (O_607,N_20788,N_20975);
nor UO_608 (O_608,N_24503,N_21554);
nor UO_609 (O_609,N_22005,N_22522);
nand UO_610 (O_610,N_24307,N_21295);
nand UO_611 (O_611,N_21624,N_20723);
nor UO_612 (O_612,N_23181,N_23195);
nor UO_613 (O_613,N_23709,N_20839);
or UO_614 (O_614,N_24440,N_23584);
nand UO_615 (O_615,N_20495,N_24816);
nor UO_616 (O_616,N_23294,N_21761);
or UO_617 (O_617,N_21359,N_20556);
and UO_618 (O_618,N_23939,N_23753);
and UO_619 (O_619,N_20031,N_23797);
and UO_620 (O_620,N_22905,N_21355);
nand UO_621 (O_621,N_23408,N_20713);
or UO_622 (O_622,N_23842,N_20100);
xor UO_623 (O_623,N_21839,N_23255);
nor UO_624 (O_624,N_20186,N_20011);
xnor UO_625 (O_625,N_24527,N_20396);
and UO_626 (O_626,N_21854,N_21697);
nor UO_627 (O_627,N_21863,N_24633);
nand UO_628 (O_628,N_22916,N_21795);
or UO_629 (O_629,N_22714,N_20415);
nand UO_630 (O_630,N_24408,N_21568);
and UO_631 (O_631,N_24340,N_23711);
nor UO_632 (O_632,N_23369,N_23794);
or UO_633 (O_633,N_22514,N_21827);
xnor UO_634 (O_634,N_23210,N_21663);
nor UO_635 (O_635,N_23558,N_20378);
nor UO_636 (O_636,N_22900,N_21199);
and UO_637 (O_637,N_22721,N_24375);
nand UO_638 (O_638,N_23742,N_20888);
and UO_639 (O_639,N_23743,N_20103);
or UO_640 (O_640,N_24915,N_20980);
nor UO_641 (O_641,N_21356,N_21587);
or UO_642 (O_642,N_22351,N_20174);
and UO_643 (O_643,N_20271,N_22179);
nor UO_644 (O_644,N_22046,N_20137);
nand UO_645 (O_645,N_23793,N_22529);
nor UO_646 (O_646,N_24113,N_24402);
nor UO_647 (O_647,N_24826,N_21832);
nand UO_648 (O_648,N_21912,N_22383);
or UO_649 (O_649,N_24231,N_20454);
or UO_650 (O_650,N_24539,N_21001);
or UO_651 (O_651,N_21981,N_23263);
nand UO_652 (O_652,N_24609,N_22629);
nor UO_653 (O_653,N_24066,N_21907);
and UO_654 (O_654,N_23033,N_22231);
nor UO_655 (O_655,N_22174,N_20244);
nor UO_656 (O_656,N_23690,N_23635);
and UO_657 (O_657,N_22927,N_22148);
and UO_658 (O_658,N_21605,N_24291);
nor UO_659 (O_659,N_21115,N_22765);
and UO_660 (O_660,N_21793,N_22066);
nand UO_661 (O_661,N_22879,N_23476);
and UO_662 (O_662,N_22119,N_23149);
nand UO_663 (O_663,N_23200,N_20299);
and UO_664 (O_664,N_24720,N_22812);
nand UO_665 (O_665,N_20734,N_22078);
nand UO_666 (O_666,N_24175,N_21617);
nand UO_667 (O_667,N_24264,N_21881);
and UO_668 (O_668,N_23615,N_24755);
or UO_669 (O_669,N_20076,N_24219);
and UO_670 (O_670,N_24712,N_21690);
nor UO_671 (O_671,N_20710,N_21813);
or UO_672 (O_672,N_21009,N_20827);
nor UO_673 (O_673,N_23861,N_23429);
or UO_674 (O_674,N_20273,N_21607);
and UO_675 (O_675,N_21880,N_24099);
nand UO_676 (O_676,N_20118,N_21157);
nand UO_677 (O_677,N_22271,N_20472);
nand UO_678 (O_678,N_24922,N_21286);
and UO_679 (O_679,N_24107,N_22317);
or UO_680 (O_680,N_22605,N_21853);
or UO_681 (O_681,N_21281,N_23526);
and UO_682 (O_682,N_20818,N_20909);
or UO_683 (O_683,N_22195,N_21915);
nor UO_684 (O_684,N_20727,N_24695);
xor UO_685 (O_685,N_24323,N_24727);
or UO_686 (O_686,N_22913,N_20708);
and UO_687 (O_687,N_20126,N_22849);
nor UO_688 (O_688,N_22320,N_21413);
and UO_689 (O_689,N_22257,N_24126);
nor UO_690 (O_690,N_23090,N_23158);
or UO_691 (O_691,N_21198,N_23219);
and UO_692 (O_692,N_22211,N_23783);
and UO_693 (O_693,N_23396,N_21784);
nor UO_694 (O_694,N_24891,N_21409);
nor UO_695 (O_695,N_22199,N_23024);
and UO_696 (O_696,N_22254,N_20058);
nor UO_697 (O_697,N_23363,N_23375);
or UO_698 (O_698,N_24957,N_20736);
xor UO_699 (O_699,N_22624,N_21225);
nand UO_700 (O_700,N_22104,N_20289);
nand UO_701 (O_701,N_21973,N_22516);
or UO_702 (O_702,N_22090,N_22039);
or UO_703 (O_703,N_24937,N_23288);
nor UO_704 (O_704,N_20777,N_23348);
nor UO_705 (O_705,N_22040,N_20636);
or UO_706 (O_706,N_21446,N_22220);
or UO_707 (O_707,N_23461,N_23236);
or UO_708 (O_708,N_20733,N_23450);
nand UO_709 (O_709,N_23911,N_21194);
nor UO_710 (O_710,N_20284,N_20506);
nand UO_711 (O_711,N_24417,N_21481);
or UO_712 (O_712,N_20518,N_21971);
or UO_713 (O_713,N_20318,N_22310);
nand UO_714 (O_714,N_20787,N_24432);
nand UO_715 (O_715,N_23154,N_24159);
nor UO_716 (O_716,N_20405,N_23855);
nor UO_717 (O_717,N_24686,N_22914);
nand UO_718 (O_718,N_24017,N_22476);
or UO_719 (O_719,N_21922,N_21344);
nand UO_720 (O_720,N_23004,N_23738);
or UO_721 (O_721,N_20490,N_20275);
and UO_722 (O_722,N_20462,N_22144);
and UO_723 (O_723,N_23890,N_23585);
nor UO_724 (O_724,N_20251,N_21178);
nor UO_725 (O_725,N_24051,N_21996);
and UO_726 (O_726,N_23027,N_20453);
nand UO_727 (O_727,N_21232,N_21369);
xor UO_728 (O_728,N_20486,N_23953);
or UO_729 (O_729,N_22551,N_22177);
nand UO_730 (O_730,N_21994,N_24920);
nor UO_731 (O_731,N_22084,N_23562);
nand UO_732 (O_732,N_23691,N_20091);
nand UO_733 (O_733,N_23035,N_24378);
or UO_734 (O_734,N_23130,N_22108);
nor UO_735 (O_735,N_21556,N_23629);
nand UO_736 (O_736,N_23151,N_23287);
nand UO_737 (O_737,N_21057,N_24668);
nor UO_738 (O_738,N_23173,N_23755);
or UO_739 (O_739,N_22187,N_23829);
and UO_740 (O_740,N_20860,N_20147);
nor UO_741 (O_741,N_21885,N_23716);
nand UO_742 (O_742,N_20531,N_23621);
nand UO_743 (O_743,N_20399,N_20544);
or UO_744 (O_744,N_20552,N_21695);
or UO_745 (O_745,N_21340,N_22398);
nor UO_746 (O_746,N_22163,N_22829);
nand UO_747 (O_747,N_23481,N_20439);
or UO_748 (O_748,N_22862,N_24262);
nor UO_749 (O_749,N_22653,N_24563);
nand UO_750 (O_750,N_20633,N_23214);
nand UO_751 (O_751,N_21195,N_24317);
nor UO_752 (O_752,N_22968,N_22607);
nand UO_753 (O_753,N_24685,N_24109);
or UO_754 (O_754,N_20237,N_21809);
and UO_755 (O_755,N_21354,N_20502);
or UO_756 (O_756,N_22867,N_23866);
nor UO_757 (O_757,N_24336,N_21715);
or UO_758 (O_758,N_24090,N_20021);
nor UO_759 (O_759,N_22052,N_21626);
or UO_760 (O_760,N_24892,N_21390);
nand UO_761 (O_761,N_20104,N_23593);
or UO_762 (O_762,N_24857,N_23744);
nor UO_763 (O_763,N_21660,N_21474);
nand UO_764 (O_764,N_22861,N_23175);
nor UO_765 (O_765,N_22826,N_24184);
nand UO_766 (O_766,N_22408,N_20882);
nor UO_767 (O_767,N_24135,N_23818);
nand UO_768 (O_768,N_22600,N_24660);
or UO_769 (O_769,N_22264,N_22225);
nand UO_770 (O_770,N_20437,N_24649);
xnor UO_771 (O_771,N_23246,N_21942);
nand UO_772 (O_772,N_21932,N_22755);
nand UO_773 (O_773,N_23955,N_21796);
and UO_774 (O_774,N_22246,N_23202);
and UO_775 (O_775,N_21664,N_23303);
nand UO_776 (O_776,N_24089,N_23948);
nor UO_777 (O_777,N_22112,N_23929);
nor UO_778 (O_778,N_23109,N_21140);
or UO_779 (O_779,N_23860,N_20613);
nand UO_780 (O_780,N_20272,N_23568);
xnor UO_781 (O_781,N_21790,N_20986);
or UO_782 (O_782,N_24723,N_23951);
or UO_783 (O_783,N_23768,N_22864);
nor UO_784 (O_784,N_22306,N_22201);
nand UO_785 (O_785,N_23451,N_21751);
and UO_786 (O_786,N_23034,N_24611);
and UO_787 (O_787,N_20483,N_20200);
or UO_788 (O_788,N_22325,N_23561);
nand UO_789 (O_789,N_24204,N_23543);
nor UO_790 (O_790,N_22926,N_20952);
nand UO_791 (O_791,N_21467,N_22319);
nor UO_792 (O_792,N_20341,N_22345);
or UO_793 (O_793,N_21569,N_20858);
and UO_794 (O_794,N_22859,N_20221);
and UO_795 (O_795,N_21647,N_23325);
nand UO_796 (O_796,N_23540,N_21077);
nor UO_797 (O_797,N_23567,N_23519);
nand UO_798 (O_798,N_24177,N_22870);
and UO_799 (O_799,N_24155,N_23581);
nand UO_800 (O_800,N_22131,N_22801);
or UO_801 (O_801,N_24680,N_22153);
and UO_802 (O_802,N_20353,N_21292);
and UO_803 (O_803,N_23789,N_23594);
nand UO_804 (O_804,N_21769,N_22734);
nand UO_805 (O_805,N_22675,N_23804);
or UO_806 (O_806,N_24318,N_23495);
and UO_807 (O_807,N_21027,N_22671);
or UO_808 (O_808,N_22815,N_24224);
nand UO_809 (O_809,N_22115,N_24622);
nor UO_810 (O_810,N_22452,N_22138);
or UO_811 (O_811,N_24544,N_20931);
and UO_812 (O_812,N_20340,N_20297);
nand UO_813 (O_813,N_21261,N_21091);
and UO_814 (O_814,N_20321,N_23537);
nand UO_815 (O_815,N_22508,N_20312);
or UO_816 (O_816,N_20780,N_24048);
nor UO_817 (O_817,N_22695,N_20116);
nand UO_818 (O_818,N_23266,N_20608);
nor UO_819 (O_819,N_23283,N_20243);
or UO_820 (O_820,N_24162,N_20142);
nor UO_821 (O_821,N_22258,N_21514);
nand UO_822 (O_822,N_21258,N_24112);
nor UO_823 (O_823,N_22352,N_21120);
or UO_824 (O_824,N_23486,N_20238);
nor UO_825 (O_825,N_20242,N_20301);
or UO_826 (O_826,N_21262,N_24457);
and UO_827 (O_827,N_20898,N_20413);
or UO_828 (O_828,N_24745,N_24188);
or UO_829 (O_829,N_24459,N_22035);
nand UO_830 (O_830,N_20233,N_20113);
and UO_831 (O_831,N_21476,N_22923);
nor UO_832 (O_832,N_23647,N_22816);
and UO_833 (O_833,N_20328,N_23290);
nor UO_834 (O_834,N_23970,N_22247);
nand UO_835 (O_835,N_21630,N_24431);
nor UO_836 (O_836,N_20370,N_20181);
nand UO_837 (O_837,N_20676,N_20088);
nand UO_838 (O_838,N_22842,N_24383);
nor UO_839 (O_839,N_22798,N_24632);
nor UO_840 (O_840,N_23997,N_20743);
nor UO_841 (O_841,N_21331,N_23603);
and UO_842 (O_842,N_22450,N_22361);
and UO_843 (O_843,N_22111,N_21530);
xor UO_844 (O_844,N_22227,N_20784);
and UO_845 (O_845,N_24971,N_21381);
nand UO_846 (O_846,N_20555,N_24942);
and UO_847 (O_847,N_20128,N_24044);
nor UO_848 (O_848,N_23305,N_20958);
or UO_849 (O_849,N_20867,N_24653);
nor UO_850 (O_850,N_22693,N_20746);
or UO_851 (O_851,N_22959,N_20029);
and UO_852 (O_852,N_23235,N_22348);
nor UO_853 (O_853,N_24068,N_23541);
or UO_854 (O_854,N_23335,N_20152);
nand UO_855 (O_855,N_22216,N_21213);
nor UO_856 (O_856,N_22709,N_21177);
and UO_857 (O_857,N_23088,N_20627);
nor UO_858 (O_858,N_23197,N_22082);
and UO_859 (O_859,N_24308,N_23411);
nand UO_860 (O_860,N_21760,N_24615);
or UO_861 (O_861,N_24205,N_21596);
nand UO_862 (O_862,N_23196,N_22668);
nor UO_863 (O_863,N_21457,N_22963);
or UO_864 (O_864,N_21227,N_22396);
nor UO_865 (O_865,N_24039,N_21749);
nor UO_866 (O_866,N_21255,N_21410);
nand UO_867 (O_867,N_23981,N_20145);
and UO_868 (O_868,N_23873,N_20973);
and UO_869 (O_869,N_24981,N_22394);
nand UO_870 (O_870,N_24022,N_22580);
xor UO_871 (O_871,N_23669,N_20198);
and UO_872 (O_872,N_21405,N_22149);
and UO_873 (O_873,N_20517,N_23905);
and UO_874 (O_874,N_24377,N_21263);
nand UO_875 (O_875,N_21890,N_24548);
nor UO_876 (O_876,N_21239,N_24993);
nor UO_877 (O_877,N_21221,N_21998);
or UO_878 (O_878,N_22713,N_22190);
nor UO_879 (O_879,N_22730,N_24004);
or UO_880 (O_880,N_21829,N_21739);
and UO_881 (O_881,N_23770,N_24196);
and UO_882 (O_882,N_22681,N_21397);
nor UO_883 (O_883,N_21722,N_24225);
nor UO_884 (O_884,N_22513,N_24245);
or UO_885 (O_885,N_24573,N_21282);
or UO_886 (O_886,N_23935,N_22089);
nor UO_887 (O_887,N_24194,N_20648);
nor UO_888 (O_888,N_22595,N_24773);
or UO_889 (O_889,N_21190,N_22771);
nor UO_890 (O_890,N_23617,N_20886);
or UO_891 (O_891,N_20035,N_21818);
or UO_892 (O_892,N_23269,N_21508);
or UO_893 (O_893,N_24492,N_21072);
nand UO_894 (O_894,N_20182,N_24154);
or UO_895 (O_895,N_21226,N_24423);
xor UO_896 (O_896,N_24889,N_23796);
nand UO_897 (O_897,N_22996,N_21085);
nor UO_898 (O_898,N_20322,N_22750);
and UO_899 (O_899,N_20822,N_24933);
nor UO_900 (O_900,N_24169,N_21005);
nor UO_901 (O_901,N_24497,N_20115);
or UO_902 (O_902,N_22301,N_22764);
nand UO_903 (O_903,N_21291,N_20205);
nand UO_904 (O_904,N_23419,N_21657);
nor UO_905 (O_905,N_23439,N_23410);
nand UO_906 (O_906,N_21655,N_22967);
or UO_907 (O_907,N_21891,N_23525);
and UO_908 (O_908,N_20294,N_23094);
or UO_909 (O_909,N_20865,N_22277);
nor UO_910 (O_910,N_22983,N_23731);
and UO_911 (O_911,N_22347,N_23022);
xor UO_912 (O_912,N_22749,N_24923);
nand UO_913 (O_913,N_21745,N_23814);
nand UO_914 (O_914,N_21092,N_23907);
or UO_915 (O_915,N_24391,N_24658);
and UO_916 (O_916,N_24754,N_20329);
nand UO_917 (O_917,N_23528,N_21724);
nor UO_918 (O_918,N_22742,N_20102);
or UO_919 (O_919,N_23910,N_20737);
nor UO_920 (O_920,N_21332,N_22922);
or UO_921 (O_921,N_22679,N_20385);
nor UO_922 (O_922,N_21643,N_20225);
nand UO_923 (O_923,N_22140,N_23632);
nor UO_924 (O_924,N_24722,N_24310);
and UO_925 (O_925,N_20607,N_23539);
nor UO_926 (O_926,N_22327,N_23551);
or UO_927 (O_927,N_20202,N_21021);
nor UO_928 (O_928,N_21349,N_20658);
or UO_929 (O_929,N_21959,N_24118);
or UO_930 (O_930,N_24863,N_21889);
nor UO_931 (O_931,N_23967,N_21058);
or UO_932 (O_932,N_21557,N_20179);
nand UO_933 (O_933,N_24830,N_22223);
and UO_934 (O_934,N_22760,N_23538);
or UO_935 (O_935,N_22880,N_20815);
and UO_936 (O_936,N_23465,N_21787);
nand UO_937 (O_937,N_23227,N_24930);
and UO_938 (O_938,N_22008,N_24413);
nor UO_939 (O_939,N_23293,N_24505);
or UO_940 (O_940,N_21965,N_22102);
and UO_941 (O_941,N_20287,N_22541);
nand UO_942 (O_942,N_24312,N_24428);
nand UO_943 (O_943,N_23717,N_23453);
nor UO_944 (O_944,N_21394,N_20212);
xor UO_945 (O_945,N_22222,N_22156);
and UO_946 (O_946,N_23591,N_21165);
or UO_947 (O_947,N_23998,N_23351);
or UO_948 (O_948,N_22560,N_20487);
nor UO_949 (O_949,N_23098,N_20361);
xor UO_950 (O_950,N_20754,N_23424);
or UO_951 (O_951,N_23605,N_22791);
or UO_952 (O_952,N_21280,N_23648);
nand UO_953 (O_953,N_21338,N_23501);
or UO_954 (O_954,N_23464,N_22995);
and UO_955 (O_955,N_20591,N_24882);
nand UO_956 (O_956,N_21738,N_21192);
or UO_957 (O_957,N_22651,N_22794);
or UO_958 (O_958,N_22109,N_22631);
and UO_959 (O_959,N_24751,N_20863);
or UO_960 (O_960,N_24081,N_21639);
nand UO_961 (O_961,N_20793,N_24407);
nand UO_962 (O_962,N_20571,N_22439);
or UO_963 (O_963,N_23277,N_20606);
or UO_964 (O_964,N_23675,N_23553);
nor UO_965 (O_965,N_22772,N_20596);
or UO_966 (O_966,N_21193,N_21586);
nand UO_967 (O_967,N_24216,N_20379);
nor UO_968 (O_968,N_21939,N_23820);
nor UO_969 (O_969,N_21138,N_23882);
nor UO_970 (O_970,N_24552,N_23961);
or UO_971 (O_971,N_22678,N_22457);
and UO_972 (O_972,N_23748,N_20226);
xnor UO_973 (O_973,N_21600,N_22422);
xor UO_974 (O_974,N_24602,N_20105);
nand UO_975 (O_975,N_20444,N_20055);
nand UO_976 (O_976,N_22451,N_23320);
nand UO_977 (O_977,N_21377,N_20220);
or UO_978 (O_978,N_22462,N_24580);
and UO_979 (O_979,N_23028,N_21402);
or UO_980 (O_980,N_22321,N_20456);
and UO_981 (O_981,N_24211,N_22097);
nand UO_982 (O_982,N_24862,N_24776);
and UO_983 (O_983,N_20398,N_24125);
or UO_984 (O_984,N_22537,N_24536);
or UO_985 (O_985,N_23864,N_23745);
or UO_986 (O_986,N_20363,N_22542);
and UO_987 (O_987,N_21869,N_21828);
or UO_988 (O_988,N_23229,N_23531);
and UO_989 (O_989,N_24639,N_23853);
nor UO_990 (O_990,N_24269,N_21416);
and UO_991 (O_991,N_22023,N_22575);
or UO_992 (O_992,N_20703,N_21646);
and UO_993 (O_993,N_24719,N_21531);
nor UO_994 (O_994,N_23706,N_23708);
and UO_995 (O_995,N_24832,N_23095);
nand UO_996 (O_996,N_24758,N_23906);
nand UO_997 (O_997,N_20654,N_24820);
or UO_998 (O_998,N_23097,N_20388);
nand UO_999 (O_999,N_21515,N_24618);
and UO_1000 (O_1000,N_23844,N_23713);
nor UO_1001 (O_1001,N_24996,N_20706);
nand UO_1002 (O_1002,N_23140,N_22357);
or UO_1003 (O_1003,N_20262,N_22504);
nand UO_1004 (O_1004,N_24963,N_21389);
xor UO_1005 (O_1005,N_23412,N_21112);
nor UO_1006 (O_1006,N_20982,N_20824);
or UO_1007 (O_1007,N_21254,N_24809);
nor UO_1008 (O_1008,N_21171,N_23167);
and UO_1009 (O_1009,N_22118,N_24327);
xor UO_1010 (O_1010,N_21911,N_24351);
or UO_1011 (O_1011,N_23329,N_23901);
nand UO_1012 (O_1012,N_21342,N_24617);
nand UO_1013 (O_1013,N_24761,N_21143);
and UO_1014 (O_1014,N_24595,N_23510);
nor UO_1015 (O_1015,N_22269,N_21197);
xor UO_1016 (O_1016,N_21229,N_20870);
and UO_1017 (O_1017,N_24343,N_20099);
nand UO_1018 (O_1018,N_20130,N_23259);
and UO_1019 (O_1019,N_24885,N_20003);
nor UO_1020 (O_1020,N_23729,N_21782);
and UO_1021 (O_1021,N_23546,N_22154);
nor UO_1022 (O_1022,N_21169,N_22903);
or UO_1023 (O_1023,N_22253,N_24094);
or UO_1024 (O_1024,N_23346,N_24657);
or UO_1025 (O_1025,N_20447,N_22409);
nor UO_1026 (O_1026,N_23307,N_21082);
nor UO_1027 (O_1027,N_24880,N_23067);
nor UO_1028 (O_1028,N_22208,N_21246);
nor UO_1029 (O_1029,N_24796,N_23322);
nand UO_1030 (O_1030,N_23782,N_22406);
nor UO_1031 (O_1031,N_22311,N_22372);
nand UO_1032 (O_1032,N_23908,N_20249);
xor UO_1033 (O_1033,N_24209,N_23724);
and UO_1034 (O_1034,N_22712,N_22939);
and UO_1035 (O_1035,N_22840,N_24846);
nor UO_1036 (O_1036,N_22539,N_21371);
nand UO_1037 (O_1037,N_24344,N_23762);
or UO_1038 (O_1038,N_24158,N_23815);
or UO_1039 (O_1039,N_23671,N_24093);
and UO_1040 (O_1040,N_21297,N_20121);
and UO_1041 (O_1041,N_23712,N_24421);
and UO_1042 (O_1042,N_23286,N_21399);
and UO_1043 (O_1043,N_24938,N_23616);
or UO_1044 (O_1044,N_24230,N_23446);
or UO_1045 (O_1045,N_21168,N_23048);
nor UO_1046 (O_1046,N_23315,N_21259);
nand UO_1047 (O_1047,N_21997,N_21181);
nor UO_1048 (O_1048,N_20963,N_21967);
nor UO_1049 (O_1049,N_24041,N_20895);
and UO_1050 (O_1050,N_20257,N_20782);
nand UO_1051 (O_1051,N_20391,N_20254);
nor UO_1052 (O_1052,N_24411,N_21604);
and UO_1053 (O_1053,N_24114,N_20933);
nor UO_1054 (O_1054,N_20536,N_20354);
nand UO_1055 (O_1055,N_23300,N_20775);
xor UO_1056 (O_1056,N_21578,N_23710);
or UO_1057 (O_1057,N_24987,N_22888);
or UO_1058 (O_1058,N_20978,N_23734);
and UO_1059 (O_1059,N_20389,N_24626);
or UO_1060 (O_1060,N_23660,N_24876);
or UO_1061 (O_1061,N_21786,N_22323);
nand UO_1062 (O_1062,N_24511,N_20718);
nand UO_1063 (O_1063,N_22908,N_21896);
nand UO_1064 (O_1064,N_23365,N_22965);
xnor UO_1065 (O_1065,N_20589,N_20915);
or UO_1066 (O_1066,N_21495,N_20926);
or UO_1067 (O_1067,N_24929,N_22226);
nand UO_1068 (O_1068,N_23801,N_21276);
nand UO_1069 (O_1069,N_21417,N_21843);
nand UO_1070 (O_1070,N_23455,N_22265);
nand UO_1071 (O_1071,N_24129,N_23995);
nor UO_1072 (O_1072,N_23613,N_22780);
nor UO_1073 (O_1073,N_22332,N_21732);
nand UO_1074 (O_1074,N_20430,N_24907);
or UO_1075 (O_1075,N_23061,N_20040);
or UO_1076 (O_1076,N_21411,N_23011);
or UO_1077 (O_1077,N_24988,N_21241);
and UO_1078 (O_1078,N_20290,N_21272);
or UO_1079 (O_1079,N_20501,N_21631);
nor UO_1080 (O_1080,N_24061,N_21298);
or UO_1081 (O_1081,N_24517,N_21414);
or UO_1082 (O_1082,N_22822,N_24619);
or UO_1083 (O_1083,N_20036,N_23275);
xor UO_1084 (O_1084,N_23511,N_22204);
and UO_1085 (O_1085,N_21611,N_21778);
nand UO_1086 (O_1086,N_21914,N_24628);
and UO_1087 (O_1087,N_23787,N_22038);
or UO_1088 (O_1088,N_23060,N_24322);
and UO_1089 (O_1089,N_20772,N_21458);
nand UO_1090 (O_1090,N_24703,N_21293);
nor UO_1091 (O_1091,N_21016,N_20614);
nor UO_1092 (O_1092,N_23960,N_24543);
nand UO_1093 (O_1093,N_22315,N_20282);
nand UO_1094 (O_1094,N_24079,N_21718);
or UO_1095 (O_1095,N_21172,N_20529);
and UO_1096 (O_1096,N_24122,N_24570);
and UO_1097 (O_1097,N_21879,N_21991);
or UO_1098 (O_1098,N_20816,N_23394);
or UO_1099 (O_1099,N_20107,N_24356);
nand UO_1100 (O_1100,N_24035,N_23135);
nor UO_1101 (O_1101,N_22428,N_24812);
or UO_1102 (O_1102,N_23345,N_23441);
nor UO_1103 (O_1103,N_24947,N_22339);
or UO_1104 (O_1104,N_24338,N_21764);
nand UO_1105 (O_1105,N_20593,N_21051);
nand UO_1106 (O_1106,N_22716,N_21633);
and UO_1107 (O_1107,N_23310,N_24771);
nor UO_1108 (O_1108,N_23828,N_22694);
nor UO_1109 (O_1109,N_21430,N_23868);
and UO_1110 (O_1110,N_24145,N_20346);
and UO_1111 (O_1111,N_24024,N_24394);
or UO_1112 (O_1112,N_24509,N_22871);
nand UO_1113 (O_1113,N_20209,N_20457);
or UO_1114 (O_1114,N_22889,N_22990);
or UO_1115 (O_1115,N_20567,N_20053);
nor UO_1116 (O_1116,N_21887,N_21926);
and UO_1117 (O_1117,N_21434,N_21701);
and UO_1118 (O_1118,N_22415,N_23311);
nand UO_1119 (O_1119,N_21028,N_24924);
nor UO_1120 (O_1120,N_24215,N_21980);
and UO_1121 (O_1121,N_24156,N_24446);
nor UO_1122 (O_1122,N_22547,N_20653);
nor UO_1123 (O_1123,N_23699,N_22806);
or UO_1124 (O_1124,N_20664,N_20792);
or UO_1125 (O_1125,N_21237,N_22881);
and UO_1126 (O_1126,N_22510,N_21373);
nor UO_1127 (O_1127,N_24799,N_22895);
or UO_1128 (O_1128,N_23785,N_24281);
or UO_1129 (O_1129,N_22579,N_21883);
nor UO_1130 (O_1130,N_23547,N_21041);
nand UO_1131 (O_1131,N_20688,N_20801);
and UO_1132 (O_1132,N_21768,N_24034);
nand UO_1133 (O_1133,N_23518,N_23053);
or UO_1134 (O_1134,N_22892,N_24439);
xor UO_1135 (O_1135,N_23101,N_20938);
or UO_1136 (O_1136,N_22792,N_24513);
and UO_1137 (O_1137,N_22041,N_20570);
nor UO_1138 (O_1138,N_24524,N_23788);
nand UO_1139 (O_1139,N_22561,N_20974);
and UO_1140 (O_1140,N_21960,N_22180);
or UO_1141 (O_1141,N_24390,N_24935);
nor UO_1142 (O_1142,N_24697,N_22523);
nor UO_1143 (O_1143,N_21512,N_21398);
and UO_1144 (O_1144,N_24982,N_24788);
nand UO_1145 (O_1145,N_22431,N_20551);
nand UO_1146 (O_1146,N_20469,N_20847);
nor UO_1147 (O_1147,N_20086,N_20769);
nor UO_1148 (O_1148,N_21612,N_21203);
nand UO_1149 (O_1149,N_24139,N_23749);
or UO_1150 (O_1150,N_22985,N_22002);
nor UO_1151 (O_1151,N_24053,N_22509);
and UO_1152 (O_1152,N_22638,N_24903);
nand UO_1153 (O_1153,N_22492,N_21835);
and UO_1154 (O_1154,N_22802,N_23840);
nor UO_1155 (O_1155,N_20332,N_20885);
and UO_1156 (O_1156,N_22186,N_21278);
nand UO_1157 (O_1157,N_22761,N_20283);
nor UO_1158 (O_1158,N_23595,N_20812);
and UO_1159 (O_1159,N_22680,N_21841);
and UO_1160 (O_1160,N_20817,N_22845);
and UO_1161 (O_1161,N_21012,N_22322);
and UO_1162 (O_1162,N_24171,N_20044);
and UO_1163 (O_1163,N_23331,N_23435);
nand UO_1164 (O_1164,N_23352,N_23141);
or UO_1165 (O_1165,N_23727,N_22280);
nand UO_1166 (O_1166,N_21118,N_20559);
or UO_1167 (O_1167,N_22291,N_23550);
or UO_1168 (O_1168,N_23319,N_20206);
and UO_1169 (O_1169,N_21676,N_23282);
or UO_1170 (O_1170,N_24438,N_24366);
and UO_1171 (O_1171,N_23583,N_22848);
nor UO_1172 (O_1172,N_22648,N_24854);
or UO_1173 (O_1173,N_22044,N_21661);
nand UO_1174 (O_1174,N_23070,N_22245);
nor UO_1175 (O_1175,N_20207,N_21180);
nand UO_1176 (O_1176,N_22698,N_20874);
or UO_1177 (O_1177,N_21591,N_24825);
nor UO_1178 (O_1178,N_23159,N_22746);
nand UO_1179 (O_1179,N_21348,N_23493);
nor UO_1180 (O_1180,N_24926,N_23765);
nand UO_1181 (O_1181,N_23121,N_21111);
nor UO_1182 (O_1182,N_22308,N_21256);
nor UO_1183 (O_1183,N_22934,N_21559);
nor UO_1184 (O_1184,N_20580,N_22997);
nor UO_1185 (O_1185,N_24848,N_22920);
and UO_1186 (O_1186,N_22244,N_23838);
and UO_1187 (O_1187,N_22412,N_20525);
nand UO_1188 (O_1188,N_21752,N_22213);
or UO_1189 (O_1189,N_23367,N_20540);
nor UO_1190 (O_1190,N_24249,N_20159);
and UO_1191 (O_1191,N_21909,N_20896);
nor UO_1192 (O_1192,N_24349,N_23588);
or UO_1193 (O_1193,N_20969,N_23133);
or UO_1194 (O_1194,N_22388,N_21127);
or UO_1195 (O_1195,N_22684,N_24331);
nand UO_1196 (O_1196,N_21993,N_23619);
and UO_1197 (O_1197,N_20414,N_23808);
nand UO_1198 (O_1198,N_20851,N_23940);
or UO_1199 (O_1199,N_24789,N_21287);
and UO_1200 (O_1200,N_21325,N_21672);
nor UO_1201 (O_1201,N_24121,N_23252);
nand UO_1202 (O_1202,N_22643,N_21368);
or UO_1203 (O_1203,N_23697,N_20965);
nor UO_1204 (O_1204,N_24728,N_23183);
nor UO_1205 (O_1205,N_24714,N_21472);
nand UO_1206 (O_1206,N_22616,N_22887);
and UO_1207 (O_1207,N_22081,N_23350);
nor UO_1208 (O_1208,N_23655,N_20744);
and UO_1209 (O_1209,N_22141,N_24020);
and UO_1210 (O_1210,N_22757,N_24388);
and UO_1211 (O_1211,N_21699,N_20981);
and UO_1212 (O_1212,N_23494,N_24480);
or UO_1213 (O_1213,N_23644,N_22724);
and UO_1214 (O_1214,N_23642,N_21448);
or UO_1215 (O_1215,N_23166,N_20208);
nand UO_1216 (O_1216,N_22933,N_24707);
or UO_1217 (O_1217,N_22642,N_22609);
nor UO_1218 (O_1218,N_24477,N_23150);
nand UO_1219 (O_1219,N_22717,N_24741);
or UO_1220 (O_1220,N_21516,N_22471);
xnor UO_1221 (O_1221,N_21814,N_24807);
nor UO_1222 (O_1222,N_21480,N_21228);
nand UO_1223 (O_1223,N_20078,N_23920);
nor UO_1224 (O_1224,N_24130,N_24379);
nand UO_1225 (O_1225,N_20836,N_21183);
nand UO_1226 (O_1226,N_22564,N_21307);
nor UO_1227 (O_1227,N_20913,N_22929);
nand UO_1228 (O_1228,N_23040,N_21562);
nand UO_1229 (O_1229,N_24292,N_21719);
nand UO_1230 (O_1230,N_24664,N_24558);
nand UO_1231 (O_1231,N_24256,N_24808);
nor UO_1232 (O_1232,N_23296,N_22127);
nor UO_1233 (O_1233,N_24236,N_21964);
and UO_1234 (O_1234,N_20473,N_24471);
or UO_1235 (O_1235,N_21374,N_20349);
or UO_1236 (O_1236,N_23914,N_24285);
or UO_1237 (O_1237,N_20844,N_23068);
nand UO_1238 (O_1238,N_20582,N_20184);
or UO_1239 (O_1239,N_22318,N_22126);
or UO_1240 (O_1240,N_22122,N_24627);
and UO_1241 (O_1241,N_24623,N_24601);
and UO_1242 (O_1242,N_21538,N_20669);
nand UO_1243 (O_1243,N_21223,N_21466);
and UO_1244 (O_1244,N_21934,N_23172);
nor UO_1245 (O_1245,N_24547,N_21443);
and UO_1246 (O_1246,N_21527,N_21950);
nand UO_1247 (O_1247,N_23760,N_22443);
nor UO_1248 (O_1248,N_20156,N_20109);
nor UO_1249 (O_1249,N_20296,N_20098);
or UO_1250 (O_1250,N_21452,N_24316);
and UO_1251 (O_1251,N_21685,N_22617);
or UO_1252 (O_1252,N_24743,N_23122);
nor UO_1253 (O_1253,N_20351,N_20866);
or UO_1254 (O_1254,N_22330,N_20089);
and UO_1255 (O_1255,N_24747,N_24881);
or UO_1256 (O_1256,N_24767,N_21415);
nor UO_1257 (O_1257,N_21294,N_22116);
xnor UO_1258 (O_1258,N_21346,N_20183);
and UO_1259 (O_1259,N_21103,N_21435);
and UO_1260 (O_1260,N_23427,N_21364);
nor UO_1261 (O_1261,N_22481,N_23385);
or UO_1262 (O_1262,N_20176,N_22488);
nand UO_1263 (O_1263,N_22012,N_22809);
nor UO_1264 (O_1264,N_20489,N_23662);
nor UO_1265 (O_1265,N_24992,N_22723);
or UO_1266 (O_1266,N_20728,N_22831);
nand UO_1267 (O_1267,N_23145,N_22690);
nor UO_1268 (O_1268,N_24844,N_22844);
and UO_1269 (O_1269,N_22184,N_22524);
or UO_1270 (O_1270,N_22015,N_20700);
or UO_1271 (O_1271,N_23566,N_23026);
xnor UO_1272 (O_1272,N_24313,N_22292);
and UO_1273 (O_1273,N_24873,N_23081);
or UO_1274 (O_1274,N_22042,N_21788);
nor UO_1275 (O_1275,N_22100,N_23386);
or UO_1276 (O_1276,N_21850,N_21925);
nor UO_1277 (O_1277,N_21820,N_24901);
and UO_1278 (O_1278,N_22395,N_22050);
nor UO_1279 (O_1279,N_24679,N_22762);
xnor UO_1280 (O_1280,N_20434,N_20065);
nor UO_1281 (O_1281,N_22350,N_22268);
nor UO_1282 (O_1282,N_23316,N_22381);
nand UO_1283 (O_1283,N_24074,N_21904);
or UO_1284 (O_1284,N_23285,N_21851);
and UO_1285 (O_1285,N_23576,N_20887);
nand UO_1286 (O_1286,N_20336,N_21119);
nand UO_1287 (O_1287,N_20998,N_21754);
nand UO_1288 (O_1288,N_24483,N_20013);
and UO_1289 (O_1289,N_24870,N_23113);
and UO_1290 (O_1290,N_22763,N_23863);
or UO_1291 (O_1291,N_23384,N_23148);
nand UO_1292 (O_1292,N_23168,N_23630);
nor UO_1293 (O_1293,N_24342,N_23973);
or UO_1294 (O_1294,N_22670,N_21334);
or UO_1295 (O_1295,N_22866,N_21231);
or UO_1296 (O_1296,N_22117,N_23260);
nand UO_1297 (O_1297,N_23332,N_23751);
and UO_1298 (O_1298,N_20196,N_20767);
or UO_1299 (O_1299,N_22421,N_20600);
and UO_1300 (O_1300,N_24174,N_24069);
nor UO_1301 (O_1301,N_21668,N_22049);
or UO_1302 (O_1302,N_20028,N_20989);
and UO_1303 (O_1303,N_23610,N_20080);
and UO_1304 (O_1304,N_20154,N_24810);
and UO_1305 (O_1305,N_24865,N_24742);
and UO_1306 (O_1306,N_24795,N_22390);
or UO_1307 (O_1307,N_21744,N_21460);
nand UO_1308 (O_1308,N_20768,N_21471);
nor UO_1309 (O_1309,N_20435,N_23805);
or UO_1310 (O_1310,N_20988,N_21251);
or UO_1311 (O_1311,N_24858,N_23448);
nor UO_1312 (O_1312,N_24259,N_22885);
nor UO_1313 (O_1313,N_21806,N_24200);
nand UO_1314 (O_1314,N_21189,N_22999);
nand UO_1315 (O_1315,N_22623,N_24164);
and UO_1316 (O_1316,N_21678,N_22531);
nor UO_1317 (O_1317,N_20095,N_20619);
and UO_1318 (O_1318,N_23017,N_21090);
and UO_1319 (O_1319,N_24600,N_24499);
and UO_1320 (O_1320,N_22214,N_20624);
nand UO_1321 (O_1321,N_23934,N_20702);
nand UO_1322 (O_1322,N_20419,N_21940);
nor UO_1323 (O_1323,N_24032,N_24913);
nand UO_1324 (O_1324,N_24581,N_22860);
or UO_1325 (O_1325,N_23592,N_21265);
nor UO_1326 (O_1326,N_24782,N_22360);
nor UO_1327 (O_1327,N_24210,N_23849);
nand UO_1328 (O_1328,N_21273,N_24766);
and UO_1329 (O_1329,N_20493,N_21022);
and UO_1330 (O_1330,N_23884,N_24646);
nor UO_1331 (O_1331,N_24928,N_20392);
nor UO_1332 (O_1332,N_23684,N_24551);
nand UO_1333 (O_1333,N_20373,N_21145);
nand UO_1334 (O_1334,N_23761,N_21483);
xor UO_1335 (O_1335,N_21008,N_20309);
or UO_1336 (O_1336,N_21955,N_21366);
and UO_1337 (O_1337,N_20692,N_22011);
nand UO_1338 (O_1338,N_22091,N_24067);
nand UO_1339 (O_1339,N_21736,N_20071);
nand UO_1340 (O_1340,N_22634,N_24704);
or UO_1341 (O_1341,N_21200,N_23589);
nand UO_1342 (O_1342,N_20394,N_23924);
nand UO_1343 (O_1343,N_22434,N_20778);
and UO_1344 (O_1344,N_22468,N_21974);
and UO_1345 (O_1345,N_21665,N_20365);
or UO_1346 (O_1346,N_22482,N_22568);
or UO_1347 (O_1347,N_20823,N_23089);
nand UO_1348 (O_1348,N_23364,N_24359);
and UO_1349 (O_1349,N_21011,N_22586);
nand UO_1350 (O_1350,N_21734,N_21566);
nor UO_1351 (O_1351,N_22943,N_20281);
nand UO_1352 (O_1352,N_24101,N_24485);
and UO_1353 (O_1353,N_21696,N_24793);
nand UO_1354 (O_1354,N_21857,N_21845);
nand UO_1355 (O_1355,N_24564,N_24961);
or UO_1356 (O_1356,N_20436,N_21623);
nand UO_1357 (O_1357,N_20690,N_23856);
nor UO_1358 (O_1358,N_23046,N_21608);
or UO_1359 (O_1359,N_20445,N_20372);
nand UO_1360 (O_1360,N_22896,N_20631);
nor UO_1361 (O_1361,N_23366,N_20018);
and UO_1362 (O_1362,N_24898,N_23927);
nand UO_1363 (O_1363,N_21792,N_20366);
nor UO_1364 (O_1364,N_22240,N_21222);
nand UO_1365 (O_1365,N_24814,N_22232);
and UO_1366 (O_1366,N_20994,N_22294);
or UO_1367 (O_1367,N_22137,N_22152);
and UO_1368 (O_1368,N_20066,N_24054);
nand UO_1369 (O_1369,N_22628,N_22493);
or UO_1370 (O_1370,N_24990,N_20452);
and UO_1371 (O_1371,N_22380,N_24673);
nor UO_1372 (O_1372,N_20455,N_20260);
nor UO_1373 (O_1373,N_23128,N_23703);
or UO_1374 (O_1374,N_20500,N_24452);
nor UO_1375 (O_1375,N_24780,N_20005);
or UO_1376 (O_1376,N_22080,N_22079);
or UO_1377 (O_1377,N_20239,N_22212);
or UO_1378 (O_1378,N_21469,N_22191);
nor UO_1379 (O_1379,N_20991,N_20826);
nor UO_1380 (O_1380,N_24167,N_23778);
nor UO_1381 (O_1381,N_21047,N_23253);
or UO_1382 (O_1382,N_23031,N_23851);
nand UO_1383 (O_1383,N_24410,N_20557);
or UO_1384 (O_1384,N_23076,N_20446);
or UO_1385 (O_1385,N_21284,N_22133);
and UO_1386 (O_1386,N_22946,N_20632);
nor UO_1387 (O_1387,N_21333,N_24571);
nor UO_1388 (O_1388,N_24160,N_21179);
and UO_1389 (O_1389,N_20307,N_24272);
and UO_1390 (O_1390,N_20056,N_23809);
or UO_1391 (O_1391,N_21062,N_24638);
nor UO_1392 (O_1392,N_20231,N_24303);
or UO_1393 (O_1393,N_21671,N_22594);
nor UO_1394 (O_1394,N_21224,N_20526);
nand UO_1395 (O_1395,N_20007,N_23664);
nand UO_1396 (O_1396,N_22356,N_22535);
and UO_1397 (O_1397,N_22316,N_20401);
or UO_1398 (O_1398,N_22727,N_23273);
and UO_1399 (O_1399,N_24603,N_24538);
nor UO_1400 (O_1400,N_24691,N_23211);
nand UO_1401 (O_1401,N_20374,N_20032);
nor UO_1402 (O_1402,N_22016,N_22503);
and UO_1403 (O_1403,N_22399,N_23042);
and UO_1404 (O_1404,N_23250,N_23199);
nor UO_1405 (O_1405,N_24944,N_22543);
or UO_1406 (O_1406,N_24141,N_21496);
nor UO_1407 (O_1407,N_24398,N_22699);
nand UO_1408 (O_1408,N_22172,N_22181);
and UO_1409 (O_1409,N_20656,N_24545);
nor UO_1410 (O_1410,N_21196,N_24016);
and UO_1411 (O_1411,N_21004,N_23144);
nand UO_1412 (O_1412,N_23638,N_22945);
or UO_1413 (O_1413,N_23157,N_23602);
nand UO_1414 (O_1414,N_21109,N_20957);
nand UO_1415 (O_1415,N_24491,N_23274);
nand UO_1416 (O_1416,N_22346,N_21930);
and UO_1417 (O_1417,N_24373,N_20538);
nor UO_1418 (O_1418,N_22413,N_20716);
xor UO_1419 (O_1419,N_24111,N_24590);
or UO_1420 (O_1420,N_20097,N_20352);
and UO_1421 (O_1421,N_20448,N_20750);
nor UO_1422 (O_1422,N_24419,N_20950);
and UO_1423 (O_1423,N_21837,N_23698);
or UO_1424 (O_1424,N_21439,N_22198);
or UO_1425 (O_1425,N_23918,N_24501);
or UO_1426 (O_1426,N_24003,N_21379);
nor UO_1427 (O_1427,N_22145,N_24577);
nand UO_1428 (O_1428,N_24775,N_21962);
nor UO_1429 (O_1429,N_23010,N_23937);
nand UO_1430 (O_1430,N_21275,N_24856);
or UO_1431 (O_1431,N_21640,N_21861);
nand UO_1432 (O_1432,N_20478,N_21731);
or UO_1433 (O_1433,N_22314,N_24181);
nor UO_1434 (O_1434,N_24800,N_20421);
and UO_1435 (O_1435,N_21525,N_20303);
or UO_1436 (O_1436,N_20671,N_23725);
nor UO_1437 (O_1437,N_23877,N_21523);
nand UO_1438 (O_1438,N_21900,N_21498);
and UO_1439 (O_1439,N_24290,N_23223);
or UO_1440 (O_1440,N_23831,N_22956);
nor UO_1441 (O_1441,N_21425,N_22676);
nor UO_1442 (O_1442,N_23361,N_21507);
nor UO_1443 (O_1443,N_21770,N_24586);
or UO_1444 (O_1444,N_20590,N_22582);
xnor UO_1445 (O_1445,N_21218,N_24756);
nand UO_1446 (O_1446,N_20707,N_20681);
and UO_1447 (O_1447,N_21767,N_24833);
and UO_1448 (O_1448,N_21097,N_23707);
and UO_1449 (O_1449,N_21654,N_24309);
or UO_1450 (O_1450,N_20513,N_22455);
xor UO_1451 (O_1451,N_23688,N_21816);
nand UO_1452 (O_1452,N_24671,N_24441);
nor UO_1453 (O_1453,N_21250,N_20467);
nor UO_1454 (O_1454,N_22621,N_21037);
and UO_1455 (O_1455,N_21583,N_23646);
or UO_1456 (O_1456,N_22147,N_24940);
nor UO_1457 (O_1457,N_21395,N_20548);
or UO_1458 (O_1458,N_23779,N_24119);
nand UO_1459 (O_1459,N_24752,N_21615);
and UO_1460 (O_1460,N_20380,N_23264);
nor UO_1461 (O_1461,N_24273,N_22379);
xor UO_1462 (O_1462,N_24479,N_20134);
and UO_1463 (O_1463,N_21924,N_24575);
nand UO_1464 (O_1464,N_23545,N_24784);
nand UO_1465 (O_1465,N_20338,N_24165);
xnor UO_1466 (O_1466,N_22655,N_21535);
nand UO_1467 (O_1467,N_21755,N_23756);
nand UO_1468 (O_1468,N_20360,N_24669);
or UO_1469 (O_1469,N_23982,N_24819);
nand UO_1470 (O_1470,N_23563,N_21776);
or UO_1471 (O_1471,N_22456,N_22919);
nor UO_1472 (O_1472,N_20634,N_20670);
or UO_1473 (O_1473,N_22299,N_24949);
or UO_1474 (O_1474,N_22032,N_20757);
or UO_1475 (O_1475,N_22704,N_22053);
nand UO_1476 (O_1476,N_21089,N_21205);
or UO_1477 (O_1477,N_23395,N_22194);
nand UO_1478 (O_1478,N_22689,N_23134);
or UO_1479 (O_1479,N_21679,N_23338);
and UO_1480 (O_1480,N_23152,N_21142);
or UO_1481 (O_1481,N_23919,N_22326);
nand UO_1482 (O_1482,N_23308,N_24252);
nand UO_1483 (O_1483,N_24278,N_20745);
or UO_1484 (O_1484,N_22906,N_23513);
nand UO_1485 (O_1485,N_22274,N_22239);
nor UO_1486 (O_1486,N_21350,N_20504);
nor UO_1487 (O_1487,N_24912,N_23523);
nand UO_1488 (O_1488,N_22424,N_20843);
and UO_1489 (O_1489,N_23472,N_23996);
or UO_1490 (O_1490,N_24675,N_24092);
and UO_1491 (O_1491,N_24607,N_21504);
xor UO_1492 (O_1492,N_21975,N_21347);
nor UO_1493 (O_1493,N_20417,N_22612);
or UO_1494 (O_1494,N_22928,N_24324);
or UO_1495 (O_1495,N_22436,N_20876);
or UO_1496 (O_1496,N_21894,N_22335);
nor UO_1497 (O_1497,N_21529,N_20362);
xnor UO_1498 (O_1498,N_21794,N_24361);
or UO_1499 (O_1499,N_21079,N_24927);
and UO_1500 (O_1500,N_20047,N_22597);
nand UO_1501 (O_1501,N_24229,N_24717);
nor UO_1502 (O_1502,N_22491,N_22827);
nor UO_1503 (O_1503,N_20343,N_20789);
xnor UO_1504 (O_1504,N_20979,N_20293);
or UO_1505 (O_1505,N_22414,N_23248);
nand UO_1506 (O_1506,N_23281,N_23822);
nor UO_1507 (O_1507,N_21444,N_24461);
or UO_1508 (O_1508,N_23077,N_22697);
or UO_1509 (O_1509,N_20923,N_21187);
or UO_1510 (O_1510,N_23392,N_24656);
and UO_1511 (O_1511,N_24330,N_21006);
nand UO_1512 (O_1512,N_21933,N_22701);
and UO_1513 (O_1513,N_21182,N_20516);
or UO_1514 (O_1514,N_24886,N_22070);
nand UO_1515 (O_1515,N_23425,N_24794);
or UO_1516 (O_1516,N_23737,N_22178);
and UO_1517 (O_1517,N_20945,N_21123);
and UO_1518 (O_1518,N_20376,N_22000);
nor UO_1519 (O_1519,N_23835,N_21323);
nand UO_1520 (O_1520,N_22203,N_21951);
nand UO_1521 (O_1521,N_24418,N_23811);
or UO_1522 (O_1522,N_20572,N_20203);
nor UO_1523 (O_1523,N_20034,N_23508);
nor UO_1524 (O_1524,N_23146,N_24948);
nand UO_1525 (O_1525,N_23943,N_22278);
nor UO_1526 (O_1526,N_21105,N_22205);
nor UO_1527 (O_1527,N_20111,N_20922);
and UO_1528 (O_1528,N_24393,N_21086);
nor UO_1529 (O_1529,N_20245,N_20776);
or UO_1530 (O_1530,N_23887,N_24470);
or UO_1531 (O_1531,N_20684,N_22566);
and UO_1532 (O_1532,N_22237,N_22737);
and UO_1533 (O_1533,N_21895,N_24203);
nand UO_1534 (O_1534,N_23003,N_22159);
nor UO_1535 (O_1535,N_23879,N_21602);
nand UO_1536 (O_1536,N_23388,N_21023);
nand UO_1537 (O_1537,N_23522,N_22917);
nor UO_1538 (O_1538,N_24843,N_24084);
nor UO_1539 (O_1539,N_20794,N_24380);
nor UO_1540 (O_1540,N_20364,N_20124);
nand UO_1541 (O_1541,N_22569,N_22532);
nand UO_1542 (O_1542,N_21941,N_20027);
or UO_1543 (O_1543,N_22536,N_22001);
or UO_1544 (O_1544,N_23845,N_23883);
or UO_1545 (O_1545,N_24137,N_20643);
nor UO_1546 (O_1546,N_21038,N_20751);
and UO_1547 (O_1547,N_24213,N_23224);
and UO_1548 (O_1548,N_22577,N_20547);
nor UO_1549 (O_1549,N_21606,N_24488);
and UO_1550 (O_1550,N_23774,N_23232);
nand UO_1551 (O_1551,N_20057,N_24835);
nand UO_1552 (O_1552,N_23895,N_23191);
and UO_1553 (O_1553,N_21487,N_24589);
and UO_1554 (O_1554,N_24400,N_23091);
or UO_1555 (O_1555,N_21167,N_21555);
nor UO_1556 (O_1556,N_21547,N_24183);
and UO_1557 (O_1557,N_24082,N_20879);
and UO_1558 (O_1558,N_21735,N_23013);
and UO_1559 (O_1559,N_24427,N_23466);
and UO_1560 (O_1560,N_23721,N_23106);
and UO_1561 (O_1561,N_24007,N_20232);
nor UO_1562 (O_1562,N_21494,N_21337);
xor UO_1563 (O_1563,N_22752,N_21486);
nor UO_1564 (O_1564,N_24179,N_24136);
and UO_1565 (O_1565,N_22251,N_23972);
nand UO_1566 (O_1566,N_21191,N_21045);
nand UO_1567 (O_1567,N_23641,N_21500);
and UO_1568 (O_1568,N_23039,N_21124);
nor UO_1569 (O_1569,N_22037,N_20889);
and UO_1570 (O_1570,N_22899,N_24797);
nor UO_1571 (O_1571,N_22076,N_22756);
and UO_1572 (O_1572,N_24073,N_23104);
nand UO_1573 (O_1573,N_23271,N_22753);
nor UO_1574 (O_1574,N_20894,N_22562);
nand UO_1575 (O_1575,N_23730,N_22856);
nor UO_1576 (O_1576,N_20859,N_21288);
or UO_1577 (O_1577,N_20621,N_24178);
nor UO_1578 (O_1578,N_23372,N_20951);
and UO_1579 (O_1579,N_23652,N_21937);
or UO_1580 (O_1580,N_21048,N_22603);
and UO_1581 (O_1581,N_21682,N_20729);
and UO_1582 (O_1582,N_21054,N_20476);
or UO_1583 (O_1583,N_23397,N_21528);
or UO_1584 (O_1584,N_20809,N_21269);
or UO_1585 (O_1585,N_22632,N_23867);
or UO_1586 (O_1586,N_23100,N_22873);
or UO_1587 (O_1587,N_23317,N_23165);
nand UO_1588 (O_1588,N_22368,N_23239);
or UO_1589 (O_1589,N_21358,N_21916);
and UO_1590 (O_1590,N_24240,N_20286);
and UO_1591 (O_1591,N_21207,N_20191);
nor UO_1592 (O_1592,N_20507,N_21144);
nor UO_1593 (O_1593,N_23912,N_22548);
or UO_1594 (O_1594,N_22813,N_23380);
or UO_1595 (O_1595,N_23297,N_20573);
xor UO_1596 (O_1596,N_23218,N_23682);
nor UO_1597 (O_1597,N_24516,N_20136);
and UO_1598 (O_1598,N_23946,N_20188);
nand UO_1599 (O_1599,N_23115,N_22134);
and UO_1600 (O_1600,N_22062,N_24699);
nand UO_1601 (O_1601,N_22521,N_21519);
nor UO_1602 (O_1602,N_22576,N_20993);
nor UO_1603 (O_1603,N_20178,N_23491);
nand UO_1604 (O_1604,N_24550,N_21056);
and UO_1605 (O_1605,N_24702,N_21074);
and UO_1606 (O_1606,N_23057,N_24294);
or UO_1607 (O_1607,N_21524,N_23280);
and UO_1608 (O_1608,N_21798,N_22702);
and UO_1609 (O_1609,N_24970,N_20645);
or UO_1610 (O_1610,N_23205,N_24583);
nor UO_1611 (O_1611,N_22328,N_24005);
nor UO_1612 (O_1612,N_24587,N_20311);
nor UO_1613 (O_1613,N_20929,N_24732);
and UO_1614 (O_1614,N_21815,N_20846);
nor UO_1615 (O_1615,N_22962,N_23005);
or UO_1616 (O_1616,N_24072,N_21019);
nand UO_1617 (O_1617,N_23837,N_23391);
xor UO_1618 (O_1618,N_24237,N_22192);
nor UO_1619 (O_1619,N_23421,N_23184);
nand UO_1620 (O_1620,N_23014,N_23909);
nand UO_1621 (O_1621,N_20796,N_23871);
and UO_1622 (O_1622,N_22599,N_24613);
nand UO_1623 (O_1623,N_24718,N_20347);
nor UO_1624 (O_1624,N_20316,N_22092);
and UO_1625 (O_1625,N_24676,N_24875);
nor UO_1626 (O_1626,N_22302,N_23357);
nand UO_1627 (O_1627,N_22711,N_24667);
and UO_1628 (O_1628,N_20561,N_21156);
and UO_1629 (O_1629,N_23966,N_23816);
or UO_1630 (O_1630,N_23672,N_20871);
nor UO_1631 (O_1631,N_24279,N_22189);
nor UO_1632 (O_1632,N_24334,N_20954);
nor UO_1633 (O_1633,N_21613,N_23469);
or UO_1634 (O_1634,N_23228,N_20025);
nand UO_1635 (O_1635,N_24535,N_21327);
nand UO_1636 (O_1636,N_24458,N_20565);
nand UO_1637 (O_1637,N_22528,N_21903);
nand UO_1638 (O_1638,N_22067,N_24406);
and UO_1639 (O_1639,N_23038,N_21753);
or UO_1640 (O_1640,N_21236,N_20072);
nor UO_1641 (O_1641,N_24792,N_24433);
and UO_1642 (O_1642,N_23085,N_24908);
or UO_1643 (O_1643,N_21860,N_23843);
nand UO_1644 (O_1644,N_21083,N_22938);
or UO_1645 (O_1645,N_20162,N_23105);
nand UO_1646 (O_1646,N_20921,N_22897);
nand UO_1647 (O_1647,N_20190,N_22573);
nor UO_1648 (O_1648,N_23301,N_24841);
and UO_1649 (O_1649,N_21893,N_24689);
nor UO_1650 (O_1650,N_23162,N_21763);
nand UO_1651 (O_1651,N_23714,N_24474);
and UO_1652 (O_1652,N_20862,N_20869);
nor UO_1653 (O_1653,N_21620,N_23587);
and UO_1654 (O_1654,N_22135,N_20659);
or UO_1655 (O_1655,N_23328,N_24620);
nand UO_1656 (O_1656,N_20657,N_22028);
or UO_1657 (O_1657,N_20252,N_20675);
nor UO_1658 (O_1658,N_22355,N_22169);
and UO_1659 (O_1659,N_21049,N_20265);
or UO_1660 (O_1660,N_20229,N_23208);
nor UO_1661 (O_1661,N_21577,N_21018);
nor UO_1662 (O_1662,N_23626,N_22728);
and UO_1663 (O_1663,N_23534,N_24451);
nand UO_1664 (O_1664,N_23018,N_24244);
or UO_1665 (O_1665,N_24890,N_23482);
or UO_1666 (O_1666,N_24460,N_21318);
nand UO_1667 (O_1667,N_20765,N_22618);
nand UO_1668 (O_1668,N_22166,N_21635);
nand UO_1669 (O_1669,N_22160,N_23358);
or UO_1670 (O_1670,N_23125,N_23292);
nand UO_1671 (O_1671,N_22819,N_20665);
and UO_1672 (O_1672,N_24999,N_20106);
nor UO_1673 (O_1673,N_21540,N_21240);
and UO_1674 (O_1674,N_20403,N_21598);
nand UO_1675 (O_1675,N_20884,N_23194);
nand UO_1676 (O_1676,N_23404,N_20064);
and UO_1677 (O_1677,N_22639,N_23436);
or UO_1678 (O_1678,N_23839,N_22974);
and UO_1679 (O_1679,N_20649,N_24510);
nor UO_1680 (O_1680,N_20008,N_22252);
or UO_1681 (O_1681,N_20324,N_21553);
and UO_1682 (O_1682,N_23659,N_20479);
or UO_1683 (O_1683,N_24849,N_21666);
nor UO_1684 (O_1684,N_23237,N_24995);
nand UO_1685 (O_1685,N_23086,N_23959);
and UO_1686 (O_1686,N_20721,N_21146);
nand UO_1687 (O_1687,N_21161,N_20629);
xor UO_1688 (O_1688,N_20144,N_22696);
xnor UO_1689 (O_1689,N_20618,N_22649);
xor UO_1690 (O_1690,N_22583,N_20108);
nand UO_1691 (O_1691,N_23977,N_20192);
and UO_1692 (O_1692,N_21983,N_20230);
nand UO_1693 (O_1693,N_22453,N_24574);
nand UO_1694 (O_1694,N_23552,N_23500);
nand UO_1695 (O_1695,N_24598,N_22692);
nor UO_1696 (O_1696,N_20427,N_22559);
and UO_1697 (O_1697,N_22774,N_22026);
and UO_1698 (O_1698,N_23611,N_24659);
or UO_1699 (O_1699,N_21773,N_21270);
or UO_1700 (O_1700,N_24337,N_21886);
nor UO_1701 (O_1701,N_24821,N_20041);
and UO_1702 (O_1702,N_22236,N_24494);
or UO_1703 (O_1703,N_22984,N_23359);
nand UO_1704 (O_1704,N_20756,N_21588);
nor UO_1705 (O_1705,N_22376,N_20549);
nor UO_1706 (O_1706,N_23974,N_22799);
nor UO_1707 (O_1707,N_20288,N_24804);
and UO_1708 (O_1708,N_22725,N_22767);
nor UO_1709 (O_1709,N_24168,N_20901);
nand UO_1710 (O_1710,N_24036,N_20491);
xor UO_1711 (O_1711,N_20139,N_22611);
xor UO_1712 (O_1712,N_22743,N_22106);
and UO_1713 (O_1713,N_21482,N_22502);
and UO_1714 (O_1714,N_24247,N_23244);
and UO_1715 (O_1715,N_22958,N_20935);
and UO_1716 (O_1716,N_23978,N_23736);
nand UO_1717 (O_1717,N_21938,N_21509);
nand UO_1718 (O_1718,N_23206,N_21490);
nor UO_1719 (O_1719,N_23569,N_23324);
nand UO_1720 (O_1720,N_23279,N_24104);
and UO_1721 (O_1721,N_24608,N_20834);
nand UO_1722 (O_1722,N_20562,N_22937);
or UO_1723 (O_1723,N_20852,N_20697);
nor UO_1724 (O_1724,N_20266,N_20122);
nor UO_1725 (O_1725,N_22824,N_24900);
nor UO_1726 (O_1726,N_20155,N_22722);
nor UO_1727 (O_1727,N_22426,N_20520);
or UO_1728 (O_1728,N_22987,N_23993);
nand UO_1729 (O_1729,N_21616,N_20442);
nor UO_1730 (O_1730,N_21132,N_21810);
or UO_1731 (O_1731,N_24395,N_20758);
nor UO_1732 (O_1732,N_20635,N_21343);
nor UO_1733 (O_1733,N_23915,N_21233);
nor UO_1734 (O_1734,N_21785,N_24011);
and UO_1735 (O_1735,N_20601,N_23941);
and UO_1736 (O_1736,N_20611,N_22255);
and UO_1737 (O_1737,N_22473,N_24897);
nand UO_1738 (O_1738,N_22295,N_22342);
or UO_1739 (O_1739,N_20416,N_24941);
nand UO_1740 (O_1740,N_20227,N_22786);
nand UO_1741 (O_1741,N_22283,N_22416);
nand UO_1742 (O_1742,N_24445,N_20752);
or UO_1743 (O_1743,N_22363,N_20987);
nor UO_1744 (O_1744,N_24304,N_21131);
nand UO_1745 (O_1745,N_24700,N_21378);
and UO_1746 (O_1746,N_23058,N_21868);
nand UO_1747 (O_1747,N_21824,N_24223);
nor UO_1748 (O_1748,N_20120,N_23813);
and UO_1749 (O_1749,N_23188,N_21822);
nor UO_1750 (O_1750,N_21059,N_21704);
nand UO_1751 (O_1751,N_24352,N_22459);
or UO_1752 (O_1752,N_22304,N_23515);
or UO_1753 (O_1753,N_21762,N_23578);
nor UO_1754 (O_1754,N_24909,N_21442);
nor UO_1755 (O_1755,N_21733,N_24350);
and UO_1756 (O_1756,N_20568,N_23298);
nand UO_1757 (O_1757,N_21906,N_21312);
nand UO_1758 (O_1758,N_21847,N_21141);
nand UO_1759 (O_1759,N_24895,N_23862);
and UO_1760 (O_1760,N_22654,N_20038);
nor UO_1761 (O_1761,N_22485,N_24060);
nand UO_1762 (O_1762,N_24234,N_24238);
nor UO_1763 (O_1763,N_24838,N_24019);
or UO_1764 (O_1764,N_20762,N_21450);
or UO_1765 (O_1765,N_20218,N_21002);
nand UO_1766 (O_1766,N_24939,N_22290);
and UO_1767 (O_1767,N_22331,N_24943);
xnor UO_1768 (O_1768,N_24721,N_20163);
and UO_1769 (O_1769,N_21316,N_21341);
nor UO_1770 (O_1770,N_23689,N_21319);
nand UO_1771 (O_1771,N_23382,N_23230);
or UO_1772 (O_1772,N_24345,N_24416);
nor UO_1773 (O_1773,N_22544,N_24258);
and UO_1774 (O_1774,N_24173,N_22270);
or UO_1775 (O_1775,N_23415,N_21046);
nand UO_1776 (O_1776,N_24955,N_24083);
or UO_1777 (O_1777,N_24062,N_22486);
nand UO_1778 (O_1778,N_20236,N_20701);
nand UO_1779 (O_1779,N_23870,N_20509);
or UO_1780 (O_1780,N_23532,N_20911);
nor UO_1781 (O_1781,N_23215,N_21501);
or UO_1782 (O_1782,N_24709,N_22957);
or UO_1783 (O_1783,N_24811,N_21590);
nor UO_1784 (O_1784,N_23242,N_21404);
and UO_1785 (O_1785,N_24052,N_24149);
and UO_1786 (O_1786,N_24960,N_23850);
or UO_1787 (O_1787,N_20333,N_23268);
and UO_1788 (O_1788,N_23950,N_21107);
nand UO_1789 (O_1789,N_21706,N_21484);
nand UO_1790 (O_1790,N_21780,N_23221);
or UO_1791 (O_1791,N_21638,N_23437);
or UO_1792 (O_1792,N_23958,N_24591);
and UO_1793 (O_1793,N_20157,N_21874);
and UO_1794 (O_1794,N_24397,N_24634);
and UO_1795 (O_1795,N_21800,N_20470);
or UO_1796 (O_1796,N_22484,N_20023);
or UO_1797 (O_1797,N_22853,N_24153);
nor UO_1798 (O_1798,N_24985,N_23334);
and UO_1799 (O_1799,N_22565,N_23457);
nand UO_1800 (O_1800,N_20135,N_21464);
or UO_1801 (O_1801,N_21700,N_22883);
xnor UO_1802 (O_1802,N_23337,N_24150);
or UO_1803 (O_1803,N_21451,N_20668);
and UO_1804 (O_1804,N_20910,N_23904);
nor UO_1805 (O_1805,N_22029,N_21166);
nand UO_1806 (O_1806,N_24663,N_22902);
nand UO_1807 (O_1807,N_23071,N_23520);
nor UO_1808 (O_1808,N_20892,N_24131);
or UO_1809 (O_1809,N_24374,N_20213);
nor UO_1810 (O_1810,N_20687,N_24080);
or UO_1811 (O_1811,N_23913,N_20739);
nor UO_1812 (O_1812,N_23686,N_23572);
and UO_1813 (O_1813,N_22759,N_20523);
nand UO_1814 (O_1814,N_20936,N_24694);
nand UO_1815 (O_1815,N_21641,N_24647);
nor UO_1816 (O_1816,N_21304,N_20215);
nor UO_1817 (O_1817,N_22538,N_23169);
or UO_1818 (O_1818,N_22947,N_24706);
nand UO_1819 (O_1819,N_20158,N_20344);
or UO_1820 (O_1820,N_22196,N_23110);
nand UO_1821 (O_1821,N_24355,N_20753);
nor UO_1822 (O_1822,N_21104,N_20350);
nand UO_1823 (O_1823,N_21367,N_22324);
or UO_1824 (O_1824,N_21017,N_20893);
nor UO_1825 (O_1825,N_23153,N_21667);
or UO_1826 (O_1826,N_23008,N_20406);
nor UO_1827 (O_1827,N_24339,N_20433);
nor UO_1828 (O_1828,N_24306,N_20223);
and UO_1829 (O_1829,N_24977,N_21353);
nor UO_1830 (O_1830,N_22686,N_23962);
or UO_1831 (O_1831,N_24208,N_23754);
nor UO_1832 (O_1832,N_21595,N_20114);
nand UO_1833 (O_1833,N_23403,N_23051);
or UO_1834 (O_1834,N_24594,N_22093);
nor UO_1835 (O_1835,N_23823,N_23343);
or UO_1836 (O_1836,N_24265,N_22197);
and UO_1837 (O_1837,N_24015,N_23447);
nand UO_1838 (O_1838,N_22289,N_22494);
nand UO_1839 (O_1839,N_21163,N_21884);
and UO_1840 (O_1840,N_24333,N_24267);
nor UO_1841 (O_1841,N_23575,N_23612);
or UO_1842 (O_1842,N_21823,N_20786);
nor UO_1843 (O_1843,N_22358,N_21445);
nand UO_1844 (O_1844,N_21541,N_22803);
or UO_1845 (O_1845,N_23971,N_21025);
xnor UO_1846 (O_1846,N_24166,N_22615);
nor UO_1847 (O_1847,N_22810,N_22507);
nor UO_1848 (O_1848,N_20165,N_20189);
nand UO_1849 (O_1849,N_21517,N_22875);
nor UO_1850 (O_1850,N_24288,N_22367);
or UO_1851 (O_1851,N_20458,N_21573);
or UO_1852 (O_1852,N_23900,N_24387);
and UO_1853 (O_1853,N_20663,N_23066);
or UO_1854 (O_1854,N_23876,N_23340);
or UO_1855 (O_1855,N_21610,N_21552);
nor UO_1856 (O_1856,N_22405,N_22487);
or UO_1857 (O_1857,N_21065,N_21210);
xor UO_1858 (O_1858,N_24662,N_20953);
and UO_1859 (O_1859,N_24199,N_24444);
nor UO_1860 (O_1860,N_22931,N_23746);
and UO_1861 (O_1861,N_22950,N_21936);
or UO_1862 (O_1862,N_20699,N_23402);
nor UO_1863 (O_1863,N_24363,N_23309);
xor UO_1864 (O_1864,N_23989,N_23681);
or UO_1865 (O_1865,N_23628,N_22533);
nand UO_1866 (O_1866,N_22998,N_22592);
and UO_1867 (O_1867,N_20408,N_23470);
or UO_1868 (O_1868,N_20604,N_24010);
nand UO_1869 (O_1869,N_21522,N_24157);
and UO_1870 (O_1870,N_21849,N_20742);
and UO_1871 (O_1871,N_22665,N_21609);
or UO_1872 (O_1872,N_23463,N_22768);
nand UO_1873 (O_1873,N_21859,N_24467);
nor UO_1874 (O_1874,N_22022,N_24095);
or UO_1875 (O_1875,N_21846,N_22188);
or UO_1876 (O_1876,N_24105,N_23728);
and UO_1877 (O_1877,N_21783,N_23693);
nor UO_1878 (O_1878,N_21931,N_23480);
nand UO_1879 (O_1879,N_20581,N_21622);
nor UO_1880 (O_1880,N_22625,N_24530);
and UO_1881 (O_1881,N_24110,N_22604);
nand UO_1882 (O_1882,N_24329,N_21693);
or UO_1883 (O_1883,N_23807,N_22073);
nand UO_1884 (O_1884,N_22986,N_21066);
and UO_1885 (O_1885,N_20554,N_23049);
nand UO_1886 (O_1886,N_24630,N_23692);
nand UO_1887 (O_1887,N_23833,N_22948);
or UO_1888 (O_1888,N_22550,N_20900);
xnor UO_1889 (O_1889,N_24420,N_23683);
or UO_1890 (O_1890,N_23449,N_20382);
and UO_1891 (O_1891,N_24532,N_20553);
nor UO_1892 (O_1892,N_24284,N_20828);
nor UO_1893 (O_1893,N_21277,N_22977);
nor UO_1894 (O_1894,N_22261,N_23715);
or UO_1895 (O_1895,N_20906,N_24422);
and UO_1896 (O_1896,N_23190,N_22499);
nor UO_1897 (O_1897,N_23423,N_20807);
or UO_1898 (O_1898,N_24729,N_24202);
and UO_1899 (O_1899,N_23623,N_24802);
nand UO_1900 (O_1900,N_20532,N_20883);
nor UO_1901 (O_1901,N_20641,N_21160);
nand UO_1902 (O_1902,N_24750,N_22558);
nor UO_1903 (O_1903,N_24713,N_22796);
and UO_1904 (O_1904,N_22981,N_24096);
and UO_1905 (O_1905,N_23043,N_24059);
nor UO_1906 (O_1906,N_20052,N_22224);
nand UO_1907 (O_1907,N_23318,N_23902);
and UO_1908 (O_1908,N_24739,N_24760);
nor UO_1909 (O_1909,N_22797,N_20393);
nand UO_1910 (O_1910,N_20045,N_21244);
nand UO_1911 (O_1911,N_21804,N_23606);
or UO_1912 (O_1912,N_20902,N_23665);
and UO_1913 (O_1913,N_23952,N_21087);
and UO_1914 (O_1914,N_22909,N_23764);
nand UO_1915 (O_1915,N_23705,N_24596);
and UO_1916 (O_1916,N_23012,N_22068);
nand UO_1917 (O_1917,N_22333,N_23443);
or UO_1918 (O_1918,N_20466,N_21043);
nand UO_1919 (O_1919,N_20511,N_23108);
or UO_1920 (O_1920,N_20123,N_20564);
xnor UO_1921 (O_1921,N_23857,N_21619);
and UO_1922 (O_1922,N_21675,N_22703);
nand UO_1923 (O_1923,N_20770,N_22034);
or UO_1924 (O_1924,N_23931,N_23645);
and UO_1925 (O_1925,N_21872,N_21564);
nor UO_1926 (O_1926,N_22234,N_22942);
and UO_1927 (O_1927,N_21336,N_24064);
nand UO_1928 (O_1928,N_23459,N_21831);
or UO_1929 (O_1929,N_21317,N_20543);
or UO_1930 (O_1930,N_21571,N_23556);
nand UO_1931 (O_1931,N_21306,N_23757);
or UO_1932 (O_1932,N_24206,N_20875);
or UO_1933 (O_1933,N_23178,N_20791);
or UO_1934 (O_1934,N_23586,N_21260);
and UO_1935 (O_1935,N_24076,N_24855);
or UO_1936 (O_1936,N_20625,N_23330);
and UO_1937 (O_1937,N_22096,N_21797);
nand UO_1938 (O_1938,N_23875,N_20761);
nor UO_1939 (O_1939,N_20263,N_24354);
nand UO_1940 (O_1940,N_23374,N_20069);
nor UO_1941 (O_1941,N_21406,N_22340);
nand UO_1942 (O_1942,N_21953,N_23198);
or UO_1943 (O_1943,N_20463,N_23405);
nand UO_1944 (O_1944,N_21686,N_21730);
nor UO_1945 (O_1945,N_21420,N_23848);
and UO_1946 (O_1946,N_21396,N_24759);
and UO_1947 (O_1947,N_20465,N_24887);
nor UO_1948 (O_1948,N_21707,N_20609);
or UO_1949 (O_1949,N_21216,N_24540);
or UO_1950 (O_1950,N_23123,N_21329);
or UO_1951 (O_1951,N_24991,N_24192);
nand UO_1952 (O_1952,N_20285,N_20093);
nor UO_1953 (O_1953,N_23772,N_21497);
nand UO_1954 (O_1954,N_21035,N_21242);
or UO_1955 (O_1955,N_20806,N_20524);
nor UO_1956 (O_1956,N_21266,N_23917);
and UO_1957 (O_1957,N_23083,N_21632);
nor UO_1958 (O_1958,N_24565,N_24403);
and UO_1959 (O_1959,N_22182,N_23685);
or UO_1960 (O_1960,N_24953,N_22585);
nor UO_1961 (O_1961,N_21978,N_23442);
nor UO_1962 (O_1962,N_22228,N_20059);
and UO_1963 (O_1963,N_20305,N_20024);
nand UO_1964 (O_1964,N_23922,N_22336);
and UO_1965 (O_1965,N_21454,N_22136);
and UO_1966 (O_1966,N_24353,N_23942);
nor UO_1967 (O_1967,N_24275,N_20537);
or UO_1968 (O_1968,N_23916,N_23314);
nor UO_1969 (O_1969,N_22823,N_24655);
nand UO_1970 (O_1970,N_21479,N_20234);
nand UO_1971 (O_1971,N_23245,N_24562);
nand UO_1972 (O_1972,N_24579,N_22530);
nor UO_1973 (O_1973,N_24341,N_20651);
nor UO_1974 (O_1974,N_23825,N_20766);
or UO_1975 (O_1975,N_24057,N_23409);
nor UO_1976 (O_1976,N_21644,N_21629);
and UO_1977 (O_1977,N_22785,N_23111);
nand UO_1978 (O_1978,N_22218,N_20569);
and UO_1979 (O_1979,N_24482,N_20424);
nor UO_1980 (O_1980,N_24319,N_21949);
nand UO_1981 (O_1981,N_20335,N_22645);
nand UO_1982 (O_1982,N_22549,N_24508);
nand UO_1983 (O_1983,N_20397,N_20566);
nor UO_1984 (O_1984,N_20781,N_20094);
and UO_1985 (O_1985,N_21628,N_22217);
nor UO_1986 (O_1986,N_20074,N_21637);
or UO_1987 (O_1987,N_20070,N_24295);
nor UO_1988 (O_1988,N_21308,N_21848);
and UO_1989 (O_1989,N_21502,N_22769);
nor UO_1990 (O_1990,N_21505,N_22139);
nand UO_1991 (O_1991,N_23930,N_20177);
and UO_1992 (O_1992,N_21648,N_22279);
nand UO_1993 (O_1993,N_22893,N_24027);
nand UO_1994 (O_1994,N_21921,N_22461);
nor UO_1995 (O_1995,N_20443,N_23186);
or UO_1996 (O_1996,N_23006,N_21159);
nand UO_1997 (O_1997,N_22418,N_21137);
or UO_1998 (O_1998,N_23625,N_23037);
nor UO_1999 (O_1999,N_20409,N_20166);
nand UO_2000 (O_2000,N_22472,N_22463);
or UO_2001 (O_2001,N_22123,N_22312);
and UO_2002 (O_2002,N_23059,N_21689);
and UO_2003 (O_2003,N_23238,N_22132);
nor UO_2004 (O_2004,N_24254,N_21740);
or UO_2005 (O_2005,N_21314,N_22954);
nor UO_2006 (O_2006,N_22498,N_21175);
and UO_2007 (O_2007,N_24612,N_22588);
nand UO_2008 (O_2008,N_20400,N_20292);
nand UO_2009 (O_2009,N_24537,N_21499);
nand UO_2010 (O_2010,N_24749,N_24506);
nand UO_2011 (O_2011,N_21873,N_23064);
or UO_2012 (O_2012,N_24077,N_20197);
and UO_2013 (O_2013,N_23643,N_23075);
nor UO_2014 (O_2014,N_23460,N_23029);
nor UO_2015 (O_2015,N_24392,N_20995);
xor UO_2016 (O_2016,N_20228,N_21188);
nand UO_2017 (O_2017,N_20749,N_24233);
nand UO_2018 (O_2018,N_20210,N_23527);
and UO_2019 (O_2019,N_20043,N_20298);
nor UO_2020 (O_2020,N_21393,N_22272);
nand UO_2021 (O_2021,N_20488,N_21945);
and UO_2022 (O_2022,N_21834,N_20760);
and UO_2023 (O_2023,N_24806,N_21206);
or UO_2024 (O_2024,N_22602,N_22930);
nor UO_2025 (O_2025,N_24757,N_24357);
xnor UO_2026 (O_2026,N_21898,N_20808);
nand UO_2027 (O_2027,N_21117,N_23555);
or UO_2028 (O_2028,N_24186,N_21692);
or UO_2029 (O_2029,N_21015,N_22043);
or UO_2030 (O_2030,N_22614,N_22387);
nor UO_2031 (O_2031,N_23903,N_24629);
and UO_2032 (O_2032,N_21913,N_22790);
and UO_2033 (O_2033,N_22811,N_21703);
and UO_2034 (O_2034,N_22206,N_20857);
and UO_2035 (O_2035,N_22557,N_23438);
nor UO_2036 (O_2036,N_22433,N_20854);
and UO_2037 (O_2037,N_21988,N_23107);
nor UO_2038 (O_2038,N_21116,N_23932);
nand UO_2039 (O_2039,N_22890,N_23963);
or UO_2040 (O_2040,N_22898,N_22837);
nand UO_2041 (O_2041,N_22249,N_21427);
nand UO_2042 (O_2042,N_23182,N_20800);
or UO_2043 (O_2043,N_24301,N_21388);
nor UO_2044 (O_2044,N_22465,N_23777);
nor UO_2045 (O_2045,N_20211,N_23792);
nand UO_2046 (O_2046,N_22708,N_23985);
nand UO_2047 (O_2047,N_22732,N_23164);
and UO_2048 (O_2048,N_21918,N_24521);
nor UO_2049 (O_2049,N_23056,N_24023);
nor UO_2050 (O_2050,N_21470,N_21683);
and UO_2051 (O_2051,N_20545,N_21618);
nor UO_2052 (O_2052,N_21249,N_20101);
nand UO_2053 (O_2053,N_20914,N_24731);
nor UO_2054 (O_2054,N_20774,N_23251);
or UO_2055 (O_2055,N_22243,N_24643);
xor UO_2056 (O_2056,N_22353,N_23323);
nand UO_2057 (O_2057,N_20015,N_22056);
and UO_2058 (O_2058,N_22303,N_24645);
and UO_2059 (O_2059,N_23512,N_20422);
nand UO_2060 (O_2060,N_24705,N_20267);
nor UO_2061 (O_2061,N_20291,N_21943);
and UO_2062 (O_2062,N_23923,N_20171);
and UO_2063 (O_2063,N_20084,N_22970);
nand UO_2064 (O_2064,N_23735,N_24781);
nor UO_2065 (O_2065,N_24894,N_22440);
and UO_2066 (O_2066,N_23475,N_24919);
nand UO_2067 (O_2067,N_21360,N_22589);
nor UO_2068 (O_2068,N_22685,N_21990);
nor UO_2069 (O_2069,N_22020,N_22961);
nand UO_2070 (O_2070,N_22120,N_24321);
and UO_2071 (O_2071,N_22256,N_22121);
and UO_2072 (O_2072,N_22518,N_24528);
nand UO_2073 (O_2073,N_22309,N_20012);
nand UO_2074 (O_2074,N_22010,N_21296);
and UO_2075 (O_2075,N_22403,N_23302);
nand UO_2076 (O_2076,N_21431,N_23598);
nand UO_2077 (O_2077,N_20587,N_21000);
nand UO_2078 (O_2078,N_24201,N_21069);
xnor UO_2079 (O_2079,N_21958,N_22054);
and UO_2080 (O_2080,N_20924,N_21003);
nand UO_2081 (O_2081,N_20855,N_21956);
nand UO_2082 (O_2082,N_24429,N_20073);
nor UO_2083 (O_2083,N_23019,N_21436);
or UO_2084 (O_2084,N_23349,N_20030);
and UO_2085 (O_2085,N_20450,N_21746);
nor UO_2086 (O_2086,N_21088,N_21148);
and UO_2087 (O_2087,N_24631,N_22846);
and UO_2088 (O_2088,N_21363,N_23956);
nor UO_2089 (O_2089,N_20247,N_20150);
and UO_2090 (O_2090,N_20799,N_21491);
nor UO_2091 (O_2091,N_20997,N_23398);
nor UO_2092 (O_2092,N_24726,N_24185);
and UO_2093 (O_2093,N_20942,N_23656);
nor UO_2094 (O_2094,N_21014,N_23132);
nor UO_2095 (O_2095,N_20825,N_22935);
nor UO_2096 (O_2096,N_22847,N_20173);
nor UO_2097 (O_2097,N_24293,N_23719);
and UO_2098 (O_2098,N_23854,N_22660);
nor UO_2099 (O_2099,N_23687,N_23600);
xnor UO_2100 (O_2100,N_22515,N_24605);
or UO_2101 (O_2101,N_23036,N_24531);
xor UO_2102 (O_2102,N_23265,N_24868);
nor UO_2103 (O_2103,N_23991,N_21201);
nor UO_2104 (O_2104,N_22128,N_23987);
or UO_2105 (O_2105,N_24724,N_21303);
and UO_2106 (O_2106,N_24614,N_20250);
nor UO_2107 (O_2107,N_20474,N_22833);
nor UO_2108 (O_2108,N_22644,N_24001);
nand UO_2109 (O_2109,N_21582,N_20268);
nor UO_2110 (O_2110,N_24584,N_24443);
and UO_2111 (O_2111,N_23573,N_20738);
xnor UO_2112 (O_2112,N_21208,N_23773);
nand UO_2113 (O_2113,N_23201,N_21067);
xor UO_2114 (O_2114,N_22241,N_24711);
and UO_2115 (O_2115,N_20928,N_20575);
and UO_2116 (O_2116,N_22392,N_24447);
nand UO_2117 (O_2117,N_23327,N_20820);
or UO_2118 (O_2118,N_20201,N_23889);
nand UO_2119 (O_2119,N_20067,N_20219);
nand UO_2120 (O_2120,N_21579,N_21653);
nand UO_2121 (O_2121,N_21982,N_22882);
and UO_2122 (O_2122,N_24382,N_21920);
and UO_2123 (O_2123,N_21526,N_22994);
or UO_2124 (O_2124,N_21247,N_21315);
and UO_2125 (O_2125,N_24896,N_22077);
and UO_2126 (O_2126,N_21310,N_22057);
nand UO_2127 (O_2127,N_23560,N_24326);
or UO_2128 (O_2128,N_23304,N_21597);
or UO_2129 (O_2129,N_20679,N_23213);
nor UO_2130 (O_2130,N_23832,N_22915);
nor UO_2131 (O_2131,N_20918,N_23821);
nand UO_2132 (O_2132,N_20004,N_23355);
nor UO_2133 (O_2133,N_24654,N_21153);
or UO_2134 (O_2134,N_24449,N_23356);
nor UO_2135 (O_2135,N_20720,N_21217);
or UO_2136 (O_2136,N_20644,N_21352);
nand UO_2137 (O_2137,N_22656,N_23841);
or UO_2138 (O_2138,N_21919,N_20725);
nand UO_2139 (O_2139,N_23827,N_22501);
and UO_2140 (O_2140,N_22664,N_23800);
or UO_2141 (O_2141,N_22207,N_20961);
and UO_2142 (O_2142,N_22584,N_21468);
and UO_2143 (O_2143,N_22391,N_22209);
nand UO_2144 (O_2144,N_24217,N_20384);
or UO_2145 (O_2145,N_22427,N_22099);
nor UO_2146 (O_2146,N_20711,N_24270);
and UO_2147 (O_2147,N_22171,N_20674);
nand UO_2148 (O_2148,N_20077,N_22411);
and UO_2149 (O_2149,N_22031,N_23416);
xnor UO_2150 (O_2150,N_23278,N_23207);
and UO_2151 (O_2151,N_21592,N_23938);
and UO_2152 (O_2152,N_21376,N_23607);
and UO_2153 (O_2153,N_21362,N_20667);
and UO_2154 (O_2154,N_22626,N_22019);
or UO_2155 (O_2155,N_21365,N_22666);
and UO_2156 (O_2156,N_21253,N_22789);
or UO_2157 (O_2157,N_22161,N_20300);
and UO_2158 (O_2158,N_22647,N_21113);
nor UO_2159 (O_2159,N_23980,N_20169);
or UO_2160 (O_2160,N_24842,N_23120);
nand UO_2161 (O_2161,N_23852,N_24143);
and UO_2162 (O_2162,N_24888,N_20967);
and UO_2163 (O_2163,N_20246,N_20811);
or UO_2164 (O_2164,N_21264,N_20149);
nand UO_2165 (O_2165,N_24239,N_23401);
nor UO_2166 (O_2166,N_24576,N_20897);
or UO_2167 (O_2167,N_20640,N_24134);
xnor UO_2168 (O_2168,N_24847,N_22715);
or UO_2169 (O_2169,N_23241,N_24071);
nand UO_2170 (O_2170,N_24401,N_20971);
nor UO_2171 (O_2171,N_21462,N_23489);
nand UO_2172 (O_2172,N_23226,N_21039);
or UO_2173 (O_2173,N_23933,N_24674);
nor UO_2174 (O_2174,N_21727,N_24476);
or UO_2175 (O_2175,N_24056,N_24921);
nand UO_2176 (O_2176,N_24585,N_23116);
or UO_2177 (O_2177,N_24191,N_23099);
and UO_2178 (O_2178,N_22059,N_22110);
nand UO_2179 (O_2179,N_22876,N_22293);
and UO_2180 (O_2180,N_24918,N_24648);
nor UO_2181 (O_2181,N_20280,N_20000);
or UO_2182 (O_2182,N_24945,N_24769);
nor UO_2183 (O_2183,N_22105,N_20402);
nand UO_2184 (O_2184,N_23073,N_23888);
and UO_2185 (O_2185,N_22740,N_23021);
nand UO_2186 (O_2186,N_24768,N_21147);
nand UO_2187 (O_2187,N_23637,N_24346);
or UO_2188 (O_2188,N_24672,N_21565);
and UO_2189 (O_2189,N_21662,N_23171);
nand UO_2190 (O_2190,N_24976,N_20325);
nor UO_2191 (O_2191,N_23389,N_24828);
and UO_2192 (O_2192,N_22669,N_24786);
and UO_2193 (O_2193,N_23752,N_21299);
nor UO_2194 (O_2194,N_20222,N_24232);
and UO_2195 (O_2195,N_21110,N_20471);
or UO_2196 (O_2196,N_24753,N_24043);
nand UO_2197 (O_2197,N_22758,N_22993);
nor UO_2198 (O_2198,N_20146,N_22298);
nand UO_2199 (O_2199,N_22979,N_22344);
or UO_2200 (O_2200,N_20010,N_24801);
nor UO_2201 (O_2201,N_20342,N_22571);
or UO_2202 (O_2202,N_20949,N_20404);
or UO_2203 (O_2203,N_20541,N_22506);
nor UO_2204 (O_2204,N_23896,N_20878);
and UO_2205 (O_2205,N_21537,N_22027);
nor UO_2206 (O_2206,N_20096,N_20235);
or UO_2207 (O_2207,N_22707,N_22971);
and UO_2208 (O_2208,N_22420,N_22447);
or UO_2209 (O_2209,N_20339,N_20383);
nand UO_2210 (O_2210,N_23784,N_23414);
xnor UO_2211 (O_2211,N_21456,N_23824);
nand UO_2212 (O_2212,N_22086,N_22238);
nor UO_2213 (O_2213,N_21440,N_20615);
nor UO_2214 (O_2214,N_24740,N_22094);
xnor UO_2215 (O_2215,N_22918,N_20496);
xor UO_2216 (O_2216,N_21064,N_24462);
nand UO_2217 (O_2217,N_20927,N_21709);
nor UO_2218 (O_2218,N_20617,N_22329);
nor UO_2219 (O_2219,N_24845,N_22904);
nor UO_2220 (O_2220,N_22808,N_20534);
nor UO_2221 (O_2221,N_24298,N_20864);
xnor UO_2222 (O_2222,N_23812,N_22021);
nor UO_2223 (O_2223,N_23434,N_23957);
nand UO_2224 (O_2224,N_20934,N_23517);
nor UO_2225 (O_2225,N_21759,N_23220);
or UO_2226 (O_2226,N_23428,N_24228);
and UO_2227 (O_2227,N_23426,N_24453);
nor UO_2228 (O_2228,N_24314,N_23965);
and UO_2229 (O_2229,N_20628,N_24533);
or UO_2230 (O_2230,N_24046,N_20132);
nor UO_2231 (O_2231,N_22474,N_23432);
nor UO_2232 (O_2232,N_20719,N_23379);
and UO_2233 (O_2233,N_23163,N_24851);
and UO_2234 (O_2234,N_20357,N_22567);
nor UO_2235 (O_2235,N_24567,N_23726);
or UO_2236 (O_2236,N_21164,N_23704);
and UO_2237 (O_2237,N_21326,N_21033);
nor UO_2238 (O_2238,N_20962,N_24193);
nor UO_2239 (O_2239,N_24399,N_24091);
nand UO_2240 (O_2240,N_20845,N_20480);
and UO_2241 (O_2241,N_23767,N_21546);
nand UO_2242 (O_2242,N_24983,N_22825);
or UO_2243 (O_2243,N_24475,N_20512);
nor UO_2244 (O_2244,N_24009,N_20499);
and UO_2245 (O_2245,N_24221,N_23079);
nor UO_2246 (O_2246,N_23234,N_23487);
and UO_2247 (O_2247,N_21441,N_21669);
nor UO_2248 (O_2248,N_23604,N_22606);
nor UO_2249 (O_2249,N_22941,N_24085);
or UO_2250 (O_2250,N_22519,N_21202);
or UO_2251 (O_2251,N_20849,N_20620);
and UO_2252 (O_2252,N_21384,N_22964);
nor UO_2253 (O_2253,N_20327,N_24682);
nor UO_2254 (O_2254,N_21461,N_20319);
nand UO_2255 (O_2255,N_23179,N_22173);
or UO_2256 (O_2256,N_23722,N_23490);
nor UO_2257 (O_2257,N_22661,N_21658);
and UO_2258 (O_2258,N_24360,N_24763);
nand UO_2259 (O_2259,N_22932,N_23514);
nand UO_2260 (O_2260,N_21659,N_21513);
xor UO_2261 (O_2261,N_23817,N_22526);
or UO_2262 (O_2262,N_24774,N_23631);
or UO_2263 (O_2263,N_24815,N_20314);
nand UO_2264 (O_2264,N_23326,N_24610);
nand UO_2265 (O_2265,N_21151,N_21510);
and UO_2266 (O_2266,N_21642,N_24984);
or UO_2267 (O_2267,N_20492,N_24730);
nand UO_2268 (O_2268,N_22520,N_21134);
and UO_2269 (O_2269,N_24243,N_24962);
nor UO_2270 (O_2270,N_21694,N_24490);
nand UO_2271 (O_2271,N_20666,N_24556);
or UO_2272 (O_2272,N_22058,N_21811);
nor UO_2273 (O_2273,N_23634,N_20623);
xnor UO_2274 (O_2274,N_20274,N_20204);
and UO_2275 (O_2275,N_21108,N_24320);
nand UO_2276 (O_2276,N_22200,N_22952);
nor UO_2277 (O_2277,N_24415,N_21935);
xnor UO_2278 (O_2278,N_24033,N_24287);
nand UO_2279 (O_2279,N_22425,N_21267);
and UO_2280 (O_2280,N_21234,N_22735);
and UO_2281 (O_2281,N_24572,N_23666);
or UO_2282 (O_2282,N_23458,N_23608);
nand UO_2283 (O_2283,N_22745,N_22175);
nand UO_2284 (O_2284,N_22004,N_24002);
nor UO_2285 (O_2285,N_23420,N_24871);
nand UO_2286 (O_2286,N_23741,N_23418);
nand UO_2287 (O_2287,N_21791,N_23497);
nor UO_2288 (O_2288,N_20001,N_24207);
or UO_2289 (O_2289,N_20755,N_20164);
nand UO_2290 (O_2290,N_24455,N_24047);
nand UO_2291 (O_2291,N_21757,N_20985);
and UO_2292 (O_2292,N_20964,N_24151);
nor UO_2293 (O_2293,N_20358,N_22297);
or UO_2294 (O_2294,N_20138,N_22496);
nor UO_2295 (O_2295,N_24902,N_23204);
nor UO_2296 (O_2296,N_22741,N_22423);
or UO_2297 (O_2297,N_24965,N_24437);
nor UO_2298 (O_2298,N_20583,N_23559);
nor UO_2299 (O_2299,N_23225,N_24381);
nor UO_2300 (O_2300,N_23504,N_21539);
and UO_2301 (O_2301,N_20061,N_22608);
and UO_2302 (O_2302,N_24872,N_20598);
nand UO_2303 (O_2303,N_24302,N_20652);
xor UO_2304 (O_2304,N_20255,N_20932);
or UO_2305 (O_2305,N_22674,N_23732);
and UO_2306 (O_2306,N_24152,N_22366);
and UO_2307 (O_2307,N_21426,N_20110);
and UO_2308 (O_2308,N_22446,N_23353);
or UO_2309 (O_2309,N_22555,N_24116);
nand UO_2310 (O_2310,N_22193,N_20919);
nor UO_2311 (O_2311,N_23276,N_20558);
nand UO_2312 (O_2312,N_20143,N_24542);
and UO_2313 (O_2313,N_24959,N_21651);
nand UO_2314 (O_2314,N_23354,N_21777);
or UO_2315 (O_2315,N_23945,N_24404);
nor UO_2316 (O_2316,N_23084,N_24973);
or UO_2317 (O_2317,N_24348,N_24874);
nand UO_2318 (O_2318,N_22202,N_20968);
nand UO_2319 (O_2319,N_23542,N_20087);
xnor UO_2320 (O_2320,N_24864,N_20140);
nand UO_2321 (O_2321,N_20129,N_22183);
nand UO_2322 (O_2322,N_20375,N_23791);
or UO_2323 (O_2323,N_22820,N_20348);
nand UO_2324 (O_2324,N_20735,N_24040);
nand UO_2325 (O_2325,N_24678,N_21081);
nor UO_2326 (O_2326,N_24578,N_24478);
and UO_2327 (O_2327,N_24604,N_22754);
or UO_2328 (O_2328,N_24248,N_20279);
or UO_2329 (O_2329,N_23947,N_24396);
xor UO_2330 (O_2330,N_24693,N_20717);
nand UO_2331 (O_2331,N_21842,N_21128);
nand UO_2332 (O_2332,N_21492,N_22988);
or UO_2333 (O_2333,N_23417,N_22788);
and UO_2334 (O_2334,N_20940,N_24170);
nand UO_2335 (O_2335,N_21585,N_20678);
nor UO_2336 (O_2336,N_22286,N_24504);
xor UO_2337 (O_2337,N_24744,N_23456);
and UO_2338 (O_2338,N_20947,N_21139);
nand UO_2339 (O_2339,N_23718,N_21705);
and UO_2340 (O_2340,N_23579,N_21545);
nand UO_2341 (O_2341,N_20655,N_21570);
nor UO_2342 (O_2342,N_20420,N_22167);
nand UO_2343 (O_2343,N_22944,N_24251);
and UO_2344 (O_2344,N_23696,N_23072);
and UO_2345 (O_2345,N_22545,N_23847);
nand UO_2346 (O_2346,N_20194,N_22884);
nor UO_2347 (O_2347,N_20673,N_23695);
nand UO_2348 (O_2348,N_20946,N_21807);
nor UO_2349 (O_2349,N_22556,N_22662);
or UO_2350 (O_2350,N_24701,N_23257);
xor UO_2351 (O_2351,N_21551,N_20672);
nor UO_2352 (O_2352,N_20425,N_23673);
nand UO_2353 (O_2353,N_24910,N_22483);
or UO_2354 (O_2354,N_20009,N_23694);
or UO_2355 (O_2355,N_21130,N_23103);
xor UO_2356 (O_2356,N_22095,N_22490);
nor UO_2357 (O_2357,N_21076,N_21084);
or UO_2358 (O_2358,N_20440,N_21126);
nor UO_2359 (O_2359,N_24367,N_24805);
or UO_2360 (O_2360,N_22143,N_20832);
or UO_2361 (O_2361,N_21135,N_23994);
nor UO_2362 (O_2362,N_24088,N_23233);
and UO_2363 (O_2363,N_22633,N_22869);
nor UO_2364 (O_2364,N_24837,N_21549);
nor UO_2365 (O_2365,N_24978,N_21096);
and UO_2366 (O_2366,N_23988,N_24748);
nand UO_2367 (O_2367,N_21550,N_20771);
nor UO_2368 (O_2368,N_24031,N_23044);
and UO_2369 (O_2369,N_24905,N_22407);
nor UO_2370 (O_2370,N_24276,N_23802);
xnor UO_2371 (O_2371,N_21102,N_22378);
nor UO_2372 (O_2372,N_22738,N_22341);
and UO_2373 (O_2373,N_24045,N_23795);
nor UO_2374 (O_2374,N_22168,N_20216);
xnor UO_2375 (O_2375,N_23422,N_20371);
nor UO_2376 (O_2376,N_23529,N_20861);
and UO_2377 (O_2377,N_23676,N_22417);
and UO_2378 (O_2378,N_22404,N_20908);
nand UO_2379 (O_2379,N_22449,N_21313);
and UO_2380 (O_2380,N_22164,N_21952);
or UO_2381 (O_2381,N_20899,N_21838);
and UO_2382 (O_2382,N_20359,N_22266);
or UO_2383 (O_2383,N_21878,N_22610);
nor UO_2384 (O_2384,N_24925,N_23119);
nor UO_2385 (O_2385,N_23047,N_20326);
nor UO_2386 (O_2386,N_24616,N_24078);
or UO_2387 (O_2387,N_21864,N_22337);
nor UO_2388 (O_2388,N_20660,N_24257);
nor UO_2389 (O_2389,N_20639,N_20082);
or UO_2390 (O_2390,N_22402,N_24008);
nand UO_2391 (O_2391,N_20647,N_23114);
or UO_2392 (O_2392,N_21186,N_21459);
nand UO_2393 (O_2393,N_24277,N_24484);
nand UO_2394 (O_2394,N_24972,N_20193);
and UO_2395 (O_2395,N_23156,N_20741);
nor UO_2396 (O_2396,N_20698,N_24212);
or UO_2397 (O_2397,N_22778,N_20320);
and UO_2398 (O_2398,N_22221,N_24450);
xnor UO_2399 (O_2399,N_24117,N_22129);
nand UO_2400 (O_2400,N_20515,N_24625);
or UO_2401 (O_2401,N_22657,N_21711);
and UO_2402 (O_2402,N_23702,N_22593);
and UO_2403 (O_2403,N_20468,N_24142);
nand UO_2404 (O_2404,N_23733,N_22430);
and UO_2405 (O_2405,N_22441,N_24466);
and UO_2406 (O_2406,N_24456,N_23878);
or UO_2407 (O_2407,N_20377,N_21713);
or UO_2408 (O_2408,N_21075,N_21152);
or UO_2409 (O_2409,N_22025,N_20429);
nand UO_2410 (O_2410,N_23052,N_22045);
nor UO_2411 (O_2411,N_20595,N_20063);
and UO_2412 (O_2412,N_20368,N_22525);
nand UO_2413 (O_2413,N_23557,N_20694);
nor UO_2414 (O_2414,N_22975,N_24555);
nand UO_2415 (O_2415,N_23819,N_21830);
and UO_2416 (O_2416,N_22165,N_21185);
xnor UO_2417 (O_2417,N_24146,N_23136);
and UO_2418 (O_2418,N_23368,N_20461);
and UO_2419 (O_2419,N_21305,N_23564);
and UO_2420 (O_2420,N_21716,N_22691);
or UO_2421 (O_2421,N_23894,N_24100);
nor UO_2422 (O_2422,N_20682,N_22305);
or UO_2423 (O_2423,N_22747,N_24496);
nor UO_2424 (O_2424,N_20269,N_22635);
nand UO_2425 (O_2425,N_21387,N_21856);
nor UO_2426 (O_2426,N_21473,N_22991);
or UO_2427 (O_2427,N_22650,N_24268);
and UO_2428 (O_2428,N_20494,N_20054);
or UO_2429 (O_2429,N_20726,N_20510);
nand UO_2430 (O_2430,N_20062,N_23390);
nand UO_2431 (O_2431,N_20917,N_20317);
or UO_2432 (O_2432,N_20386,N_22807);
or UO_2433 (O_2433,N_21328,N_22098);
and UO_2434 (O_2434,N_20905,N_22085);
and UO_2435 (O_2435,N_22834,N_24692);
or UO_2436 (O_2436,N_23092,N_22505);
nor UO_2437 (O_2437,N_24358,N_20856);
or UO_2438 (O_2438,N_23212,N_20331);
xor UO_2439 (O_2439,N_20258,N_22375);
nor UO_2440 (O_2440,N_20814,N_20850);
nand UO_2441 (O_2441,N_23639,N_24893);
nand UO_2442 (O_2442,N_22627,N_21984);
nand UO_2443 (O_2443,N_24906,N_22659);
nor UO_2444 (O_2444,N_20610,N_20217);
xnor UO_2445 (O_2445,N_22489,N_23999);
nand UO_2446 (O_2446,N_20185,N_20731);
or UO_2447 (O_2447,N_22162,N_21386);
nand UO_2448 (O_2448,N_22248,N_20790);
or UO_2449 (O_2449,N_24599,N_24042);
or UO_2450 (O_2450,N_23590,N_21407);
and UO_2451 (O_2451,N_24189,N_23535);
and UO_2452 (O_2452,N_20685,N_23668);
and UO_2453 (O_2453,N_24914,N_20395);
or UO_2454 (O_2454,N_21095,N_23826);
and UO_2455 (O_2455,N_22907,N_24371);
or UO_2456 (O_2456,N_23093,N_22230);
or UO_2457 (O_2457,N_21149,N_23055);
or UO_2458 (O_2458,N_21645,N_24582);
or UO_2459 (O_2459,N_24541,N_22479);
and UO_2460 (O_2460,N_23376,N_20261);
nand UO_2461 (O_2461,N_20637,N_21802);
nor UO_2462 (O_2462,N_23258,N_21424);
or UO_2463 (O_2463,N_20407,N_20612);
nand UO_2464 (O_2464,N_23407,N_22596);
or UO_2465 (O_2465,N_20925,N_21063);
and UO_2466 (O_2466,N_23203,N_20943);
and UO_2467 (O_2467,N_23869,N_24831);
nand UO_2468 (O_2468,N_23341,N_24197);
or UO_2469 (O_2469,N_24829,N_24883);
xor UO_2470 (O_2470,N_22874,N_22470);
and UO_2471 (O_2471,N_22287,N_21401);
nor UO_2472 (O_2472,N_24968,N_21825);
nor UO_2473 (O_2473,N_20168,N_22663);
or UO_2474 (O_2474,N_22362,N_22064);
or UO_2475 (O_2475,N_24364,N_24642);
or UO_2476 (O_2476,N_21391,N_24227);
nand UO_2477 (O_2477,N_24650,N_20759);
or UO_2478 (O_2478,N_23836,N_22636);
or UO_2479 (O_2479,N_20966,N_21068);
or UO_2480 (O_2480,N_24559,N_23160);
nor UO_2481 (O_2481,N_23954,N_24376);
or UO_2482 (O_2482,N_24097,N_20830);
nand UO_2483 (O_2483,N_20539,N_20833);
nor UO_2484 (O_2484,N_22563,N_22868);
nor UO_2485 (O_2485,N_22854,N_22672);
and UO_2486 (O_2486,N_23771,N_23360);
nor UO_2487 (O_2487,N_24424,N_20704);
or UO_2488 (O_2488,N_24250,N_24966);
nor UO_2489 (O_2489,N_24127,N_20696);
or UO_2490 (O_2490,N_24006,N_20992);
and UO_2491 (O_2491,N_21599,N_23893);
and UO_2492 (O_2492,N_24557,N_22377);
and UO_2493 (O_2493,N_20195,N_21125);
nand UO_2494 (O_2494,N_20019,N_21684);
nor UO_2495 (O_2495,N_23478,N_24588);
and UO_2496 (O_2496,N_20418,N_23467);
or UO_2497 (O_2497,N_24778,N_23023);
and UO_2498 (O_2498,N_24641,N_21972);
nand UO_2499 (O_2499,N_24086,N_24553);
or UO_2500 (O_2500,N_20931,N_21540);
and UO_2501 (O_2501,N_22437,N_22832);
or UO_2502 (O_2502,N_22104,N_20884);
and UO_2503 (O_2503,N_24980,N_21002);
or UO_2504 (O_2504,N_20161,N_22961);
or UO_2505 (O_2505,N_20041,N_20710);
and UO_2506 (O_2506,N_22889,N_23448);
nor UO_2507 (O_2507,N_24626,N_20909);
nand UO_2508 (O_2508,N_21090,N_20208);
or UO_2509 (O_2509,N_21045,N_23585);
nand UO_2510 (O_2510,N_22461,N_21303);
and UO_2511 (O_2511,N_20656,N_22765);
or UO_2512 (O_2512,N_20661,N_24235);
nand UO_2513 (O_2513,N_22880,N_24086);
nand UO_2514 (O_2514,N_22925,N_22473);
nor UO_2515 (O_2515,N_20070,N_22233);
or UO_2516 (O_2516,N_20053,N_24892);
or UO_2517 (O_2517,N_21593,N_21873);
and UO_2518 (O_2518,N_23326,N_22583);
and UO_2519 (O_2519,N_22328,N_22363);
nor UO_2520 (O_2520,N_22191,N_20165);
nand UO_2521 (O_2521,N_21129,N_23693);
nand UO_2522 (O_2522,N_20599,N_21173);
or UO_2523 (O_2523,N_23718,N_20988);
nand UO_2524 (O_2524,N_23676,N_20106);
nand UO_2525 (O_2525,N_23960,N_21144);
nand UO_2526 (O_2526,N_24702,N_21693);
nand UO_2527 (O_2527,N_22338,N_24307);
nor UO_2528 (O_2528,N_20715,N_20546);
nor UO_2529 (O_2529,N_20558,N_22126);
or UO_2530 (O_2530,N_21431,N_24892);
nand UO_2531 (O_2531,N_20459,N_24093);
nand UO_2532 (O_2532,N_20613,N_23291);
and UO_2533 (O_2533,N_23908,N_22173);
nor UO_2534 (O_2534,N_21019,N_21660);
nor UO_2535 (O_2535,N_24537,N_22280);
nor UO_2536 (O_2536,N_23061,N_23421);
and UO_2537 (O_2537,N_24346,N_20547);
nor UO_2538 (O_2538,N_23186,N_23769);
or UO_2539 (O_2539,N_24260,N_23172);
or UO_2540 (O_2540,N_20049,N_21632);
and UO_2541 (O_2541,N_23264,N_22551);
nor UO_2542 (O_2542,N_21424,N_21998);
and UO_2543 (O_2543,N_20799,N_23129);
and UO_2544 (O_2544,N_24522,N_20506);
and UO_2545 (O_2545,N_22557,N_20955);
and UO_2546 (O_2546,N_21989,N_21416);
and UO_2547 (O_2547,N_20467,N_22844);
or UO_2548 (O_2548,N_22021,N_20895);
and UO_2549 (O_2549,N_22234,N_21036);
and UO_2550 (O_2550,N_20027,N_21842);
nor UO_2551 (O_2551,N_20263,N_23614);
and UO_2552 (O_2552,N_21481,N_24371);
or UO_2553 (O_2553,N_20920,N_21665);
or UO_2554 (O_2554,N_24067,N_20383);
nand UO_2555 (O_2555,N_24253,N_22160);
and UO_2556 (O_2556,N_23186,N_23773);
xnor UO_2557 (O_2557,N_23638,N_23912);
and UO_2558 (O_2558,N_21707,N_22708);
nand UO_2559 (O_2559,N_24658,N_24544);
or UO_2560 (O_2560,N_22216,N_20413);
nand UO_2561 (O_2561,N_21251,N_20378);
nand UO_2562 (O_2562,N_20025,N_21557);
nor UO_2563 (O_2563,N_21178,N_23411);
and UO_2564 (O_2564,N_20483,N_21995);
nor UO_2565 (O_2565,N_21023,N_22495);
and UO_2566 (O_2566,N_23754,N_22785);
xor UO_2567 (O_2567,N_20573,N_20858);
and UO_2568 (O_2568,N_23201,N_24009);
or UO_2569 (O_2569,N_20434,N_20204);
or UO_2570 (O_2570,N_20762,N_21940);
or UO_2571 (O_2571,N_20429,N_23477);
nor UO_2572 (O_2572,N_22233,N_23537);
nor UO_2573 (O_2573,N_20906,N_21479);
and UO_2574 (O_2574,N_20589,N_20998);
nand UO_2575 (O_2575,N_23414,N_23662);
nand UO_2576 (O_2576,N_24201,N_22318);
nor UO_2577 (O_2577,N_23002,N_23805);
xor UO_2578 (O_2578,N_20014,N_22407);
or UO_2579 (O_2579,N_24963,N_21938);
and UO_2580 (O_2580,N_20404,N_24349);
nor UO_2581 (O_2581,N_20529,N_21256);
nor UO_2582 (O_2582,N_22283,N_21472);
and UO_2583 (O_2583,N_21418,N_20900);
nor UO_2584 (O_2584,N_22211,N_21239);
or UO_2585 (O_2585,N_22080,N_20444);
or UO_2586 (O_2586,N_21870,N_23915);
nand UO_2587 (O_2587,N_24628,N_21896);
or UO_2588 (O_2588,N_21609,N_24160);
nor UO_2589 (O_2589,N_22787,N_22329);
nor UO_2590 (O_2590,N_23962,N_24311);
or UO_2591 (O_2591,N_23323,N_21726);
and UO_2592 (O_2592,N_23593,N_23974);
or UO_2593 (O_2593,N_20057,N_21867);
nor UO_2594 (O_2594,N_20080,N_23590);
and UO_2595 (O_2595,N_20281,N_23487);
xor UO_2596 (O_2596,N_23425,N_23006);
nor UO_2597 (O_2597,N_21895,N_24633);
and UO_2598 (O_2598,N_21154,N_21444);
and UO_2599 (O_2599,N_24055,N_23377);
and UO_2600 (O_2600,N_21653,N_23427);
nand UO_2601 (O_2601,N_23951,N_24914);
nor UO_2602 (O_2602,N_21738,N_20781);
or UO_2603 (O_2603,N_23103,N_20185);
nor UO_2604 (O_2604,N_23402,N_23746);
nor UO_2605 (O_2605,N_24179,N_24982);
nor UO_2606 (O_2606,N_23856,N_20380);
and UO_2607 (O_2607,N_23721,N_22380);
or UO_2608 (O_2608,N_21648,N_21523);
and UO_2609 (O_2609,N_22271,N_21125);
or UO_2610 (O_2610,N_24901,N_20750);
and UO_2611 (O_2611,N_24305,N_21670);
nor UO_2612 (O_2612,N_22564,N_21681);
nand UO_2613 (O_2613,N_21685,N_20180);
and UO_2614 (O_2614,N_21134,N_23498);
nand UO_2615 (O_2615,N_21608,N_20824);
nor UO_2616 (O_2616,N_21537,N_20677);
or UO_2617 (O_2617,N_24750,N_23754);
and UO_2618 (O_2618,N_24073,N_22630);
nor UO_2619 (O_2619,N_21950,N_21761);
or UO_2620 (O_2620,N_21095,N_23596);
nand UO_2621 (O_2621,N_22233,N_24798);
nand UO_2622 (O_2622,N_23611,N_20056);
nor UO_2623 (O_2623,N_23822,N_21395);
nand UO_2624 (O_2624,N_22594,N_24400);
or UO_2625 (O_2625,N_22803,N_23841);
nand UO_2626 (O_2626,N_23036,N_22787);
nor UO_2627 (O_2627,N_23991,N_23769);
or UO_2628 (O_2628,N_22447,N_21207);
and UO_2629 (O_2629,N_24257,N_22249);
xnor UO_2630 (O_2630,N_22510,N_24993);
nand UO_2631 (O_2631,N_20157,N_22007);
nand UO_2632 (O_2632,N_23890,N_24084);
and UO_2633 (O_2633,N_23909,N_23841);
or UO_2634 (O_2634,N_20243,N_23115);
nand UO_2635 (O_2635,N_20129,N_21577);
nor UO_2636 (O_2636,N_24601,N_23927);
and UO_2637 (O_2637,N_24902,N_21630);
and UO_2638 (O_2638,N_24308,N_20967);
nor UO_2639 (O_2639,N_24829,N_21586);
or UO_2640 (O_2640,N_22500,N_21900);
nand UO_2641 (O_2641,N_22553,N_20156);
and UO_2642 (O_2642,N_24838,N_23512);
nand UO_2643 (O_2643,N_20694,N_24178);
or UO_2644 (O_2644,N_22577,N_24883);
nand UO_2645 (O_2645,N_20378,N_22087);
and UO_2646 (O_2646,N_24247,N_24217);
nor UO_2647 (O_2647,N_24052,N_22065);
nand UO_2648 (O_2648,N_24749,N_22105);
nor UO_2649 (O_2649,N_20368,N_22549);
or UO_2650 (O_2650,N_24300,N_23285);
or UO_2651 (O_2651,N_22599,N_23885);
or UO_2652 (O_2652,N_24504,N_20441);
or UO_2653 (O_2653,N_22429,N_23128);
or UO_2654 (O_2654,N_21804,N_23673);
or UO_2655 (O_2655,N_20376,N_21695);
or UO_2656 (O_2656,N_23984,N_22552);
xnor UO_2657 (O_2657,N_20567,N_24752);
and UO_2658 (O_2658,N_24204,N_22158);
and UO_2659 (O_2659,N_22760,N_23259);
nand UO_2660 (O_2660,N_24984,N_22783);
or UO_2661 (O_2661,N_23789,N_22771);
and UO_2662 (O_2662,N_22614,N_23406);
and UO_2663 (O_2663,N_24188,N_21166);
nor UO_2664 (O_2664,N_20407,N_24852);
nor UO_2665 (O_2665,N_21489,N_24486);
and UO_2666 (O_2666,N_20054,N_23982);
or UO_2667 (O_2667,N_24947,N_22542);
and UO_2668 (O_2668,N_21664,N_22872);
or UO_2669 (O_2669,N_22936,N_20664);
or UO_2670 (O_2670,N_22296,N_24284);
and UO_2671 (O_2671,N_21663,N_23297);
nor UO_2672 (O_2672,N_20307,N_21621);
and UO_2673 (O_2673,N_22081,N_22735);
and UO_2674 (O_2674,N_20207,N_22633);
nor UO_2675 (O_2675,N_22314,N_23411);
and UO_2676 (O_2676,N_23307,N_23022);
nand UO_2677 (O_2677,N_24386,N_24145);
nor UO_2678 (O_2678,N_23766,N_22812);
nand UO_2679 (O_2679,N_23773,N_23352);
nand UO_2680 (O_2680,N_24149,N_22753);
or UO_2681 (O_2681,N_24346,N_24930);
nor UO_2682 (O_2682,N_24825,N_24920);
xnor UO_2683 (O_2683,N_21530,N_24439);
and UO_2684 (O_2684,N_22395,N_21475);
nand UO_2685 (O_2685,N_22708,N_24156);
nor UO_2686 (O_2686,N_21520,N_23895);
nor UO_2687 (O_2687,N_21213,N_22165);
nor UO_2688 (O_2688,N_22601,N_21672);
nand UO_2689 (O_2689,N_24793,N_21174);
nand UO_2690 (O_2690,N_21232,N_20838);
nand UO_2691 (O_2691,N_21267,N_20015);
nor UO_2692 (O_2692,N_23824,N_21509);
nand UO_2693 (O_2693,N_23587,N_24292);
nand UO_2694 (O_2694,N_24406,N_20382);
nor UO_2695 (O_2695,N_23035,N_20022);
or UO_2696 (O_2696,N_22934,N_22092);
or UO_2697 (O_2697,N_21240,N_23034);
or UO_2698 (O_2698,N_20469,N_21419);
nor UO_2699 (O_2699,N_24640,N_21038);
or UO_2700 (O_2700,N_24661,N_20594);
and UO_2701 (O_2701,N_22237,N_23916);
or UO_2702 (O_2702,N_20383,N_22513);
nor UO_2703 (O_2703,N_20448,N_23252);
nor UO_2704 (O_2704,N_20760,N_21518);
nor UO_2705 (O_2705,N_24272,N_24286);
or UO_2706 (O_2706,N_21144,N_20493);
nand UO_2707 (O_2707,N_21207,N_22911);
or UO_2708 (O_2708,N_21803,N_20478);
nor UO_2709 (O_2709,N_24151,N_24875);
nand UO_2710 (O_2710,N_20476,N_24224);
and UO_2711 (O_2711,N_22271,N_23995);
or UO_2712 (O_2712,N_21947,N_21494);
xnor UO_2713 (O_2713,N_20434,N_21294);
and UO_2714 (O_2714,N_23793,N_20631);
nand UO_2715 (O_2715,N_23894,N_24584);
or UO_2716 (O_2716,N_24572,N_21780);
and UO_2717 (O_2717,N_22947,N_21416);
nor UO_2718 (O_2718,N_21918,N_21136);
or UO_2719 (O_2719,N_23847,N_21170);
nand UO_2720 (O_2720,N_23812,N_22007);
nand UO_2721 (O_2721,N_24210,N_24308);
nand UO_2722 (O_2722,N_21937,N_20522);
nand UO_2723 (O_2723,N_22513,N_24142);
nand UO_2724 (O_2724,N_24289,N_24433);
nand UO_2725 (O_2725,N_24281,N_21680);
nor UO_2726 (O_2726,N_21608,N_22549);
or UO_2727 (O_2727,N_21417,N_23175);
xor UO_2728 (O_2728,N_20887,N_21496);
nor UO_2729 (O_2729,N_22668,N_23984);
nor UO_2730 (O_2730,N_24331,N_23133);
or UO_2731 (O_2731,N_21095,N_23143);
nand UO_2732 (O_2732,N_24748,N_23614);
and UO_2733 (O_2733,N_22290,N_24457);
nor UO_2734 (O_2734,N_24580,N_20357);
nor UO_2735 (O_2735,N_22169,N_22241);
and UO_2736 (O_2736,N_23707,N_22039);
xor UO_2737 (O_2737,N_22526,N_22832);
nand UO_2738 (O_2738,N_20857,N_23441);
or UO_2739 (O_2739,N_20225,N_24526);
or UO_2740 (O_2740,N_24834,N_24013);
or UO_2741 (O_2741,N_23456,N_24229);
and UO_2742 (O_2742,N_24697,N_20990);
and UO_2743 (O_2743,N_20797,N_20231);
nor UO_2744 (O_2744,N_23231,N_21547);
and UO_2745 (O_2745,N_24812,N_22512);
and UO_2746 (O_2746,N_21799,N_22015);
nor UO_2747 (O_2747,N_22697,N_23111);
or UO_2748 (O_2748,N_24719,N_20146);
nand UO_2749 (O_2749,N_22267,N_20510);
nand UO_2750 (O_2750,N_20092,N_24345);
nand UO_2751 (O_2751,N_21348,N_23965);
and UO_2752 (O_2752,N_20296,N_23790);
and UO_2753 (O_2753,N_21321,N_20562);
or UO_2754 (O_2754,N_20048,N_22045);
nor UO_2755 (O_2755,N_21598,N_23531);
and UO_2756 (O_2756,N_24210,N_22350);
nor UO_2757 (O_2757,N_22650,N_21845);
nor UO_2758 (O_2758,N_21908,N_23559);
and UO_2759 (O_2759,N_20441,N_22530);
nand UO_2760 (O_2760,N_22995,N_21959);
or UO_2761 (O_2761,N_21412,N_20564);
or UO_2762 (O_2762,N_20840,N_20445);
nand UO_2763 (O_2763,N_20974,N_22034);
xnor UO_2764 (O_2764,N_20712,N_22744);
nor UO_2765 (O_2765,N_24442,N_21768);
and UO_2766 (O_2766,N_21766,N_24187);
nor UO_2767 (O_2767,N_23563,N_21711);
nand UO_2768 (O_2768,N_24576,N_22783);
nor UO_2769 (O_2769,N_24357,N_24641);
nor UO_2770 (O_2770,N_23995,N_21636);
nor UO_2771 (O_2771,N_21439,N_23020);
nor UO_2772 (O_2772,N_23142,N_22578);
nor UO_2773 (O_2773,N_22315,N_22879);
nand UO_2774 (O_2774,N_24026,N_23281);
nor UO_2775 (O_2775,N_23934,N_20981);
nor UO_2776 (O_2776,N_21931,N_22144);
and UO_2777 (O_2777,N_22776,N_20600);
or UO_2778 (O_2778,N_22950,N_24894);
nor UO_2779 (O_2779,N_21010,N_20256);
and UO_2780 (O_2780,N_22938,N_22805);
nand UO_2781 (O_2781,N_24447,N_24743);
or UO_2782 (O_2782,N_20570,N_23952);
and UO_2783 (O_2783,N_23096,N_23699);
nor UO_2784 (O_2784,N_22691,N_21849);
nor UO_2785 (O_2785,N_24306,N_24171);
nor UO_2786 (O_2786,N_24311,N_20714);
or UO_2787 (O_2787,N_20951,N_22580);
nor UO_2788 (O_2788,N_22588,N_21107);
nand UO_2789 (O_2789,N_23026,N_22138);
xor UO_2790 (O_2790,N_21995,N_22335);
nor UO_2791 (O_2791,N_23951,N_20632);
and UO_2792 (O_2792,N_22250,N_21360);
nor UO_2793 (O_2793,N_22734,N_20978);
nor UO_2794 (O_2794,N_22330,N_24150);
and UO_2795 (O_2795,N_21544,N_23674);
or UO_2796 (O_2796,N_20988,N_24426);
and UO_2797 (O_2797,N_21333,N_23636);
and UO_2798 (O_2798,N_20089,N_22717);
nand UO_2799 (O_2799,N_20368,N_23222);
or UO_2800 (O_2800,N_24374,N_23163);
nor UO_2801 (O_2801,N_23897,N_23456);
nand UO_2802 (O_2802,N_22560,N_24749);
nand UO_2803 (O_2803,N_20429,N_24626);
and UO_2804 (O_2804,N_21133,N_24521);
or UO_2805 (O_2805,N_23348,N_22725);
nor UO_2806 (O_2806,N_24221,N_22630);
and UO_2807 (O_2807,N_24846,N_23021);
and UO_2808 (O_2808,N_21724,N_23509);
and UO_2809 (O_2809,N_23233,N_21119);
and UO_2810 (O_2810,N_22698,N_24298);
nor UO_2811 (O_2811,N_24141,N_21011);
nor UO_2812 (O_2812,N_20619,N_23793);
xor UO_2813 (O_2813,N_23649,N_24450);
nand UO_2814 (O_2814,N_24963,N_21405);
or UO_2815 (O_2815,N_24819,N_22440);
and UO_2816 (O_2816,N_24852,N_20583);
nor UO_2817 (O_2817,N_20461,N_22851);
and UO_2818 (O_2818,N_22195,N_22047);
nor UO_2819 (O_2819,N_20453,N_20370);
nor UO_2820 (O_2820,N_21092,N_22318);
nor UO_2821 (O_2821,N_22027,N_24534);
nor UO_2822 (O_2822,N_21133,N_23871);
xnor UO_2823 (O_2823,N_22643,N_20401);
nor UO_2824 (O_2824,N_20378,N_21592);
nor UO_2825 (O_2825,N_23023,N_23413);
or UO_2826 (O_2826,N_20482,N_20229);
or UO_2827 (O_2827,N_23013,N_23043);
xor UO_2828 (O_2828,N_22142,N_23697);
and UO_2829 (O_2829,N_21852,N_23507);
nand UO_2830 (O_2830,N_24457,N_21790);
nor UO_2831 (O_2831,N_23200,N_20871);
or UO_2832 (O_2832,N_22406,N_20538);
or UO_2833 (O_2833,N_24655,N_21173);
nor UO_2834 (O_2834,N_24626,N_23513);
and UO_2835 (O_2835,N_23096,N_24331);
xor UO_2836 (O_2836,N_24739,N_22916);
and UO_2837 (O_2837,N_20762,N_21872);
nor UO_2838 (O_2838,N_21222,N_21140);
or UO_2839 (O_2839,N_21385,N_24158);
nor UO_2840 (O_2840,N_20449,N_21377);
and UO_2841 (O_2841,N_21944,N_24015);
or UO_2842 (O_2842,N_23335,N_22717);
and UO_2843 (O_2843,N_21366,N_24324);
or UO_2844 (O_2844,N_21412,N_21389);
nand UO_2845 (O_2845,N_21400,N_22835);
nand UO_2846 (O_2846,N_20617,N_24688);
nor UO_2847 (O_2847,N_22116,N_21431);
or UO_2848 (O_2848,N_21109,N_20976);
nor UO_2849 (O_2849,N_24955,N_20719);
nor UO_2850 (O_2850,N_21724,N_24108);
nand UO_2851 (O_2851,N_21129,N_23311);
nand UO_2852 (O_2852,N_21173,N_22465);
nor UO_2853 (O_2853,N_21520,N_24935);
nor UO_2854 (O_2854,N_21075,N_20493);
or UO_2855 (O_2855,N_20283,N_23906);
nor UO_2856 (O_2856,N_24012,N_22889);
or UO_2857 (O_2857,N_23161,N_22275);
nor UO_2858 (O_2858,N_22676,N_24128);
or UO_2859 (O_2859,N_23376,N_24830);
nand UO_2860 (O_2860,N_23197,N_21426);
and UO_2861 (O_2861,N_22796,N_20360);
nor UO_2862 (O_2862,N_21745,N_21378);
or UO_2863 (O_2863,N_24059,N_23228);
or UO_2864 (O_2864,N_20167,N_22912);
and UO_2865 (O_2865,N_21097,N_21465);
nand UO_2866 (O_2866,N_22328,N_22077);
or UO_2867 (O_2867,N_24855,N_22476);
or UO_2868 (O_2868,N_21950,N_21544);
nor UO_2869 (O_2869,N_22021,N_24900);
nor UO_2870 (O_2870,N_20505,N_22757);
and UO_2871 (O_2871,N_22721,N_24185);
nand UO_2872 (O_2872,N_20145,N_24582);
and UO_2873 (O_2873,N_21477,N_22153);
or UO_2874 (O_2874,N_22392,N_24471);
and UO_2875 (O_2875,N_20572,N_22526);
and UO_2876 (O_2876,N_20022,N_23701);
nor UO_2877 (O_2877,N_24620,N_22227);
nor UO_2878 (O_2878,N_24111,N_21891);
or UO_2879 (O_2879,N_22070,N_21862);
nand UO_2880 (O_2880,N_24596,N_22996);
or UO_2881 (O_2881,N_20877,N_21850);
nand UO_2882 (O_2882,N_21364,N_21708);
nand UO_2883 (O_2883,N_24340,N_20110);
xnor UO_2884 (O_2884,N_21428,N_21884);
nor UO_2885 (O_2885,N_23131,N_22752);
nor UO_2886 (O_2886,N_22655,N_23151);
or UO_2887 (O_2887,N_22607,N_21558);
nor UO_2888 (O_2888,N_22903,N_20866);
nor UO_2889 (O_2889,N_21725,N_21706);
or UO_2890 (O_2890,N_21026,N_20851);
nor UO_2891 (O_2891,N_22123,N_24533);
nand UO_2892 (O_2892,N_23017,N_22309);
or UO_2893 (O_2893,N_23977,N_22052);
nor UO_2894 (O_2894,N_20710,N_20230);
or UO_2895 (O_2895,N_24048,N_21094);
nand UO_2896 (O_2896,N_21578,N_21594);
or UO_2897 (O_2897,N_20707,N_21375);
nand UO_2898 (O_2898,N_23976,N_21952);
nor UO_2899 (O_2899,N_24773,N_22617);
nor UO_2900 (O_2900,N_20655,N_22889);
and UO_2901 (O_2901,N_21943,N_20532);
and UO_2902 (O_2902,N_24298,N_21323);
and UO_2903 (O_2903,N_20986,N_20791);
nand UO_2904 (O_2904,N_21538,N_24215);
or UO_2905 (O_2905,N_22967,N_21984);
nand UO_2906 (O_2906,N_20542,N_21180);
and UO_2907 (O_2907,N_24520,N_21292);
xnor UO_2908 (O_2908,N_23861,N_22243);
or UO_2909 (O_2909,N_21446,N_24279);
and UO_2910 (O_2910,N_21636,N_23785);
and UO_2911 (O_2911,N_23786,N_24145);
and UO_2912 (O_2912,N_20188,N_22603);
or UO_2913 (O_2913,N_21983,N_20307);
nand UO_2914 (O_2914,N_22096,N_22534);
nor UO_2915 (O_2915,N_21824,N_20449);
or UO_2916 (O_2916,N_21315,N_23035);
and UO_2917 (O_2917,N_24143,N_24797);
or UO_2918 (O_2918,N_22724,N_20258);
nor UO_2919 (O_2919,N_21961,N_22294);
and UO_2920 (O_2920,N_22207,N_24537);
nor UO_2921 (O_2921,N_24404,N_21571);
nand UO_2922 (O_2922,N_24568,N_23549);
and UO_2923 (O_2923,N_21493,N_21886);
nand UO_2924 (O_2924,N_22610,N_21382);
nand UO_2925 (O_2925,N_23908,N_23664);
nor UO_2926 (O_2926,N_24904,N_22414);
xor UO_2927 (O_2927,N_20610,N_21603);
nand UO_2928 (O_2928,N_20165,N_24226);
and UO_2929 (O_2929,N_22256,N_23062);
or UO_2930 (O_2930,N_24918,N_20211);
nand UO_2931 (O_2931,N_20809,N_21676);
or UO_2932 (O_2932,N_24971,N_20665);
and UO_2933 (O_2933,N_23109,N_23791);
and UO_2934 (O_2934,N_22786,N_23536);
and UO_2935 (O_2935,N_22066,N_23847);
nor UO_2936 (O_2936,N_24438,N_20499);
nor UO_2937 (O_2937,N_21055,N_22131);
and UO_2938 (O_2938,N_20871,N_22188);
nand UO_2939 (O_2939,N_24171,N_22530);
or UO_2940 (O_2940,N_21818,N_21724);
nand UO_2941 (O_2941,N_23572,N_22618);
nor UO_2942 (O_2942,N_24071,N_24167);
nor UO_2943 (O_2943,N_20378,N_21115);
nand UO_2944 (O_2944,N_21131,N_24094);
or UO_2945 (O_2945,N_21146,N_20629);
or UO_2946 (O_2946,N_24274,N_20651);
nor UO_2947 (O_2947,N_20436,N_23339);
nand UO_2948 (O_2948,N_22645,N_20184);
nor UO_2949 (O_2949,N_21065,N_20664);
and UO_2950 (O_2950,N_21317,N_22579);
and UO_2951 (O_2951,N_20651,N_23058);
nor UO_2952 (O_2952,N_23843,N_24932);
nor UO_2953 (O_2953,N_21246,N_20131);
nor UO_2954 (O_2954,N_21401,N_22419);
nand UO_2955 (O_2955,N_20711,N_23374);
nand UO_2956 (O_2956,N_20681,N_24268);
and UO_2957 (O_2957,N_20129,N_22216);
nand UO_2958 (O_2958,N_23265,N_24188);
nor UO_2959 (O_2959,N_24390,N_20084);
xor UO_2960 (O_2960,N_22061,N_22062);
or UO_2961 (O_2961,N_22003,N_24660);
and UO_2962 (O_2962,N_20143,N_22822);
nand UO_2963 (O_2963,N_23699,N_21003);
nand UO_2964 (O_2964,N_23708,N_22855);
and UO_2965 (O_2965,N_22662,N_22724);
or UO_2966 (O_2966,N_20168,N_24589);
or UO_2967 (O_2967,N_23089,N_20586);
and UO_2968 (O_2968,N_24664,N_24218);
or UO_2969 (O_2969,N_20112,N_21131);
or UO_2970 (O_2970,N_23751,N_22880);
and UO_2971 (O_2971,N_23340,N_21432);
and UO_2972 (O_2972,N_21508,N_21278);
and UO_2973 (O_2973,N_21913,N_21135);
or UO_2974 (O_2974,N_20919,N_24330);
nand UO_2975 (O_2975,N_21095,N_24046);
nor UO_2976 (O_2976,N_20706,N_23659);
nand UO_2977 (O_2977,N_21738,N_20252);
nand UO_2978 (O_2978,N_23588,N_21961);
or UO_2979 (O_2979,N_24363,N_23643);
nand UO_2980 (O_2980,N_22952,N_24067);
or UO_2981 (O_2981,N_24949,N_20677);
and UO_2982 (O_2982,N_24734,N_23445);
or UO_2983 (O_2983,N_22944,N_23908);
nor UO_2984 (O_2984,N_23122,N_23576);
nand UO_2985 (O_2985,N_23591,N_21140);
nand UO_2986 (O_2986,N_22828,N_24795);
or UO_2987 (O_2987,N_23488,N_23806);
and UO_2988 (O_2988,N_21915,N_22589);
or UO_2989 (O_2989,N_24206,N_24227);
and UO_2990 (O_2990,N_21719,N_24303);
nor UO_2991 (O_2991,N_24783,N_20063);
or UO_2992 (O_2992,N_20021,N_24504);
nand UO_2993 (O_2993,N_22380,N_20775);
or UO_2994 (O_2994,N_21619,N_20616);
and UO_2995 (O_2995,N_23294,N_20299);
nand UO_2996 (O_2996,N_24522,N_20123);
nor UO_2997 (O_2997,N_22256,N_23268);
nor UO_2998 (O_2998,N_24803,N_22347);
or UO_2999 (O_2999,N_21266,N_21506);
endmodule