module basic_5000_50000_5000_100_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_123,In_490);
nor U1 (N_1,In_803,In_4026);
or U2 (N_2,In_2166,In_2750);
nor U3 (N_3,In_2381,In_228);
nand U4 (N_4,In_694,In_3678);
nand U5 (N_5,In_3377,In_2911);
xnor U6 (N_6,In_2553,In_518);
nand U7 (N_7,In_2415,In_1035);
and U8 (N_8,In_4655,In_4436);
nand U9 (N_9,In_1371,In_1025);
xnor U10 (N_10,In_4785,In_3545);
nand U11 (N_11,In_3772,In_1037);
or U12 (N_12,In_873,In_336);
nor U13 (N_13,In_1871,In_1794);
and U14 (N_14,In_2391,In_677);
and U15 (N_15,In_3927,In_3355);
and U16 (N_16,In_974,In_4013);
xnor U17 (N_17,In_4608,In_2136);
and U18 (N_18,In_1459,In_23);
xnor U19 (N_19,In_4181,In_4313);
and U20 (N_20,In_1415,In_2384);
xnor U21 (N_21,In_1096,In_4184);
nor U22 (N_22,In_4534,In_4176);
nor U23 (N_23,In_1433,In_81);
nor U24 (N_24,In_2301,In_369);
nand U25 (N_25,In_4247,In_1229);
nor U26 (N_26,In_3963,In_1666);
nand U27 (N_27,In_4759,In_1768);
xor U28 (N_28,In_4398,In_362);
nor U29 (N_29,In_1596,In_3117);
and U30 (N_30,In_831,In_4798);
or U31 (N_31,In_2722,In_3968);
or U32 (N_32,In_3697,In_4673);
and U33 (N_33,In_4606,In_4022);
nand U34 (N_34,In_2247,In_4169);
xor U35 (N_35,In_132,In_3386);
or U36 (N_36,In_243,In_3908);
and U37 (N_37,In_1609,In_442);
xnor U38 (N_38,In_2386,In_3566);
nand U39 (N_39,In_2290,In_660);
nor U40 (N_40,In_3380,In_3374);
or U41 (N_41,In_594,In_2965);
nor U42 (N_42,In_954,In_882);
or U43 (N_43,In_3174,In_4119);
nand U44 (N_44,In_1112,In_1687);
and U45 (N_45,In_4154,In_2871);
nand U46 (N_46,In_2907,In_799);
and U47 (N_47,In_1838,In_2571);
and U48 (N_48,In_4469,In_2476);
or U49 (N_49,In_3334,In_4381);
and U50 (N_50,In_4165,In_4599);
nor U51 (N_51,In_3241,In_517);
nor U52 (N_52,In_2206,In_2398);
nand U53 (N_53,In_1006,In_2685);
nand U54 (N_54,In_3417,In_2740);
nor U55 (N_55,In_4416,In_1142);
and U56 (N_56,In_3115,In_959);
xor U57 (N_57,In_3606,In_927);
or U58 (N_58,In_2835,In_4190);
and U59 (N_59,In_1542,In_2489);
nand U60 (N_60,In_3257,In_4405);
and U61 (N_61,In_352,In_3654);
or U62 (N_62,In_1749,In_2847);
nor U63 (N_63,In_2117,In_4576);
or U64 (N_64,In_2648,In_1535);
nor U65 (N_65,In_977,In_1547);
and U66 (N_66,In_3224,In_560);
nand U67 (N_67,In_996,In_1360);
nand U68 (N_68,In_4720,In_118);
nand U69 (N_69,In_774,In_4246);
nor U70 (N_70,In_1225,In_1247);
xnor U71 (N_71,In_740,In_1237);
or U72 (N_72,In_2978,In_3580);
or U73 (N_73,In_1321,In_3325);
nor U74 (N_74,In_2987,In_110);
nand U75 (N_75,In_1361,In_3114);
nor U76 (N_76,In_334,In_1526);
xor U77 (N_77,In_4049,In_173);
and U78 (N_78,In_1414,In_4009);
and U79 (N_79,In_2914,In_1695);
xor U80 (N_80,In_1844,In_1391);
nor U81 (N_81,In_3581,In_468);
or U82 (N_82,In_2281,In_271);
nand U83 (N_83,In_170,In_3290);
and U84 (N_84,In_3037,In_2097);
nor U85 (N_85,In_1746,In_2518);
nor U86 (N_86,In_2974,In_3322);
or U87 (N_87,In_3902,In_3877);
nor U88 (N_88,In_19,In_1705);
and U89 (N_89,In_471,In_4306);
nand U90 (N_90,In_3160,In_3672);
xnor U91 (N_91,In_4039,In_3266);
or U92 (N_92,In_1818,In_3424);
and U93 (N_93,In_16,In_1207);
and U94 (N_94,In_3401,In_868);
and U95 (N_95,In_2155,In_934);
nor U96 (N_96,In_2278,In_864);
nand U97 (N_97,In_1032,In_2182);
or U98 (N_98,In_2851,In_4986);
and U99 (N_99,In_436,In_1560);
nor U100 (N_100,In_567,In_2880);
xor U101 (N_101,In_4484,In_3707);
nand U102 (N_102,In_2115,In_2929);
nor U103 (N_103,In_2869,In_1545);
nand U104 (N_104,In_4538,In_3218);
and U105 (N_105,In_4308,In_345);
nand U106 (N_106,In_1990,In_3625);
or U107 (N_107,In_230,In_218);
nor U108 (N_108,In_366,In_1500);
nand U109 (N_109,In_1453,In_3157);
nor U110 (N_110,In_2579,In_991);
nor U111 (N_111,In_1743,In_2064);
nand U112 (N_112,In_968,In_41);
nor U113 (N_113,In_154,In_3120);
nor U114 (N_114,In_1304,In_2540);
xor U115 (N_115,In_4153,In_2797);
or U116 (N_116,In_1355,In_4767);
nand U117 (N_117,In_2282,In_542);
nand U118 (N_118,In_669,In_666);
nand U119 (N_119,In_3652,In_4228);
or U120 (N_120,In_2331,In_4323);
or U121 (N_121,In_3835,In_426);
nor U122 (N_122,In_2569,In_950);
nand U123 (N_123,In_4114,In_3070);
nand U124 (N_124,In_446,In_2525);
nand U125 (N_125,In_2801,In_4668);
nor U126 (N_126,In_1062,In_4685);
and U127 (N_127,In_4595,In_1719);
xnor U128 (N_128,In_4096,In_358);
nor U129 (N_129,In_693,In_116);
and U130 (N_130,In_3867,In_800);
and U131 (N_131,In_1063,In_1823);
or U132 (N_132,In_2782,In_1981);
xnor U133 (N_133,In_1150,In_4556);
xnor U134 (N_134,In_2095,In_53);
or U135 (N_135,In_4806,In_4085);
and U136 (N_136,In_95,In_3512);
or U137 (N_137,In_1479,In_1727);
xnor U138 (N_138,In_1893,In_651);
nor U139 (N_139,In_3599,In_3893);
or U140 (N_140,In_3454,In_618);
xor U141 (N_141,In_3880,In_4237);
nand U142 (N_142,In_3742,In_3913);
nor U143 (N_143,In_1486,In_2304);
or U144 (N_144,In_1344,In_4990);
or U145 (N_145,In_3118,In_4264);
nor U146 (N_146,In_3941,In_1730);
and U147 (N_147,In_4743,In_2169);
or U148 (N_148,In_3737,In_2335);
or U149 (N_149,In_2733,In_2165);
and U150 (N_150,In_2626,In_4255);
and U151 (N_151,In_3222,In_4771);
and U152 (N_152,In_2709,In_531);
or U153 (N_153,In_2421,In_1357);
and U154 (N_154,In_696,In_1303);
nor U155 (N_155,In_854,In_4582);
nand U156 (N_156,In_569,In_681);
or U157 (N_157,In_2590,In_1909);
xnor U158 (N_158,In_3148,In_248);
nor U159 (N_159,In_1863,In_2046);
and U160 (N_160,In_1791,In_2890);
nor U161 (N_161,In_4651,In_4631);
nand U162 (N_162,In_3031,In_1916);
nand U163 (N_163,In_4280,In_1275);
nand U164 (N_164,In_3244,In_4678);
nor U165 (N_165,In_4338,In_3998);
xnor U166 (N_166,In_1552,In_689);
nor U167 (N_167,In_1358,In_732);
or U168 (N_168,In_2359,In_4523);
xor U169 (N_169,In_3951,In_4440);
and U170 (N_170,In_2234,In_1272);
and U171 (N_171,In_3048,In_4777);
or U172 (N_172,In_3069,In_3799);
nor U173 (N_173,In_4449,In_2804);
and U174 (N_174,In_4768,In_22);
or U175 (N_175,In_1093,In_2082);
and U176 (N_176,In_1216,In_2758);
and U177 (N_177,In_615,In_4647);
or U178 (N_178,In_4648,In_4772);
and U179 (N_179,In_746,In_4645);
nor U180 (N_180,In_3590,In_1720);
or U181 (N_181,In_1245,In_308);
nor U182 (N_182,In_26,In_441);
nand U183 (N_183,In_1997,In_3574);
or U184 (N_184,In_3495,In_3211);
xnor U185 (N_185,In_4949,In_3427);
or U186 (N_186,In_2466,In_2402);
nor U187 (N_187,In_1809,In_4628);
nand U188 (N_188,In_2334,In_1228);
nor U189 (N_189,In_3777,In_190);
or U190 (N_190,In_4840,In_2267);
xnor U191 (N_191,In_2495,In_4404);
nor U192 (N_192,In_3614,In_611);
and U193 (N_193,In_3766,In_2603);
and U194 (N_194,In_313,In_891);
nor U195 (N_195,In_2811,In_1369);
and U196 (N_196,In_760,In_2490);
and U197 (N_197,In_4197,In_4187);
or U198 (N_198,In_668,In_2452);
and U199 (N_199,In_4590,In_1378);
nor U200 (N_200,In_4396,In_4042);
nor U201 (N_201,In_4159,In_926);
or U202 (N_202,In_1167,In_1205);
and U203 (N_203,In_4964,In_4135);
or U204 (N_204,In_226,In_3932);
nor U205 (N_205,In_4142,In_4295);
and U206 (N_206,In_1038,In_4683);
or U207 (N_207,In_3936,In_1024);
nor U208 (N_208,In_1034,In_1302);
nor U209 (N_209,In_2455,In_3004);
xor U210 (N_210,In_4212,In_3522);
and U211 (N_211,In_2552,In_2408);
or U212 (N_212,In_4289,In_4468);
and U213 (N_213,In_3461,In_2539);
nor U214 (N_214,In_2017,In_2680);
and U215 (N_215,In_1004,In_3516);
and U216 (N_216,In_4411,In_4883);
nor U217 (N_217,In_1269,In_3188);
and U218 (N_218,In_4109,In_2870);
or U219 (N_219,In_3565,In_2118);
or U220 (N_220,In_2312,In_2152);
nand U221 (N_221,In_1769,In_2993);
nor U222 (N_222,In_4494,In_2706);
or U223 (N_223,In_4605,In_2);
or U224 (N_224,In_305,In_1536);
nor U225 (N_225,In_4170,In_3588);
or U226 (N_226,In_1690,In_3747);
nor U227 (N_227,In_3882,In_1496);
nand U228 (N_228,In_995,In_1194);
nand U229 (N_229,In_2394,In_3820);
nand U230 (N_230,In_4562,In_4200);
and U231 (N_231,In_4307,In_1723);
xnor U232 (N_232,In_1694,In_559);
and U233 (N_233,In_1429,In_802);
and U234 (N_234,In_2034,In_4579);
or U235 (N_235,In_300,In_674);
nor U236 (N_236,In_410,In_4133);
nand U237 (N_237,In_3662,In_250);
and U238 (N_238,In_1508,In_2293);
or U239 (N_239,In_3217,In_853);
nor U240 (N_240,In_379,In_2143);
and U241 (N_241,In_2008,In_79);
xnor U242 (N_242,In_4000,In_3367);
and U243 (N_243,In_855,In_2717);
xnor U244 (N_244,In_734,In_144);
nand U245 (N_245,In_4898,In_4058);
nand U246 (N_246,In_1485,In_3277);
nor U247 (N_247,In_3783,In_4808);
nand U248 (N_248,In_290,In_820);
nor U249 (N_249,In_4548,In_1072);
or U250 (N_250,In_4732,In_826);
and U251 (N_251,In_667,In_4707);
or U252 (N_252,In_4378,In_908);
and U253 (N_253,In_3883,In_119);
and U254 (N_254,In_2789,In_4310);
nand U255 (N_255,In_470,In_2736);
nor U256 (N_256,In_1370,In_916);
nor U257 (N_257,In_4445,In_3492);
xor U258 (N_258,In_1789,In_4101);
and U259 (N_259,In_1095,In_9);
nor U260 (N_260,In_627,In_1382);
nor U261 (N_261,In_215,In_398);
and U262 (N_262,In_1330,In_121);
nor U263 (N_263,In_1270,In_3842);
nand U264 (N_264,In_1439,In_2371);
and U265 (N_265,In_4791,In_4331);
and U266 (N_266,In_166,In_384);
nor U267 (N_267,In_3043,In_1885);
or U268 (N_268,In_1550,In_1111);
nor U269 (N_269,In_2537,In_3579);
xor U270 (N_270,In_1423,In_3317);
nand U271 (N_271,In_3119,In_4691);
or U272 (N_272,In_4254,In_637);
nor U273 (N_273,In_2682,In_1153);
nand U274 (N_274,In_4792,In_2388);
and U275 (N_275,In_3987,In_2816);
xor U276 (N_276,In_3035,In_2439);
or U277 (N_277,In_4884,In_3901);
xor U278 (N_278,In_874,In_3716);
nand U279 (N_279,In_315,In_214);
nand U280 (N_280,In_3628,In_256);
or U281 (N_281,In_4415,In_1677);
or U282 (N_282,In_133,In_2419);
nor U283 (N_283,In_2461,In_1267);
or U284 (N_284,In_688,In_2689);
or U285 (N_285,In_437,In_3226);
nor U286 (N_286,In_2201,In_3291);
or U287 (N_287,In_4361,In_1926);
xnor U288 (N_288,In_946,In_2776);
and U289 (N_289,In_1193,In_4367);
nor U290 (N_290,In_2948,In_425);
or U291 (N_291,In_993,In_113);
and U292 (N_292,In_2265,In_4906);
or U293 (N_293,In_3866,In_3409);
and U294 (N_294,In_3456,In_2001);
and U295 (N_295,In_100,In_4850);
nand U296 (N_296,In_1957,In_1758);
xor U297 (N_297,In_4118,In_4419);
or U298 (N_298,In_3520,In_2954);
nand U299 (N_299,In_3139,In_1036);
nand U300 (N_300,In_307,In_3832);
nand U301 (N_301,In_3145,In_449);
nor U302 (N_302,In_2385,In_804);
nor U303 (N_303,In_487,In_4196);
nand U304 (N_304,In_1709,In_2751);
and U305 (N_305,In_911,In_70);
or U306 (N_306,In_310,In_3650);
or U307 (N_307,In_4745,In_3900);
nor U308 (N_308,In_4446,In_3939);
xnor U309 (N_309,In_3863,In_4554);
or U310 (N_310,In_2109,In_3972);
and U311 (N_311,In_3423,In_1203);
and U312 (N_312,In_767,In_4193);
and U313 (N_313,In_335,In_287);
and U314 (N_314,In_4565,In_2876);
xor U315 (N_315,In_4974,In_1314);
or U316 (N_316,In_1230,In_2899);
xnor U317 (N_317,In_2777,In_1611);
nor U318 (N_318,In_687,In_4868);
nor U319 (N_319,In_4509,In_2240);
and U320 (N_320,In_4048,In_810);
nand U321 (N_321,In_2977,In_3519);
nor U322 (N_322,In_2687,In_1886);
and U323 (N_323,In_1455,In_2846);
nor U324 (N_324,In_1122,In_3234);
or U325 (N_325,In_4129,In_2674);
and U326 (N_326,In_4244,In_2767);
xnor U327 (N_327,In_2494,In_1837);
or U328 (N_328,In_1223,In_3833);
nand U329 (N_329,In_1359,In_2252);
and U330 (N_330,In_3812,In_3845);
nor U331 (N_331,In_435,In_2796);
nor U332 (N_332,In_4724,In_3757);
and U333 (N_333,In_2129,In_540);
nand U334 (N_334,In_3978,In_3916);
and U335 (N_335,In_2465,In_2480);
nor U336 (N_336,In_4741,In_199);
nand U337 (N_337,In_4010,In_2612);
xnor U338 (N_338,In_4662,In_929);
nand U339 (N_339,In_2052,In_3705);
nand U340 (N_340,In_4708,In_3743);
or U341 (N_341,In_2633,In_1989);
nor U342 (N_342,In_3432,In_4168);
or U343 (N_343,In_3817,In_4991);
nand U344 (N_344,In_3989,In_4750);
or U345 (N_345,In_4158,In_84);
nand U346 (N_346,In_3138,In_1379);
or U347 (N_347,In_4797,In_4814);
or U348 (N_348,In_661,In_500);
nand U349 (N_349,In_2319,In_4150);
nand U350 (N_350,In_2238,In_238);
and U351 (N_351,In_1450,In_4624);
and U352 (N_352,In_3959,In_3762);
and U353 (N_353,In_2351,In_3155);
nor U354 (N_354,In_201,In_4033);
and U355 (N_355,In_3072,In_102);
nor U356 (N_356,In_1440,In_4302);
nand U357 (N_357,In_3256,In_1435);
and U358 (N_358,In_1045,In_3789);
nor U359 (N_359,In_1441,In_1775);
nor U360 (N_360,In_3352,In_4177);
xor U361 (N_361,In_1334,In_3894);
xor U362 (N_362,In_2272,In_3230);
or U363 (N_363,In_4065,In_2865);
nand U364 (N_364,In_1891,In_3164);
or U365 (N_365,In_1353,In_2275);
nor U366 (N_366,In_4387,In_1143);
or U367 (N_367,In_4551,In_1876);
nand U368 (N_368,In_2326,In_2330);
or U369 (N_369,In_1742,In_4123);
nand U370 (N_370,In_2288,In_148);
and U371 (N_371,In_2262,In_3017);
nor U372 (N_372,In_4564,In_4373);
and U373 (N_373,In_4781,In_3929);
nor U374 (N_374,In_3755,In_671);
nor U375 (N_375,In_4427,In_3607);
nor U376 (N_376,In_2181,In_4896);
or U377 (N_377,In_564,In_3602);
nand U378 (N_378,In_2891,In_3810);
xor U379 (N_379,In_3233,In_4443);
or U380 (N_380,In_1315,In_706);
or U381 (N_381,In_3295,In_985);
or U382 (N_382,In_1983,In_2597);
nor U383 (N_383,In_4339,In_3064);
nor U384 (N_384,In_2347,In_2396);
xnor U385 (N_385,In_1023,In_1868);
nand U386 (N_386,In_1310,In_3521);
xor U387 (N_387,In_1186,In_1985);
nand U388 (N_388,In_935,In_1057);
and U389 (N_389,In_97,In_3045);
nand U390 (N_390,In_1800,In_1930);
xor U391 (N_391,In_2091,In_1832);
nor U392 (N_392,In_2053,In_1388);
and U393 (N_393,In_2089,In_327);
or U394 (N_394,In_3675,In_3736);
nor U395 (N_395,In_3729,In_638);
nand U396 (N_396,In_3919,In_3370);
nand U397 (N_397,In_1603,In_3977);
nor U398 (N_398,In_511,In_2227);
xnor U399 (N_399,In_3659,In_1759);
or U400 (N_400,In_1470,In_39);
and U401 (N_401,In_1480,In_922);
and U402 (N_402,In_1195,In_1491);
or U403 (N_403,In_1962,In_1325);
or U404 (N_404,In_2210,In_4968);
or U405 (N_405,In_1668,In_4652);
nand U406 (N_406,In_406,In_3105);
xor U407 (N_407,In_3215,In_1444);
or U408 (N_408,In_964,In_5);
nand U409 (N_409,In_1646,In_2069);
nand U410 (N_410,In_2827,In_1208);
and U411 (N_411,In_2039,In_3931);
nand U412 (N_412,In_8,In_3054);
nand U413 (N_413,In_349,In_3273);
nand U414 (N_414,In_2690,In_2170);
nor U415 (N_415,In_3760,In_2711);
and U416 (N_416,In_2470,In_1171);
and U417 (N_417,In_4262,In_172);
xnor U418 (N_418,In_2497,In_4452);
nand U419 (N_419,In_4594,In_4183);
and U420 (N_420,In_3798,In_3554);
xnor U421 (N_421,In_4689,In_3227);
and U422 (N_422,In_2176,In_3128);
or U423 (N_423,In_4575,In_1890);
nand U424 (N_424,In_2418,In_2045);
and U425 (N_425,In_2560,In_4438);
and U426 (N_426,In_2822,In_790);
nand U427 (N_427,In_3744,In_3408);
nand U428 (N_428,In_4297,In_2973);
or U429 (N_429,In_1389,In_1722);
and U430 (N_430,In_285,In_850);
or U431 (N_431,In_145,In_1580);
or U432 (N_432,In_701,In_719);
or U433 (N_433,In_1406,In_888);
nand U434 (N_434,In_2931,In_2239);
nand U435 (N_435,In_259,In_4904);
or U436 (N_436,In_4859,In_1638);
or U437 (N_437,In_3245,In_2456);
xnor U438 (N_438,In_4189,In_1704);
or U439 (N_439,In_4722,In_455);
nor U440 (N_440,In_3410,In_549);
nor U441 (N_441,In_4945,In_3240);
nor U442 (N_442,In_3484,In_466);
and U443 (N_443,In_2500,In_4700);
and U444 (N_444,In_3437,In_4081);
nor U445 (N_445,In_780,In_2493);
nor U446 (N_446,In_3618,In_4047);
nand U447 (N_447,In_4340,In_4574);
or U448 (N_448,In_2984,In_754);
and U449 (N_449,In_2988,In_3061);
and U450 (N_450,In_1784,In_3903);
xnor U451 (N_451,In_952,In_3156);
nand U452 (N_452,In_1577,In_2852);
xor U453 (N_453,In_1711,In_4076);
nand U454 (N_454,In_2764,In_955);
nand U455 (N_455,In_2557,In_4681);
or U456 (N_456,In_2369,In_3028);
nor U457 (N_457,In_2739,In_1628);
nor U458 (N_458,In_2694,In_1101);
nor U459 (N_459,In_3020,In_2932);
nand U460 (N_460,In_4229,In_141);
or U461 (N_461,In_4252,In_1110);
nand U462 (N_462,In_1472,In_2507);
or U463 (N_463,In_72,In_1263);
nand U464 (N_464,In_3311,In_4265);
nor U465 (N_465,In_3236,In_4656);
and U466 (N_466,In_2892,In_4971);
nand U467 (N_467,In_295,In_1581);
nor U468 (N_468,In_2757,In_2018);
or U469 (N_469,In_3771,In_348);
nor U470 (N_470,In_4210,In_3385);
or U471 (N_471,In_3421,In_4935);
nand U472 (N_472,In_477,In_2520);
and U473 (N_473,In_3875,In_4434);
and U474 (N_474,In_2729,In_304);
nand U475 (N_475,In_3981,In_2619);
or U476 (N_476,In_2230,In_3947);
nand U477 (N_477,In_3807,In_1168);
nand U478 (N_478,In_2236,In_2642);
and U479 (N_479,In_645,In_1220);
or U480 (N_480,In_4890,In_3605);
nor U481 (N_481,In_1113,In_2270);
nand U482 (N_482,In_1123,In_1614);
nor U483 (N_483,In_4638,In_3557);
nor U484 (N_484,In_4386,In_476);
nor U485 (N_485,In_1060,In_3725);
nand U486 (N_486,In_1907,In_3319);
nor U487 (N_487,In_1495,In_227);
or U488 (N_488,In_3753,In_3076);
or U489 (N_489,In_4248,In_4223);
nor U490 (N_490,In_3383,In_883);
and U491 (N_491,In_2881,In_2550);
or U492 (N_492,In_83,In_3000);
nand U493 (N_493,In_270,In_4976);
nand U494 (N_494,In_3252,In_3976);
nand U495 (N_495,In_1086,In_522);
nand U496 (N_496,In_2287,In_3369);
xor U497 (N_497,In_3831,In_3970);
or U498 (N_498,In_2924,In_1965);
and U499 (N_499,In_4395,In_2073);
xor U500 (N_500,In_1179,In_856);
nor U501 (N_501,In_4105,In_4028);
nor U502 (N_502,In_4211,In_2504);
or U503 (N_503,In_1601,In_262);
nor U504 (N_504,In_1154,In_1428);
or U505 (N_505,In_3668,In_907);
nand U506 (N_506,In_3123,In_4241);
nor U507 (N_507,In_1676,In_2445);
and U508 (N_508,In_3053,In_2409);
or U509 (N_509,In_465,In_4222);
or U510 (N_510,In_990,In_443);
and U511 (N_511,In_1782,In_3400);
nand U512 (N_512,In_3336,In_858);
nand U513 (N_513,In_833,In_2228);
or U514 (N_514,In_4359,In_1944);
and U515 (N_515,In_4642,In_1982);
nor U516 (N_516,N_330,In_328);
nor U517 (N_517,In_3356,In_623);
or U518 (N_518,In_4205,In_2033);
xor U519 (N_519,In_2141,In_1814);
xor U520 (N_520,In_3805,In_1517);
or U521 (N_521,In_128,In_3542);
nand U522 (N_522,In_127,In_4173);
nor U523 (N_523,In_2337,In_3523);
or U524 (N_524,In_4510,In_2483);
nor U525 (N_525,In_4847,In_2621);
nor U526 (N_526,In_581,In_3300);
and U527 (N_527,In_1820,In_4186);
and U528 (N_528,In_2077,N_52);
or U529 (N_529,N_34,In_2066);
nand U530 (N_530,In_634,In_2231);
xnor U531 (N_531,In_3100,In_3003);
or U532 (N_532,In_67,In_1731);
or U533 (N_533,In_2375,In_2332);
nand U534 (N_534,In_4334,In_2510);
nand U535 (N_535,In_197,In_401);
nand U536 (N_536,In_4863,N_33);
nand U537 (N_537,In_3040,In_2131);
xor U538 (N_538,In_4011,In_2156);
nor U539 (N_539,In_1795,In_3622);
nor U540 (N_540,In_727,In_3459);
nand U541 (N_541,In_1588,N_406);
or U542 (N_542,In_2083,In_1816);
xor U543 (N_543,In_456,In_3429);
nor U544 (N_544,In_1793,In_724);
or U545 (N_545,In_2198,In_1657);
nor U546 (N_546,In_1710,In_376);
and U547 (N_547,In_779,In_1578);
xor U548 (N_548,N_212,In_444);
nor U549 (N_549,In_1853,In_3026);
nor U550 (N_550,In_733,In_2966);
nand U551 (N_551,In_1328,In_3485);
nand U552 (N_552,In_2926,In_1128);
xor U553 (N_553,N_480,In_3480);
nand U554 (N_554,In_4922,N_58);
nand U555 (N_555,In_3814,In_1329);
or U556 (N_556,In_2828,In_363);
nand U557 (N_557,In_432,In_795);
nand U558 (N_558,In_1082,In_2468);
nand U559 (N_559,In_3535,In_4131);
nor U560 (N_560,In_2605,In_1978);
nand U561 (N_561,In_1796,In_4143);
nor U562 (N_562,In_4912,In_3996);
nor U563 (N_563,N_415,In_2716);
xor U564 (N_564,In_2449,In_3089);
and U565 (N_565,In_2889,In_2204);
or U566 (N_566,In_3463,In_3125);
xnor U567 (N_567,In_1014,In_520);
and U568 (N_568,In_344,In_2615);
and U569 (N_569,In_4283,In_3841);
or U570 (N_570,In_3656,In_825);
nor U571 (N_571,In_2641,In_3238);
or U572 (N_572,In_2661,In_546);
nand U573 (N_573,N_120,In_4905);
nor U574 (N_574,In_4287,N_446);
xor U575 (N_575,In_4275,In_4122);
nor U576 (N_576,In_1170,In_1187);
nor U577 (N_577,In_341,N_397);
nor U578 (N_578,In_4845,In_2424);
and U579 (N_579,In_3464,In_3392);
nor U580 (N_580,In_3691,N_493);
and U581 (N_581,In_1282,In_454);
nand U582 (N_582,In_759,In_509);
nand U583 (N_583,In_4356,In_2883);
or U584 (N_584,In_3517,In_3284);
and U585 (N_585,In_194,In_4008);
nand U586 (N_586,In_4774,In_2505);
and U587 (N_587,In_1531,In_3220);
and U588 (N_588,In_263,In_3112);
nand U589 (N_589,In_3730,In_3184);
nor U590 (N_590,In_4382,In_3062);
or U591 (N_591,In_2382,In_3710);
nand U592 (N_592,In_167,In_2982);
nor U593 (N_593,In_1394,N_196);
or U594 (N_594,N_84,In_139);
nor U595 (N_595,In_1482,In_4420);
nand U596 (N_596,In_956,N_190);
nand U597 (N_597,In_2607,In_1689);
nand U598 (N_598,In_1770,In_2019);
and U599 (N_599,In_1176,N_348);
nor U600 (N_600,In_4640,In_4711);
xor U601 (N_601,In_871,N_81);
and U602 (N_602,In_4269,In_4267);
xor U603 (N_603,In_3379,In_1373);
xnor U604 (N_604,In_684,In_4240);
and U605 (N_605,In_1684,In_2354);
and U606 (N_606,In_3474,In_3102);
and U607 (N_607,In_1049,In_2416);
or U608 (N_608,In_2655,In_3056);
nor U609 (N_609,In_1262,In_4513);
or U610 (N_610,In_3734,In_1172);
nand U611 (N_611,In_140,In_3924);
or U612 (N_612,In_3250,In_592);
nor U613 (N_613,In_3660,In_4588);
and U614 (N_614,N_275,In_1341);
nand U615 (N_615,In_3134,N_180);
xor U616 (N_616,In_1632,N_82);
and U617 (N_617,In_1084,In_1674);
or U618 (N_618,In_1539,In_2813);
nand U619 (N_619,In_1738,In_3195);
nand U620 (N_620,In_1280,In_2208);
and U621 (N_621,N_163,In_4451);
nor U622 (N_622,N_460,In_4734);
nor U623 (N_623,N_471,In_1409);
nor U624 (N_624,In_663,In_3508);
and U625 (N_625,In_7,In_2395);
nor U626 (N_626,In_984,In_1265);
or U627 (N_627,In_4633,In_3288);
and U628 (N_628,In_4972,In_402);
and U629 (N_629,In_403,In_2915);
or U630 (N_630,In_2316,N_256);
nor U631 (N_631,In_630,N_16);
xnor U632 (N_632,In_2631,In_863);
xor U633 (N_633,In_322,In_4512);
and U634 (N_634,In_338,In_1197);
nand U635 (N_635,In_784,In_3286);
or U636 (N_636,N_417,In_1018);
or U637 (N_637,In_2310,In_2488);
and U638 (N_638,N_83,In_2454);
xor U639 (N_639,In_2686,N_125);
and U640 (N_640,In_2837,In_3039);
and U641 (N_641,In_4162,In_3425);
nor U642 (N_642,In_2844,In_246);
nor U643 (N_643,In_2738,In_589);
or U644 (N_644,N_124,In_1050);
or U645 (N_645,In_1565,In_3342);
or U646 (N_646,In_115,N_235);
nand U647 (N_647,N_472,In_1697);
nor U648 (N_648,In_4729,In_2617);
xnor U649 (N_649,In_2241,In_4999);
nand U650 (N_650,In_2684,In_3131);
nor U651 (N_651,In_828,N_138);
nand U652 (N_652,In_1297,In_711);
nand U653 (N_653,In_460,In_3462);
and U654 (N_654,In_1227,In_1288);
nor U655 (N_655,N_207,In_3268);
nor U656 (N_656,In_1412,In_111);
or U657 (N_657,In_4946,In_2766);
nor U658 (N_658,In_2216,In_4414);
or U659 (N_659,In_457,In_1156);
or U660 (N_660,In_2538,In_2158);
and U661 (N_661,In_3333,In_3768);
and U662 (N_662,In_3731,In_453);
or U663 (N_663,In_2110,In_2584);
xnor U664 (N_664,In_4149,In_47);
nor U665 (N_665,In_3345,In_2258);
or U666 (N_666,In_2487,In_1664);
nand U667 (N_667,In_2574,In_3578);
and U668 (N_668,In_1102,In_3878);
nand U669 (N_669,In_2087,In_3569);
and U670 (N_670,In_1942,In_4107);
or U671 (N_671,In_3065,In_3327);
nand U672 (N_672,In_3988,In_3872);
xor U673 (N_673,In_4916,In_3177);
nor U674 (N_674,In_999,In_1892);
and U675 (N_675,In_4095,In_2566);
nor U676 (N_676,In_483,In_419);
nand U677 (N_677,In_182,In_4439);
nand U678 (N_678,In_2908,In_4881);
nor U679 (N_679,In_1839,N_458);
nand U680 (N_680,N_292,N_318);
xor U681 (N_681,In_1963,In_3183);
or U682 (N_682,In_3600,In_4994);
nor U683 (N_683,In_3819,In_1860);
xnor U684 (N_684,N_238,In_2486);
or U685 (N_685,In_3792,N_189);
or U686 (N_686,N_26,N_398);
or U687 (N_687,In_3852,In_2010);
nand U688 (N_688,In_2645,N_116);
nand U689 (N_689,In_3001,In_1575);
or U690 (N_690,In_2100,In_4023);
nand U691 (N_691,In_3640,In_835);
and U692 (N_692,In_2744,In_1872);
and U693 (N_693,In_4764,In_629);
xnor U694 (N_694,In_422,In_1144);
nor U695 (N_695,In_3358,In_830);
or U696 (N_696,In_3381,In_936);
or U697 (N_697,In_680,In_1248);
nand U698 (N_698,In_4349,In_2765);
nand U699 (N_699,In_1094,In_940);
nand U700 (N_700,In_4475,In_707);
or U701 (N_701,In_554,In_4755);
nor U702 (N_702,In_1925,In_729);
nor U703 (N_703,In_4397,In_1938);
nand U704 (N_704,In_332,In_2446);
or U705 (N_705,In_152,In_2596);
xnor U706 (N_706,In_2791,N_298);
nor U707 (N_707,In_705,N_178);
or U708 (N_708,In_3204,In_2457);
nand U709 (N_709,In_1008,In_1556);
and U710 (N_710,In_4032,N_290);
nor U711 (N_711,In_1913,In_628);
or U712 (N_712,In_2320,In_1033);
nor U713 (N_713,In_2997,In_3752);
or U714 (N_714,N_134,In_3365);
and U715 (N_715,N_429,In_555);
nor U716 (N_716,In_4823,In_309);
or U717 (N_717,In_122,In_2779);
or U718 (N_718,In_3797,In_2372);
and U719 (N_719,In_3967,In_4675);
xor U720 (N_720,In_819,In_756);
or U721 (N_721,In_2610,N_210);
nand U722 (N_722,In_2874,In_2122);
or U723 (N_723,In_3922,In_3851);
nor U724 (N_724,In_114,In_4544);
or U725 (N_725,N_461,In_4341);
and U726 (N_726,In_776,In_4684);
or U727 (N_727,In_945,In_4717);
and U728 (N_728,In_1622,In_3434);
nor U729 (N_729,In_3098,In_2121);
nor U730 (N_730,In_885,In_3687);
and U731 (N_731,In_4923,In_3940);
and U732 (N_732,In_3315,In_360);
nor U733 (N_733,In_1337,In_893);
nor U734 (N_734,N_324,In_3185);
and U735 (N_735,In_4329,In_2970);
nand U736 (N_736,In_2922,In_4784);
or U737 (N_737,In_4666,In_1798);
nor U738 (N_738,In_4347,In_876);
or U739 (N_739,In_1069,In_1858);
nand U740 (N_740,In_608,In_333);
and U741 (N_741,In_258,N_162);
nand U742 (N_742,In_3677,In_2675);
nand U743 (N_743,In_4852,N_423);
nand U744 (N_744,In_2795,In_463);
and U745 (N_745,In_3524,In_1780);
and U746 (N_746,In_4182,In_1100);
nand U747 (N_747,In_1562,In_1501);
nand U748 (N_748,In_2530,In_771);
or U749 (N_749,In_4163,In_1534);
or U750 (N_750,In_2853,N_281);
and U751 (N_751,In_4489,In_4456);
or U752 (N_752,In_1984,In_1005);
or U753 (N_753,In_2000,In_2047);
and U754 (N_754,In_4071,In_4132);
nor U755 (N_755,In_4502,In_4238);
or U756 (N_756,In_1098,In_1680);
or U757 (N_757,In_3868,In_2271);
and U758 (N_758,In_464,In_292);
nand U759 (N_759,In_4524,In_3096);
and U760 (N_760,In_142,In_1642);
or U761 (N_761,In_4903,In_27);
nor U762 (N_762,In_3075,In_2492);
or U763 (N_763,In_1318,N_387);
xnor U764 (N_764,In_4503,In_1299);
nor U765 (N_765,In_3873,In_3198);
or U766 (N_766,In_4615,In_1620);
or U767 (N_767,N_205,In_1867);
or U768 (N_768,In_2377,In_4498);
and U769 (N_769,In_1090,In_3391);
or U770 (N_770,In_3394,In_4927);
xor U771 (N_771,In_3280,N_434);
xnor U772 (N_772,N_490,N_277);
and U773 (N_773,In_4932,In_1960);
and U774 (N_774,In_3682,In_1767);
nand U775 (N_775,In_1996,N_174);
xor U776 (N_776,N_363,In_4253);
nand U777 (N_777,In_3717,In_61);
nor U778 (N_778,In_3354,In_2094);
and U779 (N_779,In_786,In_1012);
or U780 (N_780,In_2072,In_4145);
xor U781 (N_781,In_3749,In_2971);
and U782 (N_782,In_601,In_595);
and U783 (N_783,N_495,In_2154);
and U784 (N_784,In_1055,In_14);
or U785 (N_785,In_3975,In_3500);
nor U786 (N_786,In_1326,In_3860);
nor U787 (N_787,In_4885,In_3144);
or U788 (N_788,In_3644,In_4084);
xnor U789 (N_789,In_2514,In_2266);
nand U790 (N_790,N_231,In_1192);
xnor U791 (N_791,In_3671,In_764);
xnor U792 (N_792,In_3570,In_4731);
nor U793 (N_793,In_3231,In_320);
and U794 (N_794,In_2338,N_46);
and U795 (N_795,In_526,In_1068);
xor U796 (N_796,In_3150,In_4568);
nand U797 (N_797,In_1551,In_1636);
and U798 (N_798,In_2781,In_4120);
nor U799 (N_799,In_2336,In_4679);
or U800 (N_800,In_4790,In_302);
nand U801 (N_801,In_4887,In_2437);
nand U802 (N_802,In_3491,In_458);
and U803 (N_803,N_267,In_2392);
or U804 (N_804,In_4172,In_354);
nor U805 (N_805,In_626,In_699);
or U806 (N_806,N_409,In_274);
and U807 (N_807,N_215,N_271);
nor U808 (N_808,In_1623,In_1349);
or U809 (N_809,In_4141,In_4518);
nor U810 (N_810,In_387,In_4217);
nor U811 (N_811,In_2957,In_781);
and U812 (N_812,In_1502,In_2964);
and U813 (N_813,In_4225,In_2450);
nor U814 (N_814,In_4718,In_982);
xnor U815 (N_815,In_3670,In_4460);
nand U816 (N_816,In_2070,In_3326);
nor U817 (N_817,In_1013,In_599);
or U818 (N_818,N_76,In_4947);
xor U819 (N_819,In_1828,In_223);
nand U820 (N_820,In_583,In_4546);
or U821 (N_821,In_1713,In_3175);
xor U822 (N_822,In_633,In_391);
xor U823 (N_823,In_25,In_3285);
xor U824 (N_824,In_2213,In_1259);
xnor U825 (N_825,In_2834,In_4563);
and U826 (N_826,In_267,In_1273);
nand U827 (N_827,In_3551,In_2534);
and U828 (N_828,In_1476,In_962);
and U829 (N_829,In_153,In_2783);
and U830 (N_830,In_496,In_4899);
nand U831 (N_831,In_1211,In_867);
nor U832 (N_832,In_4908,In_2030);
nor U833 (N_833,In_566,In_1515);
nand U834 (N_834,In_461,In_1283);
nor U835 (N_835,In_2602,N_402);
and U836 (N_836,In_4242,In_389);
or U837 (N_837,In_1157,In_4474);
nor U838 (N_838,In_2063,In_3024);
nand U839 (N_839,In_1729,In_3700);
and U840 (N_840,In_1855,In_1070);
or U841 (N_841,In_1519,In_1923);
nor U842 (N_842,In_3774,In_129);
nand U843 (N_843,In_2820,In_1665);
nand U844 (N_844,In_2991,In_4027);
and U845 (N_845,In_4422,In_3920);
xnor U846 (N_846,In_4151,N_44);
xnor U847 (N_847,N_2,In_4324);
nor U848 (N_848,In_3692,In_2927);
xnor U849 (N_849,In_3915,In_1530);
nand U850 (N_850,In_2235,In_534);
nor U851 (N_851,In_1803,In_3741);
or U852 (N_852,In_1324,In_1712);
xor U853 (N_853,In_1972,In_4206);
or U854 (N_854,In_2180,In_2079);
nor U855 (N_855,In_1507,In_1801);
nand U856 (N_856,In_1762,In_545);
nand U857 (N_857,In_1781,In_675);
nor U858 (N_858,In_1879,In_1579);
and U859 (N_859,In_3759,In_3068);
and U860 (N_860,In_2565,In_3207);
or U861 (N_861,In_3642,In_3166);
and U862 (N_862,In_836,In_3824);
nor U863 (N_863,In_4889,In_2637);
or U864 (N_864,N_384,In_2692);
nand U865 (N_865,In_371,In_4639);
nor U866 (N_866,In_93,In_2303);
or U867 (N_867,In_2189,In_4559);
and U868 (N_868,In_2699,In_1017);
nand U869 (N_869,In_1079,In_2654);
and U870 (N_870,In_3776,In_4960);
or U871 (N_871,In_1910,In_1678);
or U872 (N_872,In_4566,In_704);
and U873 (N_873,In_4104,In_1660);
or U874 (N_874,In_2586,In_1572);
nand U875 (N_875,In_735,In_434);
and U876 (N_876,In_3708,N_114);
nor U877 (N_877,In_4842,In_2936);
and U878 (N_878,In_2591,In_4113);
or U879 (N_879,In_4315,In_3419);
xor U880 (N_880,In_3107,In_4726);
nor U881 (N_881,In_2667,In_2426);
nand U882 (N_882,In_4432,In_3086);
or U883 (N_883,In_1418,In_4379);
xor U884 (N_884,In_3255,In_3839);
or U885 (N_885,In_4857,In_2283);
and U886 (N_886,In_1806,In_2345);
nor U887 (N_887,In_588,In_4388);
or U888 (N_888,In_768,In_695);
nand U889 (N_889,In_31,In_4822);
nand U890 (N_890,In_3499,In_812);
nor U891 (N_891,N_135,In_942);
and U892 (N_892,In_1825,In_600);
nand U893 (N_893,N_479,In_407);
nor U894 (N_894,In_2088,In_1419);
or U895 (N_895,N_399,In_3239);
and U896 (N_896,N_492,In_4291);
nand U897 (N_897,In_284,In_340);
and U898 (N_898,In_4128,In_2824);
nand U899 (N_899,In_3550,In_1404);
nor U900 (N_900,In_897,In_3084);
xnor U901 (N_901,In_3047,In_4486);
and U902 (N_902,In_2501,In_2358);
nor U903 (N_903,In_4620,In_737);
and U904 (N_904,In_1261,In_4051);
nor U905 (N_905,In_1492,In_656);
and U906 (N_906,In_4499,In_3782);
or U907 (N_907,In_2663,In_539);
nor U908 (N_908,In_3349,In_2226);
xnor U909 (N_909,In_4216,In_1617);
nor U910 (N_910,In_2286,In_3971);
or U911 (N_911,In_2879,In_1214);
and U912 (N_912,In_3828,N_25);
or U913 (N_913,In_3541,In_4230);
nand U914 (N_914,In_2868,In_1380);
nor U915 (N_915,In_4801,In_4844);
nor U916 (N_916,In_3203,In_2904);
or U917 (N_917,N_243,In_2042);
nor U918 (N_918,In_4312,In_2255);
nor U919 (N_919,In_3711,In_3553);
or U920 (N_920,In_138,In_2509);
and U921 (N_921,In_3027,In_3090);
or U922 (N_922,In_4602,In_951);
nand U923 (N_923,N_443,N_131);
or U924 (N_924,In_2616,In_1136);
and U925 (N_925,In_4059,In_1483);
nand U926 (N_926,In_4441,In_1692);
or U927 (N_927,In_1673,In_1952);
and U928 (N_928,N_192,In_198);
xor U929 (N_929,In_3548,In_1043);
or U930 (N_930,In_3169,In_717);
and U931 (N_931,In_2009,In_3648);
or U932 (N_932,In_1618,In_1740);
xor U933 (N_933,In_2946,In_4703);
and U934 (N_934,In_3679,In_537);
nor U935 (N_935,In_842,In_2313);
nand U936 (N_936,In_1606,In_889);
nand U937 (N_937,In_1613,In_4335);
nand U938 (N_938,In_2273,In_722);
or U939 (N_939,N_226,N_478);
and U940 (N_940,In_3205,In_4644);
and U941 (N_941,In_2443,N_0);
nand U942 (N_942,In_1629,In_2650);
nor U943 (N_943,In_312,In_4266);
nor U944 (N_944,In_4231,In_4570);
or U945 (N_945,In_574,In_1783);
xor U946 (N_946,In_52,In_762);
nor U947 (N_947,In_2894,N_5);
and U948 (N_948,In_958,N_454);
nand U949 (N_949,In_355,In_4550);
nor U950 (N_950,N_260,N_47);
or U951 (N_951,In_1725,In_782);
nor U952 (N_952,N_432,In_2023);
and U953 (N_953,In_4549,In_2762);
nand U954 (N_954,In_3630,In_4117);
and U955 (N_955,In_1298,In_98);
and U956 (N_956,In_2639,In_2996);
or U957 (N_957,In_4661,In_2364);
xnor U958 (N_958,In_777,In_2149);
nand U959 (N_959,In_4977,In_3518);
and U960 (N_960,In_2126,In_2498);
nand U961 (N_961,In_2535,In_1466);
nor U962 (N_962,In_2994,In_3809);
xnor U963 (N_963,In_670,In_736);
nor U964 (N_964,In_3483,In_813);
or U965 (N_965,In_2028,In_847);
or U966 (N_966,In_3332,In_4598);
xor U967 (N_967,In_672,In_3683);
and U968 (N_968,In_3021,In_3674);
nand U969 (N_969,In_3296,In_2567);
and U970 (N_970,In_4194,In_2203);
or U971 (N_971,In_257,In_2350);
and U972 (N_972,In_1571,In_2370);
nor U973 (N_973,In_4517,In_1718);
and U974 (N_974,In_3214,In_1231);
or U975 (N_975,In_700,In_451);
nor U976 (N_976,In_1778,In_791);
nor U977 (N_977,In_2918,In_4547);
and U978 (N_978,In_4426,In_1434);
nor U979 (N_979,In_3303,In_975);
or U980 (N_980,In_2517,In_3136);
nor U981 (N_981,In_2438,N_380);
xnor U982 (N_982,In_2950,In_1351);
and U983 (N_983,In_1593,In_213);
or U984 (N_984,In_1175,In_3984);
nand U985 (N_985,N_386,In_2473);
nand U986 (N_986,In_1319,In_1835);
or U987 (N_987,In_452,In_1597);
nand U988 (N_988,In_1644,In_1384);
nand U989 (N_989,N_8,In_4985);
nand U990 (N_990,In_4973,In_2207);
nand U991 (N_991,In_2323,In_4067);
and U992 (N_992,In_1232,In_2527);
and U993 (N_993,In_861,In_4988);
and U994 (N_994,In_1065,In_1640);
nor U995 (N_995,In_1212,In_3360);
nor U996 (N_996,In_294,In_3830);
or U997 (N_997,In_1833,In_3122);
or U998 (N_998,In_1129,In_1658);
xor U999 (N_999,In_4592,In_917);
xnor U1000 (N_1000,N_880,In_903);
nor U1001 (N_1001,In_3246,In_4530);
nor U1002 (N_1002,In_523,In_519);
and U1003 (N_1003,N_811,In_3208);
or U1004 (N_1004,In_159,In_2576);
nor U1005 (N_1005,In_4607,In_4969);
nand U1006 (N_1006,In_3813,In_2589);
xor U1007 (N_1007,In_4515,In_4089);
nor U1008 (N_1008,In_2274,N_222);
or U1009 (N_1009,In_4866,In_1268);
nor U1010 (N_1010,In_2400,In_515);
and U1011 (N_1011,In_2613,N_715);
nand U1012 (N_1012,In_2972,N_810);
nand U1013 (N_1013,In_3995,In_2594);
and U1014 (N_1014,In_3728,In_252);
or U1015 (N_1015,In_3885,In_3348);
or U1016 (N_1016,N_403,N_500);
nand U1017 (N_1017,In_3925,N_7);
and U1018 (N_1018,In_2506,In_3750);
or U1019 (N_1019,In_3376,In_45);
or U1020 (N_1020,N_885,N_297);
nand U1021 (N_1021,In_846,In_2697);
and U1022 (N_1022,In_642,N_430);
nor U1023 (N_1023,In_1922,In_3532);
and U1024 (N_1024,N_629,In_527);
and U1025 (N_1025,In_3962,In_2442);
nand U1026 (N_1026,In_1250,In_193);
nand U1027 (N_1027,In_1458,In_2944);
and U1028 (N_1028,N_305,In_2662);
or U1029 (N_1029,In_3658,In_4636);
and U1030 (N_1030,In_4093,N_136);
or U1031 (N_1031,N_12,N_608);
xor U1032 (N_1032,In_2665,In_4021);
and U1033 (N_1033,In_2634,N_283);
and U1034 (N_1034,N_50,In_428);
nand U1035 (N_1035,In_814,In_3979);
nor U1036 (N_1036,In_2725,In_3176);
nor U1037 (N_1037,In_703,In_1792);
or U1038 (N_1038,In_3586,In_1908);
nor U1039 (N_1039,In_4616,In_1896);
nand U1040 (N_1040,In_2952,In_109);
and U1041 (N_1041,In_4377,In_3631);
or U1042 (N_1042,In_1878,N_110);
and U1043 (N_1043,N_542,In_479);
or U1044 (N_1044,N_965,In_3993);
or U1045 (N_1045,N_758,In_4727);
nor U1046 (N_1046,In_708,N_476);
and U1047 (N_1047,In_183,N_928);
or U1048 (N_1048,In_720,In_938);
nor U1049 (N_1049,In_2340,In_4304);
and U1050 (N_1050,In_2775,In_886);
nor U1051 (N_1051,In_2138,N_704);
nand U1052 (N_1052,In_1750,In_3754);
and U1053 (N_1053,In_4271,In_4044);
and U1054 (N_1054,In_233,In_3910);
and U1055 (N_1055,N_609,N_588);
nor U1056 (N_1056,In_2886,In_3272);
nor U1057 (N_1057,N_691,In_1066);
nor U1058 (N_1058,In_2195,In_3044);
nand U1059 (N_1059,In_103,In_189);
and U1060 (N_1060,N_862,In_3651);
nand U1061 (N_1061,In_3281,In_3387);
xnor U1062 (N_1062,N_164,In_2373);
and U1063 (N_1063,In_1685,N_547);
and U1064 (N_1064,N_183,In_3263);
or U1065 (N_1065,In_2098,N_589);
xor U1066 (N_1066,In_2660,N_543);
nor U1067 (N_1067,In_2845,In_1141);
or U1068 (N_1068,In_3458,In_3726);
nor U1069 (N_1069,In_4195,In_2593);
or U1070 (N_1070,In_1160,In_136);
nor U1071 (N_1071,In_4100,In_890);
nor U1072 (N_1072,In_1537,N_481);
nor U1073 (N_1073,In_1308,In_892);
or U1074 (N_1074,In_4940,In_4914);
nor U1075 (N_1075,In_1736,In_1188);
and U1076 (N_1076,N_791,In_529);
or U1077 (N_1077,N_869,N_278);
nor U1078 (N_1078,N_669,In_3494);
or U1079 (N_1079,In_4939,In_4293);
and U1080 (N_1080,N_565,In_3645);
nand U1081 (N_1081,In_4034,In_4412);
and U1082 (N_1082,In_1201,In_1754);
and U1083 (N_1083,N_622,In_2896);
and U1084 (N_1084,In_1967,N_325);
nor U1085 (N_1085,In_2389,In_77);
nand U1086 (N_1086,In_357,In_380);
and U1087 (N_1087,In_343,In_135);
nor U1088 (N_1088,In_89,N_567);
xor U1089 (N_1089,In_2058,In_4713);
and U1090 (N_1090,N_477,In_2572);
xor U1091 (N_1091,N_505,In_1089);
nand U1092 (N_1092,In_4783,In_204);
nand U1093 (N_1093,In_4540,In_2333);
nand U1094 (N_1094,In_1041,In_1251);
nor U1095 (N_1095,In_2666,In_2838);
or U1096 (N_1096,In_3396,In_551);
or U1097 (N_1097,In_796,In_4090);
nand U1098 (N_1098,N_30,In_4357);
nand U1099 (N_1099,In_2020,In_1799);
nor U1100 (N_1100,In_1881,N_605);
or U1101 (N_1101,In_2737,In_3861);
or U1102 (N_1102,In_3412,In_1140);
nand U1103 (N_1103,In_4055,In_1988);
and U1104 (N_1104,In_4958,In_74);
nor U1105 (N_1105,N_659,N_332);
and U1106 (N_1106,N_329,In_400);
nor U1107 (N_1107,In_3058,In_650);
or U1108 (N_1108,In_4748,In_493);
nand U1109 (N_1109,In_393,In_2044);
nor U1110 (N_1110,In_1289,In_4780);
or U1111 (N_1111,In_2163,In_254);
and U1112 (N_1112,In_766,In_3918);
nand U1113 (N_1113,In_932,N_51);
nand U1114 (N_1114,In_3899,In_2659);
nor U1115 (N_1115,In_1924,In_1377);
nor U1116 (N_1116,N_654,N_530);
nor U1117 (N_1117,In_4827,In_2627);
or U1118 (N_1118,In_4245,In_2036);
nand U1119 (N_1119,N_798,In_1198);
or U1120 (N_1120,In_3906,In_718);
or U1121 (N_1121,In_4127,N_650);
nor U1122 (N_1122,In_3689,In_4836);
or U1123 (N_1123,In_3507,In_772);
nand U1124 (N_1124,In_3896,In_1975);
xnor U1125 (N_1125,N_160,In_481);
nand U1126 (N_1126,In_3953,In_2691);
nand U1127 (N_1127,N_118,In_2959);
or U1128 (N_1128,In_2544,N_894);
or U1129 (N_1129,In_1714,N_75);
nor U1130 (N_1130,In_3323,In_598);
nand U1131 (N_1131,In_1859,In_1760);
nor U1132 (N_1132,In_4429,In_2212);
and U1133 (N_1133,In_4937,N_556);
xnor U1134 (N_1134,N_952,In_413);
nor U1135 (N_1135,In_117,In_2012);
nor U1136 (N_1136,In_4112,In_2397);
or U1137 (N_1137,In_408,In_2413);
and U1138 (N_1138,N_835,In_4865);
or U1139 (N_1139,In_2471,N_122);
and U1140 (N_1140,In_104,N_70);
nor U1141 (N_1141,In_3299,N_308);
nor U1142 (N_1142,In_484,In_306);
and U1143 (N_1143,In_1777,In_1939);
xor U1144 (N_1144,N_921,In_94);
xnor U1145 (N_1145,In_337,In_467);
nor U1146 (N_1146,In_4625,In_2916);
or U1147 (N_1147,In_255,N_717);
nand U1148 (N_1148,In_4477,In_4496);
or U1149 (N_1149,In_1797,In_612);
and U1150 (N_1150,In_4893,N_637);
and U1151 (N_1151,In_1538,N_857);
nand U1152 (N_1152,In_640,In_1612);
or U1153 (N_1153,In_521,In_4161);
xor U1154 (N_1154,In_1020,In_3337);
nand U1155 (N_1155,N_672,N_321);
nor U1156 (N_1156,In_3399,In_160);
and U1157 (N_1157,In_1987,In_24);
or U1158 (N_1158,In_4569,In_4389);
nand U1159 (N_1159,In_1887,In_1257);
and U1160 (N_1160,In_4045,In_1445);
nand U1161 (N_1161,N_944,N_141);
nor U1162 (N_1162,In_2194,In_34);
xor U1163 (N_1163,N_453,In_1804);
or U1164 (N_1164,In_3684,In_2746);
nor U1165 (N_1165,In_99,N_126);
nand U1166 (N_1166,In_2632,In_1931);
or U1167 (N_1167,In_1080,In_3837);
nor U1168 (N_1168,In_1387,In_4016);
and U1169 (N_1169,In_2007,In_1745);
nand U1170 (N_1170,In_725,In_448);
xnor U1171 (N_1171,In_1374,In_4075);
and U1172 (N_1172,N_379,In_429);
nand U1173 (N_1173,N_489,In_3638);
nand U1174 (N_1174,N_724,In_844);
or U1175 (N_1175,N_249,In_2638);
nor U1176 (N_1176,In_1594,N_223);
nand U1177 (N_1177,In_1854,In_4778);
or U1178 (N_1178,N_48,In_1234);
or U1179 (N_1179,In_887,In_2412);
xor U1180 (N_1180,N_550,In_1264);
or U1181 (N_1181,In_1696,N_587);
nand U1182 (N_1182,In_563,In_216);
and U1183 (N_1183,In_1635,In_69);
nand U1184 (N_1184,In_3067,In_3191);
xnor U1185 (N_1185,In_3663,In_4688);
and U1186 (N_1186,N_179,N_496);
nor U1187 (N_1187,In_4680,N_546);
nor U1188 (N_1188,In_1817,N_416);
nand U1189 (N_1189,In_3676,In_4054);
and U1190 (N_1190,In_3864,In_1895);
or U1191 (N_1191,In_1637,In_2958);
or U1192 (N_1192,In_4867,N_979);
or U1193 (N_1193,In_3478,In_2636);
and U1194 (N_1194,In_1992,N_978);
nor U1195 (N_1195,In_3871,In_2752);
or U1196 (N_1196,N_840,In_4705);
nor U1197 (N_1197,In_4328,In_2429);
nand U1198 (N_1198,In_2732,In_245);
and U1199 (N_1199,N_346,In_390);
nor U1200 (N_1200,In_3702,N_357);
and U1201 (N_1201,N_670,In_1621);
nand U1202 (N_1202,In_4878,In_370);
xnor U1203 (N_1203,In_3223,In_3153);
or U1204 (N_1204,N_299,N_145);
xnor U1205 (N_1205,In_1576,In_3368);
or U1206 (N_1206,In_2724,In_325);
or U1207 (N_1207,N_743,In_4701);
or U1208 (N_1208,In_783,In_2960);
xnor U1209 (N_1209,In_3973,N_827);
or U1210 (N_1210,In_3960,N_864);
nor U1211 (N_1211,In_4204,In_497);
and U1212 (N_1212,In_3398,In_3598);
nor U1213 (N_1213,N_382,In_2872);
or U1214 (N_1214,In_1532,In_4910);
and U1215 (N_1215,In_1274,In_3567);
nor U1216 (N_1216,In_2218,In_4955);
nand U1217 (N_1217,N_316,In_4874);
nor U1218 (N_1218,In_2953,In_1691);
xor U1219 (N_1219,N_731,In_2482);
or U1220 (N_1220,N_43,In_609);
and U1221 (N_1221,In_730,In_2162);
or U1222 (N_1222,In_4374,In_2150);
nor U1223 (N_1223,In_4888,In_1513);
or U1224 (N_1224,In_4796,In_1356);
nand U1225 (N_1225,N_739,In_2132);
or U1226 (N_1226,In_619,In_3071);
nor U1227 (N_1227,In_2363,In_823);
or U1228 (N_1228,In_4728,In_2321);
or U1229 (N_1229,In_4318,N_331);
and U1230 (N_1230,N_711,In_2893);
and U1231 (N_1231,In_4488,In_2856);
nor U1232 (N_1232,In_4522,N_538);
and U1233 (N_1233,In_1381,N_581);
or U1234 (N_1234,N_747,In_2799);
or U1235 (N_1235,In_2431,N_897);
nor U1236 (N_1236,In_2202,N_778);
or U1237 (N_1237,In_203,In_3344);
nand U1238 (N_1238,In_899,N_832);
nand U1239 (N_1239,In_3964,N_60);
nand U1240 (N_1240,In_4099,In_3632);
nor U1241 (N_1241,In_2792,In_4589);
xnor U1242 (N_1242,In_2962,In_1058);
nor U1243 (N_1243,In_1392,In_191);
nand U1244 (N_1244,In_1149,In_2577);
and U1245 (N_1245,In_4980,In_2774);
nand U1246 (N_1246,N_583,In_3686);
nand U1247 (N_1247,In_4521,In_1053);
nand U1248 (N_1248,N_211,In_3077);
nor U1249 (N_1249,In_1332,In_57);
and U1250 (N_1250,In_1919,In_4462);
or U1251 (N_1251,In_3735,In_3106);
and U1252 (N_1252,N_27,N_948);
nor U1253 (N_1253,In_4126,N_915);
nor U1254 (N_1254,N_170,In_4715);
and U1255 (N_1255,In_4155,In_4053);
nor U1256 (N_1256,N_400,In_2885);
or U1257 (N_1257,In_3639,In_507);
xor U1258 (N_1258,In_1648,In_1790);
and U1259 (N_1259,In_205,In_3073);
xor U1260 (N_1260,In_4671,In_2656);
and U1261 (N_1261,In_2107,In_4815);
and U1262 (N_1262,In_44,In_2362);
nand U1263 (N_1263,In_3216,In_2747);
or U1264 (N_1264,N_815,N_537);
nor U1265 (N_1265,In_2919,N_28);
or U1266 (N_1266,In_3426,N_552);
nor U1267 (N_1267,N_232,N_956);
or U1268 (N_1268,In_1278,In_748);
and U1269 (N_1269,In_1498,N_312);
or U1270 (N_1270,N_236,N_941);
or U1271 (N_1271,N_29,In_4816);
nor U1272 (N_1272,In_2968,In_4393);
xnor U1273 (N_1273,In_4336,In_816);
or U1274 (N_1274,N_504,In_4799);
and U1275 (N_1275,N_177,In_1085);
and U1276 (N_1276,In_1540,In_76);
and U1277 (N_1277,N_889,N_133);
nor U1278 (N_1278,In_162,N_674);
nand U1279 (N_1279,N_826,In_4754);
and U1280 (N_1280,In_4060,In_350);
and U1281 (N_1281,N_819,N_718);
and U1282 (N_1282,N_660,In_4069);
or U1283 (N_1283,In_1313,In_3343);
nand U1284 (N_1284,N_759,In_3465);
nor U1285 (N_1285,In_4239,In_4723);
xnor U1286 (N_1286,In_1411,In_4403);
nor U1287 (N_1287,In_1130,N_790);
nand U1288 (N_1288,In_3986,In_3132);
or U1289 (N_1289,In_4481,In_240);
xnor U1290 (N_1290,In_297,In_1311);
nand U1291 (N_1291,In_43,In_3746);
or U1292 (N_1292,N_18,N_792);
or U1293 (N_1293,In_1475,In_10);
nor U1294 (N_1294,In_655,In_1469);
nand U1295 (N_1295,In_957,N_855);
or U1296 (N_1296,In_3167,N_176);
and U1297 (N_1297,In_2200,In_1243);
nand U1298 (N_1298,In_773,In_1015);
nor U1299 (N_1299,In_3945,N_173);
nor U1300 (N_1300,N_515,N_877);
or U1301 (N_1301,In_4716,In_508);
and U1302 (N_1302,In_2024,N_483);
or U1303 (N_1303,In_3816,In_2976);
nor U1304 (N_1304,N_377,In_3560);
and U1305 (N_1305,In_3887,In_3363);
and U1306 (N_1306,In_4213,In_3011);
nor U1307 (N_1307,In_1772,N_982);
and U1308 (N_1308,In_3146,In_373);
nand U1309 (N_1309,In_3339,In_1461);
and U1310 (N_1310,In_757,N_457);
or U1311 (N_1311,N_777,In_3078);
nand U1312 (N_1312,In_4424,In_4461);
nor U1313 (N_1313,In_2983,N_590);
xnor U1314 (N_1314,N_927,In_808);
and U1315 (N_1315,In_3846,In_1307);
nand U1316 (N_1316,In_914,N_286);
nand U1317 (N_1317,In_2512,N_825);
nand U1318 (N_1318,In_787,In_4721);
and U1319 (N_1319,In_4719,In_211);
and U1320 (N_1320,In_4736,N_766);
nor U1321 (N_1321,In_4830,In_1290);
nor U1322 (N_1322,In_3504,N_441);
nor U1323 (N_1323,In_3584,In_978);
xor U1324 (N_1324,In_572,In_3892);
nand U1325 (N_1325,In_3858,In_532);
and U1326 (N_1326,In_1518,In_2898);
or U1327 (N_1327,In_1209,In_918);
and U1328 (N_1328,In_3992,In_2551);
and U1329 (N_1329,In_4285,In_1401);
and U1330 (N_1330,In_55,In_3080);
nand U1331 (N_1331,In_1845,In_3572);
nand U1332 (N_1332,In_3301,N_866);
nor U1333 (N_1333,In_3052,In_4346);
and U1334 (N_1334,In_4943,In_4350);
and U1335 (N_1335,In_4139,In_3407);
or U1336 (N_1336,In_3793,N_69);
and U1337 (N_1337,In_2742,In_1564);
or U1338 (N_1338,N_793,In_207);
or U1339 (N_1339,N_961,In_1044);
and U1340 (N_1340,In_1703,In_3473);
xor U1341 (N_1341,In_178,N_706);
nand U1342 (N_1342,In_3453,In_676);
nand U1343 (N_1343,In_793,In_3912);
nand U1344 (N_1344,In_2985,In_2910);
xor U1345 (N_1345,In_2469,In_2588);
or U1346 (N_1346,N_72,N_740);
and U1347 (N_1347,In_3442,In_2878);
nand U1348 (N_1348,In_3613,In_2294);
nand U1349 (N_1349,In_4858,In_2411);
and U1350 (N_1350,N_279,In_486);
and U1351 (N_1351,N_719,In_3690);
xnor U1352 (N_1352,In_405,In_4851);
and U1353 (N_1353,In_298,In_3141);
nor U1354 (N_1354,N_404,N_770);
or U1355 (N_1355,In_1226,In_2859);
xnor U1356 (N_1356,N_115,In_2346);
nand U1357 (N_1357,N_314,In_2888);
nor U1358 (N_1358,In_168,In_4261);
or U1359 (N_1359,In_3050,N_765);
nand U1360 (N_1360,In_2728,In_78);
and U1361 (N_1361,N_705,In_4950);
and U1362 (N_1362,In_794,N_698);
nand U1363 (N_1363,In_4455,In_2349);
xor U1364 (N_1364,In_1413,In_2628);
nand U1365 (N_1365,In_4533,In_4459);
and U1366 (N_1366,In_4601,In_1116);
nand U1367 (N_1367,In_3821,In_1751);
or U1368 (N_1368,In_450,N_491);
or U1369 (N_1369,In_4435,In_1748);
or U1370 (N_1370,In_4541,In_570);
nand U1371 (N_1371,N_690,In_4752);
nand U1372 (N_1372,N_560,In_1679);
nor U1373 (N_1373,In_1301,In_4632);
nand U1374 (N_1374,In_3482,In_1039);
nand U1375 (N_1375,In_1641,In_3849);
nor U1376 (N_1376,N_807,In_2830);
nor U1377 (N_1377,In_862,In_1776);
or U1378 (N_1378,In_2217,In_440);
and U1379 (N_1379,In_2081,In_3293);
nand U1380 (N_1380,N_597,In_2295);
nor U1381 (N_1381,N_92,In_2254);
or U1382 (N_1382,In_2269,In_2324);
nand U1383 (N_1383,N_241,In_1920);
or U1384 (N_1384,In_3247,N_562);
and U1385 (N_1385,In_528,In_967);
nand U1386 (N_1386,In_3706,N_37);
xnor U1387 (N_1387,In_4064,In_1497);
nand U1388 (N_1388,In_3790,In_4358);
nor U1389 (N_1389,N_549,In_2858);
nand U1390 (N_1390,In_4174,In_3669);
or U1391 (N_1391,N_32,N_344);
nand U1392 (N_1392,N_974,N_943);
xor U1393 (N_1393,In_1076,In_1582);
xor U1394 (N_1394,In_2168,In_3219);
or U1395 (N_1395,N_370,In_2041);
nor U1396 (N_1396,N_464,In_3320);
xnor U1397 (N_1397,In_1276,In_3447);
or U1398 (N_1398,In_3949,In_902);
xnor U1399 (N_1399,In_1650,In_805);
nand U1400 (N_1400,In_2570,In_1587);
and U1401 (N_1401,In_130,In_3808);
nand U1402 (N_1402,N_262,In_915);
and U1403 (N_1403,In_2934,In_1222);
and U1404 (N_1404,In_2681,In_3151);
nor U1405 (N_1405,In_4941,N_112);
nor U1406 (N_1406,N_914,In_3597);
nor U1407 (N_1407,N_800,In_2147);
or U1408 (N_1408,In_137,N_929);
and U1409 (N_1409,In_3079,In_2630);
or U1410 (N_1410,In_1327,In_1688);
nor U1411 (N_1411,N_679,In_4106);
nor U1412 (N_1412,N_572,N_742);
xor U1413 (N_1413,N_62,In_3623);
nor U1414 (N_1414,In_38,In_3297);
or U1415 (N_1415,In_4967,In_4087);
nor U1416 (N_1416,N_153,N_699);
nor U1417 (N_1417,N_300,N_20);
nand U1418 (N_1418,In_3375,In_606);
nor U1419 (N_1419,In_2836,N_217);
nor U1420 (N_1420,N_317,N_687);
or U1421 (N_1421,In_2496,In_303);
nor U1422 (N_1422,In_3212,In_4876);
and U1423 (N_1423,In_120,In_4537);
nand U1424 (N_1424,In_4005,In_4040);
nand U1425 (N_1425,In_1917,In_1585);
nor U1426 (N_1426,In_2434,In_1639);
nor U1427 (N_1427,In_91,In_1785);
nand U1428 (N_1428,In_2862,In_4061);
and U1429 (N_1429,In_505,N_465);
nor U1430 (N_1430,In_4672,In_2587);
nor U1431 (N_1431,In_2329,In_3418);
nand U1432 (N_1432,In_3905,In_1350);
nand U1433 (N_1433,In_4235,In_2559);
and U1434 (N_1434,In_3187,In_2135);
nand U1435 (N_1435,N_119,In_2707);
nor U1436 (N_1436,In_392,In_2368);
and U1437 (N_1437,In_2939,In_1427);
xor U1438 (N_1438,In_1367,In_3811);
nor U1439 (N_1439,In_709,In_1127);
nand U1440 (N_1440,In_2704,In_4082);
nor U1441 (N_1441,In_3149,In_4760);
nand U1442 (N_1442,In_3108,In_3116);
or U1443 (N_1443,In_657,In_603);
or U1444 (N_1444,In_158,In_80);
nand U1445 (N_1445,In_1773,In_3854);
and U1446 (N_1446,In_4696,In_1682);
nand U1447 (N_1447,In_2243,In_1204);
nor U1448 (N_1448,In_4399,In_147);
nand U1449 (N_1449,In_2909,In_1511);
or U1450 (N_1450,In_928,N_517);
nand U1451 (N_1451,In_2062,N_182);
or U1452 (N_1452,In_323,In_3013);
or U1453 (N_1453,In_2833,In_584);
or U1454 (N_1454,In_3455,N_159);
nand U1455 (N_1455,In_36,In_1752);
or U1456 (N_1456,In_2523,In_1808);
and U1457 (N_1457,N_892,In_4849);
nor U1458 (N_1458,In_1543,N_154);
or U1459 (N_1459,In_682,N_615);
and U1460 (N_1460,N_522,In_3433);
and U1461 (N_1461,In_568,In_1559);
xor U1462 (N_1462,In_3826,In_3667);
nand U1463 (N_1463,N_431,In_2067);
or U1464 (N_1464,In_264,In_3917);
or U1465 (N_1465,In_4332,In_3582);
xor U1466 (N_1466,N_712,In_4337);
or U1467 (N_1467,In_4892,N_584);
and U1468 (N_1468,In_4560,In_2826);
nand U1469 (N_1469,In_1481,In_42);
and U1470 (N_1470,N_853,In_2171);
and U1471 (N_1471,In_2417,In_1819);
nor U1472 (N_1472,In_2229,In_1528);
nor U1473 (N_1473,In_2676,In_4989);
or U1474 (N_1474,In_1146,In_3196);
or U1475 (N_1475,In_1812,In_2348);
nand U1476 (N_1476,N_306,In_2116);
xor U1477 (N_1477,In_3324,In_278);
xor U1478 (N_1478,N_445,N_918);
nand U1479 (N_1479,N_455,In_558);
nand U1480 (N_1480,In_1503,In_1771);
and U1481 (N_1481,N_882,In_504);
xnor U1482 (N_1482,In_4966,N_697);
and U1483 (N_1483,In_4491,In_3232);
nor U1484 (N_1484,In_1698,N_566);
nand U1485 (N_1485,In_2941,In_1763);
and U1486 (N_1486,N_303,N_801);
nor U1487 (N_1487,In_981,In_1277);
or U1488 (N_1488,N_794,In_1061);
xor U1489 (N_1489,In_2211,N_591);
and U1490 (N_1490,In_3909,In_4921);
nand U1491 (N_1491,N_269,In_269);
and U1492 (N_1492,N_64,In_2921);
xnor U1493 (N_1493,In_2625,In_1788);
xnor U1494 (N_1494,N_959,In_4848);
xor U1495 (N_1495,In_4553,In_3353);
nand U1496 (N_1496,N_518,In_4191);
or U1497 (N_1497,N_88,N_161);
xnor U1498 (N_1498,In_2101,In_2127);
nor U1499 (N_1499,In_3534,N_639);
nor U1500 (N_1500,In_1945,In_2817);
nand U1501 (N_1501,In_1131,In_1557);
nor U1502 (N_1502,N_1467,N_59);
nor U1503 (N_1503,N_665,In_4224);
nor U1504 (N_1504,In_3038,In_4092);
nand U1505 (N_1505,In_2111,In_3634);
xor U1506 (N_1506,In_4454,In_2296);
xnor U1507 (N_1507,N_438,N_1430);
nor U1508 (N_1508,In_11,N_833);
nand U1509 (N_1509,In_2139,In_2651);
and U1510 (N_1510,N_87,N_1426);
and U1511 (N_1511,In_3999,In_202);
nand U1512 (N_1512,In_494,N_830);
xor U1513 (N_1513,In_743,N_1355);
nand U1514 (N_1514,In_1584,In_4931);
and U1515 (N_1515,In_2657,In_604);
nand U1516 (N_1516,In_1164,In_3641);
nor U1517 (N_1517,In_4098,N_1429);
nor U1518 (N_1518,In_3431,N_1063);
and U1519 (N_1519,In_857,N_1365);
or U1520 (N_1520,N_1062,In_597);
or U1521 (N_1521,N_1142,In_3180);
nand U1522 (N_1522,In_2526,N_763);
xnor U1523 (N_1523,In_3308,In_1661);
nor U1524 (N_1524,In_775,N_452);
and U1525 (N_1525,N_1084,In_602);
nand U1526 (N_1526,N_939,N_227);
nand U1527 (N_1527,N_646,N_1267);
nand U1528 (N_1528,In_3275,In_4603);
nand U1529 (N_1529,In_1955,In_941);
and U1530 (N_1530,N_799,In_1395);
and U1531 (N_1531,In_4391,In_4762);
or U1532 (N_1532,In_4202,In_2242);
nor U1533 (N_1533,N_1381,In_3193);
and U1534 (N_1534,In_3944,N_1330);
nor U1535 (N_1535,In_2022,In_3647);
and U1536 (N_1536,In_3055,In_4036);
and U1537 (N_1537,In_2112,In_4809);
nor U1538 (N_1538,In_1520,In_4585);
nor U1539 (N_1539,N_926,In_2187);
nor U1540 (N_1540,In_4476,In_3787);
nor U1541 (N_1541,N_636,In_3954);
or U1542 (N_1542,In_1173,In_1134);
and U1543 (N_1543,N_228,In_2832);
nand U1544 (N_1544,N_632,In_395);
or U1545 (N_1545,N_534,In_3346);
or U1546 (N_1546,In_1161,In_281);
nand U1547 (N_1547,In_3827,In_2773);
and U1548 (N_1548,In_2635,In_2289);
and U1549 (N_1549,In_840,In_12);
xor U1550 (N_1550,In_1974,In_1031);
and U1551 (N_1551,In_3443,N_1274);
and U1552 (N_1552,In_3655,In_3778);
nor U1553 (N_1553,N_356,In_4057);
nor U1554 (N_1554,In_3389,In_4765);
nand U1555 (N_1555,In_1733,In_1929);
or U1556 (N_1556,N_355,In_2937);
or U1557 (N_1557,In_4428,In_4580);
or U1558 (N_1558,In_2311,In_691);
nand U1559 (N_1559,N_1037,In_2679);
nor U1560 (N_1560,In_541,In_293);
nand U1561 (N_1561,N_1030,In_960);
and U1562 (N_1562,In_3775,In_2814);
and U1563 (N_1563,In_164,In_2209);
xor U1564 (N_1564,N_1017,N_847);
xor U1565 (N_1565,In_2564,In_4953);
or U1566 (N_1566,In_4298,In_3626);
nand U1567 (N_1567,In_54,N_1372);
or U1568 (N_1568,N_41,In_3636);
nor U1569 (N_1569,In_1728,N_1145);
and U1570 (N_1570,In_4687,In_1386);
nor U1571 (N_1571,In_265,In_4431);
and U1572 (N_1572,In_2173,N_996);
nor U1573 (N_1573,In_385,N_268);
nor U1574 (N_1574,In_3393,N_510);
or U1575 (N_1575,In_3178,N_1285);
nand U1576 (N_1576,In_2259,N_364);
nand U1577 (N_1577,In_251,In_1901);
and U1578 (N_1578,In_4818,N_375);
and U1579 (N_1579,N_1471,In_610);
nor U1580 (N_1580,N_1247,N_6);
or U1581 (N_1581,In_3262,In_2011);
or U1582 (N_1582,N_206,In_788);
and U1583 (N_1583,In_2843,N_1048);
nor U1584 (N_1584,N_99,In_2841);
or U1585 (N_1585,N_1415,In_3712);
or U1586 (N_1586,In_1385,In_2618);
and U1587 (N_1587,In_1372,In_1105);
nor U1588 (N_1588,In_3287,In_3306);
or U1589 (N_1589,In_2481,In_1969);
nor U1590 (N_1590,In_2344,In_620);
xnor U1591 (N_1591,In_4654,In_2220);
nand U1592 (N_1592,N_1302,In_1019);
nor U1593 (N_1593,In_3673,N_797);
and U1594 (N_1594,N_1451,N_319);
and U1595 (N_1595,In_88,In_1398);
or U1596 (N_1596,In_3404,In_1457);
nand U1597 (N_1597,In_4573,N_1173);
and U1598 (N_1598,In_1889,N_508);
or U1599 (N_1599,In_4342,In_3254);
xnor U1600 (N_1600,In_4417,N_94);
nor U1601 (N_1601,N_749,N_374);
nand U1602 (N_1602,N_401,In_2280);
nand U1603 (N_1603,In_2673,In_4003);
xor U1604 (N_1604,In_4018,In_3748);
and U1605 (N_1605,In_4981,In_4511);
nor U1606 (N_1606,N_848,In_1734);
nor U1607 (N_1607,N_1153,In_421);
or U1608 (N_1608,In_4526,In_2475);
nor U1609 (N_1609,In_4220,In_3490);
xor U1610 (N_1610,In_2646,In_3411);
nand U1611 (N_1611,In_3985,In_2519);
nor U1612 (N_1612,In_2491,In_4062);
nand U1613 (N_1613,In_3980,N_251);
nor U1614 (N_1614,N_1368,In_4505);
or U1615 (N_1615,In_2678,In_3046);
xor U1616 (N_1616,In_225,N_422);
nor U1617 (N_1617,In_4872,In_2407);
or U1618 (N_1618,In_2533,In_2048);
and U1619 (N_1619,In_3937,In_3587);
xnor U1620 (N_1620,In_291,In_4739);
nand U1621 (N_1621,In_2339,In_438);
and U1622 (N_1622,In_59,In_3415);
nand U1623 (N_1623,In_879,N_1440);
or U1624 (N_1624,In_4629,In_4770);
nand U1625 (N_1625,In_2153,N_787);
and U1626 (N_1626,In_4385,In_753);
or U1627 (N_1627,In_321,In_1054);
and U1628 (N_1628,N_708,N_1271);
or U1629 (N_1629,N_1016,In_4278);
nand U1630 (N_1630,In_491,N_548);
and U1631 (N_1631,N_388,N_773);
and U1632 (N_1632,In_3251,N_352);
and U1633 (N_1633,In_3635,N_872);
and U1634 (N_1634,In_4766,N_1449);
nand U1635 (N_1635,In_649,N_1251);
or U1636 (N_1636,In_3025,N_274);
and U1637 (N_1637,N_288,In_3543);
nand U1638 (N_1638,In_1424,N_459);
nand U1639 (N_1639,In_326,In_2992);
and U1640 (N_1640,In_1118,In_980);
nand U1641 (N_1641,N_999,In_552);
nand U1642 (N_1642,In_3298,In_4353);
nor U1643 (N_1643,In_2882,In_3173);
nor U1644 (N_1644,N_103,In_3926);
nand U1645 (N_1645,In_3701,In_3722);
or U1646 (N_1646,In_1242,N_751);
xor U1647 (N_1647,In_1490,N_1116);
nand U1648 (N_1648,N_1281,N_675);
nand U1649 (N_1649,N_157,In_2753);
nand U1650 (N_1650,In_1615,In_2425);
nand U1651 (N_1651,In_1460,N_1199);
or U1652 (N_1652,N_618,In_2499);
and U1653 (N_1653,In_939,N_1110);
or U1654 (N_1654,In_1994,In_1042);
or U1655 (N_1655,N_786,In_3884);
and U1656 (N_1656,In_2849,In_837);
and U1657 (N_1657,N_1079,In_1958);
nor U1658 (N_1658,In_4492,N_485);
and U1659 (N_1659,In_1408,In_4604);
and U1660 (N_1660,N_1184,In_2383);
and U1661 (N_1661,N_167,In_234);
nand U1662 (N_1662,In_415,In_697);
nand U1663 (N_1663,N_954,In_3439);
nand U1664 (N_1664,In_4869,N_333);
nand U1665 (N_1665,In_4175,N_554);
nand U1666 (N_1666,In_1339,In_3664);
nand U1667 (N_1667,In_4646,N_514);
xor U1668 (N_1668,In_3487,N_845);
and U1669 (N_1669,In_1331,In_356);
nand U1670 (N_1670,In_351,N_1495);
xnor U1671 (N_1671,N_466,In_654);
nand U1672 (N_1672,N_1160,In_3397);
and U1673 (N_1673,N_805,N_1323);
xor U1674 (N_1674,In_644,In_3696);
nor U1675 (N_1675,N_916,In_3276);
nand U1676 (N_1676,In_2920,In_3886);
nor U1677 (N_1677,In_2123,N_1064);
nand U1678 (N_1678,N_868,N_796);
and U1679 (N_1679,In_905,In_2124);
nor U1680 (N_1680,N_651,In_4507);
and U1681 (N_1681,In_751,In_1254);
nor U1682 (N_1682,N_713,N_140);
and U1683 (N_1683,In_1125,N_68);
nand U1684 (N_1684,N_1273,In_4097);
and U1685 (N_1685,N_456,In_557);
or U1686 (N_1686,N_390,In_4166);
nand U1687 (N_1687,In_607,N_202);
nor U1688 (N_1688,In_503,In_714);
nor U1689 (N_1689,N_1301,In_4343);
or U1690 (N_1690,In_3589,N_1039);
and U1691 (N_1691,N_863,In_904);
or U1692 (N_1692,In_3505,In_3);
nor U1693 (N_1693,N_343,In_3780);
and U1694 (N_1694,N_1335,N_1339);
and U1695 (N_1695,In_4495,In_4470);
nand U1696 (N_1696,In_2902,N_972);
nor U1697 (N_1697,In_712,In_75);
and U1698 (N_1698,N_412,In_4360);
or U1699 (N_1699,In_2720,In_3564);
and U1700 (N_1700,In_949,In_4433);
nor U1701 (N_1701,In_150,N_449);
nor U1702 (N_1702,In_1815,N_1259);
and U1703 (N_1703,In_4188,In_4596);
nand U1704 (N_1704,In_4962,In_2151);
nor U1705 (N_1705,N_482,N_1374);
and U1706 (N_1706,N_1045,In_1779);
or U1707 (N_1707,N_1375,N_1484);
or U1708 (N_1708,In_1083,In_4037);
xor U1709 (N_1709,In_1590,In_2803);
nand U1710 (N_1710,In_4352,N_568);
nor U1711 (N_1711,In_3384,In_2802);
xor U1712 (N_1712,In_3958,In_3803);
nor U1713 (N_1713,N_239,In_3329);
nand U1714 (N_1714,In_2877,In_1425);
nand U1715 (N_1715,N_365,In_1716);
xnor U1716 (N_1716,In_478,In_4993);
or U1717 (N_1717,N_1183,N_1065);
nand U1718 (N_1718,In_1097,N_320);
nor U1719 (N_1719,In_4951,In_4641);
nor U1720 (N_1720,N_1013,In_3802);
or U1721 (N_1721,In_988,In_2912);
nand U1722 (N_1722,In_4627,In_2260);
or U1723 (N_1723,In_3351,N_529);
or U1724 (N_1724,N_1320,In_3294);
and U1725 (N_1725,In_3897,N_1370);
nor U1726 (N_1726,In_896,In_3063);
nor U1727 (N_1727,In_236,N_166);
or U1728 (N_1728,In_4794,In_3271);
nor U1729 (N_1729,In_1663,In_1655);
or U1730 (N_1730,In_3794,In_2768);
nor U1731 (N_1731,In_761,In_690);
and U1732 (N_1732,In_2542,In_4406);
nor U1733 (N_1733,N_470,N_1445);
nor U1734 (N_1734,N_975,In_1087);
nor U1735 (N_1735,In_3476,N_169);
and U1736 (N_1736,N_1341,In_3621);
nor U1737 (N_1737,In_3133,N_1326);
nand U1738 (N_1738,In_664,In_247);
nor U1739 (N_1739,In_4525,N_1284);
or U1740 (N_1740,N_1444,N_1476);
and U1741 (N_1741,In_3163,In_3767);
nand U1742 (N_1742,In_1073,In_4052);
or U1743 (N_1743,In_1869,In_1494);
and U1744 (N_1744,In_4501,N_1366);
nand U1745 (N_1745,In_3321,In_3441);
nand U1746 (N_1746,N_906,In_4326);
and U1747 (N_1747,N_1425,In_4611);
nor U1748 (N_1748,N_667,In_798);
nor U1749 (N_1749,In_4094,In_1416);
nor U1750 (N_1750,In_976,In_4001);
and U1751 (N_1751,In_3930,In_1654);
nand U1752 (N_1752,In_206,In_2923);
nand U1753 (N_1753,N_524,N_337);
xnor U1754 (N_1754,In_4273,In_2731);
nor U1755 (N_1755,In_3991,In_586);
nor U1756 (N_1756,N_733,In_2901);
nand U1757 (N_1757,In_1905,N_203);
nand U1758 (N_1758,N_896,In_4485);
nor U1759 (N_1759,N_309,In_4704);
xor U1760 (N_1760,In_4928,N_229);
and U1761 (N_1761,In_1224,In_495);
xor U1762 (N_1762,N_528,In_4437);
nor U1763 (N_1763,In_1431,In_1563);
xnor U1764 (N_1764,In_1956,N_946);
nand U1765 (N_1765,N_1443,N_425);
and U1766 (N_1766,In_3558,In_1437);
nand U1767 (N_1767,N_1362,In_1851);
nand U1768 (N_1768,N_1113,N_938);
and U1769 (N_1769,In_3022,In_4712);
and U1770 (N_1770,In_3237,In_3420);
nand U1771 (N_1771,N_1230,In_1555);
xor U1772 (N_1772,N_1058,In_2743);
nor U1773 (N_1773,In_4063,In_4208);
or U1774 (N_1774,In_1980,N_1298);
nor U1775 (N_1775,N_506,N_168);
nand U1776 (N_1776,In_1888,N_302);
or U1777 (N_1777,In_1856,In_3016);
nor U1778 (N_1778,In_4578,In_3537);
xnor U1779 (N_1779,In_46,In_2050);
or U1780 (N_1780,In_2086,In_1959);
nand U1781 (N_1781,N_585,N_707);
nor U1782 (N_1782,N_361,N_1399);
and U1783 (N_1783,In_1732,In_4886);
nand U1784 (N_1784,In_4747,In_4199);
and U1785 (N_1785,In_3571,In_2485);
nand U1786 (N_1786,N_1308,In_2322);
or U1787 (N_1787,In_3758,N_893);
nor U1788 (N_1788,In_2298,In_2479);
and U1789 (N_1789,In_2975,In_3585);
nand U1790 (N_1790,N_976,N_1423);
nand U1791 (N_1791,In_3416,In_2812);
or U1792 (N_1792,In_1940,N_264);
nand U1793 (N_1793,In_702,In_4649);
nand U1794 (N_1794,N_193,In_678);
and U1795 (N_1795,In_841,N_613);
or U1796 (N_1796,In_2672,In_2508);
and U1797 (N_1797,N_1119,In_3402);
nand U1798 (N_1798,In_3448,N_1288);
nand U1799 (N_1799,In_4710,N_682);
xor U1800 (N_1800,In_1631,In_1046);
nor U1801 (N_1801,In_3994,In_3225);
xor U1802 (N_1802,N_463,In_4557);
nor U1803 (N_1803,In_4012,In_241);
or U1804 (N_1804,In_3933,In_739);
nor U1805 (N_1805,In_2448,In_2106);
xor U1806 (N_1806,In_4508,In_1882);
or U1807 (N_1807,In_4125,N_593);
nor U1808 (N_1808,In_4516,N_1161);
nor U1809 (N_1809,In_3033,In_580);
or U1810 (N_1810,In_2199,In_3403);
nand U1811 (N_1811,In_3446,N_571);
nand U1812 (N_1812,In_4952,In_3186);
nor U1813 (N_1813,In_1757,In_2793);
xnor U1814 (N_1814,N_1384,N_1272);
nor U1815 (N_1815,In_1399,In_2712);
nor U1816 (N_1816,In_506,N_1499);
nor U1817 (N_1817,N_1367,In_1510);
nand U1818 (N_1818,In_561,In_2137);
and U1819 (N_1819,N_1117,In_2357);
nand U1820 (N_1820,In_2410,In_3990);
nor U1821 (N_1821,In_2253,N_1241);
nand U1822 (N_1822,In_4124,N_951);
nand U1823 (N_1823,N_444,N_829);
nand U1824 (N_1824,In_2059,In_4152);
nand U1825 (N_1825,In_4178,In_1527);
xnor U1826 (N_1826,N_342,N_358);
nand U1827 (N_1827,In_577,In_4902);
or U1828 (N_1828,N_424,In_2819);
nor U1829 (N_1829,In_875,N_1277);
nand U1830 (N_1830,In_3804,N_776);
xnor U1831 (N_1831,N_101,N_494);
and U1832 (N_1832,N_723,In_2543);
nor U1833 (N_1833,In_2104,In_1322);
nor U1834 (N_1834,In_937,In_1249);
nor U1835 (N_1835,In_1364,In_538);
or U1836 (N_1836,N_1373,In_4725);
or U1837 (N_1837,In_3103,N_1453);
nor U1838 (N_1838,In_2342,In_2545);
nand U1839 (N_1839,N_1211,In_4657);
or U1840 (N_1840,In_3261,In_3091);
or U1841 (N_1841,N_451,In_4970);
nor U1842 (N_1842,N_962,In_548);
nor U1843 (N_1843,N_1316,In_1529);
and U1844 (N_1844,N_638,In_212);
and U1845 (N_1845,In_1569,In_3561);
nand U1846 (N_1846,N_512,N_1477);
and U1847 (N_1847,In_2478,In_3034);
and U1848 (N_1848,N_1138,In_1934);
and U1849 (N_1849,In_3014,N_336);
or U1850 (N_1850,In_3330,In_2969);
nand U1851 (N_1851,N_701,N_994);
xnor U1852 (N_1852,N_1433,In_1279);
or U1853 (N_1853,N_1254,In_195);
nor U1854 (N_1854,In_4810,In_1735);
nand U1855 (N_1855,In_1071,In_3661);
nand U1856 (N_1856,In_2995,In_972);
xor U1857 (N_1857,In_4004,N_647);
nand U1858 (N_1858,In_3549,In_4243);
nand U1859 (N_1859,In_961,N_1157);
or U1860 (N_1860,In_575,In_763);
nand U1861 (N_1861,In_1949,N_439);
or U1862 (N_1862,N_191,In_4787);
nand U1863 (N_1863,N_354,In_3154);
nor U1864 (N_1864,In_1300,In_3435);
xnor U1865 (N_1865,In_3005,In_1951);
nor U1866 (N_1866,In_3680,In_4363);
nor U1867 (N_1867,In_339,N_1360);
nor U1868 (N_1868,In_789,N_1469);
or U1869 (N_1869,In_4900,N_1387);
nor U1870 (N_1870,N_410,In_616);
or U1871 (N_1871,In_4618,N_610);
nand U1872 (N_1872,In_4677,In_1936);
or U1873 (N_1873,N_1470,In_3591);
nor U1874 (N_1874,In_1260,In_1619);
or U1875 (N_1875,In_1937,N_924);
or U1876 (N_1876,N_953,In_4879);
and U1877 (N_1877,In_1320,In_4171);
xor U1878 (N_1878,In_686,In_2696);
xor U1879 (N_1879,In_3469,In_530);
nor U1880 (N_1880,In_2951,In_750);
and U1881 (N_1881,N_935,N_668);
nand U1882 (N_1882,N_735,N_607);
or U1883 (N_1883,N_15,In_2698);
nand U1884 (N_1884,In_4079,N_230);
or U1885 (N_1885,In_547,N_413);
and U1886 (N_1886,In_1670,In_3822);
nor U1887 (N_1887,N_555,In_797);
nor U1888 (N_1888,N_901,In_3862);
and U1889 (N_1889,N_1325,In_324);
or U1890 (N_1890,In_4539,N_1276);
xor U1891 (N_1891,In_2735,N_1086);
nand U1892 (N_1892,In_4583,In_4233);
nand U1893 (N_1893,In_4944,In_2760);
and U1894 (N_1894,N_1005,In_1484);
nand U1895 (N_1895,In_2355,N_1106);
nand U1896 (N_1896,In_4083,In_20);
or U1897 (N_1897,In_1287,In_2580);
nor U1898 (N_1898,N_716,N_258);
nand U1899 (N_1899,In_4841,In_2562);
xnor U1900 (N_1900,In_744,N_536);
and U1901 (N_1901,N_1095,In_643);
nand U1902 (N_1902,In_4824,In_1028);
or U1903 (N_1903,In_4108,In_3612);
xor U1904 (N_1904,In_4466,N_1280);
nand U1905 (N_1905,N_643,In_1206);
and U1906 (N_1906,N_255,N_1307);
or U1907 (N_1907,In_3206,In_3982);
nand U1908 (N_1908,In_2695,In_622);
xnor U1909 (N_1909,N_1485,In_4354);
and U1910 (N_1910,In_749,In_524);
or U1911 (N_1911,N_781,In_4621);
nor U1912 (N_1912,In_1420,In_3646);
or U1913 (N_1913,N_1431,In_3643);
or U1914 (N_1914,In_4664,N_85);
and U1915 (N_1915,In_2054,In_2945);
xnor U1916 (N_1916,In_1506,N_1092);
and U1917 (N_1917,N_541,In_1468);
nand U1918 (N_1918,N_780,In_4862);
xnor U1919 (N_1919,In_2573,N_1025);
or U1920 (N_1920,In_1656,In_2608);
nor U1921 (N_1921,In_342,In_107);
nand U1922 (N_1922,N_1201,N_750);
nand U1923 (N_1923,In_3405,N_767);
or U1924 (N_1924,N_376,N_284);
nor U1925 (N_1925,In_4924,In_2414);
or U1926 (N_1926,N_102,In_37);
or U1927 (N_1927,In_4805,N_874);
xnor U1928 (N_1928,In_2374,In_106);
nand U1929 (N_1929,N_932,N_535);
nand U1930 (N_1930,In_1436,N_579);
and U1931 (N_1931,N_890,N_677);
and U1932 (N_1932,N_1198,In_2074);
and U1933 (N_1933,N_1406,N_969);
or U1934 (N_1934,In_769,N_1023);
or U1935 (N_1935,In_1180,N_266);
xnor U1936 (N_1936,In_1236,N_89);
or U1937 (N_1937,In_1443,In_60);
or U1938 (N_1938,In_1902,N_1177);
and U1939 (N_1939,In_3818,In_4531);
nand U1940 (N_1940,In_1196,In_2787);
nor U1941 (N_1941,In_232,N_925);
or U1942 (N_1942,In_1973,N_1409);
and U1943 (N_1943,N_1283,In_4219);
or U1944 (N_1944,N_1098,In_4137);
or U1945 (N_1945,In_3341,N_383);
nand U1946 (N_1946,In_3844,N_1279);
nor U1947 (N_1947,In_1707,N_1450);
and U1948 (N_1948,In_2815,In_3907);
nand U1949 (N_1949,In_472,In_1410);
and U1950 (N_1950,N_887,In_4371);
nor U1951 (N_1951,In_3784,In_4593);
xor U1952 (N_1952,In_3172,In_605);
and U1953 (N_1953,N_435,In_2021);
and U1954 (N_1954,In_3848,In_4146);
nand U1955 (N_1955,In_966,In_3843);
and U1956 (N_1956,N_1100,N_1006);
nor U1957 (N_1957,N_1234,N_371);
nand U1958 (N_1958,N_860,N_1394);
or U1959 (N_1959,In_1124,In_1717);
or U1960 (N_1960,In_827,N_109);
or U1961 (N_1961,In_1558,In_3546);
and U1962 (N_1962,In_209,In_4198);
xnor U1963 (N_1963,In_3514,In_48);
nor U1964 (N_1964,In_4394,In_3594);
and U1965 (N_1965,In_2179,In_2575);
and U1966 (N_1966,In_4077,In_1604);
nor U1967 (N_1967,In_698,In_536);
or U1968 (N_1968,N_1227,In_2464);
or U1969 (N_1969,In_71,N_551);
or U1970 (N_1970,In_4584,N_426);
nor U1971 (N_1971,In_1432,In_565);
nor U1972 (N_1972,In_397,In_1715);
and U1973 (N_1973,In_4401,N_557);
and U1974 (N_1974,In_4658,In_4025);
nor U1975 (N_1975,N_1231,In_4846);
and U1976 (N_1976,In_1390,N_1289);
nand U1977 (N_1977,N_1209,In_3788);
nand U1978 (N_1978,In_3720,In_1546);
and U1979 (N_1979,In_4138,In_925);
or U1980 (N_1980,In_1946,In_4933);
or U1981 (N_1981,In_4110,N_1);
nor U1982 (N_1982,In_196,In_4407);
nand U1983 (N_1983,In_4073,N_678);
and U1984 (N_1984,N_186,In_1181);
or U1985 (N_1985,In_2831,In_3460);
xor U1986 (N_1986,In_1914,N_729);
or U1987 (N_1987,In_979,In_4299);
or U1988 (N_1988,N_1412,In_2192);
nand U1989 (N_1989,In_2399,In_1600);
nor U1990 (N_1990,In_1824,N_338);
nand U1991 (N_1991,In_2582,In_4322);
nand U1992 (N_1992,In_510,N_487);
nor U1993 (N_1993,In_2703,N_1439);
nand U1994 (N_1994,In_3611,In_742);
nor U1995 (N_1995,N_1269,In_3006);
nand U1996 (N_1996,In_3573,In_3583);
and U1997 (N_1997,N_756,N_688);
or U1998 (N_1998,N_1488,N_310);
and U1999 (N_1999,In_3739,In_1151);
nor U2000 (N_2000,N_574,In_1215);
and U2001 (N_2001,N_1981,In_279);
or U2002 (N_2002,In_1075,In_4148);
or U2003 (N_2003,N_1487,In_96);
nand U2004 (N_2004,N_1958,N_1250);
nand U2005 (N_2005,N_850,In_3110);
or U2006 (N_2006,In_1219,N_1625);
or U2007 (N_2007,In_4478,N_54);
or U2008 (N_2008,In_3952,In_3087);
or U2009 (N_2009,N_1896,N_1882);
nor U2010 (N_2010,N_1849,N_151);
or U2011 (N_2011,In_3769,In_2769);
nand U2012 (N_2012,N_1038,In_2353);
nand U2013 (N_2013,N_1783,In_445);
and U2014 (N_2014,In_383,In_4543);
nor U2015 (N_2015,In_3051,In_2806);
or U2016 (N_2016,In_3733,N_1459);
and U2017 (N_2017,In_785,In_143);
and U2018 (N_2018,In_2913,In_3688);
xor U2019 (N_2019,In_3097,N_936);
nor U2020 (N_2020,N_1660,N_1557);
or U2021 (N_2021,N_1612,N_1737);
or U2022 (N_2022,In_4227,In_913);
or U2023 (N_2023,In_3761,N_879);
and U2024 (N_2024,N_1801,In_3221);
or U2025 (N_2025,In_4529,N_420);
or U2026 (N_2026,N_844,In_2078);
nor U2027 (N_2027,In_4871,N_1246);
nand U2028 (N_2028,In_288,N_137);
and U2029 (N_2029,In_3533,N_1441);
nor U2030 (N_2030,In_1693,In_2620);
or U2031 (N_2031,N_1950,In_1651);
or U2032 (N_2032,N_1057,In_2839);
nor U2033 (N_2033,N_1750,In_1067);
and U2034 (N_2034,N_57,N_841);
nand U2035 (N_2035,In_2561,In_2343);
or U2036 (N_2036,In_4882,In_2146);
and U2037 (N_2037,N_1893,In_3270);
and U2038 (N_2038,In_1884,N_1505);
xnor U2039 (N_2039,N_1353,N_1711);
nor U2040 (N_2040,N_1964,N_1514);
or U2041 (N_2041,In_2327,In_124);
nor U2042 (N_2042,In_3057,N_1171);
or U2043 (N_2043,In_535,N_1747);
or U2044 (N_2044,N_1233,In_1662);
nand U2045 (N_2045,N_171,In_1343);
nand U2046 (N_2046,In_872,In_1027);
nor U2047 (N_2047,In_2963,In_1761);
or U2048 (N_2048,In_2701,In_2177);
nand U2049 (N_2049,N_1634,N_817);
nand U2050 (N_2050,In_2906,N_873);
and U2051 (N_2051,N_1224,N_185);
nor U2052 (N_2052,In_3165,In_4444);
nand U2053 (N_2053,N_437,In_4274);
xnor U2054 (N_2054,N_1344,N_1359);
and U2055 (N_2055,N_1738,N_373);
or U2056 (N_2056,In_3127,N_1813);
nor U2057 (N_2057,In_2875,N_641);
xnor U2058 (N_2058,N_1836,N_958);
or U2059 (N_2059,N_36,In_3855);
xor U2060 (N_2060,In_1724,In_3665);
nand U2061 (N_2061,In_3510,N_1497);
or U2062 (N_2062,In_3278,In_658);
and U2063 (N_2063,In_4920,N_1486);
nor U2064 (N_2064,N_1114,N_891);
and U2065 (N_2065,N_405,N_366);
nand U2066 (N_2066,In_970,In_613);
and U2067 (N_2067,In_3121,N_1946);
nor U2068 (N_2068,N_1826,N_24);
xor U2069 (N_2069,N_931,N_1935);
and U2070 (N_2070,In_1335,In_1645);
xor U2071 (N_2071,In_2693,In_1686);
or U2072 (N_2072,In_4690,N_272);
or U2073 (N_2073,In_852,N_617);
nor U2074 (N_2074,In_2071,In_68);
nor U2075 (N_2075,In_3617,N_448);
and U2076 (N_2076,N_1034,N_1489);
or U2077 (N_2077,In_878,In_2366);
or U2078 (N_2078,N_1297,N_1725);
nor U2079 (N_2079,In_1977,In_4366);
and U2080 (N_2080,N_1202,In_1286);
nor U2081 (N_2081,N_1675,N_501);
nand U2082 (N_2082,N_66,N_1601);
nand U2083 (N_2083,In_3359,In_2075);
nand U2084 (N_2084,In_817,N_1069);
nand U2085 (N_2085,N_955,N_1892);
or U2086 (N_2086,In_4758,In_2546);
or U2087 (N_2087,N_1570,In_1836);
nand U2088 (N_2088,N_1723,N_486);
nand U2089 (N_2089,N_1393,In_2134);
or U2090 (N_2090,N_1943,In_3032);
and U2091 (N_2091,In_1570,In_1185);
xor U2092 (N_2092,In_821,N_823);
or U2093 (N_2093,N_1524,N_1448);
and U2094 (N_2094,In_2108,N_1204);
or U2095 (N_2095,In_1137,In_2623);
and U2096 (N_2096,In_498,In_3479);
and U2097 (N_2097,N_1758,N_1434);
nor U2098 (N_2098,N_1350,N_1475);
or U2099 (N_2099,N_1756,In_1217);
nand U2100 (N_2100,In_3615,N_1884);
nor U2101 (N_2101,In_4918,N_1383);
nand U2102 (N_2102,N_1595,In_965);
nand U2103 (N_2103,N_1240,N_997);
and U2104 (N_2104,N_1551,In_512);
nand U2105 (N_2105,In_3715,In_277);
nor U2106 (N_2106,N_1024,N_1546);
xnor U2107 (N_2107,In_2161,In_4413);
nor U2108 (N_2108,In_2897,N_74);
and U2109 (N_2109,In_2060,In_2683);
nand U2110 (N_2110,In_268,N_1510);
and U2111 (N_2111,In_1447,N_1797);
nand U2112 (N_2112,N_1096,N_1651);
and U2113 (N_2113,In_3350,In_4030);
nor U2114 (N_2114,In_4996,In_4147);
nor U2115 (N_2115,N_837,In_3773);
nand U2116 (N_2116,N_645,N_1237);
or U2117 (N_2117,In_2037,In_829);
and U2118 (N_2118,In_1605,N_1457);
nand U2119 (N_2119,In_1077,In_2257);
nor U2120 (N_2120,N_1938,N_1670);
nor U2121 (N_2121,In_2967,In_1421);
or U2122 (N_2122,N_1094,In_3060);
or U2123 (N_2123,N_1127,In_4467);
nor U2124 (N_2124,N_812,N_1729);
nand U2125 (N_2125,N_1312,In_4514);
nand U2126 (N_2126,In_3911,N_1293);
nor U2127 (N_2127,N_1754,In_4670);
or U2128 (N_2128,In_1986,In_3182);
xor U2129 (N_2129,N_1292,N_1784);
nand U2130 (N_2130,In_3113,In_4804);
or U2131 (N_2131,In_2903,In_869);
nor U2132 (N_2132,N_96,In_2026);
and U2133 (N_2133,N_1692,In_3791);
and U2134 (N_2134,N_1822,N_1733);
or U2135 (N_2135,In_573,N_1073);
nor U2136 (N_2136,In_1478,N_1043);
nand U2137 (N_2137,In_4418,In_2451);
nor U2138 (N_2138,In_4402,N_428);
or U2139 (N_2139,In_2056,In_3593);
and U2140 (N_2140,In_721,N_1984);
or U2141 (N_2141,In_1681,In_1081);
and U2142 (N_2142,In_924,N_440);
or U2143 (N_2143,In_2460,In_3390);
nand U2144 (N_2144,In_4561,N_655);
xnor U2145 (N_2145,In_485,N_1914);
and U2146 (N_2146,In_4134,N_1974);
and U2147 (N_2147,In_1971,In_1295);
xor U2148 (N_2148,In_1107,N_1763);
nand U2149 (N_2149,In_3289,N_414);
nand U2150 (N_2150,In_394,In_1148);
or U2151 (N_2151,In_3506,N_1888);
or U2152 (N_2152,In_155,N_1081);
and U2153 (N_2153,In_4660,In_2595);
nor U2154 (N_2154,In_3556,In_3158);
xor U2155 (N_2155,In_187,In_4987);
nor U2156 (N_2156,In_2873,In_1166);
and U2157 (N_2157,In_1011,In_2609);
and U2158 (N_2158,In_244,In_3304);
or U2159 (N_2159,In_488,In_314);
and U2160 (N_2160,N_1258,N_1159);
nor U2161 (N_2161,N_1877,N_1697);
nand U2162 (N_2162,N_408,N_1340);
nor U2163 (N_2163,N_1195,In_1786);
or U2164 (N_2164,In_4457,N_1713);
nand U2165 (N_2165,N_1111,N_1552);
nor U2166 (N_2166,In_4775,In_1953);
and U2167 (N_2167,In_1874,N_737);
nand U2168 (N_2168,N_23,N_130);
and U2169 (N_2169,In_4504,N_369);
nor U2170 (N_2170,N_1987,In_3228);
nand U2171 (N_2171,N_1704,In_4258);
nor U2172 (N_2172,In_2981,N_1508);
and U2173 (N_2173,In_2175,In_1700);
nand U2174 (N_2174,In_266,In_3723);
or U2175 (N_2175,In_15,N_1369);
nand U2176 (N_2176,N_858,In_4279);
nor U2177 (N_2177,In_2763,In_4074);
or U2178 (N_2178,In_3955,N_296);
nand U2179 (N_2179,In_4218,N_1389);
nor U2180 (N_2180,N_569,N_967);
nand U2181 (N_2181,In_809,N_601);
xor U2182 (N_2182,In_1659,N_389);
or U2183 (N_2183,In_3382,In_4930);
or U2184 (N_2184,In_2780,N_86);
nor U2185 (N_2185,In_2745,In_296);
nor U2186 (N_2186,N_1175,In_1266);
and U2187 (N_2187,N_611,N_849);
and U2188 (N_2188,In_3126,In_4984);
xor U2189 (N_2189,In_1463,N_1975);
nand U2190 (N_2190,In_1852,In_4458);
nand U2191 (N_2191,In_1548,In_3422);
nor U2192 (N_2192,N_1135,In_2653);
nor U2193 (N_2193,In_1281,In_4835);
nand U2194 (N_2194,N_1238,In_4236);
nand U2195 (N_2195,N_1579,In_4542);
or U2196 (N_2196,In_1741,In_4303);
and U2197 (N_2197,N_1846,In_4782);
or U2198 (N_2198,N_1108,N_734);
nor U2199 (N_2199,N_488,In_4421);
nor U2200 (N_2200,In_2367,N_1068);
nor U2201 (N_2201,In_3036,N_1908);
or U2202 (N_2202,In_807,N_1709);
nand U2203 (N_2203,N_392,N_1363);
or U2204 (N_2204,In_3627,In_4207);
nand U2205 (N_2205,In_404,In_353);
nand U2206 (N_2206,In_260,N_1594);
and U2207 (N_2207,N_65,N_1788);
nor U2208 (N_2208,In_1052,N_1796);
and U2209 (N_2209,In_4915,In_2133);
or U2210 (N_2210,In_4201,N_987);
nand U2211 (N_2211,N_1155,N_1627);
xor U2212 (N_2212,N_1158,In_2585);
or U2213 (N_2213,In_4753,N_252);
nor U2214 (N_2214,In_1522,N_875);
nand U2215 (N_2215,N_1746,N_1591);
nand U2216 (N_2216,In_662,In_4963);
nor U2217 (N_2217,In_2700,N_1921);
and U2218 (N_2218,N_1203,In_1499);
nor U2219 (N_2219,N_1219,N_1834);
nor U2220 (N_2220,N_595,In_1189);
or U2221 (N_2221,N_968,N_132);
nor U2222 (N_2222,N_313,In_2306);
nor U2223 (N_2223,In_3685,N_695);
or U2224 (N_2224,In_3152,N_1932);
and U2225 (N_2225,N_67,In_1726);
nand U2226 (N_2226,N_1656,In_1826);
nand U2227 (N_2227,In_3099,N_156);
nor U2228 (N_2228,N_1926,N_1855);
xnor U2229 (N_2229,In_4519,N_1575);
xor U2230 (N_2230,N_1550,In_4497);
nor U2231 (N_2231,N_1973,In_1446);
nor U2232 (N_2232,In_4637,In_1898);
or U2233 (N_2233,In_2930,In_4041);
or U2234 (N_2234,In_1099,N_843);
nor U2235 (N_2235,In_1964,In_1928);
nor U2236 (N_2236,N_1042,In_18);
nor U2237 (N_2237,N_1952,In_3879);
nor U2238 (N_2238,In_4832,In_973);
nor U2239 (N_2239,N_1694,In_35);
nor U2240 (N_2240,In_4942,In_3559);
nand U2241 (N_2241,In_1285,In_1000);
and U2242 (N_2242,N_600,In_1183);
and U2243 (N_2243,In_411,N_1534);
or U2244 (N_2244,In_4829,N_219);
nand U2245 (N_2245,In_4314,In_971);
and U2246 (N_2246,N_1646,In_4746);
and U2247 (N_2247,In_3825,In_382);
or U2248 (N_2248,In_101,In_587);
and U2249 (N_2249,In_3957,In_1912);
nand U2250 (N_2250,N_1221,N_1971);
and U2251 (N_2251,In_3608,In_4130);
nor U2252 (N_2252,In_673,In_3544);
or U2253 (N_2253,In_4786,N_526);
or U2254 (N_2254,N_1821,N_1574);
and U2255 (N_2255,N_1194,In_4909);
and U2256 (N_2256,N_696,In_2705);
nand U2257 (N_2257,In_2474,In_224);
nand U2258 (N_2258,N_19,N_273);
and U2259 (N_2259,In_1702,N_1236);
or U2260 (N_2260,In_51,In_1383);
or U2261 (N_2261,In_3921,In_3140);
and U2262 (N_2262,In_1862,N_73);
nand U2263 (N_2263,In_3002,In_2503);
nand U2264 (N_2264,N_1120,N_1056);
and U2265 (N_2265,N_1395,N_1011);
nand U2266 (N_2266,In_1312,In_4080);
nand U2267 (N_2267,N_1408,In_2895);
xnor U2268 (N_2268,N_1131,In_3983);
nor U2269 (N_2269,In_591,In_948);
nand U2270 (N_2270,In_731,In_3338);
nor U2271 (N_2271,In_3310,In_4453);
nor U2272 (N_2272,In_1549,In_2393);
or U2273 (N_2273,In_1352,N_100);
xnor U2274 (N_2274,N_1416,N_1863);
nor U2275 (N_2275,N_433,N_353);
or U2276 (N_2276,In_4500,N_90);
nor U2277 (N_2277,In_3501,N_900);
nor U2278 (N_2278,In_4017,In_3881);
nand U2279 (N_2279,N_1872,In_1866);
xor U2280 (N_2280,N_1352,N_293);
xor U2281 (N_2281,In_492,In_4024);
xor U2282 (N_2282,In_3279,In_2599);
nor U2283 (N_2283,In_921,In_4179);
nor U2284 (N_2284,In_3213,In_2809);
nor U2285 (N_2285,N_1876,N_1206);
nor U2286 (N_2286,N_1040,N_1886);
or U2287 (N_2287,N_1789,N_540);
nor U2288 (N_2288,N_40,N_681);
and U2289 (N_2289,N_1585,N_1956);
nand U2290 (N_2290,In_2035,In_685);
xor U2291 (N_2291,N_663,In_4954);
or U2292 (N_2292,In_4802,N_1410);
nand U2293 (N_2293,N_559,N_1641);
and U2294 (N_2294,In_1051,N_1396);
and U2295 (N_2295,In_3406,In_4319);
nand U2296 (N_2296,In_1451,N_1182);
nor U2297 (N_2297,N_1957,In_2352);
nor U2298 (N_2298,N_774,In_4221);
nor U2299 (N_2299,N_1351,In_4998);
or U2300 (N_2300,In_4471,In_1477);
or U2301 (N_2301,N_1681,In_3440);
nor U2302 (N_2302,N_214,N_1222);
nor U2303 (N_2303,In_378,N_1507);
and U2304 (N_2304,N_1839,N_1382);
nor U2305 (N_2305,In_2248,In_4380);
and U2306 (N_2306,In_3210,In_1218);
nand U2307 (N_2307,N_1511,N_1319);
nor U2308 (N_2308,N_1603,N_1604);
nand U2309 (N_2309,In_2049,N_1519);
or U2310 (N_2310,In_3331,In_884);
nor U2311 (N_2311,In_2317,N_722);
nor U2312 (N_2312,In_4376,N_1193);
and U2313 (N_2313,In_2647,In_745);
or U2314 (N_2314,N_525,In_4600);
and U2315 (N_2315,N_1731,In_4877);
or U2316 (N_2316,In_29,N_1152);
nor U2317 (N_2317,In_2528,N_1531);
xnor U2318 (N_2318,In_289,In_4880);
or U2319 (N_2319,N_1895,N_604);
nand U2320 (N_2320,In_1870,N_1945);
xor U2321 (N_2321,In_513,N_1532);
nand U2322 (N_2322,N_1808,In_1162);
nand U2323 (N_2323,In_3130,In_3413);
nand U2324 (N_2324,In_1843,In_2420);
nand U2325 (N_2325,N_656,N_1792);
nand U2326 (N_2326,N_253,In_2713);
nand U2327 (N_2327,In_2531,In_219);
or U2328 (N_2328,In_3889,N_1210);
xor U2329 (N_2329,N_1838,In_367);
nor U2330 (N_2330,In_2818,In_3018);
or U2331 (N_2331,N_580,In_2422);
or U2332 (N_2332,N_1047,In_3302);
and U2333 (N_2333,In_2719,In_417);
nor U2334 (N_2334,N_1684,In_4263);
xnor U2335 (N_2335,N_1866,N_1176);
or U2336 (N_2336,In_859,In_1452);
or U2337 (N_2337,N_1611,In_571);
and U2338 (N_2338,In_174,In_3637);
nor U2339 (N_2339,In_1589,N_920);
or U2340 (N_2340,N_871,N_1414);
and U2341 (N_2341,In_1756,In_2477);
nor U2342 (N_2342,In_3732,N_1590);
and U2343 (N_2343,In_3092,N_1481);
or U2344 (N_2344,In_3515,In_4864);
or U2345 (N_2345,In_2942,N_1154);
or U2346 (N_2346,In_4038,N_1167);
or U2347 (N_2347,N_1148,In_1875);
and U2348 (N_2348,In_2511,In_3629);
and U2349 (N_2349,In_3378,N_21);
nand U2350 (N_2350,In_2251,N_1463);
or U2351 (N_2351,N_378,N_662);
and U2352 (N_2352,In_1566,In_848);
and U2353 (N_2353,In_3023,N_1516);
nand U2354 (N_2354,In_692,In_2884);
nor U2355 (N_2355,N_261,N_1252);
nor U2356 (N_2356,In_4272,N_1392);
and U2357 (N_2357,In_4232,N_1816);
or U2358 (N_2358,In_2606,In_4891);
nand U2359 (N_2359,In_3258,N_516);
or U2360 (N_2360,In_1163,In_2671);
nand U2361 (N_2361,N_1715,N_1906);
and U2362 (N_2362,In_108,N_1712);
xor U2363 (N_2363,N_1588,N_1417);
or U2364 (N_2364,In_3745,In_4779);
xnor U2365 (N_2365,In_4450,In_1104);
and U2366 (N_2366,N_93,N_1407);
nand U2367 (N_2367,In_635,N_1530);
or U2368 (N_2368,In_4423,N_1480);
and U2369 (N_2369,In_4643,In_361);
nand U2370 (N_2370,N_142,N_1730);
and U2371 (N_2371,In_3965,In_4982);
and U2372 (N_2372,In_2061,N_816);
nand U2373 (N_2373,In_2515,In_851);
nor U2374 (N_2374,In_3015,In_4465);
nor U2375 (N_2375,In_1009,In_923);
and U2376 (N_2376,N_738,N_511);
nor U2377 (N_2377,In_4121,N_467);
nor U2378 (N_2378,N_78,In_4738);
and U2379 (N_2379,In_3452,N_1889);
or U2380 (N_2380,In_3436,In_482);
or U2381 (N_2381,In_3243,N_1883);
nand U2382 (N_2382,In_1583,In_838);
and U2383 (N_2383,N_1850,In_912);
or U2384 (N_2384,In_2292,In_778);
nor U2385 (N_2385,N_242,N_779);
nand U2386 (N_2386,In_3890,In_4214);
nand U2387 (N_2387,N_1275,N_1347);
nor U2388 (N_2388,N_187,N_1667);
and U2389 (N_2389,In_2232,In_4390);
and U2390 (N_2390,N_1266,In_1126);
and U2391 (N_2391,N_1494,In_3486);
nor U2392 (N_2392,In_416,In_474);
nand U2393 (N_2393,N_1770,In_4383);
nor U2394 (N_2394,In_2785,In_3620);
nor U2395 (N_2395,N_1164,N_1857);
nor U2396 (N_2396,In_1669,N_1637);
and U2397 (N_2397,N_1286,N_1020);
nand U2398 (N_2398,N_814,In_2423);
and U2399 (N_2399,N_1336,N_393);
nand U2400 (N_2400,N_813,In_2917);
xnor U2401 (N_2401,In_1608,In_3961);
nor U2402 (N_2402,N_746,In_4997);
or U2403 (N_2403,N_703,N_1951);
and U2404 (N_2404,In_1147,In_185);
or U2405 (N_2405,In_1774,N_883);
and U2406 (N_2406,In_4020,In_1541);
or U2407 (N_2407,In_2222,In_4934);
nor U2408 (N_2408,N_1529,In_1021);
and U2409 (N_2409,N_1767,In_4626);
and U2410 (N_2410,N_741,In_624);
nand U2411 (N_2411,N_1676,N_692);
xnor U2412 (N_2412,N_1815,N_970);
or U2413 (N_2413,In_758,N_148);
and U2414 (N_2414,N_1705,N_1125);
nor U2415 (N_2415,In_909,N_1891);
nand U2416 (N_2416,N_981,N_1602);
and U2417 (N_2417,N_1584,N_1188);
and U2418 (N_2418,In_3633,N_1418);
xnor U2419 (N_2419,In_4763,In_3457);
nor U2420 (N_2420,In_184,In_1091);
and U2421 (N_2421,In_4825,N_304);
nand U2422 (N_2422,In_1239,In_3948);
nand U2423 (N_2423,N_821,In_2279);
or U2424 (N_2424,In_997,In_1918);
xnor U2425 (N_2425,N_1215,In_983);
nand U2426 (N_2426,N_1693,In_3796);
nand U2427 (N_2427,In_2225,In_683);
nor U2428 (N_2428,In_1602,N_1536);
or U2429 (N_2429,In_1108,N_818);
nand U2430 (N_2430,N_1940,N_1379);
nor U2431 (N_2431,N_1055,N_1504);
nand U2432 (N_2432,In_1400,In_2640);
nor U2433 (N_2433,N_1028,N_1012);
or U2434 (N_2434,In_4733,N_1991);
and U2435 (N_2435,In_4301,N_1650);
nor U2436 (N_2436,N_1698,N_1960);
nand U2437 (N_2437,In_2848,N_1004);
and U2438 (N_2438,N_248,In_2842);
nor U2439 (N_2439,In_3307,In_4425);
and U2440 (N_2440,In_3019,In_2297);
nand U2441 (N_2441,N_795,N_1314);
or U2442 (N_2442,N_1721,In_2103);
and U2443 (N_2443,N_971,In_3318);
nor U2444 (N_2444,N_720,In_4260);
nand U2445 (N_2445,In_4875,N_158);
nor U2446 (N_2446,N_1755,In_4612);
or U2447 (N_2447,N_1572,N_1169);
xnor U2448 (N_2448,N_1539,In_2223);
or U2449 (N_2449,N_233,N_498);
xnor U2450 (N_2450,In_1568,In_716);
and U2451 (N_2451,In_163,N_1832);
nor U2452 (N_2452,In_3800,In_3142);
and U2453 (N_2453,In_4284,N_1232);
and U2454 (N_2454,In_2197,N_1420);
and U2455 (N_2455,In_1616,N_1749);
or U2456 (N_2456,N_1490,In_386);
or U2457 (N_2457,N_905,N_803);
nor U2458 (N_2458,N_519,N_1088);
and U2459 (N_2459,In_2472,N_683);
xnor U2460 (N_2460,In_1721,In_2032);
nand U2461 (N_2461,In_3179,In_329);
and U2462 (N_2462,N_326,In_3170);
or U2463 (N_2463,In_3135,N_1151);
nand U2464 (N_2464,In_1966,In_1880);
nor U2465 (N_2465,In_2114,In_1599);
nor U2466 (N_2466,In_66,N_1223);
nor U2467 (N_2467,In_579,In_2441);
nor U2468 (N_2468,In_3895,N_1898);
nor U2469 (N_2469,N_627,N_1007);
nor U2470 (N_2470,In_3974,In_3801);
and U2471 (N_2471,N_1993,In_2428);
nor U2472 (N_2472,N_1482,In_4370);
or U2473 (N_2473,In_4493,N_558);
and U2474 (N_2474,In_4697,In_3609);
nand U2475 (N_2475,In_3202,N_1636);
or U2476 (N_2476,N_1829,In_822);
or U2477 (N_2477,N_254,In_4088);
nor U2478 (N_2478,N_934,In_2341);
nand U2479 (N_2479,In_2855,In_2006);
nand U2480 (N_2480,In_4854,N_1190);
nor U2481 (N_2481,In_1516,N_1115);
and U2482 (N_2482,In_4744,In_2085);
nor U2483 (N_2483,N_362,In_1627);
nand U2484 (N_2484,In_217,In_3704);
nand U2485 (N_2485,N_1847,In_1906);
nand U2486 (N_2486,N_1290,In_590);
nand U2487 (N_2487,In_414,In_4749);
and U2488 (N_2488,In_3171,In_516);
nor U2489 (N_2489,N_859,In_4581);
nor U2490 (N_2490,In_4800,In_2940);
and U2491 (N_2491,In_4856,In_843);
xnor U2492 (N_2492,N_61,In_4831);
nor U2493 (N_2493,In_3395,N_1680);
nor U2494 (N_2494,In_2840,In_4789);
or U2495 (N_2495,In_1342,In_4617);
and U2496 (N_2496,In_1241,In_1);
nor U2497 (N_2497,In_4300,In_3604);
nor U2498 (N_2498,N_1809,In_2328);
or U2499 (N_2499,N_1947,In_2378);
xor U2500 (N_2500,N_2091,N_1720);
nor U2501 (N_2501,In_4919,In_1365);
and U2502 (N_2502,In_865,N_977);
or U2503 (N_2503,In_2191,N_2261);
nand U2504 (N_2504,In_3129,N_785);
xor U2505 (N_2505,N_1969,In_2554);
or U2506 (N_2506,In_1155,In_631);
nand U2507 (N_2507,In_2361,In_1396);
or U2508 (N_2508,In_1340,N_2215);
nor U2509 (N_2509,N_1027,N_1128);
and U2510 (N_2510,N_2180,N_2331);
nand U2511 (N_2511,N_1003,N_1775);
and U2512 (N_2512,N_1166,N_341);
nand U2513 (N_2513,N_2127,N_930);
and U2514 (N_2514,In_4277,In_2244);
or U2515 (N_2515,In_157,In_4667);
or U2516 (N_2516,N_2463,In_3467);
nand U2517 (N_2517,In_2405,In_2741);
nor U2518 (N_2518,N_2318,In_4843);
nor U2519 (N_2519,N_2207,In_2928);
nand U2520 (N_2520,In_659,N_1424);
or U2521 (N_2521,N_539,N_246);
nor U2522 (N_2522,N_188,In_4327);
and U2523 (N_2523,N_620,N_294);
and U2524 (N_2524,In_1883,In_3502);
or U2525 (N_2525,N_2290,In_2989);
nor U2526 (N_2526,In_1737,In_3041);
nor U2527 (N_2527,In_3083,In_2029);
nand U2528 (N_2528,N_2395,N_671);
or U2529 (N_2529,In_2622,N_350);
and U2530 (N_2530,N_276,N_1565);
or U2531 (N_2531,In_1169,N_1690);
or U2532 (N_2532,N_2041,In_1454);
and U2533 (N_2533,N_1626,N_1294);
nor U2534 (N_2534,In_4813,N_2134);
xnor U2535 (N_2535,N_1710,N_2048);
nor U2536 (N_2536,In_3260,N_2419);
nand U2537 (N_2537,N_1535,In_3475);
or U2538 (N_2538,In_2761,In_4442);
or U2539 (N_2539,N_2292,In_4706);
nand U2540 (N_2540,N_1582,N_1869);
or U2541 (N_2541,N_2240,In_3904);
nand U2542 (N_2542,N_2073,N_1054);
or U2543 (N_2543,In_3898,N_1515);
or U2544 (N_2544,In_1376,In_2160);
nand U2545 (N_2545,In_433,N_2248);
nand U2546 (N_2546,In_4663,N_2279);
nand U2547 (N_2547,In_1145,N_1483);
or U2548 (N_2548,N_1740,N_828);
nand U2549 (N_2549,In_1813,In_998);
or U2550 (N_2550,In_4665,N_98);
nand U2551 (N_2551,In_1841,N_2295);
or U2552 (N_2552,N_1909,N_1419);
and U2553 (N_2553,In_171,In_906);
nand U2554 (N_2554,In_2829,N_1657);
nand U2555 (N_2555,N_1200,N_1178);
nand U2556 (N_2556,N_2359,In_86);
or U2557 (N_2557,In_1417,In_3347);
or U2558 (N_2558,In_1624,In_1834);
and U2559 (N_2559,N_1703,N_1599);
or U2560 (N_2560,N_2308,In_3007);
nand U2561 (N_2561,In_1348,N_1343);
and U2562 (N_2562,In_4610,N_2204);
and U2563 (N_2563,In_1190,N_1456);
and U2564 (N_2564,N_1976,In_3509);
xor U2565 (N_2565,In_713,N_1070);
nand U2566 (N_2566,N_1773,N_1076);
xnor U2567 (N_2567,N_1002,In_3445);
or U2568 (N_2568,N_2214,N_1695);
nand U2569 (N_2569,In_3552,N_2407);
and U2570 (N_2570,In_2185,N_2130);
nand U2571 (N_2571,In_2084,In_2309);
and U2572 (N_2572,N_247,In_2721);
and U2573 (N_2573,In_4545,N_2222);
and U2574 (N_2574,In_3192,In_420);
nor U2575 (N_2575,In_2556,N_1318);
and U2576 (N_2576,In_3888,N_1804);
nor U2577 (N_2577,N_2296,N_917);
xor U2578 (N_2578,In_1525,N_861);
or U2579 (N_2579,In_49,In_4959);
and U2580 (N_2580,N_2254,N_2351);
nand U2581 (N_2581,N_2312,In_2291);
and U2582 (N_2582,N_2156,In_596);
or U2583 (N_2583,In_2380,N_768);
or U2584 (N_2584,N_1955,In_4296);
nand U2585 (N_2585,N_2045,N_2281);
or U2586 (N_2586,In_62,N_2287);
nor U2587 (N_2587,In_1810,In_1857);
nand U2588 (N_2588,In_4086,N_2498);
nor U2589 (N_2589,In_2935,N_1328);
and U2590 (N_2590,N_1109,N_2455);
nand U2591 (N_2591,N_2316,N_1085);
xnor U2592 (N_2592,N_1606,N_1257);
or U2593 (N_2593,N_1010,N_1873);
nand U2594 (N_2594,N_1376,In_1284);
nor U2595 (N_2595,N_55,In_388);
or U2596 (N_2596,In_1030,N_1716);
and U2597 (N_2597,In_866,N_523);
and U2598 (N_2598,N_1248,N_870);
or U2599 (N_2599,In_4215,In_3197);
nand U2600 (N_2600,N_2424,N_989);
nor U2601 (N_2601,In_220,N_732);
and U2602 (N_2602,N_218,N_947);
nor U2603 (N_2603,In_2268,In_1235);
nor U2604 (N_2604,N_809,N_194);
and U2605 (N_2605,N_113,N_1661);
nor U2606 (N_2606,In_2710,N_1580);
nor U2607 (N_2607,In_1256,In_2125);
nand U2608 (N_2608,N_2243,In_3610);
and U2609 (N_2609,In_4490,In_2800);
and U2610 (N_2610,In_1354,N_2411);
nor U2611 (N_2611,In_3181,In_316);
nor U2612 (N_2612,N_1771,N_2483);
nand U2613 (N_2613,N_1683,In_3357);
or U2614 (N_2614,In_2219,In_614);
nand U2615 (N_2615,In_4979,N_2428);
nand U2616 (N_2616,N_986,In_180);
nor U2617 (N_2617,In_2999,In_2863);
nor U2618 (N_2618,In_261,N_760);
nor U2619 (N_2619,N_824,N_1912);
and U2620 (N_2620,N_2006,N_804);
and U2621 (N_2621,In_4634,N_1781);
or U2622 (N_2622,N_985,N_1858);
nand U2623 (N_2623,In_1865,N_1968);
nand U2624 (N_2624,In_1393,N_1736);
xor U2625 (N_2625,N_1920,In_1626);
nand U2626 (N_2626,N_1701,N_625);
and U2627 (N_2627,In_1246,N_1179);
nand U2628 (N_2628,N_447,N_2039);
or U2629 (N_2629,In_933,N_2220);
nor U2630 (N_2630,In_1078,In_3935);
xor U2631 (N_2631,N_1622,N_2036);
nor U2632 (N_2632,N_1549,N_983);
nand U2633 (N_2633,N_1875,N_2349);
or U2634 (N_2634,N_280,In_459);
nor U2635 (N_2635,N_991,N_2229);
nor U2636 (N_2636,N_2037,In_90);
or U2637 (N_2637,N_257,N_111);
xor U2638 (N_2638,N_2178,N_2051);
xor U2639 (N_2639,In_2376,In_4757);
or U2640 (N_2640,In_3472,In_3601);
and U2641 (N_2641,N_1904,N_902);
xor U2642 (N_2642,N_1066,In_920);
nor U2643 (N_2643,In_2990,In_2148);
nor U2644 (N_2644,N_2472,N_854);
or U2645 (N_2645,N_2101,In_1109);
nor U2646 (N_2646,In_2979,N_1890);
nand U2647 (N_2647,N_221,In_1426);
and U2648 (N_2648,N_1970,In_40);
and U2649 (N_2649,N_1666,N_1853);
nor U2650 (N_2650,In_4983,N_865);
or U2651 (N_2651,In_1943,In_4408);
nand U2652 (N_2652,N_1944,In_1921);
xor U2653 (N_2653,N_2343,N_1305);
nand U2654 (N_2654,In_169,In_21);
nand U2655 (N_2655,N_2228,In_2196);
nor U2656 (N_2656,N_599,N_2244);
nor U2657 (N_2657,In_2284,In_4737);
and U2658 (N_2658,In_1903,In_4674);
nand U2659 (N_2659,In_648,In_1970);
nand U2660 (N_2660,In_1088,N_995);
or U2661 (N_2661,In_4567,N_1630);
nand U2662 (N_2662,N_898,In_2521);
nor U2663 (N_2663,N_1075,N_2413);
or U2664 (N_2664,In_4325,N_2192);
nor U2665 (N_2665,N_2137,N_2093);
and U2666 (N_2666,N_744,N_2205);
or U2667 (N_2667,In_4926,N_2384);
or U2668 (N_2668,In_2120,In_4290);
and U2669 (N_2669,In_1489,N_497);
nor U2670 (N_2670,N_2421,In_3283);
nor U2671 (N_2671,N_1150,N_1346);
xor U2672 (N_2672,In_2798,N_1766);
and U2673 (N_2673,N_2181,N_2015);
xor U2674 (N_2674,In_3265,In_1553);
and U2675 (N_2675,N_1617,N_2010);
nor U2676 (N_2676,In_1598,N_1300);
nand U2677 (N_2677,N_1571,N_1102);
nand U2678 (N_2678,N_1146,In_4288);
xor U2679 (N_2679,In_652,In_4364);
nand U2680 (N_2680,N_757,N_1256);
nand U2681 (N_2681,In_276,N_2206);
nand U2682 (N_2682,In_1240,In_3763);
xor U2683 (N_2683,In_1900,In_2016);
or U2684 (N_2684,In_2285,N_1438);
and U2685 (N_2685,N_2477,N_2126);
nand U2686 (N_2686,N_42,N_2451);
nand U2687 (N_2687,N_2059,In_4591);
nor U2688 (N_2688,N_1998,N_1999);
nor U2689 (N_2689,In_4056,In_1979);
nand U2690 (N_2690,In_4714,N_1435);
or U2691 (N_2691,In_2677,N_736);
nand U2692 (N_2692,In_943,N_2258);
or U2693 (N_2693,In_4776,N_598);
nand U2694 (N_2694,N_2155,N_1919);
nor U2695 (N_2695,In_1074,N_2386);
and U2696 (N_2696,N_2393,N_39);
nand U2697 (N_2697,In_4630,N_2160);
or U2698 (N_2698,In_4281,N_2022);
or U2699 (N_2699,In_4091,N_1718);
and U2700 (N_2700,N_1812,N_2389);
and U2701 (N_2701,In_3740,N_964);
and U2702 (N_2702,In_424,N_1442);
nor U2703 (N_2703,In_1850,N_117);
nor U2704 (N_2704,N_2415,N_831);
nand U2705 (N_2705,In_3201,In_409);
and U2706 (N_2706,In_931,N_1819);
or U2707 (N_2707,In_3159,N_2147);
xnor U2708 (N_2708,N_1708,In_2090);
xor U2709 (N_2709,In_1296,In_4520);
nor U2710 (N_2710,In_4695,N_1885);
or U2711 (N_2711,N_710,In_3012);
or U2712 (N_2712,N_13,N_216);
nor U2713 (N_2713,N_2400,N_2361);
nor U2714 (N_2714,N_1561,N_2448);
xor U2715 (N_2715,In_2484,N_2271);
nand U2716 (N_2716,In_765,N_2333);
nand U2717 (N_2717,N_95,N_1607);
and U2718 (N_2718,In_4282,In_3124);
nor U2719 (N_2719,N_2434,N_2327);
and U2720 (N_2720,N_2046,N_1197);
nor U2721 (N_2721,N_2139,N_1633);
and U2722 (N_2722,N_1583,In_4464);
nor U2723 (N_2723,In_1643,N_1963);
or U2724 (N_2724,N_2390,N_2376);
or U2725 (N_2725,N_2191,In_4333);
and U2726 (N_2726,N_1245,N_1865);
or U2727 (N_2727,In_272,N_128);
nand U2728 (N_2728,N_761,N_1757);
and U2729 (N_2729,N_2304,N_1787);
and U2730 (N_2730,In_4819,N_1397);
nor U2731 (N_2731,N_1555,In_4268);
or U2732 (N_2732,In_3305,In_2772);
nand U2733 (N_2733,In_2947,N_602);
and U2734 (N_2734,N_1049,In_2563);
or U2735 (N_2735,In_1397,N_1009);
xnor U2736 (N_2736,N_2438,In_2601);
nand U2737 (N_2737,In_1133,N_2198);
nor U2738 (N_2738,N_2221,In_3451);
nor U2739 (N_2739,N_2202,In_4111);
and U2740 (N_2740,N_2476,In_4276);
nor U2741 (N_2741,N_1540,In_4769);
and U2742 (N_2742,In_4820,N_265);
nor U2743 (N_2743,N_919,N_2042);
and U2744 (N_2744,In_3248,In_4209);
xnor U2745 (N_2745,In_399,N_1338);
and U2746 (N_2746,In_112,In_3364);
or U2747 (N_2747,N_1180,N_1983);
or U2748 (N_2748,In_1135,N_2236);
nor U2749 (N_2749,In_4555,In_1787);
nor U2750 (N_2750,N_1313,N_673);
and U2751 (N_2751,In_4735,In_3503);
nor U2752 (N_2752,In_3624,N_2239);
and U2753 (N_2753,In_4006,N_527);
nand U2754 (N_2754,In_6,N_2398);
or U2755 (N_2755,In_1811,In_2887);
and U2756 (N_2756,N_2372,N_2146);
and U2757 (N_2757,In_3313,In_177);
nand U2758 (N_2758,In_632,N_881);
nand U2759 (N_2759,N_1933,In_3709);
xnor U2760 (N_2760,N_1523,N_2196);
nor U2761 (N_2761,In_653,N_2169);
or U2762 (N_2762,In_3946,N_1644);
nand U2763 (N_2763,N_2002,In_1488);
or U2764 (N_2764,N_2025,In_165);
nor U2765 (N_2765,In_1442,In_4698);
or U2766 (N_2766,N_846,In_462);
nor U2767 (N_2767,N_2185,N_2352);
and U2768 (N_2768,N_621,N_842);
nor U2769 (N_2769,In_3540,In_4614);
nand U2770 (N_2770,N_2427,N_1428);
nor U2771 (N_2771,In_3719,In_4375);
and U2772 (N_2772,In_3756,In_544);
nand U2773 (N_2773,In_32,N_2355);
nand U2774 (N_2774,N_1966,N_2484);
and U2775 (N_2775,N_2263,In_231);
or U2776 (N_2776,N_664,N_2061);
nand U2777 (N_2777,N_1460,N_2364);
nand U2778 (N_2778,In_2600,In_4400);
and U2779 (N_2779,In_4528,In_1948);
nand U2780 (N_2780,N_1498,In_1864);
nor U2781 (N_2781,In_4,In_2038);
and U2782 (N_2782,In_2754,N_2114);
nor U2783 (N_2783,N_1554,N_1172);
nand U2784 (N_2784,N_2200,N_484);
nor U2785 (N_2785,In_4136,In_4917);
and U2786 (N_2786,In_752,N_1518);
or U2787 (N_2787,N_1464,N_1793);
or U2788 (N_2788,N_2350,N_1867);
nand U2789 (N_2789,In_992,N_1123);
and U2790 (N_2790,In_4897,In_365);
or U2791 (N_2791,N_822,In_2356);
and U2792 (N_2792,N_2371,In_126);
nand U2793 (N_2793,N_2096,In_1291);
nor U2794 (N_2794,N_2430,N_2280);
nor U2795 (N_2795,N_2035,N_2011);
or U2796 (N_2796,In_3249,N_1528);
nand U2797 (N_2797,N_903,N_2033);
and U2798 (N_2798,In_1221,N_2443);
or U2799 (N_2799,N_1823,In_1633);
nand U2800 (N_2800,In_4164,N_1967);
and U2801 (N_2801,In_2644,N_213);
xnor U2802 (N_2802,N_2195,In_4572);
nand U2803 (N_2803,N_1093,N_2138);
and U2804 (N_2804,In_3388,N_1401);
nor U2805 (N_2805,N_289,N_2122);
or U2806 (N_2806,N_1544,N_2283);
nor U2807 (N_2807,In_3857,N_1287);
and U2808 (N_2808,In_4938,In_3562);
nor U2809 (N_2809,In_1848,N_1899);
nor U2810 (N_2810,In_1933,In_200);
xor U2811 (N_2811,N_1807,In_4014);
nand U2812 (N_2812,In_4895,N_2285);
and U2813 (N_2813,In_3577,In_282);
nand U2814 (N_2814,N_77,N_2245);
nand U2815 (N_2815,N_335,N_1446);
nand U2816 (N_2816,N_1840,In_2188);
or U2817 (N_2817,In_770,In_283);
nand U2818 (N_2818,N_1619,In_3340);
nand U2819 (N_2819,N_2057,N_2230);
nor U2820 (N_2820,N_1015,In_895);
nand U2821 (N_2821,N_754,In_646);
xnor U2822 (N_2822,N_564,N_2397);
or U2823 (N_2823,N_1799,N_806);
nor U2824 (N_2824,In_1422,N_1934);
or U2825 (N_2825,N_2306,N_2403);
nand U2826 (N_2826,In_4532,In_1954);
or U2827 (N_2827,In_1993,In_4853);
or U2828 (N_2828,In_4911,N_2163);
nand U2829 (N_2829,N_2092,N_395);
and U2830 (N_2830,N_2129,N_1562);
or U2831 (N_2831,N_2074,N_2123);
nand U2832 (N_2832,N_752,N_10);
nor U2833 (N_2833,N_1986,In_3488);
and U2834 (N_2834,In_556,In_1119);
nand U2835 (N_2835,In_3823,In_4992);
nand U2836 (N_2836,N_2422,N_2217);
nor U2837 (N_2837,N_2370,N_1835);
and U2838 (N_2838,In_3209,N_1129);
xor U2839 (N_2839,N_904,N_106);
or U2840 (N_2840,In_4473,N_1937);
nand U2841 (N_2841,N_836,In_3010);
and U2842 (N_2842,In_2938,N_1824);
nand U2843 (N_2843,N_1124,N_1400);
nor U2844 (N_2844,N_2334,In_4586);
nand U2845 (N_2845,In_4669,N_2465);
or U2846 (N_2846,N_1790,N_1707);
nor U2847 (N_2847,N_1593,N_1765);
nor U2848 (N_2848,N_945,In_849);
and U2849 (N_2849,In_1683,N_2284);
and U2850 (N_2850,N_152,N_2009);
nor U2851 (N_2851,N_2264,In_1177);
or U2852 (N_2852,In_2233,N_2282);
xor U2853 (N_2853,N_1862,N_2336);
nand U2854 (N_2854,In_3066,N_1520);
nor U2855 (N_2855,N_1295,N_1036);
nor U2856 (N_2856,In_1935,N_1018);
and U2857 (N_2857,N_992,N_2262);
nand U2858 (N_2858,In_3449,N_2479);
or U2859 (N_2859,N_1614,N_1837);
and U2860 (N_2860,N_2293,In_412);
and U2861 (N_2861,N_1144,In_582);
nand U2862 (N_2862,N_2193,In_4031);
nand U2863 (N_2863,N_1385,N_960);
nor U2864 (N_2864,N_658,In_156);
nor U2865 (N_2865,In_2002,In_2318);
nand U2866 (N_2866,In_815,N_2249);
xnor U2867 (N_2867,In_1368,N_631);
xor U2868 (N_2868,In_4309,In_3714);
or U2869 (N_2869,N_937,In_2808);
and U2870 (N_2870,N_1727,In_3529);
xor U2871 (N_2871,In_3493,N_2342);
nor U2872 (N_2872,In_1509,N_1491);
and U2873 (N_2873,N_2068,In_1138);
and U2874 (N_2874,In_2718,N_1229);
and U2875 (N_2875,N_2357,In_4817);
nand U2876 (N_2876,In_2093,N_2432);
nand U2877 (N_2877,N_1029,N_1978);
or U2878 (N_2878,In_2167,In_146);
nand U2879 (N_2879,N_2154,N_427);
xnor U2880 (N_2880,N_2081,In_2532);
and U2881 (N_2881,In_4694,N_2474);
or U2882 (N_2882,N_2450,N_442);
nand U2883 (N_2883,In_4102,N_2375);
nor U2884 (N_2884,In_4803,In_1362);
nor U2885 (N_2885,N_1682,N_1982);
nor U2886 (N_2886,N_1686,N_1742);
nor U2887 (N_2887,N_2170,In_3657);
nand U2888 (N_2888,N_208,N_1610);
and U2889 (N_2889,In_1822,In_514);
or U2890 (N_2890,N_1216,N_1759);
and U2891 (N_2891,In_4650,In_4558);
nand U2892 (N_2892,In_4956,N_204);
and U2893 (N_2893,In_4837,In_3856);
or U2894 (N_2894,N_993,In_1904);
nand U2895 (N_2895,N_503,N_2362);
or U2896 (N_2896,N_2358,N_1868);
nor U2897 (N_2897,N_839,N_2153);
nand U2898 (N_2898,In_4050,N_702);
or U2899 (N_2899,In_2598,N_2148);
xnor U2900 (N_2900,N_909,N_2072);
or U2901 (N_2901,In_3876,In_1827);
nand U2902 (N_2902,N_2054,N_2102);
or U2903 (N_2903,N_2183,N_2019);
and U2904 (N_2904,In_1029,N_1691);
and U2905 (N_2905,In_2436,N_2256);
nand U2906 (N_2906,N_1880,In_2825);
nor U2907 (N_2907,In_105,N_1089);
nor U2908 (N_2908,N_1078,N_2016);
or U2909 (N_2909,In_3834,N_2462);
nand U2910 (N_2910,N_2300,N_340);
or U2911 (N_2911,In_4483,In_4330);
and U2912 (N_2912,N_2247,N_2199);
nand U2913 (N_2913,N_1186,N_1304);
nand U2914 (N_2914,In_877,In_418);
nor U2915 (N_2915,In_4838,In_1366);
or U2916 (N_2916,N_2454,N_1798);
and U2917 (N_2917,N_2203,In_4692);
xor U2918 (N_2918,N_1848,In_2453);
nor U2919 (N_2919,N_1980,N_1901);
xor U2920 (N_2920,N_1255,In_747);
nand U2921 (N_2921,N_1472,In_3847);
and U2922 (N_2922,N_2001,In_1932);
nor U2923 (N_2923,N_907,N_1997);
nor U2924 (N_2924,N_2186,N_1143);
nor U2925 (N_2925,In_1003,In_2664);
or U2926 (N_2926,N_1139,N_755);
and U2927 (N_2927,N_2272,In_1407);
nand U2928 (N_2928,N_2062,In_0);
or U2929 (N_2929,N_2008,In_3466);
or U2930 (N_2930,N_544,N_1261);
xnor U2931 (N_2931,In_4552,N_2447);
nor U2932 (N_2932,N_1687,In_3815);
xnor U2933 (N_2933,In_4015,N_1608);
and U2934 (N_2934,N_1577,In_1671);
nand U2935 (N_2935,N_2223,In_2308);
and U2936 (N_2936,In_880,N_263);
xor U2937 (N_2937,In_3253,N_2497);
or U2938 (N_2938,N_2143,In_1634);
xor U2939 (N_2939,N_1743,In_1191);
or U2940 (N_2940,In_1059,N_220);
nand U2941 (N_2941,N_2289,N_175);
or U2942 (N_2942,N_1503,N_368);
nor U2943 (N_2943,N_1268,In_710);
nor U2944 (N_2944,N_963,N_1244);
and U2945 (N_2945,N_2329,N_908);
nand U2946 (N_2946,N_2227,N_2473);
or U2947 (N_2947,N_1662,N_2315);
and U2948 (N_2948,N_1994,In_2065);
nand U2949 (N_2949,In_3699,In_2043);
nand U2950 (N_2950,N_1500,N_2431);
or U2951 (N_2951,In_210,N_721);
xor U2952 (N_2952,N_2103,In_17);
nor U2953 (N_2953,N_1674,N_1371);
and U2954 (N_2954,N_2380,N_45);
xnor U2955 (N_2955,In_64,In_4185);
or U2956 (N_2956,N_2087,In_4348);
or U2957 (N_2957,In_4362,In_1533);
and U2958 (N_2958,N_2162,In_4676);
nor U2959 (N_2959,N_250,N_1046);
nand U2960 (N_2960,N_2365,In_870);
or U2961 (N_2961,N_642,N_624);
or U2962 (N_2962,In_2669,In_2102);
xor U2963 (N_2963,In_944,N_2338);
or U2964 (N_2964,In_1159,N_748);
or U2965 (N_2965,In_2522,N_2286);
or U2966 (N_2966,N_2482,N_285);
nor U2967 (N_2967,In_4192,N_1479);
or U2968 (N_2968,N_1714,N_1132);
nor U2969 (N_2969,In_1464,In_3695);
nor U2970 (N_2970,In_3137,N_2084);
nand U2971 (N_2971,N_2426,In_4365);
nand U2972 (N_2972,N_2456,N_1985);
nand U2973 (N_2973,N_1825,N_2322);
nor U2974 (N_2974,N_2324,In_4855);
nor U2975 (N_2975,N_2471,In_368);
and U2976 (N_2976,N_1905,N_2166);
nor U2977 (N_2977,In_1625,N_307);
nand U2978 (N_2978,In_2866,In_2502);
or U2979 (N_2979,N_1427,N_2383);
or U2980 (N_2980,In_3269,In_2998);
or U2981 (N_2981,N_1249,In_1523);
xnor U2982 (N_2982,N_685,N_1735);
nor U2983 (N_2983,In_4070,N_2151);
and U2984 (N_2984,In_1672,In_3199);
nor U2985 (N_2985,N_351,N_2056);
xor U2986 (N_2986,In_1877,N_1080);
or U2987 (N_2987,In_553,In_4002);
xor U2988 (N_2988,N_2120,In_3531);
and U2989 (N_2989,N_2392,N_1732);
or U2990 (N_2990,In_4482,N_1688);
nor U2991 (N_2991,In_1699,N_1564);
xor U2992 (N_2992,In_1114,In_4007);
and U2993 (N_2993,N_635,N_1745);
nand U2994 (N_2994,In_641,In_208);
or U2995 (N_2995,In_647,In_2536);
and U2996 (N_2996,N_1033,In_1630);
nor U2997 (N_2997,In_3724,In_2057);
and U2998 (N_2998,In_3328,N_2090);
nand U2999 (N_2999,In_2315,In_1473);
nor U3000 (N_3000,In_1941,N_2332);
nand U3001 (N_3001,N_532,N_1860);
nand U3002 (N_3002,In_1744,N_2960);
and U3003 (N_3003,N_984,N_181);
nor U3004 (N_3004,In_4250,N_1642);
or U3005 (N_3005,N_2678,N_2614);
or U3006 (N_3006,N_2373,In_2516);
nor U3007 (N_3007,In_3527,N_1752);
and U3008 (N_3008,N_121,N_2291);
nand U3009 (N_3009,N_2152,In_2986);
xor U3010 (N_3010,In_617,N_2496);
and U3011 (N_3011,N_1726,N_2854);
nand U3012 (N_3012,N_1191,N_878);
xnor U3013 (N_3013,N_1345,N_1831);
nand U3014 (N_3014,N_2545,In_593);
and U3015 (N_3015,N_2704,N_886);
or U3016 (N_3016,In_375,N_1324);
nor U3017 (N_3017,N_2989,In_4167);
or U3018 (N_3018,In_1846,N_2814);
nor U3019 (N_3019,N_2491,N_2328);
or U3020 (N_3020,N_2378,N_2337);
or U3021 (N_3021,N_2317,N_2866);
nor U3022 (N_3022,N_2550,In_1293);
xor U3023 (N_3023,N_1954,N_2601);
nand U3024 (N_3024,N_2341,N_2060);
nor U3025 (N_3025,N_2732,In_4480);
nor U3026 (N_3026,N_2527,N_2837);
and U3027 (N_3027,In_4795,N_2957);
nand U3028 (N_3028,In_3838,N_1871);
nor U3029 (N_3029,N_2174,N_2563);
nor U3030 (N_3030,N_419,N_2636);
and U3031 (N_3031,N_1242,In_2004);
and U3032 (N_3032,N_2739,N_1639);
or U3033 (N_3033,N_2741,N_2420);
and U3034 (N_3034,In_3101,N_2159);
and U3035 (N_3035,N_2696,N_1218);
or U3036 (N_3036,N_197,N_1506);
or U3037 (N_3037,N_2505,N_2698);
or U3038 (N_3038,N_2676,N_1391);
or U3039 (N_3039,N_1805,N_2526);
nand U3040 (N_3040,N_2569,N_2548);
xnor U3041 (N_3041,N_1948,N_2609);
nand U3042 (N_3042,In_3235,N_851);
xnor U3043 (N_3043,In_3563,In_726);
and U3044 (N_3044,In_2263,N_1192);
and U3045 (N_3045,In_792,N_2165);
nor U3046 (N_3046,N_616,N_2797);
or U3047 (N_3047,In_3161,N_2367);
xnor U3048 (N_3048,In_3727,N_1728);
or U3049 (N_3049,N_2790,N_2514);
nor U3050 (N_3050,N_2775,N_2785);
nand U3051 (N_3051,In_4965,N_2445);
nand U3052 (N_3052,N_1533,N_2882);
nor U3053 (N_3053,In_2096,In_3938);
or U3054 (N_3054,N_507,N_49);
or U3055 (N_3055,N_2624,In_3008);
xnor U3056 (N_3056,N_147,In_3786);
nor U3057 (N_3057,N_1035,In_3093);
and U3058 (N_3058,N_1334,N_2515);
and U3059 (N_3059,N_949,N_2974);
and U3060 (N_3060,N_1087,N_2855);
xor U3061 (N_3061,N_1212,In_447);
xnor U3062 (N_3062,N_2973,N_381);
and U3063 (N_3063,In_3649,N_2194);
nor U3064 (N_3064,In_1915,In_2860);
and U3065 (N_3065,In_473,In_3366);
nor U3066 (N_3066,N_1598,N_2485);
and U3067 (N_3067,N_2530,N_2353);
and U3068 (N_3068,N_2209,N_1189);
nor U3069 (N_3069,In_1807,In_331);
and U3070 (N_3070,N_2547,In_1829);
and U3071 (N_3071,N_2903,N_2297);
nand U3072 (N_3072,In_4536,In_2581);
and U3073 (N_3073,In_489,In_1165);
and U3074 (N_3074,N_2881,In_423);
nand U3075 (N_3075,N_2277,N_2310);
xnor U3076 (N_3076,In_2013,N_2736);
nor U3077 (N_3077,N_2738,N_2347);
or U3078 (N_3078,In_2157,In_381);
and U3079 (N_3079,N_1454,In_4740);
nor U3080 (N_3080,N_2664,N_912);
nand U3081 (N_3081,N_998,In_3795);
and U3082 (N_3082,In_636,In_2144);
xnor U3083 (N_3083,N_2187,In_2529);
xor U3084 (N_3084,In_3538,In_4368);
nor U3085 (N_3085,In_273,In_2164);
nand U3086 (N_3086,N_2274,N_726);
and U3087 (N_3087,N_2119,N_592);
nand U3088 (N_3088,In_4901,In_2031);
or U3089 (N_3089,In_2055,N_1647);
or U3090 (N_3090,N_107,In_1840);
nand U3091 (N_3091,N_2840,N_509);
or U3092 (N_3092,N_2612,N_1782);
and U3093 (N_3093,N_1364,N_2313);
nor U3094 (N_3094,N_2339,N_2117);
nand U3095 (N_3095,N_888,N_2546);
nor U3096 (N_3096,N_1361,N_2786);
and U3097 (N_3097,N_2591,N_1466);
or U3098 (N_3098,N_2553,N_2662);
nor U3099 (N_3099,N_2288,In_2040);
nor U3100 (N_3100,N_694,N_2675);
nor U3101 (N_3101,In_1092,N_1762);
nor U3102 (N_3102,In_4344,In_832);
and U3103 (N_3103,N_2733,N_2730);
nand U3104 (N_3104,N_2053,N_1493);
nand U3105 (N_3105,N_2003,N_2604);
and U3106 (N_3106,N_2769,N_2919);
nor U3107 (N_3107,In_1514,N_2125);
xnor U3108 (N_3108,N_2959,N_35);
and U3109 (N_3109,N_2097,N_2029);
nor U3110 (N_3110,In_1305,N_2499);
nor U3111 (N_3111,In_898,In_2759);
and U3112 (N_3112,N_2537,N_2627);
nor U3113 (N_3113,In_2810,In_1174);
nand U3114 (N_3114,N_2630,In_1449);
or U3115 (N_3115,In_4693,N_2177);
or U3116 (N_3116,In_2702,N_940);
and U3117 (N_3117,N_2475,N_2985);
or U3118 (N_3118,In_4046,In_2401);
nand U3119 (N_3119,N_2921,N_2737);
nor U3120 (N_3120,N_1881,In_3168);
or U3121 (N_3121,N_1019,N_957);
nor U3122 (N_3122,N_127,N_2314);
and U3123 (N_3123,In_3934,N_1156);
xnor U3124 (N_3124,In_2174,N_2708);
nand U3125 (N_3125,N_2320,In_1117);
nand U3126 (N_3126,In_1448,In_1316);
and U3127 (N_3127,N_2772,In_3481);
and U3128 (N_3128,In_222,N_2575);
nand U3129 (N_3129,In_1471,N_2818);
nand U3130 (N_3130,N_1052,In_1753);
and U3131 (N_3131,N_973,N_612);
nand U3132 (N_3132,N_2622,N_1386);
and U3133 (N_3133,N_2746,In_963);
and U3134 (N_3134,N_2596,N_2616);
or U3135 (N_3135,In_2624,In_2652);
and U3136 (N_3136,N_1894,In_3372);
xnor U3137 (N_3137,N_1008,N_2374);
nor U3138 (N_3138,N_2175,N_1828);
or U3139 (N_3139,In_1873,N_2613);
nand U3140 (N_3140,N_2858,N_2140);
and U3141 (N_3141,In_2734,N_1060);
or U3142 (N_3142,N_2954,In_2771);
or U3143 (N_3143,In_4839,N_2345);
xor U3144 (N_3144,N_2441,N_2998);
or U3145 (N_3145,N_2213,In_4622);
nor U3146 (N_3146,N_2007,N_1455);
nand U3147 (N_3147,N_2595,N_2416);
nor U3148 (N_3148,N_1299,In_989);
nor U3149 (N_3149,In_1805,In_175);
xnor U3150 (N_3150,N_2510,In_2723);
nand U3151 (N_3151,In_4320,In_4487);
nor U3152 (N_3152,N_11,In_475);
nor U3153 (N_3153,N_2150,In_4019);
and U3154 (N_3154,N_2673,N_2815);
and U3155 (N_3155,N_2765,N_1050);
and U3156 (N_3156,In_2748,In_741);
nand U3157 (N_3157,In_2458,N_2860);
nand U3158 (N_3158,N_2780,N_1101);
nor U3159 (N_3159,N_2109,In_1016);
nor U3160 (N_3160,In_2237,In_818);
nand U3161 (N_3161,In_1462,N_2326);
nand U3162 (N_3162,N_22,In_430);
and U3163 (N_3163,N_2650,N_2939);
nand U3164 (N_3164,N_2394,N_1887);
and U3165 (N_3165,N_2265,N_2799);
and U3166 (N_3166,N_2911,In_2249);
nand U3167 (N_3167,N_2864,In_3497);
nand U3168 (N_3168,N_2767,N_349);
and U3169 (N_3169,N_2651,N_1748);
or U3170 (N_3170,In_3666,N_2648);
and U3171 (N_3171,N_1861,N_2684);
and U3172 (N_3172,N_628,N_2665);
or U3173 (N_3173,In_3430,In_1238);
and U3174 (N_3174,In_4828,N_545);
nand U3175 (N_3175,N_334,N_2124);
and U3176 (N_3176,N_2190,In_4078);
or U3177 (N_3177,N_1278,N_630);
or U3178 (N_3178,N_1764,N_2133);
nor U3179 (N_3179,N_2085,In_1493);
or U3180 (N_3180,In_1897,N_2838);
nand U3181 (N_3181,In_4659,In_1199);
nand U3182 (N_3182,N_2525,N_2623);
or U3183 (N_3183,In_3869,N_2834);
xnor U3184 (N_3184,N_980,N_2625);
or U3185 (N_3185,N_270,N_1930);
nand U3186 (N_3186,N_2590,In_179);
and U3187 (N_3187,N_2760,In_3966);
nand U3188 (N_3188,N_2880,In_3088);
nand U3189 (N_3189,N_2783,In_4773);
or U3190 (N_3190,N_2995,In_3513);
xor U3191 (N_3191,N_2851,In_4751);
nor U3192 (N_3192,In_181,In_151);
or U3193 (N_3193,In_4479,In_3693);
nand U3194 (N_3194,N_1672,N_2711);
xnor U3195 (N_3195,N_1329,N_2559);
nor U3196 (N_3196,In_1139,In_3414);
nor U3197 (N_3197,N_2926,In_3526);
or U3198 (N_3198,N_2823,In_3162);
nor U3199 (N_3199,N_2218,N_1979);
and U3200 (N_3200,N_56,In_3785);
or U3201 (N_3201,N_14,N_1311);
or U3202 (N_3202,N_295,N_2076);
or U3203 (N_3203,N_2049,N_2870);
xnor U3204 (N_3204,N_2955,In_3694);
and U3205 (N_3205,N_2246,In_1842);
xnor U3206 (N_3206,N_1671,N_1196);
nor U3207 (N_3207,N_1421,N_2493);
xor U3208 (N_3208,In_3942,In_1524);
and U3209 (N_3209,In_2524,N_2705);
or U3210 (N_3210,N_1310,In_311);
nor U3211 (N_3211,N_1473,N_2094);
or U3212 (N_3212,N_2901,In_1022);
nor U3213 (N_3213,N_38,In_3074);
xor U3214 (N_3214,In_73,In_1252);
or U3215 (N_3215,In_3095,N_2587);
nand U3216 (N_3216,N_2747,N_2889);
nor U3217 (N_3217,In_2770,N_2887);
or U3218 (N_3218,N_2461,N_2902);
nand U3219 (N_3219,In_1253,In_2867);
and U3220 (N_3220,N_2961,N_1107);
or U3221 (N_3221,In_4103,N_2157);
nor U3222 (N_3222,N_1953,N_2429);
nor U3223 (N_3223,N_2107,In_4686);
xnor U3224 (N_3224,In_4311,N_394);
xnor U3225 (N_3225,N_1569,N_1845);
nor U3226 (N_3226,In_4384,In_2611);
and U3227 (N_3227,N_149,N_2298);
nor U3228 (N_3228,N_2558,N_2744);
xnor U3229 (N_3229,N_2044,N_1140);
nand U3230 (N_3230,In_860,N_2577);
and U3231 (N_3231,N_2801,N_2778);
nor U3232 (N_3232,N_1053,N_1543);
nor U3233 (N_3233,N_2584,N_634);
and U3234 (N_3234,N_686,N_2714);
or U3235 (N_3235,N_2252,N_2210);
nand U3236 (N_3236,In_621,N_1851);
nor U3237 (N_3237,N_2894,N_2633);
nor U3238 (N_3238,N_2539,N_2774);
nand U3239 (N_3239,N_1000,N_1623);
nand U3240 (N_3240,N_899,N_640);
or U3241 (N_3241,N_1977,N_2131);
xor U3242 (N_3242,In_1056,N_1615);
and U3243 (N_3243,N_563,In_4995);
nor U3244 (N_3244,In_2790,N_1722);
and U3245 (N_3245,In_2786,N_1436);
or U3246 (N_3246,N_2947,N_63);
and U3247 (N_3247,In_4256,In_738);
and U3248 (N_3248,N_1621,N_1700);
nor U3249 (N_3249,In_2668,In_2805);
and U3250 (N_3250,N_644,N_1929);
nand U3251 (N_3251,N_1001,N_1992);
or U3252 (N_3252,N_2551,N_391);
and U3253 (N_3253,N_2906,In_2245);
and U3254 (N_3254,In_4066,N_1768);
nand U3255 (N_3255,In_4115,In_1764);
xnor U3256 (N_3256,In_4653,N_1349);
nand U3257 (N_3257,In_1158,N_2861);
and U3258 (N_3258,In_1244,N_2164);
nor U3259 (N_3259,N_1910,In_242);
nor U3260 (N_3260,In_2184,N_2892);
or U3261 (N_3261,N_2619,In_1115);
or U3262 (N_3262,N_1818,In_930);
and U3263 (N_3263,In_4929,N_2405);
nand U3264 (N_3264,In_1591,N_1842);
nor U3265 (N_3265,N_2663,In_1894);
and U3266 (N_3266,In_4788,N_2417);
or U3267 (N_3267,N_2690,N_1097);
xnor U3268 (N_3268,N_2418,N_2523);
or U3269 (N_3269,N_2568,In_3653);
nand U3270 (N_3270,In_4535,N_575);
and U3271 (N_3271,In_1430,N_2808);
nor U3272 (N_3272,In_625,In_4609);
nand U3273 (N_3273,N_2924,In_33);
nand U3274 (N_3274,N_2682,N_1928);
nand U3275 (N_3275,N_396,In_2130);
or U3276 (N_3276,N_2030,N_2745);
nor U3277 (N_3277,N_469,N_2171);
nand U3278 (N_3278,In_2714,In_3596);
or U3279 (N_3279,In_947,N_684);
or U3280 (N_3280,N_2843,N_2984);
xnor U3281 (N_3281,In_1574,N_2791);
or U3282 (N_3282,N_1181,In_3282);
or U3283 (N_3283,N_2798,N_2695);
and U3284 (N_3284,In_1047,In_1706);
nor U3285 (N_3285,N_2401,N_1751);
and U3286 (N_3286,N_2020,In_2555);
nor U3287 (N_3287,In_3914,In_2178);
nor U3288 (N_3288,In_2142,N_1348);
xor U3289 (N_3289,N_2560,In_1766);
nor U3290 (N_3290,N_680,In_4506);
or U3291 (N_3291,In_4463,N_2588);
nand U3292 (N_3292,In_1120,N_2034);
nand U3293 (N_3293,In_585,In_3471);
nand U3294 (N_3294,In_502,N_728);
nor U3295 (N_3295,N_2406,N_1653);
or U3296 (N_3296,N_2912,N_2172);
and U3297 (N_3297,N_1492,N_2807);
nor U3298 (N_3298,In_2688,N_1404);
nand U3299 (N_3299,In_1512,In_1561);
nor U3300 (N_3300,In_2003,In_3770);
or U3301 (N_3301,N_1791,N_1843);
nor U3302 (N_3302,In_839,N_2212);
and U3303 (N_3303,In_1927,N_2874);
nand U3304 (N_3304,In_1405,N_2436);
or U3305 (N_3305,In_4372,N_2071);
xnor U3306 (N_3306,N_2972,N_2752);
nand U3307 (N_3307,N_784,N_201);
or U3308 (N_3308,In_4234,N_753);
or U3309 (N_3309,In_3681,N_2694);
and U3310 (N_3310,N_129,N_17);
or U3311 (N_3311,N_1432,In_2427);
nand U3312 (N_3312,N_2991,In_2299);
nor U3313 (N_3313,N_2573,N_2078);
nor U3314 (N_3314,N_2999,In_2435);
and U3315 (N_3315,N_1051,N_2653);
nor U3316 (N_3316,N_2824,N_1800);
or U3317 (N_3317,N_2869,N_1654);
nor U3318 (N_3318,In_3470,In_28);
nand U3319 (N_3319,N_1496,N_2835);
or U3320 (N_3320,N_2224,N_2992);
nor U3321 (N_3321,N_287,In_4068);
and U3322 (N_3322,N_2917,In_1573);
and U3323 (N_3323,N_1021,N_2743);
or U3324 (N_3324,N_1566,N_1931);
nand U3325 (N_3325,In_1007,N_1303);
and U3326 (N_3326,N_2532,N_2883);
nand U3327 (N_3327,N_1553,In_2277);
xor U3328 (N_3328,In_4826,N_2453);
or U3329 (N_3329,N_2900,In_3143);
or U3330 (N_3330,In_1995,N_2877);
and U3331 (N_3331,In_2592,In_639);
and U3332 (N_3332,In_2956,In_4286);
nand U3333 (N_3333,In_2314,N_614);
or U3334 (N_3334,N_1105,N_2751);
nand U3335 (N_3335,N_2830,In_1456);
nand U3336 (N_3336,In_2649,N_1044);
and U3337 (N_3337,N_2031,N_2968);
and U3338 (N_3338,N_1941,In_2302);
nor U3339 (N_3339,In_2778,N_2937);
nor U3340 (N_3340,N_2399,N_2610);
and U3341 (N_3341,In_4409,N_2089);
nor U3342 (N_3342,N_2885,In_1831);
or U3343 (N_3343,N_2793,N_2982);
and U3344 (N_3344,N_1077,In_3085);
nand U3345 (N_3345,N_499,In_13);
or U3346 (N_3346,In_3309,In_1653);
and U3347 (N_3347,N_1526,N_2520);
nor U3348 (N_3348,N_144,N_2026);
nand U3349 (N_3349,In_4709,N_2275);
and U3350 (N_3350,N_436,N_2773);
nand U3351 (N_3351,N_1990,N_2161);
and U3352 (N_3352,N_700,In_1402);
nand U3353 (N_3353,In_176,N_2606);
and U3354 (N_3354,In_3109,N_1724);
or U3355 (N_3355,In_253,N_2077);
nand U3356 (N_3356,N_2857,N_2439);
and U3357 (N_3357,N_2608,N_1817);
nand U3358 (N_3358,In_2755,N_2949);
nor U3359 (N_3359,N_2729,In_4321);
or U3360 (N_3360,N_2032,N_2534);
nand U3361 (N_3361,N_2391,In_2670);
nor U3362 (N_3362,In_910,N_950);
and U3363 (N_3363,In_301,N_2875);
nand U3364 (N_3364,In_2092,N_1411);
and U3365 (N_3365,N_2776,In_4160);
or U3366 (N_3366,N_2712,N_2934);
nand U3367 (N_3367,In_2578,N_475);
nand U3368 (N_3368,In_562,N_1547);
or U3369 (N_3369,In_4613,N_195);
or U3370 (N_3370,In_4294,N_808);
nand U3371 (N_3371,N_2023,N_2423);
and U3372 (N_3372,In_2925,N_2580);
nand U3373 (N_3373,N_1802,In_1675);
and U3374 (N_3374,N_2916,N_2014);
or U3375 (N_3375,In_1048,In_4702);
and U3376 (N_3376,N_2142,N_2652);
nand U3377 (N_3377,N_626,In_679);
nand U3378 (N_3378,In_2788,In_2900);
or U3379 (N_3379,In_4948,N_2516);
and U3380 (N_3380,N_2255,N_2859);
and U3381 (N_3381,N_1972,N_2710);
and U3382 (N_3382,N_2997,N_2585);
or U3383 (N_3383,In_1821,In_1950);
and U3384 (N_3384,N_2253,In_3264);
and U3385 (N_3385,N_1776,N_573);
or U3386 (N_3386,N_2589,In_221);
nand U3387 (N_3387,N_2388,In_543);
or U3388 (N_3388,In_2365,N_2467);
xnor U3389 (N_3389,N_2723,N_2554);
xnor U3390 (N_3390,N_1624,N_2920);
nor U3391 (N_3391,In_4472,In_2215);
nor U3392 (N_3392,In_1103,N_1649);
nand U3393 (N_3393,N_2829,In_845);
xnor U3394 (N_3394,In_4730,N_2728);
or U3395 (N_3395,N_2945,N_1916);
and U3396 (N_3396,N_2490,N_1959);
xor U3397 (N_3397,In_1152,N_2971);
and U3398 (N_3398,In_4043,N_2344);
and U3399 (N_3399,N_2535,N_1309);
xor U3400 (N_3400,In_3009,N_1942);
or U3401 (N_3401,N_2079,N_2144);
nor U3402 (N_3402,N_2862,N_1874);
nor U3403 (N_3403,N_2771,N_1918);
nand U3404 (N_3404,N_2492,N_2368);
and U3405 (N_3405,N_884,In_3943);
nor U3406 (N_3406,N_2909,N_2135);
nand U3407 (N_3407,N_200,In_3950);
nor U3408 (N_3408,In_4527,N_1501);
or U3409 (N_3409,N_2599,N_2540);
nand U3410 (N_3410,N_1134,In_1002);
nor U3411 (N_3411,N_2931,In_2955);
or U3412 (N_3412,N_2270,N_1174);
nor U3413 (N_3413,N_1103,N_2907);
nor U3414 (N_3414,N_2976,N_2457);
nand U3415 (N_3415,In_1336,In_1667);
xnor U3416 (N_3416,N_1922,In_2905);
nand U3417 (N_3417,In_1830,N_2309);
nor U3418 (N_3418,N_2895,N_1072);
nor U3419 (N_3419,In_396,N_291);
nand U3420 (N_3420,N_2672,In_427);
and U3421 (N_3421,In_4369,In_2113);
and U3422 (N_3422,In_149,In_728);
and U3423 (N_3423,In_4270,In_4345);
and U3424 (N_3424,N_745,N_4);
nor U3425 (N_3425,In_1544,In_1213);
or U3426 (N_3426,N_2301,N_2259);
or U3427 (N_3427,N_2890,In_3450);
nor U3428 (N_3428,N_2586,In_4936);
nand U3429 (N_3429,In_2933,N_2066);
nor U3430 (N_3430,In_2715,N_462);
or U3431 (N_3431,N_3,N_1541);
and U3432 (N_3432,In_1363,N_2458);
nand U3433 (N_3433,In_2025,N_1631);
xor U3434 (N_3434,In_4144,In_4249);
and U3435 (N_3435,N_2437,N_2566);
xor U3436 (N_3436,In_4861,In_4860);
nor U3437 (N_3437,N_502,N_1806);
and U3438 (N_3438,N_1936,In_2190);
nor U3439 (N_3439,In_131,N_2531);
and U3440 (N_3440,N_2446,N_143);
nor U3441 (N_3441,N_2028,N_1739);
and U3442 (N_3442,N_2552,N_315);
xnor U3443 (N_3443,N_1112,In_3361);
and U3444 (N_3444,In_1345,N_2940);
or U3445 (N_3445,N_1059,N_1031);
xor U3446 (N_3446,N_2038,In_2404);
xnor U3447 (N_3447,N_2768,N_1380);
and U3448 (N_3448,In_2513,N_966);
and U3449 (N_3449,In_1294,N_1878);
xnor U3450 (N_3450,In_3969,N_2749);
nor U3451 (N_3451,N_2679,In_1292);
nor U3452 (N_3452,N_867,N_2668);
or U3453 (N_3453,In_3539,N_1573);
nor U3454 (N_3454,N_1648,N_2702);
nor U3455 (N_3455,In_4226,In_3030);
nand U3456 (N_3456,N_2444,In_1438);
nand U3457 (N_3457,N_838,N_2758);
xnor U3458 (N_3458,N_2952,N_139);
and U3459 (N_3459,In_2447,N_1468);
nand U3460 (N_3460,N_1567,In_4203);
and U3461 (N_3461,N_2176,N_2602);
nand U3462 (N_3462,N_727,N_2043);
nand U3463 (N_3463,N_339,N_2656);
nor U3464 (N_3464,N_2899,In_4913);
nor U3465 (N_3465,N_1645,N_2409);
xnor U3466 (N_3466,N_1673,In_1586);
and U3467 (N_3467,N_2833,N_2757);
nor U3468 (N_3468,N_2543,N_1665);
nand U3469 (N_3469,N_2788,N_820);
and U3470 (N_3470,N_259,In_1847);
nand U3471 (N_3471,N_146,In_58);
or U3472 (N_3472,N_2052,N_1327);
and U3473 (N_3473,N_1679,N_2118);
and U3474 (N_3474,N_1118,N_1925);
xnor U3475 (N_3475,N_2617,N_2522);
nand U3476 (N_3476,N_2179,In_1010);
nand U3477 (N_3477,N_2914,N_2459);
nand U3478 (N_3478,In_2159,N_2740);
xor U3479 (N_3479,N_2211,N_2943);
xnor U3480 (N_3480,In_1317,In_2080);
nand U3481 (N_3481,In_4619,N_385);
xnor U3482 (N_3482,N_1525,N_2250);
nor U3483 (N_3483,N_2478,N_782);
or U3484 (N_3484,N_2167,In_953);
nand U3485 (N_3485,In_63,N_2764);
or U3486 (N_3486,N_2561,In_3525);
xor U3487 (N_3487,N_2626,N_788);
and U3488 (N_3488,In_2300,In_2246);
or U3489 (N_3489,N_714,N_1213);
or U3490 (N_3490,In_1911,N_789);
nor U3491 (N_3491,In_2430,N_2583);
nand U3492 (N_3492,N_2518,N_2820);
or U3493 (N_3493,N_1810,In_3373);
nand U3494 (N_3494,N_2000,N_1149);
or U3495 (N_3495,N_1578,N_2075);
nand U3496 (N_3496,N_2929,N_2888);
nand U3497 (N_3497,N_1014,N_533);
nor U3498 (N_3498,N_2556,N_1678);
nand U3499 (N_3499,N_1264,In_1064);
and U3500 (N_3500,N_3375,N_623);
or U3501 (N_3501,N_3063,N_1502);
or U3502 (N_3502,N_1903,In_1968);
nand U3503 (N_3503,N_2727,N_2509);
nor U3504 (N_3504,In_4957,N_553);
or U3505 (N_3505,N_2942,N_3024);
nand U3506 (N_3506,N_172,In_2658);
xor U3507 (N_3507,In_372,N_3138);
and U3508 (N_3508,N_2396,N_2064);
and U3509 (N_3509,N_3343,N_2635);
nor U3510 (N_3510,N_1628,N_3378);
nor U3511 (N_3511,N_2618,N_3048);
or U3512 (N_3512,N_3436,N_3178);
nor U3513 (N_3513,N_2994,N_1911);
and U3514 (N_3514,N_3182,N_2382);
or U3515 (N_3515,N_1220,N_3491);
or U3516 (N_3516,N_2237,N_1844);
nor U3517 (N_3517,N_3324,N_2302);
xnor U3518 (N_3518,N_3265,N_3194);
nand U3519 (N_3519,N_3073,In_2727);
xnor U3520 (N_3520,N_3101,N_301);
or U3521 (N_3521,N_3159,N_1071);
nand U3522 (N_3522,In_2027,N_3007);
nand U3523 (N_3523,N_2506,N_3109);
xnor U3524 (N_3524,N_245,N_3311);
and U3525 (N_3525,N_2188,N_2047);
xor U3526 (N_3526,N_2065,In_665);
or U3527 (N_3527,N_3074,N_2878);
nor U3528 (N_3528,N_3360,In_3200);
or U3529 (N_3529,N_2628,N_407);
nor U3530 (N_3530,N_104,In_4821);
xor U3531 (N_3531,N_79,N_1413);
nand U3532 (N_3532,N_3302,N_1777);
or U3533 (N_3533,N_578,N_3249);
and U3534 (N_3534,N_3191,N_3288);
nor U3535 (N_3535,N_2754,N_2115);
or U3536 (N_3536,N_3463,N_3117);
nor U3537 (N_3537,N_3467,In_2387);
and U3538 (N_3538,In_3190,N_2410);
and U3539 (N_3539,In_1947,N_3286);
and U3540 (N_3540,N_3499,N_3030);
or U3541 (N_3541,N_2680,N_3268);
or U3542 (N_3542,N_2978,N_3089);
and U3543 (N_3543,N_2719,N_1864);
nor U3544 (N_3544,N_3243,N_3216);
nor U3545 (N_3545,N_3331,N_3424);
and U3546 (N_3546,N_3239,N_2825);
or U3547 (N_3547,N_3257,N_895);
or U3548 (N_3548,N_3457,In_994);
nand U3549 (N_3549,In_4894,N_2876);
nand U3550 (N_3550,N_3435,N_772);
and U3551 (N_3551,In_2463,N_2241);
or U3552 (N_3552,N_2442,N_3279);
nand U3553 (N_3553,N_3422,N_2544);
or U3554 (N_3554,N_1669,N_3021);
nor U3555 (N_3555,N_3460,N_2260);
or U3556 (N_3556,N_3221,In_3147);
nor U3557 (N_3557,N_2242,N_3472);
or U3558 (N_3558,N_3176,N_3177);
nor U3559 (N_3559,N_1225,N_657);
and U3560 (N_3560,In_1595,N_2642);
xnor U3561 (N_3561,N_2104,In_1652);
nand U3562 (N_3562,N_582,N_2639);
or U3563 (N_3563,N_3461,N_1452);
or U3564 (N_3564,In_3619,N_2149);
and U3565 (N_3565,N_1989,In_3547);
nand U3566 (N_3566,N_594,N_80);
nand U3567 (N_3567,N_1677,N_1133);
xor U3568 (N_3568,N_3130,In_987);
xor U3569 (N_3569,In_3362,N_184);
and U3570 (N_3570,N_2233,N_3372);
nand U3571 (N_3571,N_2988,N_1596);
nor U3572 (N_3572,N_913,N_2655);
and U3573 (N_3573,N_852,N_2716);
or U3574 (N_3574,N_1521,N_3044);
and U3575 (N_3575,In_2360,N_2641);
or U3576 (N_3576,N_2321,N_473);
or U3577 (N_3577,N_2963,N_1265);
nor U3578 (N_3578,N_3273,N_3416);
and U3579 (N_3579,N_411,N_1422);
nor U3580 (N_3580,N_3059,In_249);
or U3581 (N_3581,In_1347,N_2781);
or U3582 (N_3582,In_4292,N_2597);
and U3583 (N_3583,In_4623,In_2276);
and U3584 (N_3584,In_286,N_3437);
or U3585 (N_3585,In_3511,In_134);
nor U3586 (N_3586,N_1388,N_2363);
xor U3587 (N_3587,N_3125,N_725);
nand U3588 (N_3588,N_31,N_1091);
nor U3589 (N_3589,N_3084,In_377);
or U3590 (N_3590,N_3404,N_1104);
nor U3591 (N_3591,N_3040,N_3202);
or U3592 (N_3592,N_3248,N_418);
nor U3593 (N_3593,N_2503,N_2184);
nor U3594 (N_3594,In_3703,N_2987);
nand U3595 (N_3595,N_2564,N_2273);
or U3596 (N_3596,N_2936,In_1106);
nand U3597 (N_3597,N_3152,N_2826);
nand U3598 (N_3598,N_2802,N_3026);
and U3599 (N_3599,In_2857,N_3384);
nor U3600 (N_3600,N_2021,N_1923);
or U3601 (N_3601,In_3781,N_2480);
nor U3602 (N_3602,N_3079,N_2225);
or U3603 (N_3603,N_3261,N_3471);
nand U3604 (N_3604,N_1605,In_1747);
nand U3605 (N_3605,N_1613,N_2879);
or U3606 (N_3606,In_3316,In_318);
nand U3607 (N_3607,N_3396,N_1780);
or U3608 (N_3608,N_3284,In_4156);
and U3609 (N_3609,N_150,In_4072);
xnor U3610 (N_3610,N_3344,N_3185);
or U3611 (N_3611,In_2807,N_3345);
or U3612 (N_3612,In_3836,N_3387);
and U3613 (N_3613,N_2905,In_894);
or U3614 (N_3614,N_2570,In_2980);
or U3615 (N_3615,N_2750,N_3038);
and U3616 (N_3616,N_2958,N_834);
or U3617 (N_3617,N_520,N_2488);
or U3618 (N_3618,N_3095,In_2548);
or U3619 (N_3619,N_1214,In_439);
or U3620 (N_3620,N_2922,N_3015);
nor U3621 (N_3621,In_2708,N_2755);
or U3622 (N_3622,N_3359,N_2643);
nand U3623 (N_3623,N_2850,N_1461);
nor U3624 (N_3624,N_3153,In_92);
nor U3625 (N_3625,N_3490,N_2925);
and U3626 (N_3626,N_1689,N_775);
xor U3627 (N_3627,N_1785,N_1856);
nand U3628 (N_3628,In_525,In_3568);
or U3629 (N_3629,N_1640,In_3721);
nand U3630 (N_3630,N_1165,N_3293);
nor U3631 (N_3631,N_3212,In_4811);
xnor U3632 (N_3632,N_3025,N_1509);
nand U3633 (N_3633,N_2966,In_2794);
or U3634 (N_3634,N_1854,N_3318);
and U3635 (N_3635,N_3033,N_2671);
and U3636 (N_3636,N_1390,In_3528);
xnor U3637 (N_3637,N_3004,N_1811);
nor U3638 (N_3638,N_3148,N_3126);
nand U3639 (N_3639,N_2717,N_2234);
xnor U3640 (N_3640,N_2720,N_3215);
nor U3641 (N_3641,N_1778,N_3381);
or U3642 (N_3642,N_3433,In_2440);
nor U3643 (N_3643,N_2809,N_311);
or U3644 (N_3644,In_237,In_3059);
nand U3645 (N_3645,N_3190,N_3136);
or U3646 (N_3646,In_2749,N_3393);
or U3647 (N_3647,N_3327,N_1147);
nor U3648 (N_3648,In_3292,N_3298);
or U3649 (N_3649,N_3162,N_3081);
nand U3650 (N_3650,N_1126,In_3555);
nand U3651 (N_3651,N_3401,N_3366);
xnor U3652 (N_3652,N_199,N_3354);
or U3653 (N_3653,N_3304,N_1458);
and U3654 (N_3654,N_3458,In_1610);
nand U3655 (N_3655,N_1378,N_666);
or U3656 (N_3656,N_2069,N_3093);
nand U3657 (N_3657,N_2360,N_2354);
xnor U3658 (N_3658,N_2693,N_2951);
or U3659 (N_3659,N_2621,N_652);
or U3660 (N_3660,N_2735,In_85);
or U3661 (N_3661,N_3488,In_4392);
and U3662 (N_3662,N_2756,N_1927);
nand U3663 (N_3663,In_2861,N_3452);
nor U3664 (N_3664,In_2250,N_2969);
and U3665 (N_3665,N_2782,N_2965);
or U3666 (N_3666,N_2311,N_2967);
nor U3667 (N_3667,N_586,In_1040);
and U3668 (N_3668,In_2604,N_2779);
xnor U3669 (N_3669,N_2086,N_3484);
and U3670 (N_3670,N_3385,N_2173);
and U3671 (N_3671,N_603,N_3277);
nand U3672 (N_3672,N_3353,N_3080);
nand U3673 (N_3673,N_2521,N_3468);
or U3674 (N_3674,N_2494,N_3065);
and U3675 (N_3675,N_1337,N_2821);
and U3676 (N_3676,N_2897,N_1226);
nor U3677 (N_3677,N_3407,N_2842);
nor U3678 (N_3678,In_4756,In_1255);
and U3679 (N_3679,N_1859,In_824);
or U3680 (N_3680,N_2603,N_1760);
or U3681 (N_3681,In_2949,In_2307);
and U3682 (N_3682,In_919,In_1306);
nor U3683 (N_3683,N_1652,N_3189);
nand U3684 (N_3684,N_3266,In_1333);
and U3685 (N_3685,In_2459,N_3446);
nand U3686 (N_3686,N_3195,In_4410);
nand U3687 (N_3687,In_3029,In_1504);
nand U3688 (N_3688,N_3037,N_3132);
nand U3689 (N_3689,N_3290,N_2425);
nor U3690 (N_3690,In_3592,N_3019);
nand U3691 (N_3691,N_3192,N_942);
and U3692 (N_3692,N_1067,N_2677);
xnor U3693 (N_3693,N_1522,In_1649);
nor U3694 (N_3694,In_4316,N_3333);
nor U3695 (N_3695,In_3840,N_3218);
or U3696 (N_3696,N_2099,N_3225);
xor U3697 (N_3697,N_2819,In_3094);
nand U3698 (N_3698,N_2763,N_1090);
nand U3699 (N_3699,N_2024,N_3146);
and U3700 (N_3700,N_2893,N_3113);
nor U3701 (N_3701,N_1563,N_2469);
and U3702 (N_3702,N_3423,N_3200);
nor U3703 (N_3703,N_3390,N_2795);
nand U3704 (N_3704,N_2683,N_1513);
nand U3705 (N_3705,N_3272,N_3172);
or U3706 (N_3706,N_3069,N_2307);
nor U3707 (N_3707,N_2528,N_648);
nand U3708 (N_3708,In_125,N_1306);
xor U3709 (N_3709,N_2121,In_4140);
nand U3710 (N_3710,N_1253,In_1202);
and U3711 (N_3711,N_3443,N_2784);
xnor U3712 (N_3712,In_881,N_2853);
and U3713 (N_3713,N_2970,N_1377);
nand U3714 (N_3714,N_3233,N_2841);
or U3715 (N_3715,N_3320,N_1517);
and U3716 (N_3716,In_2128,In_2568);
nand U3717 (N_3717,N_3456,In_1802);
nand U3718 (N_3718,In_2756,N_2565);
nor U3719 (N_3719,N_3164,N_3009);
and U3720 (N_3720,N_3431,N_2257);
xnor U3721 (N_3721,N_3292,N_3205);
and U3722 (N_3722,N_3028,N_2822);
nor U3723 (N_3723,N_3474,N_1961);
nor U3724 (N_3724,N_3029,N_3271);
nor U3725 (N_3725,N_2629,N_2132);
or U3726 (N_3726,N_2541,In_2261);
and U3727 (N_3727,N_3322,In_1991);
or U3728 (N_3728,N_2731,N_3156);
or U3729 (N_3729,In_4812,In_2305);
and U3730 (N_3730,N_2100,N_225);
or U3731 (N_3731,N_1915,N_3196);
or U3732 (N_3732,N_3434,N_531);
nand U3733 (N_3733,N_3493,In_3616);
or U3734 (N_3734,N_2105,N_3294);
or U3735 (N_3735,In_1271,In_3314);
and U3736 (N_3736,N_3447,N_1719);
or U3737 (N_3737,N_802,N_1638);
or U3738 (N_3738,N_2863,N_3008);
nand U3739 (N_3739,N_3180,N_3076);
and U3740 (N_3740,N_2299,N_1879);
or U3741 (N_3741,N_372,In_4180);
xnor U3742 (N_3742,N_3131,N_2670);
nand U3743 (N_3743,N_3251,N_2805);
nand U3744 (N_3744,In_4873,N_347);
nand U3745 (N_3745,N_2692,In_2105);
or U3746 (N_3746,N_3157,N_2050);
nor U3747 (N_3747,N_2789,N_2871);
and U3748 (N_3748,In_1210,N_3313);
nor U3749 (N_3749,In_4447,N_3319);
and U3750 (N_3750,N_1548,In_3428);
nand U3751 (N_3751,N_2703,N_3203);
nor U3752 (N_3752,N_3105,N_3274);
and U3753 (N_3753,N_2637,In_3468);
nand U3754 (N_3754,N_633,N_2278);
or U3755 (N_3755,In_1467,N_2504);
nor U3756 (N_3756,N_3350,N_3480);
nor U3757 (N_3757,N_3250,N_3479);
and U3758 (N_3758,N_1317,In_469);
or U3759 (N_3759,N_2579,N_2904);
or U3760 (N_3760,N_3349,In_3806);
nand U3761 (N_3761,In_3698,In_1592);
and U3762 (N_3762,N_3486,N_1913);
xor U3763 (N_3763,N_3264,N_3301);
and U3764 (N_3764,In_2784,N_2058);
nor U3765 (N_3765,N_2844,N_2027);
and U3766 (N_3766,N_1803,N_3428);
nand U3767 (N_3767,N_3227,In_3267);
nor U3768 (N_3768,N_2533,In_2629);
and U3769 (N_3769,N_3418,N_2557);
or U3770 (N_3770,N_2713,N_2012);
nand U3771 (N_3771,In_2444,In_347);
nand U3772 (N_3772,N_1270,In_1739);
nand U3773 (N_3773,N_3309,N_3374);
nor U3774 (N_3774,N_2724,N_933);
xor U3775 (N_3775,N_2197,N_1795);
and U3776 (N_3776,In_1998,N_1659);
and U3777 (N_3777,N_3377,In_1521);
nor U3778 (N_3778,N_3388,N_123);
nor U3779 (N_3779,N_1741,N_1786);
or U3780 (N_3780,N_2369,In_1976);
nor U3781 (N_3781,In_1309,N_2113);
and U3782 (N_3782,N_2886,N_3380);
nand U3783 (N_3783,N_2524,N_1600);
nor U3784 (N_3784,In_3242,N_468);
nor U3785 (N_3785,N_2513,N_3235);
nand U3786 (N_3786,N_2865,N_2634);
nand U3787 (N_3787,N_2412,N_3209);
and U3788 (N_3788,In_330,N_2847);
nand U3789 (N_3789,N_3072,N_2082);
and U3790 (N_3790,N_771,N_3145);
nand U3791 (N_3791,N_3016,N_2018);
nand U3792 (N_3792,N_2701,N_2106);
xor U3793 (N_3793,In_235,N_1820);
nand U3794 (N_3794,N_1402,N_3438);
and U3795 (N_3795,N_2219,N_421);
and U3796 (N_3796,N_3451,N_2811);
nand U3797 (N_3797,N_3241,In_3194);
or U3798 (N_3798,N_3077,N_1717);
or U3799 (N_3799,N_3012,N_2495);
or U3800 (N_3800,N_1917,N_856);
xor U3801 (N_3801,N_2873,N_1779);
and U3802 (N_3802,N_1162,N_1296);
nor U3803 (N_3803,N_2852,N_1658);
and U3804 (N_3804,N_3121,N_3259);
nand U3805 (N_3805,N_2571,N_2112);
nand U3806 (N_3806,N_3364,N_3419);
and U3807 (N_3807,N_3245,N_3230);
nand U3808 (N_3808,N_764,In_4448);
nand U3809 (N_3809,N_3269,N_2828);
or U3810 (N_3810,N_3295,In_2943);
nand U3811 (N_3811,In_2583,N_1897);
nand U3812 (N_3812,N_3238,N_2661);
nor U3813 (N_3813,N_2993,N_2231);
and U3814 (N_3814,N_198,In_280);
or U3815 (N_3815,N_3183,N_3347);
or U3816 (N_3816,N_3303,In_2433);
nand U3817 (N_3817,N_1356,N_2832);
or U3818 (N_3818,N_1965,In_4742);
and U3819 (N_3819,N_3222,N_3092);
nand U3820 (N_3820,In_3779,N_3338);
or U3821 (N_3821,N_3351,N_2722);
and U3822 (N_3822,N_2080,N_3469);
and U3823 (N_3823,N_3386,N_3362);
nor U3824 (N_3824,In_2205,N_2810);
or U3825 (N_3825,In_1132,In_900);
nand U3826 (N_3826,N_2145,N_3001);
and U3827 (N_3827,N_3470,N_2387);
or U3828 (N_3828,N_1699,N_3106);
nor U3829 (N_3829,In_4925,N_2605);
nand U3830 (N_3830,In_533,N_1586);
nand U3831 (N_3831,N_345,N_1702);
xnor U3832 (N_3832,N_3155,In_239);
nor U3833 (N_3833,N_3128,N_1321);
xnor U3834 (N_3834,N_3011,N_3006);
nand U3835 (N_3835,N_521,N_165);
or U3836 (N_3836,N_2979,N_689);
nor U3837 (N_3837,N_3232,N_237);
nand U3838 (N_3838,N_3442,N_2464);
and U3839 (N_3839,N_1643,N_2055);
or U3840 (N_3840,N_2576,N_3409);
nand U3841 (N_3841,N_3465,N_1587);
nor U3842 (N_3842,In_346,N_1537);
nand U3843 (N_3843,N_2770,N_3482);
or U3844 (N_3844,N_1331,N_1403);
or U3845 (N_3845,N_2512,In_2726);
nand U3846 (N_3846,N_1833,N_2435);
or U3847 (N_3847,N_3166,In_1465);
and U3848 (N_3848,N_2182,In_3859);
and U3849 (N_3849,N_2685,N_3036);
xor U3850 (N_3850,In_2186,N_2611);
nand U3851 (N_3851,N_3102,N_2268);
xor U3852 (N_3852,N_3321,N_3291);
nand U3853 (N_3853,N_2468,N_2686);
and U3854 (N_3854,N_3118,N_2340);
or U3855 (N_3855,In_275,N_3315);
or U3856 (N_3856,N_1852,N_3169);
nand U3857 (N_3857,N_2408,N_2519);
nor U3858 (N_3858,N_3379,N_108);
nand U3859 (N_3859,N_2654,N_2063);
and U3860 (N_3860,N_2083,N_2511);
nand U3861 (N_3861,N_3317,N_1263);
xnor U3862 (N_3862,N_2017,N_3439);
and U3863 (N_3863,In_3765,In_834);
or U3864 (N_3864,N_3252,N_3187);
nor U3865 (N_3865,In_2643,N_3420);
nor U3866 (N_3866,In_901,N_2645);
or U3867 (N_3867,N_1924,N_359);
xor U3868 (N_3868,N_2941,N_1939);
or U3869 (N_3869,N_3258,N_3088);
nand U3870 (N_3870,N_1243,N_3263);
xor U3871 (N_3871,N_1609,In_2140);
or U3872 (N_3872,N_2578,In_3498);
and U3873 (N_3873,N_327,In_2961);
and U3874 (N_3874,N_3476,N_1618);
nand U3875 (N_3875,In_1701,N_3275);
and U3876 (N_3876,N_2927,N_2748);
nor U3877 (N_3877,N_3285,N_3497);
nand U3878 (N_3878,N_3229,N_3056);
nor U3879 (N_3879,N_3237,N_322);
xor U3880 (N_3880,N_2953,N_3489);
and U3881 (N_3881,In_1647,N_762);
nand U3882 (N_3882,N_2839,In_1505);
or U3883 (N_3883,In_2864,In_374);
and U3884 (N_3884,N_3341,N_3085);
or U3885 (N_3885,In_501,N_3256);
nand U3886 (N_3886,N_577,N_2660);
or U3887 (N_3887,In_1755,N_3071);
or U3888 (N_3888,N_3244,N_3158);
and U3889 (N_3889,In_3111,N_3141);
nor U3890 (N_3890,N_1559,N_2108);
nor U3891 (N_3891,N_3184,N_2812);
nor U3892 (N_3892,N_9,In_2172);
or U3893 (N_3893,N_3450,N_3368);
nand U3894 (N_3894,N_3492,N_2555);
and U3895 (N_3895,N_3403,In_1765);
nand U3896 (N_3896,N_1696,In_4355);
nor U3897 (N_3897,N_2581,N_3070);
and U3898 (N_3898,In_4761,N_2734);
nor U3899 (N_3899,N_2915,N_649);
nor U3900 (N_3900,N_2697,In_4351);
nand U3901 (N_3901,N_3032,N_3335);
and U3902 (N_3902,N_1207,N_3336);
or U3903 (N_3903,N_367,N_2715);
nor U3904 (N_3904,N_2088,N_3361);
xnor U3905 (N_3905,N_2414,N_1282);
or U3906 (N_3906,In_1899,N_2607);
nand U3907 (N_3907,N_1322,N_576);
nor U3908 (N_3908,N_3425,N_911);
xor U3909 (N_3909,In_2614,N_2269);
and U3910 (N_3910,N_1949,N_3013);
nor U3911 (N_3911,N_3464,N_2848);
xor U3912 (N_3912,N_3091,N_3287);
nand U3913 (N_3913,N_3140,In_4430);
and U3914 (N_3914,N_3035,In_3536);
nor U3915 (N_3915,In_4305,N_1902);
nor U3916 (N_3916,N_2356,N_3415);
nand U3917 (N_3917,In_1554,N_2632);
nand U3918 (N_3918,N_3305,N_450);
or U3919 (N_3919,N_2896,N_1841);
and U3920 (N_3920,N_2930,In_161);
or U3921 (N_3921,N_2948,N_1734);
or U3922 (N_3922,N_2718,N_2804);
nand U3923 (N_3923,N_3055,N_2542);
or U3924 (N_3924,N_2983,N_1900);
and U3925 (N_3925,In_1184,In_4577);
nand U3926 (N_3926,N_1099,N_3139);
nand U3927 (N_3927,N_661,N_2667);
and U3928 (N_3928,N_155,N_3297);
nor U3929 (N_3929,In_2015,N_3242);
or U3930 (N_3930,N_3391,In_3853);
nor U3931 (N_3931,In_1200,N_3163);
nand U3932 (N_3932,In_1474,N_3188);
and U3933 (N_3933,N_1774,In_229);
nor U3934 (N_3934,N_3097,N_3394);
nand U3935 (N_3935,N_3165,In_3042);
or U3936 (N_3936,In_56,In_3081);
or U3937 (N_3937,In_82,N_2817);
nor U3938 (N_3938,N_2303,N_2884);
and U3939 (N_3939,N_2792,N_234);
or U3940 (N_3940,In_4317,In_4682);
or U3941 (N_3941,N_2440,N_3061);
or U3942 (N_3942,In_2014,N_3031);
and U3943 (N_3943,In_3764,N_3129);
nor U3944 (N_3944,In_1861,N_3276);
or U3945 (N_3945,N_1560,N_3412);
or U3946 (N_3946,N_3058,N_990);
and U3947 (N_3947,N_3137,In_4571);
nand U3948 (N_3948,In_2214,N_2996);
and U3949 (N_3949,N_1558,N_3135);
or U3950 (N_3950,N_2266,N_3150);
and U3951 (N_3951,N_3173,N_282);
or U3952 (N_3952,N_3120,N_3094);
xnor U3953 (N_3953,N_2323,N_3478);
nand U3954 (N_3954,N_3096,N_3363);
or U3955 (N_3955,In_319,N_2669);
nor U3956 (N_3956,In_3956,In_3874);
and U3957 (N_3957,In_1338,N_2657);
xnor U3958 (N_3958,N_1026,In_2224);
nand U3959 (N_3959,N_1962,N_2004);
nand U3960 (N_3960,N_676,In_3229);
or U3961 (N_3961,N_3346,N_3370);
nor U3962 (N_3962,N_3283,N_1592);
or U3963 (N_3963,N_3127,N_2836);
or U3964 (N_3964,N_3111,In_4870);
or U3965 (N_3965,N_2267,N_3116);
nand U3966 (N_3966,In_87,In_2541);
nand U3967 (N_3967,N_2466,N_3207);
nor U3968 (N_3968,N_2699,In_2432);
nor U3969 (N_3969,N_3086,N_1163);
nand U3970 (N_3970,N_1556,N_3154);
xnor U3971 (N_3971,N_1538,N_3042);
or U3972 (N_3972,N_2700,N_3171);
or U3973 (N_3973,N_3199,In_1487);
and U3974 (N_3974,N_3223,In_4807);
or U3975 (N_3975,In_3923,N_2707);
or U3976 (N_3976,N_1581,N_3481);
and U3977 (N_3977,In_2549,N_2956);
or U3978 (N_3978,In_2403,N_1405);
nand U3979 (N_3979,N_3314,N_2593);
and U3980 (N_3980,N_2592,N_2481);
nor U3981 (N_3981,N_2803,N_2385);
and U3982 (N_3982,N_2813,N_709);
nand U3983 (N_3983,N_3220,N_2487);
nand U3984 (N_3984,In_2823,N_2647);
xnor U3985 (N_3985,N_3206,In_1233);
or U3986 (N_3986,In_715,N_3051);
nand U3987 (N_3987,N_2348,N_1629);
nor U3988 (N_3988,N_2977,N_2452);
nand U3989 (N_3989,In_2264,N_3485);
nor U3990 (N_3990,N_1597,N_783);
xor U3991 (N_3991,N_1205,N_3473);
nor U3992 (N_3992,N_2631,In_1567);
and U3993 (N_3993,N_3358,N_2753);
nor U3994 (N_3994,N_1235,N_3201);
and U3995 (N_3995,N_3181,N_2726);
and U3996 (N_3996,N_2687,N_2898);
nor U3997 (N_3997,N_3454,N_105);
nor U3998 (N_3998,N_3373,N_910);
xnor U3999 (N_3999,N_3316,In_431);
or U4000 (N_4000,N_2981,N_3383);
xnor U4001 (N_4001,N_3684,N_3687);
nor U4002 (N_4002,N_3829,N_2168);
and U4003 (N_4003,N_3830,N_3726);
or U4004 (N_4004,N_2891,N_2688);
nand U4005 (N_4005,N_3657,N_3964);
nor U4006 (N_4006,N_3495,N_1185);
xor U4007 (N_4007,N_1260,N_3805);
xnor U4008 (N_4008,N_3785,N_3611);
nand U4009 (N_4009,N_3449,N_2932);
nand U4010 (N_4010,N_3983,N_2646);
xor U4011 (N_4011,N_1870,N_3701);
or U4012 (N_4012,N_3665,N_3369);
or U4013 (N_4013,N_3897,N_3924);
nor U4014 (N_4014,N_3776,N_3860);
nand U4015 (N_4015,N_3432,N_3588);
nand U4016 (N_4016,N_3532,N_3820);
nand U4017 (N_4017,N_3427,In_3371);
and U4018 (N_4018,N_3554,N_3445);
xnor U4019 (N_4019,N_3893,N_2379);
xor U4020 (N_4020,N_2944,N_3255);
and U4021 (N_4021,N_3610,N_3618);
nor U4022 (N_4022,N_3936,In_4975);
nor U4023 (N_4023,N_3709,N_3832);
or U4024 (N_4024,N_3942,N_3247);
and U4025 (N_4025,N_2404,N_3546);
and U4026 (N_4026,N_2501,N_3605);
xnor U4027 (N_4027,N_2950,N_3650);
nand U4028 (N_4028,N_2787,In_65);
nand U4029 (N_4029,N_3578,N_3867);
and U4030 (N_4030,N_2766,N_3975);
nand U4031 (N_4031,N_2276,N_3045);
and U4032 (N_4032,N_3067,N_3110);
nand U4033 (N_4033,N_1568,N_3859);
nand U4034 (N_4034,N_3943,N_3767);
nor U4035 (N_4035,N_3598,N_3340);
and U4036 (N_4036,N_3977,N_3167);
or U4037 (N_4037,N_3795,N_3552);
nand U4038 (N_4038,N_2538,N_3838);
or U4039 (N_4039,N_3667,N_3542);
xor U4040 (N_4040,N_3865,In_2068);
nand U4041 (N_4041,N_3633,N_1187);
or U4042 (N_4042,N_3822,N_3296);
or U4043 (N_4043,N_2598,N_3475);
and U4044 (N_4044,In_4961,N_3824);
xor U4045 (N_4045,N_3995,N_3544);
nand U4046 (N_4046,N_3898,N_3402);
nand U4047 (N_4047,N_3161,N_3312);
and U4048 (N_4048,N_3536,N_3804);
nor U4049 (N_4049,N_3857,N_3041);
nand U4050 (N_4050,N_3104,N_3591);
and U4051 (N_4051,N_3782,N_3976);
xor U4052 (N_4052,N_3984,N_3880);
xnor U4053 (N_4053,N_3912,N_3054);
xor U4054 (N_4054,N_3945,N_3962);
nand U4055 (N_4055,N_2110,N_1616);
or U4056 (N_4056,N_3920,N_988);
nand U4057 (N_4057,N_561,N_1576);
xor U4058 (N_4058,In_3530,N_3453);
and U4059 (N_4059,N_3039,In_550);
nand U4060 (N_4060,N_2572,N_3604);
and U4061 (N_4061,N_3090,N_3540);
or U4062 (N_4062,N_3240,N_3555);
nor U4063 (N_4063,N_3729,N_1668);
nor U4064 (N_4064,N_3310,N_2433);
xnor U4065 (N_4065,N_3623,In_2256);
nor U4066 (N_4066,N_1907,N_2918);
nand U4067 (N_4067,N_3950,N_3689);
nand U4068 (N_4068,N_3047,N_3325);
xnor U4069 (N_4069,N_3739,N_3873);
or U4070 (N_4070,N_3632,N_1620);
or U4071 (N_4071,N_3990,N_1474);
nor U4072 (N_4072,N_2849,In_1375);
and U4073 (N_4073,N_3763,N_1794);
or U4074 (N_4074,N_3557,N_3864);
xnor U4075 (N_4075,N_3204,In_3496);
nor U4076 (N_4076,N_3955,N_3810);
nor U4077 (N_4077,N_3625,N_3330);
and U4078 (N_4078,N_3927,N_2644);
xor U4079 (N_4079,N_3334,N_3837);
or U4080 (N_4080,N_619,N_3594);
nor U4081 (N_4081,In_4116,N_3680);
and U4082 (N_4082,N_3147,N_3848);
nand U4083 (N_4083,N_3828,N_3376);
or U4084 (N_4084,In_4978,N_3708);
and U4085 (N_4085,N_2990,N_3355);
nand U4086 (N_4086,N_3811,In_969);
nor U4087 (N_4087,N_3064,N_3466);
and U4088 (N_4088,N_3332,N_3537);
nor U4089 (N_4089,N_3603,N_3959);
nor U4090 (N_4090,N_3902,N_2536);
and U4091 (N_4091,N_3986,N_3669);
or U4092 (N_4092,In_1182,N_3891);
nand U4093 (N_4093,In_2099,N_3716);
xnor U4094 (N_4094,N_3749,In_723);
nand U4095 (N_4095,N_3548,N_3149);
nand U4096 (N_4096,N_2910,N_3328);
nor U4097 (N_4097,N_3768,In_3891);
and U4098 (N_4098,N_1527,N_3168);
or U4099 (N_4099,N_3112,N_2913);
or U4100 (N_4100,N_3807,N_2517);
nand U4101 (N_4101,N_3855,N_3808);
and U4102 (N_4102,N_3918,N_3921);
xor U4103 (N_4103,N_3231,N_3721);
nor U4104 (N_4104,N_2235,N_3602);
and U4105 (N_4105,N_1995,N_2529);
nor U4106 (N_4106,N_3890,N_2933);
or U4107 (N_4107,N_3958,N_3946);
xnor U4108 (N_4108,N_3727,N_3649);
nor U4109 (N_4109,N_3699,N_2816);
or U4110 (N_4110,N_3658,N_3919);
xnor U4111 (N_4111,N_91,N_3694);
nand U4112 (N_4112,N_3909,N_3569);
and U4113 (N_4113,N_3590,N_3735);
and U4114 (N_4114,In_3477,N_3883);
nand U4115 (N_4115,N_2946,In_3870);
and U4116 (N_4116,N_2067,N_2567);
nor U4117 (N_4117,N_3801,N_224);
xor U4118 (N_4118,N_3018,N_3062);
and U4119 (N_4119,N_3046,N_3020);
nand U4120 (N_4120,In_3438,N_1354);
nor U4121 (N_4121,N_3392,N_3186);
or U4122 (N_4122,N_3553,N_3515);
or U4123 (N_4123,N_3724,N_1744);
nand U4124 (N_4124,N_3791,N_3956);
and U4125 (N_4125,N_1769,N_3780);
nand U4126 (N_4126,N_3957,N_3908);
or U4127 (N_4127,N_3520,N_2502);
and U4128 (N_4128,N_2709,N_3947);
or U4129 (N_4129,N_3119,N_3993);
nor U4130 (N_4130,N_53,N_3802);
nand U4131 (N_4131,N_3809,N_3690);
nand U4132 (N_4132,N_3884,N_3814);
or U4133 (N_4133,N_1357,N_3886);
and U4134 (N_4134,In_2005,In_2145);
nand U4135 (N_4135,N_3747,N_3799);
and U4136 (N_4136,N_3888,N_3010);
and U4137 (N_4137,N_3707,N_3757);
nor U4138 (N_4138,N_3965,N_3681);
and U4139 (N_4139,N_2201,N_3617);
nor U4140 (N_4140,N_3348,N_2725);
nand U4141 (N_4141,N_3533,N_3925);
and U4142 (N_4142,N_3043,In_1121);
nor U4143 (N_4143,N_3448,N_3960);
or U4144 (N_4144,N_209,N_2294);
or U4145 (N_4145,N_1130,In_3082);
nor U4146 (N_4146,N_3840,In_30);
nand U4147 (N_4147,N_1437,N_3899);
or U4148 (N_4148,N_2975,N_3710);
or U4149 (N_4149,N_2226,N_2449);
and U4150 (N_4150,N_3663,In_2854);
or U4151 (N_4151,In_4834,N_3827);
nand U4152 (N_4152,In_4259,N_3570);
xnor U4153 (N_4153,N_3750,In_4907);
or U4154 (N_4154,N_3133,N_3528);
xnor U4155 (N_4155,N_2594,N_3744);
nand U4156 (N_4156,N_3929,N_3686);
nand U4157 (N_4157,N_3389,N_3691);
nor U4158 (N_4158,N_3879,N_3267);
and U4159 (N_4159,N_2402,N_3027);
and U4160 (N_4160,N_2013,N_3882);
nor U4161 (N_4161,N_3430,N_3794);
or U4162 (N_4162,N_2141,N_3798);
nand U4163 (N_4163,N_3737,N_1814);
or U4164 (N_4164,N_3526,N_3507);
nand U4165 (N_4165,N_3483,N_3697);
and U4166 (N_4166,N_3108,N_2232);
or U4167 (N_4167,In_4587,In_2051);
and U4168 (N_4168,In_192,N_2827);
or U4169 (N_4169,N_1753,In_3444);
and U4170 (N_4170,N_3440,In_4035);
or U4171 (N_4171,N_3597,N_3903);
nor U4172 (N_4172,N_3523,N_3678);
and U4173 (N_4173,N_3892,N_3787);
nand U4174 (N_4174,N_3397,N_3967);
and U4175 (N_4175,N_3500,N_3997);
nand U4176 (N_4176,N_3529,N_3099);
nand U4177 (N_4177,N_1465,N_3939);
or U4178 (N_4178,N_3940,In_2193);
or U4179 (N_4179,N_3211,N_3262);
or U4180 (N_4180,In_1323,In_3595);
and U4181 (N_4181,N_3645,N_3224);
and U4182 (N_4182,N_3784,In_499);
or U4183 (N_4183,N_3103,N_3406);
nor U4184 (N_4184,N_3871,N_2216);
nand U4185 (N_4185,N_3660,N_3151);
or U4186 (N_4186,N_3728,In_1403);
xnor U4187 (N_4187,N_3733,In_806);
nand U4188 (N_4188,N_3659,In_4029);
and U4189 (N_4189,N_3600,N_3299);
nand U4190 (N_4190,N_2761,N_3175);
and U4191 (N_4191,N_3608,N_3589);
nand U4192 (N_4192,N_2136,N_3289);
xnor U4193 (N_4193,N_2638,N_3753);
and U4194 (N_4194,N_3115,N_3280);
nor U4195 (N_4195,N_3561,N_1083);
or U4196 (N_4196,N_1137,N_1462);
nor U4197 (N_4197,N_3601,N_3410);
nand U4198 (N_4198,N_3408,N_3835);
nor U4199 (N_4199,N_2923,N_1664);
nor U4200 (N_4200,N_3661,N_3613);
nand U4201 (N_4201,N_3651,N_3713);
or U4202 (N_4202,N_3836,N_3866);
nand U4203 (N_4203,N_2928,N_1830);
and U4204 (N_4204,In_3576,N_3429);
or U4205 (N_4205,N_3550,N_3644);
and U4206 (N_4206,N_3577,N_3852);
xnor U4207 (N_4207,In_2379,N_3668);
or U4208 (N_4208,In_1999,N_1315);
and U4209 (N_4209,N_3723,N_3278);
nor U4210 (N_4210,N_3741,In_2119);
and U4211 (N_4211,N_3124,N_3516);
xnor U4212 (N_4212,N_3254,N_2507);
nor U4213 (N_4213,N_3246,N_3797);
nor U4214 (N_4214,N_3720,N_3556);
nor U4215 (N_4215,N_3922,N_2938);
or U4216 (N_4216,N_3307,N_3198);
and U4217 (N_4217,N_3869,N_2689);
nor U4218 (N_4218,N_3868,N_3834);
and U4219 (N_4219,N_3781,N_2508);
xor U4220 (N_4220,N_3586,N_3881);
or U4221 (N_4221,In_2850,N_3505);
nor U4222 (N_4222,N_3545,In_4597);
nor U4223 (N_4223,In_755,N_3614);
or U4224 (N_4224,N_3521,N_1170);
nor U4225 (N_4225,N_3911,N_3932);
and U4226 (N_4226,N_3253,N_3398);
xor U4227 (N_4227,N_3653,N_3904);
nand U4228 (N_4228,N_3014,N_3923);
xnor U4229 (N_4229,In_50,N_3582);
nand U4230 (N_4230,N_3504,N_360);
or U4231 (N_4231,In_4635,N_3512);
nand U4232 (N_4232,N_2158,N_3214);
xnor U4233 (N_4233,In_3928,N_97);
and U4234 (N_4234,N_3719,N_3455);
nand U4235 (N_4235,N_3944,N_3282);
nand U4236 (N_4236,N_2846,N_3839);
nor U4237 (N_4237,N_2615,N_3996);
nand U4238 (N_4238,N_3496,N_3740);
nor U4239 (N_4239,N_3326,N_3875);
or U4240 (N_4240,N_3365,N_3522);
and U4241 (N_4241,N_3664,N_3575);
nor U4242 (N_4242,N_3952,N_2674);
and U4243 (N_4243,In_1346,N_3992);
xor U4244 (N_4244,In_986,N_3637);
nand U4245 (N_4245,In_2221,N_3511);
nand U4246 (N_4246,N_3560,N_244);
nand U4247 (N_4247,N_3991,In_4251);
nor U4248 (N_4248,N_3718,N_3833);
nor U4249 (N_4249,In_1849,N_3648);
nor U4250 (N_4250,N_3052,N_2574);
nor U4251 (N_4251,N_2831,N_2128);
nand U4252 (N_4252,N_2721,N_3685);
nor U4253 (N_4253,In_4699,N_3571);
and U4254 (N_4254,N_1635,N_3980);
nand U4255 (N_4255,In_186,N_3844);
or U4256 (N_4256,In_4793,N_3049);
and U4257 (N_4257,N_2600,N_3619);
nand U4258 (N_4258,N_2208,N_3329);
nor U4259 (N_4259,N_3765,N_3583);
nor U4260 (N_4260,N_3973,N_2620);
nand U4261 (N_4261,In_2730,N_3563);
or U4262 (N_4262,N_3573,N_3444);
or U4263 (N_4263,In_2183,N_2005);
nor U4264 (N_4264,N_3700,N_2319);
nand U4265 (N_4265,N_2659,N_3702);
nand U4266 (N_4266,In_3865,In_1178);
or U4267 (N_4267,N_3974,N_3851);
or U4268 (N_4268,N_2691,N_3579);
or U4269 (N_4269,N_3654,N_3527);
nor U4270 (N_4270,N_3541,N_3764);
or U4271 (N_4271,N_1291,N_3395);
and U4272 (N_4272,N_3862,N_1706);
and U4273 (N_4273,N_3426,In_1607);
xor U4274 (N_4274,N_3635,In_3104);
or U4275 (N_4275,N_1121,N_3717);
or U4276 (N_4276,N_3655,N_3854);
and U4277 (N_4277,N_3761,N_3978);
and U4278 (N_4278,N_3656,N_1655);
nor U4279 (N_4279,In_3489,In_3850);
nor U4280 (N_4280,In_1258,N_3308);
or U4281 (N_4281,N_2935,N_1342);
or U4282 (N_4282,N_3107,N_1632);
nand U4283 (N_4283,N_3825,N_3677);
xnor U4284 (N_4284,N_3777,N_3652);
or U4285 (N_4285,In_3718,In_2547);
and U4286 (N_4286,N_3926,N_2706);
or U4287 (N_4287,N_2098,In_4157);
nand U4288 (N_4288,N_2908,N_3306);
nand U4289 (N_4289,N_2796,N_3751);
and U4290 (N_4290,N_3281,N_3405);
nor U4291 (N_4291,N_1827,N_3969);
or U4292 (N_4292,In_3575,N_2335);
and U4293 (N_4293,N_2759,N_3812);
nor U4294 (N_4294,N_2856,N_570);
and U4295 (N_4295,N_3773,N_3647);
xor U4296 (N_4296,N_1082,N_3574);
or U4297 (N_4297,N_3863,N_693);
nor U4298 (N_4298,N_3622,N_3770);
and U4299 (N_4299,N_3411,N_3671);
and U4300 (N_4300,N_3954,N_3774);
nor U4301 (N_4301,N_3503,N_3615);
nor U4302 (N_4302,N_3510,N_3621);
nor U4303 (N_4303,In_4257,N_3966);
nor U4304 (N_4304,N_3683,In_2076);
nor U4305 (N_4305,N_3585,N_3581);
nor U4306 (N_4306,N_730,N_3606);
nor U4307 (N_4307,N_3565,N_3748);
or U4308 (N_4308,N_1772,N_2649);
or U4309 (N_4309,N_3771,N_3817);
nor U4310 (N_4310,N_3738,N_3901);
or U4311 (N_4311,N_3698,N_1022);
nor U4312 (N_4312,N_3937,N_3023);
xor U4313 (N_4313,N_513,N_3760);
or U4314 (N_4314,N_3083,N_922);
nand U4315 (N_4315,N_3323,N_2366);
nand U4316 (N_4316,N_3792,N_3519);
nor U4317 (N_4317,N_240,N_3612);
or U4318 (N_4318,N_2794,N_3123);
or U4319 (N_4319,N_3421,N_1542);
and U4320 (N_4320,N_3907,N_3337);
nor U4321 (N_4321,N_1589,In_2558);
xor U4322 (N_4322,N_323,N_3742);
nand U4323 (N_4323,N_474,In_3738);
nor U4324 (N_4324,N_3640,In_3189);
nand U4325 (N_4325,N_3098,In_578);
or U4326 (N_4326,N_1262,N_3217);
xnor U4327 (N_4327,N_653,N_3693);
or U4328 (N_4328,N_2346,N_3895);
xnor U4329 (N_4329,N_3968,N_3914);
nor U4330 (N_4330,N_3122,N_3706);
nand U4331 (N_4331,N_3535,N_1122);
xnor U4332 (N_4332,In_359,N_3916);
nor U4333 (N_4333,N_3352,N_3981);
and U4334 (N_4334,N_3236,N_3134);
nand U4335 (N_4335,N_3371,N_3642);
nand U4336 (N_4336,N_3075,N_3772);
or U4337 (N_4337,N_3087,In_2462);
and U4338 (N_4338,N_3144,N_3756);
or U4339 (N_4339,N_2806,N_3786);
and U4340 (N_4340,N_3714,N_923);
or U4341 (N_4341,N_3210,N_3459);
or U4342 (N_4342,N_3228,In_3049);
nand U4343 (N_4343,N_2040,N_2962);
and U4344 (N_4344,N_3413,N_3896);
nor U4345 (N_4345,N_3775,N_2377);
nor U4346 (N_4346,N_3213,N_328);
nor U4347 (N_4347,N_3704,N_1358);
nand U4348 (N_4348,N_3549,N_3160);
nand U4349 (N_4349,N_3587,N_3595);
xnor U4350 (N_4350,N_3872,N_3736);
nand U4351 (N_4351,N_1332,N_3462);
nor U4352 (N_4352,N_3858,N_3643);
xnor U4353 (N_4353,N_3620,N_3998);
nand U4354 (N_4354,N_3856,N_3796);
nand U4355 (N_4355,N_876,In_576);
nand U4356 (N_4356,N_2251,N_2116);
and U4357 (N_4357,N_3999,In_317);
or U4358 (N_4358,N_3531,N_1217);
or U4359 (N_4359,N_606,N_3831);
nor U4360 (N_4360,N_3745,N_3580);
or U4361 (N_4361,N_3778,N_3711);
and U4362 (N_4362,N_3003,N_3963);
and U4363 (N_4363,N_3906,N_3193);
or U4364 (N_4364,N_1398,N_3813);
or U4365 (N_4365,N_3938,N_3971);
and U4366 (N_4366,In_188,N_3987);
nand U4367 (N_4367,N_3951,N_3675);
and U4368 (N_4368,N_3501,N_3979);
and U4369 (N_4369,N_1168,N_3688);
xor U4370 (N_4370,N_3517,N_3731);
or U4371 (N_4371,N_3818,N_3845);
nor U4372 (N_4372,N_3988,N_2800);
or U4373 (N_4373,N_3592,N_3518);
nor U4374 (N_4374,N_3562,N_3679);
nand U4375 (N_4375,N_3551,N_3638);
nor U4376 (N_4376,N_3695,In_3312);
nor U4377 (N_4377,N_3961,N_3841);
nor U4378 (N_4378,In_299,N_3078);
or U4379 (N_4379,N_3630,N_3970);
or U4380 (N_4380,N_3877,N_3752);
or U4381 (N_4381,N_3788,In_3274);
nor U4382 (N_4382,N_3170,N_3949);
xor U4383 (N_4383,N_3743,N_3887);
nor U4384 (N_4384,N_3626,N_3754);
or U4385 (N_4385,N_2562,N_3823);
or U4386 (N_4386,N_3734,N_2500);
or U4387 (N_4387,N_3367,N_3628);
or U4388 (N_4388,N_3017,N_3599);
nor U4389 (N_4389,In_2390,N_3226);
nor U4390 (N_4390,N_2640,N_3539);
nor U4391 (N_4391,N_3803,N_3682);
and U4392 (N_4392,N_2189,N_3850);
nor U4393 (N_4393,N_3715,N_2868);
and U4394 (N_4394,N_2867,N_1061);
and U4395 (N_4395,N_3766,N_1136);
and U4396 (N_4396,N_3513,N_3558);
nand U4397 (N_4397,N_3174,N_2070);
nor U4398 (N_4398,N_2325,N_3874);
and U4399 (N_4399,N_3616,N_3568);
or U4400 (N_4400,N_3900,N_3985);
nor U4401 (N_4401,N_2330,N_1074);
or U4402 (N_4402,In_1001,N_3639);
nand U4403 (N_4403,N_3530,N_3972);
or U4404 (N_4404,N_3399,In_1026);
nor U4405 (N_4405,N_3050,In_2406);
nand U4406 (N_4406,N_3769,N_2742);
nor U4407 (N_4407,N_3755,N_3524);
nand U4408 (N_4408,N_3356,N_3631);
nand U4409 (N_4409,N_3759,N_3889);
or U4410 (N_4410,N_3082,N_3382);
nand U4411 (N_4411,In_3603,N_3624);
or U4412 (N_4412,N_1478,N_3509);
nand U4413 (N_4413,N_3636,N_3878);
or U4414 (N_4414,N_596,In_2325);
nor U4415 (N_4415,N_2762,N_1447);
or U4416 (N_4416,N_3270,N_3815);
and U4417 (N_4417,N_3826,N_3234);
nand U4418 (N_4418,N_3068,N_3861);
xnor U4419 (N_4419,N_3609,N_3002);
or U4420 (N_4420,N_3779,N_3417);
or U4421 (N_4421,In_2467,In_1961);
nand U4422 (N_4422,N_1141,N_2489);
and U4423 (N_4423,N_3596,N_3670);
and U4424 (N_4424,N_3342,N_3928);
nor U4425 (N_4425,N_3843,N_1041);
and U4426 (N_4426,N_3414,N_3260);
or U4427 (N_4427,N_3870,N_2381);
nor U4428 (N_4428,N_3725,N_3722);
or U4429 (N_4429,N_3933,In_801);
xnor U4430 (N_4430,N_2111,N_3989);
and U4431 (N_4431,N_2305,N_3477);
or U4432 (N_4432,N_3853,N_1996);
nor U4433 (N_4433,N_3646,N_2460);
and U4434 (N_4434,N_3696,N_3525);
nand U4435 (N_4435,N_3905,N_3806);
and U4436 (N_4436,N_3584,N_769);
or U4437 (N_4437,N_3607,N_3666);
nand U4438 (N_4438,N_71,N_3534);
or U4439 (N_4439,N_3793,N_2872);
or U4440 (N_4440,N_3641,N_3538);
nand U4441 (N_4441,N_2681,N_1988);
xor U4442 (N_4442,N_3931,N_1761);
and U4443 (N_4443,N_3000,N_3953);
and U4444 (N_4444,N_2582,N_3502);
nor U4445 (N_4445,N_3543,N_3053);
and U4446 (N_4446,N_2964,In_364);
nand U4447 (N_4447,In_3335,N_2549);
and U4448 (N_4448,N_3508,N_3662);
and U4449 (N_4449,N_3564,N_1228);
or U4450 (N_4450,In_3829,N_3179);
nand U4451 (N_4451,N_3849,In_2821);
or U4452 (N_4452,N_3634,N_3143);
or U4453 (N_4453,N_3441,N_3758);
and U4454 (N_4454,N_2666,N_2095);
and U4455 (N_4455,In_3713,N_3790);
nand U4456 (N_4456,N_3692,N_3816);
nor U4457 (N_4457,N_3800,N_3917);
nor U4458 (N_4458,N_1545,N_1333);
nand U4459 (N_4459,N_3847,N_3732);
or U4460 (N_4460,In_3751,N_3913);
or U4461 (N_4461,N_3762,N_3300);
nand U4462 (N_4462,N_3066,N_3057);
or U4463 (N_4463,N_3712,N_3934);
nor U4464 (N_4464,N_3339,N_2658);
nor U4465 (N_4465,N_3506,N_3672);
or U4466 (N_4466,N_3219,N_1685);
nor U4467 (N_4467,N_3994,N_3060);
nand U4468 (N_4468,N_3842,N_3948);
nor U4469 (N_4469,N_3034,N_3494);
xnor U4470 (N_4470,N_2238,N_3876);
nand U4471 (N_4471,N_3915,N_3783);
and U4472 (N_4472,N_3819,N_3941);
nand U4473 (N_4473,N_3572,N_3703);
and U4474 (N_4474,N_2845,N_3627);
or U4475 (N_4475,N_3100,N_3559);
nor U4476 (N_4476,N_3142,N_3629);
nand U4477 (N_4477,N_3547,N_3846);
xor U4478 (N_4478,N_3593,N_3566);
nand U4479 (N_4479,N_3676,N_1663);
and U4480 (N_4480,N_3022,N_1512);
and U4481 (N_4481,N_1032,N_3114);
or U4482 (N_4482,N_3208,N_3821);
nor U4483 (N_4483,N_3730,N_3982);
nand U4484 (N_4484,N_3746,In_811);
nand U4485 (N_4485,In_1708,N_3673);
or U4486 (N_4486,N_3487,N_2777);
nand U4487 (N_4487,N_3674,In_3259);
and U4488 (N_4488,N_3705,N_2980);
nand U4489 (N_4489,N_1208,N_2486);
or U4490 (N_4490,In_3997,N_3576);
nand U4491 (N_4491,N_3935,In_4833);
nand U4492 (N_4492,N_3197,N_3357);
nor U4493 (N_4493,N_3567,N_3885);
nor U4494 (N_4494,N_3514,N_2470);
and U4495 (N_4495,N_3894,N_3789);
and U4496 (N_4496,N_1239,In_480);
nand U4497 (N_4497,N_2986,N_3910);
or U4498 (N_4498,N_3498,N_3400);
nand U4499 (N_4499,N_3930,N_3005);
or U4500 (N_4500,N_4268,N_4234);
xnor U4501 (N_4501,N_4044,N_4046);
xor U4502 (N_4502,N_4127,N_4397);
nor U4503 (N_4503,N_4100,N_4342);
or U4504 (N_4504,N_4084,N_4463);
and U4505 (N_4505,N_4261,N_4144);
or U4506 (N_4506,N_4070,N_4211);
and U4507 (N_4507,N_4034,N_4159);
nand U4508 (N_4508,N_4078,N_4407);
or U4509 (N_4509,N_4200,N_4208);
and U4510 (N_4510,N_4202,N_4298);
nand U4511 (N_4511,N_4102,N_4314);
xnor U4512 (N_4512,N_4014,N_4187);
nand U4513 (N_4513,N_4056,N_4170);
nand U4514 (N_4514,N_4233,N_4137);
or U4515 (N_4515,N_4467,N_4009);
or U4516 (N_4516,N_4385,N_4461);
xor U4517 (N_4517,N_4262,N_4321);
and U4518 (N_4518,N_4072,N_4418);
nand U4519 (N_4519,N_4090,N_4382);
and U4520 (N_4520,N_4344,N_4332);
and U4521 (N_4521,N_4057,N_4316);
or U4522 (N_4522,N_4391,N_4053);
and U4523 (N_4523,N_4259,N_4171);
or U4524 (N_4524,N_4381,N_4319);
or U4525 (N_4525,N_4177,N_4188);
and U4526 (N_4526,N_4452,N_4213);
or U4527 (N_4527,N_4021,N_4293);
nor U4528 (N_4528,N_4371,N_4436);
or U4529 (N_4529,N_4284,N_4026);
nand U4530 (N_4530,N_4096,N_4449);
nor U4531 (N_4531,N_4160,N_4274);
or U4532 (N_4532,N_4176,N_4460);
and U4533 (N_4533,N_4236,N_4041);
nor U4534 (N_4534,N_4282,N_4412);
and U4535 (N_4535,N_4334,N_4326);
nand U4536 (N_4536,N_4083,N_4087);
or U4537 (N_4537,N_4290,N_4360);
nand U4538 (N_4538,N_4434,N_4349);
nand U4539 (N_4539,N_4311,N_4424);
and U4540 (N_4540,N_4351,N_4099);
and U4541 (N_4541,N_4441,N_4199);
nand U4542 (N_4542,N_4266,N_4367);
nand U4543 (N_4543,N_4362,N_4337);
and U4544 (N_4544,N_4347,N_4495);
nand U4545 (N_4545,N_4086,N_4092);
or U4546 (N_4546,N_4076,N_4069);
nor U4547 (N_4547,N_4228,N_4359);
nand U4548 (N_4548,N_4483,N_4297);
nand U4549 (N_4549,N_4364,N_4440);
nand U4550 (N_4550,N_4417,N_4478);
and U4551 (N_4551,N_4263,N_4265);
nand U4552 (N_4552,N_4062,N_4198);
nor U4553 (N_4553,N_4308,N_4378);
nor U4554 (N_4554,N_4398,N_4329);
and U4555 (N_4555,N_4167,N_4355);
nor U4556 (N_4556,N_4366,N_4112);
nand U4557 (N_4557,N_4264,N_4317);
or U4558 (N_4558,N_4027,N_4130);
nand U4559 (N_4559,N_4439,N_4286);
or U4560 (N_4560,N_4250,N_4303);
nand U4561 (N_4561,N_4377,N_4001);
and U4562 (N_4562,N_4346,N_4458);
and U4563 (N_4563,N_4050,N_4134);
and U4564 (N_4564,N_4003,N_4142);
nor U4565 (N_4565,N_4283,N_4153);
nand U4566 (N_4566,N_4012,N_4331);
nand U4567 (N_4567,N_4114,N_4037);
xnor U4568 (N_4568,N_4244,N_4361);
or U4569 (N_4569,N_4287,N_4481);
and U4570 (N_4570,N_4085,N_4411);
and U4571 (N_4571,N_4428,N_4493);
nand U4572 (N_4572,N_4150,N_4402);
nand U4573 (N_4573,N_4182,N_4444);
nor U4574 (N_4574,N_4479,N_4138);
nand U4575 (N_4575,N_4291,N_4248);
xnor U4576 (N_4576,N_4074,N_4232);
or U4577 (N_4577,N_4107,N_4272);
nand U4578 (N_4578,N_4082,N_4011);
nand U4579 (N_4579,N_4241,N_4466);
and U4580 (N_4580,N_4431,N_4443);
nor U4581 (N_4581,N_4005,N_4141);
nand U4582 (N_4582,N_4052,N_4343);
or U4583 (N_4583,N_4222,N_4183);
nand U4584 (N_4584,N_4327,N_4075);
nor U4585 (N_4585,N_4437,N_4051);
or U4586 (N_4586,N_4013,N_4108);
nor U4587 (N_4587,N_4235,N_4128);
nand U4588 (N_4588,N_4492,N_4476);
or U4589 (N_4589,N_4019,N_4470);
nor U4590 (N_4590,N_4038,N_4065);
nor U4591 (N_4591,N_4219,N_4393);
xnor U4592 (N_4592,N_4471,N_4406);
xnor U4593 (N_4593,N_4116,N_4191);
nand U4594 (N_4594,N_4031,N_4455);
nor U4595 (N_4595,N_4295,N_4457);
xnor U4596 (N_4596,N_4077,N_4194);
and U4597 (N_4597,N_4210,N_4110);
xor U4598 (N_4598,N_4140,N_4474);
or U4599 (N_4599,N_4469,N_4067);
nand U4600 (N_4600,N_4043,N_4464);
nand U4601 (N_4601,N_4215,N_4193);
nor U4602 (N_4602,N_4473,N_4433);
or U4603 (N_4603,N_4126,N_4275);
or U4604 (N_4604,N_4358,N_4118);
nor U4605 (N_4605,N_4029,N_4098);
xor U4606 (N_4606,N_4223,N_4459);
or U4607 (N_4607,N_4256,N_4498);
or U4608 (N_4608,N_4305,N_4320);
and U4609 (N_4609,N_4273,N_4489);
or U4610 (N_4610,N_4093,N_4022);
or U4611 (N_4611,N_4094,N_4073);
or U4612 (N_4612,N_4363,N_4106);
nor U4613 (N_4613,N_4354,N_4136);
or U4614 (N_4614,N_4373,N_4312);
or U4615 (N_4615,N_4288,N_4310);
or U4616 (N_4616,N_4294,N_4227);
xnor U4617 (N_4617,N_4400,N_4081);
xor U4618 (N_4618,N_4416,N_4447);
nor U4619 (N_4619,N_4174,N_4451);
xor U4620 (N_4620,N_4068,N_4122);
nand U4621 (N_4621,N_4404,N_4119);
nand U4622 (N_4622,N_4220,N_4230);
and U4623 (N_4623,N_4484,N_4237);
nand U4624 (N_4624,N_4209,N_4190);
nor U4625 (N_4625,N_4135,N_4401);
xnor U4626 (N_4626,N_4023,N_4318);
or U4627 (N_4627,N_4386,N_4482);
xor U4628 (N_4628,N_4179,N_4004);
or U4629 (N_4629,N_4278,N_4335);
or U4630 (N_4630,N_4323,N_4207);
nor U4631 (N_4631,N_4429,N_4338);
nand U4632 (N_4632,N_4375,N_4405);
and U4633 (N_4633,N_4025,N_4060);
nor U4634 (N_4634,N_4020,N_4379);
xor U4635 (N_4635,N_4267,N_4131);
nand U4636 (N_4636,N_4205,N_4413);
and U4637 (N_4637,N_4339,N_4061);
nand U4638 (N_4638,N_4221,N_4423);
nand U4639 (N_4639,N_4462,N_4139);
nor U4640 (N_4640,N_4269,N_4178);
nand U4641 (N_4641,N_4480,N_4330);
xnor U4642 (N_4642,N_4164,N_4113);
and U4643 (N_4643,N_4324,N_4356);
or U4644 (N_4644,N_4152,N_4111);
xor U4645 (N_4645,N_4255,N_4292);
nor U4646 (N_4646,N_4350,N_4496);
nand U4647 (N_4647,N_4105,N_4180);
nand U4648 (N_4648,N_4477,N_4097);
nor U4649 (N_4649,N_4218,N_4030);
xor U4650 (N_4650,N_4487,N_4066);
or U4651 (N_4651,N_4499,N_4438);
nor U4652 (N_4652,N_4166,N_4442);
and U4653 (N_4653,N_4225,N_4403);
nor U4654 (N_4654,N_4206,N_4195);
nand U4655 (N_4655,N_4184,N_4432);
or U4656 (N_4656,N_4063,N_4032);
nor U4657 (N_4657,N_4071,N_4054);
nand U4658 (N_4658,N_4485,N_4216);
or U4659 (N_4659,N_4425,N_4427);
nand U4660 (N_4660,N_4392,N_4079);
and U4661 (N_4661,N_4189,N_4380);
nor U4662 (N_4662,N_4059,N_4388);
nor U4663 (N_4663,N_4133,N_4247);
xor U4664 (N_4664,N_4280,N_4456);
or U4665 (N_4665,N_4162,N_4124);
and U4666 (N_4666,N_4175,N_4115);
and U4667 (N_4667,N_4145,N_4204);
and U4668 (N_4668,N_4390,N_4396);
and U4669 (N_4669,N_4475,N_4486);
nand U4670 (N_4670,N_4309,N_4465);
nor U4671 (N_4671,N_4374,N_4018);
nand U4672 (N_4672,N_4217,N_4251);
nor U4673 (N_4673,N_4448,N_4289);
nor U4674 (N_4674,N_4008,N_4148);
nor U4675 (N_4675,N_4299,N_4033);
nand U4676 (N_4676,N_4414,N_4049);
and U4677 (N_4677,N_4016,N_4491);
and U4678 (N_4678,N_4196,N_4254);
or U4679 (N_4679,N_4226,N_4168);
nor U4680 (N_4680,N_4121,N_4095);
or U4681 (N_4681,N_4010,N_4408);
and U4682 (N_4682,N_4315,N_4157);
or U4683 (N_4683,N_4389,N_4253);
and U4684 (N_4684,N_4281,N_4224);
and U4685 (N_4685,N_4242,N_4333);
xnor U4686 (N_4686,N_4245,N_4123);
or U4687 (N_4687,N_4002,N_4120);
and U4688 (N_4688,N_4306,N_4277);
xnor U4689 (N_4689,N_4048,N_4246);
nand U4690 (N_4690,N_4240,N_4322);
or U4691 (N_4691,N_4426,N_4101);
or U4692 (N_4692,N_4352,N_4125);
or U4693 (N_4693,N_4169,N_4421);
nand U4694 (N_4694,N_4357,N_4007);
nor U4695 (N_4695,N_4345,N_4192);
and U4696 (N_4696,N_4201,N_4185);
and U4697 (N_4697,N_4036,N_4369);
nand U4698 (N_4698,N_4422,N_4304);
nor U4699 (N_4699,N_4300,N_4419);
or U4700 (N_4700,N_4387,N_4472);
and U4701 (N_4701,N_4155,N_4383);
nand U4702 (N_4702,N_4158,N_4197);
nand U4703 (N_4703,N_4340,N_4181);
or U4704 (N_4704,N_4173,N_4257);
nand U4705 (N_4705,N_4271,N_4146);
nand U4706 (N_4706,N_4231,N_4129);
xnor U4707 (N_4707,N_4494,N_4258);
nor U4708 (N_4708,N_4450,N_4276);
or U4709 (N_4709,N_4446,N_4058);
or U4710 (N_4710,N_4229,N_4104);
and U4711 (N_4711,N_4328,N_4420);
nand U4712 (N_4712,N_4395,N_4488);
nand U4713 (N_4713,N_4239,N_4147);
nand U4714 (N_4714,N_4017,N_4410);
or U4715 (N_4715,N_4279,N_4040);
or U4716 (N_4716,N_4028,N_4117);
and U4717 (N_4717,N_4302,N_4435);
or U4718 (N_4718,N_4006,N_4325);
nand U4719 (N_4719,N_4430,N_4154);
or U4720 (N_4720,N_4238,N_4270);
or U4721 (N_4721,N_4109,N_4348);
nand U4722 (N_4722,N_4336,N_4370);
nand U4723 (N_4723,N_4445,N_4409);
nor U4724 (N_4724,N_4353,N_4260);
xnor U4725 (N_4725,N_4394,N_4064);
and U4726 (N_4726,N_4368,N_4089);
nor U4727 (N_4727,N_4468,N_4163);
nand U4728 (N_4728,N_4103,N_4497);
nand U4729 (N_4729,N_4055,N_4047);
or U4730 (N_4730,N_4203,N_4214);
nor U4731 (N_4731,N_4415,N_4042);
or U4732 (N_4732,N_4399,N_4285);
and U4733 (N_4733,N_4132,N_4384);
or U4734 (N_4734,N_4156,N_4000);
or U4735 (N_4735,N_4372,N_4149);
or U4736 (N_4736,N_4454,N_4165);
nor U4737 (N_4737,N_4151,N_4252);
or U4738 (N_4738,N_4045,N_4143);
and U4739 (N_4739,N_4365,N_4172);
nor U4740 (N_4740,N_4341,N_4212);
or U4741 (N_4741,N_4249,N_4015);
and U4742 (N_4742,N_4307,N_4313);
xnor U4743 (N_4743,N_4088,N_4091);
and U4744 (N_4744,N_4039,N_4301);
nand U4745 (N_4745,N_4186,N_4161);
or U4746 (N_4746,N_4035,N_4024);
nand U4747 (N_4747,N_4490,N_4453);
nand U4748 (N_4748,N_4243,N_4296);
or U4749 (N_4749,N_4376,N_4080);
or U4750 (N_4750,N_4015,N_4260);
nand U4751 (N_4751,N_4372,N_4319);
nand U4752 (N_4752,N_4429,N_4141);
nor U4753 (N_4753,N_4024,N_4007);
and U4754 (N_4754,N_4051,N_4404);
xor U4755 (N_4755,N_4338,N_4346);
nand U4756 (N_4756,N_4352,N_4023);
nand U4757 (N_4757,N_4382,N_4123);
nand U4758 (N_4758,N_4245,N_4135);
or U4759 (N_4759,N_4062,N_4470);
nor U4760 (N_4760,N_4365,N_4371);
nand U4761 (N_4761,N_4022,N_4492);
or U4762 (N_4762,N_4263,N_4382);
and U4763 (N_4763,N_4424,N_4431);
nor U4764 (N_4764,N_4181,N_4407);
nor U4765 (N_4765,N_4131,N_4193);
nor U4766 (N_4766,N_4081,N_4017);
nand U4767 (N_4767,N_4337,N_4026);
nor U4768 (N_4768,N_4058,N_4366);
xnor U4769 (N_4769,N_4056,N_4103);
and U4770 (N_4770,N_4497,N_4137);
nor U4771 (N_4771,N_4060,N_4159);
or U4772 (N_4772,N_4471,N_4370);
or U4773 (N_4773,N_4189,N_4238);
nand U4774 (N_4774,N_4152,N_4107);
or U4775 (N_4775,N_4149,N_4109);
or U4776 (N_4776,N_4240,N_4454);
and U4777 (N_4777,N_4170,N_4007);
nor U4778 (N_4778,N_4133,N_4207);
or U4779 (N_4779,N_4035,N_4369);
nor U4780 (N_4780,N_4409,N_4126);
or U4781 (N_4781,N_4468,N_4287);
xnor U4782 (N_4782,N_4407,N_4094);
and U4783 (N_4783,N_4415,N_4189);
xnor U4784 (N_4784,N_4162,N_4335);
nand U4785 (N_4785,N_4277,N_4034);
or U4786 (N_4786,N_4221,N_4236);
nand U4787 (N_4787,N_4336,N_4430);
nor U4788 (N_4788,N_4143,N_4193);
nand U4789 (N_4789,N_4400,N_4249);
nand U4790 (N_4790,N_4053,N_4208);
and U4791 (N_4791,N_4051,N_4120);
nand U4792 (N_4792,N_4172,N_4385);
nand U4793 (N_4793,N_4389,N_4069);
nand U4794 (N_4794,N_4038,N_4481);
nor U4795 (N_4795,N_4045,N_4327);
nand U4796 (N_4796,N_4265,N_4162);
and U4797 (N_4797,N_4139,N_4089);
nand U4798 (N_4798,N_4204,N_4152);
nor U4799 (N_4799,N_4177,N_4047);
nor U4800 (N_4800,N_4378,N_4497);
xnor U4801 (N_4801,N_4089,N_4187);
nor U4802 (N_4802,N_4383,N_4294);
and U4803 (N_4803,N_4350,N_4328);
and U4804 (N_4804,N_4028,N_4162);
or U4805 (N_4805,N_4378,N_4233);
or U4806 (N_4806,N_4213,N_4210);
nand U4807 (N_4807,N_4488,N_4429);
nor U4808 (N_4808,N_4370,N_4358);
and U4809 (N_4809,N_4241,N_4059);
xor U4810 (N_4810,N_4012,N_4234);
or U4811 (N_4811,N_4417,N_4383);
or U4812 (N_4812,N_4117,N_4489);
nand U4813 (N_4813,N_4387,N_4206);
and U4814 (N_4814,N_4211,N_4144);
nor U4815 (N_4815,N_4325,N_4086);
nand U4816 (N_4816,N_4131,N_4012);
and U4817 (N_4817,N_4314,N_4390);
nor U4818 (N_4818,N_4470,N_4310);
nor U4819 (N_4819,N_4087,N_4018);
and U4820 (N_4820,N_4381,N_4273);
or U4821 (N_4821,N_4225,N_4247);
or U4822 (N_4822,N_4382,N_4238);
xor U4823 (N_4823,N_4149,N_4205);
or U4824 (N_4824,N_4179,N_4295);
nor U4825 (N_4825,N_4237,N_4244);
nand U4826 (N_4826,N_4245,N_4419);
and U4827 (N_4827,N_4042,N_4487);
or U4828 (N_4828,N_4062,N_4094);
or U4829 (N_4829,N_4169,N_4085);
nand U4830 (N_4830,N_4462,N_4070);
nor U4831 (N_4831,N_4452,N_4313);
nor U4832 (N_4832,N_4290,N_4224);
nor U4833 (N_4833,N_4364,N_4026);
nand U4834 (N_4834,N_4133,N_4340);
or U4835 (N_4835,N_4297,N_4107);
xor U4836 (N_4836,N_4386,N_4272);
xor U4837 (N_4837,N_4178,N_4232);
or U4838 (N_4838,N_4276,N_4492);
and U4839 (N_4839,N_4376,N_4290);
nor U4840 (N_4840,N_4091,N_4185);
xnor U4841 (N_4841,N_4425,N_4331);
and U4842 (N_4842,N_4019,N_4409);
nor U4843 (N_4843,N_4051,N_4107);
nand U4844 (N_4844,N_4001,N_4383);
nor U4845 (N_4845,N_4005,N_4459);
nor U4846 (N_4846,N_4354,N_4405);
nor U4847 (N_4847,N_4455,N_4437);
and U4848 (N_4848,N_4230,N_4010);
and U4849 (N_4849,N_4335,N_4317);
nand U4850 (N_4850,N_4429,N_4380);
nand U4851 (N_4851,N_4011,N_4287);
and U4852 (N_4852,N_4140,N_4287);
nor U4853 (N_4853,N_4322,N_4038);
nand U4854 (N_4854,N_4066,N_4364);
nand U4855 (N_4855,N_4243,N_4414);
nand U4856 (N_4856,N_4405,N_4295);
and U4857 (N_4857,N_4346,N_4473);
or U4858 (N_4858,N_4358,N_4265);
xor U4859 (N_4859,N_4270,N_4275);
nand U4860 (N_4860,N_4051,N_4230);
nor U4861 (N_4861,N_4137,N_4204);
and U4862 (N_4862,N_4124,N_4345);
or U4863 (N_4863,N_4464,N_4135);
nand U4864 (N_4864,N_4012,N_4226);
or U4865 (N_4865,N_4408,N_4181);
and U4866 (N_4866,N_4319,N_4382);
and U4867 (N_4867,N_4493,N_4471);
nor U4868 (N_4868,N_4217,N_4361);
xor U4869 (N_4869,N_4319,N_4406);
and U4870 (N_4870,N_4194,N_4113);
nand U4871 (N_4871,N_4244,N_4315);
and U4872 (N_4872,N_4439,N_4125);
nand U4873 (N_4873,N_4146,N_4212);
or U4874 (N_4874,N_4152,N_4390);
and U4875 (N_4875,N_4303,N_4006);
and U4876 (N_4876,N_4089,N_4444);
and U4877 (N_4877,N_4410,N_4465);
nor U4878 (N_4878,N_4389,N_4209);
or U4879 (N_4879,N_4485,N_4271);
or U4880 (N_4880,N_4394,N_4322);
nor U4881 (N_4881,N_4253,N_4118);
nor U4882 (N_4882,N_4176,N_4259);
nor U4883 (N_4883,N_4073,N_4103);
nand U4884 (N_4884,N_4137,N_4251);
nand U4885 (N_4885,N_4251,N_4065);
nor U4886 (N_4886,N_4117,N_4276);
nor U4887 (N_4887,N_4458,N_4370);
nor U4888 (N_4888,N_4186,N_4267);
nand U4889 (N_4889,N_4178,N_4008);
xnor U4890 (N_4890,N_4091,N_4452);
and U4891 (N_4891,N_4264,N_4133);
xor U4892 (N_4892,N_4004,N_4020);
or U4893 (N_4893,N_4069,N_4054);
nor U4894 (N_4894,N_4167,N_4448);
and U4895 (N_4895,N_4085,N_4139);
or U4896 (N_4896,N_4092,N_4354);
nor U4897 (N_4897,N_4372,N_4467);
nor U4898 (N_4898,N_4163,N_4177);
or U4899 (N_4899,N_4106,N_4453);
nand U4900 (N_4900,N_4002,N_4426);
or U4901 (N_4901,N_4260,N_4147);
and U4902 (N_4902,N_4468,N_4222);
or U4903 (N_4903,N_4081,N_4219);
and U4904 (N_4904,N_4349,N_4495);
nor U4905 (N_4905,N_4270,N_4004);
and U4906 (N_4906,N_4202,N_4275);
nand U4907 (N_4907,N_4238,N_4314);
nor U4908 (N_4908,N_4360,N_4384);
nand U4909 (N_4909,N_4411,N_4082);
nor U4910 (N_4910,N_4441,N_4089);
and U4911 (N_4911,N_4336,N_4193);
nand U4912 (N_4912,N_4110,N_4377);
nor U4913 (N_4913,N_4255,N_4264);
or U4914 (N_4914,N_4134,N_4459);
nand U4915 (N_4915,N_4486,N_4065);
or U4916 (N_4916,N_4338,N_4280);
and U4917 (N_4917,N_4096,N_4238);
or U4918 (N_4918,N_4335,N_4239);
nand U4919 (N_4919,N_4016,N_4123);
and U4920 (N_4920,N_4173,N_4225);
xnor U4921 (N_4921,N_4372,N_4155);
nand U4922 (N_4922,N_4063,N_4264);
xnor U4923 (N_4923,N_4389,N_4418);
and U4924 (N_4924,N_4342,N_4084);
or U4925 (N_4925,N_4233,N_4443);
nor U4926 (N_4926,N_4011,N_4147);
xor U4927 (N_4927,N_4270,N_4446);
or U4928 (N_4928,N_4240,N_4114);
and U4929 (N_4929,N_4056,N_4358);
and U4930 (N_4930,N_4097,N_4080);
nor U4931 (N_4931,N_4449,N_4412);
nor U4932 (N_4932,N_4242,N_4287);
nand U4933 (N_4933,N_4248,N_4048);
or U4934 (N_4934,N_4303,N_4060);
or U4935 (N_4935,N_4243,N_4210);
nand U4936 (N_4936,N_4490,N_4039);
and U4937 (N_4937,N_4348,N_4131);
nor U4938 (N_4938,N_4438,N_4378);
and U4939 (N_4939,N_4089,N_4285);
or U4940 (N_4940,N_4176,N_4376);
and U4941 (N_4941,N_4292,N_4090);
nor U4942 (N_4942,N_4268,N_4370);
and U4943 (N_4943,N_4396,N_4191);
and U4944 (N_4944,N_4417,N_4427);
nand U4945 (N_4945,N_4261,N_4124);
nor U4946 (N_4946,N_4303,N_4368);
xor U4947 (N_4947,N_4089,N_4100);
nor U4948 (N_4948,N_4230,N_4040);
or U4949 (N_4949,N_4306,N_4445);
and U4950 (N_4950,N_4414,N_4185);
and U4951 (N_4951,N_4049,N_4125);
and U4952 (N_4952,N_4183,N_4485);
and U4953 (N_4953,N_4332,N_4090);
nor U4954 (N_4954,N_4373,N_4121);
xor U4955 (N_4955,N_4215,N_4295);
nand U4956 (N_4956,N_4093,N_4422);
and U4957 (N_4957,N_4314,N_4403);
nor U4958 (N_4958,N_4467,N_4497);
and U4959 (N_4959,N_4174,N_4455);
nor U4960 (N_4960,N_4021,N_4416);
and U4961 (N_4961,N_4471,N_4147);
nor U4962 (N_4962,N_4147,N_4153);
nand U4963 (N_4963,N_4299,N_4318);
nor U4964 (N_4964,N_4406,N_4126);
and U4965 (N_4965,N_4080,N_4417);
nor U4966 (N_4966,N_4247,N_4348);
nand U4967 (N_4967,N_4347,N_4352);
nand U4968 (N_4968,N_4067,N_4054);
and U4969 (N_4969,N_4140,N_4388);
nor U4970 (N_4970,N_4471,N_4312);
and U4971 (N_4971,N_4039,N_4235);
xor U4972 (N_4972,N_4199,N_4322);
nor U4973 (N_4973,N_4403,N_4411);
nor U4974 (N_4974,N_4056,N_4459);
and U4975 (N_4975,N_4125,N_4364);
xor U4976 (N_4976,N_4071,N_4243);
and U4977 (N_4977,N_4060,N_4439);
or U4978 (N_4978,N_4270,N_4208);
or U4979 (N_4979,N_4316,N_4499);
or U4980 (N_4980,N_4098,N_4333);
xor U4981 (N_4981,N_4067,N_4097);
or U4982 (N_4982,N_4489,N_4020);
and U4983 (N_4983,N_4273,N_4344);
nor U4984 (N_4984,N_4382,N_4383);
nor U4985 (N_4985,N_4329,N_4119);
or U4986 (N_4986,N_4301,N_4332);
nand U4987 (N_4987,N_4097,N_4475);
and U4988 (N_4988,N_4203,N_4413);
xnor U4989 (N_4989,N_4170,N_4319);
nand U4990 (N_4990,N_4228,N_4465);
and U4991 (N_4991,N_4441,N_4228);
or U4992 (N_4992,N_4306,N_4206);
or U4993 (N_4993,N_4252,N_4479);
or U4994 (N_4994,N_4099,N_4286);
or U4995 (N_4995,N_4089,N_4109);
or U4996 (N_4996,N_4380,N_4217);
and U4997 (N_4997,N_4220,N_4448);
nor U4998 (N_4998,N_4209,N_4307);
nand U4999 (N_4999,N_4162,N_4063);
nand U5000 (N_5000,N_4925,N_4563);
and U5001 (N_5001,N_4592,N_4725);
nor U5002 (N_5002,N_4971,N_4529);
and U5003 (N_5003,N_4933,N_4798);
nor U5004 (N_5004,N_4964,N_4961);
or U5005 (N_5005,N_4810,N_4537);
nor U5006 (N_5006,N_4712,N_4610);
and U5007 (N_5007,N_4700,N_4621);
nand U5008 (N_5008,N_4675,N_4573);
nand U5009 (N_5009,N_4570,N_4574);
xor U5010 (N_5010,N_4702,N_4545);
or U5011 (N_5011,N_4557,N_4784);
xnor U5012 (N_5012,N_4704,N_4865);
xnor U5013 (N_5013,N_4636,N_4951);
nor U5014 (N_5014,N_4821,N_4902);
or U5015 (N_5015,N_4713,N_4834);
and U5016 (N_5016,N_4604,N_4802);
nand U5017 (N_5017,N_4851,N_4750);
nor U5018 (N_5018,N_4624,N_4891);
nor U5019 (N_5019,N_4653,N_4658);
or U5020 (N_5020,N_4631,N_4895);
and U5021 (N_5021,N_4830,N_4781);
nor U5022 (N_5022,N_4936,N_4500);
nor U5023 (N_5023,N_4663,N_4870);
nand U5024 (N_5024,N_4540,N_4647);
or U5025 (N_5025,N_4643,N_4849);
or U5026 (N_5026,N_4659,N_4648);
nand U5027 (N_5027,N_4703,N_4609);
nor U5028 (N_5028,N_4950,N_4603);
and U5029 (N_5029,N_4728,N_4769);
nor U5030 (N_5030,N_4792,N_4770);
and U5031 (N_5031,N_4579,N_4926);
nor U5032 (N_5032,N_4789,N_4715);
xnor U5033 (N_5033,N_4670,N_4980);
nor U5034 (N_5034,N_4701,N_4732);
or U5035 (N_5035,N_4650,N_4800);
or U5036 (N_5036,N_4657,N_4873);
or U5037 (N_5037,N_4710,N_4743);
and U5038 (N_5038,N_4942,N_4917);
and U5039 (N_5039,N_4921,N_4782);
nand U5040 (N_5040,N_4813,N_4503);
nor U5041 (N_5041,N_4694,N_4930);
or U5042 (N_5042,N_4940,N_4958);
nand U5043 (N_5043,N_4556,N_4887);
or U5044 (N_5044,N_4542,N_4916);
nor U5045 (N_5045,N_4823,N_4532);
or U5046 (N_5046,N_4538,N_4594);
nor U5047 (N_5047,N_4763,N_4688);
and U5048 (N_5048,N_4667,N_4736);
xnor U5049 (N_5049,N_4999,N_4780);
and U5050 (N_5050,N_4669,N_4837);
and U5051 (N_5051,N_4854,N_4939);
nor U5052 (N_5052,N_4833,N_4880);
nor U5053 (N_5053,N_4533,N_4777);
nor U5054 (N_5054,N_4524,N_4518);
and U5055 (N_5055,N_4505,N_4581);
nor U5056 (N_5056,N_4835,N_4909);
or U5057 (N_5057,N_4779,N_4906);
or U5058 (N_5058,N_4944,N_4879);
and U5059 (N_5059,N_4672,N_4735);
or U5060 (N_5060,N_4730,N_4831);
or U5061 (N_5061,N_4978,N_4765);
and U5062 (N_5062,N_4803,N_4892);
and U5063 (N_5063,N_4908,N_4539);
nor U5064 (N_5064,N_4739,N_4508);
or U5065 (N_5065,N_4857,N_4741);
and U5066 (N_5066,N_4602,N_4668);
nand U5067 (N_5067,N_4824,N_4904);
xnor U5068 (N_5068,N_4787,N_4559);
or U5069 (N_5069,N_4804,N_4749);
xor U5070 (N_5070,N_4558,N_4501);
nor U5071 (N_5071,N_4687,N_4861);
nand U5072 (N_5072,N_4826,N_4593);
nor U5073 (N_5073,N_4948,N_4740);
and U5074 (N_5074,N_4774,N_4589);
nor U5075 (N_5075,N_4811,N_4843);
xor U5076 (N_5076,N_4981,N_4756);
xor U5077 (N_5077,N_4918,N_4967);
and U5078 (N_5078,N_4884,N_4711);
nor U5079 (N_5079,N_4796,N_4963);
nand U5080 (N_5080,N_4850,N_4731);
nand U5081 (N_5081,N_4753,N_4677);
nand U5082 (N_5082,N_4893,N_4869);
and U5083 (N_5083,N_4859,N_4615);
nor U5084 (N_5084,N_4896,N_4852);
or U5085 (N_5085,N_4528,N_4514);
nor U5086 (N_5086,N_4635,N_4520);
nand U5087 (N_5087,N_4553,N_4552);
and U5088 (N_5088,N_4513,N_4790);
nand U5089 (N_5089,N_4771,N_4973);
or U5090 (N_5090,N_4561,N_4705);
nor U5091 (N_5091,N_4760,N_4716);
nor U5092 (N_5092,N_4699,N_4901);
nor U5093 (N_5093,N_4706,N_4651);
or U5094 (N_5094,N_4630,N_4584);
nor U5095 (N_5095,N_4510,N_4975);
nand U5096 (N_5096,N_4633,N_4872);
nor U5097 (N_5097,N_4516,N_4686);
nand U5098 (N_5098,N_4748,N_4642);
or U5099 (N_5099,N_4759,N_4776);
and U5100 (N_5100,N_4847,N_4751);
nor U5101 (N_5101,N_4690,N_4511);
nor U5102 (N_5102,N_4785,N_4646);
nand U5103 (N_5103,N_4882,N_4761);
nand U5104 (N_5104,N_4995,N_4805);
or U5105 (N_5105,N_4640,N_4745);
nor U5106 (N_5106,N_4839,N_4827);
or U5107 (N_5107,N_4565,N_4877);
and U5108 (N_5108,N_4674,N_4814);
or U5109 (N_5109,N_4899,N_4866);
nor U5110 (N_5110,N_4575,N_4985);
and U5111 (N_5111,N_4838,N_4645);
nor U5112 (N_5112,N_4949,N_4519);
nor U5113 (N_5113,N_4543,N_4578);
and U5114 (N_5114,N_4910,N_4692);
and U5115 (N_5115,N_4606,N_4585);
or U5116 (N_5116,N_4591,N_4817);
and U5117 (N_5117,N_4938,N_4608);
and U5118 (N_5118,N_4729,N_4637);
xnor U5119 (N_5119,N_4816,N_4541);
or U5120 (N_5120,N_4620,N_4548);
nor U5121 (N_5121,N_4734,N_4726);
or U5122 (N_5122,N_4970,N_4569);
or U5123 (N_5123,N_4932,N_4818);
nor U5124 (N_5124,N_4587,N_4864);
nand U5125 (N_5125,N_4795,N_4616);
nand U5126 (N_5126,N_4515,N_4867);
nor U5127 (N_5127,N_4890,N_4812);
nand U5128 (N_5128,N_4502,N_4622);
and U5129 (N_5129,N_4571,N_4625);
and U5130 (N_5130,N_4664,N_4521);
or U5131 (N_5131,N_4959,N_4928);
nand U5132 (N_5132,N_4707,N_4860);
nor U5133 (N_5133,N_4517,N_4952);
xor U5134 (N_5134,N_4504,N_4768);
or U5135 (N_5135,N_4937,N_4871);
or U5136 (N_5136,N_4825,N_4568);
nor U5137 (N_5137,N_4679,N_4946);
and U5138 (N_5138,N_4927,N_4874);
xnor U5139 (N_5139,N_4644,N_4722);
or U5140 (N_5140,N_4767,N_4634);
xnor U5141 (N_5141,N_4778,N_4724);
nor U5142 (N_5142,N_4666,N_4684);
or U5143 (N_5143,N_4875,N_4691);
xor U5144 (N_5144,N_4992,N_4998);
nand U5145 (N_5145,N_4984,N_4689);
and U5146 (N_5146,N_4956,N_4526);
xor U5147 (N_5147,N_4791,N_4619);
xnor U5148 (N_5148,N_4617,N_4954);
nor U5149 (N_5149,N_4966,N_4661);
nor U5150 (N_5150,N_4993,N_4786);
nand U5151 (N_5151,N_4747,N_4986);
nand U5152 (N_5152,N_4962,N_4605);
nor U5153 (N_5153,N_4566,N_4564);
nor U5154 (N_5154,N_4754,N_4693);
nor U5155 (N_5155,N_4819,N_4652);
or U5156 (N_5156,N_4919,N_4885);
nor U5157 (N_5157,N_4665,N_4853);
nand U5158 (N_5158,N_4547,N_4947);
or U5159 (N_5159,N_4709,N_4590);
nand U5160 (N_5160,N_4912,N_4614);
or U5161 (N_5161,N_4828,N_4582);
nand U5162 (N_5162,N_4969,N_4600);
nand U5163 (N_5163,N_4613,N_4897);
and U5164 (N_5164,N_4595,N_4922);
nand U5165 (N_5165,N_4898,N_4836);
nor U5166 (N_5166,N_4611,N_4717);
xnor U5167 (N_5167,N_4876,N_4530);
or U5168 (N_5168,N_4991,N_4738);
nand U5169 (N_5169,N_4721,N_4943);
nand U5170 (N_5170,N_4878,N_4957);
nand U5171 (N_5171,N_4863,N_4913);
or U5172 (N_5172,N_4806,N_4977);
and U5173 (N_5173,N_4845,N_4746);
nor U5174 (N_5174,N_4755,N_4737);
or U5175 (N_5175,N_4960,N_4685);
xor U5176 (N_5176,N_4972,N_4544);
xnor U5177 (N_5177,N_4607,N_4588);
nor U5178 (N_5178,N_4742,N_4868);
and U5179 (N_5179,N_4577,N_4560);
xnor U5180 (N_5180,N_4920,N_4714);
and U5181 (N_5181,N_4822,N_4846);
xor U5182 (N_5182,N_4583,N_4994);
xnor U5183 (N_5183,N_4911,N_4979);
and U5184 (N_5184,N_4996,N_4681);
and U5185 (N_5185,N_4903,N_4723);
nand U5186 (N_5186,N_4799,N_4698);
and U5187 (N_5187,N_4881,N_4809);
or U5188 (N_5188,N_4509,N_4931);
nand U5189 (N_5189,N_4567,N_4976);
nand U5190 (N_5190,N_4599,N_4649);
and U5191 (N_5191,N_4989,N_4757);
nand U5192 (N_5192,N_4929,N_4934);
or U5193 (N_5193,N_4695,N_4546);
nor U5194 (N_5194,N_4855,N_4923);
or U5195 (N_5195,N_4525,N_4856);
nand U5196 (N_5196,N_4848,N_4788);
nand U5197 (N_5197,N_4900,N_4889);
nand U5198 (N_5198,N_4678,N_4844);
nor U5199 (N_5199,N_4727,N_4842);
and U5200 (N_5200,N_4586,N_4983);
nor U5201 (N_5201,N_4829,N_4550);
and U5202 (N_5202,N_4953,N_4862);
and U5203 (N_5203,N_4536,N_4820);
nor U5204 (N_5204,N_4627,N_4562);
and U5205 (N_5205,N_4907,N_4974);
nor U5206 (N_5206,N_4883,N_4612);
nand U5207 (N_5207,N_4965,N_4793);
nand U5208 (N_5208,N_4982,N_4534);
nor U5209 (N_5209,N_4915,N_4719);
nor U5210 (N_5210,N_4682,N_4894);
and U5211 (N_5211,N_4708,N_4758);
xnor U5212 (N_5212,N_4764,N_4801);
nand U5213 (N_5213,N_4718,N_4654);
nand U5214 (N_5214,N_4886,N_4914);
nor U5215 (N_5215,N_4531,N_4580);
nand U5216 (N_5216,N_4535,N_4744);
nand U5217 (N_5217,N_4945,N_4527);
and U5218 (N_5218,N_4680,N_4506);
nand U5219 (N_5219,N_4697,N_4696);
xnor U5220 (N_5220,N_4618,N_4572);
or U5221 (N_5221,N_4597,N_4671);
and U5222 (N_5222,N_4766,N_4840);
xor U5223 (N_5223,N_4673,N_4794);
and U5224 (N_5224,N_4752,N_4628);
nand U5225 (N_5225,N_4808,N_4997);
nor U5226 (N_5226,N_4555,N_4623);
nor U5227 (N_5227,N_4941,N_4655);
nor U5228 (N_5228,N_4639,N_4662);
nor U5229 (N_5229,N_4773,N_4775);
xnor U5230 (N_5230,N_4720,N_4832);
or U5231 (N_5231,N_4858,N_4598);
nand U5232 (N_5232,N_4807,N_4683);
nand U5233 (N_5233,N_4641,N_4783);
or U5234 (N_5234,N_4990,N_4762);
or U5235 (N_5235,N_4549,N_4955);
or U5236 (N_5236,N_4988,N_4924);
and U5237 (N_5237,N_4797,N_4601);
xnor U5238 (N_5238,N_4522,N_4888);
and U5239 (N_5239,N_4629,N_4638);
xor U5240 (N_5240,N_4632,N_4841);
nand U5241 (N_5241,N_4576,N_4656);
or U5242 (N_5242,N_4733,N_4968);
nor U5243 (N_5243,N_4987,N_4676);
and U5244 (N_5244,N_4596,N_4512);
nand U5245 (N_5245,N_4815,N_4554);
nor U5246 (N_5246,N_4551,N_4626);
or U5247 (N_5247,N_4772,N_4905);
and U5248 (N_5248,N_4523,N_4660);
xor U5249 (N_5249,N_4935,N_4507);
and U5250 (N_5250,N_4567,N_4864);
nand U5251 (N_5251,N_4979,N_4882);
nand U5252 (N_5252,N_4795,N_4741);
or U5253 (N_5253,N_4665,N_4762);
nor U5254 (N_5254,N_4783,N_4861);
xor U5255 (N_5255,N_4819,N_4566);
nand U5256 (N_5256,N_4577,N_4844);
xnor U5257 (N_5257,N_4656,N_4971);
or U5258 (N_5258,N_4668,N_4685);
nor U5259 (N_5259,N_4976,N_4646);
nand U5260 (N_5260,N_4539,N_4543);
nand U5261 (N_5261,N_4642,N_4555);
and U5262 (N_5262,N_4537,N_4687);
nand U5263 (N_5263,N_4787,N_4938);
nor U5264 (N_5264,N_4657,N_4938);
and U5265 (N_5265,N_4735,N_4664);
nand U5266 (N_5266,N_4739,N_4604);
nand U5267 (N_5267,N_4568,N_4786);
xnor U5268 (N_5268,N_4862,N_4952);
or U5269 (N_5269,N_4686,N_4800);
or U5270 (N_5270,N_4601,N_4788);
nand U5271 (N_5271,N_4546,N_4583);
and U5272 (N_5272,N_4504,N_4794);
nand U5273 (N_5273,N_4608,N_4553);
or U5274 (N_5274,N_4658,N_4971);
or U5275 (N_5275,N_4988,N_4765);
nand U5276 (N_5276,N_4601,N_4676);
nand U5277 (N_5277,N_4999,N_4975);
or U5278 (N_5278,N_4994,N_4802);
nand U5279 (N_5279,N_4568,N_4672);
nand U5280 (N_5280,N_4820,N_4774);
or U5281 (N_5281,N_4882,N_4948);
xor U5282 (N_5282,N_4894,N_4597);
or U5283 (N_5283,N_4887,N_4526);
and U5284 (N_5284,N_4768,N_4708);
or U5285 (N_5285,N_4714,N_4623);
or U5286 (N_5286,N_4764,N_4859);
nand U5287 (N_5287,N_4899,N_4562);
and U5288 (N_5288,N_4997,N_4573);
nor U5289 (N_5289,N_4586,N_4987);
nor U5290 (N_5290,N_4661,N_4595);
nor U5291 (N_5291,N_4861,N_4619);
nand U5292 (N_5292,N_4732,N_4995);
or U5293 (N_5293,N_4569,N_4724);
nor U5294 (N_5294,N_4851,N_4597);
and U5295 (N_5295,N_4565,N_4751);
nor U5296 (N_5296,N_4731,N_4846);
nor U5297 (N_5297,N_4510,N_4630);
and U5298 (N_5298,N_4753,N_4905);
or U5299 (N_5299,N_4787,N_4755);
or U5300 (N_5300,N_4968,N_4814);
xnor U5301 (N_5301,N_4716,N_4581);
or U5302 (N_5302,N_4790,N_4639);
nand U5303 (N_5303,N_4755,N_4811);
or U5304 (N_5304,N_4547,N_4886);
or U5305 (N_5305,N_4752,N_4601);
and U5306 (N_5306,N_4511,N_4869);
nand U5307 (N_5307,N_4641,N_4622);
or U5308 (N_5308,N_4595,N_4827);
nand U5309 (N_5309,N_4940,N_4819);
nor U5310 (N_5310,N_4705,N_4932);
and U5311 (N_5311,N_4574,N_4724);
nor U5312 (N_5312,N_4560,N_4767);
nor U5313 (N_5313,N_4508,N_4663);
and U5314 (N_5314,N_4609,N_4690);
and U5315 (N_5315,N_4751,N_4853);
and U5316 (N_5316,N_4834,N_4522);
nand U5317 (N_5317,N_4544,N_4518);
nor U5318 (N_5318,N_4825,N_4995);
or U5319 (N_5319,N_4768,N_4794);
and U5320 (N_5320,N_4925,N_4810);
nor U5321 (N_5321,N_4702,N_4961);
nand U5322 (N_5322,N_4697,N_4609);
or U5323 (N_5323,N_4743,N_4552);
nor U5324 (N_5324,N_4778,N_4846);
nand U5325 (N_5325,N_4538,N_4901);
nor U5326 (N_5326,N_4833,N_4678);
and U5327 (N_5327,N_4718,N_4910);
xor U5328 (N_5328,N_4629,N_4748);
and U5329 (N_5329,N_4668,N_4504);
nand U5330 (N_5330,N_4689,N_4892);
nand U5331 (N_5331,N_4829,N_4888);
and U5332 (N_5332,N_4608,N_4749);
and U5333 (N_5333,N_4686,N_4754);
nand U5334 (N_5334,N_4728,N_4505);
nor U5335 (N_5335,N_4951,N_4750);
and U5336 (N_5336,N_4573,N_4601);
nand U5337 (N_5337,N_4632,N_4926);
and U5338 (N_5338,N_4869,N_4914);
nand U5339 (N_5339,N_4777,N_4682);
and U5340 (N_5340,N_4992,N_4966);
nand U5341 (N_5341,N_4767,N_4814);
xnor U5342 (N_5342,N_4646,N_4925);
or U5343 (N_5343,N_4766,N_4871);
nor U5344 (N_5344,N_4863,N_4984);
nand U5345 (N_5345,N_4919,N_4720);
nand U5346 (N_5346,N_4884,N_4714);
nand U5347 (N_5347,N_4895,N_4787);
and U5348 (N_5348,N_4843,N_4823);
and U5349 (N_5349,N_4577,N_4836);
xnor U5350 (N_5350,N_4530,N_4885);
nor U5351 (N_5351,N_4716,N_4704);
or U5352 (N_5352,N_4940,N_4516);
nor U5353 (N_5353,N_4716,N_4684);
nor U5354 (N_5354,N_4955,N_4715);
nor U5355 (N_5355,N_4661,N_4938);
nand U5356 (N_5356,N_4849,N_4862);
xnor U5357 (N_5357,N_4685,N_4509);
and U5358 (N_5358,N_4873,N_4684);
or U5359 (N_5359,N_4559,N_4705);
xor U5360 (N_5360,N_4908,N_4510);
or U5361 (N_5361,N_4997,N_4598);
nor U5362 (N_5362,N_4938,N_4875);
and U5363 (N_5363,N_4925,N_4704);
nand U5364 (N_5364,N_4913,N_4611);
and U5365 (N_5365,N_4559,N_4704);
nand U5366 (N_5366,N_4687,N_4854);
xnor U5367 (N_5367,N_4607,N_4846);
or U5368 (N_5368,N_4867,N_4791);
and U5369 (N_5369,N_4765,N_4647);
nor U5370 (N_5370,N_4788,N_4722);
nand U5371 (N_5371,N_4544,N_4706);
nand U5372 (N_5372,N_4991,N_4944);
or U5373 (N_5373,N_4855,N_4777);
and U5374 (N_5374,N_4735,N_4958);
nor U5375 (N_5375,N_4739,N_4678);
and U5376 (N_5376,N_4887,N_4740);
xor U5377 (N_5377,N_4695,N_4616);
nor U5378 (N_5378,N_4570,N_4798);
and U5379 (N_5379,N_4648,N_4842);
nor U5380 (N_5380,N_4700,N_4753);
and U5381 (N_5381,N_4859,N_4820);
or U5382 (N_5382,N_4549,N_4975);
nand U5383 (N_5383,N_4596,N_4986);
nand U5384 (N_5384,N_4891,N_4712);
nor U5385 (N_5385,N_4672,N_4563);
nor U5386 (N_5386,N_4655,N_4756);
xor U5387 (N_5387,N_4895,N_4904);
and U5388 (N_5388,N_4648,N_4834);
or U5389 (N_5389,N_4515,N_4883);
nand U5390 (N_5390,N_4578,N_4573);
or U5391 (N_5391,N_4841,N_4993);
or U5392 (N_5392,N_4622,N_4646);
nor U5393 (N_5393,N_4921,N_4573);
and U5394 (N_5394,N_4744,N_4819);
and U5395 (N_5395,N_4869,N_4809);
nand U5396 (N_5396,N_4876,N_4573);
xor U5397 (N_5397,N_4953,N_4990);
and U5398 (N_5398,N_4999,N_4952);
or U5399 (N_5399,N_4830,N_4696);
nor U5400 (N_5400,N_4786,N_4506);
or U5401 (N_5401,N_4758,N_4833);
or U5402 (N_5402,N_4828,N_4876);
nor U5403 (N_5403,N_4823,N_4878);
and U5404 (N_5404,N_4569,N_4643);
and U5405 (N_5405,N_4881,N_4922);
or U5406 (N_5406,N_4716,N_4810);
and U5407 (N_5407,N_4711,N_4721);
and U5408 (N_5408,N_4905,N_4981);
xnor U5409 (N_5409,N_4502,N_4581);
or U5410 (N_5410,N_4775,N_4741);
or U5411 (N_5411,N_4966,N_4567);
nand U5412 (N_5412,N_4902,N_4654);
or U5413 (N_5413,N_4648,N_4552);
nand U5414 (N_5414,N_4914,N_4713);
nor U5415 (N_5415,N_4570,N_4619);
nor U5416 (N_5416,N_4731,N_4955);
or U5417 (N_5417,N_4564,N_4797);
and U5418 (N_5418,N_4608,N_4915);
xnor U5419 (N_5419,N_4999,N_4628);
nand U5420 (N_5420,N_4505,N_4731);
nand U5421 (N_5421,N_4893,N_4766);
and U5422 (N_5422,N_4910,N_4777);
or U5423 (N_5423,N_4515,N_4697);
nand U5424 (N_5424,N_4501,N_4968);
and U5425 (N_5425,N_4788,N_4910);
nor U5426 (N_5426,N_4592,N_4726);
nor U5427 (N_5427,N_4998,N_4820);
nand U5428 (N_5428,N_4593,N_4683);
or U5429 (N_5429,N_4976,N_4968);
nor U5430 (N_5430,N_4594,N_4552);
or U5431 (N_5431,N_4848,N_4664);
and U5432 (N_5432,N_4593,N_4751);
and U5433 (N_5433,N_4756,N_4874);
or U5434 (N_5434,N_4979,N_4645);
nor U5435 (N_5435,N_4577,N_4692);
and U5436 (N_5436,N_4874,N_4657);
or U5437 (N_5437,N_4645,N_4688);
xor U5438 (N_5438,N_4572,N_4606);
nand U5439 (N_5439,N_4881,N_4926);
nand U5440 (N_5440,N_4504,N_4775);
and U5441 (N_5441,N_4590,N_4829);
nor U5442 (N_5442,N_4653,N_4643);
nand U5443 (N_5443,N_4935,N_4541);
nor U5444 (N_5444,N_4966,N_4923);
and U5445 (N_5445,N_4754,N_4667);
and U5446 (N_5446,N_4699,N_4649);
or U5447 (N_5447,N_4740,N_4805);
nor U5448 (N_5448,N_4949,N_4520);
nand U5449 (N_5449,N_4824,N_4885);
nor U5450 (N_5450,N_4783,N_4621);
and U5451 (N_5451,N_4993,N_4618);
and U5452 (N_5452,N_4783,N_4505);
nor U5453 (N_5453,N_4679,N_4754);
nand U5454 (N_5454,N_4517,N_4831);
xor U5455 (N_5455,N_4585,N_4634);
xnor U5456 (N_5456,N_4665,N_4939);
and U5457 (N_5457,N_4865,N_4782);
nand U5458 (N_5458,N_4536,N_4557);
or U5459 (N_5459,N_4872,N_4754);
nand U5460 (N_5460,N_4773,N_4835);
or U5461 (N_5461,N_4845,N_4596);
or U5462 (N_5462,N_4585,N_4564);
nor U5463 (N_5463,N_4559,N_4925);
and U5464 (N_5464,N_4825,N_4782);
nand U5465 (N_5465,N_4544,N_4637);
nand U5466 (N_5466,N_4900,N_4855);
or U5467 (N_5467,N_4739,N_4547);
or U5468 (N_5468,N_4795,N_4860);
or U5469 (N_5469,N_4621,N_4920);
xnor U5470 (N_5470,N_4838,N_4936);
or U5471 (N_5471,N_4884,N_4575);
or U5472 (N_5472,N_4886,N_4850);
and U5473 (N_5473,N_4642,N_4750);
nand U5474 (N_5474,N_4754,N_4550);
or U5475 (N_5475,N_4632,N_4707);
nand U5476 (N_5476,N_4504,N_4544);
and U5477 (N_5477,N_4752,N_4591);
and U5478 (N_5478,N_4925,N_4697);
or U5479 (N_5479,N_4617,N_4734);
or U5480 (N_5480,N_4506,N_4876);
xnor U5481 (N_5481,N_4889,N_4806);
nor U5482 (N_5482,N_4967,N_4544);
nand U5483 (N_5483,N_4934,N_4984);
and U5484 (N_5484,N_4593,N_4942);
nand U5485 (N_5485,N_4950,N_4802);
nand U5486 (N_5486,N_4720,N_4963);
and U5487 (N_5487,N_4792,N_4700);
nor U5488 (N_5488,N_4548,N_4854);
or U5489 (N_5489,N_4651,N_4792);
and U5490 (N_5490,N_4743,N_4901);
nand U5491 (N_5491,N_4569,N_4607);
or U5492 (N_5492,N_4572,N_4672);
nand U5493 (N_5493,N_4821,N_4781);
and U5494 (N_5494,N_4846,N_4777);
nand U5495 (N_5495,N_4783,N_4642);
or U5496 (N_5496,N_4784,N_4895);
nor U5497 (N_5497,N_4744,N_4714);
and U5498 (N_5498,N_4580,N_4677);
nand U5499 (N_5499,N_4582,N_4524);
and U5500 (N_5500,N_5332,N_5218);
nand U5501 (N_5501,N_5117,N_5273);
nor U5502 (N_5502,N_5100,N_5188);
nor U5503 (N_5503,N_5392,N_5461);
nor U5504 (N_5504,N_5370,N_5413);
and U5505 (N_5505,N_5038,N_5293);
or U5506 (N_5506,N_5208,N_5079);
nand U5507 (N_5507,N_5118,N_5399);
and U5508 (N_5508,N_5158,N_5252);
xnor U5509 (N_5509,N_5357,N_5396);
xor U5510 (N_5510,N_5334,N_5155);
nor U5511 (N_5511,N_5416,N_5395);
or U5512 (N_5512,N_5466,N_5437);
and U5513 (N_5513,N_5064,N_5050);
nand U5514 (N_5514,N_5485,N_5260);
nand U5515 (N_5515,N_5164,N_5135);
nand U5516 (N_5516,N_5367,N_5228);
nor U5517 (N_5517,N_5402,N_5156);
nand U5518 (N_5518,N_5148,N_5033);
or U5519 (N_5519,N_5318,N_5199);
nand U5520 (N_5520,N_5363,N_5078);
nor U5521 (N_5521,N_5207,N_5283);
nand U5522 (N_5522,N_5264,N_5397);
and U5523 (N_5523,N_5234,N_5274);
and U5524 (N_5524,N_5312,N_5240);
xnor U5525 (N_5525,N_5376,N_5464);
and U5526 (N_5526,N_5123,N_5230);
nor U5527 (N_5527,N_5095,N_5315);
nor U5528 (N_5528,N_5089,N_5458);
and U5529 (N_5529,N_5422,N_5446);
or U5530 (N_5530,N_5069,N_5119);
xor U5531 (N_5531,N_5304,N_5111);
or U5532 (N_5532,N_5390,N_5006);
xnor U5533 (N_5533,N_5453,N_5190);
or U5534 (N_5534,N_5270,N_5113);
nor U5535 (N_5535,N_5369,N_5206);
and U5536 (N_5536,N_5091,N_5420);
nor U5537 (N_5537,N_5114,N_5306);
and U5538 (N_5538,N_5452,N_5439);
and U5539 (N_5539,N_5349,N_5434);
nand U5540 (N_5540,N_5368,N_5484);
nor U5541 (N_5541,N_5298,N_5398);
and U5542 (N_5542,N_5233,N_5125);
or U5543 (N_5543,N_5300,N_5004);
nor U5544 (N_5544,N_5179,N_5441);
nor U5545 (N_5545,N_5407,N_5449);
or U5546 (N_5546,N_5163,N_5442);
nand U5547 (N_5547,N_5198,N_5284);
and U5548 (N_5548,N_5126,N_5140);
or U5549 (N_5549,N_5288,N_5018);
or U5550 (N_5550,N_5122,N_5302);
nand U5551 (N_5551,N_5007,N_5251);
and U5552 (N_5552,N_5154,N_5428);
nand U5553 (N_5553,N_5189,N_5301);
nor U5554 (N_5554,N_5328,N_5414);
nor U5555 (N_5555,N_5450,N_5011);
nor U5556 (N_5556,N_5237,N_5292);
or U5557 (N_5557,N_5146,N_5393);
or U5558 (N_5558,N_5058,N_5444);
nand U5559 (N_5559,N_5480,N_5287);
nor U5560 (N_5560,N_5411,N_5039);
or U5561 (N_5561,N_5223,N_5265);
or U5562 (N_5562,N_5020,N_5204);
nand U5563 (N_5563,N_5305,N_5098);
xnor U5564 (N_5564,N_5329,N_5102);
and U5565 (N_5565,N_5291,N_5219);
or U5566 (N_5566,N_5105,N_5025);
and U5567 (N_5567,N_5479,N_5253);
nor U5568 (N_5568,N_5465,N_5350);
and U5569 (N_5569,N_5391,N_5195);
nor U5570 (N_5570,N_5131,N_5296);
nor U5571 (N_5571,N_5436,N_5250);
xnor U5572 (N_5572,N_5375,N_5055);
nor U5573 (N_5573,N_5435,N_5071);
and U5574 (N_5574,N_5415,N_5462);
nand U5575 (N_5575,N_5157,N_5335);
nand U5576 (N_5576,N_5197,N_5244);
nor U5577 (N_5577,N_5320,N_5322);
and U5578 (N_5578,N_5331,N_5389);
nand U5579 (N_5579,N_5262,N_5343);
xnor U5580 (N_5580,N_5333,N_5239);
xnor U5581 (N_5581,N_5068,N_5168);
nand U5582 (N_5582,N_5307,N_5238);
xor U5583 (N_5583,N_5259,N_5232);
or U5584 (N_5584,N_5088,N_5133);
and U5585 (N_5585,N_5182,N_5371);
and U5586 (N_5586,N_5108,N_5077);
nor U5587 (N_5587,N_5241,N_5027);
or U5588 (N_5588,N_5203,N_5001);
nor U5589 (N_5589,N_5115,N_5213);
or U5590 (N_5590,N_5438,N_5469);
nand U5591 (N_5591,N_5495,N_5021);
or U5592 (N_5592,N_5431,N_5445);
or U5593 (N_5593,N_5215,N_5366);
nor U5594 (N_5594,N_5022,N_5073);
or U5595 (N_5595,N_5016,N_5483);
nor U5596 (N_5596,N_5472,N_5120);
nor U5597 (N_5597,N_5171,N_5187);
nor U5598 (N_5598,N_5319,N_5498);
nor U5599 (N_5599,N_5344,N_5191);
and U5600 (N_5600,N_5165,N_5267);
nor U5601 (N_5601,N_5476,N_5327);
and U5602 (N_5602,N_5192,N_5275);
nor U5603 (N_5603,N_5005,N_5013);
or U5604 (N_5604,N_5268,N_5426);
nor U5605 (N_5605,N_5217,N_5003);
and U5606 (N_5606,N_5432,N_5070);
or U5607 (N_5607,N_5324,N_5104);
and U5608 (N_5608,N_5072,N_5227);
or U5609 (N_5609,N_5053,N_5313);
and U5610 (N_5610,N_5258,N_5385);
nand U5611 (N_5611,N_5460,N_5271);
nor U5612 (N_5612,N_5345,N_5030);
or U5613 (N_5613,N_5099,N_5184);
nand U5614 (N_5614,N_5356,N_5201);
and U5615 (N_5615,N_5278,N_5294);
nand U5616 (N_5616,N_5497,N_5346);
nand U5617 (N_5617,N_5037,N_5257);
nor U5618 (N_5618,N_5311,N_5143);
and U5619 (N_5619,N_5170,N_5412);
and U5620 (N_5620,N_5128,N_5051);
or U5621 (N_5621,N_5137,N_5153);
or U5622 (N_5622,N_5010,N_5121);
nand U5623 (N_5623,N_5196,N_5085);
and U5624 (N_5624,N_5309,N_5231);
or U5625 (N_5625,N_5417,N_5277);
and U5626 (N_5626,N_5295,N_5242);
nor U5627 (N_5627,N_5372,N_5141);
and U5628 (N_5628,N_5289,N_5193);
and U5629 (N_5629,N_5377,N_5132);
nor U5630 (N_5630,N_5008,N_5235);
nor U5631 (N_5631,N_5029,N_5222);
nand U5632 (N_5632,N_5477,N_5167);
and U5633 (N_5633,N_5076,N_5359);
or U5634 (N_5634,N_5427,N_5059);
and U5635 (N_5635,N_5381,N_5379);
or U5636 (N_5636,N_5116,N_5134);
and U5637 (N_5637,N_5430,N_5127);
and U5638 (N_5638,N_5130,N_5418);
xor U5639 (N_5639,N_5455,N_5488);
nor U5640 (N_5640,N_5012,N_5202);
nor U5641 (N_5641,N_5049,N_5405);
nor U5642 (N_5642,N_5063,N_5310);
nor U5643 (N_5643,N_5026,N_5378);
or U5644 (N_5644,N_5261,N_5360);
and U5645 (N_5645,N_5496,N_5145);
nor U5646 (N_5646,N_5124,N_5400);
nor U5647 (N_5647,N_5308,N_5220);
or U5648 (N_5648,N_5280,N_5348);
nand U5649 (N_5649,N_5406,N_5245);
nor U5650 (N_5650,N_5107,N_5110);
or U5651 (N_5651,N_5106,N_5173);
nor U5652 (N_5652,N_5354,N_5282);
xnor U5653 (N_5653,N_5060,N_5478);
nand U5654 (N_5654,N_5456,N_5314);
nor U5655 (N_5655,N_5249,N_5044);
and U5656 (N_5656,N_5255,N_5093);
or U5657 (N_5657,N_5246,N_5052);
nand U5658 (N_5658,N_5474,N_5147);
nor U5659 (N_5659,N_5419,N_5440);
and U5660 (N_5660,N_5303,N_5321);
nor U5661 (N_5661,N_5347,N_5338);
xnor U5662 (N_5662,N_5224,N_5373);
and U5663 (N_5663,N_5183,N_5162);
or U5664 (N_5664,N_5180,N_5457);
xor U5665 (N_5665,N_5243,N_5043);
xnor U5666 (N_5666,N_5225,N_5185);
xor U5667 (N_5667,N_5355,N_5035);
nor U5668 (N_5668,N_5492,N_5087);
nand U5669 (N_5669,N_5097,N_5149);
or U5670 (N_5670,N_5493,N_5212);
nor U5671 (N_5671,N_5263,N_5177);
nand U5672 (N_5672,N_5086,N_5279);
or U5673 (N_5673,N_5172,N_5388);
nand U5674 (N_5674,N_5297,N_5139);
xor U5675 (N_5675,N_5336,N_5205);
nand U5676 (N_5676,N_5254,N_5491);
or U5677 (N_5677,N_5341,N_5017);
or U5678 (N_5678,N_5326,N_5423);
and U5679 (N_5679,N_5383,N_5463);
xor U5680 (N_5680,N_5339,N_5160);
nand U5681 (N_5681,N_5403,N_5325);
nor U5682 (N_5682,N_5019,N_5054);
xor U5683 (N_5683,N_5286,N_5210);
and U5684 (N_5684,N_5353,N_5061);
nor U5685 (N_5685,N_5216,N_5066);
xor U5686 (N_5686,N_5090,N_5394);
and U5687 (N_5687,N_5045,N_5150);
nand U5688 (N_5688,N_5015,N_5358);
or U5689 (N_5689,N_5136,N_5481);
or U5690 (N_5690,N_5074,N_5471);
nand U5691 (N_5691,N_5384,N_5489);
or U5692 (N_5692,N_5151,N_5009);
nand U5693 (N_5693,N_5083,N_5459);
nor U5694 (N_5694,N_5036,N_5034);
or U5695 (N_5695,N_5214,N_5057);
nor U5696 (N_5696,N_5386,N_5065);
nand U5697 (N_5697,N_5067,N_5032);
nand U5698 (N_5698,N_5424,N_5129);
or U5699 (N_5699,N_5473,N_5159);
and U5700 (N_5700,N_5142,N_5092);
and U5701 (N_5701,N_5028,N_5194);
or U5702 (N_5702,N_5200,N_5443);
nand U5703 (N_5703,N_5340,N_5316);
or U5704 (N_5704,N_5175,N_5075);
xnor U5705 (N_5705,N_5425,N_5330);
nand U5706 (N_5706,N_5209,N_5081);
xnor U5707 (N_5707,N_5490,N_5470);
nand U5708 (N_5708,N_5031,N_5002);
nand U5709 (N_5709,N_5364,N_5062);
nor U5710 (N_5710,N_5352,N_5323);
xnor U5711 (N_5711,N_5176,N_5454);
and U5712 (N_5712,N_5221,N_5266);
and U5713 (N_5713,N_5467,N_5211);
xnor U5714 (N_5714,N_5236,N_5361);
and U5715 (N_5715,N_5109,N_5144);
and U5716 (N_5716,N_5169,N_5112);
or U5717 (N_5717,N_5276,N_5451);
xor U5718 (N_5718,N_5408,N_5024);
and U5719 (N_5719,N_5166,N_5499);
and U5720 (N_5720,N_5101,N_5269);
or U5721 (N_5721,N_5401,N_5014);
or U5722 (N_5722,N_5048,N_5365);
nor U5723 (N_5723,N_5475,N_5421);
nand U5724 (N_5724,N_5299,N_5337);
nor U5725 (N_5725,N_5174,N_5447);
or U5726 (N_5726,N_5256,N_5103);
or U5727 (N_5727,N_5161,N_5494);
and U5728 (N_5728,N_5023,N_5290);
nand U5729 (N_5729,N_5186,N_5486);
or U5730 (N_5730,N_5042,N_5468);
xnor U5731 (N_5731,N_5433,N_5281);
or U5732 (N_5732,N_5084,N_5317);
or U5733 (N_5733,N_5047,N_5096);
and U5734 (N_5734,N_5248,N_5152);
and U5735 (N_5735,N_5046,N_5374);
nor U5736 (N_5736,N_5387,N_5272);
or U5737 (N_5737,N_5181,N_5362);
nand U5738 (N_5738,N_5229,N_5482);
nor U5739 (N_5739,N_5226,N_5080);
or U5740 (N_5740,N_5138,N_5448);
nor U5741 (N_5741,N_5285,N_5040);
nand U5742 (N_5742,N_5247,N_5056);
nor U5743 (N_5743,N_5178,N_5000);
and U5744 (N_5744,N_5409,N_5382);
nand U5745 (N_5745,N_5082,N_5404);
or U5746 (N_5746,N_5094,N_5410);
nand U5747 (N_5747,N_5429,N_5342);
or U5748 (N_5748,N_5380,N_5487);
nand U5749 (N_5749,N_5041,N_5351);
and U5750 (N_5750,N_5484,N_5033);
nor U5751 (N_5751,N_5389,N_5077);
or U5752 (N_5752,N_5212,N_5030);
xnor U5753 (N_5753,N_5113,N_5011);
nor U5754 (N_5754,N_5193,N_5005);
or U5755 (N_5755,N_5307,N_5275);
and U5756 (N_5756,N_5399,N_5100);
nor U5757 (N_5757,N_5454,N_5453);
and U5758 (N_5758,N_5394,N_5488);
and U5759 (N_5759,N_5145,N_5142);
nor U5760 (N_5760,N_5115,N_5496);
or U5761 (N_5761,N_5271,N_5372);
nor U5762 (N_5762,N_5198,N_5333);
and U5763 (N_5763,N_5400,N_5492);
xor U5764 (N_5764,N_5411,N_5485);
or U5765 (N_5765,N_5478,N_5305);
nor U5766 (N_5766,N_5382,N_5383);
nor U5767 (N_5767,N_5259,N_5086);
xor U5768 (N_5768,N_5094,N_5269);
and U5769 (N_5769,N_5462,N_5061);
nand U5770 (N_5770,N_5227,N_5025);
nand U5771 (N_5771,N_5105,N_5229);
nor U5772 (N_5772,N_5499,N_5006);
and U5773 (N_5773,N_5086,N_5450);
nand U5774 (N_5774,N_5463,N_5232);
nand U5775 (N_5775,N_5296,N_5137);
nor U5776 (N_5776,N_5019,N_5136);
and U5777 (N_5777,N_5353,N_5410);
nor U5778 (N_5778,N_5204,N_5109);
nor U5779 (N_5779,N_5177,N_5447);
nor U5780 (N_5780,N_5389,N_5335);
xnor U5781 (N_5781,N_5338,N_5197);
or U5782 (N_5782,N_5197,N_5194);
nand U5783 (N_5783,N_5088,N_5105);
or U5784 (N_5784,N_5124,N_5100);
or U5785 (N_5785,N_5481,N_5322);
or U5786 (N_5786,N_5468,N_5109);
nor U5787 (N_5787,N_5178,N_5294);
and U5788 (N_5788,N_5186,N_5049);
or U5789 (N_5789,N_5272,N_5245);
or U5790 (N_5790,N_5469,N_5288);
nand U5791 (N_5791,N_5447,N_5286);
nor U5792 (N_5792,N_5225,N_5409);
xor U5793 (N_5793,N_5496,N_5385);
or U5794 (N_5794,N_5073,N_5275);
and U5795 (N_5795,N_5354,N_5080);
and U5796 (N_5796,N_5115,N_5311);
and U5797 (N_5797,N_5007,N_5299);
nand U5798 (N_5798,N_5124,N_5019);
or U5799 (N_5799,N_5467,N_5113);
nor U5800 (N_5800,N_5024,N_5232);
nor U5801 (N_5801,N_5448,N_5488);
nor U5802 (N_5802,N_5248,N_5085);
nand U5803 (N_5803,N_5296,N_5008);
nand U5804 (N_5804,N_5436,N_5067);
nor U5805 (N_5805,N_5291,N_5188);
or U5806 (N_5806,N_5364,N_5239);
or U5807 (N_5807,N_5204,N_5021);
nand U5808 (N_5808,N_5433,N_5405);
or U5809 (N_5809,N_5271,N_5231);
or U5810 (N_5810,N_5215,N_5418);
or U5811 (N_5811,N_5446,N_5211);
nor U5812 (N_5812,N_5372,N_5230);
nor U5813 (N_5813,N_5238,N_5203);
nand U5814 (N_5814,N_5217,N_5398);
nand U5815 (N_5815,N_5176,N_5035);
and U5816 (N_5816,N_5348,N_5460);
or U5817 (N_5817,N_5262,N_5017);
nor U5818 (N_5818,N_5333,N_5156);
and U5819 (N_5819,N_5392,N_5044);
nand U5820 (N_5820,N_5360,N_5456);
nand U5821 (N_5821,N_5474,N_5107);
nand U5822 (N_5822,N_5073,N_5214);
nand U5823 (N_5823,N_5111,N_5094);
nor U5824 (N_5824,N_5001,N_5445);
nor U5825 (N_5825,N_5498,N_5137);
nand U5826 (N_5826,N_5303,N_5499);
nor U5827 (N_5827,N_5187,N_5369);
nor U5828 (N_5828,N_5373,N_5238);
nand U5829 (N_5829,N_5022,N_5321);
or U5830 (N_5830,N_5189,N_5328);
nand U5831 (N_5831,N_5164,N_5443);
nand U5832 (N_5832,N_5463,N_5015);
and U5833 (N_5833,N_5100,N_5297);
nor U5834 (N_5834,N_5115,N_5486);
or U5835 (N_5835,N_5291,N_5118);
or U5836 (N_5836,N_5444,N_5245);
xor U5837 (N_5837,N_5022,N_5290);
or U5838 (N_5838,N_5074,N_5277);
and U5839 (N_5839,N_5029,N_5169);
or U5840 (N_5840,N_5292,N_5408);
or U5841 (N_5841,N_5260,N_5387);
nand U5842 (N_5842,N_5385,N_5001);
xor U5843 (N_5843,N_5452,N_5333);
nand U5844 (N_5844,N_5243,N_5086);
nor U5845 (N_5845,N_5316,N_5222);
or U5846 (N_5846,N_5495,N_5155);
nor U5847 (N_5847,N_5185,N_5244);
and U5848 (N_5848,N_5268,N_5309);
or U5849 (N_5849,N_5415,N_5113);
or U5850 (N_5850,N_5364,N_5455);
or U5851 (N_5851,N_5401,N_5333);
nand U5852 (N_5852,N_5246,N_5268);
nor U5853 (N_5853,N_5420,N_5416);
nand U5854 (N_5854,N_5370,N_5148);
or U5855 (N_5855,N_5274,N_5440);
nor U5856 (N_5856,N_5184,N_5487);
nand U5857 (N_5857,N_5197,N_5233);
and U5858 (N_5858,N_5396,N_5382);
nor U5859 (N_5859,N_5423,N_5353);
and U5860 (N_5860,N_5076,N_5167);
nand U5861 (N_5861,N_5244,N_5474);
or U5862 (N_5862,N_5019,N_5482);
nor U5863 (N_5863,N_5459,N_5016);
nor U5864 (N_5864,N_5211,N_5483);
or U5865 (N_5865,N_5428,N_5454);
nand U5866 (N_5866,N_5327,N_5379);
nor U5867 (N_5867,N_5283,N_5384);
nand U5868 (N_5868,N_5025,N_5225);
nand U5869 (N_5869,N_5099,N_5054);
nand U5870 (N_5870,N_5448,N_5279);
and U5871 (N_5871,N_5093,N_5364);
nor U5872 (N_5872,N_5404,N_5192);
and U5873 (N_5873,N_5490,N_5334);
xnor U5874 (N_5874,N_5136,N_5229);
and U5875 (N_5875,N_5004,N_5417);
nand U5876 (N_5876,N_5493,N_5403);
and U5877 (N_5877,N_5064,N_5252);
and U5878 (N_5878,N_5377,N_5042);
or U5879 (N_5879,N_5284,N_5057);
nand U5880 (N_5880,N_5096,N_5210);
nand U5881 (N_5881,N_5038,N_5334);
or U5882 (N_5882,N_5160,N_5484);
or U5883 (N_5883,N_5400,N_5377);
nor U5884 (N_5884,N_5049,N_5028);
or U5885 (N_5885,N_5039,N_5252);
and U5886 (N_5886,N_5357,N_5226);
or U5887 (N_5887,N_5486,N_5216);
nand U5888 (N_5888,N_5446,N_5358);
and U5889 (N_5889,N_5047,N_5452);
xnor U5890 (N_5890,N_5406,N_5254);
xnor U5891 (N_5891,N_5081,N_5265);
or U5892 (N_5892,N_5447,N_5142);
and U5893 (N_5893,N_5333,N_5369);
nor U5894 (N_5894,N_5408,N_5315);
and U5895 (N_5895,N_5062,N_5194);
and U5896 (N_5896,N_5370,N_5241);
nand U5897 (N_5897,N_5222,N_5294);
xnor U5898 (N_5898,N_5086,N_5064);
nor U5899 (N_5899,N_5005,N_5194);
or U5900 (N_5900,N_5202,N_5242);
and U5901 (N_5901,N_5278,N_5313);
nand U5902 (N_5902,N_5480,N_5026);
nor U5903 (N_5903,N_5398,N_5253);
and U5904 (N_5904,N_5252,N_5166);
and U5905 (N_5905,N_5434,N_5440);
xnor U5906 (N_5906,N_5288,N_5229);
nor U5907 (N_5907,N_5463,N_5330);
nand U5908 (N_5908,N_5424,N_5156);
nand U5909 (N_5909,N_5130,N_5098);
xor U5910 (N_5910,N_5205,N_5282);
or U5911 (N_5911,N_5136,N_5360);
nand U5912 (N_5912,N_5081,N_5282);
nor U5913 (N_5913,N_5236,N_5274);
nand U5914 (N_5914,N_5168,N_5222);
and U5915 (N_5915,N_5287,N_5477);
nor U5916 (N_5916,N_5352,N_5036);
and U5917 (N_5917,N_5182,N_5179);
nand U5918 (N_5918,N_5235,N_5111);
xnor U5919 (N_5919,N_5032,N_5407);
or U5920 (N_5920,N_5217,N_5218);
xnor U5921 (N_5921,N_5079,N_5451);
xor U5922 (N_5922,N_5263,N_5184);
and U5923 (N_5923,N_5302,N_5339);
nor U5924 (N_5924,N_5027,N_5293);
nand U5925 (N_5925,N_5153,N_5218);
nand U5926 (N_5926,N_5379,N_5323);
and U5927 (N_5927,N_5202,N_5254);
and U5928 (N_5928,N_5016,N_5463);
and U5929 (N_5929,N_5467,N_5436);
and U5930 (N_5930,N_5126,N_5358);
xnor U5931 (N_5931,N_5321,N_5147);
nor U5932 (N_5932,N_5162,N_5471);
nor U5933 (N_5933,N_5150,N_5464);
or U5934 (N_5934,N_5221,N_5465);
and U5935 (N_5935,N_5389,N_5233);
and U5936 (N_5936,N_5480,N_5324);
nor U5937 (N_5937,N_5481,N_5460);
nor U5938 (N_5938,N_5159,N_5330);
nor U5939 (N_5939,N_5308,N_5482);
nand U5940 (N_5940,N_5268,N_5422);
and U5941 (N_5941,N_5285,N_5093);
or U5942 (N_5942,N_5353,N_5464);
nor U5943 (N_5943,N_5384,N_5214);
and U5944 (N_5944,N_5010,N_5090);
and U5945 (N_5945,N_5239,N_5291);
nand U5946 (N_5946,N_5121,N_5315);
xor U5947 (N_5947,N_5101,N_5000);
xor U5948 (N_5948,N_5084,N_5269);
and U5949 (N_5949,N_5398,N_5025);
nand U5950 (N_5950,N_5116,N_5401);
nor U5951 (N_5951,N_5354,N_5281);
or U5952 (N_5952,N_5272,N_5141);
nand U5953 (N_5953,N_5400,N_5379);
nor U5954 (N_5954,N_5164,N_5416);
nor U5955 (N_5955,N_5322,N_5222);
and U5956 (N_5956,N_5312,N_5423);
nor U5957 (N_5957,N_5326,N_5219);
nor U5958 (N_5958,N_5182,N_5016);
nand U5959 (N_5959,N_5308,N_5261);
or U5960 (N_5960,N_5222,N_5114);
nand U5961 (N_5961,N_5455,N_5102);
nand U5962 (N_5962,N_5277,N_5409);
and U5963 (N_5963,N_5085,N_5309);
and U5964 (N_5964,N_5016,N_5264);
or U5965 (N_5965,N_5319,N_5152);
or U5966 (N_5966,N_5270,N_5211);
xnor U5967 (N_5967,N_5162,N_5105);
and U5968 (N_5968,N_5224,N_5288);
xnor U5969 (N_5969,N_5380,N_5259);
nor U5970 (N_5970,N_5193,N_5160);
or U5971 (N_5971,N_5120,N_5186);
nand U5972 (N_5972,N_5380,N_5464);
nor U5973 (N_5973,N_5102,N_5412);
nor U5974 (N_5974,N_5276,N_5201);
nand U5975 (N_5975,N_5219,N_5095);
nor U5976 (N_5976,N_5233,N_5245);
nand U5977 (N_5977,N_5406,N_5306);
or U5978 (N_5978,N_5156,N_5076);
nor U5979 (N_5979,N_5145,N_5283);
and U5980 (N_5980,N_5456,N_5311);
and U5981 (N_5981,N_5230,N_5213);
xor U5982 (N_5982,N_5206,N_5213);
nor U5983 (N_5983,N_5310,N_5105);
nand U5984 (N_5984,N_5315,N_5254);
or U5985 (N_5985,N_5404,N_5280);
nor U5986 (N_5986,N_5443,N_5252);
and U5987 (N_5987,N_5040,N_5134);
or U5988 (N_5988,N_5471,N_5207);
nand U5989 (N_5989,N_5026,N_5431);
nor U5990 (N_5990,N_5048,N_5346);
xor U5991 (N_5991,N_5114,N_5409);
or U5992 (N_5992,N_5041,N_5065);
nand U5993 (N_5993,N_5362,N_5075);
nand U5994 (N_5994,N_5440,N_5112);
and U5995 (N_5995,N_5329,N_5120);
nor U5996 (N_5996,N_5417,N_5317);
xor U5997 (N_5997,N_5156,N_5134);
xnor U5998 (N_5998,N_5206,N_5097);
nor U5999 (N_5999,N_5001,N_5479);
or U6000 (N_6000,N_5658,N_5524);
nand U6001 (N_6001,N_5593,N_5928);
or U6002 (N_6002,N_5621,N_5839);
and U6003 (N_6003,N_5823,N_5574);
or U6004 (N_6004,N_5889,N_5773);
or U6005 (N_6005,N_5608,N_5627);
and U6006 (N_6006,N_5921,N_5724);
nand U6007 (N_6007,N_5519,N_5675);
and U6008 (N_6008,N_5596,N_5742);
nand U6009 (N_6009,N_5576,N_5886);
nand U6010 (N_6010,N_5753,N_5704);
and U6011 (N_6011,N_5984,N_5965);
and U6012 (N_6012,N_5817,N_5547);
or U6013 (N_6013,N_5580,N_5629);
and U6014 (N_6014,N_5783,N_5535);
or U6015 (N_6015,N_5611,N_5897);
nor U6016 (N_6016,N_5991,N_5835);
or U6017 (N_6017,N_5791,N_5689);
xnor U6018 (N_6018,N_5843,N_5782);
and U6019 (N_6019,N_5625,N_5642);
nand U6020 (N_6020,N_5802,N_5931);
nor U6021 (N_6021,N_5855,N_5529);
nand U6022 (N_6022,N_5618,N_5761);
or U6023 (N_6023,N_5614,N_5899);
or U6024 (N_6024,N_5944,N_5867);
and U6025 (N_6025,N_5640,N_5940);
nor U6026 (N_6026,N_5901,N_5883);
or U6027 (N_6027,N_5764,N_5787);
nor U6028 (N_6028,N_5669,N_5657);
nor U6029 (N_6029,N_5846,N_5792);
nor U6030 (N_6030,N_5954,N_5795);
nor U6031 (N_6031,N_5875,N_5805);
nand U6032 (N_6032,N_5896,N_5863);
or U6033 (N_6033,N_5918,N_5832);
nor U6034 (N_6034,N_5985,N_5654);
and U6035 (N_6035,N_5544,N_5912);
or U6036 (N_6036,N_5868,N_5793);
nand U6037 (N_6037,N_5874,N_5520);
and U6038 (N_6038,N_5962,N_5968);
or U6039 (N_6039,N_5756,N_5553);
nand U6040 (N_6040,N_5610,N_5938);
or U6041 (N_6041,N_5927,N_5722);
nand U6042 (N_6042,N_5757,N_5684);
and U6043 (N_6043,N_5528,N_5691);
and U6044 (N_6044,N_5507,N_5545);
nand U6045 (N_6045,N_5973,N_5633);
nor U6046 (N_6046,N_5934,N_5646);
nor U6047 (N_6047,N_5649,N_5884);
xor U6048 (N_6048,N_5799,N_5981);
nand U6049 (N_6049,N_5905,N_5502);
nand U6050 (N_6050,N_5930,N_5683);
nand U6051 (N_6051,N_5915,N_5916);
nand U6052 (N_6052,N_5759,N_5650);
nor U6053 (N_6053,N_5810,N_5564);
and U6054 (N_6054,N_5549,N_5837);
nand U6055 (N_6055,N_5754,N_5775);
nor U6056 (N_6056,N_5721,N_5589);
and U6057 (N_6057,N_5869,N_5917);
and U6058 (N_6058,N_5733,N_5630);
nor U6059 (N_6059,N_5676,N_5537);
nor U6060 (N_6060,N_5623,N_5508);
nand U6061 (N_6061,N_5853,N_5577);
nand U6062 (N_6062,N_5840,N_5975);
nand U6063 (N_6063,N_5786,N_5804);
and U6064 (N_6064,N_5612,N_5609);
nand U6065 (N_6065,N_5734,N_5711);
and U6066 (N_6066,N_5989,N_5878);
nand U6067 (N_6067,N_5737,N_5700);
nor U6068 (N_6068,N_5741,N_5638);
nand U6069 (N_6069,N_5750,N_5513);
xnor U6070 (N_6070,N_5966,N_5562);
nor U6071 (N_6071,N_5800,N_5946);
or U6072 (N_6072,N_5813,N_5748);
nand U6073 (N_6073,N_5635,N_5821);
and U6074 (N_6074,N_5871,N_5616);
or U6075 (N_6075,N_5746,N_5725);
xnor U6076 (N_6076,N_5602,N_5988);
or U6077 (N_6077,N_5718,N_5941);
or U6078 (N_6078,N_5955,N_5661);
xnor U6079 (N_6079,N_5866,N_5824);
nor U6080 (N_6080,N_5844,N_5913);
nor U6081 (N_6081,N_5847,N_5951);
or U6082 (N_6082,N_5767,N_5557);
nor U6083 (N_6083,N_5876,N_5515);
or U6084 (N_6084,N_5690,N_5849);
or U6085 (N_6085,N_5807,N_5864);
nand U6086 (N_6086,N_5812,N_5703);
and U6087 (N_6087,N_5970,N_5958);
or U6088 (N_6088,N_5829,N_5879);
nand U6089 (N_6089,N_5882,N_5815);
or U6090 (N_6090,N_5816,N_5579);
nand U6091 (N_6091,N_5587,N_5932);
nor U6092 (N_6092,N_5851,N_5527);
nor U6093 (N_6093,N_5662,N_5933);
nor U6094 (N_6094,N_5893,N_5729);
and U6095 (N_6095,N_5588,N_5701);
or U6096 (N_6096,N_5667,N_5987);
nor U6097 (N_6097,N_5891,N_5752);
nand U6098 (N_6098,N_5826,N_5518);
or U6099 (N_6099,N_5862,N_5536);
or U6100 (N_6100,N_5719,N_5809);
xnor U6101 (N_6101,N_5842,N_5573);
nor U6102 (N_6102,N_5914,N_5695);
and U6103 (N_6103,N_5626,N_5776);
or U6104 (N_6104,N_5670,N_5825);
or U6105 (N_6105,N_5600,N_5990);
or U6106 (N_6106,N_5796,N_5762);
and U6107 (N_6107,N_5926,N_5881);
and U6108 (N_6108,N_5584,N_5976);
or U6109 (N_6109,N_5909,N_5993);
nand U6110 (N_6110,N_5890,N_5850);
nor U6111 (N_6111,N_5705,N_5929);
xor U6112 (N_6112,N_5902,N_5861);
or U6113 (N_6113,N_5935,N_5790);
nand U6114 (N_6114,N_5709,N_5925);
or U6115 (N_6115,N_5738,N_5643);
xnor U6116 (N_6116,N_5628,N_5660);
and U6117 (N_6117,N_5509,N_5950);
or U6118 (N_6118,N_5983,N_5677);
xnor U6119 (N_6119,N_5665,N_5525);
nand U6120 (N_6120,N_5583,N_5644);
nand U6121 (N_6121,N_5877,N_5533);
nor U6122 (N_6122,N_5641,N_5679);
or U6123 (N_6123,N_5768,N_5672);
nand U6124 (N_6124,N_5910,N_5598);
or U6125 (N_6125,N_5586,N_5624);
xor U6126 (N_6126,N_5971,N_5828);
nor U6127 (N_6127,N_5595,N_5594);
nor U6128 (N_6128,N_5606,N_5906);
nand U6129 (N_6129,N_5781,N_5561);
nor U6130 (N_6130,N_5702,N_5911);
nand U6131 (N_6131,N_5834,N_5723);
xnor U6132 (N_6132,N_5634,N_5590);
and U6133 (N_6133,N_5994,N_5870);
nand U6134 (N_6134,N_5511,N_5998);
nand U6135 (N_6135,N_5539,N_5637);
and U6136 (N_6136,N_5997,N_5728);
or U6137 (N_6137,N_5698,N_5697);
nor U6138 (N_6138,N_5500,N_5727);
and U6139 (N_6139,N_5585,N_5960);
nand U6140 (N_6140,N_5653,N_5555);
or U6141 (N_6141,N_5845,N_5710);
nor U6142 (N_6142,N_5563,N_5522);
nand U6143 (N_6143,N_5542,N_5622);
or U6144 (N_6144,N_5992,N_5751);
and U6145 (N_6145,N_5922,N_5953);
or U6146 (N_6146,N_5977,N_5655);
and U6147 (N_6147,N_5613,N_5948);
or U6148 (N_6148,N_5924,N_5771);
and U6149 (N_6149,N_5732,N_5720);
and U6150 (N_6150,N_5963,N_5521);
and U6151 (N_6151,N_5666,N_5707);
nor U6152 (N_6152,N_5789,N_5591);
and U6153 (N_6153,N_5856,N_5673);
nand U6154 (N_6154,N_5664,N_5900);
nand U6155 (N_6155,N_5551,N_5716);
nand U6156 (N_6156,N_5560,N_5731);
nand U6157 (N_6157,N_5706,N_5831);
nand U6158 (N_6158,N_5747,N_5540);
nand U6159 (N_6159,N_5601,N_5696);
xor U6160 (N_6160,N_5546,N_5819);
nand U6161 (N_6161,N_5659,N_5801);
nand U6162 (N_6162,N_5514,N_5713);
nor U6163 (N_6163,N_5964,N_5957);
nor U6164 (N_6164,N_5923,N_5686);
or U6165 (N_6165,N_5543,N_5833);
or U6166 (N_6166,N_5999,N_5699);
xor U6167 (N_6167,N_5575,N_5503);
and U6168 (N_6168,N_5569,N_5956);
nand U6169 (N_6169,N_5532,N_5943);
nand U6170 (N_6170,N_5920,N_5603);
xor U6171 (N_6171,N_5694,N_5979);
nand U6172 (N_6172,N_5652,N_5501);
or U6173 (N_6173,N_5505,N_5974);
and U6174 (N_6174,N_5581,N_5766);
or U6175 (N_6175,N_5692,N_5740);
nand U6176 (N_6176,N_5937,N_5744);
nand U6177 (N_6177,N_5648,N_5541);
nor U6178 (N_6178,N_5571,N_5599);
and U6179 (N_6179,N_5784,N_5760);
nand U6180 (N_6180,N_5632,N_5749);
nor U6181 (N_6181,N_5523,N_5919);
nor U6182 (N_6182,N_5671,N_5567);
nand U6183 (N_6183,N_5769,N_5619);
nand U6184 (N_6184,N_5592,N_5811);
nor U6185 (N_6185,N_5739,N_5548);
nor U6186 (N_6186,N_5554,N_5681);
or U6187 (N_6187,N_5693,N_5639);
xnor U6188 (N_6188,N_5651,N_5857);
nand U6189 (N_6189,N_5772,N_5888);
xor U6190 (N_6190,N_5730,N_5903);
and U6191 (N_6191,N_5848,N_5818);
nand U6192 (N_6192,N_5647,N_5656);
or U6193 (N_6193,N_5777,N_5887);
or U6194 (N_6194,N_5794,N_5512);
nor U6195 (N_6195,N_5770,N_5758);
or U6196 (N_6196,N_5880,N_5604);
or U6197 (N_6197,N_5530,N_5617);
or U6198 (N_6198,N_5895,N_5854);
xor U6199 (N_6199,N_5996,N_5827);
nor U6200 (N_6200,N_5531,N_5566);
or U6201 (N_6201,N_5568,N_5552);
xor U6202 (N_6202,N_5830,N_5806);
nor U6203 (N_6203,N_5570,N_5526);
nor U6204 (N_6204,N_5945,N_5745);
or U6205 (N_6205,N_5788,N_5504);
xnor U6206 (N_6206,N_5860,N_5808);
or U6207 (N_6207,N_5517,N_5678);
or U6208 (N_6208,N_5885,N_5726);
xnor U6209 (N_6209,N_5582,N_5822);
or U6210 (N_6210,N_5865,N_5952);
nand U6211 (N_6211,N_5763,N_5814);
nor U6212 (N_6212,N_5785,N_5717);
nor U6213 (N_6213,N_5668,N_5708);
and U6214 (N_6214,N_5838,N_5735);
and U6215 (N_6215,N_5986,N_5506);
or U6216 (N_6216,N_5620,N_5715);
or U6217 (N_6217,N_5980,N_5550);
xnor U6218 (N_6218,N_5836,N_5967);
nand U6219 (N_6219,N_5972,N_5685);
nand U6220 (N_6220,N_5858,N_5820);
xor U6221 (N_6221,N_5898,N_5873);
xnor U6222 (N_6222,N_5894,N_5947);
nor U6223 (N_6223,N_5687,N_5995);
and U6224 (N_6224,N_5674,N_5607);
xor U6225 (N_6225,N_5803,N_5565);
or U6226 (N_6226,N_5743,N_5859);
or U6227 (N_6227,N_5765,N_5682);
nor U6228 (N_6228,N_5959,N_5907);
xor U6229 (N_6229,N_5558,N_5780);
nor U6230 (N_6230,N_5969,N_5755);
xor U6231 (N_6231,N_5712,N_5645);
and U6232 (N_6232,N_5631,N_5797);
and U6233 (N_6233,N_5841,N_5779);
and U6234 (N_6234,N_5942,N_5534);
nand U6235 (N_6235,N_5949,N_5636);
nor U6236 (N_6236,N_5978,N_5852);
nand U6237 (N_6237,N_5936,N_5578);
or U6238 (N_6238,N_5892,N_5982);
xnor U6239 (N_6239,N_5516,N_5961);
xor U6240 (N_6240,N_5510,N_5597);
or U6241 (N_6241,N_5736,N_5904);
or U6242 (N_6242,N_5774,N_5615);
or U6243 (N_6243,N_5939,N_5538);
nor U6244 (N_6244,N_5714,N_5688);
or U6245 (N_6245,N_5778,N_5798);
xnor U6246 (N_6246,N_5556,N_5572);
or U6247 (N_6247,N_5680,N_5908);
or U6248 (N_6248,N_5559,N_5872);
nor U6249 (N_6249,N_5605,N_5663);
and U6250 (N_6250,N_5727,N_5665);
or U6251 (N_6251,N_5737,N_5851);
and U6252 (N_6252,N_5947,N_5969);
nand U6253 (N_6253,N_5559,N_5542);
nand U6254 (N_6254,N_5674,N_5847);
nand U6255 (N_6255,N_5688,N_5744);
nor U6256 (N_6256,N_5690,N_5505);
and U6257 (N_6257,N_5955,N_5732);
nand U6258 (N_6258,N_5896,N_5669);
nor U6259 (N_6259,N_5699,N_5994);
nand U6260 (N_6260,N_5676,N_5878);
nand U6261 (N_6261,N_5904,N_5906);
and U6262 (N_6262,N_5746,N_5597);
and U6263 (N_6263,N_5936,N_5713);
nor U6264 (N_6264,N_5812,N_5808);
xor U6265 (N_6265,N_5904,N_5851);
nand U6266 (N_6266,N_5838,N_5899);
nor U6267 (N_6267,N_5824,N_5881);
nand U6268 (N_6268,N_5541,N_5722);
xor U6269 (N_6269,N_5858,N_5698);
or U6270 (N_6270,N_5930,N_5907);
nor U6271 (N_6271,N_5962,N_5741);
and U6272 (N_6272,N_5630,N_5737);
or U6273 (N_6273,N_5586,N_5659);
xnor U6274 (N_6274,N_5581,N_5886);
or U6275 (N_6275,N_5715,N_5501);
or U6276 (N_6276,N_5698,N_5938);
nor U6277 (N_6277,N_5562,N_5626);
or U6278 (N_6278,N_5613,N_5584);
and U6279 (N_6279,N_5858,N_5999);
or U6280 (N_6280,N_5754,N_5942);
and U6281 (N_6281,N_5614,N_5609);
or U6282 (N_6282,N_5622,N_5767);
and U6283 (N_6283,N_5999,N_5653);
or U6284 (N_6284,N_5840,N_5826);
nand U6285 (N_6285,N_5903,N_5852);
xnor U6286 (N_6286,N_5561,N_5833);
xnor U6287 (N_6287,N_5671,N_5715);
nand U6288 (N_6288,N_5675,N_5827);
nor U6289 (N_6289,N_5657,N_5702);
and U6290 (N_6290,N_5989,N_5848);
or U6291 (N_6291,N_5906,N_5578);
or U6292 (N_6292,N_5951,N_5771);
nor U6293 (N_6293,N_5801,N_5607);
nand U6294 (N_6294,N_5921,N_5996);
xnor U6295 (N_6295,N_5634,N_5586);
nor U6296 (N_6296,N_5891,N_5796);
and U6297 (N_6297,N_5767,N_5792);
xor U6298 (N_6298,N_5723,N_5932);
or U6299 (N_6299,N_5606,N_5874);
nor U6300 (N_6300,N_5924,N_5665);
or U6301 (N_6301,N_5674,N_5718);
xor U6302 (N_6302,N_5555,N_5996);
nor U6303 (N_6303,N_5767,N_5634);
and U6304 (N_6304,N_5792,N_5715);
nor U6305 (N_6305,N_5945,N_5974);
and U6306 (N_6306,N_5564,N_5888);
or U6307 (N_6307,N_5649,N_5743);
nand U6308 (N_6308,N_5639,N_5539);
and U6309 (N_6309,N_5538,N_5581);
nor U6310 (N_6310,N_5848,N_5981);
and U6311 (N_6311,N_5939,N_5897);
nor U6312 (N_6312,N_5502,N_5935);
and U6313 (N_6313,N_5638,N_5836);
nand U6314 (N_6314,N_5883,N_5727);
nand U6315 (N_6315,N_5975,N_5504);
or U6316 (N_6316,N_5585,N_5732);
nor U6317 (N_6317,N_5675,N_5741);
or U6318 (N_6318,N_5990,N_5595);
nand U6319 (N_6319,N_5890,N_5739);
nor U6320 (N_6320,N_5539,N_5922);
xnor U6321 (N_6321,N_5706,N_5745);
and U6322 (N_6322,N_5689,N_5833);
or U6323 (N_6323,N_5810,N_5814);
or U6324 (N_6324,N_5774,N_5544);
nor U6325 (N_6325,N_5782,N_5996);
and U6326 (N_6326,N_5828,N_5599);
xnor U6327 (N_6327,N_5771,N_5860);
or U6328 (N_6328,N_5755,N_5584);
nor U6329 (N_6329,N_5786,N_5724);
and U6330 (N_6330,N_5752,N_5572);
xnor U6331 (N_6331,N_5774,N_5715);
or U6332 (N_6332,N_5997,N_5689);
or U6333 (N_6333,N_5572,N_5730);
and U6334 (N_6334,N_5751,N_5933);
nand U6335 (N_6335,N_5852,N_5771);
nand U6336 (N_6336,N_5535,N_5629);
and U6337 (N_6337,N_5781,N_5503);
nor U6338 (N_6338,N_5573,N_5683);
nand U6339 (N_6339,N_5651,N_5686);
nor U6340 (N_6340,N_5654,N_5548);
or U6341 (N_6341,N_5891,N_5927);
xnor U6342 (N_6342,N_5759,N_5688);
xor U6343 (N_6343,N_5892,N_5572);
and U6344 (N_6344,N_5609,N_5554);
nor U6345 (N_6345,N_5845,N_5996);
xor U6346 (N_6346,N_5553,N_5983);
and U6347 (N_6347,N_5969,N_5560);
and U6348 (N_6348,N_5786,N_5831);
or U6349 (N_6349,N_5514,N_5622);
or U6350 (N_6350,N_5608,N_5522);
or U6351 (N_6351,N_5954,N_5909);
and U6352 (N_6352,N_5957,N_5950);
or U6353 (N_6353,N_5770,N_5820);
or U6354 (N_6354,N_5681,N_5592);
and U6355 (N_6355,N_5594,N_5602);
xor U6356 (N_6356,N_5785,N_5755);
and U6357 (N_6357,N_5713,N_5765);
nand U6358 (N_6358,N_5576,N_5719);
xnor U6359 (N_6359,N_5755,N_5995);
nor U6360 (N_6360,N_5687,N_5879);
or U6361 (N_6361,N_5974,N_5807);
nor U6362 (N_6362,N_5644,N_5591);
or U6363 (N_6363,N_5843,N_5750);
nand U6364 (N_6364,N_5660,N_5754);
xor U6365 (N_6365,N_5645,N_5631);
and U6366 (N_6366,N_5818,N_5968);
xnor U6367 (N_6367,N_5877,N_5922);
nand U6368 (N_6368,N_5639,N_5954);
nor U6369 (N_6369,N_5563,N_5665);
or U6370 (N_6370,N_5870,N_5764);
nor U6371 (N_6371,N_5885,N_5888);
nand U6372 (N_6372,N_5522,N_5515);
xor U6373 (N_6373,N_5651,N_5829);
nor U6374 (N_6374,N_5601,N_5954);
and U6375 (N_6375,N_5869,N_5932);
or U6376 (N_6376,N_5720,N_5664);
xnor U6377 (N_6377,N_5869,N_5940);
nand U6378 (N_6378,N_5859,N_5543);
nand U6379 (N_6379,N_5619,N_5523);
nor U6380 (N_6380,N_5611,N_5736);
and U6381 (N_6381,N_5986,N_5861);
or U6382 (N_6382,N_5571,N_5528);
and U6383 (N_6383,N_5550,N_5898);
nand U6384 (N_6384,N_5744,N_5919);
or U6385 (N_6385,N_5993,N_5964);
nand U6386 (N_6386,N_5565,N_5725);
nor U6387 (N_6387,N_5596,N_5590);
nand U6388 (N_6388,N_5776,N_5878);
nand U6389 (N_6389,N_5506,N_5750);
or U6390 (N_6390,N_5631,N_5657);
nor U6391 (N_6391,N_5570,N_5755);
and U6392 (N_6392,N_5790,N_5776);
xor U6393 (N_6393,N_5755,N_5818);
and U6394 (N_6394,N_5879,N_5645);
or U6395 (N_6395,N_5521,N_5678);
nor U6396 (N_6396,N_5867,N_5571);
and U6397 (N_6397,N_5697,N_5573);
nand U6398 (N_6398,N_5798,N_5508);
or U6399 (N_6399,N_5755,N_5594);
xnor U6400 (N_6400,N_5736,N_5815);
and U6401 (N_6401,N_5874,N_5776);
nand U6402 (N_6402,N_5502,N_5820);
and U6403 (N_6403,N_5547,N_5598);
nand U6404 (N_6404,N_5755,N_5981);
or U6405 (N_6405,N_5792,N_5607);
or U6406 (N_6406,N_5776,N_5592);
or U6407 (N_6407,N_5732,N_5848);
nor U6408 (N_6408,N_5773,N_5972);
and U6409 (N_6409,N_5897,N_5796);
nand U6410 (N_6410,N_5769,N_5617);
or U6411 (N_6411,N_5871,N_5839);
or U6412 (N_6412,N_5780,N_5762);
nand U6413 (N_6413,N_5912,N_5640);
and U6414 (N_6414,N_5827,N_5824);
or U6415 (N_6415,N_5834,N_5900);
nor U6416 (N_6416,N_5819,N_5576);
xnor U6417 (N_6417,N_5714,N_5930);
or U6418 (N_6418,N_5505,N_5876);
nor U6419 (N_6419,N_5704,N_5636);
and U6420 (N_6420,N_5770,N_5859);
and U6421 (N_6421,N_5517,N_5787);
nand U6422 (N_6422,N_5736,N_5972);
nand U6423 (N_6423,N_5907,N_5919);
and U6424 (N_6424,N_5659,N_5664);
and U6425 (N_6425,N_5885,N_5708);
and U6426 (N_6426,N_5858,N_5671);
nand U6427 (N_6427,N_5965,N_5941);
xnor U6428 (N_6428,N_5777,N_5592);
or U6429 (N_6429,N_5771,N_5564);
nand U6430 (N_6430,N_5823,N_5882);
or U6431 (N_6431,N_5903,N_5517);
or U6432 (N_6432,N_5763,N_5517);
or U6433 (N_6433,N_5691,N_5995);
nor U6434 (N_6434,N_5648,N_5989);
and U6435 (N_6435,N_5746,N_5924);
and U6436 (N_6436,N_5841,N_5992);
or U6437 (N_6437,N_5832,N_5913);
nand U6438 (N_6438,N_5623,N_5516);
or U6439 (N_6439,N_5894,N_5678);
or U6440 (N_6440,N_5566,N_5625);
nor U6441 (N_6441,N_5574,N_5871);
and U6442 (N_6442,N_5863,N_5607);
or U6443 (N_6443,N_5923,N_5998);
nor U6444 (N_6444,N_5843,N_5648);
and U6445 (N_6445,N_5974,N_5817);
nor U6446 (N_6446,N_5949,N_5627);
and U6447 (N_6447,N_5631,N_5859);
nand U6448 (N_6448,N_5610,N_5645);
nand U6449 (N_6449,N_5895,N_5583);
xnor U6450 (N_6450,N_5763,N_5783);
nor U6451 (N_6451,N_5641,N_5694);
or U6452 (N_6452,N_5716,N_5642);
xor U6453 (N_6453,N_5647,N_5899);
nor U6454 (N_6454,N_5673,N_5512);
or U6455 (N_6455,N_5825,N_5647);
and U6456 (N_6456,N_5701,N_5657);
and U6457 (N_6457,N_5601,N_5905);
and U6458 (N_6458,N_5557,N_5846);
nand U6459 (N_6459,N_5970,N_5974);
nand U6460 (N_6460,N_5838,N_5959);
nor U6461 (N_6461,N_5642,N_5976);
nand U6462 (N_6462,N_5878,N_5840);
and U6463 (N_6463,N_5644,N_5555);
nand U6464 (N_6464,N_5865,N_5982);
and U6465 (N_6465,N_5928,N_5631);
nand U6466 (N_6466,N_5991,N_5538);
and U6467 (N_6467,N_5849,N_5628);
or U6468 (N_6468,N_5873,N_5772);
xor U6469 (N_6469,N_5876,N_5930);
and U6470 (N_6470,N_5689,N_5901);
xor U6471 (N_6471,N_5830,N_5948);
nor U6472 (N_6472,N_5724,N_5792);
and U6473 (N_6473,N_5640,N_5910);
and U6474 (N_6474,N_5692,N_5578);
nor U6475 (N_6475,N_5506,N_5758);
or U6476 (N_6476,N_5867,N_5994);
or U6477 (N_6477,N_5615,N_5638);
nor U6478 (N_6478,N_5767,N_5625);
nand U6479 (N_6479,N_5596,N_5647);
nor U6480 (N_6480,N_5970,N_5992);
nor U6481 (N_6481,N_5580,N_5549);
nand U6482 (N_6482,N_5871,N_5600);
nor U6483 (N_6483,N_5754,N_5589);
xnor U6484 (N_6484,N_5886,N_5546);
nor U6485 (N_6485,N_5738,N_5886);
xnor U6486 (N_6486,N_5679,N_5653);
and U6487 (N_6487,N_5731,N_5804);
xor U6488 (N_6488,N_5550,N_5764);
xor U6489 (N_6489,N_5862,N_5938);
or U6490 (N_6490,N_5578,N_5865);
nor U6491 (N_6491,N_5548,N_5601);
and U6492 (N_6492,N_5502,N_5830);
and U6493 (N_6493,N_5725,N_5982);
nor U6494 (N_6494,N_5779,N_5820);
nand U6495 (N_6495,N_5705,N_5538);
nor U6496 (N_6496,N_5728,N_5628);
nand U6497 (N_6497,N_5768,N_5854);
and U6498 (N_6498,N_5663,N_5782);
or U6499 (N_6499,N_5863,N_5519);
and U6500 (N_6500,N_6254,N_6205);
and U6501 (N_6501,N_6165,N_6308);
nand U6502 (N_6502,N_6143,N_6261);
nand U6503 (N_6503,N_6303,N_6293);
and U6504 (N_6504,N_6444,N_6184);
or U6505 (N_6505,N_6135,N_6053);
and U6506 (N_6506,N_6074,N_6405);
nand U6507 (N_6507,N_6140,N_6124);
nor U6508 (N_6508,N_6339,N_6100);
nand U6509 (N_6509,N_6017,N_6012);
nand U6510 (N_6510,N_6079,N_6276);
and U6511 (N_6511,N_6183,N_6451);
or U6512 (N_6512,N_6358,N_6332);
nand U6513 (N_6513,N_6433,N_6419);
or U6514 (N_6514,N_6327,N_6044);
nor U6515 (N_6515,N_6016,N_6494);
nor U6516 (N_6516,N_6076,N_6023);
nor U6517 (N_6517,N_6265,N_6066);
nor U6518 (N_6518,N_6243,N_6226);
nor U6519 (N_6519,N_6214,N_6200);
or U6520 (N_6520,N_6031,N_6316);
and U6521 (N_6521,N_6445,N_6310);
or U6522 (N_6522,N_6356,N_6292);
nand U6523 (N_6523,N_6319,N_6375);
nor U6524 (N_6524,N_6467,N_6450);
nand U6525 (N_6525,N_6109,N_6164);
xnor U6526 (N_6526,N_6177,N_6090);
nand U6527 (N_6527,N_6203,N_6370);
nand U6528 (N_6528,N_6378,N_6418);
or U6529 (N_6529,N_6286,N_6487);
and U6530 (N_6530,N_6294,N_6034);
nand U6531 (N_6531,N_6070,N_6238);
nand U6532 (N_6532,N_6134,N_6481);
xor U6533 (N_6533,N_6122,N_6432);
xnor U6534 (N_6534,N_6406,N_6386);
and U6535 (N_6535,N_6448,N_6175);
nand U6536 (N_6536,N_6056,N_6281);
and U6537 (N_6537,N_6251,N_6300);
or U6538 (N_6538,N_6367,N_6366);
nor U6539 (N_6539,N_6010,N_6230);
nor U6540 (N_6540,N_6427,N_6298);
nor U6541 (N_6541,N_6312,N_6402);
nand U6542 (N_6542,N_6289,N_6463);
nand U6543 (N_6543,N_6035,N_6264);
nor U6544 (N_6544,N_6178,N_6244);
and U6545 (N_6545,N_6403,N_6201);
xor U6546 (N_6546,N_6065,N_6197);
or U6547 (N_6547,N_6239,N_6496);
nor U6548 (N_6548,N_6227,N_6499);
and U6549 (N_6549,N_6085,N_6045);
xnor U6550 (N_6550,N_6145,N_6409);
and U6551 (N_6551,N_6020,N_6147);
nor U6552 (N_6552,N_6137,N_6417);
nand U6553 (N_6553,N_6422,N_6221);
or U6554 (N_6554,N_6229,N_6054);
and U6555 (N_6555,N_6340,N_6395);
nor U6556 (N_6556,N_6062,N_6036);
and U6557 (N_6557,N_6260,N_6170);
or U6558 (N_6558,N_6410,N_6118);
nand U6559 (N_6559,N_6058,N_6389);
and U6560 (N_6560,N_6462,N_6470);
xor U6561 (N_6561,N_6159,N_6234);
nand U6562 (N_6562,N_6345,N_6443);
and U6563 (N_6563,N_6133,N_6083);
and U6564 (N_6564,N_6228,N_6192);
xnor U6565 (N_6565,N_6051,N_6088);
nand U6566 (N_6566,N_6005,N_6277);
nand U6567 (N_6567,N_6461,N_6232);
nor U6568 (N_6568,N_6441,N_6262);
or U6569 (N_6569,N_6093,N_6460);
or U6570 (N_6570,N_6105,N_6430);
nand U6571 (N_6571,N_6196,N_6231);
and U6572 (N_6572,N_6362,N_6325);
xor U6573 (N_6573,N_6369,N_6220);
nand U6574 (N_6574,N_6453,N_6007);
nor U6575 (N_6575,N_6314,N_6296);
or U6576 (N_6576,N_6149,N_6364);
nor U6577 (N_6577,N_6104,N_6275);
and U6578 (N_6578,N_6152,N_6163);
xnor U6579 (N_6579,N_6235,N_6299);
nor U6580 (N_6580,N_6471,N_6492);
nand U6581 (N_6581,N_6162,N_6155);
nand U6582 (N_6582,N_6285,N_6048);
nand U6583 (N_6583,N_6157,N_6042);
nand U6584 (N_6584,N_6290,N_6047);
or U6585 (N_6585,N_6334,N_6287);
xnor U6586 (N_6586,N_6028,N_6321);
nor U6587 (N_6587,N_6263,N_6166);
or U6588 (N_6588,N_6429,N_6046);
xor U6589 (N_6589,N_6390,N_6349);
and U6590 (N_6590,N_6361,N_6127);
and U6591 (N_6591,N_6457,N_6101);
nand U6592 (N_6592,N_6039,N_6297);
nand U6593 (N_6593,N_6397,N_6216);
nand U6594 (N_6594,N_6497,N_6439);
nor U6595 (N_6595,N_6156,N_6181);
or U6596 (N_6596,N_6317,N_6411);
and U6597 (N_6597,N_6040,N_6377);
nor U6598 (N_6598,N_6412,N_6438);
nor U6599 (N_6599,N_6218,N_6078);
and U6600 (N_6600,N_6307,N_6211);
xnor U6601 (N_6601,N_6027,N_6456);
nor U6602 (N_6602,N_6237,N_6119);
or U6603 (N_6603,N_6038,N_6338);
nand U6604 (N_6604,N_6486,N_6291);
or U6605 (N_6605,N_6142,N_6015);
and U6606 (N_6606,N_6049,N_6011);
nand U6607 (N_6607,N_6279,N_6102);
or U6608 (N_6608,N_6350,N_6120);
nor U6609 (N_6609,N_6013,N_6274);
xnor U6610 (N_6610,N_6404,N_6014);
nor U6611 (N_6611,N_6153,N_6212);
or U6612 (N_6612,N_6478,N_6075);
nor U6613 (N_6613,N_6380,N_6019);
or U6614 (N_6614,N_6415,N_6283);
nor U6615 (N_6615,N_6252,N_6333);
and U6616 (N_6616,N_6324,N_6139);
nand U6617 (N_6617,N_6222,N_6305);
nand U6618 (N_6618,N_6191,N_6179);
xnor U6619 (N_6619,N_6326,N_6037);
or U6620 (N_6620,N_6344,N_6131);
and U6621 (N_6621,N_6257,N_6396);
xor U6622 (N_6622,N_6382,N_6446);
nand U6623 (N_6623,N_6067,N_6468);
nor U6624 (N_6624,N_6425,N_6442);
or U6625 (N_6625,N_6328,N_6084);
and U6626 (N_6626,N_6117,N_6416);
nand U6627 (N_6627,N_6169,N_6111);
and U6628 (N_6628,N_6107,N_6082);
or U6629 (N_6629,N_6435,N_6190);
xnor U6630 (N_6630,N_6077,N_6158);
and U6631 (N_6631,N_6144,N_6401);
nor U6632 (N_6632,N_6288,N_6272);
nand U6633 (N_6633,N_6346,N_6223);
xnor U6634 (N_6634,N_6173,N_6154);
nand U6635 (N_6635,N_6168,N_6360);
or U6636 (N_6636,N_6474,N_6434);
and U6637 (N_6637,N_6353,N_6110);
nor U6638 (N_6638,N_6204,N_6393);
nor U6639 (N_6639,N_6342,N_6247);
nand U6640 (N_6640,N_6259,N_6391);
nand U6641 (N_6641,N_6304,N_6069);
and U6642 (N_6642,N_6407,N_6186);
xnor U6643 (N_6643,N_6026,N_6225);
and U6644 (N_6644,N_6138,N_6399);
or U6645 (N_6645,N_6302,N_6113);
nand U6646 (N_6646,N_6309,N_6413);
nor U6647 (N_6647,N_6343,N_6213);
or U6648 (N_6648,N_6002,N_6236);
xnor U6649 (N_6649,N_6320,N_6379);
and U6650 (N_6650,N_6482,N_6207);
or U6651 (N_6651,N_6136,N_6387);
and U6652 (N_6652,N_6388,N_6268);
nand U6653 (N_6653,N_6423,N_6357);
xnor U6654 (N_6654,N_6021,N_6215);
nor U6655 (N_6655,N_6171,N_6001);
xor U6656 (N_6656,N_6025,N_6195);
or U6657 (N_6657,N_6055,N_6428);
or U6658 (N_6658,N_6041,N_6485);
nor U6659 (N_6659,N_6484,N_6477);
and U6660 (N_6660,N_6004,N_6267);
and U6661 (N_6661,N_6081,N_6273);
nor U6662 (N_6662,N_6488,N_6099);
or U6663 (N_6663,N_6018,N_6420);
xor U6664 (N_6664,N_6098,N_6359);
or U6665 (N_6665,N_6278,N_6210);
nand U6666 (N_6666,N_6202,N_6176);
and U6667 (N_6667,N_6050,N_6029);
nand U6668 (N_6668,N_6452,N_6003);
nand U6669 (N_6669,N_6491,N_6365);
and U6670 (N_6670,N_6248,N_6282);
and U6671 (N_6671,N_6246,N_6063);
nor U6672 (N_6672,N_6061,N_6189);
xor U6673 (N_6673,N_6006,N_6114);
nand U6674 (N_6674,N_6495,N_6129);
nand U6675 (N_6675,N_6475,N_6187);
and U6676 (N_6676,N_6141,N_6126);
nor U6677 (N_6677,N_6198,N_6455);
nor U6678 (N_6678,N_6096,N_6449);
xnor U6679 (N_6679,N_6458,N_6383);
or U6680 (N_6680,N_6341,N_6008);
or U6681 (N_6681,N_6091,N_6022);
and U6682 (N_6682,N_6271,N_6330);
or U6683 (N_6683,N_6347,N_6414);
nand U6684 (N_6684,N_6266,N_6348);
and U6685 (N_6685,N_6249,N_6431);
and U6686 (N_6686,N_6121,N_6033);
and U6687 (N_6687,N_6241,N_6080);
nand U6688 (N_6688,N_6352,N_6043);
and U6689 (N_6689,N_6489,N_6351);
and U6690 (N_6690,N_6284,N_6060);
or U6691 (N_6691,N_6384,N_6363);
and U6692 (N_6692,N_6424,N_6151);
and U6693 (N_6693,N_6132,N_6466);
or U6694 (N_6694,N_6250,N_6188);
nor U6695 (N_6695,N_6318,N_6024);
nor U6696 (N_6696,N_6150,N_6269);
and U6697 (N_6697,N_6087,N_6112);
xnor U6698 (N_6698,N_6146,N_6180);
xor U6699 (N_6699,N_6465,N_6301);
nand U6700 (N_6700,N_6400,N_6329);
xor U6701 (N_6701,N_6374,N_6454);
and U6702 (N_6702,N_6493,N_6224);
or U6703 (N_6703,N_6064,N_6280);
nand U6704 (N_6704,N_6371,N_6209);
and U6705 (N_6705,N_6240,N_6219);
nand U6706 (N_6706,N_6295,N_6071);
or U6707 (N_6707,N_6167,N_6381);
or U6708 (N_6708,N_6030,N_6483);
and U6709 (N_6709,N_6373,N_6057);
nand U6710 (N_6710,N_6490,N_6476);
nand U6711 (N_6711,N_6459,N_6421);
or U6712 (N_6712,N_6128,N_6354);
or U6713 (N_6713,N_6108,N_6473);
xnor U6714 (N_6714,N_6199,N_6089);
and U6715 (N_6715,N_6336,N_6372);
nand U6716 (N_6716,N_6095,N_6331);
xnor U6717 (N_6717,N_6255,N_6469);
or U6718 (N_6718,N_6052,N_6313);
or U6719 (N_6719,N_6161,N_6009);
or U6720 (N_6720,N_6073,N_6000);
and U6721 (N_6721,N_6032,N_6160);
or U6722 (N_6722,N_6479,N_6174);
nand U6723 (N_6723,N_6480,N_6072);
and U6724 (N_6724,N_6086,N_6472);
nor U6725 (N_6725,N_6306,N_6068);
nor U6726 (N_6726,N_6440,N_6464);
nor U6727 (N_6727,N_6206,N_6185);
nand U6728 (N_6728,N_6245,N_6130);
or U6729 (N_6729,N_6394,N_6172);
nor U6730 (N_6730,N_6368,N_6103);
nor U6731 (N_6731,N_6437,N_6208);
or U6732 (N_6732,N_6355,N_6270);
or U6733 (N_6733,N_6315,N_6094);
and U6734 (N_6734,N_6337,N_6253);
or U6735 (N_6735,N_6125,N_6242);
nand U6736 (N_6736,N_6258,N_6322);
or U6737 (N_6737,N_6092,N_6182);
nor U6738 (N_6738,N_6335,N_6256);
and U6739 (N_6739,N_6392,N_6148);
nand U6740 (N_6740,N_6217,N_6385);
xnor U6741 (N_6741,N_6194,N_6097);
and U6742 (N_6742,N_6408,N_6115);
nor U6743 (N_6743,N_6193,N_6376);
nand U6744 (N_6744,N_6426,N_6436);
nor U6745 (N_6745,N_6116,N_6106);
xnor U6746 (N_6746,N_6323,N_6123);
xnor U6747 (N_6747,N_6059,N_6498);
nand U6748 (N_6748,N_6447,N_6311);
nand U6749 (N_6749,N_6233,N_6398);
nor U6750 (N_6750,N_6160,N_6180);
and U6751 (N_6751,N_6065,N_6346);
and U6752 (N_6752,N_6404,N_6000);
xnor U6753 (N_6753,N_6021,N_6321);
nor U6754 (N_6754,N_6479,N_6035);
and U6755 (N_6755,N_6354,N_6480);
or U6756 (N_6756,N_6410,N_6269);
and U6757 (N_6757,N_6435,N_6038);
or U6758 (N_6758,N_6170,N_6011);
and U6759 (N_6759,N_6375,N_6480);
xnor U6760 (N_6760,N_6026,N_6407);
or U6761 (N_6761,N_6364,N_6152);
nor U6762 (N_6762,N_6159,N_6397);
or U6763 (N_6763,N_6403,N_6239);
xor U6764 (N_6764,N_6478,N_6340);
nand U6765 (N_6765,N_6001,N_6429);
nor U6766 (N_6766,N_6236,N_6021);
nor U6767 (N_6767,N_6201,N_6166);
nor U6768 (N_6768,N_6295,N_6468);
nor U6769 (N_6769,N_6442,N_6182);
nor U6770 (N_6770,N_6073,N_6316);
nor U6771 (N_6771,N_6467,N_6418);
nand U6772 (N_6772,N_6111,N_6206);
nand U6773 (N_6773,N_6409,N_6375);
or U6774 (N_6774,N_6160,N_6087);
or U6775 (N_6775,N_6112,N_6394);
nand U6776 (N_6776,N_6101,N_6032);
and U6777 (N_6777,N_6300,N_6464);
or U6778 (N_6778,N_6005,N_6421);
and U6779 (N_6779,N_6269,N_6407);
nor U6780 (N_6780,N_6208,N_6231);
nand U6781 (N_6781,N_6085,N_6400);
nor U6782 (N_6782,N_6241,N_6483);
xnor U6783 (N_6783,N_6348,N_6184);
and U6784 (N_6784,N_6102,N_6422);
or U6785 (N_6785,N_6264,N_6218);
nor U6786 (N_6786,N_6059,N_6057);
and U6787 (N_6787,N_6412,N_6170);
nor U6788 (N_6788,N_6079,N_6142);
and U6789 (N_6789,N_6454,N_6183);
nand U6790 (N_6790,N_6124,N_6028);
nand U6791 (N_6791,N_6399,N_6328);
or U6792 (N_6792,N_6167,N_6054);
or U6793 (N_6793,N_6364,N_6384);
and U6794 (N_6794,N_6479,N_6478);
and U6795 (N_6795,N_6476,N_6087);
and U6796 (N_6796,N_6472,N_6175);
nor U6797 (N_6797,N_6335,N_6093);
and U6798 (N_6798,N_6470,N_6429);
and U6799 (N_6799,N_6388,N_6026);
nor U6800 (N_6800,N_6350,N_6070);
xor U6801 (N_6801,N_6410,N_6035);
nand U6802 (N_6802,N_6130,N_6006);
xor U6803 (N_6803,N_6210,N_6034);
and U6804 (N_6804,N_6380,N_6021);
nand U6805 (N_6805,N_6015,N_6151);
nor U6806 (N_6806,N_6048,N_6142);
and U6807 (N_6807,N_6032,N_6005);
nor U6808 (N_6808,N_6347,N_6078);
nand U6809 (N_6809,N_6288,N_6438);
nor U6810 (N_6810,N_6262,N_6408);
xor U6811 (N_6811,N_6293,N_6026);
and U6812 (N_6812,N_6305,N_6141);
nor U6813 (N_6813,N_6362,N_6403);
nand U6814 (N_6814,N_6333,N_6151);
or U6815 (N_6815,N_6235,N_6113);
nand U6816 (N_6816,N_6154,N_6360);
nand U6817 (N_6817,N_6285,N_6395);
nand U6818 (N_6818,N_6208,N_6227);
or U6819 (N_6819,N_6337,N_6243);
or U6820 (N_6820,N_6450,N_6126);
and U6821 (N_6821,N_6181,N_6302);
and U6822 (N_6822,N_6450,N_6055);
nand U6823 (N_6823,N_6421,N_6461);
xnor U6824 (N_6824,N_6095,N_6027);
xnor U6825 (N_6825,N_6072,N_6313);
xnor U6826 (N_6826,N_6249,N_6433);
and U6827 (N_6827,N_6419,N_6455);
xnor U6828 (N_6828,N_6419,N_6180);
or U6829 (N_6829,N_6028,N_6178);
nand U6830 (N_6830,N_6499,N_6065);
or U6831 (N_6831,N_6051,N_6340);
nand U6832 (N_6832,N_6174,N_6466);
xnor U6833 (N_6833,N_6025,N_6096);
or U6834 (N_6834,N_6326,N_6400);
or U6835 (N_6835,N_6375,N_6188);
nor U6836 (N_6836,N_6226,N_6208);
nand U6837 (N_6837,N_6280,N_6306);
nor U6838 (N_6838,N_6080,N_6387);
and U6839 (N_6839,N_6026,N_6463);
nand U6840 (N_6840,N_6395,N_6308);
nor U6841 (N_6841,N_6360,N_6264);
or U6842 (N_6842,N_6359,N_6145);
or U6843 (N_6843,N_6495,N_6281);
nand U6844 (N_6844,N_6343,N_6079);
nand U6845 (N_6845,N_6190,N_6478);
and U6846 (N_6846,N_6447,N_6349);
nand U6847 (N_6847,N_6444,N_6495);
nand U6848 (N_6848,N_6004,N_6430);
nor U6849 (N_6849,N_6000,N_6072);
or U6850 (N_6850,N_6401,N_6493);
nand U6851 (N_6851,N_6250,N_6114);
or U6852 (N_6852,N_6218,N_6063);
nand U6853 (N_6853,N_6496,N_6340);
nand U6854 (N_6854,N_6032,N_6427);
and U6855 (N_6855,N_6281,N_6130);
or U6856 (N_6856,N_6337,N_6496);
and U6857 (N_6857,N_6362,N_6064);
nand U6858 (N_6858,N_6253,N_6333);
and U6859 (N_6859,N_6263,N_6176);
nand U6860 (N_6860,N_6241,N_6101);
and U6861 (N_6861,N_6107,N_6170);
nor U6862 (N_6862,N_6384,N_6264);
nor U6863 (N_6863,N_6005,N_6384);
nand U6864 (N_6864,N_6045,N_6241);
nand U6865 (N_6865,N_6441,N_6381);
nor U6866 (N_6866,N_6322,N_6199);
or U6867 (N_6867,N_6336,N_6220);
nand U6868 (N_6868,N_6253,N_6497);
nor U6869 (N_6869,N_6090,N_6299);
and U6870 (N_6870,N_6468,N_6385);
or U6871 (N_6871,N_6348,N_6186);
xnor U6872 (N_6872,N_6156,N_6211);
nand U6873 (N_6873,N_6436,N_6432);
nand U6874 (N_6874,N_6323,N_6442);
nor U6875 (N_6875,N_6062,N_6042);
nand U6876 (N_6876,N_6077,N_6207);
nor U6877 (N_6877,N_6366,N_6190);
and U6878 (N_6878,N_6000,N_6262);
xnor U6879 (N_6879,N_6100,N_6379);
or U6880 (N_6880,N_6448,N_6478);
or U6881 (N_6881,N_6162,N_6097);
or U6882 (N_6882,N_6048,N_6368);
or U6883 (N_6883,N_6408,N_6388);
and U6884 (N_6884,N_6215,N_6467);
and U6885 (N_6885,N_6318,N_6184);
or U6886 (N_6886,N_6305,N_6456);
xnor U6887 (N_6887,N_6051,N_6390);
and U6888 (N_6888,N_6070,N_6427);
and U6889 (N_6889,N_6350,N_6048);
xor U6890 (N_6890,N_6477,N_6330);
nor U6891 (N_6891,N_6244,N_6051);
xnor U6892 (N_6892,N_6337,N_6289);
nor U6893 (N_6893,N_6021,N_6292);
nor U6894 (N_6894,N_6097,N_6051);
nor U6895 (N_6895,N_6157,N_6451);
nor U6896 (N_6896,N_6255,N_6472);
xor U6897 (N_6897,N_6488,N_6217);
or U6898 (N_6898,N_6393,N_6302);
nand U6899 (N_6899,N_6009,N_6213);
nor U6900 (N_6900,N_6327,N_6340);
and U6901 (N_6901,N_6373,N_6385);
and U6902 (N_6902,N_6353,N_6480);
and U6903 (N_6903,N_6275,N_6117);
or U6904 (N_6904,N_6450,N_6412);
nor U6905 (N_6905,N_6310,N_6099);
xnor U6906 (N_6906,N_6184,N_6209);
or U6907 (N_6907,N_6248,N_6389);
and U6908 (N_6908,N_6124,N_6221);
xnor U6909 (N_6909,N_6043,N_6471);
nor U6910 (N_6910,N_6432,N_6370);
nand U6911 (N_6911,N_6277,N_6201);
nor U6912 (N_6912,N_6001,N_6093);
nor U6913 (N_6913,N_6129,N_6103);
and U6914 (N_6914,N_6482,N_6295);
nor U6915 (N_6915,N_6475,N_6004);
nand U6916 (N_6916,N_6471,N_6217);
or U6917 (N_6917,N_6207,N_6258);
nor U6918 (N_6918,N_6110,N_6416);
and U6919 (N_6919,N_6077,N_6176);
and U6920 (N_6920,N_6268,N_6248);
nor U6921 (N_6921,N_6212,N_6288);
nor U6922 (N_6922,N_6377,N_6060);
nand U6923 (N_6923,N_6344,N_6493);
or U6924 (N_6924,N_6144,N_6490);
or U6925 (N_6925,N_6360,N_6237);
and U6926 (N_6926,N_6272,N_6440);
nor U6927 (N_6927,N_6333,N_6363);
xor U6928 (N_6928,N_6226,N_6499);
and U6929 (N_6929,N_6411,N_6145);
or U6930 (N_6930,N_6342,N_6383);
and U6931 (N_6931,N_6434,N_6347);
nand U6932 (N_6932,N_6105,N_6447);
nand U6933 (N_6933,N_6296,N_6143);
or U6934 (N_6934,N_6038,N_6180);
and U6935 (N_6935,N_6222,N_6476);
or U6936 (N_6936,N_6039,N_6078);
xnor U6937 (N_6937,N_6292,N_6351);
nor U6938 (N_6938,N_6017,N_6191);
nand U6939 (N_6939,N_6401,N_6462);
and U6940 (N_6940,N_6058,N_6322);
and U6941 (N_6941,N_6340,N_6468);
nand U6942 (N_6942,N_6317,N_6468);
nor U6943 (N_6943,N_6039,N_6212);
nand U6944 (N_6944,N_6385,N_6202);
nor U6945 (N_6945,N_6188,N_6359);
or U6946 (N_6946,N_6416,N_6333);
nand U6947 (N_6947,N_6406,N_6346);
nor U6948 (N_6948,N_6309,N_6459);
nor U6949 (N_6949,N_6494,N_6438);
or U6950 (N_6950,N_6429,N_6286);
nor U6951 (N_6951,N_6444,N_6430);
nor U6952 (N_6952,N_6252,N_6288);
and U6953 (N_6953,N_6479,N_6397);
nand U6954 (N_6954,N_6333,N_6377);
or U6955 (N_6955,N_6023,N_6154);
nor U6956 (N_6956,N_6099,N_6295);
xnor U6957 (N_6957,N_6337,N_6421);
and U6958 (N_6958,N_6042,N_6459);
or U6959 (N_6959,N_6301,N_6413);
nor U6960 (N_6960,N_6039,N_6337);
and U6961 (N_6961,N_6392,N_6346);
or U6962 (N_6962,N_6399,N_6127);
nand U6963 (N_6963,N_6331,N_6242);
and U6964 (N_6964,N_6121,N_6417);
or U6965 (N_6965,N_6221,N_6149);
and U6966 (N_6966,N_6075,N_6295);
nand U6967 (N_6967,N_6137,N_6394);
nand U6968 (N_6968,N_6093,N_6103);
and U6969 (N_6969,N_6100,N_6034);
nand U6970 (N_6970,N_6144,N_6095);
or U6971 (N_6971,N_6278,N_6445);
and U6972 (N_6972,N_6268,N_6272);
or U6973 (N_6973,N_6216,N_6201);
nand U6974 (N_6974,N_6438,N_6348);
or U6975 (N_6975,N_6164,N_6101);
or U6976 (N_6976,N_6245,N_6324);
and U6977 (N_6977,N_6196,N_6228);
nand U6978 (N_6978,N_6012,N_6185);
and U6979 (N_6979,N_6219,N_6212);
nor U6980 (N_6980,N_6290,N_6014);
xnor U6981 (N_6981,N_6423,N_6325);
or U6982 (N_6982,N_6218,N_6479);
nand U6983 (N_6983,N_6145,N_6213);
nor U6984 (N_6984,N_6409,N_6288);
and U6985 (N_6985,N_6318,N_6396);
xor U6986 (N_6986,N_6212,N_6364);
and U6987 (N_6987,N_6374,N_6287);
nor U6988 (N_6988,N_6242,N_6192);
or U6989 (N_6989,N_6497,N_6215);
nand U6990 (N_6990,N_6433,N_6218);
nor U6991 (N_6991,N_6328,N_6396);
and U6992 (N_6992,N_6380,N_6476);
nand U6993 (N_6993,N_6020,N_6065);
or U6994 (N_6994,N_6134,N_6086);
and U6995 (N_6995,N_6022,N_6048);
nor U6996 (N_6996,N_6133,N_6156);
nor U6997 (N_6997,N_6430,N_6200);
or U6998 (N_6998,N_6278,N_6176);
and U6999 (N_6999,N_6012,N_6342);
and U7000 (N_7000,N_6889,N_6680);
nor U7001 (N_7001,N_6526,N_6840);
xnor U7002 (N_7002,N_6542,N_6850);
and U7003 (N_7003,N_6654,N_6651);
xor U7004 (N_7004,N_6825,N_6833);
nor U7005 (N_7005,N_6975,N_6997);
xnor U7006 (N_7006,N_6613,N_6964);
and U7007 (N_7007,N_6712,N_6696);
nor U7008 (N_7008,N_6928,N_6940);
xor U7009 (N_7009,N_6871,N_6950);
nor U7010 (N_7010,N_6703,N_6609);
nor U7011 (N_7011,N_6934,N_6784);
and U7012 (N_7012,N_6540,N_6993);
or U7013 (N_7013,N_6633,N_6755);
and U7014 (N_7014,N_6661,N_6734);
nand U7015 (N_7015,N_6990,N_6608);
and U7016 (N_7016,N_6805,N_6679);
or U7017 (N_7017,N_6702,N_6557);
or U7018 (N_7018,N_6709,N_6801);
or U7019 (N_7019,N_6845,N_6626);
or U7020 (N_7020,N_6598,N_6969);
or U7021 (N_7021,N_6830,N_6777);
nand U7022 (N_7022,N_6795,N_6501);
or U7023 (N_7023,N_6583,N_6731);
or U7024 (N_7024,N_6924,N_6819);
nand U7025 (N_7025,N_6506,N_6809);
nor U7026 (N_7026,N_6509,N_6797);
xnor U7027 (N_7027,N_6650,N_6658);
xnor U7028 (N_7028,N_6808,N_6848);
nand U7029 (N_7029,N_6925,N_6725);
or U7030 (N_7030,N_6959,N_6511);
xnor U7031 (N_7031,N_6705,N_6793);
and U7032 (N_7032,N_6656,N_6592);
nor U7033 (N_7033,N_6645,N_6541);
or U7034 (N_7034,N_6896,N_6919);
nor U7035 (N_7035,N_6647,N_6868);
or U7036 (N_7036,N_6977,N_6922);
and U7037 (N_7037,N_6595,N_6707);
nand U7038 (N_7038,N_6728,N_6552);
xnor U7039 (N_7039,N_6691,N_6740);
and U7040 (N_7040,N_6972,N_6682);
nand U7041 (N_7041,N_6527,N_6739);
nand U7042 (N_7042,N_6687,N_6835);
and U7043 (N_7043,N_6756,N_6502);
nand U7044 (N_7044,N_6638,N_6737);
or U7045 (N_7045,N_6779,N_6824);
nand U7046 (N_7046,N_6617,N_6996);
nor U7047 (N_7047,N_6535,N_6718);
xor U7048 (N_7048,N_6674,N_6981);
nand U7049 (N_7049,N_6634,N_6872);
xor U7050 (N_7050,N_6546,N_6876);
or U7051 (N_7051,N_6998,N_6800);
nand U7052 (N_7052,N_6758,N_6841);
nor U7053 (N_7053,N_6565,N_6544);
and U7054 (N_7054,N_6909,N_6512);
or U7055 (N_7055,N_6867,N_6560);
nor U7056 (N_7056,N_6746,N_6986);
xnor U7057 (N_7057,N_6956,N_6937);
nor U7058 (N_7058,N_6521,N_6816);
or U7059 (N_7059,N_6750,N_6607);
and U7060 (N_7060,N_6878,N_6846);
or U7061 (N_7061,N_6792,N_6568);
nor U7062 (N_7062,N_6523,N_6810);
or U7063 (N_7063,N_6615,N_6672);
and U7064 (N_7064,N_6945,N_6515);
or U7065 (N_7065,N_6858,N_6524);
nand U7066 (N_7066,N_6643,N_6500);
nor U7067 (N_7067,N_6605,N_6630);
nor U7068 (N_7068,N_6735,N_6620);
and U7069 (N_7069,N_6891,N_6985);
nand U7070 (N_7070,N_6563,N_6628);
xor U7071 (N_7071,N_6806,N_6843);
nor U7072 (N_7072,N_6721,N_6855);
nor U7073 (N_7073,N_6893,N_6936);
xor U7074 (N_7074,N_6538,N_6839);
and U7075 (N_7075,N_6545,N_6591);
nand U7076 (N_7076,N_6899,N_6914);
nor U7077 (N_7077,N_6549,N_6988);
nand U7078 (N_7078,N_6804,N_6765);
or U7079 (N_7079,N_6791,N_6602);
or U7080 (N_7080,N_6958,N_6917);
nand U7081 (N_7081,N_6743,N_6686);
nand U7082 (N_7082,N_6773,N_6948);
nor U7083 (N_7083,N_6522,N_6790);
or U7084 (N_7084,N_6852,N_6724);
xnor U7085 (N_7085,N_6699,N_6828);
and U7086 (N_7086,N_6769,N_6762);
nand U7087 (N_7087,N_6982,N_6890);
or U7088 (N_7088,N_6796,N_6597);
and U7089 (N_7089,N_6518,N_6955);
nand U7090 (N_7090,N_6688,N_6660);
nand U7091 (N_7091,N_6967,N_6904);
or U7092 (N_7092,N_6717,N_6741);
nand U7093 (N_7093,N_6973,N_6851);
nor U7094 (N_7094,N_6774,N_6822);
and U7095 (N_7095,N_6856,N_6820);
and U7096 (N_7096,N_6865,N_6794);
nand U7097 (N_7097,N_6869,N_6847);
nand U7098 (N_7098,N_6838,N_6564);
xor U7099 (N_7099,N_6579,N_6670);
nand U7100 (N_7100,N_6907,N_6772);
nand U7101 (N_7101,N_6775,N_6749);
nand U7102 (N_7102,N_6788,N_6732);
or U7103 (N_7103,N_6836,N_6926);
or U7104 (N_7104,N_6561,N_6757);
and U7105 (N_7105,N_6652,N_6811);
and U7106 (N_7106,N_6547,N_6786);
nand U7107 (N_7107,N_6970,N_6533);
and U7108 (N_7108,N_6995,N_6516);
xnor U7109 (N_7109,N_6823,N_6752);
nor U7110 (N_7110,N_6920,N_6514);
nand U7111 (N_7111,N_6649,N_6979);
or U7112 (N_7112,N_6723,N_6653);
nand U7113 (N_7113,N_6528,N_6803);
and U7114 (N_7114,N_6625,N_6778);
nand U7115 (N_7115,N_6677,N_6974);
nor U7116 (N_7116,N_6505,N_6763);
nor U7117 (N_7117,N_6873,N_6837);
nand U7118 (N_7118,N_6905,N_6764);
or U7119 (N_7119,N_6954,N_6553);
and U7120 (N_7120,N_6681,N_6957);
nor U7121 (N_7121,N_6994,N_6751);
nor U7122 (N_7122,N_6943,N_6678);
nor U7123 (N_7123,N_6903,N_6578);
nand U7124 (N_7124,N_6644,N_6676);
nand U7125 (N_7125,N_6657,N_6881);
and U7126 (N_7126,N_6636,N_6714);
xnor U7127 (N_7127,N_6713,N_6738);
nor U7128 (N_7128,N_6508,N_6874);
and U7129 (N_7129,N_6548,N_6968);
or U7130 (N_7130,N_6572,N_6612);
nor U7131 (N_7131,N_6554,N_6517);
or U7132 (N_7132,N_6927,N_6567);
or U7133 (N_7133,N_6991,N_6770);
xor U7134 (N_7134,N_6671,N_6556);
and U7135 (N_7135,N_6888,N_6611);
nand U7136 (N_7136,N_6892,N_6621);
nand U7137 (N_7137,N_6923,N_6949);
xor U7138 (N_7138,N_6627,N_6933);
nor U7139 (N_7139,N_6853,N_6733);
or U7140 (N_7140,N_6610,N_6946);
and U7141 (N_7141,N_6711,N_6659);
xnor U7142 (N_7142,N_6722,N_6673);
and U7143 (N_7143,N_6537,N_6675);
nand U7144 (N_7144,N_6503,N_6832);
nor U7145 (N_7145,N_6558,N_6887);
nand U7146 (N_7146,N_6601,N_6866);
nor U7147 (N_7147,N_6551,N_6619);
nand U7148 (N_7148,N_6895,N_6629);
and U7149 (N_7149,N_6827,N_6555);
nand U7150 (N_7150,N_6701,N_6727);
or U7151 (N_7151,N_6963,N_6594);
and U7152 (N_7152,N_6942,N_6759);
nor U7153 (N_7153,N_6886,N_6692);
xnor U7154 (N_7154,N_6776,N_6864);
or U7155 (N_7155,N_6921,N_6894);
and U7156 (N_7156,N_6879,N_6736);
nand U7157 (N_7157,N_6520,N_6513);
or U7158 (N_7158,N_6953,N_6861);
or U7159 (N_7159,N_6562,N_6916);
xnor U7160 (N_7160,N_6664,N_6599);
or U7161 (N_7161,N_6510,N_6531);
and U7162 (N_7162,N_6992,N_6593);
nand U7163 (N_7163,N_6665,N_6589);
or U7164 (N_7164,N_6960,N_6566);
nor U7165 (N_7165,N_6685,N_6813);
nand U7166 (N_7166,N_6821,N_6834);
or U7167 (N_7167,N_6781,N_6815);
nand U7168 (N_7168,N_6559,N_6623);
nand U7169 (N_7169,N_6761,N_6947);
nand U7170 (N_7170,N_6571,N_6951);
nand U7171 (N_7171,N_6704,N_6906);
nand U7172 (N_7172,N_6882,N_6569);
and U7173 (N_7173,N_6596,N_6577);
or U7174 (N_7174,N_6900,N_6600);
nor U7175 (N_7175,N_6965,N_6844);
and U7176 (N_7176,N_6978,N_6639);
or U7177 (N_7177,N_6938,N_6799);
and U7178 (N_7178,N_6880,N_6863);
and U7179 (N_7179,N_6780,N_6663);
and U7180 (N_7180,N_6587,N_6550);
nor U7181 (N_7181,N_6532,N_6668);
xnor U7182 (N_7182,N_6883,N_6507);
nor U7183 (N_7183,N_6989,N_6829);
nor U7184 (N_7184,N_6708,N_6669);
and U7185 (N_7185,N_6729,N_6754);
nand U7186 (N_7186,N_6831,N_6910);
and U7187 (N_7187,N_6902,N_6716);
nand U7188 (N_7188,N_6525,N_6939);
nor U7189 (N_7189,N_6908,N_6935);
nor U7190 (N_7190,N_6530,N_6860);
or U7191 (N_7191,N_6854,N_6573);
or U7192 (N_7192,N_6606,N_6574);
nand U7193 (N_7193,N_6529,N_6585);
nor U7194 (N_7194,N_6697,N_6767);
or U7195 (N_7195,N_6603,N_6966);
or U7196 (N_7196,N_6710,N_6536);
or U7197 (N_7197,N_6582,N_6575);
and U7198 (N_7198,N_6884,N_6826);
nor U7199 (N_7199,N_6849,N_6766);
and U7200 (N_7200,N_6747,N_6918);
or U7201 (N_7201,N_6760,N_6842);
nand U7202 (N_7202,N_6753,N_6616);
or U7203 (N_7203,N_6667,N_6662);
nor U7204 (N_7204,N_6862,N_6980);
or U7205 (N_7205,N_6930,N_6534);
or U7206 (N_7206,N_6877,N_6952);
nand U7207 (N_7207,N_6787,N_6987);
or U7208 (N_7208,N_6962,N_6817);
or U7209 (N_7209,N_6604,N_6932);
xnor U7210 (N_7210,N_6875,N_6912);
nand U7211 (N_7211,N_6745,N_6576);
nand U7212 (N_7212,N_6614,N_6812);
nand U7213 (N_7213,N_6693,N_6539);
and U7214 (N_7214,N_6519,N_6570);
or U7215 (N_7215,N_6655,N_6818);
and U7216 (N_7216,N_6798,N_6807);
nand U7217 (N_7217,N_6637,N_6789);
nor U7218 (N_7218,N_6586,N_6684);
nor U7219 (N_7219,N_6941,N_6929);
and U7220 (N_7220,N_6870,N_6700);
and U7221 (N_7221,N_6983,N_6543);
xor U7222 (N_7222,N_6584,N_6944);
nor U7223 (N_7223,N_6689,N_6976);
nand U7224 (N_7224,N_6690,N_6744);
nor U7225 (N_7225,N_6590,N_6897);
and U7226 (N_7226,N_6785,N_6726);
nor U7227 (N_7227,N_6715,N_6631);
nor U7228 (N_7228,N_6911,N_6504);
nor U7229 (N_7229,N_6641,N_6632);
and U7230 (N_7230,N_6748,N_6694);
xnor U7231 (N_7231,N_6771,N_6984);
nand U7232 (N_7232,N_6719,N_6783);
and U7233 (N_7233,N_6901,N_6720);
and U7234 (N_7234,N_6814,N_6588);
and U7235 (N_7235,N_6885,N_6618);
xnor U7236 (N_7236,N_6706,N_6580);
nor U7237 (N_7237,N_6857,N_6635);
nand U7238 (N_7238,N_6931,N_6802);
and U7239 (N_7239,N_6915,N_6971);
nor U7240 (N_7240,N_6624,N_6648);
and U7241 (N_7241,N_6961,N_6581);
nand U7242 (N_7242,N_6683,N_6695);
or U7243 (N_7243,N_6640,N_6646);
or U7244 (N_7244,N_6768,N_6782);
and U7245 (N_7245,N_6913,N_6999);
and U7246 (N_7246,N_6742,N_6859);
or U7247 (N_7247,N_6622,N_6698);
xor U7248 (N_7248,N_6898,N_6642);
nor U7249 (N_7249,N_6666,N_6730);
or U7250 (N_7250,N_6745,N_6897);
and U7251 (N_7251,N_6961,N_6512);
nand U7252 (N_7252,N_6570,N_6731);
xor U7253 (N_7253,N_6788,N_6782);
nor U7254 (N_7254,N_6752,N_6686);
nor U7255 (N_7255,N_6707,N_6938);
nor U7256 (N_7256,N_6663,N_6947);
nor U7257 (N_7257,N_6966,N_6537);
nor U7258 (N_7258,N_6826,N_6942);
nand U7259 (N_7259,N_6594,N_6637);
xnor U7260 (N_7260,N_6657,N_6587);
nor U7261 (N_7261,N_6991,N_6920);
and U7262 (N_7262,N_6528,N_6745);
nor U7263 (N_7263,N_6966,N_6631);
nor U7264 (N_7264,N_6760,N_6807);
and U7265 (N_7265,N_6897,N_6958);
nor U7266 (N_7266,N_6931,N_6899);
nand U7267 (N_7267,N_6648,N_6642);
nor U7268 (N_7268,N_6711,N_6807);
or U7269 (N_7269,N_6671,N_6929);
nand U7270 (N_7270,N_6551,N_6942);
xnor U7271 (N_7271,N_6595,N_6677);
or U7272 (N_7272,N_6705,N_6692);
nand U7273 (N_7273,N_6677,N_6753);
nor U7274 (N_7274,N_6887,N_6881);
nand U7275 (N_7275,N_6799,N_6914);
or U7276 (N_7276,N_6708,N_6598);
and U7277 (N_7277,N_6910,N_6992);
and U7278 (N_7278,N_6881,N_6962);
and U7279 (N_7279,N_6635,N_6813);
or U7280 (N_7280,N_6800,N_6775);
nand U7281 (N_7281,N_6627,N_6856);
or U7282 (N_7282,N_6640,N_6557);
or U7283 (N_7283,N_6996,N_6598);
nand U7284 (N_7284,N_6997,N_6937);
nand U7285 (N_7285,N_6612,N_6702);
nand U7286 (N_7286,N_6662,N_6527);
and U7287 (N_7287,N_6579,N_6546);
or U7288 (N_7288,N_6652,N_6690);
nand U7289 (N_7289,N_6808,N_6658);
or U7290 (N_7290,N_6782,N_6888);
or U7291 (N_7291,N_6852,N_6735);
nor U7292 (N_7292,N_6560,N_6881);
or U7293 (N_7293,N_6582,N_6651);
or U7294 (N_7294,N_6733,N_6565);
and U7295 (N_7295,N_6746,N_6920);
nand U7296 (N_7296,N_6542,N_6775);
and U7297 (N_7297,N_6681,N_6910);
and U7298 (N_7298,N_6650,N_6680);
nor U7299 (N_7299,N_6909,N_6510);
xnor U7300 (N_7300,N_6698,N_6502);
and U7301 (N_7301,N_6980,N_6563);
nand U7302 (N_7302,N_6934,N_6600);
and U7303 (N_7303,N_6904,N_6878);
or U7304 (N_7304,N_6552,N_6821);
and U7305 (N_7305,N_6817,N_6709);
and U7306 (N_7306,N_6971,N_6980);
nor U7307 (N_7307,N_6623,N_6645);
and U7308 (N_7308,N_6948,N_6755);
nor U7309 (N_7309,N_6538,N_6879);
nor U7310 (N_7310,N_6810,N_6919);
and U7311 (N_7311,N_6922,N_6825);
or U7312 (N_7312,N_6848,N_6633);
xnor U7313 (N_7313,N_6958,N_6989);
nor U7314 (N_7314,N_6713,N_6511);
nor U7315 (N_7315,N_6975,N_6823);
and U7316 (N_7316,N_6731,N_6847);
xnor U7317 (N_7317,N_6503,N_6742);
or U7318 (N_7318,N_6934,N_6868);
or U7319 (N_7319,N_6966,N_6507);
or U7320 (N_7320,N_6824,N_6971);
nor U7321 (N_7321,N_6811,N_6920);
nor U7322 (N_7322,N_6870,N_6817);
and U7323 (N_7323,N_6947,N_6705);
and U7324 (N_7324,N_6874,N_6807);
or U7325 (N_7325,N_6796,N_6647);
xor U7326 (N_7326,N_6822,N_6903);
nand U7327 (N_7327,N_6757,N_6924);
xor U7328 (N_7328,N_6679,N_6895);
and U7329 (N_7329,N_6719,N_6651);
and U7330 (N_7330,N_6843,N_6898);
nand U7331 (N_7331,N_6587,N_6933);
and U7332 (N_7332,N_6869,N_6785);
nand U7333 (N_7333,N_6753,N_6761);
and U7334 (N_7334,N_6906,N_6729);
and U7335 (N_7335,N_6822,N_6509);
xnor U7336 (N_7336,N_6746,N_6963);
nor U7337 (N_7337,N_6647,N_6703);
nand U7338 (N_7338,N_6515,N_6624);
or U7339 (N_7339,N_6543,N_6505);
xor U7340 (N_7340,N_6561,N_6798);
nand U7341 (N_7341,N_6789,N_6523);
or U7342 (N_7342,N_6823,N_6969);
and U7343 (N_7343,N_6798,N_6621);
nor U7344 (N_7344,N_6715,N_6504);
or U7345 (N_7345,N_6824,N_6981);
nor U7346 (N_7346,N_6502,N_6814);
and U7347 (N_7347,N_6636,N_6503);
nand U7348 (N_7348,N_6884,N_6936);
xor U7349 (N_7349,N_6666,N_6927);
nand U7350 (N_7350,N_6628,N_6716);
or U7351 (N_7351,N_6639,N_6575);
xor U7352 (N_7352,N_6654,N_6875);
and U7353 (N_7353,N_6750,N_6873);
or U7354 (N_7354,N_6903,N_6865);
or U7355 (N_7355,N_6572,N_6658);
or U7356 (N_7356,N_6849,N_6753);
nor U7357 (N_7357,N_6874,N_6621);
or U7358 (N_7358,N_6572,N_6751);
or U7359 (N_7359,N_6610,N_6988);
nor U7360 (N_7360,N_6697,N_6595);
nand U7361 (N_7361,N_6851,N_6978);
nor U7362 (N_7362,N_6955,N_6916);
nand U7363 (N_7363,N_6558,N_6859);
nand U7364 (N_7364,N_6777,N_6931);
xor U7365 (N_7365,N_6645,N_6517);
or U7366 (N_7366,N_6600,N_6946);
xor U7367 (N_7367,N_6935,N_6545);
and U7368 (N_7368,N_6637,N_6833);
or U7369 (N_7369,N_6581,N_6630);
nand U7370 (N_7370,N_6546,N_6708);
nand U7371 (N_7371,N_6787,N_6958);
nand U7372 (N_7372,N_6780,N_6626);
xnor U7373 (N_7373,N_6884,N_6960);
or U7374 (N_7374,N_6793,N_6531);
and U7375 (N_7375,N_6504,N_6561);
and U7376 (N_7376,N_6554,N_6547);
or U7377 (N_7377,N_6831,N_6890);
and U7378 (N_7378,N_6580,N_6972);
nor U7379 (N_7379,N_6765,N_6575);
or U7380 (N_7380,N_6611,N_6585);
and U7381 (N_7381,N_6594,N_6850);
or U7382 (N_7382,N_6617,N_6849);
or U7383 (N_7383,N_6585,N_6849);
nand U7384 (N_7384,N_6961,N_6716);
or U7385 (N_7385,N_6845,N_6941);
or U7386 (N_7386,N_6737,N_6995);
nand U7387 (N_7387,N_6927,N_6862);
nor U7388 (N_7388,N_6656,N_6639);
or U7389 (N_7389,N_6622,N_6767);
nor U7390 (N_7390,N_6764,N_6632);
and U7391 (N_7391,N_6681,N_6554);
and U7392 (N_7392,N_6913,N_6502);
nand U7393 (N_7393,N_6841,N_6839);
nand U7394 (N_7394,N_6707,N_6990);
and U7395 (N_7395,N_6971,N_6876);
nor U7396 (N_7396,N_6757,N_6862);
and U7397 (N_7397,N_6505,N_6776);
nor U7398 (N_7398,N_6785,N_6731);
nor U7399 (N_7399,N_6711,N_6650);
and U7400 (N_7400,N_6737,N_6761);
nor U7401 (N_7401,N_6500,N_6607);
nand U7402 (N_7402,N_6911,N_6813);
nand U7403 (N_7403,N_6966,N_6738);
nor U7404 (N_7404,N_6615,N_6871);
xor U7405 (N_7405,N_6932,N_6684);
xnor U7406 (N_7406,N_6791,N_6847);
and U7407 (N_7407,N_6690,N_6903);
nand U7408 (N_7408,N_6975,N_6932);
xor U7409 (N_7409,N_6774,N_6514);
or U7410 (N_7410,N_6508,N_6961);
nand U7411 (N_7411,N_6821,N_6705);
nand U7412 (N_7412,N_6830,N_6658);
nand U7413 (N_7413,N_6981,N_6620);
and U7414 (N_7414,N_6793,N_6715);
and U7415 (N_7415,N_6834,N_6500);
nand U7416 (N_7416,N_6956,N_6687);
nand U7417 (N_7417,N_6958,N_6818);
nor U7418 (N_7418,N_6970,N_6511);
and U7419 (N_7419,N_6999,N_6686);
nand U7420 (N_7420,N_6854,N_6746);
xor U7421 (N_7421,N_6834,N_6981);
nand U7422 (N_7422,N_6846,N_6624);
nor U7423 (N_7423,N_6847,N_6945);
nand U7424 (N_7424,N_6775,N_6902);
xor U7425 (N_7425,N_6771,N_6526);
and U7426 (N_7426,N_6966,N_6888);
and U7427 (N_7427,N_6964,N_6801);
xor U7428 (N_7428,N_6757,N_6686);
and U7429 (N_7429,N_6907,N_6700);
nor U7430 (N_7430,N_6843,N_6522);
nor U7431 (N_7431,N_6589,N_6530);
nand U7432 (N_7432,N_6825,N_6614);
or U7433 (N_7433,N_6569,N_6847);
or U7434 (N_7434,N_6659,N_6640);
nand U7435 (N_7435,N_6673,N_6879);
and U7436 (N_7436,N_6726,N_6695);
nor U7437 (N_7437,N_6535,N_6548);
nand U7438 (N_7438,N_6502,N_6517);
nor U7439 (N_7439,N_6913,N_6622);
or U7440 (N_7440,N_6579,N_6513);
and U7441 (N_7441,N_6544,N_6898);
or U7442 (N_7442,N_6847,N_6755);
nor U7443 (N_7443,N_6510,N_6890);
nand U7444 (N_7444,N_6511,N_6637);
nor U7445 (N_7445,N_6582,N_6906);
or U7446 (N_7446,N_6589,N_6540);
nand U7447 (N_7447,N_6508,N_6824);
and U7448 (N_7448,N_6807,N_6674);
nand U7449 (N_7449,N_6640,N_6853);
nand U7450 (N_7450,N_6882,N_6604);
and U7451 (N_7451,N_6819,N_6913);
and U7452 (N_7452,N_6734,N_6860);
or U7453 (N_7453,N_6970,N_6882);
xor U7454 (N_7454,N_6782,N_6572);
or U7455 (N_7455,N_6819,N_6502);
and U7456 (N_7456,N_6818,N_6716);
nand U7457 (N_7457,N_6960,N_6504);
nand U7458 (N_7458,N_6600,N_6673);
nand U7459 (N_7459,N_6833,N_6966);
nand U7460 (N_7460,N_6972,N_6708);
and U7461 (N_7461,N_6592,N_6574);
nor U7462 (N_7462,N_6675,N_6699);
nand U7463 (N_7463,N_6760,N_6791);
or U7464 (N_7464,N_6813,N_6656);
or U7465 (N_7465,N_6838,N_6732);
xnor U7466 (N_7466,N_6946,N_6683);
or U7467 (N_7467,N_6923,N_6992);
xnor U7468 (N_7468,N_6837,N_6971);
or U7469 (N_7469,N_6931,N_6689);
and U7470 (N_7470,N_6732,N_6985);
and U7471 (N_7471,N_6707,N_6858);
and U7472 (N_7472,N_6928,N_6840);
nor U7473 (N_7473,N_6614,N_6949);
nor U7474 (N_7474,N_6576,N_6752);
or U7475 (N_7475,N_6722,N_6904);
nand U7476 (N_7476,N_6859,N_6969);
nor U7477 (N_7477,N_6595,N_6823);
xnor U7478 (N_7478,N_6607,N_6737);
nor U7479 (N_7479,N_6853,N_6652);
or U7480 (N_7480,N_6826,N_6531);
nor U7481 (N_7481,N_6849,N_6958);
and U7482 (N_7482,N_6959,N_6633);
and U7483 (N_7483,N_6636,N_6702);
nor U7484 (N_7484,N_6945,N_6815);
and U7485 (N_7485,N_6508,N_6725);
nor U7486 (N_7486,N_6768,N_6664);
nand U7487 (N_7487,N_6966,N_6544);
and U7488 (N_7488,N_6717,N_6526);
or U7489 (N_7489,N_6793,N_6848);
nor U7490 (N_7490,N_6849,N_6505);
and U7491 (N_7491,N_6514,N_6869);
nand U7492 (N_7492,N_6673,N_6740);
nor U7493 (N_7493,N_6550,N_6556);
nor U7494 (N_7494,N_6991,N_6968);
nor U7495 (N_7495,N_6832,N_6944);
nor U7496 (N_7496,N_6924,N_6566);
and U7497 (N_7497,N_6787,N_6588);
or U7498 (N_7498,N_6808,N_6636);
nand U7499 (N_7499,N_6899,N_6559);
or U7500 (N_7500,N_7400,N_7487);
nor U7501 (N_7501,N_7468,N_7100);
nor U7502 (N_7502,N_7301,N_7423);
nor U7503 (N_7503,N_7040,N_7257);
nor U7504 (N_7504,N_7348,N_7180);
or U7505 (N_7505,N_7153,N_7323);
and U7506 (N_7506,N_7005,N_7162);
xor U7507 (N_7507,N_7430,N_7288);
nor U7508 (N_7508,N_7366,N_7344);
nor U7509 (N_7509,N_7345,N_7135);
xor U7510 (N_7510,N_7273,N_7491);
or U7511 (N_7511,N_7432,N_7433);
xor U7512 (N_7512,N_7281,N_7374);
nor U7513 (N_7513,N_7058,N_7083);
xor U7514 (N_7514,N_7370,N_7128);
nand U7515 (N_7515,N_7034,N_7462);
nor U7516 (N_7516,N_7316,N_7396);
nor U7517 (N_7517,N_7327,N_7193);
or U7518 (N_7518,N_7269,N_7466);
nand U7519 (N_7519,N_7410,N_7268);
or U7520 (N_7520,N_7174,N_7495);
xor U7521 (N_7521,N_7170,N_7026);
nor U7522 (N_7522,N_7217,N_7156);
and U7523 (N_7523,N_7074,N_7061);
and U7524 (N_7524,N_7096,N_7161);
or U7525 (N_7525,N_7009,N_7132);
nor U7526 (N_7526,N_7299,N_7238);
nor U7527 (N_7527,N_7008,N_7391);
or U7528 (N_7528,N_7032,N_7244);
and U7529 (N_7529,N_7020,N_7151);
and U7530 (N_7530,N_7051,N_7091);
nor U7531 (N_7531,N_7414,N_7191);
and U7532 (N_7532,N_7159,N_7305);
nor U7533 (N_7533,N_7160,N_7110);
nor U7534 (N_7534,N_7263,N_7496);
or U7535 (N_7535,N_7250,N_7176);
nor U7536 (N_7536,N_7480,N_7108);
nand U7537 (N_7537,N_7007,N_7282);
xor U7538 (N_7538,N_7329,N_7489);
xor U7539 (N_7539,N_7200,N_7425);
nor U7540 (N_7540,N_7078,N_7314);
nor U7541 (N_7541,N_7056,N_7066);
nor U7542 (N_7542,N_7278,N_7377);
nand U7543 (N_7543,N_7295,N_7077);
nand U7544 (N_7544,N_7421,N_7006);
or U7545 (N_7545,N_7057,N_7230);
and U7546 (N_7546,N_7279,N_7086);
or U7547 (N_7547,N_7261,N_7267);
nand U7548 (N_7548,N_7118,N_7138);
or U7549 (N_7549,N_7014,N_7319);
or U7550 (N_7550,N_7208,N_7227);
nand U7551 (N_7551,N_7420,N_7039);
nand U7552 (N_7552,N_7052,N_7334);
and U7553 (N_7553,N_7064,N_7140);
and U7554 (N_7554,N_7486,N_7456);
and U7555 (N_7555,N_7399,N_7408);
nor U7556 (N_7556,N_7081,N_7233);
nor U7557 (N_7557,N_7458,N_7497);
and U7558 (N_7558,N_7249,N_7087);
and U7559 (N_7559,N_7405,N_7248);
and U7560 (N_7560,N_7333,N_7098);
nand U7561 (N_7561,N_7048,N_7229);
xnor U7562 (N_7562,N_7145,N_7136);
nand U7563 (N_7563,N_7201,N_7464);
nor U7564 (N_7564,N_7447,N_7380);
nor U7565 (N_7565,N_7041,N_7265);
and U7566 (N_7566,N_7474,N_7188);
and U7567 (N_7567,N_7451,N_7127);
or U7568 (N_7568,N_7050,N_7341);
and U7569 (N_7569,N_7084,N_7463);
or U7570 (N_7570,N_7363,N_7076);
nor U7571 (N_7571,N_7046,N_7452);
and U7572 (N_7572,N_7115,N_7352);
and U7573 (N_7573,N_7179,N_7178);
nor U7574 (N_7574,N_7362,N_7092);
nor U7575 (N_7575,N_7484,N_7166);
or U7576 (N_7576,N_7418,N_7122);
nor U7577 (N_7577,N_7382,N_7429);
nand U7578 (N_7578,N_7417,N_7221);
nand U7579 (N_7579,N_7002,N_7024);
and U7580 (N_7580,N_7394,N_7053);
nor U7581 (N_7581,N_7252,N_7297);
nand U7582 (N_7582,N_7088,N_7449);
and U7583 (N_7583,N_7303,N_7318);
nor U7584 (N_7584,N_7448,N_7321);
xnor U7585 (N_7585,N_7183,N_7389);
nand U7586 (N_7586,N_7371,N_7167);
and U7587 (N_7587,N_7253,N_7171);
nand U7588 (N_7588,N_7182,N_7353);
or U7589 (N_7589,N_7205,N_7476);
or U7590 (N_7590,N_7435,N_7307);
and U7591 (N_7591,N_7398,N_7375);
nor U7592 (N_7592,N_7231,N_7383);
nand U7593 (N_7593,N_7422,N_7367);
nor U7594 (N_7594,N_7120,N_7388);
or U7595 (N_7595,N_7202,N_7472);
nand U7596 (N_7596,N_7356,N_7097);
xor U7597 (N_7597,N_7017,N_7402);
nor U7598 (N_7598,N_7428,N_7241);
and U7599 (N_7599,N_7075,N_7190);
nand U7600 (N_7600,N_7222,N_7450);
nor U7601 (N_7601,N_7337,N_7290);
and U7602 (N_7602,N_7245,N_7335);
or U7603 (N_7603,N_7016,N_7199);
nor U7604 (N_7604,N_7256,N_7492);
and U7605 (N_7605,N_7237,N_7325);
nor U7606 (N_7606,N_7315,N_7226);
and U7607 (N_7607,N_7045,N_7387);
and U7608 (N_7608,N_7234,N_7246);
or U7609 (N_7609,N_7114,N_7471);
or U7610 (N_7610,N_7123,N_7274);
nand U7611 (N_7611,N_7310,N_7047);
or U7612 (N_7612,N_7029,N_7173);
nand U7613 (N_7613,N_7384,N_7073);
nand U7614 (N_7614,N_7266,N_7021);
and U7615 (N_7615,N_7350,N_7102);
or U7616 (N_7616,N_7094,N_7296);
or U7617 (N_7617,N_7089,N_7477);
or U7618 (N_7618,N_7139,N_7194);
and U7619 (N_7619,N_7001,N_7042);
or U7620 (N_7620,N_7072,N_7124);
nor U7621 (N_7621,N_7372,N_7411);
xnor U7622 (N_7622,N_7004,N_7436);
or U7623 (N_7623,N_7393,N_7460);
nand U7624 (N_7624,N_7499,N_7481);
and U7625 (N_7625,N_7444,N_7454);
nor U7626 (N_7626,N_7442,N_7494);
nand U7627 (N_7627,N_7211,N_7258);
or U7628 (N_7628,N_7185,N_7163);
nand U7629 (N_7629,N_7473,N_7206);
or U7630 (N_7630,N_7298,N_7106);
or U7631 (N_7631,N_7158,N_7364);
and U7632 (N_7632,N_7453,N_7232);
and U7633 (N_7633,N_7030,N_7025);
or U7634 (N_7634,N_7311,N_7378);
xnor U7635 (N_7635,N_7457,N_7441);
nor U7636 (N_7636,N_7483,N_7479);
nand U7637 (N_7637,N_7060,N_7272);
and U7638 (N_7638,N_7037,N_7289);
or U7639 (N_7639,N_7031,N_7104);
nor U7640 (N_7640,N_7446,N_7349);
nor U7641 (N_7641,N_7331,N_7216);
and U7642 (N_7642,N_7338,N_7080);
xnor U7643 (N_7643,N_7482,N_7130);
nor U7644 (N_7644,N_7461,N_7359);
nand U7645 (N_7645,N_7079,N_7220);
nor U7646 (N_7646,N_7099,N_7198);
nand U7647 (N_7647,N_7044,N_7152);
or U7648 (N_7648,N_7240,N_7141);
nor U7649 (N_7649,N_7493,N_7129);
nand U7650 (N_7650,N_7413,N_7235);
or U7651 (N_7651,N_7035,N_7023);
and U7652 (N_7652,N_7068,N_7144);
nand U7653 (N_7653,N_7228,N_7390);
xor U7654 (N_7654,N_7459,N_7142);
nand U7655 (N_7655,N_7340,N_7131);
nand U7656 (N_7656,N_7304,N_7117);
or U7657 (N_7657,N_7186,N_7286);
or U7658 (N_7658,N_7470,N_7243);
and U7659 (N_7659,N_7070,N_7109);
and U7660 (N_7660,N_7424,N_7165);
nand U7661 (N_7661,N_7284,N_7093);
or U7662 (N_7662,N_7067,N_7443);
and U7663 (N_7663,N_7415,N_7134);
nand U7664 (N_7664,N_7225,N_7440);
or U7665 (N_7665,N_7369,N_7154);
nand U7666 (N_7666,N_7059,N_7177);
nand U7667 (N_7667,N_7022,N_7426);
nand U7668 (N_7668,N_7342,N_7309);
nor U7669 (N_7669,N_7300,N_7328);
nor U7670 (N_7670,N_7085,N_7105);
or U7671 (N_7671,N_7285,N_7113);
nor U7672 (N_7672,N_7385,N_7197);
xor U7673 (N_7673,N_7090,N_7407);
and U7674 (N_7674,N_7330,N_7065);
or U7675 (N_7675,N_7347,N_7419);
or U7676 (N_7676,N_7003,N_7195);
or U7677 (N_7677,N_7168,N_7416);
or U7678 (N_7678,N_7439,N_7187);
nor U7679 (N_7679,N_7101,N_7033);
and U7680 (N_7680,N_7339,N_7336);
or U7681 (N_7681,N_7346,N_7172);
nand U7682 (N_7682,N_7143,N_7397);
or U7683 (N_7683,N_7287,N_7027);
or U7684 (N_7684,N_7116,N_7062);
and U7685 (N_7685,N_7251,N_7351);
and U7686 (N_7686,N_7326,N_7275);
or U7687 (N_7687,N_7204,N_7445);
and U7688 (N_7688,N_7386,N_7147);
nand U7689 (N_7689,N_7150,N_7488);
xor U7690 (N_7690,N_7189,N_7055);
nand U7691 (N_7691,N_7465,N_7038);
or U7692 (N_7692,N_7054,N_7373);
and U7693 (N_7693,N_7317,N_7207);
and U7694 (N_7694,N_7069,N_7107);
and U7695 (N_7695,N_7467,N_7155);
nor U7696 (N_7696,N_7320,N_7018);
xor U7697 (N_7697,N_7112,N_7121);
nor U7698 (N_7698,N_7438,N_7343);
nor U7699 (N_7699,N_7213,N_7146);
and U7700 (N_7700,N_7175,N_7313);
nand U7701 (N_7701,N_7361,N_7431);
nor U7702 (N_7702,N_7490,N_7149);
nand U7703 (N_7703,N_7291,N_7036);
nand U7704 (N_7704,N_7239,N_7095);
nor U7705 (N_7705,N_7028,N_7126);
nand U7706 (N_7706,N_7071,N_7049);
xor U7707 (N_7707,N_7412,N_7355);
nor U7708 (N_7708,N_7360,N_7395);
nor U7709 (N_7709,N_7437,N_7427);
nor U7710 (N_7710,N_7306,N_7011);
nand U7711 (N_7711,N_7255,N_7485);
nor U7712 (N_7712,N_7434,N_7013);
nor U7713 (N_7713,N_7324,N_7312);
or U7714 (N_7714,N_7498,N_7148);
nand U7715 (N_7715,N_7392,N_7270);
nor U7716 (N_7716,N_7302,N_7403);
xnor U7717 (N_7717,N_7214,N_7264);
nor U7718 (N_7718,N_7276,N_7280);
and U7719 (N_7719,N_7137,N_7010);
nor U7720 (N_7720,N_7219,N_7236);
nand U7721 (N_7721,N_7294,N_7322);
nor U7722 (N_7722,N_7293,N_7376);
and U7723 (N_7723,N_7365,N_7332);
nand U7724 (N_7724,N_7212,N_7455);
nor U7725 (N_7725,N_7223,N_7184);
nand U7726 (N_7726,N_7357,N_7224);
nand U7727 (N_7727,N_7247,N_7203);
and U7728 (N_7728,N_7218,N_7254);
and U7729 (N_7729,N_7379,N_7262);
nor U7730 (N_7730,N_7354,N_7157);
nand U7731 (N_7731,N_7283,N_7242);
and U7732 (N_7732,N_7015,N_7409);
or U7733 (N_7733,N_7196,N_7259);
xor U7734 (N_7734,N_7478,N_7000);
nor U7735 (N_7735,N_7169,N_7475);
or U7736 (N_7736,N_7292,N_7103);
nor U7737 (N_7737,N_7043,N_7063);
and U7738 (N_7738,N_7209,N_7019);
and U7739 (N_7739,N_7210,N_7012);
nand U7740 (N_7740,N_7401,N_7260);
or U7741 (N_7741,N_7181,N_7125);
or U7742 (N_7742,N_7215,N_7271);
nor U7743 (N_7743,N_7119,N_7368);
xnor U7744 (N_7744,N_7192,N_7277);
or U7745 (N_7745,N_7133,N_7404);
nor U7746 (N_7746,N_7381,N_7406);
nand U7747 (N_7747,N_7469,N_7308);
nand U7748 (N_7748,N_7358,N_7111);
or U7749 (N_7749,N_7082,N_7164);
nor U7750 (N_7750,N_7113,N_7027);
nand U7751 (N_7751,N_7195,N_7029);
or U7752 (N_7752,N_7366,N_7243);
nor U7753 (N_7753,N_7158,N_7117);
and U7754 (N_7754,N_7101,N_7462);
and U7755 (N_7755,N_7407,N_7360);
nor U7756 (N_7756,N_7102,N_7181);
and U7757 (N_7757,N_7329,N_7144);
nor U7758 (N_7758,N_7422,N_7112);
and U7759 (N_7759,N_7212,N_7125);
nor U7760 (N_7760,N_7063,N_7399);
nand U7761 (N_7761,N_7034,N_7230);
nand U7762 (N_7762,N_7429,N_7145);
and U7763 (N_7763,N_7483,N_7093);
and U7764 (N_7764,N_7184,N_7072);
nand U7765 (N_7765,N_7495,N_7111);
or U7766 (N_7766,N_7036,N_7283);
or U7767 (N_7767,N_7350,N_7293);
and U7768 (N_7768,N_7337,N_7289);
and U7769 (N_7769,N_7006,N_7084);
and U7770 (N_7770,N_7128,N_7239);
nor U7771 (N_7771,N_7133,N_7161);
nand U7772 (N_7772,N_7203,N_7411);
nand U7773 (N_7773,N_7251,N_7018);
and U7774 (N_7774,N_7284,N_7054);
or U7775 (N_7775,N_7321,N_7311);
xnor U7776 (N_7776,N_7061,N_7041);
or U7777 (N_7777,N_7165,N_7376);
nor U7778 (N_7778,N_7014,N_7104);
nand U7779 (N_7779,N_7361,N_7329);
nor U7780 (N_7780,N_7105,N_7035);
or U7781 (N_7781,N_7173,N_7143);
nand U7782 (N_7782,N_7072,N_7033);
nand U7783 (N_7783,N_7481,N_7293);
or U7784 (N_7784,N_7366,N_7444);
and U7785 (N_7785,N_7049,N_7087);
and U7786 (N_7786,N_7444,N_7062);
xnor U7787 (N_7787,N_7322,N_7481);
or U7788 (N_7788,N_7294,N_7484);
and U7789 (N_7789,N_7184,N_7109);
nor U7790 (N_7790,N_7418,N_7420);
and U7791 (N_7791,N_7460,N_7353);
or U7792 (N_7792,N_7112,N_7326);
nor U7793 (N_7793,N_7177,N_7384);
or U7794 (N_7794,N_7128,N_7495);
and U7795 (N_7795,N_7426,N_7069);
or U7796 (N_7796,N_7372,N_7146);
and U7797 (N_7797,N_7225,N_7489);
and U7798 (N_7798,N_7152,N_7416);
nor U7799 (N_7799,N_7118,N_7150);
or U7800 (N_7800,N_7033,N_7282);
and U7801 (N_7801,N_7275,N_7131);
or U7802 (N_7802,N_7342,N_7159);
nand U7803 (N_7803,N_7487,N_7153);
or U7804 (N_7804,N_7220,N_7067);
or U7805 (N_7805,N_7455,N_7024);
nand U7806 (N_7806,N_7197,N_7042);
nor U7807 (N_7807,N_7344,N_7177);
or U7808 (N_7808,N_7039,N_7321);
xor U7809 (N_7809,N_7243,N_7127);
xnor U7810 (N_7810,N_7058,N_7211);
nand U7811 (N_7811,N_7120,N_7033);
nand U7812 (N_7812,N_7294,N_7109);
and U7813 (N_7813,N_7171,N_7378);
nor U7814 (N_7814,N_7283,N_7237);
nor U7815 (N_7815,N_7405,N_7340);
nand U7816 (N_7816,N_7202,N_7283);
or U7817 (N_7817,N_7350,N_7035);
or U7818 (N_7818,N_7074,N_7496);
and U7819 (N_7819,N_7352,N_7062);
and U7820 (N_7820,N_7315,N_7065);
nand U7821 (N_7821,N_7485,N_7035);
xnor U7822 (N_7822,N_7031,N_7478);
nand U7823 (N_7823,N_7449,N_7139);
and U7824 (N_7824,N_7020,N_7492);
xnor U7825 (N_7825,N_7400,N_7360);
xnor U7826 (N_7826,N_7266,N_7250);
nor U7827 (N_7827,N_7377,N_7099);
or U7828 (N_7828,N_7171,N_7239);
and U7829 (N_7829,N_7314,N_7486);
and U7830 (N_7830,N_7295,N_7073);
xnor U7831 (N_7831,N_7036,N_7438);
nor U7832 (N_7832,N_7449,N_7243);
and U7833 (N_7833,N_7444,N_7419);
or U7834 (N_7834,N_7316,N_7223);
or U7835 (N_7835,N_7460,N_7371);
and U7836 (N_7836,N_7067,N_7428);
nand U7837 (N_7837,N_7403,N_7266);
and U7838 (N_7838,N_7183,N_7125);
or U7839 (N_7839,N_7206,N_7400);
nand U7840 (N_7840,N_7057,N_7477);
and U7841 (N_7841,N_7483,N_7113);
nor U7842 (N_7842,N_7014,N_7193);
nor U7843 (N_7843,N_7372,N_7467);
or U7844 (N_7844,N_7380,N_7188);
nand U7845 (N_7845,N_7075,N_7264);
or U7846 (N_7846,N_7253,N_7040);
nor U7847 (N_7847,N_7157,N_7383);
xor U7848 (N_7848,N_7424,N_7107);
or U7849 (N_7849,N_7228,N_7049);
and U7850 (N_7850,N_7439,N_7086);
and U7851 (N_7851,N_7313,N_7090);
nand U7852 (N_7852,N_7297,N_7061);
nor U7853 (N_7853,N_7146,N_7092);
or U7854 (N_7854,N_7240,N_7231);
and U7855 (N_7855,N_7251,N_7167);
and U7856 (N_7856,N_7362,N_7431);
xnor U7857 (N_7857,N_7041,N_7205);
and U7858 (N_7858,N_7398,N_7191);
and U7859 (N_7859,N_7143,N_7246);
and U7860 (N_7860,N_7246,N_7494);
nor U7861 (N_7861,N_7381,N_7228);
nor U7862 (N_7862,N_7170,N_7041);
nand U7863 (N_7863,N_7485,N_7122);
nor U7864 (N_7864,N_7174,N_7381);
and U7865 (N_7865,N_7339,N_7480);
or U7866 (N_7866,N_7425,N_7042);
nor U7867 (N_7867,N_7040,N_7301);
nand U7868 (N_7868,N_7252,N_7260);
nand U7869 (N_7869,N_7080,N_7000);
and U7870 (N_7870,N_7135,N_7348);
nand U7871 (N_7871,N_7179,N_7103);
or U7872 (N_7872,N_7175,N_7189);
nand U7873 (N_7873,N_7347,N_7152);
and U7874 (N_7874,N_7488,N_7231);
or U7875 (N_7875,N_7013,N_7316);
xnor U7876 (N_7876,N_7186,N_7257);
nor U7877 (N_7877,N_7114,N_7105);
xnor U7878 (N_7878,N_7250,N_7033);
nand U7879 (N_7879,N_7228,N_7421);
and U7880 (N_7880,N_7267,N_7334);
or U7881 (N_7881,N_7078,N_7119);
nor U7882 (N_7882,N_7194,N_7208);
and U7883 (N_7883,N_7175,N_7019);
and U7884 (N_7884,N_7465,N_7371);
or U7885 (N_7885,N_7444,N_7039);
or U7886 (N_7886,N_7287,N_7080);
and U7887 (N_7887,N_7390,N_7438);
nand U7888 (N_7888,N_7025,N_7127);
xnor U7889 (N_7889,N_7493,N_7176);
or U7890 (N_7890,N_7020,N_7007);
and U7891 (N_7891,N_7148,N_7313);
nor U7892 (N_7892,N_7404,N_7490);
nor U7893 (N_7893,N_7331,N_7474);
xor U7894 (N_7894,N_7454,N_7118);
or U7895 (N_7895,N_7315,N_7016);
nand U7896 (N_7896,N_7128,N_7117);
or U7897 (N_7897,N_7162,N_7307);
nor U7898 (N_7898,N_7268,N_7216);
or U7899 (N_7899,N_7052,N_7350);
nor U7900 (N_7900,N_7030,N_7231);
nor U7901 (N_7901,N_7284,N_7073);
and U7902 (N_7902,N_7435,N_7441);
nand U7903 (N_7903,N_7054,N_7154);
nand U7904 (N_7904,N_7223,N_7209);
xor U7905 (N_7905,N_7006,N_7217);
nand U7906 (N_7906,N_7466,N_7398);
and U7907 (N_7907,N_7331,N_7014);
nor U7908 (N_7908,N_7172,N_7027);
or U7909 (N_7909,N_7307,N_7104);
or U7910 (N_7910,N_7375,N_7481);
nand U7911 (N_7911,N_7153,N_7473);
and U7912 (N_7912,N_7349,N_7236);
xnor U7913 (N_7913,N_7266,N_7319);
or U7914 (N_7914,N_7358,N_7333);
and U7915 (N_7915,N_7000,N_7163);
and U7916 (N_7916,N_7006,N_7059);
nand U7917 (N_7917,N_7413,N_7100);
or U7918 (N_7918,N_7477,N_7319);
nand U7919 (N_7919,N_7441,N_7294);
or U7920 (N_7920,N_7344,N_7445);
nor U7921 (N_7921,N_7388,N_7473);
or U7922 (N_7922,N_7467,N_7273);
and U7923 (N_7923,N_7065,N_7139);
and U7924 (N_7924,N_7174,N_7369);
or U7925 (N_7925,N_7259,N_7247);
nor U7926 (N_7926,N_7084,N_7115);
nor U7927 (N_7927,N_7174,N_7000);
and U7928 (N_7928,N_7230,N_7466);
or U7929 (N_7929,N_7402,N_7063);
and U7930 (N_7930,N_7031,N_7279);
nand U7931 (N_7931,N_7426,N_7460);
xnor U7932 (N_7932,N_7359,N_7254);
xor U7933 (N_7933,N_7277,N_7234);
nand U7934 (N_7934,N_7243,N_7241);
nand U7935 (N_7935,N_7435,N_7246);
and U7936 (N_7936,N_7234,N_7402);
nand U7937 (N_7937,N_7183,N_7044);
and U7938 (N_7938,N_7498,N_7240);
nor U7939 (N_7939,N_7444,N_7478);
nor U7940 (N_7940,N_7221,N_7353);
nor U7941 (N_7941,N_7180,N_7450);
and U7942 (N_7942,N_7491,N_7063);
and U7943 (N_7943,N_7265,N_7400);
xor U7944 (N_7944,N_7186,N_7224);
nand U7945 (N_7945,N_7449,N_7126);
nand U7946 (N_7946,N_7396,N_7180);
or U7947 (N_7947,N_7310,N_7420);
or U7948 (N_7948,N_7182,N_7023);
or U7949 (N_7949,N_7481,N_7194);
nor U7950 (N_7950,N_7163,N_7363);
or U7951 (N_7951,N_7041,N_7166);
and U7952 (N_7952,N_7017,N_7386);
nor U7953 (N_7953,N_7338,N_7294);
nor U7954 (N_7954,N_7265,N_7058);
nor U7955 (N_7955,N_7468,N_7483);
or U7956 (N_7956,N_7391,N_7497);
xor U7957 (N_7957,N_7211,N_7022);
nand U7958 (N_7958,N_7218,N_7384);
nor U7959 (N_7959,N_7398,N_7139);
nor U7960 (N_7960,N_7479,N_7275);
and U7961 (N_7961,N_7216,N_7394);
nand U7962 (N_7962,N_7420,N_7250);
xnor U7963 (N_7963,N_7471,N_7075);
or U7964 (N_7964,N_7252,N_7078);
and U7965 (N_7965,N_7300,N_7238);
nand U7966 (N_7966,N_7160,N_7075);
nand U7967 (N_7967,N_7340,N_7180);
and U7968 (N_7968,N_7084,N_7126);
and U7969 (N_7969,N_7361,N_7396);
or U7970 (N_7970,N_7100,N_7205);
and U7971 (N_7971,N_7116,N_7322);
and U7972 (N_7972,N_7496,N_7185);
or U7973 (N_7973,N_7467,N_7375);
nor U7974 (N_7974,N_7088,N_7010);
and U7975 (N_7975,N_7294,N_7036);
or U7976 (N_7976,N_7073,N_7475);
or U7977 (N_7977,N_7293,N_7147);
nand U7978 (N_7978,N_7040,N_7136);
or U7979 (N_7979,N_7069,N_7282);
nor U7980 (N_7980,N_7218,N_7264);
nor U7981 (N_7981,N_7134,N_7284);
or U7982 (N_7982,N_7113,N_7226);
nand U7983 (N_7983,N_7209,N_7104);
and U7984 (N_7984,N_7178,N_7165);
nor U7985 (N_7985,N_7234,N_7041);
and U7986 (N_7986,N_7269,N_7495);
xor U7987 (N_7987,N_7223,N_7214);
and U7988 (N_7988,N_7498,N_7225);
nor U7989 (N_7989,N_7133,N_7490);
nand U7990 (N_7990,N_7086,N_7420);
or U7991 (N_7991,N_7445,N_7212);
xor U7992 (N_7992,N_7162,N_7322);
or U7993 (N_7993,N_7268,N_7447);
nor U7994 (N_7994,N_7479,N_7495);
nand U7995 (N_7995,N_7374,N_7074);
and U7996 (N_7996,N_7216,N_7395);
and U7997 (N_7997,N_7084,N_7300);
nand U7998 (N_7998,N_7013,N_7402);
nor U7999 (N_7999,N_7203,N_7442);
and U8000 (N_8000,N_7620,N_7626);
and U8001 (N_8001,N_7990,N_7945);
nor U8002 (N_8002,N_7769,N_7907);
or U8003 (N_8003,N_7759,N_7851);
and U8004 (N_8004,N_7692,N_7942);
or U8005 (N_8005,N_7522,N_7925);
or U8006 (N_8006,N_7742,N_7997);
nor U8007 (N_8007,N_7686,N_7930);
nor U8008 (N_8008,N_7782,N_7879);
nand U8009 (N_8009,N_7574,N_7526);
or U8010 (N_8010,N_7783,N_7912);
nand U8011 (N_8011,N_7811,N_7806);
or U8012 (N_8012,N_7670,N_7735);
or U8013 (N_8013,N_7656,N_7815);
nand U8014 (N_8014,N_7647,N_7602);
nor U8015 (N_8015,N_7880,N_7689);
nand U8016 (N_8016,N_7871,N_7953);
xor U8017 (N_8017,N_7565,N_7906);
and U8018 (N_8018,N_7531,N_7791);
or U8019 (N_8019,N_7619,N_7798);
nor U8020 (N_8020,N_7521,N_7895);
nand U8021 (N_8021,N_7989,N_7818);
nand U8022 (N_8022,N_7671,N_7969);
and U8023 (N_8023,N_7996,N_7785);
and U8024 (N_8024,N_7911,N_7604);
nor U8025 (N_8025,N_7527,N_7552);
xor U8026 (N_8026,N_7749,N_7714);
or U8027 (N_8027,N_7719,N_7638);
xnor U8028 (N_8028,N_7847,N_7512);
nand U8029 (N_8029,N_7795,N_7748);
nand U8030 (N_8030,N_7956,N_7534);
or U8031 (N_8031,N_7902,N_7754);
and U8032 (N_8032,N_7543,N_7805);
xor U8033 (N_8033,N_7810,N_7863);
nand U8034 (N_8034,N_7849,N_7698);
or U8035 (N_8035,N_7955,N_7684);
xor U8036 (N_8036,N_7781,N_7792);
xor U8037 (N_8037,N_7598,N_7950);
nor U8038 (N_8038,N_7694,N_7509);
nand U8039 (N_8039,N_7649,N_7774);
or U8040 (N_8040,N_7926,N_7572);
or U8041 (N_8041,N_7763,N_7508);
nor U8042 (N_8042,N_7645,N_7533);
and U8043 (N_8043,N_7983,N_7540);
nor U8044 (N_8044,N_7720,N_7903);
or U8045 (N_8045,N_7820,N_7766);
nand U8046 (N_8046,N_7535,N_7998);
or U8047 (N_8047,N_7844,N_7780);
or U8048 (N_8048,N_7741,N_7756);
or U8049 (N_8049,N_7797,N_7938);
nor U8050 (N_8050,N_7885,N_7917);
nand U8051 (N_8051,N_7853,N_7706);
nand U8052 (N_8052,N_7650,N_7519);
and U8053 (N_8053,N_7737,N_7869);
and U8054 (N_8054,N_7923,N_7623);
and U8055 (N_8055,N_7914,N_7693);
or U8056 (N_8056,N_7773,N_7652);
nor U8057 (N_8057,N_7932,N_7663);
nand U8058 (N_8058,N_7659,N_7995);
or U8059 (N_8059,N_7755,N_7948);
or U8060 (N_8060,N_7713,N_7845);
and U8061 (N_8061,N_7726,N_7547);
nand U8062 (N_8062,N_7537,N_7506);
or U8063 (N_8063,N_7965,N_7711);
or U8064 (N_8064,N_7518,N_7555);
nand U8065 (N_8065,N_7517,N_7702);
nor U8066 (N_8066,N_7979,N_7788);
or U8067 (N_8067,N_7787,N_7753);
or U8068 (N_8068,N_7883,N_7984);
nor U8069 (N_8069,N_7916,N_7515);
and U8070 (N_8070,N_7646,N_7899);
and U8071 (N_8071,N_7796,N_7590);
and U8072 (N_8072,N_7553,N_7941);
nand U8073 (N_8073,N_7961,N_7872);
or U8074 (N_8074,N_7633,N_7991);
nor U8075 (N_8075,N_7661,N_7747);
nand U8076 (N_8076,N_7700,N_7894);
or U8077 (N_8077,N_7587,N_7963);
nand U8078 (N_8078,N_7993,N_7776);
and U8079 (N_8079,N_7595,N_7709);
nor U8080 (N_8080,N_7594,N_7858);
nand U8081 (N_8081,N_7743,N_7958);
or U8082 (N_8082,N_7935,N_7688);
nor U8083 (N_8083,N_7727,N_7669);
nor U8084 (N_8084,N_7822,N_7589);
or U8085 (N_8085,N_7823,N_7952);
nor U8086 (N_8086,N_7968,N_7637);
xor U8087 (N_8087,N_7772,N_7978);
nand U8088 (N_8088,N_7761,N_7828);
and U8089 (N_8089,N_7939,N_7736);
nand U8090 (N_8090,N_7551,N_7873);
or U8091 (N_8091,N_7653,N_7651);
or U8092 (N_8092,N_7967,N_7870);
nand U8093 (N_8093,N_7542,N_7501);
nor U8094 (N_8094,N_7954,N_7850);
or U8095 (N_8095,N_7557,N_7562);
or U8096 (N_8096,N_7559,N_7502);
or U8097 (N_8097,N_7840,N_7568);
nor U8098 (N_8098,N_7745,N_7970);
nand U8099 (N_8099,N_7672,N_7944);
nor U8100 (N_8100,N_7615,N_7578);
nor U8101 (N_8101,N_7790,N_7732);
nand U8102 (N_8102,N_7800,N_7634);
and U8103 (N_8103,N_7571,N_7929);
or U8104 (N_8104,N_7994,N_7927);
or U8105 (N_8105,N_7657,N_7541);
nor U8106 (N_8106,N_7641,N_7612);
or U8107 (N_8107,N_7928,N_7708);
and U8108 (N_8108,N_7861,N_7583);
or U8109 (N_8109,N_7617,N_7814);
nor U8110 (N_8110,N_7546,N_7888);
or U8111 (N_8111,N_7528,N_7878);
xor U8112 (N_8112,N_7824,N_7585);
and U8113 (N_8113,N_7549,N_7611);
nor U8114 (N_8114,N_7830,N_7854);
or U8115 (N_8115,N_7908,N_7778);
nor U8116 (N_8116,N_7580,N_7835);
and U8117 (N_8117,N_7524,N_7616);
or U8118 (N_8118,N_7723,N_7831);
nand U8119 (N_8119,N_7740,N_7862);
xor U8120 (N_8120,N_7545,N_7505);
nor U8121 (N_8121,N_7786,N_7881);
nand U8122 (N_8122,N_7951,N_7918);
and U8123 (N_8123,N_7632,N_7975);
and U8124 (N_8124,N_7592,N_7731);
nor U8125 (N_8125,N_7609,N_7627);
or U8126 (N_8126,N_7898,N_7550);
and U8127 (N_8127,N_7974,N_7724);
or U8128 (N_8128,N_7802,N_7893);
xor U8129 (N_8129,N_7725,N_7904);
nor U8130 (N_8130,N_7697,N_7924);
nand U8131 (N_8131,N_7520,N_7721);
nor U8132 (N_8132,N_7621,N_7654);
and U8133 (N_8133,N_7890,N_7564);
nor U8134 (N_8134,N_7674,N_7596);
nand U8135 (N_8135,N_7629,N_7886);
nand U8136 (N_8136,N_7757,N_7920);
and U8137 (N_8137,N_7601,N_7964);
xnor U8138 (N_8138,N_7986,N_7771);
nor U8139 (N_8139,N_7607,N_7793);
nand U8140 (N_8140,N_7630,N_7857);
or U8141 (N_8141,N_7677,N_7576);
nand U8142 (N_8142,N_7662,N_7569);
nor U8143 (N_8143,N_7833,N_7642);
nor U8144 (N_8144,N_7525,N_7856);
nand U8145 (N_8145,N_7507,N_7566);
and U8146 (N_8146,N_7896,N_7685);
nor U8147 (N_8147,N_7503,N_7775);
and U8148 (N_8148,N_7668,N_7675);
nand U8149 (N_8149,N_7848,N_7760);
nand U8150 (N_8150,N_7915,N_7937);
and U8151 (N_8151,N_7710,N_7513);
or U8152 (N_8152,N_7746,N_7809);
nor U8153 (N_8153,N_7514,N_7919);
and U8154 (N_8154,N_7529,N_7744);
nor U8155 (N_8155,N_7789,N_7784);
or U8156 (N_8156,N_7913,N_7843);
nor U8157 (N_8157,N_7538,N_7860);
xor U8158 (N_8158,N_7981,N_7581);
xnor U8159 (N_8159,N_7764,N_7622);
nor U8160 (N_8160,N_7544,N_7768);
nand U8161 (N_8161,N_7874,N_7588);
nand U8162 (N_8162,N_7605,N_7987);
nand U8163 (N_8163,N_7799,N_7728);
or U8164 (N_8164,N_7563,N_7900);
nor U8165 (N_8165,N_7825,N_7722);
or U8166 (N_8166,N_7897,N_7839);
nor U8167 (N_8167,N_7980,N_7703);
and U8168 (N_8168,N_7631,N_7999);
xor U8169 (N_8169,N_7640,N_7584);
or U8170 (N_8170,N_7676,N_7946);
nor U8171 (N_8171,N_7624,N_7976);
and U8172 (N_8172,N_7767,N_7666);
nor U8173 (N_8173,N_7664,N_7852);
nand U8174 (N_8174,N_7794,N_7901);
nand U8175 (N_8175,N_7827,N_7730);
and U8176 (N_8176,N_7931,N_7817);
and U8177 (N_8177,N_7934,N_7838);
or U8178 (N_8178,N_7910,N_7936);
or U8179 (N_8179,N_7921,N_7597);
or U8180 (N_8180,N_7680,N_7865);
nand U8181 (N_8181,N_7579,N_7603);
or U8182 (N_8182,N_7949,N_7705);
nor U8183 (N_8183,N_7988,N_7733);
nor U8184 (N_8184,N_7687,N_7567);
or U8185 (N_8185,N_7864,N_7573);
xor U8186 (N_8186,N_7715,N_7943);
or U8187 (N_8187,N_7884,N_7834);
and U8188 (N_8188,N_7985,N_7972);
and U8189 (N_8189,N_7682,N_7752);
and U8190 (N_8190,N_7973,N_7681);
and U8191 (N_8191,N_7808,N_7570);
xor U8192 (N_8192,N_7679,N_7876);
and U8193 (N_8193,N_7947,N_7739);
nand U8194 (N_8194,N_7867,N_7614);
nor U8195 (N_8195,N_7556,N_7593);
nor U8196 (N_8196,N_7842,N_7777);
nor U8197 (N_8197,N_7716,N_7613);
and U8198 (N_8198,N_7859,N_7765);
nand U8199 (N_8199,N_7807,N_7922);
nor U8200 (N_8200,N_7819,N_7816);
and U8201 (N_8201,N_7586,N_7905);
nand U8202 (N_8202,N_7832,N_7643);
or U8203 (N_8203,N_7868,N_7548);
and U8204 (N_8204,N_7977,N_7889);
or U8205 (N_8205,N_7695,N_7667);
nand U8206 (N_8206,N_7539,N_7575);
nor U8207 (N_8207,N_7909,N_7940);
xor U8208 (N_8208,N_7751,N_7554);
nor U8209 (N_8209,N_7658,N_7636);
or U8210 (N_8210,N_7729,N_7960);
nor U8211 (N_8211,N_7523,N_7891);
and U8212 (N_8212,N_7734,N_7750);
and U8213 (N_8213,N_7826,N_7699);
nand U8214 (N_8214,N_7758,N_7560);
nand U8215 (N_8215,N_7673,N_7655);
and U8216 (N_8216,N_7606,N_7712);
and U8217 (N_8217,N_7691,N_7690);
nor U8218 (N_8218,N_7959,N_7933);
nand U8219 (N_8219,N_7639,N_7882);
nor U8220 (N_8220,N_7628,N_7683);
nor U8221 (N_8221,N_7511,N_7770);
nor U8222 (N_8222,N_7875,N_7846);
and U8223 (N_8223,N_7701,N_7644);
or U8224 (N_8224,N_7813,N_7836);
nor U8225 (N_8225,N_7803,N_7635);
and U8226 (N_8226,N_7801,N_7717);
xnor U8227 (N_8227,N_7610,N_7887);
or U8228 (N_8228,N_7648,N_7618);
or U8229 (N_8229,N_7866,N_7504);
nand U8230 (N_8230,N_7536,N_7696);
and U8231 (N_8231,N_7625,N_7599);
nand U8232 (N_8232,N_7812,N_7665);
and U8233 (N_8233,N_7608,N_7829);
nor U8234 (N_8234,N_7962,N_7821);
nand U8235 (N_8235,N_7561,N_7704);
or U8236 (N_8236,N_7718,N_7971);
nor U8237 (N_8237,N_7707,N_7532);
nor U8238 (N_8238,N_7510,N_7804);
nor U8239 (N_8239,N_7992,N_7855);
nand U8240 (N_8240,N_7966,N_7779);
nor U8241 (N_8241,N_7982,N_7841);
xnor U8242 (N_8242,N_7660,N_7892);
nor U8243 (N_8243,N_7530,N_7600);
or U8244 (N_8244,N_7678,N_7877);
and U8245 (N_8245,N_7582,N_7558);
nor U8246 (N_8246,N_7577,N_7762);
nor U8247 (N_8247,N_7516,N_7957);
nor U8248 (N_8248,N_7591,N_7500);
nor U8249 (N_8249,N_7738,N_7837);
or U8250 (N_8250,N_7746,N_7855);
nor U8251 (N_8251,N_7520,N_7607);
nor U8252 (N_8252,N_7825,N_7779);
or U8253 (N_8253,N_7634,N_7569);
or U8254 (N_8254,N_7603,N_7771);
nor U8255 (N_8255,N_7964,N_7877);
or U8256 (N_8256,N_7831,N_7572);
xor U8257 (N_8257,N_7905,N_7755);
and U8258 (N_8258,N_7987,N_7578);
or U8259 (N_8259,N_7700,N_7840);
and U8260 (N_8260,N_7541,N_7522);
or U8261 (N_8261,N_7520,N_7714);
nor U8262 (N_8262,N_7852,N_7650);
and U8263 (N_8263,N_7525,N_7945);
nand U8264 (N_8264,N_7674,N_7952);
or U8265 (N_8265,N_7828,N_7768);
nor U8266 (N_8266,N_7632,N_7618);
or U8267 (N_8267,N_7933,N_7709);
or U8268 (N_8268,N_7641,N_7871);
and U8269 (N_8269,N_7904,N_7569);
nand U8270 (N_8270,N_7704,N_7947);
and U8271 (N_8271,N_7916,N_7724);
or U8272 (N_8272,N_7967,N_7908);
or U8273 (N_8273,N_7531,N_7512);
nand U8274 (N_8274,N_7749,N_7697);
nand U8275 (N_8275,N_7635,N_7915);
and U8276 (N_8276,N_7617,N_7514);
nand U8277 (N_8277,N_7920,N_7576);
nor U8278 (N_8278,N_7682,N_7713);
or U8279 (N_8279,N_7838,N_7892);
nand U8280 (N_8280,N_7608,N_7525);
nand U8281 (N_8281,N_7844,N_7953);
nand U8282 (N_8282,N_7653,N_7652);
and U8283 (N_8283,N_7768,N_7885);
xnor U8284 (N_8284,N_7608,N_7539);
or U8285 (N_8285,N_7515,N_7935);
and U8286 (N_8286,N_7726,N_7690);
and U8287 (N_8287,N_7766,N_7869);
nand U8288 (N_8288,N_7797,N_7786);
or U8289 (N_8289,N_7526,N_7716);
nand U8290 (N_8290,N_7593,N_7915);
nor U8291 (N_8291,N_7550,N_7690);
and U8292 (N_8292,N_7711,N_7784);
nor U8293 (N_8293,N_7792,N_7501);
nor U8294 (N_8294,N_7507,N_7565);
or U8295 (N_8295,N_7604,N_7908);
and U8296 (N_8296,N_7753,N_7907);
xor U8297 (N_8297,N_7753,N_7836);
or U8298 (N_8298,N_7854,N_7555);
nor U8299 (N_8299,N_7665,N_7579);
and U8300 (N_8300,N_7976,N_7814);
or U8301 (N_8301,N_7531,N_7566);
nor U8302 (N_8302,N_7898,N_7837);
nand U8303 (N_8303,N_7886,N_7585);
nor U8304 (N_8304,N_7546,N_7952);
or U8305 (N_8305,N_7767,N_7705);
and U8306 (N_8306,N_7893,N_7944);
or U8307 (N_8307,N_7807,N_7654);
or U8308 (N_8308,N_7969,N_7516);
or U8309 (N_8309,N_7705,N_7926);
or U8310 (N_8310,N_7894,N_7720);
and U8311 (N_8311,N_7897,N_7572);
nand U8312 (N_8312,N_7677,N_7738);
nand U8313 (N_8313,N_7789,N_7567);
and U8314 (N_8314,N_7799,N_7714);
and U8315 (N_8315,N_7778,N_7983);
nand U8316 (N_8316,N_7926,N_7821);
or U8317 (N_8317,N_7582,N_7918);
nand U8318 (N_8318,N_7943,N_7743);
xnor U8319 (N_8319,N_7879,N_7956);
nor U8320 (N_8320,N_7923,N_7585);
nor U8321 (N_8321,N_7581,N_7829);
and U8322 (N_8322,N_7917,N_7975);
nor U8323 (N_8323,N_7955,N_7674);
and U8324 (N_8324,N_7974,N_7609);
nand U8325 (N_8325,N_7976,N_7984);
nor U8326 (N_8326,N_7575,N_7948);
nor U8327 (N_8327,N_7796,N_7735);
nand U8328 (N_8328,N_7924,N_7597);
nand U8329 (N_8329,N_7753,N_7567);
or U8330 (N_8330,N_7754,N_7791);
xnor U8331 (N_8331,N_7926,N_7925);
and U8332 (N_8332,N_7805,N_7995);
and U8333 (N_8333,N_7764,N_7765);
or U8334 (N_8334,N_7615,N_7648);
and U8335 (N_8335,N_7635,N_7660);
nand U8336 (N_8336,N_7760,N_7833);
and U8337 (N_8337,N_7535,N_7906);
nor U8338 (N_8338,N_7566,N_7760);
nand U8339 (N_8339,N_7808,N_7538);
or U8340 (N_8340,N_7540,N_7612);
nor U8341 (N_8341,N_7646,N_7750);
or U8342 (N_8342,N_7688,N_7729);
or U8343 (N_8343,N_7960,N_7788);
nand U8344 (N_8344,N_7567,N_7805);
xnor U8345 (N_8345,N_7527,N_7898);
nand U8346 (N_8346,N_7692,N_7669);
nor U8347 (N_8347,N_7825,N_7856);
nor U8348 (N_8348,N_7856,N_7513);
nand U8349 (N_8349,N_7693,N_7521);
nor U8350 (N_8350,N_7854,N_7704);
or U8351 (N_8351,N_7682,N_7657);
nand U8352 (N_8352,N_7728,N_7735);
nor U8353 (N_8353,N_7789,N_7671);
nand U8354 (N_8354,N_7901,N_7786);
nor U8355 (N_8355,N_7752,N_7676);
nor U8356 (N_8356,N_7560,N_7890);
nand U8357 (N_8357,N_7620,N_7628);
xnor U8358 (N_8358,N_7933,N_7828);
or U8359 (N_8359,N_7557,N_7609);
and U8360 (N_8360,N_7634,N_7681);
and U8361 (N_8361,N_7637,N_7642);
nand U8362 (N_8362,N_7711,N_7962);
xor U8363 (N_8363,N_7860,N_7905);
or U8364 (N_8364,N_7747,N_7603);
nor U8365 (N_8365,N_7519,N_7861);
nand U8366 (N_8366,N_7734,N_7738);
or U8367 (N_8367,N_7515,N_7512);
nor U8368 (N_8368,N_7743,N_7767);
nor U8369 (N_8369,N_7891,N_7996);
nor U8370 (N_8370,N_7665,N_7521);
and U8371 (N_8371,N_7632,N_7516);
or U8372 (N_8372,N_7886,N_7759);
nor U8373 (N_8373,N_7683,N_7697);
and U8374 (N_8374,N_7699,N_7964);
nor U8375 (N_8375,N_7688,N_7925);
or U8376 (N_8376,N_7540,N_7899);
xnor U8377 (N_8377,N_7797,N_7810);
or U8378 (N_8378,N_7724,N_7731);
and U8379 (N_8379,N_7804,N_7912);
or U8380 (N_8380,N_7584,N_7926);
nor U8381 (N_8381,N_7797,N_7694);
nand U8382 (N_8382,N_7719,N_7502);
and U8383 (N_8383,N_7682,N_7675);
and U8384 (N_8384,N_7887,N_7906);
nor U8385 (N_8385,N_7993,N_7921);
and U8386 (N_8386,N_7886,N_7557);
nand U8387 (N_8387,N_7645,N_7785);
nand U8388 (N_8388,N_7664,N_7946);
xnor U8389 (N_8389,N_7821,N_7537);
or U8390 (N_8390,N_7589,N_7514);
nor U8391 (N_8391,N_7844,N_7857);
and U8392 (N_8392,N_7690,N_7637);
xor U8393 (N_8393,N_7520,N_7864);
and U8394 (N_8394,N_7707,N_7546);
and U8395 (N_8395,N_7798,N_7940);
nand U8396 (N_8396,N_7861,N_7603);
nand U8397 (N_8397,N_7922,N_7574);
and U8398 (N_8398,N_7818,N_7972);
and U8399 (N_8399,N_7822,N_7974);
or U8400 (N_8400,N_7979,N_7958);
nor U8401 (N_8401,N_7587,N_7949);
xnor U8402 (N_8402,N_7621,N_7926);
and U8403 (N_8403,N_7792,N_7528);
or U8404 (N_8404,N_7969,N_7884);
nor U8405 (N_8405,N_7601,N_7703);
or U8406 (N_8406,N_7743,N_7812);
nor U8407 (N_8407,N_7559,N_7830);
or U8408 (N_8408,N_7642,N_7661);
or U8409 (N_8409,N_7713,N_7933);
or U8410 (N_8410,N_7795,N_7999);
nand U8411 (N_8411,N_7937,N_7752);
nand U8412 (N_8412,N_7537,N_7540);
xnor U8413 (N_8413,N_7835,N_7582);
and U8414 (N_8414,N_7841,N_7517);
xor U8415 (N_8415,N_7854,N_7551);
and U8416 (N_8416,N_7909,N_7564);
nor U8417 (N_8417,N_7799,N_7529);
nor U8418 (N_8418,N_7749,N_7842);
xnor U8419 (N_8419,N_7899,N_7661);
nand U8420 (N_8420,N_7551,N_7751);
and U8421 (N_8421,N_7969,N_7838);
nor U8422 (N_8422,N_7550,N_7737);
nand U8423 (N_8423,N_7666,N_7991);
or U8424 (N_8424,N_7941,N_7929);
or U8425 (N_8425,N_7522,N_7841);
xor U8426 (N_8426,N_7859,N_7921);
xor U8427 (N_8427,N_7887,N_7735);
and U8428 (N_8428,N_7957,N_7824);
or U8429 (N_8429,N_7658,N_7976);
and U8430 (N_8430,N_7831,N_7735);
and U8431 (N_8431,N_7766,N_7975);
xor U8432 (N_8432,N_7682,N_7553);
nand U8433 (N_8433,N_7994,N_7670);
xor U8434 (N_8434,N_7604,N_7991);
or U8435 (N_8435,N_7712,N_7721);
nand U8436 (N_8436,N_7565,N_7681);
and U8437 (N_8437,N_7813,N_7555);
or U8438 (N_8438,N_7666,N_7706);
and U8439 (N_8439,N_7954,N_7949);
xnor U8440 (N_8440,N_7616,N_7589);
nand U8441 (N_8441,N_7931,N_7937);
nor U8442 (N_8442,N_7951,N_7966);
and U8443 (N_8443,N_7824,N_7830);
and U8444 (N_8444,N_7586,N_7722);
nor U8445 (N_8445,N_7968,N_7940);
nor U8446 (N_8446,N_7839,N_7657);
nor U8447 (N_8447,N_7996,N_7681);
nand U8448 (N_8448,N_7575,N_7954);
nand U8449 (N_8449,N_7543,N_7798);
nor U8450 (N_8450,N_7970,N_7863);
or U8451 (N_8451,N_7502,N_7577);
or U8452 (N_8452,N_7741,N_7596);
nor U8453 (N_8453,N_7857,N_7562);
nor U8454 (N_8454,N_7890,N_7800);
nand U8455 (N_8455,N_7853,N_7680);
xor U8456 (N_8456,N_7954,N_7573);
nor U8457 (N_8457,N_7817,N_7853);
and U8458 (N_8458,N_7526,N_7957);
and U8459 (N_8459,N_7839,N_7901);
and U8460 (N_8460,N_7630,N_7841);
or U8461 (N_8461,N_7750,N_7542);
nand U8462 (N_8462,N_7663,N_7689);
nor U8463 (N_8463,N_7717,N_7890);
xnor U8464 (N_8464,N_7894,N_7627);
or U8465 (N_8465,N_7939,N_7955);
and U8466 (N_8466,N_7666,N_7677);
nor U8467 (N_8467,N_7844,N_7851);
nor U8468 (N_8468,N_7939,N_7994);
and U8469 (N_8469,N_7662,N_7965);
nor U8470 (N_8470,N_7898,N_7620);
or U8471 (N_8471,N_7904,N_7990);
or U8472 (N_8472,N_7649,N_7599);
or U8473 (N_8473,N_7641,N_7894);
nand U8474 (N_8474,N_7587,N_7999);
and U8475 (N_8475,N_7617,N_7594);
nor U8476 (N_8476,N_7637,N_7522);
and U8477 (N_8477,N_7895,N_7968);
or U8478 (N_8478,N_7702,N_7797);
nor U8479 (N_8479,N_7874,N_7692);
nor U8480 (N_8480,N_7717,N_7837);
nor U8481 (N_8481,N_7509,N_7596);
nand U8482 (N_8482,N_7770,N_7942);
xor U8483 (N_8483,N_7552,N_7662);
and U8484 (N_8484,N_7674,N_7970);
nand U8485 (N_8485,N_7822,N_7718);
or U8486 (N_8486,N_7644,N_7954);
nor U8487 (N_8487,N_7866,N_7542);
and U8488 (N_8488,N_7741,N_7986);
or U8489 (N_8489,N_7843,N_7822);
and U8490 (N_8490,N_7821,N_7628);
nand U8491 (N_8491,N_7906,N_7950);
or U8492 (N_8492,N_7813,N_7958);
and U8493 (N_8493,N_7948,N_7811);
and U8494 (N_8494,N_7578,N_7557);
or U8495 (N_8495,N_7907,N_7954);
or U8496 (N_8496,N_7500,N_7917);
nand U8497 (N_8497,N_7515,N_7966);
xor U8498 (N_8498,N_7961,N_7705);
nand U8499 (N_8499,N_7838,N_7908);
nand U8500 (N_8500,N_8130,N_8477);
or U8501 (N_8501,N_8372,N_8274);
and U8502 (N_8502,N_8175,N_8058);
nor U8503 (N_8503,N_8205,N_8098);
and U8504 (N_8504,N_8296,N_8252);
or U8505 (N_8505,N_8380,N_8177);
nand U8506 (N_8506,N_8286,N_8272);
nand U8507 (N_8507,N_8427,N_8028);
nand U8508 (N_8508,N_8492,N_8407);
nand U8509 (N_8509,N_8401,N_8195);
and U8510 (N_8510,N_8000,N_8324);
nand U8511 (N_8511,N_8390,N_8111);
nand U8512 (N_8512,N_8183,N_8473);
nand U8513 (N_8513,N_8253,N_8135);
and U8514 (N_8514,N_8320,N_8347);
xnor U8515 (N_8515,N_8336,N_8018);
and U8516 (N_8516,N_8365,N_8114);
and U8517 (N_8517,N_8491,N_8227);
xnor U8518 (N_8518,N_8465,N_8331);
xor U8519 (N_8519,N_8271,N_8005);
xnor U8520 (N_8520,N_8303,N_8223);
nor U8521 (N_8521,N_8443,N_8475);
nor U8522 (N_8522,N_8471,N_8126);
or U8523 (N_8523,N_8085,N_8106);
nand U8524 (N_8524,N_8090,N_8360);
nand U8525 (N_8525,N_8363,N_8329);
nor U8526 (N_8526,N_8042,N_8181);
or U8527 (N_8527,N_8458,N_8164);
and U8528 (N_8528,N_8495,N_8453);
nor U8529 (N_8529,N_8484,N_8304);
nand U8530 (N_8530,N_8228,N_8041);
and U8531 (N_8531,N_8062,N_8125);
nor U8532 (N_8532,N_8210,N_8101);
nand U8533 (N_8533,N_8449,N_8354);
or U8534 (N_8534,N_8386,N_8222);
and U8535 (N_8535,N_8261,N_8137);
and U8536 (N_8536,N_8486,N_8464);
nor U8537 (N_8537,N_8439,N_8088);
nand U8538 (N_8538,N_8397,N_8338);
or U8539 (N_8539,N_8207,N_8048);
nor U8540 (N_8540,N_8105,N_8235);
nand U8541 (N_8541,N_8093,N_8309);
or U8542 (N_8542,N_8422,N_8369);
nor U8543 (N_8543,N_8353,N_8379);
and U8544 (N_8544,N_8147,N_8482);
or U8545 (N_8545,N_8382,N_8499);
or U8546 (N_8546,N_8030,N_8411);
nand U8547 (N_8547,N_8202,N_8263);
or U8548 (N_8548,N_8074,N_8172);
and U8549 (N_8549,N_8371,N_8096);
and U8550 (N_8550,N_8166,N_8212);
and U8551 (N_8551,N_8128,N_8036);
and U8552 (N_8552,N_8469,N_8060);
nor U8553 (N_8553,N_8299,N_8346);
and U8554 (N_8554,N_8144,N_8383);
xnor U8555 (N_8555,N_8328,N_8203);
or U8556 (N_8556,N_8468,N_8070);
xor U8557 (N_8557,N_8281,N_8433);
nor U8558 (N_8558,N_8051,N_8257);
and U8559 (N_8559,N_8268,N_8141);
and U8560 (N_8560,N_8340,N_8014);
and U8561 (N_8561,N_8357,N_8410);
and U8562 (N_8562,N_8010,N_8277);
nor U8563 (N_8563,N_8127,N_8426);
xor U8564 (N_8564,N_8457,N_8124);
and U8565 (N_8565,N_8221,N_8109);
nor U8566 (N_8566,N_8092,N_8066);
xor U8567 (N_8567,N_8061,N_8113);
and U8568 (N_8568,N_8364,N_8431);
nor U8569 (N_8569,N_8376,N_8022);
xnor U8570 (N_8570,N_8450,N_8013);
and U8571 (N_8571,N_8091,N_8348);
or U8572 (N_8572,N_8129,N_8053);
nand U8573 (N_8573,N_8032,N_8494);
nand U8574 (N_8574,N_8103,N_8311);
or U8575 (N_8575,N_8319,N_8318);
nand U8576 (N_8576,N_8326,N_8145);
and U8577 (N_8577,N_8199,N_8073);
nand U8578 (N_8578,N_8262,N_8288);
nor U8579 (N_8579,N_8472,N_8171);
or U8580 (N_8580,N_8021,N_8341);
nand U8581 (N_8581,N_8020,N_8287);
and U8582 (N_8582,N_8415,N_8143);
and U8583 (N_8583,N_8370,N_8488);
nand U8584 (N_8584,N_8312,N_8275);
or U8585 (N_8585,N_8094,N_8050);
nand U8586 (N_8586,N_8008,N_8115);
or U8587 (N_8587,N_8442,N_8045);
nand U8588 (N_8588,N_8334,N_8155);
nand U8589 (N_8589,N_8146,N_8280);
or U8590 (N_8590,N_8279,N_8230);
nand U8591 (N_8591,N_8463,N_8149);
nand U8592 (N_8592,N_8081,N_8375);
nor U8593 (N_8593,N_8201,N_8295);
nand U8594 (N_8594,N_8409,N_8385);
or U8595 (N_8595,N_8403,N_8445);
nand U8596 (N_8596,N_8119,N_8231);
nand U8597 (N_8597,N_8241,N_8011);
or U8598 (N_8598,N_8134,N_8063);
xnor U8599 (N_8599,N_8278,N_8264);
nand U8600 (N_8600,N_8158,N_8368);
nor U8601 (N_8601,N_8460,N_8104);
or U8602 (N_8602,N_8327,N_8239);
or U8603 (N_8603,N_8220,N_8388);
and U8604 (N_8604,N_8425,N_8016);
nor U8605 (N_8605,N_8413,N_8417);
nor U8606 (N_8606,N_8497,N_8215);
xor U8607 (N_8607,N_8420,N_8291);
and U8608 (N_8608,N_8029,N_8138);
nand U8609 (N_8609,N_8352,N_8266);
nor U8610 (N_8610,N_8224,N_8232);
nand U8611 (N_8611,N_8455,N_8269);
or U8612 (N_8612,N_8498,N_8121);
xor U8613 (N_8613,N_8219,N_8082);
xor U8614 (N_8614,N_8007,N_8116);
or U8615 (N_8615,N_8440,N_8430);
and U8616 (N_8616,N_8136,N_8034);
and U8617 (N_8617,N_8349,N_8496);
or U8618 (N_8618,N_8321,N_8306);
nor U8619 (N_8619,N_8169,N_8398);
or U8620 (N_8620,N_8255,N_8071);
nor U8621 (N_8621,N_8107,N_8163);
or U8622 (N_8622,N_8024,N_8466);
or U8623 (N_8623,N_8026,N_8132);
xor U8624 (N_8624,N_8399,N_8293);
xnor U8625 (N_8625,N_8389,N_8483);
xor U8626 (N_8626,N_8474,N_8167);
nand U8627 (N_8627,N_8174,N_8402);
nand U8628 (N_8628,N_8194,N_8416);
nor U8629 (N_8629,N_8284,N_8462);
nand U8630 (N_8630,N_8187,N_8151);
or U8631 (N_8631,N_8323,N_8238);
and U8632 (N_8632,N_8226,N_8216);
nand U8633 (N_8633,N_8423,N_8017);
nor U8634 (N_8634,N_8037,N_8078);
nand U8635 (N_8635,N_8178,N_8156);
nor U8636 (N_8636,N_8308,N_8384);
nor U8637 (N_8637,N_8206,N_8432);
and U8638 (N_8638,N_8069,N_8170);
and U8639 (N_8639,N_8451,N_8095);
or U8640 (N_8640,N_8342,N_8461);
nor U8641 (N_8641,N_8487,N_8419);
or U8642 (N_8642,N_8068,N_8214);
or U8643 (N_8643,N_8260,N_8120);
or U8644 (N_8644,N_8438,N_8047);
and U8645 (N_8645,N_8240,N_8448);
and U8646 (N_8646,N_8004,N_8394);
or U8647 (N_8647,N_8002,N_8313);
nor U8648 (N_8648,N_8059,N_8229);
or U8649 (N_8649,N_8396,N_8290);
xnor U8650 (N_8650,N_8191,N_8259);
nand U8651 (N_8651,N_8421,N_8305);
nor U8652 (N_8652,N_8161,N_8412);
nand U8653 (N_8653,N_8332,N_8100);
and U8654 (N_8654,N_8055,N_8429);
nand U8655 (N_8655,N_8193,N_8079);
nor U8656 (N_8656,N_8490,N_8196);
xnor U8657 (N_8657,N_8225,N_8118);
or U8658 (N_8658,N_8454,N_8282);
xor U8659 (N_8659,N_8283,N_8400);
nand U8660 (N_8660,N_8054,N_8441);
nand U8661 (N_8661,N_8197,N_8023);
and U8662 (N_8662,N_8244,N_8168);
or U8663 (N_8663,N_8248,N_8233);
xor U8664 (N_8664,N_8192,N_8250);
or U8665 (N_8665,N_8251,N_8366);
xnor U8666 (N_8666,N_8046,N_8086);
and U8667 (N_8667,N_8148,N_8140);
nor U8668 (N_8668,N_8077,N_8276);
nor U8669 (N_8669,N_8333,N_8133);
and U8670 (N_8670,N_8356,N_8075);
nor U8671 (N_8671,N_8325,N_8456);
or U8672 (N_8672,N_8478,N_8038);
xnor U8673 (N_8673,N_8436,N_8316);
nor U8674 (N_8674,N_8150,N_8344);
or U8675 (N_8675,N_8317,N_8031);
nand U8676 (N_8676,N_8322,N_8083);
or U8677 (N_8677,N_8345,N_8182);
xnor U8678 (N_8678,N_8099,N_8447);
and U8679 (N_8679,N_8337,N_8330);
or U8680 (N_8680,N_8198,N_8246);
nand U8681 (N_8681,N_8476,N_8122);
or U8682 (N_8682,N_8355,N_8392);
xnor U8683 (N_8683,N_8404,N_8395);
and U8684 (N_8684,N_8176,N_8056);
nor U8685 (N_8685,N_8359,N_8006);
xnor U8686 (N_8686,N_8052,N_8185);
xnor U8687 (N_8687,N_8485,N_8373);
nand U8688 (N_8688,N_8097,N_8139);
nor U8689 (N_8689,N_8300,N_8180);
nand U8690 (N_8690,N_8258,N_8159);
and U8691 (N_8691,N_8200,N_8035);
xnor U8692 (N_8692,N_8391,N_8254);
nand U8693 (N_8693,N_8049,N_8160);
nor U8694 (N_8694,N_8102,N_8157);
nor U8695 (N_8695,N_8189,N_8470);
nand U8696 (N_8696,N_8315,N_8184);
nand U8697 (N_8697,N_8064,N_8236);
nand U8698 (N_8698,N_8213,N_8381);
or U8699 (N_8699,N_8285,N_8123);
or U8700 (N_8700,N_8310,N_8080);
nor U8701 (N_8701,N_8003,N_8190);
nor U8702 (N_8702,N_8493,N_8437);
nand U8703 (N_8703,N_8065,N_8173);
nand U8704 (N_8704,N_8218,N_8444);
or U8705 (N_8705,N_8467,N_8406);
nor U8706 (N_8706,N_8408,N_8179);
xnor U8707 (N_8707,N_8076,N_8234);
or U8708 (N_8708,N_8001,N_8188);
xor U8709 (N_8709,N_8084,N_8350);
xnor U8710 (N_8710,N_8245,N_8154);
or U8711 (N_8711,N_8358,N_8162);
and U8712 (N_8712,N_8211,N_8243);
or U8713 (N_8713,N_8459,N_8377);
nand U8714 (N_8714,N_8292,N_8019);
nand U8715 (N_8715,N_8393,N_8237);
nor U8716 (N_8716,N_8405,N_8152);
and U8717 (N_8717,N_8273,N_8387);
nand U8718 (N_8718,N_8367,N_8270);
nand U8719 (N_8719,N_8351,N_8057);
and U8720 (N_8720,N_8446,N_8247);
or U8721 (N_8721,N_8131,N_8480);
nor U8722 (N_8722,N_8256,N_8209);
nand U8723 (N_8723,N_8039,N_8249);
and U8724 (N_8724,N_8302,N_8025);
nand U8725 (N_8725,N_8087,N_8301);
nand U8726 (N_8726,N_8481,N_8089);
and U8727 (N_8727,N_8479,N_8297);
and U8728 (N_8728,N_8153,N_8361);
nor U8729 (N_8729,N_8374,N_8142);
nor U8730 (N_8730,N_8117,N_8110);
and U8731 (N_8731,N_8414,N_8009);
and U8732 (N_8732,N_8040,N_8165);
nand U8733 (N_8733,N_8108,N_8242);
or U8734 (N_8734,N_8072,N_8452);
xor U8735 (N_8735,N_8204,N_8314);
nor U8736 (N_8736,N_8033,N_8434);
nand U8737 (N_8737,N_8012,N_8294);
nand U8738 (N_8738,N_8265,N_8112);
nor U8739 (N_8739,N_8343,N_8015);
xor U8740 (N_8740,N_8362,N_8267);
nand U8741 (N_8741,N_8067,N_8289);
or U8742 (N_8742,N_8418,N_8186);
nand U8743 (N_8743,N_8027,N_8298);
or U8744 (N_8744,N_8335,N_8489);
nand U8745 (N_8745,N_8043,N_8378);
or U8746 (N_8746,N_8435,N_8424);
and U8747 (N_8747,N_8217,N_8208);
and U8748 (N_8748,N_8307,N_8428);
nor U8749 (N_8749,N_8044,N_8339);
and U8750 (N_8750,N_8216,N_8160);
and U8751 (N_8751,N_8222,N_8471);
nand U8752 (N_8752,N_8443,N_8497);
and U8753 (N_8753,N_8030,N_8395);
nor U8754 (N_8754,N_8202,N_8468);
and U8755 (N_8755,N_8059,N_8341);
and U8756 (N_8756,N_8106,N_8013);
and U8757 (N_8757,N_8264,N_8045);
xor U8758 (N_8758,N_8163,N_8050);
or U8759 (N_8759,N_8172,N_8295);
and U8760 (N_8760,N_8137,N_8203);
and U8761 (N_8761,N_8423,N_8375);
nor U8762 (N_8762,N_8483,N_8013);
and U8763 (N_8763,N_8210,N_8437);
nand U8764 (N_8764,N_8023,N_8172);
nor U8765 (N_8765,N_8220,N_8206);
nor U8766 (N_8766,N_8490,N_8192);
and U8767 (N_8767,N_8292,N_8074);
xnor U8768 (N_8768,N_8017,N_8434);
xnor U8769 (N_8769,N_8042,N_8407);
nor U8770 (N_8770,N_8423,N_8328);
or U8771 (N_8771,N_8381,N_8415);
or U8772 (N_8772,N_8006,N_8168);
nand U8773 (N_8773,N_8240,N_8450);
and U8774 (N_8774,N_8434,N_8491);
nor U8775 (N_8775,N_8370,N_8114);
nand U8776 (N_8776,N_8080,N_8043);
or U8777 (N_8777,N_8236,N_8461);
or U8778 (N_8778,N_8236,N_8419);
and U8779 (N_8779,N_8020,N_8317);
nor U8780 (N_8780,N_8127,N_8401);
xor U8781 (N_8781,N_8490,N_8409);
xor U8782 (N_8782,N_8315,N_8380);
or U8783 (N_8783,N_8277,N_8343);
and U8784 (N_8784,N_8396,N_8064);
nor U8785 (N_8785,N_8004,N_8228);
nor U8786 (N_8786,N_8002,N_8098);
and U8787 (N_8787,N_8339,N_8224);
nor U8788 (N_8788,N_8450,N_8384);
nor U8789 (N_8789,N_8123,N_8231);
or U8790 (N_8790,N_8449,N_8432);
nor U8791 (N_8791,N_8000,N_8493);
or U8792 (N_8792,N_8113,N_8204);
xor U8793 (N_8793,N_8375,N_8053);
or U8794 (N_8794,N_8037,N_8323);
or U8795 (N_8795,N_8086,N_8061);
nor U8796 (N_8796,N_8348,N_8269);
xnor U8797 (N_8797,N_8165,N_8081);
or U8798 (N_8798,N_8235,N_8222);
nand U8799 (N_8799,N_8255,N_8022);
xor U8800 (N_8800,N_8399,N_8316);
xnor U8801 (N_8801,N_8121,N_8361);
and U8802 (N_8802,N_8287,N_8403);
nor U8803 (N_8803,N_8067,N_8127);
nand U8804 (N_8804,N_8155,N_8255);
nand U8805 (N_8805,N_8463,N_8225);
xnor U8806 (N_8806,N_8214,N_8010);
or U8807 (N_8807,N_8364,N_8264);
nand U8808 (N_8808,N_8363,N_8413);
or U8809 (N_8809,N_8236,N_8355);
nor U8810 (N_8810,N_8088,N_8488);
nor U8811 (N_8811,N_8042,N_8343);
nor U8812 (N_8812,N_8026,N_8437);
or U8813 (N_8813,N_8090,N_8391);
nand U8814 (N_8814,N_8453,N_8076);
or U8815 (N_8815,N_8463,N_8350);
nor U8816 (N_8816,N_8131,N_8356);
and U8817 (N_8817,N_8393,N_8150);
and U8818 (N_8818,N_8276,N_8491);
and U8819 (N_8819,N_8133,N_8382);
nand U8820 (N_8820,N_8184,N_8140);
and U8821 (N_8821,N_8122,N_8142);
and U8822 (N_8822,N_8216,N_8166);
or U8823 (N_8823,N_8261,N_8277);
nand U8824 (N_8824,N_8008,N_8274);
nand U8825 (N_8825,N_8301,N_8298);
nor U8826 (N_8826,N_8312,N_8453);
nor U8827 (N_8827,N_8497,N_8284);
nor U8828 (N_8828,N_8371,N_8415);
or U8829 (N_8829,N_8270,N_8292);
and U8830 (N_8830,N_8052,N_8409);
nor U8831 (N_8831,N_8408,N_8490);
nand U8832 (N_8832,N_8063,N_8307);
or U8833 (N_8833,N_8272,N_8107);
or U8834 (N_8834,N_8441,N_8205);
nand U8835 (N_8835,N_8078,N_8497);
or U8836 (N_8836,N_8397,N_8111);
nand U8837 (N_8837,N_8397,N_8106);
and U8838 (N_8838,N_8366,N_8077);
nor U8839 (N_8839,N_8050,N_8470);
or U8840 (N_8840,N_8245,N_8170);
and U8841 (N_8841,N_8478,N_8425);
or U8842 (N_8842,N_8404,N_8108);
nand U8843 (N_8843,N_8015,N_8231);
or U8844 (N_8844,N_8084,N_8034);
nor U8845 (N_8845,N_8460,N_8461);
nand U8846 (N_8846,N_8430,N_8166);
and U8847 (N_8847,N_8175,N_8266);
nand U8848 (N_8848,N_8222,N_8015);
nor U8849 (N_8849,N_8228,N_8307);
and U8850 (N_8850,N_8418,N_8069);
or U8851 (N_8851,N_8300,N_8404);
or U8852 (N_8852,N_8403,N_8361);
nand U8853 (N_8853,N_8020,N_8318);
nand U8854 (N_8854,N_8284,N_8063);
nor U8855 (N_8855,N_8112,N_8207);
nand U8856 (N_8856,N_8245,N_8076);
or U8857 (N_8857,N_8334,N_8465);
nor U8858 (N_8858,N_8022,N_8208);
or U8859 (N_8859,N_8291,N_8413);
nor U8860 (N_8860,N_8385,N_8071);
and U8861 (N_8861,N_8195,N_8015);
or U8862 (N_8862,N_8090,N_8489);
and U8863 (N_8863,N_8372,N_8015);
nor U8864 (N_8864,N_8269,N_8222);
or U8865 (N_8865,N_8436,N_8029);
or U8866 (N_8866,N_8164,N_8452);
nor U8867 (N_8867,N_8283,N_8301);
and U8868 (N_8868,N_8004,N_8124);
and U8869 (N_8869,N_8308,N_8465);
nand U8870 (N_8870,N_8076,N_8436);
xor U8871 (N_8871,N_8150,N_8475);
and U8872 (N_8872,N_8088,N_8070);
nand U8873 (N_8873,N_8273,N_8189);
nand U8874 (N_8874,N_8232,N_8242);
nand U8875 (N_8875,N_8476,N_8125);
nand U8876 (N_8876,N_8029,N_8342);
or U8877 (N_8877,N_8229,N_8323);
nor U8878 (N_8878,N_8161,N_8495);
and U8879 (N_8879,N_8097,N_8268);
and U8880 (N_8880,N_8311,N_8029);
nor U8881 (N_8881,N_8095,N_8157);
nor U8882 (N_8882,N_8175,N_8068);
or U8883 (N_8883,N_8420,N_8334);
nor U8884 (N_8884,N_8333,N_8340);
and U8885 (N_8885,N_8116,N_8023);
nand U8886 (N_8886,N_8114,N_8451);
and U8887 (N_8887,N_8012,N_8317);
and U8888 (N_8888,N_8082,N_8419);
and U8889 (N_8889,N_8201,N_8388);
nand U8890 (N_8890,N_8117,N_8168);
and U8891 (N_8891,N_8334,N_8366);
nand U8892 (N_8892,N_8011,N_8133);
or U8893 (N_8893,N_8462,N_8380);
nor U8894 (N_8894,N_8299,N_8018);
nand U8895 (N_8895,N_8098,N_8376);
nor U8896 (N_8896,N_8113,N_8371);
or U8897 (N_8897,N_8083,N_8364);
nor U8898 (N_8898,N_8428,N_8090);
or U8899 (N_8899,N_8274,N_8394);
nor U8900 (N_8900,N_8440,N_8242);
nor U8901 (N_8901,N_8143,N_8445);
and U8902 (N_8902,N_8399,N_8469);
nor U8903 (N_8903,N_8192,N_8428);
and U8904 (N_8904,N_8044,N_8448);
xor U8905 (N_8905,N_8120,N_8452);
nand U8906 (N_8906,N_8220,N_8236);
and U8907 (N_8907,N_8262,N_8266);
nand U8908 (N_8908,N_8240,N_8156);
or U8909 (N_8909,N_8373,N_8214);
xnor U8910 (N_8910,N_8231,N_8499);
or U8911 (N_8911,N_8412,N_8497);
nand U8912 (N_8912,N_8148,N_8155);
nor U8913 (N_8913,N_8297,N_8086);
nand U8914 (N_8914,N_8441,N_8310);
nand U8915 (N_8915,N_8430,N_8269);
nor U8916 (N_8916,N_8028,N_8322);
nand U8917 (N_8917,N_8151,N_8433);
or U8918 (N_8918,N_8388,N_8095);
xnor U8919 (N_8919,N_8216,N_8093);
nand U8920 (N_8920,N_8343,N_8288);
and U8921 (N_8921,N_8389,N_8498);
and U8922 (N_8922,N_8444,N_8096);
and U8923 (N_8923,N_8417,N_8017);
or U8924 (N_8924,N_8080,N_8173);
and U8925 (N_8925,N_8455,N_8111);
or U8926 (N_8926,N_8091,N_8322);
and U8927 (N_8927,N_8171,N_8452);
and U8928 (N_8928,N_8205,N_8070);
or U8929 (N_8929,N_8242,N_8181);
nor U8930 (N_8930,N_8336,N_8147);
or U8931 (N_8931,N_8200,N_8151);
or U8932 (N_8932,N_8335,N_8091);
nor U8933 (N_8933,N_8306,N_8136);
xnor U8934 (N_8934,N_8091,N_8497);
or U8935 (N_8935,N_8209,N_8078);
or U8936 (N_8936,N_8124,N_8261);
or U8937 (N_8937,N_8171,N_8234);
nand U8938 (N_8938,N_8375,N_8035);
and U8939 (N_8939,N_8388,N_8446);
or U8940 (N_8940,N_8487,N_8238);
or U8941 (N_8941,N_8007,N_8473);
nand U8942 (N_8942,N_8418,N_8081);
and U8943 (N_8943,N_8057,N_8148);
or U8944 (N_8944,N_8066,N_8085);
or U8945 (N_8945,N_8172,N_8124);
or U8946 (N_8946,N_8464,N_8191);
nand U8947 (N_8947,N_8002,N_8411);
and U8948 (N_8948,N_8490,N_8134);
nand U8949 (N_8949,N_8249,N_8344);
nand U8950 (N_8950,N_8432,N_8311);
or U8951 (N_8951,N_8127,N_8485);
nand U8952 (N_8952,N_8080,N_8225);
and U8953 (N_8953,N_8361,N_8034);
or U8954 (N_8954,N_8267,N_8057);
or U8955 (N_8955,N_8400,N_8484);
and U8956 (N_8956,N_8246,N_8388);
xor U8957 (N_8957,N_8195,N_8131);
nor U8958 (N_8958,N_8422,N_8388);
or U8959 (N_8959,N_8310,N_8304);
and U8960 (N_8960,N_8453,N_8048);
and U8961 (N_8961,N_8229,N_8273);
or U8962 (N_8962,N_8353,N_8410);
nand U8963 (N_8963,N_8017,N_8292);
and U8964 (N_8964,N_8132,N_8382);
or U8965 (N_8965,N_8277,N_8487);
or U8966 (N_8966,N_8030,N_8316);
or U8967 (N_8967,N_8440,N_8226);
and U8968 (N_8968,N_8493,N_8223);
xnor U8969 (N_8969,N_8406,N_8277);
nor U8970 (N_8970,N_8042,N_8179);
xnor U8971 (N_8971,N_8082,N_8369);
xor U8972 (N_8972,N_8233,N_8188);
nor U8973 (N_8973,N_8303,N_8083);
and U8974 (N_8974,N_8050,N_8226);
and U8975 (N_8975,N_8322,N_8078);
or U8976 (N_8976,N_8060,N_8043);
nand U8977 (N_8977,N_8243,N_8098);
and U8978 (N_8978,N_8425,N_8460);
or U8979 (N_8979,N_8466,N_8104);
nand U8980 (N_8980,N_8286,N_8227);
xor U8981 (N_8981,N_8099,N_8213);
or U8982 (N_8982,N_8016,N_8210);
nand U8983 (N_8983,N_8122,N_8454);
nor U8984 (N_8984,N_8381,N_8210);
nor U8985 (N_8985,N_8345,N_8178);
or U8986 (N_8986,N_8262,N_8111);
and U8987 (N_8987,N_8070,N_8031);
nor U8988 (N_8988,N_8471,N_8496);
nor U8989 (N_8989,N_8239,N_8187);
nor U8990 (N_8990,N_8202,N_8309);
nand U8991 (N_8991,N_8188,N_8365);
and U8992 (N_8992,N_8059,N_8132);
or U8993 (N_8993,N_8378,N_8379);
and U8994 (N_8994,N_8472,N_8475);
nand U8995 (N_8995,N_8491,N_8270);
nand U8996 (N_8996,N_8066,N_8360);
and U8997 (N_8997,N_8098,N_8385);
nor U8998 (N_8998,N_8490,N_8496);
xnor U8999 (N_8999,N_8432,N_8397);
xnor U9000 (N_9000,N_8756,N_8717);
and U9001 (N_9001,N_8951,N_8678);
and U9002 (N_9002,N_8813,N_8785);
or U9003 (N_9003,N_8591,N_8992);
nand U9004 (N_9004,N_8933,N_8626);
nor U9005 (N_9005,N_8965,N_8810);
nor U9006 (N_9006,N_8700,N_8661);
or U9007 (N_9007,N_8932,N_8574);
xnor U9008 (N_9008,N_8628,N_8924);
or U9009 (N_9009,N_8782,N_8606);
or U9010 (N_9010,N_8504,N_8572);
nand U9011 (N_9011,N_8881,N_8780);
or U9012 (N_9012,N_8950,N_8940);
nand U9013 (N_9013,N_8897,N_8788);
nor U9014 (N_9014,N_8922,N_8892);
or U9015 (N_9015,N_8869,N_8957);
and U9016 (N_9016,N_8673,N_8521);
nor U9017 (N_9017,N_8640,N_8500);
and U9018 (N_9018,N_8873,N_8835);
nand U9019 (N_9019,N_8876,N_8524);
xnor U9020 (N_9020,N_8605,N_8962);
nor U9021 (N_9021,N_8664,N_8687);
and U9022 (N_9022,N_8943,N_8989);
nor U9023 (N_9023,N_8670,N_8578);
nand U9024 (N_9024,N_8798,N_8733);
or U9025 (N_9025,N_8573,N_8783);
and U9026 (N_9026,N_8871,N_8553);
nor U9027 (N_9027,N_8637,N_8805);
xnor U9028 (N_9028,N_8523,N_8825);
nor U9029 (N_9029,N_8550,N_8784);
or U9030 (N_9030,N_8822,N_8761);
nor U9031 (N_9031,N_8826,N_8928);
xor U9032 (N_9032,N_8914,N_8773);
or U9033 (N_9033,N_8604,N_8554);
and U9034 (N_9034,N_8641,N_8985);
or U9035 (N_9035,N_8587,N_8919);
xnor U9036 (N_9036,N_8594,N_8684);
nor U9037 (N_9037,N_8565,N_8797);
or U9038 (N_9038,N_8735,N_8948);
or U9039 (N_9039,N_8693,N_8648);
or U9040 (N_9040,N_8966,N_8953);
or U9041 (N_9041,N_8958,N_8997);
nor U9042 (N_9042,N_8695,N_8839);
nand U9043 (N_9043,N_8938,N_8666);
and U9044 (N_9044,N_8506,N_8592);
xor U9045 (N_9045,N_8507,N_8724);
or U9046 (N_9046,N_8612,N_8993);
and U9047 (N_9047,N_8575,N_8767);
nand U9048 (N_9048,N_8976,N_8791);
nand U9049 (N_9049,N_8770,N_8900);
and U9050 (N_9050,N_8832,N_8636);
nor U9051 (N_9051,N_8515,N_8901);
nor U9052 (N_9052,N_8760,N_8600);
and U9053 (N_9053,N_8546,N_8580);
or U9054 (N_9054,N_8746,N_8677);
and U9055 (N_9055,N_8890,N_8833);
nand U9056 (N_9056,N_8801,N_8512);
and U9057 (N_9057,N_8729,N_8838);
and U9058 (N_9058,N_8539,N_8564);
nor U9059 (N_9059,N_8621,N_8883);
and U9060 (N_9060,N_8769,N_8759);
and U9061 (N_9061,N_8518,N_8569);
nand U9062 (N_9062,N_8669,N_8991);
or U9063 (N_9063,N_8567,N_8744);
and U9064 (N_9064,N_8638,N_8622);
nand U9065 (N_9065,N_8996,N_8541);
or U9066 (N_9066,N_8586,N_8986);
nand U9067 (N_9067,N_8676,N_8777);
nand U9068 (N_9068,N_8917,N_8624);
nor U9069 (N_9069,N_8945,N_8964);
nand U9070 (N_9070,N_8699,N_8918);
nand U9071 (N_9071,N_8821,N_8559);
nand U9072 (N_9072,N_8549,N_8776);
nor U9073 (N_9073,N_8757,N_8895);
or U9074 (N_9074,N_8696,N_8921);
nor U9075 (N_9075,N_8875,N_8834);
nor U9076 (N_9076,N_8589,N_8701);
nand U9077 (N_9077,N_8898,N_8952);
nor U9078 (N_9078,N_8905,N_8946);
nand U9079 (N_9079,N_8853,N_8610);
xor U9080 (N_9080,N_8680,N_8705);
or U9081 (N_9081,N_8625,N_8795);
xnor U9082 (N_9082,N_8845,N_8730);
nand U9083 (N_9083,N_8837,N_8796);
nand U9084 (N_9084,N_8753,N_8618);
xor U9085 (N_9085,N_8752,N_8681);
nand U9086 (N_9086,N_8935,N_8768);
nor U9087 (N_9087,N_8896,N_8887);
xor U9088 (N_9088,N_8503,N_8955);
and U9089 (N_9089,N_8536,N_8861);
nand U9090 (N_9090,N_8741,N_8979);
and U9091 (N_9091,N_8903,N_8915);
nor U9092 (N_9092,N_8601,N_8889);
xor U9093 (N_9093,N_8737,N_8763);
and U9094 (N_9094,N_8548,N_8971);
or U9095 (N_9095,N_8652,N_8519);
or U9096 (N_9096,N_8685,N_8694);
nand U9097 (N_9097,N_8584,N_8792);
nor U9098 (N_9098,N_8981,N_8959);
nand U9099 (N_9099,N_8674,N_8880);
or U9100 (N_9100,N_8818,N_8844);
nor U9101 (N_9101,N_8615,N_8501);
and U9102 (N_9102,N_8831,N_8689);
or U9103 (N_9103,N_8545,N_8806);
and U9104 (N_9104,N_8527,N_8603);
or U9105 (N_9105,N_8528,N_8639);
or U9106 (N_9106,N_8540,N_8660);
nor U9107 (N_9107,N_8855,N_8886);
and U9108 (N_9108,N_8533,N_8787);
or U9109 (N_9109,N_8929,N_8726);
and U9110 (N_9110,N_8772,N_8902);
nand U9111 (N_9111,N_8854,N_8532);
nand U9112 (N_9112,N_8894,N_8650);
or U9113 (N_9113,N_8884,N_8651);
and U9114 (N_9114,N_8697,N_8596);
and U9115 (N_9115,N_8823,N_8551);
nand U9116 (N_9116,N_8682,N_8530);
nand U9117 (N_9117,N_8631,N_8858);
or U9118 (N_9118,N_8947,N_8793);
nor U9119 (N_9119,N_8642,N_8824);
nand U9120 (N_9120,N_8885,N_8817);
nor U9121 (N_9121,N_8904,N_8585);
nor U9122 (N_9122,N_8973,N_8520);
nand U9123 (N_9123,N_8906,N_8691);
xor U9124 (N_9124,N_8653,N_8916);
xor U9125 (N_9125,N_8843,N_8703);
nor U9126 (N_9126,N_8840,N_8751);
or U9127 (N_9127,N_8960,N_8926);
and U9128 (N_9128,N_8667,N_8781);
and U9129 (N_9129,N_8830,N_8583);
nor U9130 (N_9130,N_8789,N_8702);
nor U9131 (N_9131,N_8808,N_8799);
nor U9132 (N_9132,N_8563,N_8920);
or U9133 (N_9133,N_8912,N_8942);
and U9134 (N_9134,N_8939,N_8514);
and U9135 (N_9135,N_8529,N_8850);
nand U9136 (N_9136,N_8774,N_8731);
and U9137 (N_9137,N_8516,N_8872);
nand U9138 (N_9138,N_8706,N_8613);
nor U9139 (N_9139,N_8775,N_8617);
and U9140 (N_9140,N_8627,N_8984);
nor U9141 (N_9141,N_8707,N_8794);
or U9142 (N_9142,N_8870,N_8688);
nor U9143 (N_9143,N_8629,N_8812);
or U9144 (N_9144,N_8815,N_8754);
and U9145 (N_9145,N_8925,N_8852);
or U9146 (N_9146,N_8842,N_8719);
nand U9147 (N_9147,N_8807,N_8710);
nor U9148 (N_9148,N_8786,N_8535);
nor U9149 (N_9149,N_8816,N_8597);
and U9150 (N_9150,N_8654,N_8590);
or U9151 (N_9151,N_8978,N_8848);
and U9152 (N_9152,N_8828,N_8608);
nand U9153 (N_9153,N_8690,N_8619);
and U9154 (N_9154,N_8620,N_8714);
nor U9155 (N_9155,N_8878,N_8542);
or U9156 (N_9156,N_8980,N_8593);
and U9157 (N_9157,N_8708,N_8804);
and U9158 (N_9158,N_8611,N_8561);
or U9159 (N_9159,N_8963,N_8750);
xor U9160 (N_9160,N_8909,N_8547);
or U9161 (N_9161,N_8739,N_8509);
and U9162 (N_9162,N_8709,N_8949);
nor U9163 (N_9163,N_8623,N_8930);
nand U9164 (N_9164,N_8543,N_8544);
nand U9165 (N_9165,N_8534,N_8582);
and U9166 (N_9166,N_8602,N_8647);
or U9167 (N_9167,N_8725,N_8802);
or U9168 (N_9168,N_8679,N_8556);
nor U9169 (N_9169,N_8995,N_8990);
nand U9170 (N_9170,N_8863,N_8765);
or U9171 (N_9171,N_8851,N_8982);
nor U9172 (N_9172,N_8771,N_8867);
nand U9173 (N_9173,N_8762,N_8513);
nor U9174 (N_9174,N_8662,N_8616);
or U9175 (N_9175,N_8595,N_8538);
nor U9176 (N_9176,N_8727,N_8779);
nand U9177 (N_9177,N_8931,N_8665);
nand U9178 (N_9178,N_8531,N_8923);
or U9179 (N_9179,N_8849,N_8508);
nor U9180 (N_9180,N_8809,N_8803);
or U9181 (N_9181,N_8588,N_8712);
and U9182 (N_9182,N_8656,N_8570);
nor U9183 (N_9183,N_8977,N_8899);
and U9184 (N_9184,N_8558,N_8510);
nor U9185 (N_9185,N_8755,N_8819);
and U9186 (N_9186,N_8657,N_8736);
and U9187 (N_9187,N_8658,N_8743);
or U9188 (N_9188,N_8748,N_8645);
and U9189 (N_9189,N_8599,N_8814);
nand U9190 (N_9190,N_8747,N_8841);
xor U9191 (N_9191,N_8552,N_8607);
and U9192 (N_9192,N_8882,N_8630);
xor U9193 (N_9193,N_8800,N_8745);
and U9194 (N_9194,N_8655,N_8555);
nand U9195 (N_9195,N_8633,N_8983);
xnor U9196 (N_9196,N_8864,N_8505);
or U9197 (N_9197,N_8649,N_8734);
nor U9198 (N_9198,N_8576,N_8718);
and U9199 (N_9199,N_8934,N_8988);
and U9200 (N_9200,N_8961,N_8846);
nand U9201 (N_9201,N_8723,N_8856);
nand U9202 (N_9202,N_8778,N_8738);
or U9203 (N_9203,N_8511,N_8749);
and U9204 (N_9204,N_8907,N_8634);
nand U9205 (N_9205,N_8879,N_8722);
or U9206 (N_9206,N_8632,N_8568);
or U9207 (N_9207,N_8598,N_8866);
nor U9208 (N_9208,N_8994,N_8672);
nand U9209 (N_9209,N_8865,N_8581);
or U9210 (N_9210,N_8728,N_8614);
or U9211 (N_9211,N_8937,N_8675);
nand U9212 (N_9212,N_8936,N_8713);
nor U9213 (N_9213,N_8987,N_8944);
or U9214 (N_9214,N_8663,N_8557);
nor U9215 (N_9215,N_8704,N_8891);
or U9216 (N_9216,N_8732,N_8671);
nor U9217 (N_9217,N_8659,N_8811);
nand U9218 (N_9218,N_8857,N_8954);
nand U9219 (N_9219,N_8860,N_8716);
or U9220 (N_9220,N_8790,N_8720);
nor U9221 (N_9221,N_8562,N_8566);
nand U9222 (N_9222,N_8927,N_8829);
and U9223 (N_9223,N_8571,N_8913);
or U9224 (N_9224,N_8874,N_8972);
nand U9225 (N_9225,N_8560,N_8862);
nand U9226 (N_9226,N_8969,N_8742);
and U9227 (N_9227,N_8956,N_8711);
nor U9228 (N_9228,N_8888,N_8847);
nand U9229 (N_9229,N_8836,N_8859);
or U9230 (N_9230,N_8577,N_8975);
nor U9231 (N_9231,N_8941,N_8635);
xor U9232 (N_9232,N_8766,N_8721);
and U9233 (N_9233,N_8692,N_8646);
nand U9234 (N_9234,N_8827,N_8683);
nor U9235 (N_9235,N_8998,N_8579);
nor U9236 (N_9236,N_8820,N_8502);
nand U9237 (N_9237,N_8974,N_8537);
and U9238 (N_9238,N_8643,N_8644);
nand U9239 (N_9239,N_8525,N_8698);
and U9240 (N_9240,N_8609,N_8868);
nand U9241 (N_9241,N_8686,N_8522);
or U9242 (N_9242,N_8877,N_8910);
or U9243 (N_9243,N_8999,N_8893);
and U9244 (N_9244,N_8526,N_8764);
or U9245 (N_9245,N_8967,N_8715);
or U9246 (N_9246,N_8970,N_8517);
nand U9247 (N_9247,N_8908,N_8740);
nand U9248 (N_9248,N_8968,N_8668);
and U9249 (N_9249,N_8758,N_8911);
and U9250 (N_9250,N_8616,N_8833);
nor U9251 (N_9251,N_8900,N_8511);
or U9252 (N_9252,N_8546,N_8940);
or U9253 (N_9253,N_8619,N_8751);
nor U9254 (N_9254,N_8520,N_8679);
and U9255 (N_9255,N_8607,N_8772);
nand U9256 (N_9256,N_8804,N_8940);
nor U9257 (N_9257,N_8989,N_8618);
nor U9258 (N_9258,N_8634,N_8856);
or U9259 (N_9259,N_8942,N_8594);
xor U9260 (N_9260,N_8737,N_8758);
or U9261 (N_9261,N_8961,N_8822);
or U9262 (N_9262,N_8530,N_8654);
xor U9263 (N_9263,N_8924,N_8998);
or U9264 (N_9264,N_8506,N_8562);
nand U9265 (N_9265,N_8545,N_8613);
or U9266 (N_9266,N_8851,N_8835);
nor U9267 (N_9267,N_8897,N_8791);
nor U9268 (N_9268,N_8983,N_8753);
and U9269 (N_9269,N_8662,N_8610);
and U9270 (N_9270,N_8559,N_8541);
and U9271 (N_9271,N_8846,N_8789);
nor U9272 (N_9272,N_8753,N_8649);
xor U9273 (N_9273,N_8528,N_8866);
xnor U9274 (N_9274,N_8713,N_8776);
xor U9275 (N_9275,N_8962,N_8978);
and U9276 (N_9276,N_8725,N_8795);
nand U9277 (N_9277,N_8824,N_8562);
nor U9278 (N_9278,N_8662,N_8534);
and U9279 (N_9279,N_8730,N_8564);
and U9280 (N_9280,N_8763,N_8738);
xnor U9281 (N_9281,N_8702,N_8554);
and U9282 (N_9282,N_8503,N_8664);
or U9283 (N_9283,N_8637,N_8705);
nor U9284 (N_9284,N_8869,N_8914);
and U9285 (N_9285,N_8686,N_8714);
and U9286 (N_9286,N_8949,N_8745);
or U9287 (N_9287,N_8568,N_8838);
and U9288 (N_9288,N_8722,N_8681);
and U9289 (N_9289,N_8894,N_8766);
or U9290 (N_9290,N_8695,N_8954);
or U9291 (N_9291,N_8730,N_8786);
nor U9292 (N_9292,N_8977,N_8955);
or U9293 (N_9293,N_8879,N_8573);
and U9294 (N_9294,N_8846,N_8559);
or U9295 (N_9295,N_8826,N_8859);
or U9296 (N_9296,N_8507,N_8784);
and U9297 (N_9297,N_8959,N_8903);
or U9298 (N_9298,N_8854,N_8910);
nor U9299 (N_9299,N_8715,N_8860);
and U9300 (N_9300,N_8777,N_8679);
nor U9301 (N_9301,N_8871,N_8569);
nor U9302 (N_9302,N_8846,N_8587);
and U9303 (N_9303,N_8943,N_8948);
nand U9304 (N_9304,N_8620,N_8967);
nor U9305 (N_9305,N_8765,N_8843);
or U9306 (N_9306,N_8694,N_8634);
nand U9307 (N_9307,N_8923,N_8912);
nor U9308 (N_9308,N_8678,N_8605);
and U9309 (N_9309,N_8697,N_8809);
nor U9310 (N_9310,N_8626,N_8771);
and U9311 (N_9311,N_8914,N_8550);
nor U9312 (N_9312,N_8584,N_8953);
or U9313 (N_9313,N_8867,N_8728);
and U9314 (N_9314,N_8591,N_8748);
and U9315 (N_9315,N_8548,N_8995);
nor U9316 (N_9316,N_8910,N_8784);
or U9317 (N_9317,N_8882,N_8587);
or U9318 (N_9318,N_8835,N_8570);
nand U9319 (N_9319,N_8876,N_8703);
nand U9320 (N_9320,N_8640,N_8632);
nand U9321 (N_9321,N_8641,N_8827);
and U9322 (N_9322,N_8926,N_8817);
or U9323 (N_9323,N_8722,N_8881);
or U9324 (N_9324,N_8604,N_8788);
nor U9325 (N_9325,N_8760,N_8710);
nor U9326 (N_9326,N_8968,N_8566);
and U9327 (N_9327,N_8542,N_8935);
nor U9328 (N_9328,N_8951,N_8784);
or U9329 (N_9329,N_8571,N_8850);
and U9330 (N_9330,N_8685,N_8725);
nand U9331 (N_9331,N_8978,N_8800);
nand U9332 (N_9332,N_8944,N_8583);
and U9333 (N_9333,N_8507,N_8513);
or U9334 (N_9334,N_8669,N_8898);
or U9335 (N_9335,N_8857,N_8814);
nand U9336 (N_9336,N_8984,N_8669);
nand U9337 (N_9337,N_8920,N_8685);
or U9338 (N_9338,N_8694,N_8578);
or U9339 (N_9339,N_8758,N_8808);
or U9340 (N_9340,N_8747,N_8503);
and U9341 (N_9341,N_8730,N_8793);
xnor U9342 (N_9342,N_8787,N_8931);
or U9343 (N_9343,N_8728,N_8976);
xor U9344 (N_9344,N_8823,N_8957);
nand U9345 (N_9345,N_8671,N_8559);
and U9346 (N_9346,N_8526,N_8906);
or U9347 (N_9347,N_8872,N_8515);
or U9348 (N_9348,N_8704,N_8616);
or U9349 (N_9349,N_8965,N_8707);
and U9350 (N_9350,N_8994,N_8514);
or U9351 (N_9351,N_8603,N_8670);
or U9352 (N_9352,N_8769,N_8928);
or U9353 (N_9353,N_8944,N_8661);
or U9354 (N_9354,N_8955,N_8644);
or U9355 (N_9355,N_8985,N_8970);
xor U9356 (N_9356,N_8795,N_8835);
nor U9357 (N_9357,N_8610,N_8653);
and U9358 (N_9358,N_8746,N_8642);
and U9359 (N_9359,N_8845,N_8513);
nand U9360 (N_9360,N_8829,N_8701);
and U9361 (N_9361,N_8576,N_8638);
or U9362 (N_9362,N_8792,N_8878);
nand U9363 (N_9363,N_8922,N_8963);
xor U9364 (N_9364,N_8719,N_8859);
xor U9365 (N_9365,N_8949,N_8746);
nor U9366 (N_9366,N_8710,N_8704);
xnor U9367 (N_9367,N_8579,N_8680);
and U9368 (N_9368,N_8921,N_8690);
nand U9369 (N_9369,N_8598,N_8774);
nand U9370 (N_9370,N_8614,N_8720);
nor U9371 (N_9371,N_8805,N_8645);
or U9372 (N_9372,N_8861,N_8635);
nor U9373 (N_9373,N_8676,N_8784);
nand U9374 (N_9374,N_8542,N_8709);
or U9375 (N_9375,N_8801,N_8560);
nand U9376 (N_9376,N_8833,N_8629);
nand U9377 (N_9377,N_8611,N_8938);
nand U9378 (N_9378,N_8791,N_8947);
and U9379 (N_9379,N_8935,N_8941);
xnor U9380 (N_9380,N_8813,N_8613);
and U9381 (N_9381,N_8661,N_8521);
and U9382 (N_9382,N_8688,N_8940);
nand U9383 (N_9383,N_8895,N_8889);
nand U9384 (N_9384,N_8926,N_8852);
nor U9385 (N_9385,N_8703,N_8675);
and U9386 (N_9386,N_8875,N_8636);
nor U9387 (N_9387,N_8940,N_8636);
or U9388 (N_9388,N_8521,N_8906);
or U9389 (N_9389,N_8987,N_8544);
xor U9390 (N_9390,N_8895,N_8955);
nand U9391 (N_9391,N_8627,N_8788);
and U9392 (N_9392,N_8558,N_8897);
xor U9393 (N_9393,N_8666,N_8728);
and U9394 (N_9394,N_8594,N_8510);
or U9395 (N_9395,N_8666,N_8739);
nor U9396 (N_9396,N_8815,N_8714);
nand U9397 (N_9397,N_8849,N_8504);
nor U9398 (N_9398,N_8700,N_8588);
or U9399 (N_9399,N_8872,N_8907);
xor U9400 (N_9400,N_8771,N_8892);
or U9401 (N_9401,N_8772,N_8544);
or U9402 (N_9402,N_8967,N_8534);
nor U9403 (N_9403,N_8562,N_8580);
nor U9404 (N_9404,N_8671,N_8895);
xnor U9405 (N_9405,N_8559,N_8538);
or U9406 (N_9406,N_8906,N_8558);
and U9407 (N_9407,N_8566,N_8563);
nor U9408 (N_9408,N_8616,N_8512);
and U9409 (N_9409,N_8984,N_8507);
xnor U9410 (N_9410,N_8584,N_8659);
or U9411 (N_9411,N_8520,N_8810);
or U9412 (N_9412,N_8893,N_8616);
nor U9413 (N_9413,N_8928,N_8639);
or U9414 (N_9414,N_8508,N_8644);
and U9415 (N_9415,N_8905,N_8587);
xor U9416 (N_9416,N_8951,N_8759);
nor U9417 (N_9417,N_8764,N_8500);
or U9418 (N_9418,N_8792,N_8603);
nand U9419 (N_9419,N_8673,N_8799);
nor U9420 (N_9420,N_8868,N_8790);
and U9421 (N_9421,N_8974,N_8681);
or U9422 (N_9422,N_8957,N_8965);
or U9423 (N_9423,N_8819,N_8646);
xnor U9424 (N_9424,N_8702,N_8695);
nand U9425 (N_9425,N_8611,N_8997);
and U9426 (N_9426,N_8975,N_8831);
or U9427 (N_9427,N_8573,N_8628);
nor U9428 (N_9428,N_8610,N_8712);
nor U9429 (N_9429,N_8732,N_8539);
nand U9430 (N_9430,N_8592,N_8833);
nor U9431 (N_9431,N_8551,N_8688);
nor U9432 (N_9432,N_8627,N_8849);
nand U9433 (N_9433,N_8672,N_8881);
and U9434 (N_9434,N_8930,N_8824);
nor U9435 (N_9435,N_8748,N_8973);
nand U9436 (N_9436,N_8701,N_8520);
or U9437 (N_9437,N_8941,N_8887);
nand U9438 (N_9438,N_8942,N_8617);
and U9439 (N_9439,N_8745,N_8775);
nor U9440 (N_9440,N_8710,N_8680);
or U9441 (N_9441,N_8807,N_8967);
xnor U9442 (N_9442,N_8765,N_8523);
nor U9443 (N_9443,N_8738,N_8999);
nor U9444 (N_9444,N_8947,N_8681);
and U9445 (N_9445,N_8958,N_8640);
nand U9446 (N_9446,N_8876,N_8922);
or U9447 (N_9447,N_8632,N_8854);
nand U9448 (N_9448,N_8568,N_8617);
or U9449 (N_9449,N_8658,N_8793);
nor U9450 (N_9450,N_8656,N_8583);
nor U9451 (N_9451,N_8622,N_8730);
nand U9452 (N_9452,N_8622,N_8620);
and U9453 (N_9453,N_8688,N_8939);
nor U9454 (N_9454,N_8680,N_8747);
or U9455 (N_9455,N_8987,N_8813);
nor U9456 (N_9456,N_8821,N_8503);
nand U9457 (N_9457,N_8577,N_8792);
nor U9458 (N_9458,N_8997,N_8704);
and U9459 (N_9459,N_8668,N_8946);
or U9460 (N_9460,N_8887,N_8853);
or U9461 (N_9461,N_8727,N_8844);
and U9462 (N_9462,N_8899,N_8939);
and U9463 (N_9463,N_8514,N_8614);
nand U9464 (N_9464,N_8916,N_8890);
and U9465 (N_9465,N_8884,N_8816);
and U9466 (N_9466,N_8967,N_8676);
and U9467 (N_9467,N_8768,N_8976);
and U9468 (N_9468,N_8839,N_8919);
nor U9469 (N_9469,N_8750,N_8585);
nor U9470 (N_9470,N_8549,N_8775);
xor U9471 (N_9471,N_8675,N_8830);
nor U9472 (N_9472,N_8604,N_8891);
nand U9473 (N_9473,N_8704,N_8519);
xnor U9474 (N_9474,N_8836,N_8938);
xnor U9475 (N_9475,N_8927,N_8701);
nand U9476 (N_9476,N_8943,N_8740);
or U9477 (N_9477,N_8802,N_8689);
or U9478 (N_9478,N_8525,N_8785);
or U9479 (N_9479,N_8530,N_8615);
and U9480 (N_9480,N_8541,N_8945);
or U9481 (N_9481,N_8781,N_8537);
nand U9482 (N_9482,N_8696,N_8653);
or U9483 (N_9483,N_8829,N_8939);
nand U9484 (N_9484,N_8923,N_8676);
xor U9485 (N_9485,N_8840,N_8949);
nand U9486 (N_9486,N_8539,N_8723);
nand U9487 (N_9487,N_8559,N_8511);
xor U9488 (N_9488,N_8973,N_8622);
xnor U9489 (N_9489,N_8628,N_8833);
nand U9490 (N_9490,N_8828,N_8584);
or U9491 (N_9491,N_8683,N_8755);
and U9492 (N_9492,N_8891,N_8951);
xor U9493 (N_9493,N_8607,N_8561);
and U9494 (N_9494,N_8572,N_8838);
and U9495 (N_9495,N_8865,N_8623);
and U9496 (N_9496,N_8622,N_8914);
nand U9497 (N_9497,N_8616,N_8744);
and U9498 (N_9498,N_8585,N_8865);
or U9499 (N_9499,N_8940,N_8815);
xnor U9500 (N_9500,N_9333,N_9396);
or U9501 (N_9501,N_9177,N_9226);
and U9502 (N_9502,N_9379,N_9128);
or U9503 (N_9503,N_9439,N_9077);
and U9504 (N_9504,N_9014,N_9117);
or U9505 (N_9505,N_9231,N_9266);
or U9506 (N_9506,N_9331,N_9278);
and U9507 (N_9507,N_9106,N_9461);
or U9508 (N_9508,N_9310,N_9281);
and U9509 (N_9509,N_9484,N_9162);
nor U9510 (N_9510,N_9228,N_9198);
and U9511 (N_9511,N_9058,N_9359);
and U9512 (N_9512,N_9417,N_9194);
and U9513 (N_9513,N_9195,N_9068);
nand U9514 (N_9514,N_9129,N_9233);
nand U9515 (N_9515,N_9357,N_9259);
nor U9516 (N_9516,N_9366,N_9126);
nor U9517 (N_9517,N_9090,N_9097);
nor U9518 (N_9518,N_9142,N_9133);
nor U9519 (N_9519,N_9273,N_9413);
xor U9520 (N_9520,N_9254,N_9093);
or U9521 (N_9521,N_9031,N_9025);
and U9522 (N_9522,N_9176,N_9185);
nor U9523 (N_9523,N_9237,N_9472);
nand U9524 (N_9524,N_9250,N_9471);
and U9525 (N_9525,N_9258,N_9165);
nor U9526 (N_9526,N_9317,N_9111);
nand U9527 (N_9527,N_9364,N_9491);
or U9528 (N_9528,N_9375,N_9028);
and U9529 (N_9529,N_9019,N_9066);
nand U9530 (N_9530,N_9230,N_9455);
and U9531 (N_9531,N_9270,N_9393);
nand U9532 (N_9532,N_9304,N_9116);
nand U9533 (N_9533,N_9183,N_9449);
or U9534 (N_9534,N_9168,N_9114);
xnor U9535 (N_9535,N_9264,N_9144);
and U9536 (N_9536,N_9118,N_9079);
nor U9537 (N_9537,N_9420,N_9135);
nor U9538 (N_9538,N_9403,N_9401);
and U9539 (N_9539,N_9347,N_9011);
or U9540 (N_9540,N_9202,N_9042);
nand U9541 (N_9541,N_9166,N_9425);
nor U9542 (N_9542,N_9227,N_9312);
and U9543 (N_9543,N_9432,N_9170);
nand U9544 (N_9544,N_9421,N_9400);
and U9545 (N_9545,N_9285,N_9063);
nand U9546 (N_9546,N_9109,N_9130);
xnor U9547 (N_9547,N_9002,N_9302);
nand U9548 (N_9548,N_9343,N_9414);
nor U9549 (N_9549,N_9492,N_9005);
or U9550 (N_9550,N_9416,N_9143);
or U9551 (N_9551,N_9123,N_9121);
nor U9552 (N_9552,N_9460,N_9088);
or U9553 (N_9553,N_9107,N_9277);
nor U9554 (N_9554,N_9206,N_9428);
or U9555 (N_9555,N_9294,N_9145);
and U9556 (N_9556,N_9137,N_9218);
or U9557 (N_9557,N_9221,N_9394);
nand U9558 (N_9558,N_9376,N_9173);
nand U9559 (N_9559,N_9456,N_9374);
or U9560 (N_9560,N_9023,N_9332);
or U9561 (N_9561,N_9245,N_9043);
and U9562 (N_9562,N_9015,N_9493);
nor U9563 (N_9563,N_9477,N_9050);
and U9564 (N_9564,N_9267,N_9252);
nand U9565 (N_9565,N_9054,N_9037);
nor U9566 (N_9566,N_9222,N_9136);
nor U9567 (N_9567,N_9274,N_9000);
or U9568 (N_9568,N_9365,N_9371);
nor U9569 (N_9569,N_9190,N_9290);
nor U9570 (N_9570,N_9249,N_9103);
and U9571 (N_9571,N_9214,N_9418);
xor U9572 (N_9572,N_9283,N_9030);
nand U9573 (N_9573,N_9271,N_9180);
xnor U9574 (N_9574,N_9125,N_9478);
and U9575 (N_9575,N_9036,N_9391);
xnor U9576 (N_9576,N_9016,N_9435);
or U9577 (N_9577,N_9004,N_9216);
nand U9578 (N_9578,N_9051,N_9062);
nand U9579 (N_9579,N_9167,N_9263);
xnor U9580 (N_9580,N_9355,N_9352);
and U9581 (N_9581,N_9034,N_9348);
nand U9582 (N_9582,N_9453,N_9344);
xnor U9583 (N_9583,N_9392,N_9149);
and U9584 (N_9584,N_9340,N_9299);
nor U9585 (N_9585,N_9039,N_9427);
nor U9586 (N_9586,N_9434,N_9096);
nand U9587 (N_9587,N_9268,N_9415);
nand U9588 (N_9588,N_9382,N_9069);
nand U9589 (N_9589,N_9341,N_9212);
and U9590 (N_9590,N_9409,N_9372);
or U9591 (N_9591,N_9100,N_9363);
and U9592 (N_9592,N_9261,N_9354);
nand U9593 (N_9593,N_9336,N_9032);
xnor U9594 (N_9594,N_9243,N_9065);
xnor U9595 (N_9595,N_9205,N_9012);
and U9596 (N_9596,N_9072,N_9440);
xnor U9597 (N_9597,N_9351,N_9407);
nand U9598 (N_9598,N_9248,N_9181);
nor U9599 (N_9599,N_9279,N_9380);
and U9600 (N_9600,N_9321,N_9334);
nand U9601 (N_9601,N_9269,N_9369);
nor U9602 (N_9602,N_9481,N_9055);
nor U9603 (N_9603,N_9020,N_9203);
or U9604 (N_9604,N_9303,N_9318);
or U9605 (N_9605,N_9462,N_9215);
and U9606 (N_9606,N_9139,N_9127);
and U9607 (N_9607,N_9119,N_9485);
and U9608 (N_9608,N_9211,N_9309);
or U9609 (N_9609,N_9147,N_9138);
nor U9610 (N_9610,N_9091,N_9152);
or U9611 (N_9611,N_9201,N_9469);
nand U9612 (N_9612,N_9141,N_9361);
and U9613 (N_9613,N_9213,N_9419);
nor U9614 (N_9614,N_9464,N_9148);
xor U9615 (N_9615,N_9288,N_9151);
nand U9616 (N_9616,N_9092,N_9494);
or U9617 (N_9617,N_9468,N_9071);
nand U9618 (N_9618,N_9102,N_9291);
nor U9619 (N_9619,N_9330,N_9242);
and U9620 (N_9620,N_9182,N_9158);
xor U9621 (N_9621,N_9061,N_9406);
nand U9622 (N_9622,N_9257,N_9490);
nand U9623 (N_9623,N_9008,N_9164);
or U9624 (N_9624,N_9429,N_9208);
or U9625 (N_9625,N_9498,N_9099);
and U9626 (N_9626,N_9284,N_9412);
xnor U9627 (N_9627,N_9384,N_9217);
or U9628 (N_9628,N_9251,N_9404);
and U9629 (N_9629,N_9229,N_9308);
and U9630 (N_9630,N_9006,N_9431);
or U9631 (N_9631,N_9024,N_9482);
nand U9632 (N_9632,N_9045,N_9436);
nand U9633 (N_9633,N_9398,N_9265);
and U9634 (N_9634,N_9150,N_9082);
or U9635 (N_9635,N_9297,N_9387);
or U9636 (N_9636,N_9084,N_9010);
and U9637 (N_9637,N_9064,N_9232);
or U9638 (N_9638,N_9470,N_9390);
and U9639 (N_9639,N_9465,N_9169);
or U9640 (N_9640,N_9256,N_9296);
nor U9641 (N_9641,N_9163,N_9113);
or U9642 (N_9642,N_9191,N_9209);
nor U9643 (N_9643,N_9335,N_9081);
and U9644 (N_9644,N_9463,N_9224);
nand U9645 (N_9645,N_9078,N_9199);
and U9646 (N_9646,N_9153,N_9282);
xor U9647 (N_9647,N_9373,N_9241);
or U9648 (N_9648,N_9474,N_9367);
and U9649 (N_9649,N_9467,N_9052);
nor U9650 (N_9650,N_9026,N_9235);
nor U9651 (N_9651,N_9307,N_9255);
nand U9652 (N_9652,N_9017,N_9124);
or U9653 (N_9653,N_9146,N_9076);
or U9654 (N_9654,N_9326,N_9422);
or U9655 (N_9655,N_9362,N_9300);
or U9656 (N_9656,N_9075,N_9159);
or U9657 (N_9657,N_9048,N_9377);
xnor U9658 (N_9658,N_9320,N_9188);
xnor U9659 (N_9659,N_9349,N_9174);
nand U9660 (N_9660,N_9029,N_9115);
nor U9661 (N_9661,N_9247,N_9018);
and U9662 (N_9662,N_9370,N_9293);
or U9663 (N_9663,N_9060,N_9246);
nor U9664 (N_9664,N_9360,N_9324);
nor U9665 (N_9665,N_9172,N_9197);
and U9666 (N_9666,N_9356,N_9475);
and U9667 (N_9667,N_9480,N_9386);
and U9668 (N_9668,N_9171,N_9001);
or U9669 (N_9669,N_9395,N_9383);
or U9670 (N_9670,N_9388,N_9098);
or U9671 (N_9671,N_9220,N_9175);
and U9672 (N_9672,N_9094,N_9424);
nor U9673 (N_9673,N_9155,N_9437);
nor U9674 (N_9674,N_9358,N_9479);
and U9675 (N_9675,N_9179,N_9476);
xnor U9676 (N_9676,N_9445,N_9410);
nor U9677 (N_9677,N_9049,N_9311);
and U9678 (N_9678,N_9044,N_9487);
and U9679 (N_9679,N_9423,N_9306);
nor U9680 (N_9680,N_9156,N_9192);
and U9681 (N_9681,N_9027,N_9262);
and U9682 (N_9682,N_9105,N_9013);
or U9683 (N_9683,N_9134,N_9466);
and U9684 (N_9684,N_9499,N_9085);
nor U9685 (N_9685,N_9305,N_9405);
and U9686 (N_9686,N_9298,N_9448);
nor U9687 (N_9687,N_9322,N_9047);
and U9688 (N_9688,N_9033,N_9441);
and U9689 (N_9689,N_9289,N_9337);
and U9690 (N_9690,N_9319,N_9346);
or U9691 (N_9691,N_9161,N_9328);
or U9692 (N_9692,N_9488,N_9389);
nand U9693 (N_9693,N_9399,N_9187);
xnor U9694 (N_9694,N_9292,N_9240);
xnor U9695 (N_9695,N_9315,N_9059);
and U9696 (N_9696,N_9408,N_9234);
nand U9697 (N_9697,N_9046,N_9236);
and U9698 (N_9698,N_9426,N_9323);
nor U9699 (N_9699,N_9486,N_9459);
nand U9700 (N_9700,N_9193,N_9104);
nand U9701 (N_9701,N_9411,N_9207);
or U9702 (N_9702,N_9253,N_9301);
nand U9703 (N_9703,N_9009,N_9110);
or U9704 (N_9704,N_9483,N_9313);
nand U9705 (N_9705,N_9342,N_9327);
nand U9706 (N_9706,N_9452,N_9239);
and U9707 (N_9707,N_9070,N_9353);
and U9708 (N_9708,N_9200,N_9186);
nand U9709 (N_9709,N_9350,N_9444);
or U9710 (N_9710,N_9450,N_9275);
or U9711 (N_9711,N_9381,N_9041);
nor U9712 (N_9712,N_9101,N_9108);
xor U9713 (N_9713,N_9003,N_9345);
nand U9714 (N_9714,N_9457,N_9443);
or U9715 (N_9715,N_9338,N_9276);
or U9716 (N_9716,N_9067,N_9272);
or U9717 (N_9717,N_9244,N_9140);
nor U9718 (N_9718,N_9378,N_9210);
nor U9719 (N_9719,N_9087,N_9089);
or U9720 (N_9720,N_9038,N_9368);
or U9721 (N_9721,N_9178,N_9056);
and U9722 (N_9722,N_9219,N_9286);
nand U9723 (N_9723,N_9325,N_9120);
and U9724 (N_9724,N_9086,N_9122);
nor U9725 (N_9725,N_9385,N_9316);
or U9726 (N_9726,N_9446,N_9438);
or U9727 (N_9727,N_9083,N_9442);
nand U9728 (N_9728,N_9053,N_9260);
nor U9729 (N_9729,N_9497,N_9280);
or U9730 (N_9730,N_9238,N_9035);
or U9731 (N_9731,N_9225,N_9073);
nor U9732 (N_9732,N_9204,N_9112);
nand U9733 (N_9733,N_9447,N_9189);
or U9734 (N_9734,N_9131,N_9157);
nand U9735 (N_9735,N_9184,N_9057);
or U9736 (N_9736,N_9473,N_9007);
nor U9737 (N_9737,N_9458,N_9430);
xnor U9738 (N_9738,N_9496,N_9329);
nand U9739 (N_9739,N_9080,N_9223);
nor U9740 (N_9740,N_9295,N_9495);
or U9741 (N_9741,N_9021,N_9433);
and U9742 (N_9742,N_9022,N_9154);
nor U9743 (N_9743,N_9489,N_9287);
xnor U9744 (N_9744,N_9339,N_9040);
and U9745 (N_9745,N_9314,N_9402);
or U9746 (N_9746,N_9196,N_9451);
nand U9747 (N_9747,N_9160,N_9132);
xnor U9748 (N_9748,N_9397,N_9454);
xor U9749 (N_9749,N_9095,N_9074);
nor U9750 (N_9750,N_9424,N_9407);
nand U9751 (N_9751,N_9061,N_9129);
xor U9752 (N_9752,N_9434,N_9432);
nor U9753 (N_9753,N_9321,N_9351);
nor U9754 (N_9754,N_9244,N_9050);
and U9755 (N_9755,N_9420,N_9072);
and U9756 (N_9756,N_9239,N_9000);
nor U9757 (N_9757,N_9494,N_9125);
or U9758 (N_9758,N_9477,N_9220);
and U9759 (N_9759,N_9452,N_9292);
nand U9760 (N_9760,N_9458,N_9075);
nand U9761 (N_9761,N_9495,N_9200);
and U9762 (N_9762,N_9474,N_9457);
or U9763 (N_9763,N_9388,N_9134);
nand U9764 (N_9764,N_9341,N_9487);
and U9765 (N_9765,N_9200,N_9450);
nand U9766 (N_9766,N_9330,N_9123);
nor U9767 (N_9767,N_9253,N_9071);
nor U9768 (N_9768,N_9422,N_9034);
xor U9769 (N_9769,N_9293,N_9249);
nand U9770 (N_9770,N_9048,N_9148);
nand U9771 (N_9771,N_9084,N_9483);
xnor U9772 (N_9772,N_9182,N_9093);
xor U9773 (N_9773,N_9435,N_9461);
or U9774 (N_9774,N_9468,N_9497);
and U9775 (N_9775,N_9004,N_9240);
nor U9776 (N_9776,N_9062,N_9411);
or U9777 (N_9777,N_9221,N_9074);
xor U9778 (N_9778,N_9216,N_9341);
nand U9779 (N_9779,N_9385,N_9235);
and U9780 (N_9780,N_9119,N_9231);
or U9781 (N_9781,N_9305,N_9411);
or U9782 (N_9782,N_9037,N_9351);
or U9783 (N_9783,N_9351,N_9188);
nor U9784 (N_9784,N_9307,N_9021);
and U9785 (N_9785,N_9330,N_9169);
nand U9786 (N_9786,N_9380,N_9034);
nor U9787 (N_9787,N_9062,N_9115);
xor U9788 (N_9788,N_9209,N_9342);
nor U9789 (N_9789,N_9471,N_9209);
nand U9790 (N_9790,N_9054,N_9074);
nand U9791 (N_9791,N_9479,N_9471);
or U9792 (N_9792,N_9163,N_9115);
or U9793 (N_9793,N_9418,N_9045);
and U9794 (N_9794,N_9469,N_9265);
and U9795 (N_9795,N_9416,N_9017);
xnor U9796 (N_9796,N_9343,N_9176);
nand U9797 (N_9797,N_9219,N_9392);
or U9798 (N_9798,N_9497,N_9337);
xnor U9799 (N_9799,N_9067,N_9254);
nor U9800 (N_9800,N_9303,N_9040);
nand U9801 (N_9801,N_9238,N_9482);
nor U9802 (N_9802,N_9496,N_9076);
and U9803 (N_9803,N_9426,N_9042);
nand U9804 (N_9804,N_9133,N_9247);
and U9805 (N_9805,N_9493,N_9047);
and U9806 (N_9806,N_9184,N_9080);
xor U9807 (N_9807,N_9143,N_9396);
nor U9808 (N_9808,N_9435,N_9024);
and U9809 (N_9809,N_9333,N_9388);
and U9810 (N_9810,N_9004,N_9329);
nor U9811 (N_9811,N_9111,N_9327);
and U9812 (N_9812,N_9068,N_9032);
and U9813 (N_9813,N_9228,N_9233);
nand U9814 (N_9814,N_9115,N_9421);
and U9815 (N_9815,N_9346,N_9348);
nand U9816 (N_9816,N_9468,N_9044);
xor U9817 (N_9817,N_9290,N_9430);
nor U9818 (N_9818,N_9205,N_9142);
nor U9819 (N_9819,N_9048,N_9084);
or U9820 (N_9820,N_9268,N_9090);
nor U9821 (N_9821,N_9002,N_9096);
nor U9822 (N_9822,N_9314,N_9188);
nand U9823 (N_9823,N_9000,N_9408);
nand U9824 (N_9824,N_9134,N_9277);
nor U9825 (N_9825,N_9348,N_9410);
and U9826 (N_9826,N_9259,N_9186);
xor U9827 (N_9827,N_9144,N_9429);
nand U9828 (N_9828,N_9323,N_9469);
nand U9829 (N_9829,N_9000,N_9373);
nor U9830 (N_9830,N_9499,N_9015);
nand U9831 (N_9831,N_9187,N_9445);
and U9832 (N_9832,N_9392,N_9051);
nand U9833 (N_9833,N_9160,N_9157);
and U9834 (N_9834,N_9354,N_9235);
or U9835 (N_9835,N_9439,N_9349);
and U9836 (N_9836,N_9475,N_9106);
nand U9837 (N_9837,N_9323,N_9106);
nand U9838 (N_9838,N_9291,N_9314);
and U9839 (N_9839,N_9158,N_9350);
and U9840 (N_9840,N_9406,N_9318);
or U9841 (N_9841,N_9489,N_9099);
or U9842 (N_9842,N_9273,N_9473);
nor U9843 (N_9843,N_9143,N_9047);
nor U9844 (N_9844,N_9055,N_9002);
xor U9845 (N_9845,N_9048,N_9392);
and U9846 (N_9846,N_9321,N_9116);
and U9847 (N_9847,N_9007,N_9441);
nor U9848 (N_9848,N_9201,N_9298);
xnor U9849 (N_9849,N_9242,N_9435);
and U9850 (N_9850,N_9105,N_9321);
or U9851 (N_9851,N_9117,N_9310);
or U9852 (N_9852,N_9401,N_9209);
or U9853 (N_9853,N_9003,N_9204);
nand U9854 (N_9854,N_9318,N_9180);
and U9855 (N_9855,N_9470,N_9244);
xor U9856 (N_9856,N_9304,N_9495);
or U9857 (N_9857,N_9318,N_9231);
nor U9858 (N_9858,N_9021,N_9325);
xor U9859 (N_9859,N_9058,N_9405);
nand U9860 (N_9860,N_9421,N_9032);
or U9861 (N_9861,N_9453,N_9475);
and U9862 (N_9862,N_9203,N_9450);
or U9863 (N_9863,N_9092,N_9109);
or U9864 (N_9864,N_9252,N_9225);
xor U9865 (N_9865,N_9460,N_9445);
or U9866 (N_9866,N_9162,N_9447);
nand U9867 (N_9867,N_9115,N_9081);
or U9868 (N_9868,N_9456,N_9326);
or U9869 (N_9869,N_9188,N_9265);
and U9870 (N_9870,N_9200,N_9031);
and U9871 (N_9871,N_9217,N_9488);
nor U9872 (N_9872,N_9035,N_9461);
xnor U9873 (N_9873,N_9165,N_9389);
nor U9874 (N_9874,N_9290,N_9107);
and U9875 (N_9875,N_9165,N_9199);
and U9876 (N_9876,N_9330,N_9141);
or U9877 (N_9877,N_9028,N_9377);
nor U9878 (N_9878,N_9089,N_9011);
nand U9879 (N_9879,N_9009,N_9426);
nand U9880 (N_9880,N_9167,N_9221);
and U9881 (N_9881,N_9044,N_9461);
and U9882 (N_9882,N_9419,N_9252);
nor U9883 (N_9883,N_9135,N_9198);
nand U9884 (N_9884,N_9037,N_9366);
nor U9885 (N_9885,N_9116,N_9344);
nor U9886 (N_9886,N_9131,N_9253);
and U9887 (N_9887,N_9059,N_9443);
or U9888 (N_9888,N_9002,N_9481);
and U9889 (N_9889,N_9382,N_9272);
nand U9890 (N_9890,N_9286,N_9017);
nor U9891 (N_9891,N_9034,N_9237);
nand U9892 (N_9892,N_9234,N_9101);
nor U9893 (N_9893,N_9469,N_9435);
nand U9894 (N_9894,N_9440,N_9266);
and U9895 (N_9895,N_9100,N_9039);
and U9896 (N_9896,N_9350,N_9312);
or U9897 (N_9897,N_9197,N_9195);
xor U9898 (N_9898,N_9395,N_9157);
and U9899 (N_9899,N_9440,N_9391);
xor U9900 (N_9900,N_9037,N_9186);
xnor U9901 (N_9901,N_9444,N_9033);
or U9902 (N_9902,N_9092,N_9315);
nor U9903 (N_9903,N_9432,N_9025);
or U9904 (N_9904,N_9278,N_9117);
and U9905 (N_9905,N_9396,N_9239);
and U9906 (N_9906,N_9419,N_9285);
nor U9907 (N_9907,N_9122,N_9093);
or U9908 (N_9908,N_9310,N_9289);
or U9909 (N_9909,N_9057,N_9340);
and U9910 (N_9910,N_9110,N_9344);
nand U9911 (N_9911,N_9364,N_9183);
and U9912 (N_9912,N_9231,N_9337);
nor U9913 (N_9913,N_9119,N_9343);
nand U9914 (N_9914,N_9048,N_9480);
or U9915 (N_9915,N_9102,N_9294);
and U9916 (N_9916,N_9412,N_9059);
nand U9917 (N_9917,N_9073,N_9429);
nor U9918 (N_9918,N_9107,N_9153);
nand U9919 (N_9919,N_9053,N_9169);
or U9920 (N_9920,N_9052,N_9057);
nand U9921 (N_9921,N_9368,N_9305);
or U9922 (N_9922,N_9112,N_9391);
nor U9923 (N_9923,N_9238,N_9330);
or U9924 (N_9924,N_9070,N_9249);
nand U9925 (N_9925,N_9437,N_9035);
nor U9926 (N_9926,N_9255,N_9114);
nand U9927 (N_9927,N_9203,N_9001);
nor U9928 (N_9928,N_9021,N_9206);
and U9929 (N_9929,N_9362,N_9193);
nor U9930 (N_9930,N_9431,N_9465);
nand U9931 (N_9931,N_9210,N_9230);
nand U9932 (N_9932,N_9334,N_9261);
xnor U9933 (N_9933,N_9257,N_9029);
or U9934 (N_9934,N_9253,N_9242);
nor U9935 (N_9935,N_9471,N_9333);
nand U9936 (N_9936,N_9021,N_9013);
nor U9937 (N_9937,N_9234,N_9383);
nand U9938 (N_9938,N_9013,N_9101);
or U9939 (N_9939,N_9280,N_9236);
nor U9940 (N_9940,N_9410,N_9018);
nor U9941 (N_9941,N_9372,N_9320);
xnor U9942 (N_9942,N_9071,N_9110);
or U9943 (N_9943,N_9067,N_9446);
xor U9944 (N_9944,N_9072,N_9161);
and U9945 (N_9945,N_9207,N_9493);
nand U9946 (N_9946,N_9356,N_9106);
nand U9947 (N_9947,N_9499,N_9176);
nor U9948 (N_9948,N_9153,N_9418);
and U9949 (N_9949,N_9132,N_9446);
xor U9950 (N_9950,N_9443,N_9266);
nor U9951 (N_9951,N_9205,N_9356);
nor U9952 (N_9952,N_9240,N_9480);
and U9953 (N_9953,N_9173,N_9108);
xor U9954 (N_9954,N_9420,N_9334);
or U9955 (N_9955,N_9427,N_9319);
and U9956 (N_9956,N_9024,N_9079);
nor U9957 (N_9957,N_9230,N_9003);
and U9958 (N_9958,N_9420,N_9307);
nor U9959 (N_9959,N_9120,N_9386);
nor U9960 (N_9960,N_9308,N_9108);
or U9961 (N_9961,N_9447,N_9152);
and U9962 (N_9962,N_9289,N_9099);
xnor U9963 (N_9963,N_9192,N_9193);
nor U9964 (N_9964,N_9381,N_9282);
nand U9965 (N_9965,N_9273,N_9127);
xor U9966 (N_9966,N_9494,N_9308);
nor U9967 (N_9967,N_9053,N_9004);
xor U9968 (N_9968,N_9163,N_9011);
nand U9969 (N_9969,N_9483,N_9456);
nand U9970 (N_9970,N_9149,N_9358);
or U9971 (N_9971,N_9224,N_9107);
and U9972 (N_9972,N_9122,N_9301);
xor U9973 (N_9973,N_9273,N_9003);
and U9974 (N_9974,N_9031,N_9247);
nand U9975 (N_9975,N_9289,N_9058);
or U9976 (N_9976,N_9414,N_9314);
or U9977 (N_9977,N_9442,N_9217);
nor U9978 (N_9978,N_9177,N_9007);
and U9979 (N_9979,N_9025,N_9407);
and U9980 (N_9980,N_9070,N_9068);
nor U9981 (N_9981,N_9434,N_9081);
and U9982 (N_9982,N_9355,N_9176);
nand U9983 (N_9983,N_9355,N_9229);
and U9984 (N_9984,N_9294,N_9119);
and U9985 (N_9985,N_9302,N_9077);
nand U9986 (N_9986,N_9375,N_9223);
nor U9987 (N_9987,N_9137,N_9399);
nor U9988 (N_9988,N_9186,N_9217);
nand U9989 (N_9989,N_9255,N_9354);
and U9990 (N_9990,N_9276,N_9494);
xnor U9991 (N_9991,N_9478,N_9229);
and U9992 (N_9992,N_9496,N_9154);
or U9993 (N_9993,N_9071,N_9389);
and U9994 (N_9994,N_9243,N_9125);
nand U9995 (N_9995,N_9455,N_9212);
nand U9996 (N_9996,N_9265,N_9349);
nand U9997 (N_9997,N_9428,N_9097);
or U9998 (N_9998,N_9215,N_9128);
or U9999 (N_9999,N_9013,N_9077);
nand U10000 (N_10000,N_9967,N_9708);
nand U10001 (N_10001,N_9972,N_9751);
nand U10002 (N_10002,N_9553,N_9635);
and U10003 (N_10003,N_9804,N_9607);
and U10004 (N_10004,N_9620,N_9792);
or U10005 (N_10005,N_9542,N_9691);
nand U10006 (N_10006,N_9902,N_9681);
or U10007 (N_10007,N_9923,N_9827);
and U10008 (N_10008,N_9683,N_9818);
and U10009 (N_10009,N_9664,N_9991);
or U10010 (N_10010,N_9671,N_9712);
and U10011 (N_10011,N_9739,N_9651);
xnor U10012 (N_10012,N_9770,N_9548);
and U10013 (N_10013,N_9610,N_9971);
xnor U10014 (N_10014,N_9630,N_9938);
and U10015 (N_10015,N_9809,N_9703);
nand U10016 (N_10016,N_9585,N_9511);
nand U10017 (N_10017,N_9983,N_9690);
or U10018 (N_10018,N_9919,N_9978);
nor U10019 (N_10019,N_9850,N_9942);
nor U10020 (N_10020,N_9820,N_9757);
and U10021 (N_10021,N_9912,N_9611);
nor U10022 (N_10022,N_9733,N_9649);
nand U10023 (N_10023,N_9900,N_9989);
nor U10024 (N_10024,N_9903,N_9695);
or U10025 (N_10025,N_9667,N_9526);
or U10026 (N_10026,N_9737,N_9619);
or U10027 (N_10027,N_9787,N_9622);
and U10028 (N_10028,N_9752,N_9560);
and U10029 (N_10029,N_9604,N_9678);
nor U10030 (N_10030,N_9985,N_9519);
or U10031 (N_10031,N_9552,N_9931);
or U10032 (N_10032,N_9773,N_9840);
nand U10033 (N_10033,N_9582,N_9791);
xnor U10034 (N_10034,N_9735,N_9930);
nor U10035 (N_10035,N_9617,N_9569);
nor U10036 (N_10036,N_9721,N_9935);
xnor U10037 (N_10037,N_9584,N_9709);
and U10038 (N_10038,N_9963,N_9779);
nor U10039 (N_10039,N_9878,N_9587);
and U10040 (N_10040,N_9808,N_9764);
xor U10041 (N_10041,N_9730,N_9642);
or U10042 (N_10042,N_9786,N_9964);
nor U10043 (N_10043,N_9997,N_9606);
and U10044 (N_10044,N_9600,N_9823);
and U10045 (N_10045,N_9655,N_9509);
and U10046 (N_10046,N_9716,N_9951);
nand U10047 (N_10047,N_9848,N_9563);
or U10048 (N_10048,N_9676,N_9858);
xor U10049 (N_10049,N_9952,N_9504);
nand U10050 (N_10050,N_9793,N_9713);
and U10051 (N_10051,N_9707,N_9871);
nand U10052 (N_10052,N_9992,N_9557);
nand U10053 (N_10053,N_9590,N_9535);
or U10054 (N_10054,N_9982,N_9645);
nand U10055 (N_10055,N_9595,N_9814);
or U10056 (N_10056,N_9941,N_9648);
and U10057 (N_10057,N_9945,N_9614);
nor U10058 (N_10058,N_9908,N_9566);
nand U10059 (N_10059,N_9830,N_9588);
xor U10060 (N_10060,N_9940,N_9766);
xor U10061 (N_10061,N_9788,N_9843);
and U10062 (N_10062,N_9508,N_9857);
nand U10063 (N_10063,N_9864,N_9897);
and U10064 (N_10064,N_9780,N_9828);
nor U10065 (N_10065,N_9839,N_9512);
or U10066 (N_10066,N_9925,N_9973);
nand U10067 (N_10067,N_9674,N_9568);
and U10068 (N_10068,N_9663,N_9679);
xor U10069 (N_10069,N_9835,N_9816);
xor U10070 (N_10070,N_9812,N_9847);
and U10071 (N_10071,N_9826,N_9524);
nor U10072 (N_10072,N_9892,N_9662);
and U10073 (N_10073,N_9725,N_9936);
xnor U10074 (N_10074,N_9929,N_9660);
xor U10075 (N_10075,N_9795,N_9594);
and U10076 (N_10076,N_9745,N_9920);
and U10077 (N_10077,N_9571,N_9722);
xnor U10078 (N_10078,N_9898,N_9536);
or U10079 (N_10079,N_9616,N_9728);
or U10080 (N_10080,N_9956,N_9624);
nor U10081 (N_10081,N_9530,N_9562);
nand U10082 (N_10082,N_9934,N_9567);
nand U10083 (N_10083,N_9863,N_9893);
or U10084 (N_10084,N_9669,N_9979);
or U10085 (N_10085,N_9701,N_9807);
and U10086 (N_10086,N_9692,N_9589);
and U10087 (N_10087,N_9901,N_9705);
nor U10088 (N_10088,N_9924,N_9968);
or U10089 (N_10089,N_9782,N_9798);
and U10090 (N_10090,N_9746,N_9612);
nand U10091 (N_10091,N_9921,N_9647);
or U10092 (N_10092,N_9532,N_9719);
and U10093 (N_10093,N_9514,N_9704);
nand U10094 (N_10094,N_9603,N_9693);
or U10095 (N_10095,N_9797,N_9927);
or U10096 (N_10096,N_9866,N_9926);
or U10097 (N_10097,N_9928,N_9533);
nand U10098 (N_10098,N_9506,N_9986);
or U10099 (N_10099,N_9981,N_9699);
nand U10100 (N_10100,N_9834,N_9995);
or U10101 (N_10101,N_9758,N_9883);
or U10102 (N_10102,N_9911,N_9586);
nor U10103 (N_10103,N_9784,N_9748);
nor U10104 (N_10104,N_9593,N_9640);
nor U10105 (N_10105,N_9794,N_9501);
nand U10106 (N_10106,N_9854,N_9801);
nand U10107 (N_10107,N_9672,N_9505);
nor U10108 (N_10108,N_9661,N_9613);
nor U10109 (N_10109,N_9710,N_9599);
or U10110 (N_10110,N_9761,N_9546);
and U10111 (N_10111,N_9627,N_9990);
and U10112 (N_10112,N_9700,N_9829);
and U10113 (N_10113,N_9776,N_9658);
nand U10114 (N_10114,N_9743,N_9646);
or U10115 (N_10115,N_9950,N_9682);
nor U10116 (N_10116,N_9769,N_9837);
or U10117 (N_10117,N_9714,N_9522);
nand U10118 (N_10118,N_9977,N_9799);
nand U10119 (N_10119,N_9841,N_9502);
or U10120 (N_10120,N_9747,N_9849);
nand U10121 (N_10121,N_9637,N_9790);
or U10122 (N_10122,N_9803,N_9516);
nand U10123 (N_10123,N_9583,N_9984);
or U10124 (N_10124,N_9783,N_9890);
and U10125 (N_10125,N_9538,N_9574);
nor U10126 (N_10126,N_9862,N_9726);
and U10127 (N_10127,N_9680,N_9960);
or U10128 (N_10128,N_9531,N_9634);
nor U10129 (N_10129,N_9545,N_9833);
nand U10130 (N_10130,N_9891,N_9517);
and U10131 (N_10131,N_9916,N_9954);
or U10132 (N_10132,N_9975,N_9653);
nand U10133 (N_10133,N_9592,N_9772);
or U10134 (N_10134,N_9697,N_9696);
xnor U10135 (N_10135,N_9768,N_9602);
nor U10136 (N_10136,N_9887,N_9886);
nand U10137 (N_10137,N_9621,N_9876);
nand U10138 (N_10138,N_9789,N_9760);
nor U10139 (N_10139,N_9670,N_9933);
and U10140 (N_10140,N_9970,N_9570);
xnor U10141 (N_10141,N_9915,N_9836);
or U10142 (N_10142,N_9949,N_9845);
nand U10143 (N_10143,N_9742,N_9564);
nand U10144 (N_10144,N_9980,N_9503);
or U10145 (N_10145,N_9537,N_9578);
xnor U10146 (N_10146,N_9870,N_9763);
or U10147 (N_10147,N_9944,N_9852);
or U10148 (N_10148,N_9844,N_9711);
and U10149 (N_10149,N_9528,N_9518);
nor U10150 (N_10150,N_9521,N_9889);
or U10151 (N_10151,N_9994,N_9507);
and U10152 (N_10152,N_9723,N_9555);
nor U10153 (N_10153,N_9947,N_9861);
and U10154 (N_10154,N_9631,N_9907);
and U10155 (N_10155,N_9525,N_9515);
and U10156 (N_10156,N_9948,N_9724);
and U10157 (N_10157,N_9939,N_9565);
nor U10158 (N_10158,N_9608,N_9550);
or U10159 (N_10159,N_9686,N_9744);
nand U10160 (N_10160,N_9668,N_9987);
nand U10161 (N_10161,N_9615,N_9632);
nand U10162 (N_10162,N_9846,N_9922);
or U10163 (N_10163,N_9937,N_9754);
nor U10164 (N_10164,N_9838,N_9596);
nor U10165 (N_10165,N_9759,N_9626);
nor U10166 (N_10166,N_9549,N_9961);
or U10167 (N_10167,N_9706,N_9666);
nand U10168 (N_10168,N_9554,N_9675);
and U10169 (N_10169,N_9687,N_9867);
nor U10170 (N_10170,N_9685,N_9551);
xor U10171 (N_10171,N_9729,N_9623);
nand U10172 (N_10172,N_9811,N_9962);
xor U10173 (N_10173,N_9529,N_9873);
or U10174 (N_10174,N_9643,N_9520);
and U10175 (N_10175,N_9727,N_9762);
and U10176 (N_10176,N_9625,N_9917);
or U10177 (N_10177,N_9998,N_9715);
nor U10178 (N_10178,N_9976,N_9894);
nand U10179 (N_10179,N_9800,N_9741);
nor U10180 (N_10180,N_9556,N_9832);
and U10181 (N_10181,N_9644,N_9575);
nand U10182 (N_10182,N_9918,N_9825);
nor U10183 (N_10183,N_9543,N_9999);
xor U10184 (N_10184,N_9581,N_9822);
xor U10185 (N_10185,N_9765,N_9905);
nor U10186 (N_10186,N_9572,N_9677);
and U10187 (N_10187,N_9896,N_9598);
nor U10188 (N_10188,N_9969,N_9573);
or U10189 (N_10189,N_9547,N_9698);
nor U10190 (N_10190,N_9628,N_9767);
and U10191 (N_10191,N_9539,N_9943);
nand U10192 (N_10192,N_9872,N_9510);
nor U10193 (N_10193,N_9885,N_9738);
and U10194 (N_10194,N_9534,N_9781);
nor U10195 (N_10195,N_9946,N_9753);
or U10196 (N_10196,N_9988,N_9601);
nor U10197 (N_10197,N_9734,N_9880);
nand U10198 (N_10198,N_9824,N_9884);
and U10199 (N_10199,N_9877,N_9577);
nand U10200 (N_10200,N_9815,N_9959);
or U10201 (N_10201,N_9673,N_9541);
xor U10202 (N_10202,N_9955,N_9775);
and U10203 (N_10203,N_9558,N_9875);
nand U10204 (N_10204,N_9659,N_9591);
xnor U10205 (N_10205,N_9813,N_9993);
nand U10206 (N_10206,N_9717,N_9906);
nand U10207 (N_10207,N_9500,N_9656);
and U10208 (N_10208,N_9881,N_9879);
xnor U10209 (N_10209,N_9579,N_9639);
or U10210 (N_10210,N_9720,N_9910);
and U10211 (N_10211,N_9932,N_9810);
nor U10212 (N_10212,N_9731,N_9821);
or U10213 (N_10213,N_9868,N_9540);
and U10214 (N_10214,N_9806,N_9974);
nand U10215 (N_10215,N_9851,N_9778);
or U10216 (N_10216,N_9831,N_9633);
xnor U10217 (N_10217,N_9888,N_9913);
and U10218 (N_10218,N_9774,N_9750);
nor U10219 (N_10219,N_9842,N_9771);
nand U10220 (N_10220,N_9694,N_9652);
nor U10221 (N_10221,N_9732,N_9618);
nor U10222 (N_10222,N_9689,N_9580);
nand U10223 (N_10223,N_9641,N_9638);
nor U10224 (N_10224,N_9869,N_9865);
nand U10225 (N_10225,N_9605,N_9914);
nor U10226 (N_10226,N_9654,N_9629);
or U10227 (N_10227,N_9576,N_9688);
and U10228 (N_10228,N_9965,N_9702);
and U10229 (N_10229,N_9904,N_9609);
nand U10230 (N_10230,N_9874,N_9882);
and U10231 (N_10231,N_9597,N_9718);
nor U10232 (N_10232,N_9953,N_9755);
or U10233 (N_10233,N_9860,N_9650);
nor U10234 (N_10234,N_9749,N_9957);
or U10235 (N_10235,N_9561,N_9909);
nor U10236 (N_10236,N_9665,N_9684);
nand U10237 (N_10237,N_9777,N_9740);
xnor U10238 (N_10238,N_9544,N_9527);
nand U10239 (N_10239,N_9853,N_9855);
and U10240 (N_10240,N_9817,N_9819);
xor U10241 (N_10241,N_9796,N_9513);
or U10242 (N_10242,N_9895,N_9756);
nand U10243 (N_10243,N_9958,N_9802);
and U10244 (N_10244,N_9736,N_9636);
nor U10245 (N_10245,N_9859,N_9559);
and U10246 (N_10246,N_9856,N_9657);
nor U10247 (N_10247,N_9785,N_9523);
nor U10248 (N_10248,N_9996,N_9966);
and U10249 (N_10249,N_9805,N_9899);
and U10250 (N_10250,N_9895,N_9738);
nand U10251 (N_10251,N_9671,N_9748);
nor U10252 (N_10252,N_9871,N_9873);
or U10253 (N_10253,N_9994,N_9554);
nand U10254 (N_10254,N_9754,N_9608);
and U10255 (N_10255,N_9898,N_9661);
nor U10256 (N_10256,N_9629,N_9843);
nor U10257 (N_10257,N_9842,N_9683);
and U10258 (N_10258,N_9717,N_9855);
and U10259 (N_10259,N_9884,N_9629);
nand U10260 (N_10260,N_9979,N_9952);
and U10261 (N_10261,N_9560,N_9997);
nand U10262 (N_10262,N_9611,N_9971);
xor U10263 (N_10263,N_9943,N_9962);
nand U10264 (N_10264,N_9558,N_9614);
nor U10265 (N_10265,N_9692,N_9503);
nand U10266 (N_10266,N_9717,N_9963);
and U10267 (N_10267,N_9915,N_9700);
and U10268 (N_10268,N_9724,N_9608);
or U10269 (N_10269,N_9892,N_9730);
nor U10270 (N_10270,N_9721,N_9959);
nor U10271 (N_10271,N_9852,N_9986);
xor U10272 (N_10272,N_9727,N_9566);
nor U10273 (N_10273,N_9876,N_9551);
and U10274 (N_10274,N_9971,N_9513);
nor U10275 (N_10275,N_9752,N_9734);
or U10276 (N_10276,N_9541,N_9682);
and U10277 (N_10277,N_9823,N_9583);
and U10278 (N_10278,N_9504,N_9839);
nand U10279 (N_10279,N_9997,N_9814);
xor U10280 (N_10280,N_9679,N_9914);
nand U10281 (N_10281,N_9691,N_9582);
or U10282 (N_10282,N_9802,N_9964);
nand U10283 (N_10283,N_9650,N_9902);
or U10284 (N_10284,N_9918,N_9979);
nand U10285 (N_10285,N_9718,N_9698);
or U10286 (N_10286,N_9621,N_9767);
xor U10287 (N_10287,N_9605,N_9614);
nand U10288 (N_10288,N_9784,N_9768);
nand U10289 (N_10289,N_9716,N_9696);
nor U10290 (N_10290,N_9882,N_9710);
xnor U10291 (N_10291,N_9771,N_9892);
nand U10292 (N_10292,N_9591,N_9562);
or U10293 (N_10293,N_9792,N_9619);
and U10294 (N_10294,N_9838,N_9502);
and U10295 (N_10295,N_9844,N_9668);
or U10296 (N_10296,N_9774,N_9695);
nor U10297 (N_10297,N_9608,N_9715);
nor U10298 (N_10298,N_9765,N_9990);
nand U10299 (N_10299,N_9771,N_9944);
xor U10300 (N_10300,N_9702,N_9583);
nand U10301 (N_10301,N_9917,N_9975);
xor U10302 (N_10302,N_9712,N_9862);
nor U10303 (N_10303,N_9802,N_9749);
and U10304 (N_10304,N_9836,N_9871);
or U10305 (N_10305,N_9726,N_9647);
and U10306 (N_10306,N_9621,N_9580);
nor U10307 (N_10307,N_9992,N_9616);
and U10308 (N_10308,N_9514,N_9712);
or U10309 (N_10309,N_9532,N_9632);
or U10310 (N_10310,N_9561,N_9550);
and U10311 (N_10311,N_9519,N_9820);
xnor U10312 (N_10312,N_9921,N_9852);
nor U10313 (N_10313,N_9908,N_9991);
and U10314 (N_10314,N_9571,N_9697);
or U10315 (N_10315,N_9981,N_9618);
nand U10316 (N_10316,N_9717,N_9946);
nand U10317 (N_10317,N_9766,N_9563);
xor U10318 (N_10318,N_9672,N_9609);
xnor U10319 (N_10319,N_9921,N_9614);
or U10320 (N_10320,N_9661,N_9590);
nor U10321 (N_10321,N_9638,N_9657);
and U10322 (N_10322,N_9900,N_9551);
nand U10323 (N_10323,N_9619,N_9855);
or U10324 (N_10324,N_9510,N_9748);
or U10325 (N_10325,N_9937,N_9893);
nor U10326 (N_10326,N_9571,N_9962);
and U10327 (N_10327,N_9851,N_9538);
or U10328 (N_10328,N_9524,N_9531);
or U10329 (N_10329,N_9951,N_9822);
and U10330 (N_10330,N_9768,N_9890);
or U10331 (N_10331,N_9807,N_9988);
nor U10332 (N_10332,N_9822,N_9546);
or U10333 (N_10333,N_9975,N_9940);
and U10334 (N_10334,N_9601,N_9840);
nand U10335 (N_10335,N_9910,N_9970);
nor U10336 (N_10336,N_9565,N_9964);
or U10337 (N_10337,N_9889,N_9545);
nand U10338 (N_10338,N_9587,N_9629);
nor U10339 (N_10339,N_9729,N_9758);
or U10340 (N_10340,N_9995,N_9852);
and U10341 (N_10341,N_9888,N_9717);
or U10342 (N_10342,N_9683,N_9759);
nor U10343 (N_10343,N_9802,N_9514);
and U10344 (N_10344,N_9681,N_9952);
xor U10345 (N_10345,N_9901,N_9802);
or U10346 (N_10346,N_9624,N_9971);
and U10347 (N_10347,N_9721,N_9945);
and U10348 (N_10348,N_9793,N_9630);
nand U10349 (N_10349,N_9635,N_9628);
and U10350 (N_10350,N_9870,N_9850);
or U10351 (N_10351,N_9538,N_9663);
nand U10352 (N_10352,N_9857,N_9872);
nor U10353 (N_10353,N_9945,N_9868);
and U10354 (N_10354,N_9793,N_9773);
and U10355 (N_10355,N_9851,N_9592);
nand U10356 (N_10356,N_9720,N_9923);
nand U10357 (N_10357,N_9916,N_9800);
nand U10358 (N_10358,N_9914,N_9875);
or U10359 (N_10359,N_9903,N_9980);
and U10360 (N_10360,N_9979,N_9675);
nand U10361 (N_10361,N_9683,N_9825);
nand U10362 (N_10362,N_9622,N_9829);
nand U10363 (N_10363,N_9696,N_9546);
or U10364 (N_10364,N_9542,N_9817);
or U10365 (N_10365,N_9930,N_9513);
xnor U10366 (N_10366,N_9559,N_9533);
nand U10367 (N_10367,N_9768,N_9883);
xnor U10368 (N_10368,N_9549,N_9569);
xor U10369 (N_10369,N_9835,N_9833);
and U10370 (N_10370,N_9776,N_9808);
nand U10371 (N_10371,N_9710,N_9890);
and U10372 (N_10372,N_9587,N_9526);
nand U10373 (N_10373,N_9942,N_9691);
nand U10374 (N_10374,N_9704,N_9910);
or U10375 (N_10375,N_9880,N_9751);
nor U10376 (N_10376,N_9647,N_9972);
or U10377 (N_10377,N_9555,N_9844);
and U10378 (N_10378,N_9625,N_9723);
or U10379 (N_10379,N_9693,N_9792);
nor U10380 (N_10380,N_9877,N_9747);
xnor U10381 (N_10381,N_9519,N_9886);
nor U10382 (N_10382,N_9719,N_9508);
nor U10383 (N_10383,N_9712,N_9777);
nor U10384 (N_10384,N_9766,N_9578);
and U10385 (N_10385,N_9962,N_9891);
or U10386 (N_10386,N_9894,N_9541);
nor U10387 (N_10387,N_9968,N_9844);
or U10388 (N_10388,N_9697,N_9768);
xor U10389 (N_10389,N_9916,N_9819);
nand U10390 (N_10390,N_9741,N_9894);
nand U10391 (N_10391,N_9615,N_9815);
or U10392 (N_10392,N_9750,N_9934);
xor U10393 (N_10393,N_9823,N_9741);
and U10394 (N_10394,N_9561,N_9825);
nand U10395 (N_10395,N_9701,N_9603);
or U10396 (N_10396,N_9920,N_9563);
xnor U10397 (N_10397,N_9806,N_9665);
nand U10398 (N_10398,N_9917,N_9751);
nor U10399 (N_10399,N_9632,N_9997);
nand U10400 (N_10400,N_9980,N_9992);
and U10401 (N_10401,N_9544,N_9722);
nor U10402 (N_10402,N_9824,N_9707);
nand U10403 (N_10403,N_9684,N_9846);
xnor U10404 (N_10404,N_9941,N_9794);
or U10405 (N_10405,N_9917,N_9576);
and U10406 (N_10406,N_9692,N_9724);
nor U10407 (N_10407,N_9718,N_9704);
and U10408 (N_10408,N_9595,N_9993);
or U10409 (N_10409,N_9954,N_9532);
and U10410 (N_10410,N_9888,N_9673);
nand U10411 (N_10411,N_9596,N_9725);
or U10412 (N_10412,N_9591,N_9670);
nand U10413 (N_10413,N_9957,N_9542);
and U10414 (N_10414,N_9596,N_9649);
or U10415 (N_10415,N_9969,N_9681);
xnor U10416 (N_10416,N_9661,N_9946);
nor U10417 (N_10417,N_9808,N_9716);
and U10418 (N_10418,N_9858,N_9564);
or U10419 (N_10419,N_9904,N_9965);
and U10420 (N_10420,N_9532,N_9934);
nor U10421 (N_10421,N_9815,N_9887);
nor U10422 (N_10422,N_9707,N_9548);
nor U10423 (N_10423,N_9562,N_9791);
and U10424 (N_10424,N_9675,N_9548);
nor U10425 (N_10425,N_9613,N_9780);
nand U10426 (N_10426,N_9759,N_9997);
and U10427 (N_10427,N_9948,N_9547);
nor U10428 (N_10428,N_9559,N_9657);
or U10429 (N_10429,N_9530,N_9606);
nor U10430 (N_10430,N_9965,N_9955);
xnor U10431 (N_10431,N_9607,N_9920);
and U10432 (N_10432,N_9661,N_9871);
nor U10433 (N_10433,N_9502,N_9753);
nor U10434 (N_10434,N_9864,N_9796);
nor U10435 (N_10435,N_9887,N_9809);
and U10436 (N_10436,N_9787,N_9999);
nor U10437 (N_10437,N_9733,N_9949);
and U10438 (N_10438,N_9849,N_9595);
or U10439 (N_10439,N_9518,N_9707);
and U10440 (N_10440,N_9567,N_9963);
xor U10441 (N_10441,N_9615,N_9551);
nor U10442 (N_10442,N_9885,N_9904);
and U10443 (N_10443,N_9529,N_9853);
nor U10444 (N_10444,N_9555,N_9530);
nor U10445 (N_10445,N_9509,N_9987);
nand U10446 (N_10446,N_9912,N_9661);
and U10447 (N_10447,N_9811,N_9797);
and U10448 (N_10448,N_9899,N_9764);
and U10449 (N_10449,N_9508,N_9535);
and U10450 (N_10450,N_9570,N_9976);
or U10451 (N_10451,N_9629,N_9925);
nand U10452 (N_10452,N_9862,N_9854);
and U10453 (N_10453,N_9897,N_9788);
nor U10454 (N_10454,N_9519,N_9796);
nor U10455 (N_10455,N_9520,N_9542);
nand U10456 (N_10456,N_9787,N_9916);
and U10457 (N_10457,N_9814,N_9820);
nor U10458 (N_10458,N_9778,N_9591);
or U10459 (N_10459,N_9776,N_9502);
nor U10460 (N_10460,N_9765,N_9676);
xnor U10461 (N_10461,N_9727,N_9787);
nor U10462 (N_10462,N_9951,N_9601);
or U10463 (N_10463,N_9933,N_9593);
and U10464 (N_10464,N_9545,N_9685);
nand U10465 (N_10465,N_9587,N_9822);
nor U10466 (N_10466,N_9925,N_9752);
nand U10467 (N_10467,N_9983,N_9647);
xor U10468 (N_10468,N_9678,N_9779);
xnor U10469 (N_10469,N_9600,N_9897);
or U10470 (N_10470,N_9780,N_9507);
nand U10471 (N_10471,N_9721,N_9505);
nor U10472 (N_10472,N_9504,N_9996);
nand U10473 (N_10473,N_9995,N_9526);
nor U10474 (N_10474,N_9658,N_9525);
nand U10475 (N_10475,N_9967,N_9808);
or U10476 (N_10476,N_9522,N_9908);
and U10477 (N_10477,N_9525,N_9645);
nor U10478 (N_10478,N_9858,N_9850);
or U10479 (N_10479,N_9531,N_9839);
nor U10480 (N_10480,N_9853,N_9539);
and U10481 (N_10481,N_9910,N_9630);
and U10482 (N_10482,N_9628,N_9604);
nor U10483 (N_10483,N_9794,N_9808);
or U10484 (N_10484,N_9593,N_9711);
nand U10485 (N_10485,N_9855,N_9676);
nand U10486 (N_10486,N_9863,N_9784);
nand U10487 (N_10487,N_9520,N_9841);
nor U10488 (N_10488,N_9757,N_9801);
or U10489 (N_10489,N_9685,N_9600);
nand U10490 (N_10490,N_9983,N_9991);
nor U10491 (N_10491,N_9818,N_9635);
and U10492 (N_10492,N_9706,N_9877);
nor U10493 (N_10493,N_9599,N_9644);
nand U10494 (N_10494,N_9976,N_9686);
xnor U10495 (N_10495,N_9765,N_9968);
nand U10496 (N_10496,N_9817,N_9594);
or U10497 (N_10497,N_9605,N_9581);
or U10498 (N_10498,N_9517,N_9759);
nor U10499 (N_10499,N_9584,N_9950);
nor U10500 (N_10500,N_10469,N_10118);
and U10501 (N_10501,N_10162,N_10462);
nand U10502 (N_10502,N_10359,N_10066);
or U10503 (N_10503,N_10116,N_10276);
nand U10504 (N_10504,N_10295,N_10395);
nor U10505 (N_10505,N_10358,N_10402);
or U10506 (N_10506,N_10060,N_10131);
and U10507 (N_10507,N_10144,N_10254);
or U10508 (N_10508,N_10471,N_10312);
nand U10509 (N_10509,N_10330,N_10311);
or U10510 (N_10510,N_10408,N_10445);
nor U10511 (N_10511,N_10309,N_10365);
nand U10512 (N_10512,N_10499,N_10238);
nand U10513 (N_10513,N_10009,N_10087);
nor U10514 (N_10514,N_10004,N_10290);
and U10515 (N_10515,N_10433,N_10383);
nand U10516 (N_10516,N_10049,N_10458);
and U10517 (N_10517,N_10135,N_10270);
or U10518 (N_10518,N_10297,N_10455);
nand U10519 (N_10519,N_10448,N_10089);
and U10520 (N_10520,N_10435,N_10377);
nand U10521 (N_10521,N_10424,N_10076);
nand U10522 (N_10522,N_10029,N_10476);
or U10523 (N_10523,N_10337,N_10257);
nand U10524 (N_10524,N_10228,N_10288);
xnor U10525 (N_10525,N_10179,N_10074);
and U10526 (N_10526,N_10129,N_10304);
and U10527 (N_10527,N_10474,N_10430);
nand U10528 (N_10528,N_10071,N_10081);
nor U10529 (N_10529,N_10022,N_10298);
nor U10530 (N_10530,N_10479,N_10472);
xnor U10531 (N_10531,N_10478,N_10077);
and U10532 (N_10532,N_10127,N_10230);
nor U10533 (N_10533,N_10280,N_10194);
nand U10534 (N_10534,N_10209,N_10369);
and U10535 (N_10535,N_10102,N_10157);
nor U10536 (N_10536,N_10044,N_10450);
nor U10537 (N_10537,N_10037,N_10006);
or U10538 (N_10538,N_10013,N_10193);
xnor U10539 (N_10539,N_10030,N_10176);
nand U10540 (N_10540,N_10360,N_10262);
or U10541 (N_10541,N_10196,N_10042);
nand U10542 (N_10542,N_10267,N_10082);
or U10543 (N_10543,N_10436,N_10463);
nor U10544 (N_10544,N_10405,N_10412);
and U10545 (N_10545,N_10331,N_10063);
nor U10546 (N_10546,N_10368,N_10158);
nand U10547 (N_10547,N_10454,N_10341);
and U10548 (N_10548,N_10361,N_10198);
and U10549 (N_10549,N_10021,N_10390);
nor U10550 (N_10550,N_10173,N_10495);
nand U10551 (N_10551,N_10409,N_10091);
or U10552 (N_10552,N_10114,N_10261);
nand U10553 (N_10553,N_10109,N_10352);
nor U10554 (N_10554,N_10213,N_10370);
nand U10555 (N_10555,N_10175,N_10340);
and U10556 (N_10556,N_10374,N_10200);
or U10557 (N_10557,N_10483,N_10201);
and U10558 (N_10558,N_10246,N_10317);
or U10559 (N_10559,N_10307,N_10052);
xor U10560 (N_10560,N_10229,N_10180);
and U10561 (N_10561,N_10010,N_10237);
nor U10562 (N_10562,N_10155,N_10249);
nand U10563 (N_10563,N_10014,N_10301);
and U10564 (N_10564,N_10147,N_10443);
xnor U10565 (N_10565,N_10349,N_10467);
nor U10566 (N_10566,N_10391,N_10335);
and U10567 (N_10567,N_10028,N_10453);
and U10568 (N_10568,N_10070,N_10165);
or U10569 (N_10569,N_10065,N_10036);
and U10570 (N_10570,N_10278,N_10425);
and U10571 (N_10571,N_10123,N_10199);
xnor U10572 (N_10572,N_10112,N_10417);
or U10573 (N_10573,N_10289,N_10258);
or U10574 (N_10574,N_10168,N_10452);
nand U10575 (N_10575,N_10306,N_10464);
or U10576 (N_10576,N_10303,N_10224);
nor U10577 (N_10577,N_10308,N_10061);
or U10578 (N_10578,N_10475,N_10015);
nor U10579 (N_10579,N_10273,N_10183);
and U10580 (N_10580,N_10149,N_10055);
or U10581 (N_10581,N_10414,N_10172);
and U10582 (N_10582,N_10287,N_10038);
nand U10583 (N_10583,N_10461,N_10160);
nor U10584 (N_10584,N_10053,N_10045);
nor U10585 (N_10585,N_10210,N_10411);
nor U10586 (N_10586,N_10326,N_10206);
nand U10587 (N_10587,N_10299,N_10039);
nor U10588 (N_10588,N_10367,N_10020);
xor U10589 (N_10589,N_10484,N_10470);
nor U10590 (N_10590,N_10465,N_10381);
nor U10591 (N_10591,N_10387,N_10423);
and U10592 (N_10592,N_10323,N_10342);
or U10593 (N_10593,N_10275,N_10274);
or U10594 (N_10594,N_10320,N_10001);
and U10595 (N_10595,N_10272,N_10447);
nor U10596 (N_10596,N_10388,N_10373);
nor U10597 (N_10597,N_10211,N_10148);
and U10598 (N_10598,N_10120,N_10121);
xnor U10599 (N_10599,N_10117,N_10394);
nor U10600 (N_10600,N_10185,N_10104);
and U10601 (N_10601,N_10159,N_10489);
nand U10602 (N_10602,N_10333,N_10446);
nor U10603 (N_10603,N_10018,N_10134);
nor U10604 (N_10604,N_10107,N_10332);
nand U10605 (N_10605,N_10233,N_10404);
nor U10606 (N_10606,N_10418,N_10236);
nand U10607 (N_10607,N_10043,N_10410);
nor U10608 (N_10608,N_10386,N_10354);
or U10609 (N_10609,N_10182,N_10119);
nor U10610 (N_10610,N_10439,N_10442);
nor U10611 (N_10611,N_10048,N_10217);
nor U10612 (N_10612,N_10026,N_10054);
xor U10613 (N_10613,N_10046,N_10285);
or U10614 (N_10614,N_10480,N_10145);
and U10615 (N_10615,N_10428,N_10327);
and U10616 (N_10616,N_10169,N_10313);
or U10617 (N_10617,N_10466,N_10371);
and U10618 (N_10618,N_10456,N_10041);
xnor U10619 (N_10619,N_10385,N_10392);
or U10620 (N_10620,N_10372,N_10243);
or U10621 (N_10621,N_10379,N_10449);
nor U10622 (N_10622,N_10033,N_10226);
nor U10623 (N_10623,N_10204,N_10429);
nand U10624 (N_10624,N_10079,N_10459);
or U10625 (N_10625,N_10012,N_10247);
or U10626 (N_10626,N_10032,N_10348);
or U10627 (N_10627,N_10399,N_10396);
and U10628 (N_10628,N_10178,N_10059);
xnor U10629 (N_10629,N_10259,N_10086);
and U10630 (N_10630,N_10181,N_10212);
or U10631 (N_10631,N_10232,N_10137);
and U10632 (N_10632,N_10031,N_10419);
nor U10633 (N_10633,N_10005,N_10197);
and U10634 (N_10634,N_10080,N_10207);
nand U10635 (N_10635,N_10092,N_10177);
xor U10636 (N_10636,N_10393,N_10122);
and U10637 (N_10637,N_10034,N_10490);
nand U10638 (N_10638,N_10191,N_10085);
or U10639 (N_10639,N_10110,N_10477);
or U10640 (N_10640,N_10138,N_10328);
nor U10641 (N_10641,N_10141,N_10072);
nand U10642 (N_10642,N_10253,N_10265);
or U10643 (N_10643,N_10397,N_10468);
nor U10644 (N_10644,N_10170,N_10111);
and U10645 (N_10645,N_10315,N_10353);
and U10646 (N_10646,N_10338,N_10356);
nand U10647 (N_10647,N_10345,N_10451);
and U10648 (N_10648,N_10271,N_10222);
nor U10649 (N_10649,N_10310,N_10432);
and U10650 (N_10650,N_10460,N_10318);
nand U10651 (N_10651,N_10486,N_10281);
nand U10652 (N_10652,N_10093,N_10362);
or U10653 (N_10653,N_10305,N_10140);
and U10654 (N_10654,N_10164,N_10019);
nor U10655 (N_10655,N_10167,N_10398);
and U10656 (N_10656,N_10284,N_10251);
nor U10657 (N_10657,N_10151,N_10401);
nand U10658 (N_10658,N_10203,N_10314);
nor U10659 (N_10659,N_10427,N_10067);
and U10660 (N_10660,N_10426,N_10171);
nor U10661 (N_10661,N_10047,N_10223);
nand U10662 (N_10662,N_10498,N_10344);
nand U10663 (N_10663,N_10282,N_10094);
xor U10664 (N_10664,N_10056,N_10421);
and U10665 (N_10665,N_10132,N_10139);
and U10666 (N_10666,N_10413,N_10146);
nor U10667 (N_10667,N_10336,N_10035);
nand U10668 (N_10668,N_10380,N_10062);
or U10669 (N_10669,N_10153,N_10161);
and U10670 (N_10670,N_10090,N_10441);
nand U10671 (N_10671,N_10188,N_10050);
nor U10672 (N_10672,N_10378,N_10115);
nand U10673 (N_10673,N_10103,N_10095);
nor U10674 (N_10674,N_10069,N_10269);
or U10675 (N_10675,N_10366,N_10389);
or U10676 (N_10676,N_10248,N_10126);
nand U10677 (N_10677,N_10219,N_10231);
nand U10678 (N_10678,N_10078,N_10011);
or U10679 (N_10679,N_10268,N_10420);
or U10680 (N_10680,N_10291,N_10125);
or U10681 (N_10681,N_10186,N_10255);
or U10682 (N_10682,N_10150,N_10073);
nor U10683 (N_10683,N_10218,N_10334);
or U10684 (N_10684,N_10040,N_10321);
nand U10685 (N_10685,N_10166,N_10264);
and U10686 (N_10686,N_10133,N_10189);
nor U10687 (N_10687,N_10487,N_10227);
nand U10688 (N_10688,N_10017,N_10235);
or U10689 (N_10689,N_10440,N_10375);
and U10690 (N_10690,N_10027,N_10023);
and U10691 (N_10691,N_10075,N_10491);
nand U10692 (N_10692,N_10302,N_10225);
nor U10693 (N_10693,N_10152,N_10245);
or U10694 (N_10694,N_10241,N_10494);
and U10695 (N_10695,N_10195,N_10260);
nand U10696 (N_10696,N_10357,N_10319);
xnor U10697 (N_10697,N_10286,N_10101);
nor U10698 (N_10698,N_10221,N_10143);
nor U10699 (N_10699,N_10051,N_10057);
nand U10700 (N_10700,N_10187,N_10382);
xnor U10701 (N_10701,N_10343,N_10485);
nor U10702 (N_10702,N_10277,N_10400);
and U10703 (N_10703,N_10208,N_10256);
and U10704 (N_10704,N_10482,N_10492);
nand U10705 (N_10705,N_10205,N_10124);
nand U10706 (N_10706,N_10434,N_10496);
xor U10707 (N_10707,N_10415,N_10431);
or U10708 (N_10708,N_10324,N_10350);
xnor U10709 (N_10709,N_10279,N_10016);
nand U10710 (N_10710,N_10292,N_10438);
and U10711 (N_10711,N_10215,N_10024);
nor U10712 (N_10712,N_10083,N_10136);
nor U10713 (N_10713,N_10322,N_10351);
nand U10714 (N_10714,N_10457,N_10384);
nor U10715 (N_10715,N_10244,N_10355);
nor U10716 (N_10716,N_10174,N_10250);
nand U10717 (N_10717,N_10007,N_10113);
xor U10718 (N_10718,N_10316,N_10406);
or U10719 (N_10719,N_10108,N_10163);
nor U10720 (N_10720,N_10422,N_10058);
xor U10721 (N_10721,N_10184,N_10216);
and U10722 (N_10722,N_10473,N_10096);
or U10723 (N_10723,N_10008,N_10097);
xnor U10724 (N_10724,N_10407,N_10142);
nor U10725 (N_10725,N_10002,N_10364);
nand U10726 (N_10726,N_10190,N_10220);
or U10727 (N_10727,N_10403,N_10263);
nand U10728 (N_10728,N_10329,N_10239);
and U10729 (N_10729,N_10346,N_10266);
or U10730 (N_10730,N_10234,N_10084);
nor U10731 (N_10731,N_10025,N_10416);
and U10732 (N_10732,N_10128,N_10064);
or U10733 (N_10733,N_10130,N_10497);
nor U10734 (N_10734,N_10192,N_10481);
nand U10735 (N_10735,N_10252,N_10202);
nor U10736 (N_10736,N_10098,N_10240);
nand U10737 (N_10737,N_10068,N_10156);
xor U10738 (N_10738,N_10099,N_10488);
nand U10739 (N_10739,N_10437,N_10105);
xnor U10740 (N_10740,N_10493,N_10283);
nand U10741 (N_10741,N_10003,N_10293);
and U10742 (N_10742,N_10325,N_10100);
nor U10743 (N_10743,N_10214,N_10363);
nor U10744 (N_10744,N_10296,N_10347);
or U10745 (N_10745,N_10242,N_10088);
or U10746 (N_10746,N_10000,N_10294);
and U10747 (N_10747,N_10444,N_10154);
and U10748 (N_10748,N_10376,N_10339);
xnor U10749 (N_10749,N_10300,N_10106);
nand U10750 (N_10750,N_10408,N_10211);
or U10751 (N_10751,N_10324,N_10111);
and U10752 (N_10752,N_10030,N_10377);
or U10753 (N_10753,N_10368,N_10420);
or U10754 (N_10754,N_10297,N_10026);
or U10755 (N_10755,N_10180,N_10440);
and U10756 (N_10756,N_10035,N_10309);
or U10757 (N_10757,N_10151,N_10470);
nor U10758 (N_10758,N_10473,N_10009);
nand U10759 (N_10759,N_10444,N_10176);
or U10760 (N_10760,N_10453,N_10212);
nand U10761 (N_10761,N_10115,N_10364);
or U10762 (N_10762,N_10178,N_10075);
nand U10763 (N_10763,N_10471,N_10495);
nor U10764 (N_10764,N_10448,N_10110);
nor U10765 (N_10765,N_10203,N_10466);
and U10766 (N_10766,N_10091,N_10107);
nor U10767 (N_10767,N_10270,N_10279);
nor U10768 (N_10768,N_10492,N_10324);
nand U10769 (N_10769,N_10267,N_10418);
nor U10770 (N_10770,N_10348,N_10317);
or U10771 (N_10771,N_10132,N_10436);
nor U10772 (N_10772,N_10302,N_10079);
xnor U10773 (N_10773,N_10032,N_10192);
xor U10774 (N_10774,N_10360,N_10037);
or U10775 (N_10775,N_10131,N_10205);
or U10776 (N_10776,N_10488,N_10269);
or U10777 (N_10777,N_10286,N_10141);
or U10778 (N_10778,N_10056,N_10124);
or U10779 (N_10779,N_10455,N_10444);
and U10780 (N_10780,N_10281,N_10260);
nand U10781 (N_10781,N_10136,N_10034);
and U10782 (N_10782,N_10010,N_10365);
and U10783 (N_10783,N_10376,N_10143);
nor U10784 (N_10784,N_10076,N_10086);
nand U10785 (N_10785,N_10273,N_10000);
or U10786 (N_10786,N_10348,N_10158);
nand U10787 (N_10787,N_10444,N_10315);
and U10788 (N_10788,N_10312,N_10243);
and U10789 (N_10789,N_10475,N_10280);
and U10790 (N_10790,N_10455,N_10274);
xnor U10791 (N_10791,N_10227,N_10207);
and U10792 (N_10792,N_10414,N_10347);
nand U10793 (N_10793,N_10287,N_10369);
xor U10794 (N_10794,N_10007,N_10189);
xor U10795 (N_10795,N_10306,N_10418);
or U10796 (N_10796,N_10299,N_10248);
and U10797 (N_10797,N_10416,N_10074);
nand U10798 (N_10798,N_10372,N_10496);
or U10799 (N_10799,N_10215,N_10197);
nand U10800 (N_10800,N_10441,N_10287);
and U10801 (N_10801,N_10322,N_10479);
or U10802 (N_10802,N_10352,N_10156);
or U10803 (N_10803,N_10041,N_10232);
or U10804 (N_10804,N_10315,N_10098);
and U10805 (N_10805,N_10267,N_10285);
xor U10806 (N_10806,N_10138,N_10284);
or U10807 (N_10807,N_10350,N_10298);
nand U10808 (N_10808,N_10050,N_10278);
and U10809 (N_10809,N_10082,N_10263);
nor U10810 (N_10810,N_10498,N_10046);
nand U10811 (N_10811,N_10263,N_10201);
nor U10812 (N_10812,N_10428,N_10254);
nand U10813 (N_10813,N_10108,N_10348);
and U10814 (N_10814,N_10332,N_10183);
xor U10815 (N_10815,N_10242,N_10066);
nand U10816 (N_10816,N_10397,N_10256);
and U10817 (N_10817,N_10256,N_10273);
or U10818 (N_10818,N_10240,N_10257);
nand U10819 (N_10819,N_10497,N_10272);
nor U10820 (N_10820,N_10428,N_10094);
or U10821 (N_10821,N_10072,N_10124);
and U10822 (N_10822,N_10477,N_10443);
or U10823 (N_10823,N_10141,N_10275);
and U10824 (N_10824,N_10222,N_10260);
or U10825 (N_10825,N_10260,N_10427);
or U10826 (N_10826,N_10232,N_10446);
or U10827 (N_10827,N_10079,N_10246);
or U10828 (N_10828,N_10124,N_10178);
nor U10829 (N_10829,N_10167,N_10115);
nand U10830 (N_10830,N_10467,N_10088);
nor U10831 (N_10831,N_10229,N_10449);
and U10832 (N_10832,N_10330,N_10013);
or U10833 (N_10833,N_10148,N_10132);
nor U10834 (N_10834,N_10028,N_10357);
or U10835 (N_10835,N_10299,N_10114);
or U10836 (N_10836,N_10035,N_10010);
and U10837 (N_10837,N_10497,N_10477);
and U10838 (N_10838,N_10253,N_10197);
nand U10839 (N_10839,N_10158,N_10146);
nand U10840 (N_10840,N_10269,N_10358);
xor U10841 (N_10841,N_10495,N_10118);
or U10842 (N_10842,N_10322,N_10086);
xor U10843 (N_10843,N_10151,N_10112);
xnor U10844 (N_10844,N_10147,N_10261);
nand U10845 (N_10845,N_10447,N_10287);
nand U10846 (N_10846,N_10208,N_10292);
or U10847 (N_10847,N_10381,N_10247);
nand U10848 (N_10848,N_10440,N_10412);
or U10849 (N_10849,N_10091,N_10198);
nand U10850 (N_10850,N_10438,N_10214);
nor U10851 (N_10851,N_10036,N_10262);
or U10852 (N_10852,N_10432,N_10423);
and U10853 (N_10853,N_10096,N_10493);
nor U10854 (N_10854,N_10449,N_10191);
or U10855 (N_10855,N_10386,N_10304);
or U10856 (N_10856,N_10000,N_10006);
or U10857 (N_10857,N_10171,N_10129);
nand U10858 (N_10858,N_10173,N_10022);
or U10859 (N_10859,N_10376,N_10052);
and U10860 (N_10860,N_10471,N_10443);
nor U10861 (N_10861,N_10316,N_10045);
and U10862 (N_10862,N_10389,N_10322);
or U10863 (N_10863,N_10044,N_10390);
nor U10864 (N_10864,N_10475,N_10222);
nor U10865 (N_10865,N_10081,N_10314);
nand U10866 (N_10866,N_10491,N_10294);
xnor U10867 (N_10867,N_10034,N_10383);
and U10868 (N_10868,N_10194,N_10096);
nand U10869 (N_10869,N_10120,N_10347);
or U10870 (N_10870,N_10183,N_10309);
nor U10871 (N_10871,N_10303,N_10085);
xor U10872 (N_10872,N_10151,N_10487);
nand U10873 (N_10873,N_10203,N_10125);
nand U10874 (N_10874,N_10198,N_10245);
nor U10875 (N_10875,N_10087,N_10482);
and U10876 (N_10876,N_10340,N_10483);
nand U10877 (N_10877,N_10110,N_10001);
or U10878 (N_10878,N_10259,N_10453);
and U10879 (N_10879,N_10030,N_10109);
or U10880 (N_10880,N_10430,N_10045);
and U10881 (N_10881,N_10123,N_10348);
nor U10882 (N_10882,N_10227,N_10040);
or U10883 (N_10883,N_10350,N_10432);
or U10884 (N_10884,N_10317,N_10485);
nor U10885 (N_10885,N_10414,N_10251);
and U10886 (N_10886,N_10075,N_10399);
nor U10887 (N_10887,N_10256,N_10357);
nand U10888 (N_10888,N_10288,N_10087);
or U10889 (N_10889,N_10396,N_10313);
or U10890 (N_10890,N_10343,N_10325);
nor U10891 (N_10891,N_10184,N_10053);
nand U10892 (N_10892,N_10161,N_10072);
xnor U10893 (N_10893,N_10447,N_10051);
nand U10894 (N_10894,N_10407,N_10120);
nand U10895 (N_10895,N_10270,N_10368);
nor U10896 (N_10896,N_10040,N_10443);
and U10897 (N_10897,N_10199,N_10031);
nor U10898 (N_10898,N_10303,N_10477);
and U10899 (N_10899,N_10022,N_10216);
nor U10900 (N_10900,N_10325,N_10194);
nor U10901 (N_10901,N_10224,N_10257);
nand U10902 (N_10902,N_10426,N_10289);
or U10903 (N_10903,N_10460,N_10057);
nor U10904 (N_10904,N_10280,N_10065);
and U10905 (N_10905,N_10372,N_10257);
and U10906 (N_10906,N_10127,N_10170);
xnor U10907 (N_10907,N_10045,N_10248);
and U10908 (N_10908,N_10292,N_10190);
nor U10909 (N_10909,N_10180,N_10306);
nand U10910 (N_10910,N_10163,N_10297);
nand U10911 (N_10911,N_10100,N_10208);
nor U10912 (N_10912,N_10070,N_10490);
and U10913 (N_10913,N_10195,N_10404);
and U10914 (N_10914,N_10263,N_10495);
and U10915 (N_10915,N_10138,N_10100);
or U10916 (N_10916,N_10493,N_10126);
or U10917 (N_10917,N_10331,N_10403);
and U10918 (N_10918,N_10114,N_10359);
or U10919 (N_10919,N_10397,N_10072);
and U10920 (N_10920,N_10194,N_10238);
nor U10921 (N_10921,N_10066,N_10263);
or U10922 (N_10922,N_10326,N_10451);
and U10923 (N_10923,N_10011,N_10412);
and U10924 (N_10924,N_10492,N_10348);
nand U10925 (N_10925,N_10203,N_10205);
and U10926 (N_10926,N_10401,N_10193);
nand U10927 (N_10927,N_10148,N_10442);
or U10928 (N_10928,N_10051,N_10312);
or U10929 (N_10929,N_10087,N_10051);
and U10930 (N_10930,N_10469,N_10342);
or U10931 (N_10931,N_10395,N_10133);
and U10932 (N_10932,N_10343,N_10229);
nand U10933 (N_10933,N_10217,N_10489);
nand U10934 (N_10934,N_10018,N_10024);
and U10935 (N_10935,N_10012,N_10438);
nand U10936 (N_10936,N_10041,N_10056);
nand U10937 (N_10937,N_10024,N_10099);
nand U10938 (N_10938,N_10056,N_10289);
or U10939 (N_10939,N_10323,N_10315);
and U10940 (N_10940,N_10240,N_10061);
xor U10941 (N_10941,N_10012,N_10131);
and U10942 (N_10942,N_10162,N_10358);
nand U10943 (N_10943,N_10192,N_10328);
nand U10944 (N_10944,N_10148,N_10283);
nor U10945 (N_10945,N_10404,N_10198);
nor U10946 (N_10946,N_10272,N_10201);
and U10947 (N_10947,N_10102,N_10131);
nand U10948 (N_10948,N_10254,N_10234);
nand U10949 (N_10949,N_10164,N_10182);
and U10950 (N_10950,N_10355,N_10100);
xnor U10951 (N_10951,N_10478,N_10404);
nor U10952 (N_10952,N_10319,N_10267);
or U10953 (N_10953,N_10397,N_10010);
or U10954 (N_10954,N_10325,N_10411);
nor U10955 (N_10955,N_10085,N_10290);
or U10956 (N_10956,N_10398,N_10003);
or U10957 (N_10957,N_10024,N_10148);
nand U10958 (N_10958,N_10117,N_10363);
and U10959 (N_10959,N_10366,N_10406);
or U10960 (N_10960,N_10229,N_10135);
or U10961 (N_10961,N_10011,N_10319);
nand U10962 (N_10962,N_10446,N_10182);
nand U10963 (N_10963,N_10065,N_10159);
nor U10964 (N_10964,N_10201,N_10482);
or U10965 (N_10965,N_10276,N_10319);
or U10966 (N_10966,N_10105,N_10035);
xnor U10967 (N_10967,N_10185,N_10097);
or U10968 (N_10968,N_10205,N_10223);
and U10969 (N_10969,N_10043,N_10094);
or U10970 (N_10970,N_10000,N_10454);
nor U10971 (N_10971,N_10173,N_10149);
nor U10972 (N_10972,N_10402,N_10422);
and U10973 (N_10973,N_10183,N_10174);
nor U10974 (N_10974,N_10332,N_10329);
and U10975 (N_10975,N_10306,N_10173);
xnor U10976 (N_10976,N_10136,N_10358);
nand U10977 (N_10977,N_10157,N_10138);
and U10978 (N_10978,N_10270,N_10196);
or U10979 (N_10979,N_10231,N_10343);
nor U10980 (N_10980,N_10194,N_10009);
nor U10981 (N_10981,N_10092,N_10093);
nor U10982 (N_10982,N_10004,N_10032);
nand U10983 (N_10983,N_10366,N_10312);
or U10984 (N_10984,N_10389,N_10371);
nand U10985 (N_10985,N_10409,N_10208);
and U10986 (N_10986,N_10119,N_10029);
and U10987 (N_10987,N_10285,N_10061);
and U10988 (N_10988,N_10217,N_10284);
nor U10989 (N_10989,N_10295,N_10154);
or U10990 (N_10990,N_10182,N_10058);
or U10991 (N_10991,N_10299,N_10169);
xnor U10992 (N_10992,N_10115,N_10283);
and U10993 (N_10993,N_10018,N_10274);
nor U10994 (N_10994,N_10165,N_10409);
and U10995 (N_10995,N_10021,N_10173);
or U10996 (N_10996,N_10302,N_10494);
nor U10997 (N_10997,N_10303,N_10021);
or U10998 (N_10998,N_10241,N_10210);
nor U10999 (N_10999,N_10191,N_10217);
and U11000 (N_11000,N_10879,N_10768);
and U11001 (N_11001,N_10713,N_10782);
nor U11002 (N_11002,N_10588,N_10911);
or U11003 (N_11003,N_10603,N_10545);
nor U11004 (N_11004,N_10549,N_10752);
and U11005 (N_11005,N_10820,N_10643);
xor U11006 (N_11006,N_10834,N_10716);
and U11007 (N_11007,N_10662,N_10825);
or U11008 (N_11008,N_10905,N_10990);
and U11009 (N_11009,N_10998,N_10796);
and U11010 (N_11010,N_10778,N_10684);
nor U11011 (N_11011,N_10519,N_10712);
nor U11012 (N_11012,N_10851,N_10822);
nand U11013 (N_11013,N_10528,N_10988);
nor U11014 (N_11014,N_10772,N_10582);
nor U11015 (N_11015,N_10849,N_10722);
and U11016 (N_11016,N_10762,N_10610);
and U11017 (N_11017,N_10974,N_10696);
and U11018 (N_11018,N_10885,N_10534);
nand U11019 (N_11019,N_10617,N_10732);
nand U11020 (N_11020,N_10649,N_10567);
nand U11021 (N_11021,N_10591,N_10624);
or U11022 (N_11022,N_10823,N_10593);
nor U11023 (N_11023,N_10886,N_10787);
and U11024 (N_11024,N_10869,N_10951);
nor U11025 (N_11025,N_10854,N_10580);
or U11026 (N_11026,N_10780,N_10745);
or U11027 (N_11027,N_10890,N_10570);
or U11028 (N_11028,N_10996,N_10831);
nand U11029 (N_11029,N_10868,N_10571);
and U11030 (N_11030,N_10714,N_10961);
nand U11031 (N_11031,N_10880,N_10948);
nor U11032 (N_11032,N_10638,N_10850);
and U11033 (N_11033,N_10866,N_10677);
nand U11034 (N_11034,N_10815,N_10829);
nor U11035 (N_11035,N_10864,N_10958);
or U11036 (N_11036,N_10839,N_10569);
or U11037 (N_11037,N_10992,N_10856);
nor U11038 (N_11038,N_10666,N_10899);
and U11039 (N_11039,N_10691,N_10679);
nor U11040 (N_11040,N_10784,N_10817);
and U11041 (N_11041,N_10819,N_10932);
nor U11042 (N_11042,N_10941,N_10555);
or U11043 (N_11043,N_10969,N_10604);
and U11044 (N_11044,N_10709,N_10740);
nor U11045 (N_11045,N_10997,N_10967);
nand U11046 (N_11046,N_10858,N_10922);
nor U11047 (N_11047,N_10509,N_10629);
nand U11048 (N_11048,N_10575,N_10667);
and U11049 (N_11049,N_10781,N_10611);
nand U11050 (N_11050,N_10682,N_10900);
xor U11051 (N_11051,N_10789,N_10689);
nand U11052 (N_11052,N_10701,N_10559);
and U11053 (N_11053,N_10830,N_10908);
or U11054 (N_11054,N_10517,N_10779);
nand U11055 (N_11055,N_10982,N_10862);
nand U11056 (N_11056,N_10635,N_10926);
xnor U11057 (N_11057,N_10927,N_10945);
or U11058 (N_11058,N_10512,N_10706);
nor U11059 (N_11059,N_10814,N_10672);
or U11060 (N_11060,N_10589,N_10760);
nor U11061 (N_11061,N_10553,N_10560);
nand U11062 (N_11062,N_10970,N_10770);
or U11063 (N_11063,N_10572,N_10953);
nand U11064 (N_11064,N_10964,N_10743);
nor U11065 (N_11065,N_10674,N_10594);
or U11066 (N_11066,N_10525,N_10888);
or U11067 (N_11067,N_10720,N_10749);
or U11068 (N_11068,N_10600,N_10565);
or U11069 (N_11069,N_10811,N_10526);
and U11070 (N_11070,N_10915,N_10965);
xnor U11071 (N_11071,N_10737,N_10514);
nor U11072 (N_11072,N_10901,N_10937);
nand U11073 (N_11073,N_10744,N_10801);
or U11074 (N_11074,N_10808,N_10524);
or U11075 (N_11075,N_10765,N_10841);
nand U11076 (N_11076,N_10710,N_10622);
and U11077 (N_11077,N_10754,N_10651);
nor U11078 (N_11078,N_10757,N_10826);
and U11079 (N_11079,N_10904,N_10898);
or U11080 (N_11080,N_10876,N_10935);
nand U11081 (N_11081,N_10641,N_10619);
and U11082 (N_11082,N_10753,N_10954);
nor U11083 (N_11083,N_10664,N_10746);
nand U11084 (N_11084,N_10980,N_10767);
or U11085 (N_11085,N_10747,N_10551);
nand U11086 (N_11086,N_10597,N_10596);
or U11087 (N_11087,N_10505,N_10612);
xnor U11088 (N_11088,N_10683,N_10907);
nand U11089 (N_11089,N_10521,N_10835);
or U11090 (N_11090,N_10618,N_10632);
and U11091 (N_11091,N_10605,N_10718);
or U11092 (N_11092,N_10942,N_10522);
and U11093 (N_11093,N_10538,N_10906);
and U11094 (N_11094,N_10883,N_10946);
or U11095 (N_11095,N_10995,N_10693);
and U11096 (N_11096,N_10581,N_10535);
and U11097 (N_11097,N_10697,N_10584);
and U11098 (N_11098,N_10668,N_10620);
nand U11099 (N_11099,N_10533,N_10550);
xnor U11100 (N_11100,N_10903,N_10595);
nand U11101 (N_11101,N_10977,N_10733);
and U11102 (N_11102,N_10585,N_10707);
nand U11103 (N_11103,N_10931,N_10750);
nor U11104 (N_11104,N_10985,N_10962);
xnor U11105 (N_11105,N_10810,N_10928);
and U11106 (N_11106,N_10936,N_10676);
and U11107 (N_11107,N_10968,N_10654);
nand U11108 (N_11108,N_10783,N_10529);
xnor U11109 (N_11109,N_10598,N_10671);
and U11110 (N_11110,N_10918,N_10731);
or U11111 (N_11111,N_10503,N_10518);
or U11112 (N_11112,N_10748,N_10592);
and U11113 (N_11113,N_10775,N_10633);
or U11114 (N_11114,N_10540,N_10981);
nand U11115 (N_11115,N_10914,N_10910);
nand U11116 (N_11116,N_10842,N_10944);
nor U11117 (N_11117,N_10756,N_10956);
and U11118 (N_11118,N_10728,N_10766);
nand U11119 (N_11119,N_10681,N_10871);
and U11120 (N_11120,N_10828,N_10501);
xor U11121 (N_11121,N_10566,N_10788);
nor U11122 (N_11122,N_10836,N_10516);
and U11123 (N_11123,N_10827,N_10934);
xor U11124 (N_11124,N_10721,N_10795);
or U11125 (N_11125,N_10639,N_10943);
nand U11126 (N_11126,N_10777,N_10507);
xnor U11127 (N_11127,N_10563,N_10530);
nand U11128 (N_11128,N_10705,N_10719);
nor U11129 (N_11129,N_10863,N_10602);
nand U11130 (N_11130,N_10902,N_10812);
nand U11131 (N_11131,N_10878,N_10544);
or U11132 (N_11132,N_10729,N_10966);
nor U11133 (N_11133,N_10993,N_10657);
or U11134 (N_11134,N_10930,N_10608);
and U11135 (N_11135,N_10573,N_10776);
nor U11136 (N_11136,N_10755,N_10925);
nand U11137 (N_11137,N_10665,N_10955);
nor U11138 (N_11138,N_10794,N_10735);
or U11139 (N_11139,N_10870,N_10882);
nor U11140 (N_11140,N_10813,N_10807);
or U11141 (N_11141,N_10785,N_10655);
or U11142 (N_11142,N_10558,N_10537);
nand U11143 (N_11143,N_10950,N_10646);
nand U11144 (N_11144,N_10973,N_10579);
nor U11145 (N_11145,N_10536,N_10847);
or U11146 (N_11146,N_10939,N_10508);
or U11147 (N_11147,N_10730,N_10855);
or U11148 (N_11148,N_10601,N_10702);
and U11149 (N_11149,N_10647,N_10527);
nor U11150 (N_11150,N_10896,N_10859);
nor U11151 (N_11151,N_10699,N_10874);
or U11152 (N_11152,N_10889,N_10803);
nand U11153 (N_11153,N_10848,N_10727);
nand U11154 (N_11154,N_10895,N_10546);
nor U11155 (N_11155,N_10894,N_10725);
and U11156 (N_11156,N_10845,N_10806);
and U11157 (N_11157,N_10816,N_10846);
or U11158 (N_11158,N_10541,N_10947);
nor U11159 (N_11159,N_10832,N_10989);
or U11160 (N_11160,N_10644,N_10615);
xor U11161 (N_11161,N_10704,N_10698);
and U11162 (N_11162,N_10574,N_10642);
or U11163 (N_11163,N_10645,N_10893);
nor U11164 (N_11164,N_10987,N_10675);
nor U11165 (N_11165,N_10510,N_10873);
or U11166 (N_11166,N_10991,N_10673);
nor U11167 (N_11167,N_10769,N_10532);
nor U11168 (N_11168,N_10653,N_10833);
nand U11169 (N_11169,N_10715,N_10726);
xnor U11170 (N_11170,N_10938,N_10628);
and U11171 (N_11171,N_10506,N_10837);
xnor U11172 (N_11172,N_10625,N_10636);
and U11173 (N_11173,N_10627,N_10686);
nand U11174 (N_11174,N_10844,N_10921);
nand U11175 (N_11175,N_10798,N_10678);
nand U11176 (N_11176,N_10515,N_10542);
or U11177 (N_11177,N_10568,N_10804);
nor U11178 (N_11178,N_10652,N_10786);
nor U11179 (N_11179,N_10658,N_10564);
xor U11180 (N_11180,N_10929,N_10669);
or U11181 (N_11181,N_10790,N_10650);
xor U11182 (N_11182,N_10680,N_10821);
or U11183 (N_11183,N_10917,N_10614);
and U11184 (N_11184,N_10738,N_10771);
or U11185 (N_11185,N_10703,N_10661);
or U11186 (N_11186,N_10984,N_10659);
nor U11187 (N_11187,N_10999,N_10971);
nand U11188 (N_11188,N_10861,N_10975);
or U11189 (N_11189,N_10791,N_10590);
nor U11190 (N_11190,N_10687,N_10513);
nor U11191 (N_11191,N_10578,N_10865);
nand U11192 (N_11192,N_10741,N_10663);
nor U11193 (N_11193,N_10960,N_10723);
and U11194 (N_11194,N_10805,N_10875);
nand U11195 (N_11195,N_10979,N_10576);
and U11196 (N_11196,N_10670,N_10739);
nor U11197 (N_11197,N_10852,N_10891);
and U11198 (N_11198,N_10761,N_10758);
nor U11199 (N_11199,N_10773,N_10857);
nor U11200 (N_11200,N_10976,N_10793);
nor U11201 (N_11201,N_10872,N_10708);
and U11202 (N_11202,N_10587,N_10561);
or U11203 (N_11203,N_10734,N_10923);
or U11204 (N_11204,N_10774,N_10609);
or U11205 (N_11205,N_10531,N_10809);
or U11206 (N_11206,N_10892,N_10940);
nor U11207 (N_11207,N_10759,N_10640);
nand U11208 (N_11208,N_10690,N_10952);
nor U11209 (N_11209,N_10724,N_10924);
xor U11210 (N_11210,N_10623,N_10556);
or U11211 (N_11211,N_10963,N_10557);
nor U11212 (N_11212,N_10621,N_10949);
or U11213 (N_11213,N_10539,N_10887);
or U11214 (N_11214,N_10656,N_10577);
nor U11215 (N_11215,N_10500,N_10606);
nand U11216 (N_11216,N_10881,N_10957);
nor U11217 (N_11217,N_10607,N_10978);
xor U11218 (N_11218,N_10838,N_10983);
nor U11219 (N_11219,N_10867,N_10511);
nor U11220 (N_11220,N_10751,N_10916);
nand U11221 (N_11221,N_10994,N_10764);
and U11222 (N_11222,N_10843,N_10692);
nor U11223 (N_11223,N_10799,N_10797);
or U11224 (N_11224,N_10685,N_10933);
xnor U11225 (N_11225,N_10616,N_10913);
and U11226 (N_11226,N_10972,N_10800);
nand U11227 (N_11227,N_10554,N_10688);
and U11228 (N_11228,N_10717,N_10502);
or U11229 (N_11229,N_10634,N_10562);
nand U11230 (N_11230,N_10630,N_10631);
or U11231 (N_11231,N_10711,N_10543);
and U11232 (N_11232,N_10613,N_10648);
nor U11233 (N_11233,N_10860,N_10504);
or U11234 (N_11234,N_10695,N_10920);
nor U11235 (N_11235,N_10986,N_10548);
nand U11236 (N_11236,N_10818,N_10840);
or U11237 (N_11237,N_10909,N_10523);
or U11238 (N_11238,N_10599,N_10586);
or U11239 (N_11239,N_10552,N_10877);
or U11240 (N_11240,N_10919,N_10626);
nand U11241 (N_11241,N_10792,N_10742);
and U11242 (N_11242,N_10763,N_10736);
nand U11243 (N_11243,N_10824,N_10884);
nor U11244 (N_11244,N_10802,N_10547);
nor U11245 (N_11245,N_10897,N_10912);
or U11246 (N_11246,N_10660,N_10700);
nor U11247 (N_11247,N_10520,N_10637);
or U11248 (N_11248,N_10694,N_10959);
or U11249 (N_11249,N_10583,N_10853);
and U11250 (N_11250,N_10803,N_10684);
nor U11251 (N_11251,N_10681,N_10842);
and U11252 (N_11252,N_10998,N_10928);
or U11253 (N_11253,N_10657,N_10839);
and U11254 (N_11254,N_10983,N_10926);
nand U11255 (N_11255,N_10978,N_10872);
nor U11256 (N_11256,N_10834,N_10504);
or U11257 (N_11257,N_10681,N_10727);
and U11258 (N_11258,N_10650,N_10675);
and U11259 (N_11259,N_10835,N_10971);
xor U11260 (N_11260,N_10827,N_10525);
xor U11261 (N_11261,N_10835,N_10923);
nand U11262 (N_11262,N_10938,N_10663);
nor U11263 (N_11263,N_10881,N_10960);
and U11264 (N_11264,N_10740,N_10757);
nor U11265 (N_11265,N_10836,N_10753);
nor U11266 (N_11266,N_10871,N_10572);
xnor U11267 (N_11267,N_10632,N_10920);
nor U11268 (N_11268,N_10641,N_10837);
nor U11269 (N_11269,N_10947,N_10951);
and U11270 (N_11270,N_10629,N_10647);
and U11271 (N_11271,N_10753,N_10546);
nor U11272 (N_11272,N_10861,N_10658);
and U11273 (N_11273,N_10554,N_10637);
or U11274 (N_11274,N_10756,N_10571);
and U11275 (N_11275,N_10969,N_10768);
or U11276 (N_11276,N_10537,N_10651);
nand U11277 (N_11277,N_10988,N_10540);
or U11278 (N_11278,N_10967,N_10549);
xnor U11279 (N_11279,N_10503,N_10788);
and U11280 (N_11280,N_10554,N_10901);
and U11281 (N_11281,N_10652,N_10805);
nor U11282 (N_11282,N_10606,N_10657);
or U11283 (N_11283,N_10909,N_10916);
nand U11284 (N_11284,N_10969,N_10756);
and U11285 (N_11285,N_10894,N_10505);
nand U11286 (N_11286,N_10691,N_10979);
and U11287 (N_11287,N_10738,N_10601);
and U11288 (N_11288,N_10670,N_10563);
and U11289 (N_11289,N_10591,N_10625);
nor U11290 (N_11290,N_10826,N_10625);
and U11291 (N_11291,N_10782,N_10961);
or U11292 (N_11292,N_10986,N_10781);
xnor U11293 (N_11293,N_10602,N_10929);
and U11294 (N_11294,N_10960,N_10925);
nand U11295 (N_11295,N_10946,N_10993);
or U11296 (N_11296,N_10669,N_10657);
nor U11297 (N_11297,N_10623,N_10942);
and U11298 (N_11298,N_10918,N_10867);
nor U11299 (N_11299,N_10653,N_10585);
or U11300 (N_11300,N_10786,N_10934);
nand U11301 (N_11301,N_10502,N_10955);
or U11302 (N_11302,N_10975,N_10788);
nor U11303 (N_11303,N_10609,N_10672);
xor U11304 (N_11304,N_10775,N_10598);
nand U11305 (N_11305,N_10912,N_10615);
or U11306 (N_11306,N_10966,N_10877);
and U11307 (N_11307,N_10741,N_10553);
and U11308 (N_11308,N_10759,N_10887);
nand U11309 (N_11309,N_10641,N_10513);
or U11310 (N_11310,N_10796,N_10849);
and U11311 (N_11311,N_10894,N_10977);
xnor U11312 (N_11312,N_10904,N_10572);
and U11313 (N_11313,N_10758,N_10983);
nor U11314 (N_11314,N_10803,N_10814);
nand U11315 (N_11315,N_10903,N_10611);
nand U11316 (N_11316,N_10681,N_10911);
nand U11317 (N_11317,N_10785,N_10848);
and U11318 (N_11318,N_10964,N_10669);
nor U11319 (N_11319,N_10569,N_10739);
and U11320 (N_11320,N_10547,N_10953);
and U11321 (N_11321,N_10897,N_10515);
nor U11322 (N_11322,N_10927,N_10685);
and U11323 (N_11323,N_10917,N_10662);
nor U11324 (N_11324,N_10741,N_10820);
nor U11325 (N_11325,N_10520,N_10950);
nand U11326 (N_11326,N_10651,N_10822);
nand U11327 (N_11327,N_10810,N_10796);
or U11328 (N_11328,N_10606,N_10633);
and U11329 (N_11329,N_10509,N_10598);
nand U11330 (N_11330,N_10708,N_10729);
or U11331 (N_11331,N_10882,N_10946);
nor U11332 (N_11332,N_10673,N_10805);
nand U11333 (N_11333,N_10996,N_10588);
nand U11334 (N_11334,N_10722,N_10506);
and U11335 (N_11335,N_10941,N_10764);
xor U11336 (N_11336,N_10557,N_10799);
nor U11337 (N_11337,N_10994,N_10671);
nand U11338 (N_11338,N_10854,N_10976);
xnor U11339 (N_11339,N_10840,N_10730);
nor U11340 (N_11340,N_10781,N_10559);
or U11341 (N_11341,N_10878,N_10564);
nand U11342 (N_11342,N_10918,N_10750);
nor U11343 (N_11343,N_10866,N_10650);
and U11344 (N_11344,N_10593,N_10808);
nand U11345 (N_11345,N_10690,N_10560);
nor U11346 (N_11346,N_10804,N_10653);
or U11347 (N_11347,N_10715,N_10631);
nor U11348 (N_11348,N_10636,N_10782);
nand U11349 (N_11349,N_10675,N_10917);
nand U11350 (N_11350,N_10938,N_10742);
and U11351 (N_11351,N_10876,N_10847);
or U11352 (N_11352,N_10603,N_10988);
and U11353 (N_11353,N_10574,N_10698);
and U11354 (N_11354,N_10963,N_10991);
and U11355 (N_11355,N_10524,N_10899);
and U11356 (N_11356,N_10920,N_10743);
or U11357 (N_11357,N_10883,N_10595);
or U11358 (N_11358,N_10536,N_10854);
and U11359 (N_11359,N_10657,N_10789);
or U11360 (N_11360,N_10617,N_10678);
or U11361 (N_11361,N_10619,N_10778);
nor U11362 (N_11362,N_10956,N_10594);
nor U11363 (N_11363,N_10893,N_10797);
and U11364 (N_11364,N_10852,N_10955);
nand U11365 (N_11365,N_10623,N_10893);
nor U11366 (N_11366,N_10716,N_10562);
xor U11367 (N_11367,N_10731,N_10709);
and U11368 (N_11368,N_10509,N_10966);
or U11369 (N_11369,N_10846,N_10734);
and U11370 (N_11370,N_10619,N_10852);
nand U11371 (N_11371,N_10976,N_10612);
nor U11372 (N_11372,N_10961,N_10809);
or U11373 (N_11373,N_10594,N_10842);
xnor U11374 (N_11374,N_10976,N_10620);
nor U11375 (N_11375,N_10844,N_10890);
xnor U11376 (N_11376,N_10705,N_10937);
and U11377 (N_11377,N_10579,N_10573);
and U11378 (N_11378,N_10552,N_10952);
and U11379 (N_11379,N_10751,N_10938);
xor U11380 (N_11380,N_10810,N_10761);
or U11381 (N_11381,N_10785,N_10653);
or U11382 (N_11382,N_10783,N_10606);
nand U11383 (N_11383,N_10958,N_10651);
or U11384 (N_11384,N_10679,N_10817);
and U11385 (N_11385,N_10630,N_10999);
or U11386 (N_11386,N_10859,N_10506);
nand U11387 (N_11387,N_10777,N_10613);
or U11388 (N_11388,N_10964,N_10791);
nor U11389 (N_11389,N_10673,N_10758);
nor U11390 (N_11390,N_10857,N_10939);
nand U11391 (N_11391,N_10815,N_10509);
or U11392 (N_11392,N_10627,N_10583);
nor U11393 (N_11393,N_10701,N_10795);
and U11394 (N_11394,N_10558,N_10520);
and U11395 (N_11395,N_10981,N_10804);
nand U11396 (N_11396,N_10543,N_10902);
and U11397 (N_11397,N_10528,N_10713);
nand U11398 (N_11398,N_10559,N_10724);
nor U11399 (N_11399,N_10716,N_10550);
and U11400 (N_11400,N_10679,N_10999);
nand U11401 (N_11401,N_10785,N_10920);
or U11402 (N_11402,N_10795,N_10949);
and U11403 (N_11403,N_10821,N_10942);
or U11404 (N_11404,N_10999,N_10899);
nor U11405 (N_11405,N_10601,N_10898);
and U11406 (N_11406,N_10608,N_10977);
nand U11407 (N_11407,N_10605,N_10933);
and U11408 (N_11408,N_10591,N_10633);
nor U11409 (N_11409,N_10934,N_10979);
nand U11410 (N_11410,N_10703,N_10826);
nand U11411 (N_11411,N_10630,N_10845);
or U11412 (N_11412,N_10818,N_10772);
nand U11413 (N_11413,N_10948,N_10557);
and U11414 (N_11414,N_10961,N_10552);
or U11415 (N_11415,N_10778,N_10843);
nor U11416 (N_11416,N_10901,N_10851);
nor U11417 (N_11417,N_10883,N_10865);
xor U11418 (N_11418,N_10983,N_10746);
and U11419 (N_11419,N_10700,N_10913);
nand U11420 (N_11420,N_10828,N_10870);
nand U11421 (N_11421,N_10532,N_10690);
nor U11422 (N_11422,N_10842,N_10782);
and U11423 (N_11423,N_10998,N_10958);
nand U11424 (N_11424,N_10582,N_10723);
nand U11425 (N_11425,N_10632,N_10828);
nor U11426 (N_11426,N_10990,N_10851);
or U11427 (N_11427,N_10509,N_10567);
and U11428 (N_11428,N_10974,N_10822);
and U11429 (N_11429,N_10566,N_10501);
or U11430 (N_11430,N_10626,N_10805);
and U11431 (N_11431,N_10611,N_10615);
or U11432 (N_11432,N_10523,N_10800);
nand U11433 (N_11433,N_10991,N_10795);
or U11434 (N_11434,N_10503,N_10868);
xor U11435 (N_11435,N_10858,N_10925);
and U11436 (N_11436,N_10796,N_10974);
nor U11437 (N_11437,N_10555,N_10635);
xor U11438 (N_11438,N_10958,N_10948);
nand U11439 (N_11439,N_10683,N_10688);
nand U11440 (N_11440,N_10588,N_10940);
xnor U11441 (N_11441,N_10760,N_10609);
nand U11442 (N_11442,N_10640,N_10561);
nand U11443 (N_11443,N_10542,N_10776);
nor U11444 (N_11444,N_10799,N_10735);
nor U11445 (N_11445,N_10884,N_10872);
and U11446 (N_11446,N_10994,N_10737);
and U11447 (N_11447,N_10907,N_10951);
and U11448 (N_11448,N_10691,N_10891);
nor U11449 (N_11449,N_10684,N_10867);
nand U11450 (N_11450,N_10608,N_10599);
nand U11451 (N_11451,N_10944,N_10515);
and U11452 (N_11452,N_10880,N_10509);
nand U11453 (N_11453,N_10893,N_10798);
nor U11454 (N_11454,N_10989,N_10605);
and U11455 (N_11455,N_10790,N_10663);
nand U11456 (N_11456,N_10536,N_10866);
nand U11457 (N_11457,N_10595,N_10596);
or U11458 (N_11458,N_10870,N_10763);
xor U11459 (N_11459,N_10813,N_10542);
nand U11460 (N_11460,N_10945,N_10933);
and U11461 (N_11461,N_10533,N_10538);
and U11462 (N_11462,N_10813,N_10529);
and U11463 (N_11463,N_10616,N_10917);
and U11464 (N_11464,N_10564,N_10501);
nor U11465 (N_11465,N_10975,N_10717);
or U11466 (N_11466,N_10533,N_10520);
and U11467 (N_11467,N_10705,N_10824);
nor U11468 (N_11468,N_10804,N_10518);
or U11469 (N_11469,N_10634,N_10915);
and U11470 (N_11470,N_10674,N_10998);
or U11471 (N_11471,N_10618,N_10642);
and U11472 (N_11472,N_10901,N_10661);
nand U11473 (N_11473,N_10705,N_10559);
nor U11474 (N_11474,N_10509,N_10737);
or U11475 (N_11475,N_10858,N_10731);
nor U11476 (N_11476,N_10550,N_10528);
or U11477 (N_11477,N_10770,N_10913);
nor U11478 (N_11478,N_10972,N_10978);
xor U11479 (N_11479,N_10904,N_10775);
and U11480 (N_11480,N_10502,N_10875);
and U11481 (N_11481,N_10967,N_10874);
nor U11482 (N_11482,N_10668,N_10528);
nand U11483 (N_11483,N_10530,N_10983);
nand U11484 (N_11484,N_10828,N_10959);
or U11485 (N_11485,N_10687,N_10826);
or U11486 (N_11486,N_10765,N_10595);
nand U11487 (N_11487,N_10934,N_10689);
nor U11488 (N_11488,N_10667,N_10551);
and U11489 (N_11489,N_10622,N_10599);
and U11490 (N_11490,N_10618,N_10962);
and U11491 (N_11491,N_10514,N_10809);
and U11492 (N_11492,N_10610,N_10994);
nor U11493 (N_11493,N_10550,N_10581);
xor U11494 (N_11494,N_10540,N_10976);
or U11495 (N_11495,N_10867,N_10976);
or U11496 (N_11496,N_10760,N_10515);
nand U11497 (N_11497,N_10943,N_10798);
nand U11498 (N_11498,N_10581,N_10776);
nor U11499 (N_11499,N_10870,N_10545);
nand U11500 (N_11500,N_11434,N_11376);
and U11501 (N_11501,N_11446,N_11094);
or U11502 (N_11502,N_11475,N_11226);
or U11503 (N_11503,N_11123,N_11336);
nand U11504 (N_11504,N_11021,N_11172);
or U11505 (N_11505,N_11353,N_11445);
nand U11506 (N_11506,N_11058,N_11200);
nand U11507 (N_11507,N_11401,N_11231);
nand U11508 (N_11508,N_11195,N_11252);
nor U11509 (N_11509,N_11472,N_11375);
xor U11510 (N_11510,N_11428,N_11278);
or U11511 (N_11511,N_11121,N_11089);
and U11512 (N_11512,N_11176,N_11496);
nor U11513 (N_11513,N_11298,N_11189);
or U11514 (N_11514,N_11031,N_11419);
nand U11515 (N_11515,N_11431,N_11218);
nor U11516 (N_11516,N_11161,N_11270);
nor U11517 (N_11517,N_11104,N_11179);
nor U11518 (N_11518,N_11198,N_11114);
nand U11519 (N_11519,N_11448,N_11192);
or U11520 (N_11520,N_11396,N_11090);
xor U11521 (N_11521,N_11332,N_11438);
and U11522 (N_11522,N_11288,N_11394);
nor U11523 (N_11523,N_11211,N_11246);
xnor U11524 (N_11524,N_11112,N_11441);
nor U11525 (N_11525,N_11409,N_11284);
and U11526 (N_11526,N_11378,N_11232);
or U11527 (N_11527,N_11006,N_11249);
nor U11528 (N_11528,N_11407,N_11002);
and U11529 (N_11529,N_11437,N_11462);
and U11530 (N_11530,N_11064,N_11103);
or U11531 (N_11531,N_11042,N_11337);
or U11532 (N_11532,N_11073,N_11361);
nor U11533 (N_11533,N_11435,N_11456);
nand U11534 (N_11534,N_11120,N_11321);
or U11535 (N_11535,N_11291,N_11416);
and U11536 (N_11536,N_11254,N_11322);
nand U11537 (N_11537,N_11347,N_11142);
and U11538 (N_11538,N_11373,N_11034);
or U11539 (N_11539,N_11091,N_11381);
and U11540 (N_11540,N_11335,N_11293);
and U11541 (N_11541,N_11048,N_11477);
and U11542 (N_11542,N_11329,N_11476);
or U11543 (N_11543,N_11060,N_11194);
nand U11544 (N_11544,N_11129,N_11440);
nand U11545 (N_11545,N_11264,N_11449);
or U11546 (N_11546,N_11026,N_11460);
and U11547 (N_11547,N_11481,N_11097);
or U11548 (N_11548,N_11320,N_11013);
nor U11549 (N_11549,N_11338,N_11267);
nand U11550 (N_11550,N_11275,N_11011);
or U11551 (N_11551,N_11471,N_11492);
nor U11552 (N_11552,N_11110,N_11136);
or U11553 (N_11553,N_11432,N_11137);
or U11554 (N_11554,N_11271,N_11443);
nor U11555 (N_11555,N_11241,N_11384);
nand U11556 (N_11556,N_11279,N_11317);
or U11557 (N_11557,N_11134,N_11054);
nor U11558 (N_11558,N_11163,N_11341);
nand U11559 (N_11559,N_11426,N_11356);
nor U11560 (N_11560,N_11280,N_11350);
or U11561 (N_11561,N_11285,N_11133);
nor U11562 (N_11562,N_11301,N_11036);
or U11563 (N_11563,N_11099,N_11281);
or U11564 (N_11564,N_11303,N_11015);
nor U11565 (N_11565,N_11209,N_11154);
nor U11566 (N_11566,N_11025,N_11143);
xnor U11567 (N_11567,N_11344,N_11455);
nor U11568 (N_11568,N_11342,N_11169);
or U11569 (N_11569,N_11385,N_11082);
and U11570 (N_11570,N_11107,N_11355);
or U11571 (N_11571,N_11418,N_11245);
or U11572 (N_11572,N_11044,N_11077);
or U11573 (N_11573,N_11256,N_11436);
xor U11574 (N_11574,N_11010,N_11427);
xnor U11575 (N_11575,N_11171,N_11439);
or U11576 (N_11576,N_11190,N_11258);
or U11577 (N_11577,N_11367,N_11191);
and U11578 (N_11578,N_11037,N_11174);
and U11579 (N_11579,N_11240,N_11146);
xor U11580 (N_11580,N_11022,N_11088);
or U11581 (N_11581,N_11420,N_11075);
or U11582 (N_11582,N_11108,N_11276);
and U11583 (N_11583,N_11071,N_11354);
and U11584 (N_11584,N_11483,N_11486);
nand U11585 (N_11585,N_11305,N_11020);
nor U11586 (N_11586,N_11244,N_11274);
nand U11587 (N_11587,N_11459,N_11306);
nor U11588 (N_11588,N_11028,N_11212);
nand U11589 (N_11589,N_11389,N_11186);
nor U11590 (N_11590,N_11422,N_11474);
nor U11591 (N_11591,N_11377,N_11290);
or U11592 (N_11592,N_11009,N_11387);
nand U11593 (N_11593,N_11282,N_11184);
nor U11594 (N_11594,N_11289,N_11417);
nand U11595 (N_11595,N_11323,N_11340);
and U11596 (N_11596,N_11268,N_11390);
or U11597 (N_11597,N_11315,N_11326);
nor U11598 (N_11598,N_11277,N_11248);
and U11599 (N_11599,N_11484,N_11399);
nor U11600 (N_11600,N_11468,N_11181);
and U11601 (N_11601,N_11318,N_11214);
or U11602 (N_11602,N_11408,N_11402);
xor U11603 (N_11603,N_11330,N_11380);
nor U11604 (N_11604,N_11220,N_11187);
nand U11605 (N_11605,N_11193,N_11461);
xor U11606 (N_11606,N_11442,N_11229);
or U11607 (N_11607,N_11287,N_11343);
nand U11608 (N_11608,N_11065,N_11405);
nand U11609 (N_11609,N_11109,N_11066);
nand U11610 (N_11610,N_11084,N_11062);
nand U11611 (N_11611,N_11498,N_11152);
nor U11612 (N_11612,N_11359,N_11199);
and U11613 (N_11613,N_11237,N_11069);
or U11614 (N_11614,N_11403,N_11410);
or U11615 (N_11615,N_11255,N_11223);
nand U11616 (N_11616,N_11397,N_11424);
and U11617 (N_11617,N_11238,N_11308);
and U11618 (N_11618,N_11364,N_11148);
or U11619 (N_11619,N_11464,N_11052);
nand U11620 (N_11620,N_11047,N_11222);
and U11621 (N_11621,N_11487,N_11078);
nand U11622 (N_11622,N_11072,N_11260);
nor U11623 (N_11623,N_11242,N_11300);
nand U11624 (N_11624,N_11196,N_11081);
nor U11625 (N_11625,N_11001,N_11247);
nor U11626 (N_11626,N_11352,N_11150);
nor U11627 (N_11627,N_11331,N_11140);
nand U11628 (N_11628,N_11313,N_11430);
nand U11629 (N_11629,N_11239,N_11295);
xnor U11630 (N_11630,N_11018,N_11372);
nand U11631 (N_11631,N_11087,N_11173);
nor U11632 (N_11632,N_11470,N_11139);
nand U11633 (N_11633,N_11033,N_11057);
nor U11634 (N_11634,N_11125,N_11131);
nand U11635 (N_11635,N_11213,N_11160);
nand U11636 (N_11636,N_11118,N_11312);
nor U11637 (N_11637,N_11266,N_11040);
nor U11638 (N_11638,N_11302,N_11030);
or U11639 (N_11639,N_11406,N_11243);
nor U11640 (N_11640,N_11262,N_11117);
nand U11641 (N_11641,N_11053,N_11102);
nand U11642 (N_11642,N_11032,N_11297);
or U11643 (N_11643,N_11115,N_11156);
nand U11644 (N_11644,N_11135,N_11205);
and U11645 (N_11645,N_11159,N_11415);
nor U11646 (N_11646,N_11055,N_11369);
xnor U11647 (N_11647,N_11392,N_11371);
xor U11648 (N_11648,N_11450,N_11059);
xnor U11649 (N_11649,N_11166,N_11491);
nand U11650 (N_11650,N_11316,N_11404);
and U11651 (N_11651,N_11207,N_11153);
or U11652 (N_11652,N_11273,N_11334);
or U11653 (N_11653,N_11019,N_11395);
nand U11654 (N_11654,N_11127,N_11061);
and U11655 (N_11655,N_11070,N_11309);
nor U11656 (N_11656,N_11145,N_11363);
nor U11657 (N_11657,N_11124,N_11038);
nand U11658 (N_11658,N_11259,N_11466);
or U11659 (N_11659,N_11413,N_11444);
and U11660 (N_11660,N_11157,N_11296);
nor U11661 (N_11661,N_11122,N_11368);
xnor U11662 (N_11662,N_11014,N_11233);
or U11663 (N_11663,N_11170,N_11469);
and U11664 (N_11664,N_11458,N_11228);
nor U11665 (N_11665,N_11050,N_11224);
or U11666 (N_11666,N_11265,N_11391);
or U11667 (N_11667,N_11079,N_11130);
and U11668 (N_11668,N_11314,N_11005);
or U11669 (N_11669,N_11197,N_11149);
nand U11670 (N_11670,N_11056,N_11043);
and U11671 (N_11671,N_11128,N_11017);
and U11672 (N_11672,N_11269,N_11457);
or U11673 (N_11673,N_11000,N_11219);
or U11674 (N_11674,N_11489,N_11253);
or U11675 (N_11675,N_11105,N_11294);
nor U11676 (N_11676,N_11164,N_11175);
and U11677 (N_11677,N_11482,N_11217);
nor U11678 (N_11678,N_11479,N_11185);
or U11679 (N_11679,N_11257,N_11162);
and U11680 (N_11680,N_11210,N_11348);
and U11681 (N_11681,N_11362,N_11080);
nand U11682 (N_11682,N_11051,N_11421);
or U11683 (N_11683,N_11126,N_11068);
nand U11684 (N_11684,N_11339,N_11029);
and U11685 (N_11685,N_11155,N_11182);
or U11686 (N_11686,N_11045,N_11147);
and U11687 (N_11687,N_11488,N_11012);
or U11688 (N_11688,N_11388,N_11490);
nand U11689 (N_11689,N_11180,N_11286);
and U11690 (N_11690,N_11493,N_11183);
or U11691 (N_11691,N_11379,N_11365);
and U11692 (N_11692,N_11454,N_11106);
nor U11693 (N_11693,N_11304,N_11411);
nor U11694 (N_11694,N_11357,N_11412);
nand U11695 (N_11695,N_11382,N_11007);
or U11696 (N_11696,N_11101,N_11096);
and U11697 (N_11697,N_11480,N_11345);
or U11698 (N_11698,N_11008,N_11360);
nand U11699 (N_11699,N_11386,N_11261);
or U11700 (N_11700,N_11307,N_11234);
nand U11701 (N_11701,N_11188,N_11119);
and U11702 (N_11702,N_11324,N_11311);
and U11703 (N_11703,N_11144,N_11366);
or U11704 (N_11704,N_11215,N_11497);
xnor U11705 (N_11705,N_11383,N_11023);
xor U11706 (N_11706,N_11467,N_11451);
and U11707 (N_11707,N_11319,N_11063);
and U11708 (N_11708,N_11425,N_11035);
or U11709 (N_11709,N_11039,N_11230);
or U11710 (N_11710,N_11283,N_11299);
and U11711 (N_11711,N_11098,N_11227);
and U11712 (N_11712,N_11447,N_11208);
and U11713 (N_11713,N_11167,N_11414);
and U11714 (N_11714,N_11485,N_11027);
and U11715 (N_11715,N_11400,N_11236);
nor U11716 (N_11716,N_11095,N_11235);
and U11717 (N_11717,N_11024,N_11263);
or U11718 (N_11718,N_11225,N_11473);
and U11719 (N_11719,N_11346,N_11494);
or U11720 (N_11720,N_11465,N_11141);
or U11721 (N_11721,N_11333,N_11452);
nand U11722 (N_11722,N_11216,N_11003);
and U11723 (N_11723,N_11177,N_11423);
xnor U11724 (N_11724,N_11158,N_11499);
and U11725 (N_11725,N_11478,N_11165);
and U11726 (N_11726,N_11111,N_11374);
or U11727 (N_11727,N_11113,N_11138);
xor U11728 (N_11728,N_11325,N_11076);
or U11729 (N_11729,N_11204,N_11328);
nor U11730 (N_11730,N_11433,N_11370);
nor U11731 (N_11731,N_11132,N_11453);
nor U11732 (N_11732,N_11201,N_11151);
or U11733 (N_11733,N_11085,N_11049);
nand U11734 (N_11734,N_11178,N_11046);
and U11735 (N_11735,N_11327,N_11393);
and U11736 (N_11736,N_11251,N_11463);
or U11737 (N_11737,N_11083,N_11074);
nand U11738 (N_11738,N_11429,N_11100);
nand U11739 (N_11739,N_11206,N_11272);
nand U11740 (N_11740,N_11221,N_11168);
nor U11741 (N_11741,N_11093,N_11092);
nor U11742 (N_11742,N_11202,N_11495);
nor U11743 (N_11743,N_11004,N_11292);
nor U11744 (N_11744,N_11041,N_11310);
nor U11745 (N_11745,N_11351,N_11203);
and U11746 (N_11746,N_11250,N_11067);
or U11747 (N_11747,N_11349,N_11016);
or U11748 (N_11748,N_11086,N_11116);
or U11749 (N_11749,N_11358,N_11398);
or U11750 (N_11750,N_11444,N_11063);
or U11751 (N_11751,N_11101,N_11269);
nand U11752 (N_11752,N_11299,N_11332);
and U11753 (N_11753,N_11037,N_11395);
nand U11754 (N_11754,N_11477,N_11133);
and U11755 (N_11755,N_11412,N_11191);
and U11756 (N_11756,N_11311,N_11444);
nor U11757 (N_11757,N_11203,N_11388);
and U11758 (N_11758,N_11348,N_11207);
and U11759 (N_11759,N_11050,N_11156);
and U11760 (N_11760,N_11284,N_11498);
nor U11761 (N_11761,N_11110,N_11121);
and U11762 (N_11762,N_11161,N_11067);
and U11763 (N_11763,N_11134,N_11411);
or U11764 (N_11764,N_11067,N_11194);
and U11765 (N_11765,N_11042,N_11197);
and U11766 (N_11766,N_11043,N_11471);
or U11767 (N_11767,N_11369,N_11119);
nor U11768 (N_11768,N_11046,N_11232);
xnor U11769 (N_11769,N_11266,N_11482);
and U11770 (N_11770,N_11280,N_11268);
and U11771 (N_11771,N_11151,N_11313);
nor U11772 (N_11772,N_11326,N_11053);
nor U11773 (N_11773,N_11375,N_11433);
and U11774 (N_11774,N_11414,N_11110);
or U11775 (N_11775,N_11438,N_11394);
or U11776 (N_11776,N_11239,N_11416);
nand U11777 (N_11777,N_11376,N_11373);
nor U11778 (N_11778,N_11316,N_11164);
or U11779 (N_11779,N_11057,N_11351);
or U11780 (N_11780,N_11360,N_11159);
and U11781 (N_11781,N_11238,N_11471);
nor U11782 (N_11782,N_11188,N_11087);
nand U11783 (N_11783,N_11289,N_11278);
or U11784 (N_11784,N_11178,N_11401);
xnor U11785 (N_11785,N_11137,N_11179);
and U11786 (N_11786,N_11099,N_11432);
nor U11787 (N_11787,N_11324,N_11382);
and U11788 (N_11788,N_11229,N_11221);
or U11789 (N_11789,N_11265,N_11091);
and U11790 (N_11790,N_11461,N_11166);
nor U11791 (N_11791,N_11198,N_11401);
or U11792 (N_11792,N_11159,N_11152);
or U11793 (N_11793,N_11278,N_11195);
nand U11794 (N_11794,N_11125,N_11402);
and U11795 (N_11795,N_11203,N_11056);
nor U11796 (N_11796,N_11361,N_11166);
or U11797 (N_11797,N_11426,N_11149);
nand U11798 (N_11798,N_11028,N_11471);
or U11799 (N_11799,N_11484,N_11325);
or U11800 (N_11800,N_11084,N_11493);
nand U11801 (N_11801,N_11374,N_11290);
nand U11802 (N_11802,N_11125,N_11475);
nor U11803 (N_11803,N_11054,N_11434);
and U11804 (N_11804,N_11034,N_11342);
xor U11805 (N_11805,N_11293,N_11091);
xor U11806 (N_11806,N_11333,N_11041);
nand U11807 (N_11807,N_11344,N_11262);
xor U11808 (N_11808,N_11358,N_11184);
and U11809 (N_11809,N_11412,N_11317);
and U11810 (N_11810,N_11334,N_11009);
nor U11811 (N_11811,N_11138,N_11238);
or U11812 (N_11812,N_11037,N_11453);
nand U11813 (N_11813,N_11314,N_11375);
or U11814 (N_11814,N_11421,N_11163);
and U11815 (N_11815,N_11257,N_11489);
nor U11816 (N_11816,N_11347,N_11241);
or U11817 (N_11817,N_11124,N_11293);
or U11818 (N_11818,N_11484,N_11058);
and U11819 (N_11819,N_11108,N_11163);
and U11820 (N_11820,N_11260,N_11156);
and U11821 (N_11821,N_11374,N_11124);
and U11822 (N_11822,N_11349,N_11199);
or U11823 (N_11823,N_11288,N_11395);
nand U11824 (N_11824,N_11076,N_11104);
or U11825 (N_11825,N_11161,N_11391);
nor U11826 (N_11826,N_11147,N_11498);
nand U11827 (N_11827,N_11026,N_11021);
nor U11828 (N_11828,N_11195,N_11075);
xor U11829 (N_11829,N_11163,N_11451);
nor U11830 (N_11830,N_11113,N_11026);
nor U11831 (N_11831,N_11221,N_11355);
and U11832 (N_11832,N_11154,N_11083);
nor U11833 (N_11833,N_11453,N_11257);
nand U11834 (N_11834,N_11275,N_11023);
nor U11835 (N_11835,N_11266,N_11284);
and U11836 (N_11836,N_11273,N_11421);
nand U11837 (N_11837,N_11164,N_11002);
nor U11838 (N_11838,N_11424,N_11401);
nand U11839 (N_11839,N_11050,N_11305);
or U11840 (N_11840,N_11339,N_11366);
or U11841 (N_11841,N_11287,N_11405);
or U11842 (N_11842,N_11458,N_11053);
nand U11843 (N_11843,N_11482,N_11246);
and U11844 (N_11844,N_11204,N_11127);
and U11845 (N_11845,N_11390,N_11404);
xor U11846 (N_11846,N_11051,N_11066);
or U11847 (N_11847,N_11440,N_11034);
and U11848 (N_11848,N_11176,N_11300);
or U11849 (N_11849,N_11461,N_11063);
and U11850 (N_11850,N_11183,N_11380);
nand U11851 (N_11851,N_11135,N_11347);
nor U11852 (N_11852,N_11445,N_11141);
xor U11853 (N_11853,N_11478,N_11430);
nand U11854 (N_11854,N_11294,N_11356);
and U11855 (N_11855,N_11283,N_11005);
nor U11856 (N_11856,N_11180,N_11280);
or U11857 (N_11857,N_11167,N_11261);
nand U11858 (N_11858,N_11323,N_11147);
or U11859 (N_11859,N_11120,N_11483);
and U11860 (N_11860,N_11278,N_11099);
nor U11861 (N_11861,N_11186,N_11023);
nand U11862 (N_11862,N_11015,N_11085);
xor U11863 (N_11863,N_11343,N_11359);
or U11864 (N_11864,N_11061,N_11020);
or U11865 (N_11865,N_11357,N_11350);
nor U11866 (N_11866,N_11064,N_11047);
and U11867 (N_11867,N_11183,N_11213);
nor U11868 (N_11868,N_11077,N_11001);
or U11869 (N_11869,N_11281,N_11201);
and U11870 (N_11870,N_11049,N_11202);
nor U11871 (N_11871,N_11204,N_11383);
nand U11872 (N_11872,N_11019,N_11100);
and U11873 (N_11873,N_11392,N_11080);
nand U11874 (N_11874,N_11488,N_11306);
and U11875 (N_11875,N_11486,N_11461);
and U11876 (N_11876,N_11006,N_11064);
nand U11877 (N_11877,N_11351,N_11273);
nand U11878 (N_11878,N_11217,N_11282);
or U11879 (N_11879,N_11368,N_11121);
nand U11880 (N_11880,N_11412,N_11458);
nor U11881 (N_11881,N_11459,N_11433);
nand U11882 (N_11882,N_11433,N_11319);
and U11883 (N_11883,N_11413,N_11079);
and U11884 (N_11884,N_11050,N_11106);
nand U11885 (N_11885,N_11007,N_11016);
and U11886 (N_11886,N_11332,N_11310);
nand U11887 (N_11887,N_11444,N_11492);
and U11888 (N_11888,N_11340,N_11284);
nand U11889 (N_11889,N_11479,N_11220);
xor U11890 (N_11890,N_11290,N_11013);
and U11891 (N_11891,N_11188,N_11461);
xor U11892 (N_11892,N_11113,N_11249);
nand U11893 (N_11893,N_11471,N_11368);
or U11894 (N_11894,N_11409,N_11296);
and U11895 (N_11895,N_11117,N_11151);
and U11896 (N_11896,N_11154,N_11159);
or U11897 (N_11897,N_11026,N_11379);
and U11898 (N_11898,N_11073,N_11496);
nand U11899 (N_11899,N_11295,N_11376);
and U11900 (N_11900,N_11190,N_11067);
nand U11901 (N_11901,N_11135,N_11174);
or U11902 (N_11902,N_11051,N_11049);
xor U11903 (N_11903,N_11359,N_11219);
nor U11904 (N_11904,N_11202,N_11451);
or U11905 (N_11905,N_11238,N_11352);
nand U11906 (N_11906,N_11375,N_11379);
nand U11907 (N_11907,N_11155,N_11150);
or U11908 (N_11908,N_11199,N_11164);
xnor U11909 (N_11909,N_11062,N_11012);
nand U11910 (N_11910,N_11403,N_11444);
nor U11911 (N_11911,N_11361,N_11160);
nand U11912 (N_11912,N_11200,N_11360);
xor U11913 (N_11913,N_11343,N_11355);
or U11914 (N_11914,N_11317,N_11488);
xnor U11915 (N_11915,N_11297,N_11461);
or U11916 (N_11916,N_11269,N_11366);
or U11917 (N_11917,N_11267,N_11441);
and U11918 (N_11918,N_11220,N_11107);
nand U11919 (N_11919,N_11424,N_11171);
or U11920 (N_11920,N_11029,N_11036);
and U11921 (N_11921,N_11270,N_11080);
or U11922 (N_11922,N_11497,N_11096);
nand U11923 (N_11923,N_11456,N_11293);
or U11924 (N_11924,N_11093,N_11448);
or U11925 (N_11925,N_11412,N_11384);
nand U11926 (N_11926,N_11419,N_11013);
and U11927 (N_11927,N_11078,N_11313);
and U11928 (N_11928,N_11106,N_11395);
xnor U11929 (N_11929,N_11364,N_11231);
or U11930 (N_11930,N_11101,N_11344);
nand U11931 (N_11931,N_11265,N_11107);
or U11932 (N_11932,N_11242,N_11379);
nor U11933 (N_11933,N_11264,N_11447);
nand U11934 (N_11934,N_11386,N_11052);
or U11935 (N_11935,N_11048,N_11336);
nand U11936 (N_11936,N_11062,N_11060);
and U11937 (N_11937,N_11336,N_11041);
nor U11938 (N_11938,N_11006,N_11316);
or U11939 (N_11939,N_11286,N_11453);
or U11940 (N_11940,N_11475,N_11259);
or U11941 (N_11941,N_11376,N_11282);
nor U11942 (N_11942,N_11415,N_11480);
and U11943 (N_11943,N_11342,N_11048);
nand U11944 (N_11944,N_11095,N_11072);
or U11945 (N_11945,N_11463,N_11347);
or U11946 (N_11946,N_11326,N_11185);
xor U11947 (N_11947,N_11164,N_11273);
nor U11948 (N_11948,N_11236,N_11247);
nor U11949 (N_11949,N_11159,N_11401);
or U11950 (N_11950,N_11200,N_11265);
nor U11951 (N_11951,N_11130,N_11346);
or U11952 (N_11952,N_11040,N_11196);
nand U11953 (N_11953,N_11225,N_11411);
nand U11954 (N_11954,N_11236,N_11214);
or U11955 (N_11955,N_11052,N_11134);
nor U11956 (N_11956,N_11318,N_11489);
or U11957 (N_11957,N_11467,N_11443);
and U11958 (N_11958,N_11391,N_11424);
and U11959 (N_11959,N_11156,N_11151);
or U11960 (N_11960,N_11416,N_11040);
nor U11961 (N_11961,N_11475,N_11215);
and U11962 (N_11962,N_11377,N_11218);
nor U11963 (N_11963,N_11473,N_11002);
and U11964 (N_11964,N_11260,N_11440);
or U11965 (N_11965,N_11005,N_11093);
xnor U11966 (N_11966,N_11371,N_11106);
nand U11967 (N_11967,N_11178,N_11175);
and U11968 (N_11968,N_11056,N_11227);
nand U11969 (N_11969,N_11299,N_11171);
nor U11970 (N_11970,N_11099,N_11312);
or U11971 (N_11971,N_11490,N_11257);
nand U11972 (N_11972,N_11105,N_11222);
and U11973 (N_11973,N_11205,N_11095);
and U11974 (N_11974,N_11459,N_11007);
nand U11975 (N_11975,N_11040,N_11314);
nand U11976 (N_11976,N_11048,N_11486);
nand U11977 (N_11977,N_11185,N_11325);
nand U11978 (N_11978,N_11378,N_11222);
nor U11979 (N_11979,N_11108,N_11380);
and U11980 (N_11980,N_11344,N_11166);
nand U11981 (N_11981,N_11151,N_11363);
and U11982 (N_11982,N_11419,N_11187);
nor U11983 (N_11983,N_11144,N_11075);
and U11984 (N_11984,N_11446,N_11313);
nand U11985 (N_11985,N_11137,N_11206);
or U11986 (N_11986,N_11284,N_11080);
or U11987 (N_11987,N_11394,N_11061);
and U11988 (N_11988,N_11116,N_11220);
or U11989 (N_11989,N_11100,N_11352);
and U11990 (N_11990,N_11171,N_11090);
or U11991 (N_11991,N_11009,N_11014);
or U11992 (N_11992,N_11384,N_11445);
or U11993 (N_11993,N_11125,N_11061);
or U11994 (N_11994,N_11260,N_11413);
and U11995 (N_11995,N_11106,N_11154);
and U11996 (N_11996,N_11356,N_11047);
nor U11997 (N_11997,N_11225,N_11109);
nand U11998 (N_11998,N_11268,N_11440);
or U11999 (N_11999,N_11208,N_11454);
nor U12000 (N_12000,N_11922,N_11986);
and U12001 (N_12001,N_11983,N_11745);
and U12002 (N_12002,N_11776,N_11638);
xnor U12003 (N_12003,N_11542,N_11836);
and U12004 (N_12004,N_11779,N_11686);
or U12005 (N_12005,N_11561,N_11803);
or U12006 (N_12006,N_11809,N_11866);
nand U12007 (N_12007,N_11702,N_11659);
nand U12008 (N_12008,N_11762,N_11564);
xnor U12009 (N_12009,N_11790,N_11903);
and U12010 (N_12010,N_11658,N_11877);
nor U12011 (N_12011,N_11885,N_11793);
or U12012 (N_12012,N_11910,N_11683);
xor U12013 (N_12013,N_11525,N_11596);
nor U12014 (N_12014,N_11926,N_11870);
or U12015 (N_12015,N_11919,N_11934);
nand U12016 (N_12016,N_11778,N_11573);
and U12017 (N_12017,N_11795,N_11710);
nor U12018 (N_12018,N_11559,N_11959);
or U12019 (N_12019,N_11879,N_11666);
and U12020 (N_12020,N_11580,N_11524);
or U12021 (N_12021,N_11878,N_11938);
nor U12022 (N_12022,N_11780,N_11689);
or U12023 (N_12023,N_11547,N_11656);
and U12024 (N_12024,N_11607,N_11916);
and U12025 (N_12025,N_11872,N_11904);
and U12026 (N_12026,N_11807,N_11582);
or U12027 (N_12027,N_11618,N_11847);
or U12028 (N_12028,N_11717,N_11967);
nor U12029 (N_12029,N_11798,N_11581);
or U12030 (N_12030,N_11929,N_11920);
nand U12031 (N_12031,N_11889,N_11634);
nor U12032 (N_12032,N_11534,N_11509);
nor U12033 (N_12033,N_11942,N_11535);
and U12034 (N_12034,N_11853,N_11936);
nor U12035 (N_12035,N_11801,N_11899);
and U12036 (N_12036,N_11900,N_11818);
nand U12037 (N_12037,N_11988,N_11529);
or U12038 (N_12038,N_11943,N_11980);
nor U12039 (N_12039,N_11727,N_11939);
nor U12040 (N_12040,N_11628,N_11894);
and U12041 (N_12041,N_11861,N_11987);
nor U12042 (N_12042,N_11556,N_11725);
xor U12043 (N_12043,N_11823,N_11568);
nor U12044 (N_12044,N_11517,N_11688);
nand U12045 (N_12045,N_11816,N_11852);
nor U12046 (N_12046,N_11597,N_11881);
nand U12047 (N_12047,N_11550,N_11583);
nand U12048 (N_12048,N_11921,N_11706);
or U12049 (N_12049,N_11569,N_11784);
xor U12050 (N_12050,N_11907,N_11911);
or U12051 (N_12051,N_11824,N_11845);
nand U12052 (N_12052,N_11901,N_11519);
nand U12053 (N_12053,N_11544,N_11738);
or U12054 (N_12054,N_11562,N_11546);
and U12055 (N_12055,N_11789,N_11577);
and U12056 (N_12056,N_11733,N_11575);
nand U12057 (N_12057,N_11844,N_11507);
xor U12058 (N_12058,N_11891,N_11643);
nor U12059 (N_12059,N_11591,N_11908);
nand U12060 (N_12060,N_11846,N_11874);
nand U12061 (N_12061,N_11694,N_11950);
and U12062 (N_12062,N_11704,N_11703);
and U12063 (N_12063,N_11932,N_11747);
or U12064 (N_12064,N_11746,N_11984);
nor U12065 (N_12065,N_11858,N_11671);
and U12066 (N_12066,N_11906,N_11956);
nand U12067 (N_12067,N_11636,N_11567);
nand U12068 (N_12068,N_11744,N_11917);
or U12069 (N_12069,N_11768,N_11912);
or U12070 (N_12070,N_11578,N_11810);
and U12071 (N_12071,N_11635,N_11948);
and U12072 (N_12072,N_11563,N_11715);
and U12073 (N_12073,N_11627,N_11961);
or U12074 (N_12074,N_11953,N_11979);
nand U12075 (N_12075,N_11617,N_11985);
or U12076 (N_12076,N_11679,N_11620);
nand U12077 (N_12077,N_11619,N_11832);
nor U12078 (N_12078,N_11586,N_11805);
nor U12079 (N_12079,N_11876,N_11646);
and U12080 (N_12080,N_11505,N_11705);
or U12081 (N_12081,N_11897,N_11642);
nor U12082 (N_12082,N_11735,N_11838);
xnor U12083 (N_12083,N_11608,N_11649);
nor U12084 (N_12084,N_11859,N_11696);
nor U12085 (N_12085,N_11652,N_11843);
and U12086 (N_12086,N_11662,N_11757);
nor U12087 (N_12087,N_11771,N_11572);
xor U12088 (N_12088,N_11681,N_11992);
nor U12089 (N_12089,N_11855,N_11557);
nor U12090 (N_12090,N_11684,N_11794);
or U12091 (N_12091,N_11660,N_11531);
nand U12092 (N_12092,N_11945,N_11835);
nor U12093 (N_12093,N_11740,N_11718);
nand U12094 (N_12094,N_11918,N_11522);
nor U12095 (N_12095,N_11698,N_11518);
or U12096 (N_12096,N_11962,N_11940);
xor U12097 (N_12097,N_11765,N_11654);
nand U12098 (N_12098,N_11584,N_11707);
or U12099 (N_12099,N_11975,N_11644);
and U12100 (N_12100,N_11722,N_11968);
or U12101 (N_12101,N_11763,N_11670);
xor U12102 (N_12102,N_11714,N_11630);
nor U12103 (N_12103,N_11516,N_11734);
and U12104 (N_12104,N_11501,N_11839);
nand U12105 (N_12105,N_11946,N_11842);
and U12106 (N_12106,N_11663,N_11592);
or U12107 (N_12107,N_11593,N_11817);
nand U12108 (N_12108,N_11513,N_11883);
nand U12109 (N_12109,N_11749,N_11549);
nand U12110 (N_12110,N_11570,N_11555);
or U12111 (N_12111,N_11895,N_11892);
or U12112 (N_12112,N_11554,N_11786);
and U12113 (N_12113,N_11752,N_11781);
and U12114 (N_12114,N_11840,N_11677);
and U12115 (N_12115,N_11648,N_11713);
or U12116 (N_12116,N_11792,N_11682);
and U12117 (N_12117,N_11651,N_11993);
nor U12118 (N_12118,N_11695,N_11965);
or U12119 (N_12119,N_11812,N_11724);
nand U12120 (N_12120,N_11813,N_11791);
and U12121 (N_12121,N_11873,N_11742);
and U12122 (N_12122,N_11611,N_11680);
nor U12123 (N_12123,N_11989,N_11804);
or U12124 (N_12124,N_11890,N_11761);
and U12125 (N_12125,N_11857,N_11560);
and U12126 (N_12126,N_11884,N_11782);
nand U12127 (N_12127,N_11621,N_11657);
and U12128 (N_12128,N_11665,N_11815);
and U12129 (N_12129,N_11831,N_11834);
or U12130 (N_12130,N_11772,N_11867);
nand U12131 (N_12131,N_11615,N_11783);
nand U12132 (N_12132,N_11587,N_11974);
nor U12133 (N_12133,N_11723,N_11991);
nand U12134 (N_12134,N_11741,N_11530);
xnor U12135 (N_12135,N_11588,N_11502);
nor U12136 (N_12136,N_11915,N_11520);
nor U12137 (N_12137,N_11958,N_11769);
nand U12138 (N_12138,N_11814,N_11709);
or U12139 (N_12139,N_11622,N_11601);
and U12140 (N_12140,N_11887,N_11821);
nor U12141 (N_12141,N_11811,N_11673);
nand U12142 (N_12142,N_11978,N_11537);
and U12143 (N_12143,N_11796,N_11775);
xor U12144 (N_12144,N_11650,N_11552);
nor U12145 (N_12145,N_11726,N_11655);
nand U12146 (N_12146,N_11672,N_11841);
nor U12147 (N_12147,N_11854,N_11830);
or U12148 (N_12148,N_11754,N_11758);
nor U12149 (N_12149,N_11609,N_11737);
or U12150 (N_12150,N_11914,N_11826);
or U12151 (N_12151,N_11731,N_11668);
nand U12152 (N_12152,N_11748,N_11716);
nand U12153 (N_12153,N_11849,N_11819);
or U12154 (N_12154,N_11576,N_11605);
and U12155 (N_12155,N_11977,N_11960);
nor U12156 (N_12156,N_11888,N_11641);
nor U12157 (N_12157,N_11909,N_11527);
xor U12158 (N_12158,N_11700,N_11925);
or U12159 (N_12159,N_11639,N_11699);
or U12160 (N_12160,N_11923,N_11970);
nor U12161 (N_12161,N_11541,N_11687);
xnor U12162 (N_12162,N_11598,N_11799);
nand U12163 (N_12163,N_11736,N_11949);
or U12164 (N_12164,N_11924,N_11558);
and U12165 (N_12165,N_11837,N_11603);
or U12166 (N_12166,N_11606,N_11963);
nor U12167 (N_12167,N_11508,N_11767);
nand U12168 (N_12168,N_11797,N_11701);
nand U12169 (N_12169,N_11905,N_11625);
nor U12170 (N_12170,N_11806,N_11770);
nand U12171 (N_12171,N_11711,N_11667);
nor U12172 (N_12172,N_11692,N_11935);
xnor U12173 (N_12173,N_11613,N_11594);
and U12174 (N_12174,N_11972,N_11629);
xnor U12175 (N_12175,N_11730,N_11869);
and U12176 (N_12176,N_11759,N_11633);
nand U12177 (N_12177,N_11600,N_11785);
nand U12178 (N_12178,N_11623,N_11712);
nand U12179 (N_12179,N_11676,N_11640);
xnor U12180 (N_12180,N_11982,N_11760);
or U12181 (N_12181,N_11571,N_11964);
and U12182 (N_12182,N_11875,N_11645);
and U12183 (N_12183,N_11739,N_11612);
and U12184 (N_12184,N_11957,N_11951);
nand U12185 (N_12185,N_11614,N_11595);
nand U12186 (N_12186,N_11822,N_11565);
or U12187 (N_12187,N_11825,N_11708);
and U12188 (N_12188,N_11589,N_11788);
nor U12189 (N_12189,N_11871,N_11808);
nor U12190 (N_12190,N_11976,N_11545);
xor U12191 (N_12191,N_11802,N_11928);
xor U12192 (N_12192,N_11787,N_11664);
nand U12193 (N_12193,N_11536,N_11604);
nand U12194 (N_12194,N_11902,N_11553);
nand U12195 (N_12195,N_11511,N_11675);
or U12196 (N_12196,N_11981,N_11751);
nand U12197 (N_12197,N_11721,N_11538);
or U12198 (N_12198,N_11882,N_11510);
xor U12199 (N_12199,N_11969,N_11990);
nand U12200 (N_12200,N_11863,N_11514);
nand U12201 (N_12201,N_11998,N_11856);
or U12202 (N_12202,N_11756,N_11632);
or U12203 (N_12203,N_11533,N_11674);
nand U12204 (N_12204,N_11548,N_11528);
and U12205 (N_12205,N_11868,N_11540);
or U12206 (N_12206,N_11994,N_11971);
nor U12207 (N_12207,N_11610,N_11693);
and U12208 (N_12208,N_11933,N_11820);
and U12209 (N_12209,N_11504,N_11997);
nand U12210 (N_12210,N_11503,N_11777);
or U12211 (N_12211,N_11774,N_11952);
or U12212 (N_12212,N_11637,N_11506);
nand U12213 (N_12213,N_11532,N_11973);
nor U12214 (N_12214,N_11848,N_11931);
and U12215 (N_12215,N_11690,N_11743);
nor U12216 (N_12216,N_11941,N_11697);
nor U12217 (N_12217,N_11661,N_11624);
and U12218 (N_12218,N_11893,N_11616);
and U12219 (N_12219,N_11999,N_11512);
nor U12220 (N_12220,N_11626,N_11865);
and U12221 (N_12221,N_11955,N_11574);
and U12222 (N_12222,N_11599,N_11526);
and U12223 (N_12223,N_11896,N_11579);
nor U12224 (N_12224,N_11551,N_11653);
and U12225 (N_12225,N_11764,N_11966);
nand U12226 (N_12226,N_11719,N_11631);
and U12227 (N_12227,N_11539,N_11996);
nor U12228 (N_12228,N_11543,N_11728);
nor U12229 (N_12229,N_11590,N_11829);
and U12230 (N_12230,N_11930,N_11850);
xor U12231 (N_12231,N_11937,N_11828);
nand U12232 (N_12232,N_11927,N_11750);
nor U12233 (N_12233,N_11602,N_11947);
and U12234 (N_12234,N_11864,N_11732);
nor U12235 (N_12235,N_11500,N_11566);
nand U12236 (N_12236,N_11898,N_11944);
xnor U12237 (N_12237,N_11833,N_11880);
or U12238 (N_12238,N_11585,N_11862);
or U12239 (N_12239,N_11755,N_11995);
or U12240 (N_12240,N_11860,N_11766);
nor U12241 (N_12241,N_11691,N_11800);
nand U12242 (N_12242,N_11523,N_11827);
nor U12243 (N_12243,N_11913,N_11720);
nor U12244 (N_12244,N_11647,N_11685);
nand U12245 (N_12245,N_11773,N_11851);
and U12246 (N_12246,N_11886,N_11753);
or U12247 (N_12247,N_11669,N_11729);
nor U12248 (N_12248,N_11515,N_11521);
or U12249 (N_12249,N_11954,N_11678);
and U12250 (N_12250,N_11535,N_11785);
nand U12251 (N_12251,N_11927,N_11531);
nand U12252 (N_12252,N_11740,N_11938);
or U12253 (N_12253,N_11990,N_11813);
and U12254 (N_12254,N_11664,N_11546);
nor U12255 (N_12255,N_11920,N_11734);
and U12256 (N_12256,N_11792,N_11697);
or U12257 (N_12257,N_11671,N_11795);
nand U12258 (N_12258,N_11828,N_11597);
nor U12259 (N_12259,N_11989,N_11536);
nor U12260 (N_12260,N_11811,N_11682);
and U12261 (N_12261,N_11695,N_11707);
nand U12262 (N_12262,N_11591,N_11509);
nand U12263 (N_12263,N_11961,N_11520);
nand U12264 (N_12264,N_11668,N_11727);
and U12265 (N_12265,N_11600,N_11821);
nand U12266 (N_12266,N_11572,N_11703);
nor U12267 (N_12267,N_11501,N_11888);
nor U12268 (N_12268,N_11656,N_11688);
nand U12269 (N_12269,N_11758,N_11625);
nand U12270 (N_12270,N_11993,N_11750);
nor U12271 (N_12271,N_11768,N_11897);
or U12272 (N_12272,N_11523,N_11858);
or U12273 (N_12273,N_11847,N_11791);
or U12274 (N_12274,N_11570,N_11714);
or U12275 (N_12275,N_11986,N_11533);
or U12276 (N_12276,N_11924,N_11703);
and U12277 (N_12277,N_11534,N_11833);
or U12278 (N_12278,N_11894,N_11933);
nor U12279 (N_12279,N_11631,N_11949);
and U12280 (N_12280,N_11659,N_11539);
xnor U12281 (N_12281,N_11926,N_11578);
or U12282 (N_12282,N_11771,N_11766);
and U12283 (N_12283,N_11816,N_11690);
nand U12284 (N_12284,N_11621,N_11655);
xnor U12285 (N_12285,N_11659,N_11934);
nand U12286 (N_12286,N_11569,N_11521);
and U12287 (N_12287,N_11962,N_11894);
nand U12288 (N_12288,N_11927,N_11729);
and U12289 (N_12289,N_11618,N_11588);
and U12290 (N_12290,N_11754,N_11997);
or U12291 (N_12291,N_11708,N_11515);
nand U12292 (N_12292,N_11788,N_11552);
or U12293 (N_12293,N_11739,N_11946);
and U12294 (N_12294,N_11887,N_11680);
and U12295 (N_12295,N_11784,N_11903);
or U12296 (N_12296,N_11543,N_11945);
and U12297 (N_12297,N_11925,N_11860);
or U12298 (N_12298,N_11519,N_11825);
or U12299 (N_12299,N_11808,N_11741);
nor U12300 (N_12300,N_11647,N_11610);
nand U12301 (N_12301,N_11993,N_11845);
or U12302 (N_12302,N_11926,N_11819);
nand U12303 (N_12303,N_11924,N_11779);
or U12304 (N_12304,N_11625,N_11673);
and U12305 (N_12305,N_11563,N_11639);
and U12306 (N_12306,N_11974,N_11698);
nor U12307 (N_12307,N_11619,N_11669);
nand U12308 (N_12308,N_11649,N_11791);
or U12309 (N_12309,N_11643,N_11555);
nand U12310 (N_12310,N_11603,N_11523);
nand U12311 (N_12311,N_11756,N_11589);
xor U12312 (N_12312,N_11923,N_11632);
and U12313 (N_12313,N_11541,N_11744);
xnor U12314 (N_12314,N_11534,N_11869);
and U12315 (N_12315,N_11526,N_11737);
xnor U12316 (N_12316,N_11589,N_11839);
or U12317 (N_12317,N_11904,N_11604);
or U12318 (N_12318,N_11807,N_11959);
or U12319 (N_12319,N_11844,N_11643);
or U12320 (N_12320,N_11778,N_11801);
and U12321 (N_12321,N_11935,N_11540);
or U12322 (N_12322,N_11946,N_11710);
and U12323 (N_12323,N_11680,N_11774);
and U12324 (N_12324,N_11881,N_11550);
and U12325 (N_12325,N_11886,N_11979);
nand U12326 (N_12326,N_11513,N_11570);
or U12327 (N_12327,N_11660,N_11655);
xor U12328 (N_12328,N_11747,N_11641);
nand U12329 (N_12329,N_11872,N_11826);
and U12330 (N_12330,N_11548,N_11644);
nand U12331 (N_12331,N_11519,N_11733);
and U12332 (N_12332,N_11549,N_11856);
nor U12333 (N_12333,N_11826,N_11792);
nor U12334 (N_12334,N_11797,N_11986);
or U12335 (N_12335,N_11549,N_11948);
or U12336 (N_12336,N_11877,N_11582);
nand U12337 (N_12337,N_11678,N_11965);
nand U12338 (N_12338,N_11935,N_11526);
and U12339 (N_12339,N_11692,N_11693);
and U12340 (N_12340,N_11641,N_11861);
or U12341 (N_12341,N_11823,N_11846);
nand U12342 (N_12342,N_11829,N_11995);
and U12343 (N_12343,N_11806,N_11961);
or U12344 (N_12344,N_11816,N_11836);
nor U12345 (N_12345,N_11686,N_11964);
or U12346 (N_12346,N_11759,N_11649);
and U12347 (N_12347,N_11982,N_11635);
nand U12348 (N_12348,N_11983,N_11780);
and U12349 (N_12349,N_11565,N_11926);
and U12350 (N_12350,N_11717,N_11753);
nor U12351 (N_12351,N_11783,N_11818);
and U12352 (N_12352,N_11925,N_11713);
nor U12353 (N_12353,N_11879,N_11968);
nand U12354 (N_12354,N_11846,N_11890);
and U12355 (N_12355,N_11847,N_11627);
and U12356 (N_12356,N_11737,N_11916);
nor U12357 (N_12357,N_11739,N_11971);
nor U12358 (N_12358,N_11731,N_11612);
nor U12359 (N_12359,N_11863,N_11780);
nand U12360 (N_12360,N_11578,N_11568);
and U12361 (N_12361,N_11998,N_11972);
xor U12362 (N_12362,N_11501,N_11510);
and U12363 (N_12363,N_11942,N_11792);
and U12364 (N_12364,N_11994,N_11678);
and U12365 (N_12365,N_11980,N_11532);
xor U12366 (N_12366,N_11662,N_11678);
nand U12367 (N_12367,N_11971,N_11734);
or U12368 (N_12368,N_11854,N_11590);
nor U12369 (N_12369,N_11970,N_11506);
or U12370 (N_12370,N_11597,N_11860);
nand U12371 (N_12371,N_11713,N_11879);
and U12372 (N_12372,N_11835,N_11693);
and U12373 (N_12373,N_11733,N_11722);
nand U12374 (N_12374,N_11937,N_11907);
or U12375 (N_12375,N_11562,N_11528);
xnor U12376 (N_12376,N_11983,N_11737);
and U12377 (N_12377,N_11912,N_11761);
nand U12378 (N_12378,N_11738,N_11888);
nand U12379 (N_12379,N_11681,N_11553);
or U12380 (N_12380,N_11542,N_11970);
and U12381 (N_12381,N_11618,N_11799);
and U12382 (N_12382,N_11626,N_11568);
and U12383 (N_12383,N_11560,N_11575);
nand U12384 (N_12384,N_11679,N_11933);
nand U12385 (N_12385,N_11766,N_11840);
and U12386 (N_12386,N_11634,N_11825);
nor U12387 (N_12387,N_11753,N_11721);
nor U12388 (N_12388,N_11748,N_11644);
or U12389 (N_12389,N_11924,N_11719);
xnor U12390 (N_12390,N_11821,N_11900);
nand U12391 (N_12391,N_11940,N_11578);
or U12392 (N_12392,N_11945,N_11676);
or U12393 (N_12393,N_11867,N_11756);
nand U12394 (N_12394,N_11742,N_11893);
xnor U12395 (N_12395,N_11854,N_11976);
nor U12396 (N_12396,N_11778,N_11855);
nand U12397 (N_12397,N_11999,N_11699);
or U12398 (N_12398,N_11546,N_11552);
or U12399 (N_12399,N_11876,N_11536);
nand U12400 (N_12400,N_11722,N_11748);
or U12401 (N_12401,N_11605,N_11858);
nand U12402 (N_12402,N_11721,N_11587);
or U12403 (N_12403,N_11623,N_11749);
or U12404 (N_12404,N_11649,N_11643);
xor U12405 (N_12405,N_11841,N_11888);
and U12406 (N_12406,N_11706,N_11733);
nor U12407 (N_12407,N_11723,N_11733);
nand U12408 (N_12408,N_11658,N_11798);
xor U12409 (N_12409,N_11771,N_11822);
and U12410 (N_12410,N_11501,N_11900);
and U12411 (N_12411,N_11624,N_11988);
xnor U12412 (N_12412,N_11895,N_11920);
xnor U12413 (N_12413,N_11545,N_11827);
xor U12414 (N_12414,N_11613,N_11714);
nand U12415 (N_12415,N_11935,N_11831);
or U12416 (N_12416,N_11655,N_11797);
or U12417 (N_12417,N_11595,N_11919);
nand U12418 (N_12418,N_11971,N_11833);
and U12419 (N_12419,N_11830,N_11784);
nor U12420 (N_12420,N_11564,N_11717);
nor U12421 (N_12421,N_11775,N_11783);
nand U12422 (N_12422,N_11771,N_11574);
and U12423 (N_12423,N_11647,N_11975);
or U12424 (N_12424,N_11558,N_11847);
xnor U12425 (N_12425,N_11959,N_11758);
xnor U12426 (N_12426,N_11623,N_11524);
nor U12427 (N_12427,N_11788,N_11763);
nor U12428 (N_12428,N_11637,N_11995);
or U12429 (N_12429,N_11759,N_11806);
nor U12430 (N_12430,N_11863,N_11727);
or U12431 (N_12431,N_11909,N_11633);
and U12432 (N_12432,N_11555,N_11852);
nand U12433 (N_12433,N_11896,N_11900);
or U12434 (N_12434,N_11609,N_11560);
nand U12435 (N_12435,N_11527,N_11580);
or U12436 (N_12436,N_11594,N_11551);
xnor U12437 (N_12437,N_11666,N_11543);
nor U12438 (N_12438,N_11878,N_11652);
nor U12439 (N_12439,N_11919,N_11913);
nor U12440 (N_12440,N_11825,N_11913);
and U12441 (N_12441,N_11984,N_11665);
nor U12442 (N_12442,N_11656,N_11621);
nand U12443 (N_12443,N_11612,N_11943);
or U12444 (N_12444,N_11949,N_11670);
nor U12445 (N_12445,N_11641,N_11635);
and U12446 (N_12446,N_11758,N_11917);
and U12447 (N_12447,N_11641,N_11930);
nor U12448 (N_12448,N_11695,N_11884);
and U12449 (N_12449,N_11597,N_11704);
and U12450 (N_12450,N_11740,N_11783);
nand U12451 (N_12451,N_11534,N_11628);
xor U12452 (N_12452,N_11669,N_11792);
xor U12453 (N_12453,N_11658,N_11782);
and U12454 (N_12454,N_11555,N_11687);
or U12455 (N_12455,N_11884,N_11743);
nand U12456 (N_12456,N_11836,N_11607);
or U12457 (N_12457,N_11727,N_11821);
nor U12458 (N_12458,N_11584,N_11752);
and U12459 (N_12459,N_11770,N_11643);
or U12460 (N_12460,N_11910,N_11927);
or U12461 (N_12461,N_11716,N_11622);
and U12462 (N_12462,N_11663,N_11774);
or U12463 (N_12463,N_11746,N_11797);
or U12464 (N_12464,N_11811,N_11998);
or U12465 (N_12465,N_11734,N_11687);
nand U12466 (N_12466,N_11827,N_11540);
or U12467 (N_12467,N_11936,N_11646);
or U12468 (N_12468,N_11531,N_11946);
nand U12469 (N_12469,N_11885,N_11755);
nor U12470 (N_12470,N_11779,N_11764);
xnor U12471 (N_12471,N_11919,N_11622);
or U12472 (N_12472,N_11509,N_11770);
and U12473 (N_12473,N_11524,N_11933);
or U12474 (N_12474,N_11846,N_11533);
and U12475 (N_12475,N_11960,N_11649);
nor U12476 (N_12476,N_11547,N_11990);
and U12477 (N_12477,N_11812,N_11988);
nand U12478 (N_12478,N_11817,N_11569);
xor U12479 (N_12479,N_11562,N_11652);
nand U12480 (N_12480,N_11582,N_11921);
or U12481 (N_12481,N_11539,N_11872);
and U12482 (N_12482,N_11841,N_11652);
nand U12483 (N_12483,N_11886,N_11917);
xor U12484 (N_12484,N_11905,N_11709);
nand U12485 (N_12485,N_11928,N_11810);
nor U12486 (N_12486,N_11982,N_11726);
nand U12487 (N_12487,N_11799,N_11791);
xnor U12488 (N_12488,N_11747,N_11734);
or U12489 (N_12489,N_11778,N_11746);
or U12490 (N_12490,N_11983,N_11543);
nor U12491 (N_12491,N_11990,N_11704);
nor U12492 (N_12492,N_11683,N_11609);
and U12493 (N_12493,N_11607,N_11730);
and U12494 (N_12494,N_11880,N_11594);
or U12495 (N_12495,N_11955,N_11946);
nand U12496 (N_12496,N_11504,N_11918);
xnor U12497 (N_12497,N_11809,N_11665);
or U12498 (N_12498,N_11556,N_11755);
and U12499 (N_12499,N_11696,N_11867);
or U12500 (N_12500,N_12012,N_12214);
nand U12501 (N_12501,N_12147,N_12454);
xor U12502 (N_12502,N_12165,N_12235);
or U12503 (N_12503,N_12104,N_12186);
and U12504 (N_12504,N_12305,N_12318);
and U12505 (N_12505,N_12390,N_12316);
or U12506 (N_12506,N_12334,N_12443);
nor U12507 (N_12507,N_12362,N_12450);
or U12508 (N_12508,N_12154,N_12244);
and U12509 (N_12509,N_12282,N_12021);
nand U12510 (N_12510,N_12019,N_12156);
xor U12511 (N_12511,N_12082,N_12369);
nor U12512 (N_12512,N_12432,N_12204);
or U12513 (N_12513,N_12057,N_12052);
or U12514 (N_12514,N_12304,N_12293);
or U12515 (N_12515,N_12242,N_12364);
and U12516 (N_12516,N_12459,N_12308);
and U12517 (N_12517,N_12475,N_12243);
nor U12518 (N_12518,N_12209,N_12492);
nor U12519 (N_12519,N_12105,N_12341);
or U12520 (N_12520,N_12030,N_12327);
nand U12521 (N_12521,N_12134,N_12275);
nand U12522 (N_12522,N_12382,N_12264);
nor U12523 (N_12523,N_12345,N_12295);
xor U12524 (N_12524,N_12170,N_12313);
or U12525 (N_12525,N_12425,N_12494);
nor U12526 (N_12526,N_12368,N_12284);
or U12527 (N_12527,N_12339,N_12177);
and U12528 (N_12528,N_12054,N_12053);
and U12529 (N_12529,N_12497,N_12399);
or U12530 (N_12530,N_12207,N_12413);
and U12531 (N_12531,N_12033,N_12353);
nand U12532 (N_12532,N_12039,N_12051);
nor U12533 (N_12533,N_12191,N_12452);
and U12534 (N_12534,N_12300,N_12229);
and U12535 (N_12535,N_12085,N_12438);
xnor U12536 (N_12536,N_12110,N_12137);
or U12537 (N_12537,N_12061,N_12409);
and U12538 (N_12538,N_12066,N_12289);
nor U12539 (N_12539,N_12312,N_12268);
or U12540 (N_12540,N_12167,N_12143);
nor U12541 (N_12541,N_12499,N_12011);
and U12542 (N_12542,N_12172,N_12359);
nor U12543 (N_12543,N_12258,N_12132);
or U12544 (N_12544,N_12067,N_12222);
nor U12545 (N_12545,N_12106,N_12123);
nor U12546 (N_12546,N_12480,N_12476);
nand U12547 (N_12547,N_12255,N_12153);
or U12548 (N_12548,N_12270,N_12278);
nand U12549 (N_12549,N_12280,N_12026);
nand U12550 (N_12550,N_12469,N_12001);
nand U12551 (N_12551,N_12403,N_12108);
and U12552 (N_12552,N_12371,N_12237);
or U12553 (N_12553,N_12276,N_12215);
nor U12554 (N_12554,N_12471,N_12175);
nor U12555 (N_12555,N_12113,N_12198);
nand U12556 (N_12556,N_12451,N_12197);
and U12557 (N_12557,N_12095,N_12265);
nand U12558 (N_12558,N_12365,N_12436);
and U12559 (N_12559,N_12329,N_12223);
or U12560 (N_12560,N_12093,N_12481);
or U12561 (N_12561,N_12400,N_12107);
or U12562 (N_12562,N_12047,N_12396);
and U12563 (N_12563,N_12094,N_12145);
xor U12564 (N_12564,N_12048,N_12421);
xor U12565 (N_12565,N_12079,N_12389);
nor U12566 (N_12566,N_12126,N_12383);
nor U12567 (N_12567,N_12122,N_12391);
nand U12568 (N_12568,N_12395,N_12491);
nor U12569 (N_12569,N_12091,N_12234);
nor U12570 (N_12570,N_12392,N_12354);
nor U12571 (N_12571,N_12272,N_12103);
nor U12572 (N_12572,N_12135,N_12006);
nand U12573 (N_12573,N_12424,N_12417);
or U12574 (N_12574,N_12393,N_12381);
and U12575 (N_12575,N_12457,N_12285);
nand U12576 (N_12576,N_12299,N_12325);
xnor U12577 (N_12577,N_12431,N_12183);
nor U12578 (N_12578,N_12224,N_12455);
and U12579 (N_12579,N_12343,N_12406);
nand U12580 (N_12580,N_12131,N_12462);
and U12581 (N_12581,N_12081,N_12130);
and U12582 (N_12582,N_12309,N_12068);
nor U12583 (N_12583,N_12227,N_12496);
nand U12584 (N_12584,N_12384,N_12340);
or U12585 (N_12585,N_12332,N_12031);
and U12586 (N_12586,N_12041,N_12298);
and U12587 (N_12587,N_12319,N_12337);
nand U12588 (N_12588,N_12205,N_12212);
nand U12589 (N_12589,N_12064,N_12428);
or U12590 (N_12590,N_12010,N_12490);
nand U12591 (N_12591,N_12314,N_12461);
or U12592 (N_12592,N_12083,N_12065);
nand U12593 (N_12593,N_12374,N_12114);
nor U12594 (N_12594,N_12072,N_12380);
xnor U12595 (N_12595,N_12288,N_12330);
and U12596 (N_12596,N_12144,N_12181);
xnor U12597 (N_12597,N_12296,N_12444);
or U12598 (N_12598,N_12248,N_12286);
nor U12599 (N_12599,N_12251,N_12037);
nand U12600 (N_12600,N_12097,N_12274);
nor U12601 (N_12601,N_12301,N_12283);
xnor U12602 (N_12602,N_12018,N_12044);
nand U12603 (N_12603,N_12092,N_12446);
or U12604 (N_12604,N_12166,N_12350);
xor U12605 (N_12605,N_12401,N_12324);
or U12606 (N_12606,N_12073,N_12155);
or U12607 (N_12607,N_12349,N_12281);
nor U12608 (N_12608,N_12426,N_12253);
nand U12609 (N_12609,N_12089,N_12419);
xor U12610 (N_12610,N_12291,N_12463);
xor U12611 (N_12611,N_12164,N_12404);
and U12612 (N_12612,N_12157,N_12259);
xor U12613 (N_12613,N_12146,N_12375);
nand U12614 (N_12614,N_12029,N_12009);
nor U12615 (N_12615,N_12348,N_12479);
nand U12616 (N_12616,N_12378,N_12005);
or U12617 (N_12617,N_12000,N_12239);
nor U12618 (N_12618,N_12078,N_12034);
nor U12619 (N_12619,N_12387,N_12453);
nand U12620 (N_12620,N_12199,N_12058);
xor U12621 (N_12621,N_12422,N_12493);
nor U12622 (N_12622,N_12460,N_12306);
or U12623 (N_12623,N_12184,N_12036);
nand U12624 (N_12624,N_12358,N_12331);
or U12625 (N_12625,N_12077,N_12075);
xor U12626 (N_12626,N_12323,N_12456);
nand U12627 (N_12627,N_12192,N_12003);
or U12628 (N_12628,N_12238,N_12180);
or U12629 (N_12629,N_12120,N_12260);
or U12630 (N_12630,N_12182,N_12117);
and U12631 (N_12631,N_12178,N_12467);
nand U12632 (N_12632,N_12441,N_12101);
or U12633 (N_12633,N_12379,N_12252);
nor U12634 (N_12634,N_12124,N_12007);
or U12635 (N_12635,N_12023,N_12254);
and U12636 (N_12636,N_12257,N_12179);
and U12637 (N_12637,N_12290,N_12152);
or U12638 (N_12638,N_12464,N_12326);
nor U12639 (N_12639,N_12218,N_12230);
or U12640 (N_12640,N_12335,N_12430);
and U12641 (N_12641,N_12249,N_12488);
nand U12642 (N_12642,N_12429,N_12347);
and U12643 (N_12643,N_12294,N_12038);
or U12644 (N_12644,N_12133,N_12211);
nor U12645 (N_12645,N_12096,N_12407);
and U12646 (N_12646,N_12195,N_12333);
nor U12647 (N_12647,N_12376,N_12484);
or U12648 (N_12648,N_12398,N_12473);
nand U12649 (N_12649,N_12213,N_12076);
or U12650 (N_12650,N_12161,N_12206);
nand U12651 (N_12651,N_12099,N_12344);
nor U12652 (N_12652,N_12189,N_12040);
nand U12653 (N_12653,N_12024,N_12263);
nand U12654 (N_12654,N_12112,N_12303);
nor U12655 (N_12655,N_12042,N_12159);
and U12656 (N_12656,N_12055,N_12355);
nor U12657 (N_12657,N_12250,N_12202);
nor U12658 (N_12658,N_12321,N_12489);
nor U12659 (N_12659,N_12433,N_12231);
and U12660 (N_12660,N_12140,N_12188);
nor U12661 (N_12661,N_12017,N_12025);
and U12662 (N_12662,N_12056,N_12427);
nand U12663 (N_12663,N_12098,N_12266);
nand U12664 (N_12664,N_12468,N_12013);
or U12665 (N_12665,N_12466,N_12414);
nor U12666 (N_12666,N_12228,N_12062);
nand U12667 (N_12667,N_12423,N_12472);
and U12668 (N_12668,N_12129,N_12069);
nor U12669 (N_12669,N_12201,N_12084);
nand U12670 (N_12670,N_12190,N_12267);
or U12671 (N_12671,N_12498,N_12035);
nor U12672 (N_12672,N_12437,N_12176);
xnor U12673 (N_12673,N_12236,N_12169);
or U12674 (N_12674,N_12185,N_12086);
nand U12675 (N_12675,N_12418,N_12050);
nor U12676 (N_12676,N_12118,N_12402);
nor U12677 (N_12677,N_12168,N_12063);
and U12678 (N_12678,N_12128,N_12412);
nor U12679 (N_12679,N_12351,N_12328);
or U12680 (N_12680,N_12315,N_12022);
or U12681 (N_12681,N_12148,N_12158);
nand U12682 (N_12682,N_12478,N_12317);
and U12683 (N_12683,N_12221,N_12232);
nand U12684 (N_12684,N_12142,N_12372);
nand U12685 (N_12685,N_12322,N_12482);
nand U12686 (N_12686,N_12439,N_12311);
and U12687 (N_12687,N_12015,N_12287);
or U12688 (N_12688,N_12447,N_12277);
and U12689 (N_12689,N_12032,N_12139);
nor U12690 (N_12690,N_12448,N_12151);
nor U12691 (N_12691,N_12043,N_12420);
or U12692 (N_12692,N_12302,N_12416);
nor U12693 (N_12693,N_12342,N_12028);
nor U12694 (N_12694,N_12338,N_12487);
and U12695 (N_12695,N_12100,N_12486);
nand U12696 (N_12696,N_12203,N_12495);
and U12697 (N_12697,N_12116,N_12090);
xnor U12698 (N_12698,N_12004,N_12356);
and U12699 (N_12699,N_12088,N_12174);
or U12700 (N_12700,N_12320,N_12370);
nor U12701 (N_12701,N_12138,N_12386);
or U12702 (N_12702,N_12219,N_12070);
nor U12703 (N_12703,N_12458,N_12102);
or U12704 (N_12704,N_12415,N_12173);
nor U12705 (N_12705,N_12397,N_12474);
or U12706 (N_12706,N_12435,N_12160);
xnor U12707 (N_12707,N_12136,N_12269);
nor U12708 (N_12708,N_12014,N_12240);
nor U12709 (N_12709,N_12208,N_12210);
or U12710 (N_12710,N_12119,N_12465);
and U12711 (N_12711,N_12121,N_12247);
or U12712 (N_12712,N_12162,N_12071);
and U12713 (N_12713,N_12226,N_12049);
and U12714 (N_12714,N_12225,N_12233);
nand U12715 (N_12715,N_12171,N_12394);
or U12716 (N_12716,N_12352,N_12008);
nand U12717 (N_12717,N_12477,N_12405);
and U12718 (N_12718,N_12216,N_12193);
and U12719 (N_12719,N_12262,N_12150);
nand U12720 (N_12720,N_12373,N_12279);
nand U12721 (N_12721,N_12271,N_12363);
nor U12722 (N_12722,N_12080,N_12385);
nor U12723 (N_12723,N_12109,N_12046);
nand U12724 (N_12724,N_12307,N_12346);
or U12725 (N_12725,N_12408,N_12045);
nand U12726 (N_12726,N_12360,N_12273);
nand U12727 (N_12727,N_12336,N_12256);
and U12728 (N_12728,N_12087,N_12246);
nor U12729 (N_12729,N_12297,N_12361);
or U12730 (N_12730,N_12411,N_12020);
nor U12731 (N_12731,N_12194,N_12127);
xnor U12732 (N_12732,N_12434,N_12196);
or U12733 (N_12733,N_12485,N_12187);
nand U12734 (N_12734,N_12449,N_12366);
or U12735 (N_12735,N_12483,N_12217);
nor U12736 (N_12736,N_12241,N_12445);
or U12737 (N_12737,N_12141,N_12310);
or U12738 (N_12738,N_12442,N_12367);
nor U12739 (N_12739,N_12111,N_12245);
nor U12740 (N_12740,N_12470,N_12059);
xnor U12741 (N_12741,N_12125,N_12220);
or U12742 (N_12742,N_12163,N_12440);
xnor U12743 (N_12743,N_12074,N_12149);
or U12744 (N_12744,N_12016,N_12027);
and U12745 (N_12745,N_12292,N_12410);
and U12746 (N_12746,N_12002,N_12357);
nor U12747 (N_12747,N_12115,N_12261);
and U12748 (N_12748,N_12060,N_12377);
and U12749 (N_12749,N_12388,N_12200);
xor U12750 (N_12750,N_12467,N_12317);
or U12751 (N_12751,N_12257,N_12226);
or U12752 (N_12752,N_12334,N_12157);
nor U12753 (N_12753,N_12290,N_12049);
nor U12754 (N_12754,N_12413,N_12451);
nor U12755 (N_12755,N_12108,N_12240);
nor U12756 (N_12756,N_12090,N_12140);
nor U12757 (N_12757,N_12223,N_12313);
or U12758 (N_12758,N_12416,N_12214);
or U12759 (N_12759,N_12456,N_12321);
nor U12760 (N_12760,N_12040,N_12034);
or U12761 (N_12761,N_12275,N_12357);
and U12762 (N_12762,N_12143,N_12209);
nor U12763 (N_12763,N_12117,N_12055);
and U12764 (N_12764,N_12381,N_12447);
and U12765 (N_12765,N_12031,N_12285);
or U12766 (N_12766,N_12097,N_12012);
or U12767 (N_12767,N_12033,N_12336);
xor U12768 (N_12768,N_12052,N_12060);
nand U12769 (N_12769,N_12275,N_12329);
nand U12770 (N_12770,N_12251,N_12497);
nand U12771 (N_12771,N_12390,N_12339);
nor U12772 (N_12772,N_12320,N_12042);
and U12773 (N_12773,N_12407,N_12170);
nand U12774 (N_12774,N_12178,N_12021);
nand U12775 (N_12775,N_12451,N_12085);
nor U12776 (N_12776,N_12090,N_12046);
and U12777 (N_12777,N_12087,N_12434);
and U12778 (N_12778,N_12285,N_12088);
xor U12779 (N_12779,N_12422,N_12237);
or U12780 (N_12780,N_12248,N_12309);
xnor U12781 (N_12781,N_12260,N_12367);
nand U12782 (N_12782,N_12149,N_12418);
and U12783 (N_12783,N_12082,N_12243);
nand U12784 (N_12784,N_12270,N_12329);
and U12785 (N_12785,N_12366,N_12062);
or U12786 (N_12786,N_12390,N_12207);
xnor U12787 (N_12787,N_12381,N_12132);
or U12788 (N_12788,N_12177,N_12061);
nand U12789 (N_12789,N_12327,N_12494);
nor U12790 (N_12790,N_12482,N_12487);
nor U12791 (N_12791,N_12403,N_12360);
nand U12792 (N_12792,N_12257,N_12326);
xnor U12793 (N_12793,N_12275,N_12236);
and U12794 (N_12794,N_12458,N_12440);
or U12795 (N_12795,N_12022,N_12393);
xor U12796 (N_12796,N_12096,N_12457);
and U12797 (N_12797,N_12154,N_12272);
nor U12798 (N_12798,N_12271,N_12411);
and U12799 (N_12799,N_12364,N_12266);
or U12800 (N_12800,N_12433,N_12277);
nand U12801 (N_12801,N_12471,N_12033);
or U12802 (N_12802,N_12171,N_12253);
nor U12803 (N_12803,N_12330,N_12208);
nand U12804 (N_12804,N_12344,N_12130);
or U12805 (N_12805,N_12313,N_12427);
and U12806 (N_12806,N_12375,N_12467);
and U12807 (N_12807,N_12394,N_12366);
and U12808 (N_12808,N_12136,N_12106);
nand U12809 (N_12809,N_12062,N_12006);
or U12810 (N_12810,N_12379,N_12403);
xor U12811 (N_12811,N_12285,N_12333);
or U12812 (N_12812,N_12322,N_12303);
nor U12813 (N_12813,N_12373,N_12449);
or U12814 (N_12814,N_12433,N_12056);
xor U12815 (N_12815,N_12353,N_12125);
and U12816 (N_12816,N_12128,N_12052);
nor U12817 (N_12817,N_12210,N_12398);
and U12818 (N_12818,N_12398,N_12032);
nor U12819 (N_12819,N_12085,N_12206);
nor U12820 (N_12820,N_12351,N_12046);
nor U12821 (N_12821,N_12101,N_12182);
nand U12822 (N_12822,N_12196,N_12481);
or U12823 (N_12823,N_12204,N_12214);
nor U12824 (N_12824,N_12078,N_12045);
nor U12825 (N_12825,N_12164,N_12049);
nor U12826 (N_12826,N_12189,N_12232);
nor U12827 (N_12827,N_12338,N_12316);
and U12828 (N_12828,N_12492,N_12355);
or U12829 (N_12829,N_12164,N_12198);
nor U12830 (N_12830,N_12433,N_12018);
or U12831 (N_12831,N_12371,N_12219);
or U12832 (N_12832,N_12128,N_12132);
nand U12833 (N_12833,N_12275,N_12293);
nor U12834 (N_12834,N_12218,N_12009);
or U12835 (N_12835,N_12238,N_12027);
or U12836 (N_12836,N_12059,N_12119);
and U12837 (N_12837,N_12307,N_12062);
and U12838 (N_12838,N_12269,N_12283);
nand U12839 (N_12839,N_12351,N_12250);
nand U12840 (N_12840,N_12189,N_12298);
and U12841 (N_12841,N_12120,N_12080);
and U12842 (N_12842,N_12432,N_12229);
or U12843 (N_12843,N_12295,N_12494);
nand U12844 (N_12844,N_12139,N_12244);
nor U12845 (N_12845,N_12266,N_12103);
nor U12846 (N_12846,N_12181,N_12061);
and U12847 (N_12847,N_12209,N_12199);
nand U12848 (N_12848,N_12212,N_12358);
and U12849 (N_12849,N_12124,N_12263);
xnor U12850 (N_12850,N_12004,N_12254);
nor U12851 (N_12851,N_12039,N_12002);
nand U12852 (N_12852,N_12274,N_12141);
xnor U12853 (N_12853,N_12344,N_12428);
and U12854 (N_12854,N_12156,N_12445);
or U12855 (N_12855,N_12205,N_12421);
and U12856 (N_12856,N_12477,N_12304);
nor U12857 (N_12857,N_12278,N_12091);
and U12858 (N_12858,N_12099,N_12360);
nor U12859 (N_12859,N_12284,N_12358);
nor U12860 (N_12860,N_12469,N_12327);
nand U12861 (N_12861,N_12074,N_12147);
or U12862 (N_12862,N_12401,N_12119);
nor U12863 (N_12863,N_12089,N_12280);
nand U12864 (N_12864,N_12125,N_12127);
nand U12865 (N_12865,N_12053,N_12089);
and U12866 (N_12866,N_12392,N_12153);
and U12867 (N_12867,N_12438,N_12261);
nand U12868 (N_12868,N_12045,N_12221);
nand U12869 (N_12869,N_12289,N_12296);
nand U12870 (N_12870,N_12024,N_12178);
nor U12871 (N_12871,N_12326,N_12374);
xnor U12872 (N_12872,N_12171,N_12357);
or U12873 (N_12873,N_12081,N_12267);
or U12874 (N_12874,N_12380,N_12315);
and U12875 (N_12875,N_12140,N_12065);
nand U12876 (N_12876,N_12111,N_12472);
or U12877 (N_12877,N_12280,N_12022);
or U12878 (N_12878,N_12298,N_12477);
or U12879 (N_12879,N_12266,N_12379);
and U12880 (N_12880,N_12486,N_12219);
nor U12881 (N_12881,N_12165,N_12309);
and U12882 (N_12882,N_12240,N_12153);
or U12883 (N_12883,N_12121,N_12024);
or U12884 (N_12884,N_12041,N_12285);
or U12885 (N_12885,N_12324,N_12056);
nand U12886 (N_12886,N_12148,N_12021);
and U12887 (N_12887,N_12105,N_12371);
or U12888 (N_12888,N_12040,N_12219);
or U12889 (N_12889,N_12160,N_12428);
or U12890 (N_12890,N_12412,N_12068);
nor U12891 (N_12891,N_12418,N_12126);
nor U12892 (N_12892,N_12096,N_12209);
xnor U12893 (N_12893,N_12135,N_12173);
nor U12894 (N_12894,N_12218,N_12441);
or U12895 (N_12895,N_12452,N_12016);
and U12896 (N_12896,N_12098,N_12210);
nor U12897 (N_12897,N_12328,N_12476);
nor U12898 (N_12898,N_12381,N_12234);
nand U12899 (N_12899,N_12461,N_12378);
and U12900 (N_12900,N_12317,N_12334);
nand U12901 (N_12901,N_12372,N_12286);
or U12902 (N_12902,N_12107,N_12463);
nand U12903 (N_12903,N_12000,N_12240);
and U12904 (N_12904,N_12404,N_12470);
or U12905 (N_12905,N_12253,N_12397);
or U12906 (N_12906,N_12402,N_12104);
nand U12907 (N_12907,N_12001,N_12044);
or U12908 (N_12908,N_12321,N_12114);
xnor U12909 (N_12909,N_12005,N_12234);
or U12910 (N_12910,N_12483,N_12158);
and U12911 (N_12911,N_12484,N_12023);
nor U12912 (N_12912,N_12192,N_12293);
and U12913 (N_12913,N_12213,N_12015);
nor U12914 (N_12914,N_12430,N_12268);
or U12915 (N_12915,N_12202,N_12066);
nand U12916 (N_12916,N_12271,N_12393);
nand U12917 (N_12917,N_12119,N_12266);
nor U12918 (N_12918,N_12049,N_12112);
and U12919 (N_12919,N_12149,N_12480);
and U12920 (N_12920,N_12131,N_12390);
nand U12921 (N_12921,N_12417,N_12266);
nor U12922 (N_12922,N_12370,N_12054);
or U12923 (N_12923,N_12440,N_12341);
and U12924 (N_12924,N_12310,N_12405);
xnor U12925 (N_12925,N_12282,N_12012);
nor U12926 (N_12926,N_12386,N_12361);
and U12927 (N_12927,N_12190,N_12265);
or U12928 (N_12928,N_12096,N_12072);
nand U12929 (N_12929,N_12122,N_12142);
and U12930 (N_12930,N_12346,N_12019);
nor U12931 (N_12931,N_12238,N_12008);
nand U12932 (N_12932,N_12321,N_12285);
or U12933 (N_12933,N_12418,N_12188);
or U12934 (N_12934,N_12321,N_12230);
nand U12935 (N_12935,N_12393,N_12023);
nand U12936 (N_12936,N_12432,N_12196);
nor U12937 (N_12937,N_12152,N_12379);
and U12938 (N_12938,N_12188,N_12274);
nand U12939 (N_12939,N_12089,N_12450);
or U12940 (N_12940,N_12400,N_12088);
or U12941 (N_12941,N_12305,N_12339);
nand U12942 (N_12942,N_12418,N_12457);
nand U12943 (N_12943,N_12146,N_12051);
nand U12944 (N_12944,N_12234,N_12144);
nand U12945 (N_12945,N_12193,N_12274);
and U12946 (N_12946,N_12203,N_12293);
xnor U12947 (N_12947,N_12156,N_12161);
nand U12948 (N_12948,N_12111,N_12344);
nor U12949 (N_12949,N_12107,N_12381);
nand U12950 (N_12950,N_12213,N_12157);
nand U12951 (N_12951,N_12498,N_12229);
nor U12952 (N_12952,N_12321,N_12309);
or U12953 (N_12953,N_12383,N_12400);
xor U12954 (N_12954,N_12036,N_12074);
or U12955 (N_12955,N_12248,N_12147);
nand U12956 (N_12956,N_12424,N_12354);
nand U12957 (N_12957,N_12379,N_12340);
and U12958 (N_12958,N_12141,N_12124);
or U12959 (N_12959,N_12203,N_12391);
and U12960 (N_12960,N_12380,N_12111);
nor U12961 (N_12961,N_12282,N_12242);
nor U12962 (N_12962,N_12235,N_12209);
nand U12963 (N_12963,N_12484,N_12450);
xor U12964 (N_12964,N_12281,N_12016);
nor U12965 (N_12965,N_12447,N_12011);
or U12966 (N_12966,N_12018,N_12498);
nor U12967 (N_12967,N_12118,N_12042);
and U12968 (N_12968,N_12123,N_12314);
xor U12969 (N_12969,N_12374,N_12158);
nor U12970 (N_12970,N_12499,N_12376);
nor U12971 (N_12971,N_12036,N_12162);
nor U12972 (N_12972,N_12058,N_12051);
nor U12973 (N_12973,N_12164,N_12459);
nand U12974 (N_12974,N_12080,N_12464);
or U12975 (N_12975,N_12209,N_12100);
nand U12976 (N_12976,N_12309,N_12279);
nor U12977 (N_12977,N_12024,N_12189);
nand U12978 (N_12978,N_12122,N_12285);
and U12979 (N_12979,N_12058,N_12251);
xnor U12980 (N_12980,N_12405,N_12220);
or U12981 (N_12981,N_12399,N_12193);
and U12982 (N_12982,N_12157,N_12251);
nor U12983 (N_12983,N_12189,N_12484);
and U12984 (N_12984,N_12276,N_12327);
or U12985 (N_12985,N_12435,N_12253);
or U12986 (N_12986,N_12396,N_12008);
nor U12987 (N_12987,N_12461,N_12254);
or U12988 (N_12988,N_12037,N_12244);
or U12989 (N_12989,N_12287,N_12087);
nor U12990 (N_12990,N_12423,N_12288);
and U12991 (N_12991,N_12311,N_12483);
or U12992 (N_12992,N_12493,N_12406);
nor U12993 (N_12993,N_12364,N_12059);
or U12994 (N_12994,N_12111,N_12462);
and U12995 (N_12995,N_12363,N_12427);
xnor U12996 (N_12996,N_12034,N_12221);
nor U12997 (N_12997,N_12319,N_12459);
or U12998 (N_12998,N_12211,N_12298);
and U12999 (N_12999,N_12289,N_12446);
nand U13000 (N_13000,N_12914,N_12599);
nor U13001 (N_13001,N_12697,N_12594);
nand U13002 (N_13002,N_12731,N_12506);
xor U13003 (N_13003,N_12972,N_12867);
nor U13004 (N_13004,N_12513,N_12569);
nor U13005 (N_13005,N_12684,N_12981);
nand U13006 (N_13006,N_12600,N_12648);
or U13007 (N_13007,N_12714,N_12749);
nor U13008 (N_13008,N_12609,N_12712);
and U13009 (N_13009,N_12614,N_12514);
nor U13010 (N_13010,N_12892,N_12797);
or U13011 (N_13011,N_12547,N_12852);
nand U13012 (N_13012,N_12935,N_12702);
nor U13013 (N_13013,N_12806,N_12964);
xnor U13014 (N_13014,N_12561,N_12755);
nand U13015 (N_13015,N_12817,N_12791);
nand U13016 (N_13016,N_12926,N_12652);
or U13017 (N_13017,N_12616,N_12898);
nand U13018 (N_13018,N_12532,N_12665);
and U13019 (N_13019,N_12709,N_12963);
or U13020 (N_13020,N_12801,N_12588);
nor U13021 (N_13021,N_12857,N_12668);
or U13022 (N_13022,N_12869,N_12848);
nor U13023 (N_13023,N_12654,N_12580);
nor U13024 (N_13024,N_12968,N_12582);
nor U13025 (N_13025,N_12982,N_12876);
nor U13026 (N_13026,N_12534,N_12978);
nor U13027 (N_13027,N_12761,N_12556);
nor U13028 (N_13028,N_12713,N_12944);
or U13029 (N_13029,N_12945,N_12593);
and U13030 (N_13030,N_12507,N_12786);
nor U13031 (N_13031,N_12805,N_12525);
nor U13032 (N_13032,N_12781,N_12906);
nor U13033 (N_13033,N_12780,N_12732);
and U13034 (N_13034,N_12856,N_12723);
xnor U13035 (N_13035,N_12657,N_12634);
and U13036 (N_13036,N_12790,N_12638);
xnor U13037 (N_13037,N_12728,N_12853);
nor U13038 (N_13038,N_12900,N_12842);
or U13039 (N_13039,N_12785,N_12639);
nor U13040 (N_13040,N_12585,N_12858);
and U13041 (N_13041,N_12640,N_12573);
and U13042 (N_13042,N_12773,N_12823);
xnor U13043 (N_13043,N_12918,N_12825);
nor U13044 (N_13044,N_12672,N_12976);
and U13045 (N_13045,N_12757,N_12896);
nor U13046 (N_13046,N_12596,N_12597);
xnor U13047 (N_13047,N_12895,N_12592);
nor U13048 (N_13048,N_12824,N_12940);
and U13049 (N_13049,N_12522,N_12618);
nor U13050 (N_13050,N_12501,N_12811);
or U13051 (N_13051,N_12620,N_12567);
xnor U13052 (N_13052,N_12726,N_12658);
nand U13053 (N_13053,N_12962,N_12741);
nor U13054 (N_13054,N_12645,N_12529);
or U13055 (N_13055,N_12610,N_12524);
and U13056 (N_13056,N_12576,N_12637);
nor U13057 (N_13057,N_12512,N_12903);
or U13058 (N_13058,N_12719,N_12936);
nor U13059 (N_13059,N_12676,N_12661);
xnor U13060 (N_13060,N_12743,N_12720);
nor U13061 (N_13061,N_12942,N_12535);
nor U13062 (N_13062,N_12571,N_12696);
nand U13063 (N_13063,N_12641,N_12932);
xnor U13064 (N_13064,N_12861,N_12974);
and U13065 (N_13065,N_12798,N_12839);
nand U13066 (N_13066,N_12746,N_12559);
and U13067 (N_13067,N_12540,N_12958);
and U13068 (N_13068,N_12931,N_12626);
xnor U13069 (N_13069,N_12987,N_12562);
and U13070 (N_13070,N_12538,N_12969);
nor U13071 (N_13071,N_12531,N_12815);
nor U13072 (N_13072,N_12554,N_12663);
xor U13073 (N_13073,N_12586,N_12920);
or U13074 (N_13074,N_12560,N_12998);
or U13075 (N_13075,N_12991,N_12765);
nor U13076 (N_13076,N_12893,N_12838);
xnor U13077 (N_13077,N_12802,N_12566);
or U13078 (N_13078,N_12704,N_12961);
nor U13079 (N_13079,N_12681,N_12759);
and U13080 (N_13080,N_12565,N_12787);
nor U13081 (N_13081,N_12715,N_12555);
or U13082 (N_13082,N_12691,N_12778);
or U13083 (N_13083,N_12705,N_12794);
or U13084 (N_13084,N_12740,N_12557);
or U13085 (N_13085,N_12651,N_12727);
or U13086 (N_13086,N_12776,N_12544);
nor U13087 (N_13087,N_12568,N_12748);
nand U13088 (N_13088,N_12664,N_12635);
nor U13089 (N_13089,N_12859,N_12827);
nor U13090 (N_13090,N_12623,N_12849);
nand U13091 (N_13091,N_12753,N_12701);
and U13092 (N_13092,N_12996,N_12826);
and U13093 (N_13093,N_12971,N_12647);
nor U13094 (N_13094,N_12503,N_12779);
or U13095 (N_13095,N_12624,N_12843);
xnor U13096 (N_13096,N_12572,N_12995);
nor U13097 (N_13097,N_12885,N_12927);
nand U13098 (N_13098,N_12956,N_12718);
or U13099 (N_13099,N_12934,N_12888);
or U13100 (N_13100,N_12537,N_12551);
nand U13101 (N_13101,N_12734,N_12783);
nand U13102 (N_13102,N_12882,N_12500);
nor U13103 (N_13103,N_12533,N_12679);
and U13104 (N_13104,N_12502,N_12539);
or U13105 (N_13105,N_12908,N_12793);
or U13106 (N_13106,N_12649,N_12970);
or U13107 (N_13107,N_12870,N_12751);
xor U13108 (N_13108,N_12946,N_12643);
and U13109 (N_13109,N_12916,N_12921);
or U13110 (N_13110,N_12833,N_12733);
and U13111 (N_13111,N_12683,N_12789);
and U13112 (N_13112,N_12677,N_12771);
nand U13113 (N_13113,N_12807,N_12922);
nor U13114 (N_13114,N_12541,N_12632);
and U13115 (N_13115,N_12711,N_12659);
nand U13116 (N_13116,N_12850,N_12703);
or U13117 (N_13117,N_12602,N_12605);
and U13118 (N_13118,N_12504,N_12994);
nor U13119 (N_13119,N_12716,N_12722);
and U13120 (N_13120,N_12905,N_12990);
and U13121 (N_13121,N_12980,N_12619);
nor U13122 (N_13122,N_12830,N_12788);
nand U13123 (N_13123,N_12615,N_12989);
nor U13124 (N_13124,N_12855,N_12814);
xor U13125 (N_13125,N_12965,N_12767);
nand U13126 (N_13126,N_12782,N_12685);
and U13127 (N_13127,N_12880,N_12628);
nand U13128 (N_13128,N_12510,N_12766);
xnor U13129 (N_13129,N_12873,N_12508);
nand U13130 (N_13130,N_12915,N_12772);
nand U13131 (N_13131,N_12924,N_12866);
nand U13132 (N_13132,N_12803,N_12700);
nor U13133 (N_13133,N_12774,N_12578);
nor U13134 (N_13134,N_12611,N_12997);
xnor U13135 (N_13135,N_12622,N_12505);
or U13136 (N_13136,N_12546,N_12591);
xor U13137 (N_13137,N_12947,N_12983);
nor U13138 (N_13138,N_12881,N_12836);
nor U13139 (N_13139,N_12536,N_12819);
xor U13140 (N_13140,N_12517,N_12937);
nor U13141 (N_13141,N_12577,N_12975);
nand U13142 (N_13142,N_12952,N_12690);
and U13143 (N_13143,N_12831,N_12919);
xor U13144 (N_13144,N_12758,N_12897);
or U13145 (N_13145,N_12871,N_12549);
nand U13146 (N_13146,N_12985,N_12864);
nor U13147 (N_13147,N_12912,N_12840);
nor U13148 (N_13148,N_12841,N_12519);
or U13149 (N_13149,N_12608,N_12710);
nor U13150 (N_13150,N_12707,N_12689);
xnor U13151 (N_13151,N_12959,N_12894);
and U13152 (N_13152,N_12667,N_12809);
xor U13153 (N_13153,N_12558,N_12606);
and U13154 (N_13154,N_12631,N_12550);
nand U13155 (N_13155,N_12545,N_12682);
and U13156 (N_13156,N_12692,N_12526);
xor U13157 (N_13157,N_12613,N_12511);
nand U13158 (N_13158,N_12820,N_12953);
or U13159 (N_13159,N_12589,N_12553);
and U13160 (N_13160,N_12808,N_12627);
and U13161 (N_13161,N_12832,N_12769);
and U13162 (N_13162,N_12601,N_12950);
and U13163 (N_13163,N_12941,N_12845);
nand U13164 (N_13164,N_12584,N_12694);
or U13165 (N_13165,N_12570,N_12777);
nor U13166 (N_13166,N_12754,N_12943);
or U13167 (N_13167,N_12644,N_12509);
nand U13168 (N_13168,N_12875,N_12796);
nor U13169 (N_13169,N_12949,N_12607);
and U13170 (N_13170,N_12603,N_12518);
nor U13171 (N_13171,N_12579,N_12821);
nor U13172 (N_13172,N_12829,N_12973);
nand U13173 (N_13173,N_12574,N_12939);
and U13174 (N_13174,N_12736,N_12530);
xor U13175 (N_13175,N_12868,N_12521);
nand U13176 (N_13176,N_12879,N_12523);
or U13177 (N_13177,N_12828,N_12930);
and U13178 (N_13178,N_12902,N_12999);
nand U13179 (N_13179,N_12587,N_12834);
xnor U13180 (N_13180,N_12735,N_12564);
nand U13181 (N_13181,N_12886,N_12516);
nand U13182 (N_13182,N_12674,N_12737);
nor U13183 (N_13183,N_12854,N_12977);
and U13184 (N_13184,N_12948,N_12527);
and U13185 (N_13185,N_12889,N_12954);
and U13186 (N_13186,N_12739,N_12993);
xor U13187 (N_13187,N_12636,N_12646);
and U13188 (N_13188,N_12901,N_12951);
and U13189 (N_13189,N_12581,N_12884);
nand U13190 (N_13190,N_12775,N_12650);
and U13191 (N_13191,N_12515,N_12911);
xor U13192 (N_13192,N_12816,N_12686);
and U13193 (N_13193,N_12687,N_12678);
nor U13194 (N_13194,N_12653,N_12910);
nor U13195 (N_13195,N_12837,N_12890);
nor U13196 (N_13196,N_12520,N_12675);
and U13197 (N_13197,N_12917,N_12818);
or U13198 (N_13198,N_12604,N_12621);
nand U13199 (N_13199,N_12860,N_12729);
or U13200 (N_13200,N_12928,N_12706);
nor U13201 (N_13201,N_12770,N_12957);
xor U13202 (N_13202,N_12862,N_12795);
and U13203 (N_13203,N_12738,N_12810);
nor U13204 (N_13204,N_12548,N_12760);
nor U13205 (N_13205,N_12863,N_12925);
and U13206 (N_13206,N_12552,N_12625);
and U13207 (N_13207,N_12583,N_12986);
or U13208 (N_13208,N_12656,N_12979);
or U13209 (N_13209,N_12784,N_12680);
nor U13210 (N_13210,N_12800,N_12542);
nand U13211 (N_13211,N_12878,N_12891);
and U13212 (N_13212,N_12846,N_12938);
nor U13213 (N_13213,N_12708,N_12877);
and U13214 (N_13214,N_12865,N_12747);
or U13215 (N_13215,N_12813,N_12909);
or U13216 (N_13216,N_12655,N_12744);
nor U13217 (N_13217,N_12742,N_12633);
nand U13218 (N_13218,N_12904,N_12874);
or U13219 (N_13219,N_12792,N_12847);
nand U13220 (N_13220,N_12745,N_12752);
nand U13221 (N_13221,N_12669,N_12913);
and U13222 (N_13222,N_12992,N_12804);
and U13223 (N_13223,N_12764,N_12563);
xnor U13224 (N_13224,N_12717,N_12899);
or U13225 (N_13225,N_12629,N_12750);
or U13226 (N_13226,N_12612,N_12617);
nand U13227 (N_13227,N_12699,N_12756);
nor U13228 (N_13228,N_12851,N_12725);
and U13229 (N_13229,N_12660,N_12955);
nand U13230 (N_13230,N_12595,N_12543);
or U13231 (N_13231,N_12923,N_12844);
nand U13232 (N_13232,N_12812,N_12966);
or U13233 (N_13233,N_12929,N_12984);
nand U13234 (N_13234,N_12642,N_12960);
nor U13235 (N_13235,N_12666,N_12883);
or U13236 (N_13236,N_12698,N_12590);
xor U13237 (N_13237,N_12762,N_12724);
xor U13238 (N_13238,N_12763,N_12670);
or U13239 (N_13239,N_12695,N_12730);
or U13240 (N_13240,N_12528,N_12887);
nor U13241 (N_13241,N_12721,N_12598);
nor U13242 (N_13242,N_12673,N_12872);
nor U13243 (N_13243,N_12768,N_12988);
nor U13244 (N_13244,N_12933,N_12799);
nor U13245 (N_13245,N_12693,N_12822);
xnor U13246 (N_13246,N_12662,N_12967);
or U13247 (N_13247,N_12835,N_12688);
xor U13248 (N_13248,N_12575,N_12671);
nor U13249 (N_13249,N_12630,N_12907);
and U13250 (N_13250,N_12798,N_12705);
nor U13251 (N_13251,N_12931,N_12960);
nand U13252 (N_13252,N_12915,N_12601);
xnor U13253 (N_13253,N_12508,N_12688);
or U13254 (N_13254,N_12551,N_12876);
nand U13255 (N_13255,N_12839,N_12576);
nor U13256 (N_13256,N_12879,N_12850);
and U13257 (N_13257,N_12645,N_12680);
and U13258 (N_13258,N_12986,N_12521);
or U13259 (N_13259,N_12765,N_12842);
or U13260 (N_13260,N_12895,N_12761);
or U13261 (N_13261,N_12531,N_12766);
nand U13262 (N_13262,N_12637,N_12683);
nand U13263 (N_13263,N_12712,N_12764);
and U13264 (N_13264,N_12827,N_12904);
or U13265 (N_13265,N_12639,N_12775);
or U13266 (N_13266,N_12501,N_12825);
and U13267 (N_13267,N_12936,N_12958);
or U13268 (N_13268,N_12963,N_12633);
nor U13269 (N_13269,N_12971,N_12557);
and U13270 (N_13270,N_12582,N_12731);
or U13271 (N_13271,N_12688,N_12923);
and U13272 (N_13272,N_12609,N_12582);
or U13273 (N_13273,N_12988,N_12722);
xor U13274 (N_13274,N_12648,N_12794);
nor U13275 (N_13275,N_12932,N_12954);
nand U13276 (N_13276,N_12887,N_12666);
xor U13277 (N_13277,N_12722,N_12651);
and U13278 (N_13278,N_12714,N_12935);
nand U13279 (N_13279,N_12921,N_12582);
nor U13280 (N_13280,N_12544,N_12631);
or U13281 (N_13281,N_12913,N_12742);
xnor U13282 (N_13282,N_12846,N_12813);
and U13283 (N_13283,N_12593,N_12888);
or U13284 (N_13284,N_12939,N_12531);
and U13285 (N_13285,N_12788,N_12687);
or U13286 (N_13286,N_12767,N_12913);
and U13287 (N_13287,N_12813,N_12516);
or U13288 (N_13288,N_12778,N_12844);
nand U13289 (N_13289,N_12878,N_12948);
nor U13290 (N_13290,N_12722,N_12603);
nand U13291 (N_13291,N_12691,N_12763);
nand U13292 (N_13292,N_12781,N_12521);
or U13293 (N_13293,N_12806,N_12519);
or U13294 (N_13294,N_12680,N_12791);
xor U13295 (N_13295,N_12977,N_12901);
or U13296 (N_13296,N_12907,N_12788);
and U13297 (N_13297,N_12647,N_12827);
xor U13298 (N_13298,N_12575,N_12873);
and U13299 (N_13299,N_12957,N_12971);
and U13300 (N_13300,N_12549,N_12952);
nand U13301 (N_13301,N_12849,N_12733);
nor U13302 (N_13302,N_12628,N_12734);
nor U13303 (N_13303,N_12759,N_12720);
nand U13304 (N_13304,N_12702,N_12996);
and U13305 (N_13305,N_12643,N_12670);
and U13306 (N_13306,N_12624,N_12610);
or U13307 (N_13307,N_12746,N_12963);
nor U13308 (N_13308,N_12606,N_12791);
nor U13309 (N_13309,N_12900,N_12549);
and U13310 (N_13310,N_12996,N_12918);
nor U13311 (N_13311,N_12519,N_12760);
xor U13312 (N_13312,N_12999,N_12501);
nor U13313 (N_13313,N_12701,N_12908);
xnor U13314 (N_13314,N_12626,N_12857);
nand U13315 (N_13315,N_12893,N_12771);
nand U13316 (N_13316,N_12791,N_12663);
xnor U13317 (N_13317,N_12811,N_12584);
nor U13318 (N_13318,N_12594,N_12541);
nor U13319 (N_13319,N_12865,N_12641);
and U13320 (N_13320,N_12646,N_12632);
or U13321 (N_13321,N_12688,N_12627);
xor U13322 (N_13322,N_12646,N_12991);
and U13323 (N_13323,N_12908,N_12887);
xnor U13324 (N_13324,N_12777,N_12800);
nor U13325 (N_13325,N_12963,N_12929);
or U13326 (N_13326,N_12655,N_12723);
or U13327 (N_13327,N_12817,N_12638);
and U13328 (N_13328,N_12595,N_12818);
nand U13329 (N_13329,N_12716,N_12750);
nand U13330 (N_13330,N_12896,N_12970);
or U13331 (N_13331,N_12787,N_12954);
and U13332 (N_13332,N_12683,N_12669);
nand U13333 (N_13333,N_12936,N_12701);
nand U13334 (N_13334,N_12991,N_12588);
nand U13335 (N_13335,N_12850,N_12690);
xor U13336 (N_13336,N_12638,N_12930);
nand U13337 (N_13337,N_12789,N_12519);
and U13338 (N_13338,N_12707,N_12547);
or U13339 (N_13339,N_12814,N_12553);
and U13340 (N_13340,N_12948,N_12786);
or U13341 (N_13341,N_12983,N_12875);
and U13342 (N_13342,N_12946,N_12972);
nor U13343 (N_13343,N_12746,N_12550);
nor U13344 (N_13344,N_12941,N_12968);
nor U13345 (N_13345,N_12941,N_12756);
or U13346 (N_13346,N_12844,N_12575);
nor U13347 (N_13347,N_12995,N_12659);
and U13348 (N_13348,N_12745,N_12609);
nor U13349 (N_13349,N_12955,N_12908);
and U13350 (N_13350,N_12558,N_12997);
and U13351 (N_13351,N_12987,N_12724);
and U13352 (N_13352,N_12558,N_12511);
xnor U13353 (N_13353,N_12850,N_12946);
and U13354 (N_13354,N_12580,N_12883);
or U13355 (N_13355,N_12989,N_12541);
nor U13356 (N_13356,N_12972,N_12519);
and U13357 (N_13357,N_12932,N_12924);
nand U13358 (N_13358,N_12901,N_12564);
xnor U13359 (N_13359,N_12935,N_12726);
and U13360 (N_13360,N_12786,N_12603);
or U13361 (N_13361,N_12751,N_12864);
nand U13362 (N_13362,N_12952,N_12957);
and U13363 (N_13363,N_12822,N_12781);
nor U13364 (N_13364,N_12524,N_12655);
and U13365 (N_13365,N_12515,N_12849);
nor U13366 (N_13366,N_12554,N_12764);
xor U13367 (N_13367,N_12988,N_12572);
nor U13368 (N_13368,N_12620,N_12929);
and U13369 (N_13369,N_12993,N_12740);
nor U13370 (N_13370,N_12950,N_12542);
nor U13371 (N_13371,N_12597,N_12506);
and U13372 (N_13372,N_12816,N_12930);
nor U13373 (N_13373,N_12607,N_12962);
nor U13374 (N_13374,N_12996,N_12686);
xnor U13375 (N_13375,N_12900,N_12569);
or U13376 (N_13376,N_12938,N_12817);
nand U13377 (N_13377,N_12699,N_12632);
nand U13378 (N_13378,N_12518,N_12783);
or U13379 (N_13379,N_12806,N_12830);
nor U13380 (N_13380,N_12745,N_12899);
and U13381 (N_13381,N_12781,N_12709);
nand U13382 (N_13382,N_12676,N_12516);
and U13383 (N_13383,N_12806,N_12973);
or U13384 (N_13384,N_12817,N_12526);
xor U13385 (N_13385,N_12883,N_12720);
and U13386 (N_13386,N_12535,N_12973);
nand U13387 (N_13387,N_12994,N_12829);
nor U13388 (N_13388,N_12777,N_12729);
nand U13389 (N_13389,N_12753,N_12773);
nand U13390 (N_13390,N_12908,N_12685);
nor U13391 (N_13391,N_12713,N_12800);
nor U13392 (N_13392,N_12507,N_12531);
or U13393 (N_13393,N_12531,N_12833);
nor U13394 (N_13394,N_12741,N_12776);
or U13395 (N_13395,N_12761,N_12745);
or U13396 (N_13396,N_12758,N_12916);
nand U13397 (N_13397,N_12932,N_12578);
nand U13398 (N_13398,N_12867,N_12956);
nand U13399 (N_13399,N_12749,N_12922);
nand U13400 (N_13400,N_12863,N_12945);
nor U13401 (N_13401,N_12847,N_12826);
nor U13402 (N_13402,N_12832,N_12920);
nand U13403 (N_13403,N_12700,N_12882);
and U13404 (N_13404,N_12695,N_12624);
nand U13405 (N_13405,N_12524,N_12824);
or U13406 (N_13406,N_12819,N_12824);
nand U13407 (N_13407,N_12744,N_12537);
or U13408 (N_13408,N_12967,N_12760);
nor U13409 (N_13409,N_12866,N_12641);
or U13410 (N_13410,N_12571,N_12916);
and U13411 (N_13411,N_12725,N_12519);
nand U13412 (N_13412,N_12887,N_12569);
or U13413 (N_13413,N_12807,N_12524);
or U13414 (N_13414,N_12561,N_12628);
xor U13415 (N_13415,N_12668,N_12795);
nand U13416 (N_13416,N_12832,N_12851);
xnor U13417 (N_13417,N_12929,N_12684);
and U13418 (N_13418,N_12822,N_12715);
and U13419 (N_13419,N_12990,N_12979);
nor U13420 (N_13420,N_12570,N_12776);
or U13421 (N_13421,N_12608,N_12537);
nor U13422 (N_13422,N_12957,N_12522);
nor U13423 (N_13423,N_12893,N_12698);
or U13424 (N_13424,N_12679,N_12716);
and U13425 (N_13425,N_12974,N_12557);
nand U13426 (N_13426,N_12552,N_12805);
and U13427 (N_13427,N_12635,N_12899);
nand U13428 (N_13428,N_12657,N_12991);
nand U13429 (N_13429,N_12515,N_12639);
or U13430 (N_13430,N_12730,N_12817);
nand U13431 (N_13431,N_12853,N_12693);
nor U13432 (N_13432,N_12923,N_12804);
nor U13433 (N_13433,N_12857,N_12739);
nor U13434 (N_13434,N_12583,N_12761);
nand U13435 (N_13435,N_12782,N_12789);
or U13436 (N_13436,N_12555,N_12744);
nor U13437 (N_13437,N_12538,N_12629);
and U13438 (N_13438,N_12604,N_12902);
xor U13439 (N_13439,N_12843,N_12670);
or U13440 (N_13440,N_12926,N_12577);
or U13441 (N_13441,N_12521,N_12525);
or U13442 (N_13442,N_12577,N_12888);
nor U13443 (N_13443,N_12800,N_12813);
or U13444 (N_13444,N_12806,N_12805);
and U13445 (N_13445,N_12785,N_12770);
nand U13446 (N_13446,N_12679,N_12780);
and U13447 (N_13447,N_12770,N_12958);
nor U13448 (N_13448,N_12536,N_12977);
and U13449 (N_13449,N_12863,N_12701);
nor U13450 (N_13450,N_12897,N_12956);
and U13451 (N_13451,N_12973,N_12710);
and U13452 (N_13452,N_12538,N_12997);
or U13453 (N_13453,N_12714,N_12934);
nor U13454 (N_13454,N_12829,N_12626);
or U13455 (N_13455,N_12834,N_12864);
or U13456 (N_13456,N_12687,N_12997);
and U13457 (N_13457,N_12632,N_12970);
nor U13458 (N_13458,N_12806,N_12944);
nor U13459 (N_13459,N_12946,N_12967);
or U13460 (N_13460,N_12874,N_12760);
and U13461 (N_13461,N_12876,N_12917);
or U13462 (N_13462,N_12819,N_12823);
or U13463 (N_13463,N_12555,N_12780);
and U13464 (N_13464,N_12744,N_12747);
or U13465 (N_13465,N_12511,N_12568);
and U13466 (N_13466,N_12530,N_12802);
xor U13467 (N_13467,N_12985,N_12921);
nor U13468 (N_13468,N_12954,N_12941);
nand U13469 (N_13469,N_12699,N_12697);
and U13470 (N_13470,N_12677,N_12838);
nor U13471 (N_13471,N_12796,N_12947);
and U13472 (N_13472,N_12847,N_12709);
nor U13473 (N_13473,N_12965,N_12941);
nor U13474 (N_13474,N_12686,N_12963);
or U13475 (N_13475,N_12880,N_12730);
and U13476 (N_13476,N_12506,N_12553);
xor U13477 (N_13477,N_12841,N_12883);
nand U13478 (N_13478,N_12674,N_12685);
and U13479 (N_13479,N_12511,N_12743);
nand U13480 (N_13480,N_12584,N_12940);
nand U13481 (N_13481,N_12973,N_12745);
nor U13482 (N_13482,N_12604,N_12670);
nand U13483 (N_13483,N_12849,N_12929);
or U13484 (N_13484,N_12524,N_12948);
nand U13485 (N_13485,N_12632,N_12834);
and U13486 (N_13486,N_12659,N_12634);
and U13487 (N_13487,N_12730,N_12971);
or U13488 (N_13488,N_12773,N_12655);
or U13489 (N_13489,N_12694,N_12508);
or U13490 (N_13490,N_12668,N_12978);
nor U13491 (N_13491,N_12874,N_12820);
and U13492 (N_13492,N_12500,N_12710);
xor U13493 (N_13493,N_12885,N_12912);
and U13494 (N_13494,N_12524,N_12611);
and U13495 (N_13495,N_12900,N_12835);
and U13496 (N_13496,N_12620,N_12749);
xor U13497 (N_13497,N_12958,N_12691);
xnor U13498 (N_13498,N_12761,N_12770);
nor U13499 (N_13499,N_12690,N_12596);
nor U13500 (N_13500,N_13182,N_13312);
nand U13501 (N_13501,N_13446,N_13435);
xnor U13502 (N_13502,N_13056,N_13403);
xnor U13503 (N_13503,N_13013,N_13358);
or U13504 (N_13504,N_13231,N_13443);
and U13505 (N_13505,N_13427,N_13163);
or U13506 (N_13506,N_13476,N_13139);
and U13507 (N_13507,N_13114,N_13481);
or U13508 (N_13508,N_13043,N_13214);
or U13509 (N_13509,N_13428,N_13256);
or U13510 (N_13510,N_13108,N_13130);
or U13511 (N_13511,N_13384,N_13453);
nand U13512 (N_13512,N_13237,N_13293);
nand U13513 (N_13513,N_13407,N_13316);
and U13514 (N_13514,N_13018,N_13101);
xnor U13515 (N_13515,N_13236,N_13172);
and U13516 (N_13516,N_13092,N_13194);
and U13517 (N_13517,N_13457,N_13333);
nand U13518 (N_13518,N_13153,N_13195);
and U13519 (N_13519,N_13015,N_13110);
nand U13520 (N_13520,N_13386,N_13368);
and U13521 (N_13521,N_13118,N_13210);
nand U13522 (N_13522,N_13440,N_13417);
and U13523 (N_13523,N_13259,N_13105);
or U13524 (N_13524,N_13454,N_13257);
nor U13525 (N_13525,N_13419,N_13411);
or U13526 (N_13526,N_13176,N_13267);
and U13527 (N_13527,N_13164,N_13205);
nand U13528 (N_13528,N_13337,N_13171);
and U13529 (N_13529,N_13348,N_13306);
nor U13530 (N_13530,N_13218,N_13211);
and U13531 (N_13531,N_13054,N_13044);
nand U13532 (N_13532,N_13160,N_13238);
nand U13533 (N_13533,N_13396,N_13438);
nor U13534 (N_13534,N_13288,N_13321);
nor U13535 (N_13535,N_13065,N_13280);
nand U13536 (N_13536,N_13497,N_13014);
or U13537 (N_13537,N_13351,N_13019);
and U13538 (N_13538,N_13399,N_13169);
nor U13539 (N_13539,N_13080,N_13330);
nor U13540 (N_13540,N_13212,N_13088);
and U13541 (N_13541,N_13391,N_13034);
and U13542 (N_13542,N_13048,N_13405);
or U13543 (N_13543,N_13038,N_13016);
nand U13544 (N_13544,N_13024,N_13128);
nor U13545 (N_13545,N_13416,N_13494);
nand U13546 (N_13546,N_13314,N_13303);
nor U13547 (N_13547,N_13091,N_13489);
nand U13548 (N_13548,N_13388,N_13049);
nor U13549 (N_13549,N_13402,N_13045);
nand U13550 (N_13550,N_13098,N_13145);
or U13551 (N_13551,N_13372,N_13265);
nor U13552 (N_13552,N_13243,N_13371);
nor U13553 (N_13553,N_13332,N_13469);
nor U13554 (N_13554,N_13367,N_13357);
or U13555 (N_13555,N_13126,N_13228);
nor U13556 (N_13556,N_13285,N_13463);
xnor U13557 (N_13557,N_13102,N_13241);
or U13558 (N_13558,N_13227,N_13437);
nor U13559 (N_13559,N_13274,N_13156);
and U13560 (N_13560,N_13178,N_13242);
or U13561 (N_13561,N_13203,N_13485);
nand U13562 (N_13562,N_13011,N_13269);
or U13563 (N_13563,N_13290,N_13363);
and U13564 (N_13564,N_13099,N_13030);
nand U13565 (N_13565,N_13134,N_13006);
or U13566 (N_13566,N_13374,N_13159);
nor U13567 (N_13567,N_13076,N_13150);
nand U13568 (N_13568,N_13246,N_13467);
nor U13569 (N_13569,N_13071,N_13422);
and U13570 (N_13570,N_13254,N_13359);
nand U13571 (N_13571,N_13122,N_13155);
and U13572 (N_13572,N_13345,N_13455);
xor U13573 (N_13573,N_13425,N_13042);
or U13574 (N_13574,N_13310,N_13389);
or U13575 (N_13575,N_13249,N_13410);
nor U13576 (N_13576,N_13373,N_13025);
and U13577 (N_13577,N_13050,N_13005);
nand U13578 (N_13578,N_13251,N_13202);
or U13579 (N_13579,N_13339,N_13433);
nand U13580 (N_13580,N_13199,N_13375);
and U13581 (N_13581,N_13093,N_13325);
nand U13582 (N_13582,N_13304,N_13039);
nand U13583 (N_13583,N_13127,N_13041);
or U13584 (N_13584,N_13225,N_13247);
nor U13585 (N_13585,N_13135,N_13083);
nor U13586 (N_13586,N_13335,N_13395);
xnor U13587 (N_13587,N_13142,N_13221);
and U13588 (N_13588,N_13406,N_13322);
nor U13589 (N_13589,N_13307,N_13344);
and U13590 (N_13590,N_13356,N_13215);
or U13591 (N_13591,N_13341,N_13029);
or U13592 (N_13592,N_13046,N_13033);
nand U13593 (N_13593,N_13106,N_13477);
nor U13594 (N_13594,N_13270,N_13370);
nand U13595 (N_13595,N_13378,N_13491);
or U13596 (N_13596,N_13380,N_13021);
or U13597 (N_13597,N_13097,N_13318);
and U13598 (N_13598,N_13198,N_13184);
nor U13599 (N_13599,N_13423,N_13057);
or U13600 (N_13600,N_13085,N_13327);
and U13601 (N_13601,N_13266,N_13369);
nand U13602 (N_13602,N_13229,N_13431);
xor U13603 (N_13603,N_13355,N_13008);
and U13604 (N_13604,N_13291,N_13323);
nand U13605 (N_13605,N_13354,N_13415);
and U13606 (N_13606,N_13094,N_13320);
and U13607 (N_13607,N_13051,N_13188);
or U13608 (N_13608,N_13035,N_13209);
or U13609 (N_13609,N_13460,N_13398);
nand U13610 (N_13610,N_13353,N_13474);
or U13611 (N_13611,N_13170,N_13275);
xnor U13612 (N_13612,N_13158,N_13343);
nand U13613 (N_13613,N_13179,N_13107);
nand U13614 (N_13614,N_13413,N_13003);
nand U13615 (N_13615,N_13360,N_13032);
xnor U13616 (N_13616,N_13338,N_13103);
and U13617 (N_13617,N_13404,N_13067);
or U13618 (N_13618,N_13064,N_13480);
and U13619 (N_13619,N_13223,N_13297);
or U13620 (N_13620,N_13078,N_13289);
or U13621 (N_13621,N_13424,N_13429);
nor U13622 (N_13622,N_13119,N_13408);
and U13623 (N_13623,N_13475,N_13296);
and U13624 (N_13624,N_13426,N_13100);
or U13625 (N_13625,N_13084,N_13452);
nand U13626 (N_13626,N_13295,N_13361);
nand U13627 (N_13627,N_13077,N_13448);
xnor U13628 (N_13628,N_13109,N_13272);
and U13629 (N_13629,N_13189,N_13152);
nand U13630 (N_13630,N_13020,N_13143);
nor U13631 (N_13631,N_13090,N_13409);
or U13632 (N_13632,N_13261,N_13095);
nand U13633 (N_13633,N_13492,N_13149);
nor U13634 (N_13634,N_13418,N_13141);
nand U13635 (N_13635,N_13233,N_13283);
nor U13636 (N_13636,N_13362,N_13070);
nand U13637 (N_13637,N_13204,N_13068);
nor U13638 (N_13638,N_13273,N_13493);
nor U13639 (N_13639,N_13124,N_13173);
and U13640 (N_13640,N_13074,N_13401);
nor U13641 (N_13641,N_13187,N_13089);
and U13642 (N_13642,N_13047,N_13271);
and U13643 (N_13643,N_13282,N_13447);
and U13644 (N_13644,N_13226,N_13007);
or U13645 (N_13645,N_13319,N_13311);
or U13646 (N_13646,N_13287,N_13420);
nand U13647 (N_13647,N_13326,N_13400);
nor U13648 (N_13648,N_13393,N_13352);
and U13649 (N_13649,N_13430,N_13060);
or U13650 (N_13650,N_13000,N_13444);
and U13651 (N_13651,N_13436,N_13346);
nand U13652 (N_13652,N_13234,N_13317);
or U13653 (N_13653,N_13232,N_13133);
or U13654 (N_13654,N_13462,N_13036);
and U13655 (N_13655,N_13313,N_13387);
and U13656 (N_13656,N_13115,N_13181);
and U13657 (N_13657,N_13147,N_13349);
nand U13658 (N_13658,N_13451,N_13366);
nor U13659 (N_13659,N_13309,N_13412);
or U13660 (N_13660,N_13081,N_13377);
nand U13661 (N_13661,N_13144,N_13058);
or U13662 (N_13662,N_13120,N_13157);
xnor U13663 (N_13663,N_13300,N_13031);
nand U13664 (N_13664,N_13023,N_13434);
or U13665 (N_13665,N_13059,N_13264);
xor U13666 (N_13666,N_13465,N_13298);
nand U13667 (N_13667,N_13347,N_13331);
nor U13668 (N_13668,N_13301,N_13113);
or U13669 (N_13669,N_13329,N_13220);
xnor U13670 (N_13670,N_13482,N_13383);
and U13671 (N_13671,N_13012,N_13186);
nor U13672 (N_13672,N_13161,N_13342);
nor U13673 (N_13673,N_13488,N_13162);
or U13674 (N_13674,N_13394,N_13069);
nor U13675 (N_13675,N_13487,N_13062);
nor U13676 (N_13676,N_13286,N_13255);
or U13677 (N_13677,N_13192,N_13305);
and U13678 (N_13678,N_13473,N_13166);
or U13679 (N_13679,N_13137,N_13498);
or U13680 (N_13680,N_13154,N_13117);
and U13681 (N_13681,N_13111,N_13200);
or U13682 (N_13682,N_13196,N_13483);
nand U13683 (N_13683,N_13224,N_13219);
nand U13684 (N_13684,N_13096,N_13464);
nand U13685 (N_13685,N_13365,N_13207);
xor U13686 (N_13686,N_13138,N_13441);
nand U13687 (N_13687,N_13206,N_13121);
and U13688 (N_13688,N_13063,N_13193);
and U13689 (N_13689,N_13364,N_13471);
xnor U13690 (N_13690,N_13250,N_13239);
nor U13691 (N_13691,N_13284,N_13439);
nor U13692 (N_13692,N_13116,N_13277);
and U13693 (N_13693,N_13168,N_13073);
xor U13694 (N_13694,N_13148,N_13175);
nor U13695 (N_13695,N_13328,N_13230);
nor U13696 (N_13696,N_13197,N_13449);
nand U13697 (N_13697,N_13499,N_13026);
or U13698 (N_13698,N_13129,N_13299);
nand U13699 (N_13699,N_13268,N_13140);
nand U13700 (N_13700,N_13104,N_13087);
or U13701 (N_13701,N_13478,N_13191);
and U13702 (N_13702,N_13379,N_13177);
or U13703 (N_13703,N_13132,N_13336);
and U13704 (N_13704,N_13174,N_13252);
nor U13705 (N_13705,N_13079,N_13052);
or U13706 (N_13706,N_13053,N_13442);
nor U13707 (N_13707,N_13421,N_13414);
or U13708 (N_13708,N_13082,N_13479);
and U13709 (N_13709,N_13240,N_13294);
xnor U13710 (N_13710,N_13302,N_13213);
or U13711 (N_13711,N_13496,N_13456);
nand U13712 (N_13712,N_13004,N_13468);
nor U13713 (N_13713,N_13131,N_13165);
nor U13714 (N_13714,N_13222,N_13245);
or U13715 (N_13715,N_13248,N_13263);
and U13716 (N_13716,N_13017,N_13185);
and U13717 (N_13717,N_13040,N_13180);
and U13718 (N_13718,N_13397,N_13390);
and U13719 (N_13719,N_13086,N_13385);
and U13720 (N_13720,N_13381,N_13075);
nor U13721 (N_13721,N_13125,N_13055);
and U13722 (N_13722,N_13276,N_13279);
nor U13723 (N_13723,N_13486,N_13002);
and U13724 (N_13724,N_13072,N_13190);
and U13725 (N_13725,N_13472,N_13281);
and U13726 (N_13726,N_13037,N_13262);
or U13727 (N_13727,N_13470,N_13151);
xnor U13728 (N_13728,N_13217,N_13123);
nor U13729 (N_13729,N_13382,N_13308);
or U13730 (N_13730,N_13253,N_13292);
nand U13731 (N_13731,N_13484,N_13235);
nand U13732 (N_13732,N_13258,N_13216);
or U13733 (N_13733,N_13461,N_13027);
and U13734 (N_13734,N_13458,N_13167);
or U13735 (N_13735,N_13010,N_13445);
and U13736 (N_13736,N_13340,N_13450);
and U13737 (N_13737,N_13183,N_13432);
xnor U13738 (N_13738,N_13009,N_13459);
nor U13739 (N_13739,N_13376,N_13136);
and U13740 (N_13740,N_13146,N_13022);
nand U13741 (N_13741,N_13490,N_13028);
nand U13742 (N_13742,N_13350,N_13112);
xor U13743 (N_13743,N_13201,N_13278);
or U13744 (N_13744,N_13324,N_13495);
and U13745 (N_13745,N_13244,N_13066);
nand U13746 (N_13746,N_13061,N_13392);
or U13747 (N_13747,N_13466,N_13334);
nor U13748 (N_13748,N_13260,N_13001);
or U13749 (N_13749,N_13208,N_13315);
or U13750 (N_13750,N_13177,N_13422);
or U13751 (N_13751,N_13075,N_13090);
or U13752 (N_13752,N_13216,N_13083);
or U13753 (N_13753,N_13090,N_13001);
xnor U13754 (N_13754,N_13206,N_13151);
nand U13755 (N_13755,N_13483,N_13290);
nand U13756 (N_13756,N_13019,N_13100);
nor U13757 (N_13757,N_13369,N_13077);
nor U13758 (N_13758,N_13484,N_13407);
or U13759 (N_13759,N_13136,N_13384);
and U13760 (N_13760,N_13337,N_13226);
and U13761 (N_13761,N_13115,N_13276);
nor U13762 (N_13762,N_13004,N_13267);
or U13763 (N_13763,N_13304,N_13403);
nor U13764 (N_13764,N_13465,N_13308);
nor U13765 (N_13765,N_13016,N_13418);
xor U13766 (N_13766,N_13022,N_13023);
nand U13767 (N_13767,N_13078,N_13211);
xnor U13768 (N_13768,N_13061,N_13198);
nand U13769 (N_13769,N_13122,N_13049);
and U13770 (N_13770,N_13235,N_13090);
or U13771 (N_13771,N_13498,N_13108);
and U13772 (N_13772,N_13225,N_13429);
nand U13773 (N_13773,N_13102,N_13375);
and U13774 (N_13774,N_13447,N_13005);
or U13775 (N_13775,N_13128,N_13291);
xnor U13776 (N_13776,N_13273,N_13310);
xor U13777 (N_13777,N_13045,N_13261);
nor U13778 (N_13778,N_13143,N_13299);
nor U13779 (N_13779,N_13175,N_13128);
and U13780 (N_13780,N_13006,N_13336);
nand U13781 (N_13781,N_13465,N_13335);
or U13782 (N_13782,N_13406,N_13190);
nor U13783 (N_13783,N_13261,N_13352);
and U13784 (N_13784,N_13368,N_13098);
and U13785 (N_13785,N_13299,N_13367);
and U13786 (N_13786,N_13223,N_13456);
nand U13787 (N_13787,N_13179,N_13186);
and U13788 (N_13788,N_13322,N_13378);
and U13789 (N_13789,N_13135,N_13145);
xor U13790 (N_13790,N_13267,N_13275);
nor U13791 (N_13791,N_13359,N_13069);
nor U13792 (N_13792,N_13451,N_13235);
nor U13793 (N_13793,N_13123,N_13060);
nor U13794 (N_13794,N_13087,N_13007);
nand U13795 (N_13795,N_13243,N_13480);
nand U13796 (N_13796,N_13031,N_13352);
xnor U13797 (N_13797,N_13072,N_13184);
nor U13798 (N_13798,N_13065,N_13098);
xnor U13799 (N_13799,N_13383,N_13259);
or U13800 (N_13800,N_13190,N_13187);
nand U13801 (N_13801,N_13092,N_13086);
nand U13802 (N_13802,N_13423,N_13182);
and U13803 (N_13803,N_13032,N_13054);
or U13804 (N_13804,N_13281,N_13366);
nand U13805 (N_13805,N_13335,N_13119);
or U13806 (N_13806,N_13124,N_13066);
nor U13807 (N_13807,N_13455,N_13056);
nand U13808 (N_13808,N_13221,N_13048);
xnor U13809 (N_13809,N_13405,N_13035);
or U13810 (N_13810,N_13006,N_13461);
or U13811 (N_13811,N_13401,N_13459);
nand U13812 (N_13812,N_13063,N_13173);
nor U13813 (N_13813,N_13121,N_13466);
nand U13814 (N_13814,N_13315,N_13078);
or U13815 (N_13815,N_13055,N_13193);
nand U13816 (N_13816,N_13257,N_13225);
or U13817 (N_13817,N_13040,N_13178);
nor U13818 (N_13818,N_13439,N_13382);
nand U13819 (N_13819,N_13341,N_13237);
or U13820 (N_13820,N_13470,N_13314);
nor U13821 (N_13821,N_13401,N_13328);
nor U13822 (N_13822,N_13133,N_13156);
nand U13823 (N_13823,N_13060,N_13371);
or U13824 (N_13824,N_13355,N_13025);
xnor U13825 (N_13825,N_13345,N_13416);
and U13826 (N_13826,N_13301,N_13334);
and U13827 (N_13827,N_13480,N_13438);
nand U13828 (N_13828,N_13398,N_13382);
or U13829 (N_13829,N_13210,N_13216);
nor U13830 (N_13830,N_13097,N_13246);
nand U13831 (N_13831,N_13460,N_13013);
and U13832 (N_13832,N_13287,N_13118);
and U13833 (N_13833,N_13355,N_13143);
nand U13834 (N_13834,N_13180,N_13050);
or U13835 (N_13835,N_13305,N_13165);
nor U13836 (N_13836,N_13123,N_13447);
nor U13837 (N_13837,N_13463,N_13109);
xnor U13838 (N_13838,N_13317,N_13354);
nor U13839 (N_13839,N_13016,N_13445);
xor U13840 (N_13840,N_13209,N_13317);
nand U13841 (N_13841,N_13427,N_13360);
or U13842 (N_13842,N_13476,N_13466);
nor U13843 (N_13843,N_13358,N_13307);
or U13844 (N_13844,N_13220,N_13201);
xor U13845 (N_13845,N_13224,N_13397);
xor U13846 (N_13846,N_13084,N_13304);
or U13847 (N_13847,N_13373,N_13398);
nand U13848 (N_13848,N_13208,N_13410);
and U13849 (N_13849,N_13365,N_13199);
and U13850 (N_13850,N_13078,N_13237);
and U13851 (N_13851,N_13094,N_13112);
nand U13852 (N_13852,N_13025,N_13149);
or U13853 (N_13853,N_13273,N_13166);
nor U13854 (N_13854,N_13409,N_13317);
nor U13855 (N_13855,N_13464,N_13170);
nor U13856 (N_13856,N_13452,N_13109);
xor U13857 (N_13857,N_13489,N_13032);
nor U13858 (N_13858,N_13078,N_13207);
nand U13859 (N_13859,N_13406,N_13402);
and U13860 (N_13860,N_13415,N_13459);
and U13861 (N_13861,N_13294,N_13238);
nor U13862 (N_13862,N_13288,N_13156);
nand U13863 (N_13863,N_13000,N_13098);
and U13864 (N_13864,N_13304,N_13140);
nor U13865 (N_13865,N_13155,N_13089);
nor U13866 (N_13866,N_13236,N_13048);
or U13867 (N_13867,N_13307,N_13331);
nand U13868 (N_13868,N_13170,N_13289);
or U13869 (N_13869,N_13001,N_13369);
or U13870 (N_13870,N_13242,N_13350);
or U13871 (N_13871,N_13446,N_13245);
xor U13872 (N_13872,N_13465,N_13197);
or U13873 (N_13873,N_13221,N_13115);
nand U13874 (N_13874,N_13439,N_13116);
and U13875 (N_13875,N_13299,N_13399);
nand U13876 (N_13876,N_13087,N_13234);
and U13877 (N_13877,N_13328,N_13044);
and U13878 (N_13878,N_13227,N_13006);
xor U13879 (N_13879,N_13202,N_13299);
or U13880 (N_13880,N_13448,N_13343);
nor U13881 (N_13881,N_13455,N_13306);
nand U13882 (N_13882,N_13477,N_13191);
or U13883 (N_13883,N_13214,N_13212);
and U13884 (N_13884,N_13158,N_13487);
or U13885 (N_13885,N_13436,N_13233);
nand U13886 (N_13886,N_13406,N_13015);
and U13887 (N_13887,N_13465,N_13058);
and U13888 (N_13888,N_13295,N_13071);
or U13889 (N_13889,N_13016,N_13387);
nor U13890 (N_13890,N_13295,N_13211);
xnor U13891 (N_13891,N_13468,N_13445);
nor U13892 (N_13892,N_13301,N_13036);
or U13893 (N_13893,N_13092,N_13293);
nand U13894 (N_13894,N_13366,N_13145);
nor U13895 (N_13895,N_13168,N_13042);
and U13896 (N_13896,N_13412,N_13473);
nor U13897 (N_13897,N_13167,N_13479);
or U13898 (N_13898,N_13499,N_13001);
and U13899 (N_13899,N_13089,N_13099);
or U13900 (N_13900,N_13230,N_13355);
or U13901 (N_13901,N_13079,N_13237);
nor U13902 (N_13902,N_13010,N_13182);
and U13903 (N_13903,N_13232,N_13261);
or U13904 (N_13904,N_13437,N_13360);
and U13905 (N_13905,N_13012,N_13059);
nand U13906 (N_13906,N_13111,N_13303);
or U13907 (N_13907,N_13163,N_13399);
nand U13908 (N_13908,N_13145,N_13094);
xor U13909 (N_13909,N_13156,N_13408);
and U13910 (N_13910,N_13283,N_13482);
or U13911 (N_13911,N_13322,N_13282);
nor U13912 (N_13912,N_13148,N_13118);
nand U13913 (N_13913,N_13306,N_13106);
or U13914 (N_13914,N_13021,N_13246);
and U13915 (N_13915,N_13099,N_13272);
and U13916 (N_13916,N_13354,N_13198);
nor U13917 (N_13917,N_13140,N_13029);
and U13918 (N_13918,N_13290,N_13104);
or U13919 (N_13919,N_13232,N_13284);
nor U13920 (N_13920,N_13436,N_13026);
or U13921 (N_13921,N_13363,N_13082);
or U13922 (N_13922,N_13015,N_13168);
or U13923 (N_13923,N_13087,N_13408);
or U13924 (N_13924,N_13480,N_13053);
or U13925 (N_13925,N_13420,N_13302);
and U13926 (N_13926,N_13423,N_13061);
and U13927 (N_13927,N_13143,N_13099);
nand U13928 (N_13928,N_13437,N_13380);
or U13929 (N_13929,N_13365,N_13286);
or U13930 (N_13930,N_13433,N_13357);
nor U13931 (N_13931,N_13116,N_13097);
or U13932 (N_13932,N_13247,N_13149);
and U13933 (N_13933,N_13096,N_13125);
or U13934 (N_13934,N_13050,N_13204);
nand U13935 (N_13935,N_13469,N_13105);
and U13936 (N_13936,N_13399,N_13137);
nand U13937 (N_13937,N_13271,N_13221);
and U13938 (N_13938,N_13369,N_13096);
nand U13939 (N_13939,N_13058,N_13220);
and U13940 (N_13940,N_13068,N_13106);
nand U13941 (N_13941,N_13059,N_13343);
xnor U13942 (N_13942,N_13332,N_13393);
xnor U13943 (N_13943,N_13338,N_13170);
or U13944 (N_13944,N_13323,N_13463);
nand U13945 (N_13945,N_13360,N_13200);
xor U13946 (N_13946,N_13446,N_13367);
nand U13947 (N_13947,N_13453,N_13007);
nor U13948 (N_13948,N_13223,N_13258);
nand U13949 (N_13949,N_13403,N_13469);
xor U13950 (N_13950,N_13196,N_13369);
xnor U13951 (N_13951,N_13332,N_13047);
or U13952 (N_13952,N_13001,N_13055);
nand U13953 (N_13953,N_13088,N_13471);
xnor U13954 (N_13954,N_13394,N_13329);
nand U13955 (N_13955,N_13173,N_13348);
or U13956 (N_13956,N_13195,N_13469);
and U13957 (N_13957,N_13157,N_13063);
nor U13958 (N_13958,N_13499,N_13235);
or U13959 (N_13959,N_13476,N_13004);
nor U13960 (N_13960,N_13255,N_13063);
or U13961 (N_13961,N_13443,N_13283);
or U13962 (N_13962,N_13250,N_13052);
xor U13963 (N_13963,N_13464,N_13193);
or U13964 (N_13964,N_13480,N_13418);
or U13965 (N_13965,N_13339,N_13340);
and U13966 (N_13966,N_13313,N_13370);
or U13967 (N_13967,N_13240,N_13499);
nor U13968 (N_13968,N_13444,N_13388);
nor U13969 (N_13969,N_13467,N_13121);
xor U13970 (N_13970,N_13250,N_13463);
and U13971 (N_13971,N_13101,N_13114);
nand U13972 (N_13972,N_13365,N_13476);
or U13973 (N_13973,N_13015,N_13066);
nand U13974 (N_13974,N_13349,N_13180);
nand U13975 (N_13975,N_13244,N_13250);
nand U13976 (N_13976,N_13022,N_13204);
nand U13977 (N_13977,N_13294,N_13270);
and U13978 (N_13978,N_13354,N_13146);
nand U13979 (N_13979,N_13006,N_13352);
or U13980 (N_13980,N_13060,N_13009);
and U13981 (N_13981,N_13275,N_13279);
nor U13982 (N_13982,N_13413,N_13193);
or U13983 (N_13983,N_13190,N_13059);
nor U13984 (N_13984,N_13282,N_13135);
or U13985 (N_13985,N_13155,N_13040);
and U13986 (N_13986,N_13459,N_13482);
nor U13987 (N_13987,N_13226,N_13358);
nand U13988 (N_13988,N_13492,N_13249);
or U13989 (N_13989,N_13097,N_13270);
nand U13990 (N_13990,N_13086,N_13242);
nand U13991 (N_13991,N_13146,N_13261);
nor U13992 (N_13992,N_13376,N_13076);
nor U13993 (N_13993,N_13458,N_13180);
nand U13994 (N_13994,N_13455,N_13027);
xor U13995 (N_13995,N_13212,N_13381);
and U13996 (N_13996,N_13099,N_13366);
nor U13997 (N_13997,N_13144,N_13313);
nor U13998 (N_13998,N_13067,N_13423);
xnor U13999 (N_13999,N_13011,N_13373);
nand U14000 (N_14000,N_13731,N_13863);
xor U14001 (N_14001,N_13711,N_13745);
nor U14002 (N_14002,N_13852,N_13733);
nor U14003 (N_14003,N_13803,N_13599);
nor U14004 (N_14004,N_13565,N_13897);
or U14005 (N_14005,N_13945,N_13635);
nor U14006 (N_14006,N_13646,N_13562);
xnor U14007 (N_14007,N_13984,N_13679);
nor U14008 (N_14008,N_13798,N_13630);
and U14009 (N_14009,N_13917,N_13967);
nor U14010 (N_14010,N_13796,N_13762);
and U14011 (N_14011,N_13775,N_13879);
and U14012 (N_14012,N_13842,N_13576);
xnor U14013 (N_14013,N_13765,N_13750);
nand U14014 (N_14014,N_13512,N_13979);
nor U14015 (N_14015,N_13870,N_13850);
and U14016 (N_14016,N_13608,N_13642);
nor U14017 (N_14017,N_13699,N_13986);
nor U14018 (N_14018,N_13799,N_13520);
xnor U14019 (N_14019,N_13563,N_13739);
nand U14020 (N_14020,N_13605,N_13972);
nor U14021 (N_14021,N_13684,N_13742);
nand U14022 (N_14022,N_13812,N_13991);
nor U14023 (N_14023,N_13736,N_13804);
or U14024 (N_14024,N_13516,N_13880);
or U14025 (N_14025,N_13710,N_13557);
nor U14026 (N_14026,N_13550,N_13906);
and U14027 (N_14027,N_13881,N_13696);
nand U14028 (N_14028,N_13993,N_13769);
nor U14029 (N_14029,N_13566,N_13729);
nor U14030 (N_14030,N_13839,N_13524);
nand U14031 (N_14031,N_13607,N_13657);
nor U14032 (N_14032,N_13586,N_13820);
nor U14033 (N_14033,N_13509,N_13723);
nor U14034 (N_14034,N_13521,N_13781);
nand U14035 (N_14035,N_13929,N_13921);
nor U14036 (N_14036,N_13797,N_13728);
xor U14037 (N_14037,N_13939,N_13694);
nand U14038 (N_14038,N_13584,N_13808);
or U14039 (N_14039,N_13625,N_13761);
or U14040 (N_14040,N_13636,N_13553);
nand U14041 (N_14041,N_13779,N_13743);
or U14042 (N_14042,N_13949,N_13577);
nor U14043 (N_14043,N_13958,N_13505);
nor U14044 (N_14044,N_13735,N_13827);
and U14045 (N_14045,N_13545,N_13611);
nor U14046 (N_14046,N_13994,N_13866);
and U14047 (N_14047,N_13914,N_13836);
xnor U14048 (N_14048,N_13670,N_13551);
or U14049 (N_14049,N_13574,N_13571);
nor U14050 (N_14050,N_13932,N_13946);
xor U14051 (N_14051,N_13559,N_13513);
and U14052 (N_14052,N_13746,N_13811);
nand U14053 (N_14053,N_13867,N_13717);
nand U14054 (N_14054,N_13995,N_13954);
xnor U14055 (N_14055,N_13969,N_13629);
or U14056 (N_14056,N_13789,N_13920);
nand U14057 (N_14057,N_13843,N_13594);
nor U14058 (N_14058,N_13877,N_13856);
nor U14059 (N_14059,N_13996,N_13709);
nor U14060 (N_14060,N_13772,N_13909);
nand U14061 (N_14061,N_13971,N_13885);
xnor U14062 (N_14062,N_13515,N_13755);
xor U14063 (N_14063,N_13912,N_13685);
nor U14064 (N_14064,N_13924,N_13744);
and U14065 (N_14065,N_13616,N_13673);
and U14066 (N_14066,N_13809,N_13582);
or U14067 (N_14067,N_13508,N_13928);
and U14068 (N_14068,N_13502,N_13749);
and U14069 (N_14069,N_13900,N_13716);
xor U14070 (N_14070,N_13826,N_13919);
nor U14071 (N_14071,N_13990,N_13837);
or U14072 (N_14072,N_13544,N_13999);
or U14073 (N_14073,N_13955,N_13930);
or U14074 (N_14074,N_13978,N_13876);
or U14075 (N_14075,N_13648,N_13988);
and U14076 (N_14076,N_13591,N_13507);
xnor U14077 (N_14077,N_13787,N_13795);
or U14078 (N_14078,N_13878,N_13597);
or U14079 (N_14079,N_13698,N_13848);
nor U14080 (N_14080,N_13776,N_13677);
or U14081 (N_14081,N_13894,N_13974);
or U14082 (N_14082,N_13814,N_13889);
nand U14083 (N_14083,N_13976,N_13853);
nor U14084 (N_14084,N_13585,N_13985);
nor U14085 (N_14085,N_13663,N_13624);
nand U14086 (N_14086,N_13884,N_13588);
and U14087 (N_14087,N_13943,N_13834);
nor U14088 (N_14088,N_13501,N_13707);
or U14089 (N_14089,N_13832,N_13620);
or U14090 (N_14090,N_13655,N_13802);
or U14091 (N_14091,N_13977,N_13911);
and U14092 (N_14092,N_13653,N_13609);
and U14093 (N_14093,N_13732,N_13845);
nand U14094 (N_14094,N_13874,N_13727);
nand U14095 (N_14095,N_13665,N_13973);
nor U14096 (N_14096,N_13844,N_13752);
nor U14097 (N_14097,N_13862,N_13983);
nand U14098 (N_14098,N_13989,N_13855);
and U14099 (N_14099,N_13506,N_13641);
nor U14100 (N_14100,N_13822,N_13758);
nor U14101 (N_14101,N_13805,N_13619);
or U14102 (N_14102,N_13916,N_13966);
or U14103 (N_14103,N_13531,N_13887);
and U14104 (N_14104,N_13703,N_13664);
and U14105 (N_14105,N_13666,N_13982);
or U14106 (N_14106,N_13581,N_13888);
nor U14107 (N_14107,N_13659,N_13782);
nor U14108 (N_14108,N_13676,N_13712);
or U14109 (N_14109,N_13936,N_13534);
or U14110 (N_14110,N_13774,N_13975);
nor U14111 (N_14111,N_13819,N_13719);
nand U14112 (N_14112,N_13615,N_13764);
nor U14113 (N_14113,N_13823,N_13947);
xor U14114 (N_14114,N_13552,N_13904);
nand U14115 (N_14115,N_13957,N_13838);
nand U14116 (N_14116,N_13854,N_13841);
nand U14117 (N_14117,N_13937,N_13740);
or U14118 (N_14118,N_13548,N_13672);
or U14119 (N_14119,N_13691,N_13598);
or U14120 (N_14120,N_13640,N_13700);
xor U14121 (N_14121,N_13858,N_13800);
nand U14122 (N_14122,N_13747,N_13500);
and U14123 (N_14123,N_13835,N_13788);
nor U14124 (N_14124,N_13737,N_13575);
and U14125 (N_14125,N_13859,N_13759);
xor U14126 (N_14126,N_13915,N_13627);
nor U14127 (N_14127,N_13734,N_13540);
nand U14128 (N_14128,N_13942,N_13583);
xor U14129 (N_14129,N_13721,N_13997);
and U14130 (N_14130,N_13956,N_13535);
or U14131 (N_14131,N_13918,N_13567);
and U14132 (N_14132,N_13715,N_13960);
and U14133 (N_14133,N_13938,N_13546);
xnor U14134 (N_14134,N_13517,N_13623);
and U14135 (N_14135,N_13533,N_13898);
nand U14136 (N_14136,N_13952,N_13579);
nor U14137 (N_14137,N_13671,N_13871);
nor U14138 (N_14138,N_13667,N_13543);
xnor U14139 (N_14139,N_13702,N_13893);
and U14140 (N_14140,N_13748,N_13523);
nor U14141 (N_14141,N_13777,N_13662);
or U14142 (N_14142,N_13722,N_13519);
nand U14143 (N_14143,N_13829,N_13560);
nand U14144 (N_14144,N_13526,N_13687);
nor U14145 (N_14145,N_13821,N_13525);
nand U14146 (N_14146,N_13681,N_13780);
xnor U14147 (N_14147,N_13913,N_13669);
and U14148 (N_14148,N_13651,N_13965);
or U14149 (N_14149,N_13910,N_13892);
nand U14150 (N_14150,N_13632,N_13941);
nor U14151 (N_14151,N_13961,N_13596);
and U14152 (N_14152,N_13539,N_13908);
nor U14153 (N_14153,N_13660,N_13587);
or U14154 (N_14154,N_13547,N_13697);
xnor U14155 (N_14155,N_13935,N_13896);
or U14156 (N_14156,N_13753,N_13873);
and U14157 (N_14157,N_13510,N_13869);
and U14158 (N_14158,N_13725,N_13950);
and U14159 (N_14159,N_13922,N_13868);
or U14160 (N_14160,N_13778,N_13618);
and U14161 (N_14161,N_13578,N_13963);
or U14162 (N_14162,N_13791,N_13886);
and U14163 (N_14163,N_13654,N_13639);
and U14164 (N_14164,N_13708,N_13554);
xnor U14165 (N_14165,N_13860,N_13541);
or U14166 (N_14166,N_13652,N_13953);
and U14167 (N_14167,N_13527,N_13705);
xnor U14168 (N_14168,N_13573,N_13903);
nand U14169 (N_14169,N_13741,N_13785);
or U14170 (N_14170,N_13730,N_13561);
nor U14171 (N_14171,N_13818,N_13933);
xor U14172 (N_14172,N_13828,N_13650);
or U14173 (N_14173,N_13738,N_13987);
nand U14174 (N_14174,N_13951,N_13634);
and U14175 (N_14175,N_13682,N_13621);
nor U14176 (N_14176,N_13857,N_13612);
or U14177 (N_14177,N_13564,N_13601);
or U14178 (N_14178,N_13840,N_13714);
nor U14179 (N_14179,N_13628,N_13980);
and U14180 (N_14180,N_13542,N_13792);
and U14181 (N_14181,N_13556,N_13718);
nor U14182 (N_14182,N_13645,N_13720);
or U14183 (N_14183,N_13810,N_13763);
nand U14184 (N_14184,N_13661,N_13572);
nand U14185 (N_14185,N_13693,N_13688);
nor U14186 (N_14186,N_13701,N_13830);
and U14187 (N_14187,N_13883,N_13771);
nor U14188 (N_14188,N_13726,N_13849);
and U14189 (N_14189,N_13537,N_13593);
nand U14190 (N_14190,N_13606,N_13905);
or U14191 (N_14191,N_13600,N_13783);
nand U14192 (N_14192,N_13617,N_13847);
nand U14193 (N_14193,N_13530,N_13766);
or U14194 (N_14194,N_13570,N_13724);
nor U14195 (N_14195,N_13851,N_13807);
xor U14196 (N_14196,N_13647,N_13643);
and U14197 (N_14197,N_13658,N_13503);
and U14198 (N_14198,N_13861,N_13538);
and U14199 (N_14199,N_13754,N_13686);
or U14200 (N_14200,N_13675,N_13631);
nand U14201 (N_14201,N_13626,N_13794);
nor U14202 (N_14202,N_13695,N_13760);
nor U14203 (N_14203,N_13528,N_13603);
nor U14204 (N_14204,N_13981,N_13891);
nor U14205 (N_14205,N_13959,N_13518);
or U14206 (N_14206,N_13610,N_13622);
xor U14207 (N_14207,N_13637,N_13815);
nand U14208 (N_14208,N_13602,N_13784);
nor U14209 (N_14209,N_13757,N_13925);
or U14210 (N_14210,N_13690,N_13773);
or U14211 (N_14211,N_13899,N_13580);
nand U14212 (N_14212,N_13633,N_13767);
nand U14213 (N_14213,N_13680,N_13656);
and U14214 (N_14214,N_13901,N_13902);
nor U14215 (N_14215,N_13865,N_13522);
xnor U14216 (N_14216,N_13801,N_13595);
or U14217 (N_14217,N_13558,N_13511);
nor U14218 (N_14218,N_13768,N_13875);
xnor U14219 (N_14219,N_13824,N_13786);
and U14220 (N_14220,N_13992,N_13882);
and U14221 (N_14221,N_13964,N_13907);
and U14222 (N_14222,N_13704,N_13970);
nand U14223 (N_14223,N_13770,N_13532);
xor U14224 (N_14224,N_13604,N_13713);
and U14225 (N_14225,N_13927,N_13864);
and U14226 (N_14226,N_13504,N_13948);
nand U14227 (N_14227,N_13590,N_13790);
and U14228 (N_14228,N_13683,N_13668);
nor U14229 (N_14229,N_13614,N_13968);
and U14230 (N_14230,N_13638,N_13833);
and U14231 (N_14231,N_13644,N_13692);
and U14232 (N_14232,N_13706,N_13568);
and U14233 (N_14233,N_13944,N_13806);
and U14234 (N_14234,N_13751,N_13589);
nand U14235 (N_14235,N_13940,N_13831);
xor U14236 (N_14236,N_13846,N_13756);
nor U14237 (N_14237,N_13555,N_13825);
nand U14238 (N_14238,N_13529,N_13895);
and U14239 (N_14239,N_13536,N_13569);
or U14240 (N_14240,N_13817,N_13890);
nand U14241 (N_14241,N_13549,N_13923);
nand U14242 (N_14242,N_13674,N_13931);
or U14243 (N_14243,N_13962,N_13813);
nor U14244 (N_14244,N_13793,N_13613);
nand U14245 (N_14245,N_13926,N_13872);
nor U14246 (N_14246,N_13514,N_13649);
nand U14247 (N_14247,N_13678,N_13816);
xnor U14248 (N_14248,N_13592,N_13934);
nand U14249 (N_14249,N_13998,N_13689);
xnor U14250 (N_14250,N_13999,N_13786);
nand U14251 (N_14251,N_13825,N_13519);
nand U14252 (N_14252,N_13955,N_13835);
or U14253 (N_14253,N_13891,N_13894);
nand U14254 (N_14254,N_13577,N_13869);
nor U14255 (N_14255,N_13979,N_13902);
nor U14256 (N_14256,N_13831,N_13734);
or U14257 (N_14257,N_13871,N_13922);
nand U14258 (N_14258,N_13669,N_13964);
or U14259 (N_14259,N_13577,N_13928);
or U14260 (N_14260,N_13681,N_13777);
and U14261 (N_14261,N_13784,N_13673);
nor U14262 (N_14262,N_13888,N_13941);
nor U14263 (N_14263,N_13871,N_13623);
or U14264 (N_14264,N_13760,N_13871);
and U14265 (N_14265,N_13956,N_13753);
nand U14266 (N_14266,N_13979,N_13623);
nand U14267 (N_14267,N_13544,N_13647);
nand U14268 (N_14268,N_13951,N_13564);
nor U14269 (N_14269,N_13625,N_13834);
or U14270 (N_14270,N_13611,N_13985);
nand U14271 (N_14271,N_13999,N_13808);
or U14272 (N_14272,N_13617,N_13868);
and U14273 (N_14273,N_13576,N_13783);
or U14274 (N_14274,N_13690,N_13883);
nor U14275 (N_14275,N_13846,N_13778);
xnor U14276 (N_14276,N_13638,N_13964);
and U14277 (N_14277,N_13829,N_13739);
and U14278 (N_14278,N_13685,N_13543);
and U14279 (N_14279,N_13903,N_13734);
or U14280 (N_14280,N_13841,N_13866);
and U14281 (N_14281,N_13579,N_13976);
nor U14282 (N_14282,N_13505,N_13910);
or U14283 (N_14283,N_13793,N_13998);
and U14284 (N_14284,N_13987,N_13745);
nor U14285 (N_14285,N_13520,N_13884);
and U14286 (N_14286,N_13670,N_13843);
nor U14287 (N_14287,N_13926,N_13644);
nand U14288 (N_14288,N_13890,N_13765);
nand U14289 (N_14289,N_13668,N_13755);
or U14290 (N_14290,N_13824,N_13850);
and U14291 (N_14291,N_13654,N_13717);
nand U14292 (N_14292,N_13830,N_13771);
and U14293 (N_14293,N_13970,N_13819);
and U14294 (N_14294,N_13511,N_13909);
or U14295 (N_14295,N_13691,N_13611);
or U14296 (N_14296,N_13613,N_13566);
and U14297 (N_14297,N_13607,N_13676);
and U14298 (N_14298,N_13724,N_13720);
and U14299 (N_14299,N_13786,N_13862);
nand U14300 (N_14300,N_13872,N_13695);
nand U14301 (N_14301,N_13666,N_13716);
and U14302 (N_14302,N_13514,N_13524);
or U14303 (N_14303,N_13745,N_13897);
or U14304 (N_14304,N_13908,N_13801);
nand U14305 (N_14305,N_13852,N_13736);
or U14306 (N_14306,N_13812,N_13931);
nand U14307 (N_14307,N_13578,N_13791);
and U14308 (N_14308,N_13891,N_13806);
nor U14309 (N_14309,N_13544,N_13989);
and U14310 (N_14310,N_13967,N_13938);
and U14311 (N_14311,N_13513,N_13594);
and U14312 (N_14312,N_13872,N_13884);
nand U14313 (N_14313,N_13845,N_13694);
nor U14314 (N_14314,N_13931,N_13547);
nor U14315 (N_14315,N_13537,N_13644);
nand U14316 (N_14316,N_13769,N_13962);
and U14317 (N_14317,N_13797,N_13948);
or U14318 (N_14318,N_13600,N_13934);
nor U14319 (N_14319,N_13988,N_13727);
and U14320 (N_14320,N_13802,N_13534);
and U14321 (N_14321,N_13800,N_13690);
nor U14322 (N_14322,N_13535,N_13764);
or U14323 (N_14323,N_13875,N_13705);
and U14324 (N_14324,N_13783,N_13501);
and U14325 (N_14325,N_13715,N_13629);
and U14326 (N_14326,N_13676,N_13887);
and U14327 (N_14327,N_13638,N_13690);
or U14328 (N_14328,N_13695,N_13793);
xnor U14329 (N_14329,N_13705,N_13793);
and U14330 (N_14330,N_13620,N_13562);
and U14331 (N_14331,N_13907,N_13502);
and U14332 (N_14332,N_13895,N_13531);
or U14333 (N_14333,N_13818,N_13822);
xnor U14334 (N_14334,N_13716,N_13628);
or U14335 (N_14335,N_13697,N_13779);
or U14336 (N_14336,N_13975,N_13772);
nor U14337 (N_14337,N_13634,N_13902);
xor U14338 (N_14338,N_13992,N_13597);
or U14339 (N_14339,N_13801,N_13927);
or U14340 (N_14340,N_13745,N_13539);
nand U14341 (N_14341,N_13829,N_13958);
nor U14342 (N_14342,N_13763,N_13798);
nand U14343 (N_14343,N_13894,N_13913);
and U14344 (N_14344,N_13962,N_13704);
and U14345 (N_14345,N_13835,N_13547);
nand U14346 (N_14346,N_13801,N_13542);
nand U14347 (N_14347,N_13607,N_13530);
and U14348 (N_14348,N_13505,N_13980);
nand U14349 (N_14349,N_13574,N_13583);
and U14350 (N_14350,N_13812,N_13759);
nand U14351 (N_14351,N_13784,N_13781);
and U14352 (N_14352,N_13993,N_13810);
nor U14353 (N_14353,N_13662,N_13751);
and U14354 (N_14354,N_13996,N_13574);
nand U14355 (N_14355,N_13557,N_13569);
nor U14356 (N_14356,N_13811,N_13686);
xor U14357 (N_14357,N_13550,N_13693);
xnor U14358 (N_14358,N_13905,N_13769);
nand U14359 (N_14359,N_13755,N_13733);
nand U14360 (N_14360,N_13626,N_13837);
and U14361 (N_14361,N_13609,N_13551);
nand U14362 (N_14362,N_13584,N_13513);
nand U14363 (N_14363,N_13772,N_13940);
or U14364 (N_14364,N_13560,N_13635);
nor U14365 (N_14365,N_13913,N_13869);
or U14366 (N_14366,N_13989,N_13597);
and U14367 (N_14367,N_13804,N_13889);
nand U14368 (N_14368,N_13788,N_13630);
nor U14369 (N_14369,N_13936,N_13588);
nor U14370 (N_14370,N_13835,N_13994);
and U14371 (N_14371,N_13553,N_13734);
nand U14372 (N_14372,N_13766,N_13655);
nor U14373 (N_14373,N_13787,N_13786);
xor U14374 (N_14374,N_13991,N_13511);
nand U14375 (N_14375,N_13626,N_13542);
or U14376 (N_14376,N_13728,N_13554);
and U14377 (N_14377,N_13697,N_13682);
nor U14378 (N_14378,N_13710,N_13507);
nand U14379 (N_14379,N_13996,N_13624);
or U14380 (N_14380,N_13881,N_13814);
nor U14381 (N_14381,N_13800,N_13894);
nor U14382 (N_14382,N_13599,N_13569);
or U14383 (N_14383,N_13651,N_13954);
or U14384 (N_14384,N_13590,N_13874);
nand U14385 (N_14385,N_13538,N_13947);
nand U14386 (N_14386,N_13748,N_13575);
and U14387 (N_14387,N_13960,N_13918);
and U14388 (N_14388,N_13807,N_13665);
nand U14389 (N_14389,N_13866,N_13976);
nand U14390 (N_14390,N_13566,N_13869);
and U14391 (N_14391,N_13731,N_13632);
nor U14392 (N_14392,N_13939,N_13652);
and U14393 (N_14393,N_13995,N_13767);
and U14394 (N_14394,N_13754,N_13780);
nand U14395 (N_14395,N_13672,N_13846);
xor U14396 (N_14396,N_13920,N_13961);
nand U14397 (N_14397,N_13998,N_13564);
nand U14398 (N_14398,N_13741,N_13855);
nand U14399 (N_14399,N_13753,N_13998);
or U14400 (N_14400,N_13734,N_13866);
and U14401 (N_14401,N_13875,N_13709);
xnor U14402 (N_14402,N_13588,N_13810);
and U14403 (N_14403,N_13536,N_13732);
nor U14404 (N_14404,N_13973,N_13566);
or U14405 (N_14405,N_13613,N_13583);
or U14406 (N_14406,N_13623,N_13854);
and U14407 (N_14407,N_13759,N_13740);
nor U14408 (N_14408,N_13883,N_13936);
and U14409 (N_14409,N_13701,N_13710);
and U14410 (N_14410,N_13655,N_13583);
nand U14411 (N_14411,N_13742,N_13866);
nor U14412 (N_14412,N_13668,N_13770);
nand U14413 (N_14413,N_13846,N_13751);
nor U14414 (N_14414,N_13569,N_13830);
nor U14415 (N_14415,N_13970,N_13604);
and U14416 (N_14416,N_13666,N_13834);
nand U14417 (N_14417,N_13540,N_13814);
and U14418 (N_14418,N_13605,N_13749);
and U14419 (N_14419,N_13743,N_13888);
or U14420 (N_14420,N_13549,N_13658);
nand U14421 (N_14421,N_13590,N_13842);
nor U14422 (N_14422,N_13551,N_13534);
and U14423 (N_14423,N_13857,N_13884);
nand U14424 (N_14424,N_13687,N_13722);
and U14425 (N_14425,N_13773,N_13930);
or U14426 (N_14426,N_13905,N_13848);
or U14427 (N_14427,N_13769,N_13617);
nand U14428 (N_14428,N_13982,N_13612);
nor U14429 (N_14429,N_13710,N_13846);
or U14430 (N_14430,N_13596,N_13865);
or U14431 (N_14431,N_13867,N_13823);
nand U14432 (N_14432,N_13560,N_13527);
and U14433 (N_14433,N_13706,N_13621);
nand U14434 (N_14434,N_13536,N_13561);
or U14435 (N_14435,N_13645,N_13762);
and U14436 (N_14436,N_13793,N_13694);
nand U14437 (N_14437,N_13811,N_13627);
and U14438 (N_14438,N_13739,N_13776);
nor U14439 (N_14439,N_13844,N_13880);
nor U14440 (N_14440,N_13999,N_13807);
and U14441 (N_14441,N_13880,N_13736);
nand U14442 (N_14442,N_13845,N_13896);
nand U14443 (N_14443,N_13706,N_13926);
nor U14444 (N_14444,N_13636,N_13577);
nand U14445 (N_14445,N_13634,N_13535);
xnor U14446 (N_14446,N_13992,N_13588);
nor U14447 (N_14447,N_13614,N_13989);
and U14448 (N_14448,N_13979,N_13554);
and U14449 (N_14449,N_13839,N_13854);
nor U14450 (N_14450,N_13890,N_13528);
and U14451 (N_14451,N_13795,N_13585);
nand U14452 (N_14452,N_13869,N_13833);
or U14453 (N_14453,N_13534,N_13811);
nor U14454 (N_14454,N_13610,N_13602);
nand U14455 (N_14455,N_13645,N_13736);
nand U14456 (N_14456,N_13803,N_13644);
and U14457 (N_14457,N_13654,N_13821);
or U14458 (N_14458,N_13635,N_13985);
or U14459 (N_14459,N_13637,N_13732);
nor U14460 (N_14460,N_13972,N_13876);
nor U14461 (N_14461,N_13617,N_13584);
or U14462 (N_14462,N_13569,N_13682);
and U14463 (N_14463,N_13974,N_13555);
and U14464 (N_14464,N_13650,N_13614);
nor U14465 (N_14465,N_13527,N_13706);
or U14466 (N_14466,N_13705,N_13686);
and U14467 (N_14467,N_13858,N_13862);
xor U14468 (N_14468,N_13529,N_13620);
nor U14469 (N_14469,N_13737,N_13922);
or U14470 (N_14470,N_13570,N_13930);
or U14471 (N_14471,N_13771,N_13666);
nor U14472 (N_14472,N_13812,N_13599);
nor U14473 (N_14473,N_13673,N_13813);
nand U14474 (N_14474,N_13906,N_13886);
nand U14475 (N_14475,N_13800,N_13955);
nor U14476 (N_14476,N_13615,N_13708);
nand U14477 (N_14477,N_13632,N_13643);
nor U14478 (N_14478,N_13824,N_13895);
nand U14479 (N_14479,N_13685,N_13601);
nand U14480 (N_14480,N_13567,N_13551);
nor U14481 (N_14481,N_13654,N_13785);
and U14482 (N_14482,N_13677,N_13969);
xor U14483 (N_14483,N_13777,N_13665);
nand U14484 (N_14484,N_13972,N_13667);
or U14485 (N_14485,N_13875,N_13720);
nand U14486 (N_14486,N_13527,N_13984);
nor U14487 (N_14487,N_13871,N_13666);
xnor U14488 (N_14488,N_13832,N_13506);
or U14489 (N_14489,N_13595,N_13808);
or U14490 (N_14490,N_13611,N_13550);
or U14491 (N_14491,N_13514,N_13549);
nor U14492 (N_14492,N_13587,N_13855);
or U14493 (N_14493,N_13871,N_13966);
nor U14494 (N_14494,N_13578,N_13715);
and U14495 (N_14495,N_13752,N_13877);
or U14496 (N_14496,N_13983,N_13997);
nor U14497 (N_14497,N_13734,N_13912);
or U14498 (N_14498,N_13574,N_13984);
or U14499 (N_14499,N_13652,N_13766);
xor U14500 (N_14500,N_14324,N_14456);
and U14501 (N_14501,N_14053,N_14159);
nand U14502 (N_14502,N_14007,N_14113);
and U14503 (N_14503,N_14181,N_14412);
and U14504 (N_14504,N_14028,N_14069);
and U14505 (N_14505,N_14365,N_14085);
nand U14506 (N_14506,N_14256,N_14380);
xnor U14507 (N_14507,N_14010,N_14091);
or U14508 (N_14508,N_14375,N_14071);
nor U14509 (N_14509,N_14156,N_14134);
nand U14510 (N_14510,N_14383,N_14038);
or U14511 (N_14511,N_14100,N_14180);
xor U14512 (N_14512,N_14428,N_14036);
or U14513 (N_14513,N_14473,N_14055);
and U14514 (N_14514,N_14026,N_14361);
or U14515 (N_14515,N_14228,N_14090);
or U14516 (N_14516,N_14114,N_14004);
nor U14517 (N_14517,N_14030,N_14407);
nand U14518 (N_14518,N_14045,N_14013);
or U14519 (N_14519,N_14147,N_14079);
nor U14520 (N_14520,N_14182,N_14430);
nand U14521 (N_14521,N_14040,N_14077);
nor U14522 (N_14522,N_14342,N_14291);
nor U14523 (N_14523,N_14024,N_14219);
and U14524 (N_14524,N_14230,N_14042);
and U14525 (N_14525,N_14101,N_14122);
nand U14526 (N_14526,N_14203,N_14389);
and U14527 (N_14527,N_14396,N_14478);
or U14528 (N_14528,N_14002,N_14021);
nand U14529 (N_14529,N_14083,N_14102);
nor U14530 (N_14530,N_14277,N_14311);
nand U14531 (N_14531,N_14381,N_14175);
and U14532 (N_14532,N_14312,N_14041);
or U14533 (N_14533,N_14443,N_14033);
nand U14534 (N_14534,N_14067,N_14323);
nor U14535 (N_14535,N_14484,N_14206);
xnor U14536 (N_14536,N_14223,N_14339);
nand U14537 (N_14537,N_14094,N_14264);
and U14538 (N_14538,N_14016,N_14255);
or U14539 (N_14539,N_14297,N_14358);
or U14540 (N_14540,N_14355,N_14370);
nor U14541 (N_14541,N_14179,N_14224);
nand U14542 (N_14542,N_14326,N_14427);
nor U14543 (N_14543,N_14418,N_14419);
nor U14544 (N_14544,N_14399,N_14497);
nand U14545 (N_14545,N_14317,N_14299);
or U14546 (N_14546,N_14458,N_14334);
and U14547 (N_14547,N_14359,N_14210);
nor U14548 (N_14548,N_14406,N_14214);
nor U14549 (N_14549,N_14075,N_14272);
nor U14550 (N_14550,N_14072,N_14105);
nand U14551 (N_14551,N_14405,N_14236);
or U14552 (N_14552,N_14336,N_14189);
and U14553 (N_14553,N_14322,N_14377);
nor U14554 (N_14554,N_14486,N_14271);
nor U14555 (N_14555,N_14483,N_14188);
nor U14556 (N_14556,N_14138,N_14480);
and U14557 (N_14557,N_14276,N_14052);
nand U14558 (N_14558,N_14426,N_14371);
and U14559 (N_14559,N_14227,N_14054);
or U14560 (N_14560,N_14201,N_14131);
xnor U14561 (N_14561,N_14125,N_14158);
nor U14562 (N_14562,N_14410,N_14195);
nand U14563 (N_14563,N_14460,N_14435);
nor U14564 (N_14564,N_14066,N_14328);
or U14565 (N_14565,N_14337,N_14310);
or U14566 (N_14566,N_14115,N_14395);
nor U14567 (N_14567,N_14049,N_14393);
xor U14568 (N_14568,N_14459,N_14363);
xor U14569 (N_14569,N_14307,N_14120);
nand U14570 (N_14570,N_14382,N_14379);
and U14571 (N_14571,N_14374,N_14281);
or U14572 (N_14572,N_14470,N_14218);
nor U14573 (N_14573,N_14314,N_14464);
and U14574 (N_14574,N_14466,N_14409);
xnor U14575 (N_14575,N_14130,N_14221);
xor U14576 (N_14576,N_14293,N_14047);
nor U14577 (N_14577,N_14136,N_14129);
and U14578 (N_14578,N_14239,N_14216);
nand U14579 (N_14579,N_14110,N_14099);
xor U14580 (N_14580,N_14319,N_14025);
nor U14581 (N_14581,N_14039,N_14414);
or U14582 (N_14582,N_14487,N_14243);
nor U14583 (N_14583,N_14284,N_14309);
nor U14584 (N_14584,N_14289,N_14126);
or U14585 (N_14585,N_14288,N_14367);
xor U14586 (N_14586,N_14017,N_14244);
xor U14587 (N_14587,N_14020,N_14296);
and U14588 (N_14588,N_14167,N_14265);
or U14589 (N_14589,N_14076,N_14242);
nor U14590 (N_14590,N_14263,N_14401);
and U14591 (N_14591,N_14354,N_14205);
nor U14592 (N_14592,N_14262,N_14402);
nor U14593 (N_14593,N_14250,N_14420);
nor U14594 (N_14594,N_14306,N_14422);
nor U14595 (N_14595,N_14012,N_14270);
or U14596 (N_14596,N_14434,N_14006);
and U14597 (N_14597,N_14109,N_14280);
nand U14598 (N_14598,N_14346,N_14215);
or U14599 (N_14599,N_14366,N_14490);
nand U14600 (N_14600,N_14461,N_14124);
nor U14601 (N_14601,N_14032,N_14043);
nand U14602 (N_14602,N_14169,N_14184);
nand U14603 (N_14603,N_14226,N_14247);
nand U14604 (N_14604,N_14074,N_14260);
xnor U14605 (N_14605,N_14092,N_14436);
nand U14606 (N_14606,N_14217,N_14425);
or U14607 (N_14607,N_14325,N_14408);
nand U14608 (N_14608,N_14469,N_14404);
and U14609 (N_14609,N_14485,N_14259);
or U14610 (N_14610,N_14440,N_14015);
or U14611 (N_14611,N_14064,N_14438);
nand U14612 (N_14612,N_14249,N_14157);
or U14613 (N_14613,N_14001,N_14295);
nand U14614 (N_14614,N_14357,N_14029);
or U14615 (N_14615,N_14369,N_14397);
nand U14616 (N_14616,N_14160,N_14424);
nand U14617 (N_14617,N_14137,N_14154);
nand U14618 (N_14618,N_14344,N_14390);
nor U14619 (N_14619,N_14373,N_14240);
and U14620 (N_14620,N_14011,N_14372);
and U14621 (N_14621,N_14423,N_14060);
nor U14622 (N_14622,N_14398,N_14246);
and U14623 (N_14623,N_14388,N_14467);
or U14624 (N_14624,N_14446,N_14096);
or U14625 (N_14625,N_14097,N_14302);
nor U14626 (N_14626,N_14448,N_14368);
nor U14627 (N_14627,N_14168,N_14479);
nand U14628 (N_14628,N_14347,N_14022);
nor U14629 (N_14629,N_14107,N_14148);
or U14630 (N_14630,N_14348,N_14237);
nor U14631 (N_14631,N_14447,N_14305);
and U14632 (N_14632,N_14378,N_14135);
nor U14633 (N_14633,N_14451,N_14048);
nand U14634 (N_14634,N_14274,N_14472);
nand U14635 (N_14635,N_14104,N_14251);
xor U14636 (N_14636,N_14127,N_14482);
or U14637 (N_14637,N_14498,N_14174);
or U14638 (N_14638,N_14194,N_14353);
and U14639 (N_14639,N_14121,N_14000);
and U14640 (N_14640,N_14035,N_14449);
xor U14641 (N_14641,N_14123,N_14233);
nand U14642 (N_14642,N_14304,N_14057);
and U14643 (N_14643,N_14084,N_14463);
and U14644 (N_14644,N_14394,N_14014);
nand U14645 (N_14645,N_14192,N_14253);
and U14646 (N_14646,N_14294,N_14351);
nor U14647 (N_14647,N_14177,N_14093);
or U14648 (N_14648,N_14481,N_14112);
or U14649 (N_14649,N_14301,N_14139);
nor U14650 (N_14650,N_14141,N_14178);
nor U14651 (N_14651,N_14350,N_14080);
or U14652 (N_14652,N_14300,N_14362);
or U14653 (N_14653,N_14421,N_14111);
and U14654 (N_14654,N_14453,N_14051);
and U14655 (N_14655,N_14145,N_14252);
or U14656 (N_14656,N_14208,N_14257);
nor U14657 (N_14657,N_14128,N_14429);
and U14658 (N_14658,N_14432,N_14162);
nor U14659 (N_14659,N_14003,N_14279);
nor U14660 (N_14660,N_14116,N_14212);
nand U14661 (N_14661,N_14386,N_14161);
and U14662 (N_14662,N_14176,N_14197);
xnor U14663 (N_14663,N_14153,N_14061);
or U14664 (N_14664,N_14496,N_14118);
or U14665 (N_14665,N_14384,N_14411);
and U14666 (N_14666,N_14171,N_14320);
nor U14667 (N_14667,N_14341,N_14313);
and U14668 (N_14668,N_14005,N_14098);
nor U14669 (N_14669,N_14499,N_14046);
nor U14670 (N_14670,N_14088,N_14462);
and U14671 (N_14671,N_14415,N_14119);
nand U14672 (N_14672,N_14292,N_14059);
xor U14673 (N_14673,N_14019,N_14209);
or U14674 (N_14674,N_14267,N_14170);
nor U14675 (N_14675,N_14431,N_14298);
or U14676 (N_14676,N_14282,N_14465);
and U14677 (N_14677,N_14173,N_14211);
nand U14678 (N_14678,N_14106,N_14152);
or U14679 (N_14679,N_14391,N_14331);
or U14680 (N_14680,N_14273,N_14155);
and U14681 (N_14681,N_14027,N_14023);
or U14682 (N_14682,N_14491,N_14338);
xor U14683 (N_14683,N_14349,N_14143);
nand U14684 (N_14684,N_14073,N_14050);
nor U14685 (N_14685,N_14471,N_14327);
and U14686 (N_14686,N_14321,N_14196);
nor U14687 (N_14687,N_14009,N_14031);
nor U14688 (N_14688,N_14417,N_14268);
or U14689 (N_14689,N_14364,N_14231);
nand U14690 (N_14690,N_14018,N_14454);
nor U14691 (N_14691,N_14193,N_14492);
or U14692 (N_14692,N_14034,N_14087);
and U14693 (N_14693,N_14238,N_14133);
or U14694 (N_14694,N_14254,N_14444);
and U14695 (N_14695,N_14163,N_14235);
nand U14696 (N_14696,N_14477,N_14150);
nand U14697 (N_14697,N_14278,N_14433);
xor U14698 (N_14698,N_14285,N_14283);
or U14699 (N_14699,N_14222,N_14489);
or U14700 (N_14700,N_14086,N_14199);
nor U14701 (N_14701,N_14202,N_14149);
nor U14702 (N_14702,N_14345,N_14225);
nor U14703 (N_14703,N_14008,N_14070);
or U14704 (N_14704,N_14318,N_14387);
or U14705 (N_14705,N_14385,N_14213);
and U14706 (N_14706,N_14081,N_14476);
xnor U14707 (N_14707,N_14204,N_14303);
and U14708 (N_14708,N_14333,N_14455);
and U14709 (N_14709,N_14117,N_14146);
or U14710 (N_14710,N_14063,N_14078);
nor U14711 (N_14711,N_14095,N_14494);
nor U14712 (N_14712,N_14330,N_14457);
nand U14713 (N_14713,N_14488,N_14186);
nand U14714 (N_14714,N_14392,N_14441);
and U14715 (N_14715,N_14132,N_14413);
or U14716 (N_14716,N_14315,N_14360);
nor U14717 (N_14717,N_14445,N_14335);
or U14718 (N_14718,N_14082,N_14232);
or U14719 (N_14719,N_14140,N_14185);
nor U14720 (N_14720,N_14248,N_14452);
nor U14721 (N_14721,N_14329,N_14450);
and U14722 (N_14722,N_14229,N_14286);
nor U14723 (N_14723,N_14142,N_14172);
nor U14724 (N_14724,N_14183,N_14495);
nand U14725 (N_14725,N_14068,N_14220);
and U14726 (N_14726,N_14261,N_14044);
or U14727 (N_14727,N_14356,N_14062);
nand U14728 (N_14728,N_14191,N_14151);
xor U14729 (N_14729,N_14475,N_14065);
nor U14730 (N_14730,N_14058,N_14165);
or U14731 (N_14731,N_14089,N_14103);
nor U14732 (N_14732,N_14287,N_14439);
and U14733 (N_14733,N_14245,N_14198);
xor U14734 (N_14734,N_14108,N_14144);
or U14735 (N_14735,N_14234,N_14190);
nor U14736 (N_14736,N_14207,N_14416);
nor U14737 (N_14737,N_14468,N_14266);
or U14738 (N_14738,N_14437,N_14056);
and U14739 (N_14739,N_14187,N_14308);
nor U14740 (N_14740,N_14376,N_14316);
nor U14741 (N_14741,N_14037,N_14400);
nor U14742 (N_14742,N_14352,N_14343);
nand U14743 (N_14743,N_14290,N_14493);
and U14744 (N_14744,N_14332,N_14275);
xnor U14745 (N_14745,N_14474,N_14166);
or U14746 (N_14746,N_14442,N_14258);
xnor U14747 (N_14747,N_14269,N_14340);
nor U14748 (N_14748,N_14200,N_14241);
xnor U14749 (N_14749,N_14164,N_14403);
nand U14750 (N_14750,N_14463,N_14136);
or U14751 (N_14751,N_14335,N_14145);
and U14752 (N_14752,N_14313,N_14076);
or U14753 (N_14753,N_14406,N_14164);
nor U14754 (N_14754,N_14423,N_14259);
nand U14755 (N_14755,N_14045,N_14390);
or U14756 (N_14756,N_14082,N_14098);
or U14757 (N_14757,N_14141,N_14003);
or U14758 (N_14758,N_14225,N_14057);
or U14759 (N_14759,N_14043,N_14192);
and U14760 (N_14760,N_14350,N_14115);
or U14761 (N_14761,N_14040,N_14125);
nor U14762 (N_14762,N_14339,N_14490);
xnor U14763 (N_14763,N_14341,N_14366);
and U14764 (N_14764,N_14085,N_14302);
nor U14765 (N_14765,N_14364,N_14290);
and U14766 (N_14766,N_14134,N_14120);
and U14767 (N_14767,N_14279,N_14146);
and U14768 (N_14768,N_14301,N_14417);
nor U14769 (N_14769,N_14315,N_14111);
xnor U14770 (N_14770,N_14247,N_14050);
xnor U14771 (N_14771,N_14113,N_14191);
and U14772 (N_14772,N_14108,N_14281);
nand U14773 (N_14773,N_14184,N_14241);
nor U14774 (N_14774,N_14155,N_14027);
xnor U14775 (N_14775,N_14081,N_14264);
xor U14776 (N_14776,N_14241,N_14350);
nor U14777 (N_14777,N_14445,N_14147);
nor U14778 (N_14778,N_14161,N_14478);
or U14779 (N_14779,N_14456,N_14163);
or U14780 (N_14780,N_14221,N_14036);
and U14781 (N_14781,N_14065,N_14153);
nand U14782 (N_14782,N_14007,N_14374);
nor U14783 (N_14783,N_14280,N_14441);
nand U14784 (N_14784,N_14189,N_14402);
nand U14785 (N_14785,N_14276,N_14195);
and U14786 (N_14786,N_14274,N_14054);
and U14787 (N_14787,N_14018,N_14451);
xnor U14788 (N_14788,N_14076,N_14410);
or U14789 (N_14789,N_14363,N_14233);
or U14790 (N_14790,N_14103,N_14334);
and U14791 (N_14791,N_14412,N_14423);
nand U14792 (N_14792,N_14447,N_14088);
and U14793 (N_14793,N_14381,N_14347);
xnor U14794 (N_14794,N_14256,N_14228);
and U14795 (N_14795,N_14428,N_14411);
or U14796 (N_14796,N_14231,N_14400);
nor U14797 (N_14797,N_14347,N_14269);
and U14798 (N_14798,N_14414,N_14051);
nand U14799 (N_14799,N_14480,N_14321);
nor U14800 (N_14800,N_14340,N_14376);
or U14801 (N_14801,N_14343,N_14176);
or U14802 (N_14802,N_14455,N_14488);
nor U14803 (N_14803,N_14143,N_14042);
nor U14804 (N_14804,N_14159,N_14067);
or U14805 (N_14805,N_14019,N_14135);
nor U14806 (N_14806,N_14047,N_14433);
or U14807 (N_14807,N_14431,N_14474);
nand U14808 (N_14808,N_14482,N_14349);
xnor U14809 (N_14809,N_14235,N_14178);
and U14810 (N_14810,N_14149,N_14427);
and U14811 (N_14811,N_14013,N_14231);
and U14812 (N_14812,N_14433,N_14245);
nand U14813 (N_14813,N_14267,N_14462);
nand U14814 (N_14814,N_14385,N_14246);
and U14815 (N_14815,N_14342,N_14013);
nor U14816 (N_14816,N_14332,N_14183);
nand U14817 (N_14817,N_14326,N_14478);
nor U14818 (N_14818,N_14108,N_14255);
xnor U14819 (N_14819,N_14408,N_14059);
xnor U14820 (N_14820,N_14370,N_14120);
nand U14821 (N_14821,N_14057,N_14187);
nand U14822 (N_14822,N_14414,N_14381);
nor U14823 (N_14823,N_14289,N_14190);
or U14824 (N_14824,N_14429,N_14444);
nor U14825 (N_14825,N_14109,N_14077);
or U14826 (N_14826,N_14215,N_14243);
nand U14827 (N_14827,N_14401,N_14074);
xor U14828 (N_14828,N_14078,N_14333);
nand U14829 (N_14829,N_14034,N_14082);
nor U14830 (N_14830,N_14327,N_14448);
nor U14831 (N_14831,N_14317,N_14050);
or U14832 (N_14832,N_14112,N_14020);
and U14833 (N_14833,N_14135,N_14025);
or U14834 (N_14834,N_14304,N_14229);
nor U14835 (N_14835,N_14259,N_14130);
nand U14836 (N_14836,N_14235,N_14285);
or U14837 (N_14837,N_14491,N_14274);
nor U14838 (N_14838,N_14349,N_14492);
nand U14839 (N_14839,N_14232,N_14285);
or U14840 (N_14840,N_14289,N_14259);
nor U14841 (N_14841,N_14430,N_14260);
and U14842 (N_14842,N_14192,N_14207);
nand U14843 (N_14843,N_14141,N_14102);
nand U14844 (N_14844,N_14010,N_14353);
and U14845 (N_14845,N_14134,N_14355);
nand U14846 (N_14846,N_14274,N_14248);
xor U14847 (N_14847,N_14026,N_14252);
and U14848 (N_14848,N_14164,N_14440);
nand U14849 (N_14849,N_14413,N_14118);
nand U14850 (N_14850,N_14339,N_14318);
or U14851 (N_14851,N_14273,N_14383);
and U14852 (N_14852,N_14237,N_14327);
or U14853 (N_14853,N_14242,N_14081);
nand U14854 (N_14854,N_14460,N_14020);
and U14855 (N_14855,N_14189,N_14292);
nand U14856 (N_14856,N_14348,N_14235);
or U14857 (N_14857,N_14097,N_14060);
or U14858 (N_14858,N_14152,N_14155);
nor U14859 (N_14859,N_14136,N_14439);
nor U14860 (N_14860,N_14310,N_14274);
or U14861 (N_14861,N_14010,N_14005);
nand U14862 (N_14862,N_14139,N_14211);
and U14863 (N_14863,N_14221,N_14473);
or U14864 (N_14864,N_14028,N_14181);
nor U14865 (N_14865,N_14186,N_14007);
and U14866 (N_14866,N_14437,N_14257);
or U14867 (N_14867,N_14051,N_14446);
nor U14868 (N_14868,N_14028,N_14021);
or U14869 (N_14869,N_14045,N_14295);
or U14870 (N_14870,N_14122,N_14007);
or U14871 (N_14871,N_14004,N_14182);
nand U14872 (N_14872,N_14086,N_14357);
or U14873 (N_14873,N_14153,N_14072);
nor U14874 (N_14874,N_14215,N_14087);
or U14875 (N_14875,N_14337,N_14075);
nand U14876 (N_14876,N_14274,N_14449);
nor U14877 (N_14877,N_14154,N_14050);
or U14878 (N_14878,N_14146,N_14349);
nand U14879 (N_14879,N_14411,N_14459);
and U14880 (N_14880,N_14072,N_14467);
or U14881 (N_14881,N_14182,N_14402);
nor U14882 (N_14882,N_14056,N_14480);
or U14883 (N_14883,N_14057,N_14002);
nor U14884 (N_14884,N_14147,N_14464);
and U14885 (N_14885,N_14032,N_14175);
nor U14886 (N_14886,N_14239,N_14159);
and U14887 (N_14887,N_14419,N_14431);
nor U14888 (N_14888,N_14203,N_14245);
nor U14889 (N_14889,N_14115,N_14211);
nand U14890 (N_14890,N_14494,N_14064);
or U14891 (N_14891,N_14229,N_14363);
nand U14892 (N_14892,N_14000,N_14306);
nor U14893 (N_14893,N_14080,N_14273);
and U14894 (N_14894,N_14317,N_14297);
or U14895 (N_14895,N_14426,N_14175);
nand U14896 (N_14896,N_14009,N_14029);
or U14897 (N_14897,N_14132,N_14064);
or U14898 (N_14898,N_14461,N_14175);
and U14899 (N_14899,N_14371,N_14004);
and U14900 (N_14900,N_14372,N_14267);
nor U14901 (N_14901,N_14486,N_14019);
nand U14902 (N_14902,N_14472,N_14130);
nor U14903 (N_14903,N_14265,N_14305);
nor U14904 (N_14904,N_14092,N_14075);
nor U14905 (N_14905,N_14017,N_14167);
or U14906 (N_14906,N_14136,N_14327);
or U14907 (N_14907,N_14010,N_14349);
nand U14908 (N_14908,N_14428,N_14027);
xor U14909 (N_14909,N_14178,N_14018);
nand U14910 (N_14910,N_14219,N_14489);
or U14911 (N_14911,N_14136,N_14013);
or U14912 (N_14912,N_14401,N_14170);
and U14913 (N_14913,N_14292,N_14253);
nor U14914 (N_14914,N_14449,N_14073);
xnor U14915 (N_14915,N_14331,N_14288);
nor U14916 (N_14916,N_14038,N_14103);
and U14917 (N_14917,N_14091,N_14235);
and U14918 (N_14918,N_14353,N_14030);
nor U14919 (N_14919,N_14494,N_14497);
and U14920 (N_14920,N_14048,N_14327);
xnor U14921 (N_14921,N_14390,N_14052);
nand U14922 (N_14922,N_14427,N_14094);
xnor U14923 (N_14923,N_14310,N_14497);
or U14924 (N_14924,N_14278,N_14364);
nor U14925 (N_14925,N_14236,N_14477);
and U14926 (N_14926,N_14497,N_14334);
nand U14927 (N_14927,N_14117,N_14086);
nor U14928 (N_14928,N_14262,N_14463);
nand U14929 (N_14929,N_14230,N_14201);
or U14930 (N_14930,N_14371,N_14182);
nor U14931 (N_14931,N_14162,N_14169);
and U14932 (N_14932,N_14354,N_14004);
nand U14933 (N_14933,N_14296,N_14447);
nor U14934 (N_14934,N_14364,N_14256);
nor U14935 (N_14935,N_14384,N_14373);
nand U14936 (N_14936,N_14287,N_14466);
nand U14937 (N_14937,N_14472,N_14267);
nand U14938 (N_14938,N_14114,N_14090);
nand U14939 (N_14939,N_14335,N_14072);
and U14940 (N_14940,N_14263,N_14160);
nor U14941 (N_14941,N_14163,N_14192);
and U14942 (N_14942,N_14383,N_14085);
or U14943 (N_14943,N_14025,N_14480);
and U14944 (N_14944,N_14004,N_14257);
or U14945 (N_14945,N_14469,N_14008);
nor U14946 (N_14946,N_14491,N_14256);
nand U14947 (N_14947,N_14478,N_14015);
nand U14948 (N_14948,N_14125,N_14025);
nand U14949 (N_14949,N_14026,N_14364);
and U14950 (N_14950,N_14437,N_14409);
nor U14951 (N_14951,N_14117,N_14151);
nor U14952 (N_14952,N_14272,N_14145);
nor U14953 (N_14953,N_14239,N_14404);
or U14954 (N_14954,N_14369,N_14211);
or U14955 (N_14955,N_14151,N_14287);
or U14956 (N_14956,N_14467,N_14144);
nand U14957 (N_14957,N_14382,N_14290);
nor U14958 (N_14958,N_14462,N_14474);
nor U14959 (N_14959,N_14127,N_14047);
or U14960 (N_14960,N_14373,N_14274);
nor U14961 (N_14961,N_14120,N_14020);
nand U14962 (N_14962,N_14354,N_14211);
nor U14963 (N_14963,N_14266,N_14380);
and U14964 (N_14964,N_14046,N_14031);
or U14965 (N_14965,N_14174,N_14007);
nand U14966 (N_14966,N_14126,N_14481);
nor U14967 (N_14967,N_14361,N_14263);
nor U14968 (N_14968,N_14208,N_14199);
nor U14969 (N_14969,N_14322,N_14435);
nand U14970 (N_14970,N_14075,N_14135);
and U14971 (N_14971,N_14292,N_14126);
and U14972 (N_14972,N_14252,N_14226);
or U14973 (N_14973,N_14179,N_14057);
nor U14974 (N_14974,N_14219,N_14494);
nand U14975 (N_14975,N_14228,N_14086);
or U14976 (N_14976,N_14306,N_14108);
nor U14977 (N_14977,N_14230,N_14015);
or U14978 (N_14978,N_14238,N_14322);
nor U14979 (N_14979,N_14164,N_14016);
and U14980 (N_14980,N_14156,N_14273);
and U14981 (N_14981,N_14400,N_14386);
or U14982 (N_14982,N_14245,N_14142);
or U14983 (N_14983,N_14459,N_14049);
nor U14984 (N_14984,N_14365,N_14172);
and U14985 (N_14985,N_14088,N_14321);
and U14986 (N_14986,N_14307,N_14025);
nand U14987 (N_14987,N_14011,N_14472);
and U14988 (N_14988,N_14228,N_14394);
xnor U14989 (N_14989,N_14151,N_14391);
nor U14990 (N_14990,N_14184,N_14185);
and U14991 (N_14991,N_14432,N_14139);
nand U14992 (N_14992,N_14241,N_14288);
nand U14993 (N_14993,N_14059,N_14108);
nor U14994 (N_14994,N_14032,N_14161);
xnor U14995 (N_14995,N_14281,N_14117);
nor U14996 (N_14996,N_14388,N_14091);
nand U14997 (N_14997,N_14335,N_14192);
or U14998 (N_14998,N_14486,N_14182);
nor U14999 (N_14999,N_14434,N_14214);
and U15000 (N_15000,N_14609,N_14613);
nand U15001 (N_15001,N_14932,N_14946);
nand U15002 (N_15002,N_14914,N_14598);
xnor U15003 (N_15003,N_14992,N_14817);
xnor U15004 (N_15004,N_14942,N_14680);
and U15005 (N_15005,N_14518,N_14940);
nor U15006 (N_15006,N_14569,N_14705);
and U15007 (N_15007,N_14661,N_14601);
and U15008 (N_15008,N_14894,N_14763);
or U15009 (N_15009,N_14665,N_14531);
nor U15010 (N_15010,N_14624,N_14880);
nor U15011 (N_15011,N_14808,N_14733);
nor U15012 (N_15012,N_14693,N_14989);
or U15013 (N_15013,N_14585,N_14745);
nor U15014 (N_15014,N_14538,N_14660);
nor U15015 (N_15015,N_14892,N_14699);
xnor U15016 (N_15016,N_14893,N_14859);
nand U15017 (N_15017,N_14648,N_14551);
and U15018 (N_15018,N_14750,N_14823);
and U15019 (N_15019,N_14802,N_14522);
and U15020 (N_15020,N_14643,N_14540);
and U15021 (N_15021,N_14861,N_14881);
nor U15022 (N_15022,N_14519,N_14617);
nand U15023 (N_15023,N_14959,N_14637);
or U15024 (N_15024,N_14957,N_14656);
nor U15025 (N_15025,N_14945,N_14712);
nor U15026 (N_15026,N_14931,N_14868);
nor U15027 (N_15027,N_14911,N_14824);
and U15028 (N_15028,N_14528,N_14939);
and U15029 (N_15029,N_14707,N_14595);
nor U15030 (N_15030,N_14998,N_14543);
or U15031 (N_15031,N_14575,N_14625);
and U15032 (N_15032,N_14753,N_14898);
nor U15033 (N_15033,N_14628,N_14944);
nor U15034 (N_15034,N_14830,N_14848);
nand U15035 (N_15035,N_14561,N_14798);
nor U15036 (N_15036,N_14542,N_14662);
and U15037 (N_15037,N_14696,N_14864);
nor U15038 (N_15038,N_14722,N_14935);
nand U15039 (N_15039,N_14618,N_14607);
or U15040 (N_15040,N_14626,N_14726);
nor U15041 (N_15041,N_14502,N_14651);
nor U15042 (N_15042,N_14521,N_14611);
or U15043 (N_15043,N_14579,N_14671);
xor U15044 (N_15044,N_14730,N_14586);
nor U15045 (N_15045,N_14907,N_14622);
or U15046 (N_15046,N_14866,N_14532);
or U15047 (N_15047,N_14619,N_14837);
nor U15048 (N_15048,N_14562,N_14718);
and U15049 (N_15049,N_14938,N_14860);
and U15050 (N_15050,N_14577,N_14644);
xnor U15051 (N_15051,N_14887,N_14820);
or U15052 (N_15052,N_14999,N_14772);
and U15053 (N_15053,N_14779,N_14889);
or U15054 (N_15054,N_14636,N_14714);
and U15055 (N_15055,N_14582,N_14762);
nand U15056 (N_15056,N_14571,N_14875);
nor U15057 (N_15057,N_14507,N_14663);
nand U15058 (N_15058,N_14670,N_14510);
nor U15059 (N_15059,N_14841,N_14814);
or U15060 (N_15060,N_14997,N_14771);
or U15061 (N_15061,N_14879,N_14534);
and U15062 (N_15062,N_14810,N_14621);
or U15063 (N_15063,N_14869,N_14882);
or U15064 (N_15064,N_14839,N_14685);
or U15065 (N_15065,N_14840,N_14857);
xor U15066 (N_15066,N_14947,N_14702);
or U15067 (N_15067,N_14970,N_14846);
nand U15068 (N_15068,N_14512,N_14654);
or U15069 (N_15069,N_14659,N_14977);
or U15070 (N_15070,N_14552,N_14682);
xnor U15071 (N_15071,N_14872,N_14574);
and U15072 (N_15072,N_14549,N_14533);
nand U15073 (N_15073,N_14835,N_14544);
nor U15074 (N_15074,N_14678,N_14852);
and U15075 (N_15075,N_14755,N_14732);
nand U15076 (N_15076,N_14987,N_14933);
and U15077 (N_15077,N_14941,N_14928);
nand U15078 (N_15078,N_14853,N_14728);
or U15079 (N_15079,N_14547,N_14969);
or U15080 (N_15080,N_14587,N_14976);
nand U15081 (N_15081,N_14523,N_14981);
xnor U15082 (N_15082,N_14556,N_14583);
nor U15083 (N_15083,N_14883,N_14650);
nand U15084 (N_15084,N_14641,N_14793);
nand U15085 (N_15085,N_14681,N_14600);
and U15086 (N_15086,N_14723,N_14974);
or U15087 (N_15087,N_14948,N_14535);
nor U15088 (N_15088,N_14821,N_14890);
or U15089 (N_15089,N_14781,N_14708);
or U15090 (N_15090,N_14983,N_14790);
nand U15091 (N_15091,N_14594,N_14546);
nor U15092 (N_15092,N_14843,N_14847);
nor U15093 (N_15093,N_14525,N_14689);
nand U15094 (N_15094,N_14580,N_14871);
and U15095 (N_15095,N_14952,N_14949);
nor U15096 (N_15096,N_14951,N_14891);
nand U15097 (N_15097,N_14508,N_14789);
nand U15098 (N_15098,N_14727,N_14612);
nor U15099 (N_15099,N_14829,N_14706);
nand U15100 (N_15100,N_14740,N_14627);
xor U15101 (N_15101,N_14800,N_14954);
and U15102 (N_15102,N_14501,N_14504);
or U15103 (N_15103,N_14845,N_14873);
and U15104 (N_15104,N_14675,N_14908);
xnor U15105 (N_15105,N_14895,N_14920);
xor U15106 (N_15106,N_14784,N_14704);
nand U15107 (N_15107,N_14623,N_14553);
or U15108 (N_15108,N_14710,N_14596);
xnor U15109 (N_15109,N_14917,N_14764);
or U15110 (N_15110,N_14652,N_14742);
or U15111 (N_15111,N_14673,N_14778);
and U15112 (N_15112,N_14955,N_14934);
or U15113 (N_15113,N_14903,N_14500);
or U15114 (N_15114,N_14801,N_14688);
xnor U15115 (N_15115,N_14536,N_14655);
or U15116 (N_15116,N_14642,N_14565);
and U15117 (N_15117,N_14985,N_14927);
nor U15118 (N_15118,N_14930,N_14776);
nor U15119 (N_15119,N_14990,N_14581);
xor U15120 (N_15120,N_14721,N_14608);
nor U15121 (N_15121,N_14827,N_14912);
and U15122 (N_15122,N_14819,N_14667);
nand U15123 (N_15123,N_14995,N_14876);
or U15124 (N_15124,N_14701,N_14620);
and U15125 (N_15125,N_14862,N_14804);
nand U15126 (N_15126,N_14516,N_14511);
nand U15127 (N_15127,N_14697,N_14795);
xor U15128 (N_15128,N_14765,N_14825);
nand U15129 (N_15129,N_14548,N_14967);
and U15130 (N_15130,N_14588,N_14572);
xor U15131 (N_15131,N_14921,N_14657);
or U15132 (N_15132,N_14834,N_14509);
xor U15133 (N_15133,N_14766,N_14926);
nand U15134 (N_15134,N_14878,N_14807);
or U15135 (N_15135,N_14557,N_14692);
nand U15136 (N_15136,N_14666,N_14629);
or U15137 (N_15137,N_14818,N_14683);
nor U15138 (N_15138,N_14849,N_14719);
and U15139 (N_15139,N_14972,N_14958);
and U15140 (N_15140,N_14592,N_14741);
and U15141 (N_15141,N_14785,N_14568);
or U15142 (N_15142,N_14550,N_14640);
or U15143 (N_15143,N_14811,N_14822);
nor U15144 (N_15144,N_14943,N_14828);
nor U15145 (N_15145,N_14633,N_14515);
and U15146 (N_15146,N_14774,N_14922);
nor U15147 (N_15147,N_14605,N_14555);
and U15148 (N_15148,N_14526,N_14530);
xnor U15149 (N_15149,N_14649,N_14858);
nor U15150 (N_15150,N_14724,N_14694);
nand U15151 (N_15151,N_14744,N_14677);
nand U15152 (N_15152,N_14517,N_14996);
xnor U15153 (N_15153,N_14988,N_14760);
nand U15154 (N_15154,N_14832,N_14713);
and U15155 (N_15155,N_14506,N_14539);
xnor U15156 (N_15156,N_14794,N_14953);
nand U15157 (N_15157,N_14910,N_14870);
and U15158 (N_15158,N_14799,N_14669);
xnor U15159 (N_15159,N_14756,N_14791);
nand U15160 (N_15160,N_14668,N_14691);
nand U15161 (N_15161,N_14597,N_14994);
nand U15162 (N_15162,N_14803,N_14971);
nand U15163 (N_15163,N_14913,N_14986);
nand U15164 (N_15164,N_14639,N_14615);
and U15165 (N_15165,N_14715,N_14738);
nand U15166 (N_15166,N_14720,N_14606);
or U15167 (N_15167,N_14812,N_14919);
nand U15168 (N_15168,N_14736,N_14573);
and U15169 (N_15169,N_14768,N_14918);
nor U15170 (N_15170,N_14754,N_14631);
or U15171 (N_15171,N_14747,N_14679);
nor U15172 (N_15172,N_14591,N_14560);
or U15173 (N_15173,N_14975,N_14796);
nor U15174 (N_15174,N_14962,N_14646);
nor U15175 (N_15175,N_14703,N_14960);
nor U15176 (N_15176,N_14735,N_14782);
nand U15177 (N_15177,N_14695,N_14775);
nor U15178 (N_15178,N_14602,N_14909);
nor U15179 (N_15179,N_14865,N_14980);
and U15180 (N_15180,N_14748,N_14855);
nand U15181 (N_15181,N_14505,N_14815);
or U15182 (N_15182,N_14541,N_14564);
nand U15183 (N_15183,N_14906,N_14826);
and U15184 (N_15184,N_14749,N_14513);
and U15185 (N_15185,N_14674,N_14851);
or U15186 (N_15186,N_14900,N_14916);
nand U15187 (N_15187,N_14645,N_14653);
xor U15188 (N_15188,N_14925,N_14716);
and U15189 (N_15189,N_14901,N_14520);
and U15190 (N_15190,N_14833,N_14770);
nor U15191 (N_15191,N_14936,N_14578);
or U15192 (N_15192,N_14743,N_14752);
and U15193 (N_15193,N_14758,N_14816);
nor U15194 (N_15194,N_14751,N_14966);
nor U15195 (N_15195,N_14725,N_14973);
nor U15196 (N_15196,N_14968,N_14711);
or U15197 (N_15197,N_14614,N_14731);
nand U15198 (N_15198,N_14780,N_14896);
xor U15199 (N_15199,N_14545,N_14792);
or U15200 (N_15200,N_14589,N_14570);
nand U15201 (N_15201,N_14842,N_14806);
nand U15202 (N_15202,N_14524,N_14698);
or U15203 (N_15203,N_14729,N_14937);
and U15204 (N_15204,N_14863,N_14809);
and U15205 (N_15205,N_14563,N_14739);
nor U15206 (N_15206,N_14854,N_14737);
and U15207 (N_15207,N_14632,N_14786);
nand U15208 (N_15208,N_14684,N_14899);
or U15209 (N_15209,N_14965,N_14964);
or U15210 (N_15210,N_14831,N_14503);
nand U15211 (N_15211,N_14759,N_14897);
or U15212 (N_15212,N_14761,N_14805);
nand U15213 (N_15213,N_14924,N_14690);
nor U15214 (N_15214,N_14888,N_14813);
nand U15215 (N_15215,N_14558,N_14527);
nand U15216 (N_15216,N_14635,N_14717);
and U15217 (N_15217,N_14599,N_14672);
nor U15218 (N_15218,N_14647,N_14576);
nand U15219 (N_15219,N_14978,N_14904);
xnor U15220 (N_15220,N_14856,N_14885);
or U15221 (N_15221,N_14979,N_14777);
nand U15222 (N_15222,N_14923,N_14709);
and U15223 (N_15223,N_14982,N_14797);
and U15224 (N_15224,N_14838,N_14514);
nor U15225 (N_15225,N_14993,N_14850);
or U15226 (N_15226,N_14746,N_14554);
and U15227 (N_15227,N_14593,N_14686);
and U15228 (N_15228,N_14836,N_14603);
or U15229 (N_15229,N_14604,N_14769);
nor U15230 (N_15230,N_14956,N_14537);
and U15231 (N_15231,N_14773,N_14610);
and U15232 (N_15232,N_14767,N_14700);
or U15233 (N_15233,N_14905,N_14529);
nand U15234 (N_15234,N_14559,N_14961);
or U15235 (N_15235,N_14844,N_14567);
or U15236 (N_15236,N_14584,N_14616);
nand U15237 (N_15237,N_14783,N_14788);
and U15238 (N_15238,N_14687,N_14757);
or U15239 (N_15239,N_14658,N_14590);
nor U15240 (N_15240,N_14950,N_14902);
nand U15241 (N_15241,N_14638,N_14915);
nor U15242 (N_15242,N_14991,N_14874);
nand U15243 (N_15243,N_14676,N_14963);
nor U15244 (N_15244,N_14734,N_14867);
nor U15245 (N_15245,N_14929,N_14787);
nand U15246 (N_15246,N_14884,N_14877);
and U15247 (N_15247,N_14634,N_14566);
nor U15248 (N_15248,N_14886,N_14630);
or U15249 (N_15249,N_14664,N_14984);
or U15250 (N_15250,N_14883,N_14807);
nand U15251 (N_15251,N_14989,N_14946);
nand U15252 (N_15252,N_14644,N_14988);
nor U15253 (N_15253,N_14634,N_14581);
or U15254 (N_15254,N_14853,N_14800);
nor U15255 (N_15255,N_14775,N_14779);
or U15256 (N_15256,N_14867,N_14745);
or U15257 (N_15257,N_14750,N_14931);
and U15258 (N_15258,N_14887,N_14924);
nand U15259 (N_15259,N_14823,N_14982);
nand U15260 (N_15260,N_14992,N_14896);
nor U15261 (N_15261,N_14670,N_14661);
xor U15262 (N_15262,N_14795,N_14883);
nor U15263 (N_15263,N_14943,N_14946);
nand U15264 (N_15264,N_14502,N_14949);
and U15265 (N_15265,N_14887,N_14830);
xor U15266 (N_15266,N_14627,N_14596);
nor U15267 (N_15267,N_14648,N_14550);
nor U15268 (N_15268,N_14546,N_14905);
or U15269 (N_15269,N_14936,N_14590);
nand U15270 (N_15270,N_14954,N_14730);
and U15271 (N_15271,N_14987,N_14978);
and U15272 (N_15272,N_14916,N_14954);
or U15273 (N_15273,N_14939,N_14981);
nand U15274 (N_15274,N_14779,N_14676);
and U15275 (N_15275,N_14656,N_14749);
xor U15276 (N_15276,N_14548,N_14607);
nand U15277 (N_15277,N_14555,N_14997);
xor U15278 (N_15278,N_14685,N_14687);
nor U15279 (N_15279,N_14758,N_14838);
nand U15280 (N_15280,N_14560,N_14955);
xor U15281 (N_15281,N_14519,N_14651);
or U15282 (N_15282,N_14987,N_14871);
nand U15283 (N_15283,N_14679,N_14812);
nand U15284 (N_15284,N_14530,N_14851);
nand U15285 (N_15285,N_14880,N_14697);
xor U15286 (N_15286,N_14845,N_14904);
or U15287 (N_15287,N_14554,N_14643);
nand U15288 (N_15288,N_14626,N_14529);
nor U15289 (N_15289,N_14910,N_14634);
and U15290 (N_15290,N_14796,N_14727);
or U15291 (N_15291,N_14617,N_14841);
xnor U15292 (N_15292,N_14692,N_14836);
or U15293 (N_15293,N_14718,N_14568);
xor U15294 (N_15294,N_14555,N_14503);
nor U15295 (N_15295,N_14632,N_14704);
nand U15296 (N_15296,N_14775,N_14882);
or U15297 (N_15297,N_14630,N_14976);
nand U15298 (N_15298,N_14652,N_14873);
nor U15299 (N_15299,N_14612,N_14723);
or U15300 (N_15300,N_14971,N_14879);
nand U15301 (N_15301,N_14976,N_14832);
nand U15302 (N_15302,N_14880,N_14677);
or U15303 (N_15303,N_14930,N_14864);
nor U15304 (N_15304,N_14915,N_14860);
nand U15305 (N_15305,N_14574,N_14744);
or U15306 (N_15306,N_14995,N_14965);
nand U15307 (N_15307,N_14676,N_14719);
or U15308 (N_15308,N_14715,N_14589);
nor U15309 (N_15309,N_14977,N_14516);
and U15310 (N_15310,N_14629,N_14643);
and U15311 (N_15311,N_14781,N_14846);
or U15312 (N_15312,N_14758,N_14542);
and U15313 (N_15313,N_14690,N_14596);
and U15314 (N_15314,N_14565,N_14785);
nand U15315 (N_15315,N_14547,N_14957);
or U15316 (N_15316,N_14724,N_14515);
or U15317 (N_15317,N_14794,N_14610);
nand U15318 (N_15318,N_14641,N_14657);
nor U15319 (N_15319,N_14563,N_14521);
nor U15320 (N_15320,N_14523,N_14656);
xnor U15321 (N_15321,N_14754,N_14798);
and U15322 (N_15322,N_14982,N_14731);
nand U15323 (N_15323,N_14854,N_14575);
nand U15324 (N_15324,N_14860,N_14508);
nor U15325 (N_15325,N_14842,N_14944);
nand U15326 (N_15326,N_14695,N_14508);
and U15327 (N_15327,N_14830,N_14911);
nand U15328 (N_15328,N_14950,N_14997);
nor U15329 (N_15329,N_14537,N_14932);
xnor U15330 (N_15330,N_14959,N_14524);
and U15331 (N_15331,N_14643,N_14885);
nor U15332 (N_15332,N_14860,N_14776);
and U15333 (N_15333,N_14589,N_14954);
nand U15334 (N_15334,N_14711,N_14653);
nor U15335 (N_15335,N_14615,N_14886);
nor U15336 (N_15336,N_14532,N_14549);
and U15337 (N_15337,N_14800,N_14889);
and U15338 (N_15338,N_14633,N_14720);
nand U15339 (N_15339,N_14947,N_14796);
or U15340 (N_15340,N_14688,N_14942);
or U15341 (N_15341,N_14644,N_14867);
nor U15342 (N_15342,N_14832,N_14931);
or U15343 (N_15343,N_14522,N_14837);
and U15344 (N_15344,N_14992,N_14720);
xnor U15345 (N_15345,N_14812,N_14603);
or U15346 (N_15346,N_14619,N_14862);
or U15347 (N_15347,N_14548,N_14610);
xnor U15348 (N_15348,N_14827,N_14918);
nand U15349 (N_15349,N_14666,N_14911);
xnor U15350 (N_15350,N_14593,N_14560);
or U15351 (N_15351,N_14894,N_14890);
or U15352 (N_15352,N_14858,N_14856);
nor U15353 (N_15353,N_14924,N_14759);
nand U15354 (N_15354,N_14944,N_14919);
xnor U15355 (N_15355,N_14678,N_14518);
nand U15356 (N_15356,N_14930,N_14772);
nand U15357 (N_15357,N_14822,N_14695);
xor U15358 (N_15358,N_14798,N_14760);
or U15359 (N_15359,N_14684,N_14950);
and U15360 (N_15360,N_14617,N_14940);
nor U15361 (N_15361,N_14812,N_14799);
nand U15362 (N_15362,N_14586,N_14500);
or U15363 (N_15363,N_14711,N_14961);
and U15364 (N_15364,N_14701,N_14570);
xor U15365 (N_15365,N_14838,N_14919);
and U15366 (N_15366,N_14564,N_14702);
nor U15367 (N_15367,N_14568,N_14653);
or U15368 (N_15368,N_14791,N_14764);
and U15369 (N_15369,N_14524,N_14727);
nand U15370 (N_15370,N_14776,N_14547);
nand U15371 (N_15371,N_14612,N_14755);
or U15372 (N_15372,N_14699,N_14733);
nand U15373 (N_15373,N_14741,N_14941);
nand U15374 (N_15374,N_14618,N_14562);
and U15375 (N_15375,N_14870,N_14588);
or U15376 (N_15376,N_14843,N_14888);
nand U15377 (N_15377,N_14943,N_14526);
and U15378 (N_15378,N_14890,N_14793);
nand U15379 (N_15379,N_14906,N_14601);
nor U15380 (N_15380,N_14679,N_14694);
xnor U15381 (N_15381,N_14616,N_14893);
or U15382 (N_15382,N_14576,N_14812);
nand U15383 (N_15383,N_14911,N_14861);
nor U15384 (N_15384,N_14935,N_14562);
xnor U15385 (N_15385,N_14815,N_14803);
or U15386 (N_15386,N_14556,N_14934);
nand U15387 (N_15387,N_14683,N_14836);
or U15388 (N_15388,N_14782,N_14993);
and U15389 (N_15389,N_14628,N_14745);
nor U15390 (N_15390,N_14893,N_14746);
or U15391 (N_15391,N_14908,N_14562);
or U15392 (N_15392,N_14774,N_14888);
and U15393 (N_15393,N_14794,N_14601);
nor U15394 (N_15394,N_14842,N_14633);
nand U15395 (N_15395,N_14731,N_14788);
or U15396 (N_15396,N_14939,N_14705);
and U15397 (N_15397,N_14504,N_14883);
and U15398 (N_15398,N_14548,N_14730);
or U15399 (N_15399,N_14958,N_14520);
or U15400 (N_15400,N_14521,N_14736);
nand U15401 (N_15401,N_14506,N_14565);
nor U15402 (N_15402,N_14955,N_14743);
and U15403 (N_15403,N_14577,N_14524);
and U15404 (N_15404,N_14929,N_14901);
nor U15405 (N_15405,N_14539,N_14588);
xnor U15406 (N_15406,N_14976,N_14669);
and U15407 (N_15407,N_14988,N_14854);
nor U15408 (N_15408,N_14508,N_14802);
nand U15409 (N_15409,N_14563,N_14890);
or U15410 (N_15410,N_14598,N_14970);
or U15411 (N_15411,N_14805,N_14985);
nand U15412 (N_15412,N_14706,N_14664);
and U15413 (N_15413,N_14777,N_14904);
and U15414 (N_15414,N_14513,N_14967);
and U15415 (N_15415,N_14849,N_14570);
xor U15416 (N_15416,N_14744,N_14790);
nor U15417 (N_15417,N_14649,N_14546);
or U15418 (N_15418,N_14592,N_14692);
or U15419 (N_15419,N_14562,N_14708);
and U15420 (N_15420,N_14685,N_14948);
or U15421 (N_15421,N_14776,N_14965);
nor U15422 (N_15422,N_14710,N_14885);
nor U15423 (N_15423,N_14722,N_14749);
and U15424 (N_15424,N_14810,N_14531);
nand U15425 (N_15425,N_14977,N_14856);
nand U15426 (N_15426,N_14614,N_14846);
and U15427 (N_15427,N_14577,N_14530);
or U15428 (N_15428,N_14698,N_14930);
nor U15429 (N_15429,N_14509,N_14620);
nand U15430 (N_15430,N_14877,N_14992);
or U15431 (N_15431,N_14655,N_14711);
nor U15432 (N_15432,N_14968,N_14937);
nand U15433 (N_15433,N_14792,N_14639);
and U15434 (N_15434,N_14797,N_14893);
nand U15435 (N_15435,N_14931,N_14599);
xnor U15436 (N_15436,N_14742,N_14642);
nand U15437 (N_15437,N_14979,N_14665);
nor U15438 (N_15438,N_14752,N_14542);
nand U15439 (N_15439,N_14779,N_14528);
nor U15440 (N_15440,N_14871,N_14602);
nand U15441 (N_15441,N_14665,N_14521);
or U15442 (N_15442,N_14864,N_14612);
and U15443 (N_15443,N_14583,N_14933);
or U15444 (N_15444,N_14609,N_14534);
or U15445 (N_15445,N_14993,N_14716);
and U15446 (N_15446,N_14586,N_14898);
xnor U15447 (N_15447,N_14601,N_14542);
nand U15448 (N_15448,N_14516,N_14596);
or U15449 (N_15449,N_14639,N_14585);
or U15450 (N_15450,N_14580,N_14825);
or U15451 (N_15451,N_14658,N_14682);
xnor U15452 (N_15452,N_14507,N_14867);
and U15453 (N_15453,N_14732,N_14519);
nand U15454 (N_15454,N_14766,N_14984);
nand U15455 (N_15455,N_14545,N_14517);
or U15456 (N_15456,N_14869,N_14862);
xnor U15457 (N_15457,N_14508,N_14611);
nor U15458 (N_15458,N_14569,N_14812);
nand U15459 (N_15459,N_14704,N_14776);
nand U15460 (N_15460,N_14870,N_14946);
or U15461 (N_15461,N_14742,N_14876);
and U15462 (N_15462,N_14885,N_14725);
nor U15463 (N_15463,N_14964,N_14842);
nand U15464 (N_15464,N_14735,N_14898);
or U15465 (N_15465,N_14935,N_14881);
nand U15466 (N_15466,N_14793,N_14797);
nand U15467 (N_15467,N_14660,N_14835);
nand U15468 (N_15468,N_14685,N_14964);
nor U15469 (N_15469,N_14931,N_14514);
nand U15470 (N_15470,N_14987,N_14916);
or U15471 (N_15471,N_14753,N_14525);
or U15472 (N_15472,N_14962,N_14893);
nand U15473 (N_15473,N_14543,N_14926);
nand U15474 (N_15474,N_14877,N_14750);
and U15475 (N_15475,N_14953,N_14505);
nor U15476 (N_15476,N_14610,N_14820);
or U15477 (N_15477,N_14975,N_14718);
nor U15478 (N_15478,N_14779,N_14803);
or U15479 (N_15479,N_14794,N_14600);
and U15480 (N_15480,N_14866,N_14624);
nor U15481 (N_15481,N_14564,N_14998);
and U15482 (N_15482,N_14710,N_14844);
and U15483 (N_15483,N_14897,N_14826);
and U15484 (N_15484,N_14768,N_14760);
or U15485 (N_15485,N_14935,N_14816);
nand U15486 (N_15486,N_14663,N_14930);
nand U15487 (N_15487,N_14545,N_14971);
or U15488 (N_15488,N_14634,N_14883);
nor U15489 (N_15489,N_14951,N_14902);
nand U15490 (N_15490,N_14619,N_14998);
and U15491 (N_15491,N_14629,N_14740);
or U15492 (N_15492,N_14617,N_14648);
nor U15493 (N_15493,N_14748,N_14923);
nor U15494 (N_15494,N_14506,N_14683);
nor U15495 (N_15495,N_14801,N_14887);
or U15496 (N_15496,N_14674,N_14614);
nand U15497 (N_15497,N_14545,N_14711);
and U15498 (N_15498,N_14638,N_14566);
and U15499 (N_15499,N_14577,N_14699);
xnor U15500 (N_15500,N_15300,N_15322);
or U15501 (N_15501,N_15410,N_15425);
or U15502 (N_15502,N_15053,N_15350);
nand U15503 (N_15503,N_15383,N_15213);
nand U15504 (N_15504,N_15420,N_15223);
nand U15505 (N_15505,N_15407,N_15156);
nand U15506 (N_15506,N_15480,N_15179);
or U15507 (N_15507,N_15470,N_15263);
nand U15508 (N_15508,N_15095,N_15105);
and U15509 (N_15509,N_15332,N_15282);
nand U15510 (N_15510,N_15180,N_15098);
and U15511 (N_15511,N_15488,N_15139);
and U15512 (N_15512,N_15284,N_15008);
and U15513 (N_15513,N_15477,N_15352);
or U15514 (N_15514,N_15133,N_15230);
nand U15515 (N_15515,N_15247,N_15195);
xnor U15516 (N_15516,N_15413,N_15244);
nand U15517 (N_15517,N_15146,N_15398);
or U15518 (N_15518,N_15038,N_15191);
and U15519 (N_15519,N_15475,N_15082);
or U15520 (N_15520,N_15207,N_15074);
or U15521 (N_15521,N_15461,N_15439);
nor U15522 (N_15522,N_15498,N_15323);
and U15523 (N_15523,N_15443,N_15108);
nand U15524 (N_15524,N_15453,N_15170);
nand U15525 (N_15525,N_15217,N_15204);
or U15526 (N_15526,N_15142,N_15232);
or U15527 (N_15527,N_15335,N_15456);
nor U15528 (N_15528,N_15444,N_15062);
and U15529 (N_15529,N_15483,N_15325);
or U15530 (N_15530,N_15474,N_15399);
nor U15531 (N_15531,N_15248,N_15137);
xnor U15532 (N_15532,N_15120,N_15035);
or U15533 (N_15533,N_15274,N_15406);
xnor U15534 (N_15534,N_15411,N_15491);
and U15535 (N_15535,N_15097,N_15434);
nor U15536 (N_15536,N_15058,N_15397);
nor U15537 (N_15537,N_15451,N_15345);
and U15538 (N_15538,N_15216,N_15200);
and U15539 (N_15539,N_15455,N_15479);
or U15540 (N_15540,N_15418,N_15319);
nand U15541 (N_15541,N_15476,N_15002);
nand U15542 (N_15542,N_15310,N_15360);
xor U15543 (N_15543,N_15061,N_15011);
and U15544 (N_15544,N_15029,N_15103);
or U15545 (N_15545,N_15018,N_15070);
and U15546 (N_15546,N_15184,N_15405);
nor U15547 (N_15547,N_15093,N_15465);
nor U15548 (N_15548,N_15177,N_15329);
and U15549 (N_15549,N_15452,N_15346);
and U15550 (N_15550,N_15118,N_15203);
or U15551 (N_15551,N_15412,N_15013);
nor U15552 (N_15552,N_15327,N_15076);
xnor U15553 (N_15553,N_15492,N_15250);
and U15554 (N_15554,N_15404,N_15078);
or U15555 (N_15555,N_15010,N_15127);
nor U15556 (N_15556,N_15278,N_15303);
or U15557 (N_15557,N_15027,N_15054);
or U15558 (N_15558,N_15471,N_15432);
nand U15559 (N_15559,N_15158,N_15342);
xor U15560 (N_15560,N_15004,N_15264);
and U15561 (N_15561,N_15429,N_15026);
xnor U15562 (N_15562,N_15286,N_15424);
and U15563 (N_15563,N_15427,N_15005);
and U15564 (N_15564,N_15357,N_15355);
xnor U15565 (N_15565,N_15311,N_15140);
nor U15566 (N_15566,N_15386,N_15065);
or U15567 (N_15567,N_15241,N_15238);
and U15568 (N_15568,N_15132,N_15292);
nand U15569 (N_15569,N_15481,N_15153);
nand U15570 (N_15570,N_15317,N_15122);
and U15571 (N_15571,N_15090,N_15316);
nor U15572 (N_15572,N_15369,N_15421);
and U15573 (N_15573,N_15163,N_15275);
and U15574 (N_15574,N_15089,N_15116);
and U15575 (N_15575,N_15102,N_15440);
nand U15576 (N_15576,N_15447,N_15025);
and U15577 (N_15577,N_15178,N_15099);
or U15578 (N_15578,N_15057,N_15148);
and U15579 (N_15579,N_15245,N_15436);
and U15580 (N_15580,N_15437,N_15174);
xor U15581 (N_15581,N_15121,N_15144);
or U15582 (N_15582,N_15258,N_15151);
and U15583 (N_15583,N_15277,N_15229);
xnor U15584 (N_15584,N_15171,N_15273);
nand U15585 (N_15585,N_15254,N_15106);
or U15586 (N_15586,N_15150,N_15086);
nand U15587 (N_15587,N_15463,N_15496);
or U15588 (N_15588,N_15462,N_15364);
or U15589 (N_15589,N_15333,N_15305);
nor U15590 (N_15590,N_15377,N_15012);
or U15591 (N_15591,N_15014,N_15285);
nor U15592 (N_15592,N_15110,N_15215);
or U15593 (N_15593,N_15314,N_15324);
and U15594 (N_15594,N_15166,N_15194);
xor U15595 (N_15595,N_15081,N_15395);
nor U15596 (N_15596,N_15328,N_15354);
and U15597 (N_15597,N_15157,N_15376);
nand U15598 (N_15598,N_15448,N_15192);
nand U15599 (N_15599,N_15188,N_15490);
xnor U15600 (N_15600,N_15290,N_15403);
or U15601 (N_15601,N_15445,N_15365);
nand U15602 (N_15602,N_15276,N_15270);
xnor U15603 (N_15603,N_15234,N_15176);
nor U15604 (N_15604,N_15006,N_15287);
nand U15605 (N_15605,N_15293,N_15031);
nor U15606 (N_15606,N_15123,N_15391);
nand U15607 (N_15607,N_15467,N_15366);
nand U15608 (N_15608,N_15077,N_15288);
nor U15609 (N_15609,N_15349,N_15092);
nor U15610 (N_15610,N_15155,N_15128);
nand U15611 (N_15611,N_15225,N_15181);
or U15612 (N_15612,N_15469,N_15135);
nor U15613 (N_15613,N_15392,N_15104);
or U15614 (N_15614,N_15036,N_15279);
nand U15615 (N_15615,N_15396,N_15208);
or U15616 (N_15616,N_15214,N_15473);
or U15617 (N_15617,N_15302,N_15117);
nor U15618 (N_15618,N_15037,N_15197);
and U15619 (N_15619,N_15338,N_15400);
or U15620 (N_15620,N_15115,N_15206);
nor U15621 (N_15621,N_15222,N_15199);
nor U15622 (N_15622,N_15262,N_15382);
or U15623 (N_15623,N_15259,N_15107);
nor U15624 (N_15624,N_15172,N_15007);
and U15625 (N_15625,N_15347,N_15313);
and U15626 (N_15626,N_15266,N_15186);
nor U15627 (N_15627,N_15064,N_15240);
or U15628 (N_15628,N_15066,N_15318);
nor U15629 (N_15629,N_15435,N_15417);
nand U15630 (N_15630,N_15226,N_15353);
xor U15631 (N_15631,N_15472,N_15138);
and U15632 (N_15632,N_15009,N_15367);
or U15633 (N_15633,N_15201,N_15051);
or U15634 (N_15634,N_15205,N_15049);
nor U15635 (N_15635,N_15315,N_15246);
nor U15636 (N_15636,N_15450,N_15283);
nor U15637 (N_15637,N_15019,N_15260);
nor U15638 (N_15638,N_15046,N_15265);
or U15639 (N_15639,N_15164,N_15209);
nor U15640 (N_15640,N_15084,N_15261);
nor U15641 (N_15641,N_15182,N_15457);
nand U15642 (N_15642,N_15017,N_15141);
and U15643 (N_15643,N_15296,N_15361);
nand U15644 (N_15644,N_15045,N_15096);
xor U15645 (N_15645,N_15190,N_15175);
nor U15646 (N_15646,N_15268,N_15060);
nor U15647 (N_15647,N_15001,N_15301);
nand U15648 (N_15648,N_15034,N_15289);
or U15649 (N_15649,N_15071,N_15087);
xnor U15650 (N_15650,N_15373,N_15372);
nor U15651 (N_15651,N_15252,N_15485);
or U15652 (N_15652,N_15210,N_15196);
nor U15653 (N_15653,N_15253,N_15295);
or U15654 (N_15654,N_15494,N_15080);
nand U15655 (N_15655,N_15402,N_15185);
or U15656 (N_15656,N_15446,N_15042);
xnor U15657 (N_15657,N_15239,N_15000);
xor U15658 (N_15658,N_15114,N_15454);
nand U15659 (N_15659,N_15337,N_15330);
and U15660 (N_15660,N_15079,N_15242);
and U15661 (N_15661,N_15458,N_15497);
and U15662 (N_15662,N_15183,N_15272);
nor U15663 (N_15663,N_15433,N_15257);
nor U15664 (N_15664,N_15040,N_15339);
nor U15665 (N_15665,N_15236,N_15228);
or U15666 (N_15666,N_15218,N_15160);
xor U15667 (N_15667,N_15023,N_15161);
nor U15668 (N_15668,N_15358,N_15052);
nand U15669 (N_15669,N_15393,N_15168);
and U15670 (N_15670,N_15466,N_15422);
and U15671 (N_15671,N_15423,N_15482);
nand U15672 (N_15672,N_15237,N_15028);
nor U15673 (N_15673,N_15309,N_15388);
nor U15674 (N_15674,N_15020,N_15131);
nor U15675 (N_15675,N_15484,N_15033);
and U15676 (N_15676,N_15362,N_15370);
nand U15677 (N_15677,N_15428,N_15464);
or U15678 (N_15678,N_15359,N_15063);
or U15679 (N_15679,N_15231,N_15438);
nand U15680 (N_15680,N_15130,N_15032);
or U15681 (N_15681,N_15387,N_15016);
and U15682 (N_15682,N_15100,N_15235);
nor U15683 (N_15683,N_15224,N_15220);
nand U15684 (N_15684,N_15389,N_15489);
nand U15685 (N_15685,N_15430,N_15459);
or U15686 (N_15686,N_15415,N_15304);
or U15687 (N_15687,N_15147,N_15441);
nor U15688 (N_15688,N_15047,N_15055);
nand U15689 (N_15689,N_15426,N_15022);
nand U15690 (N_15690,N_15416,N_15212);
or U15691 (N_15691,N_15003,N_15308);
xnor U15692 (N_15692,N_15134,N_15041);
nor U15693 (N_15693,N_15075,N_15299);
nand U15694 (N_15694,N_15101,N_15294);
nand U15695 (N_15695,N_15380,N_15129);
and U15696 (N_15696,N_15401,N_15379);
nand U15697 (N_15697,N_15321,N_15149);
nand U15698 (N_15698,N_15187,N_15039);
nor U15699 (N_15699,N_15143,N_15243);
or U15700 (N_15700,N_15384,N_15291);
nor U15701 (N_15701,N_15043,N_15312);
nor U15702 (N_15702,N_15271,N_15189);
or U15703 (N_15703,N_15169,N_15331);
and U15704 (N_15704,N_15341,N_15371);
nand U15705 (N_15705,N_15162,N_15059);
or U15706 (N_15706,N_15499,N_15091);
nor U15707 (N_15707,N_15113,N_15340);
and U15708 (N_15708,N_15486,N_15109);
or U15709 (N_15709,N_15211,N_15085);
or U15710 (N_15710,N_15281,N_15449);
nor U15711 (N_15711,N_15326,N_15044);
xor U15712 (N_15712,N_15173,N_15126);
nor U15713 (N_15713,N_15348,N_15249);
or U15714 (N_15714,N_15255,N_15297);
xor U15715 (N_15715,N_15269,N_15021);
or U15716 (N_15716,N_15111,N_15154);
and U15717 (N_15717,N_15056,N_15320);
nand U15718 (N_15718,N_15374,N_15152);
and U15719 (N_15719,N_15159,N_15112);
or U15720 (N_15720,N_15306,N_15015);
or U15721 (N_15721,N_15094,N_15495);
nor U15722 (N_15722,N_15267,N_15219);
nand U15723 (N_15723,N_15073,N_15414);
nand U15724 (N_15724,N_15307,N_15487);
nor U15725 (N_15725,N_15493,N_15165);
and U15726 (N_15726,N_15381,N_15390);
nor U15727 (N_15727,N_15119,N_15048);
nor U15728 (N_15728,N_15068,N_15136);
nor U15729 (N_15729,N_15385,N_15334);
and U15730 (N_15730,N_15227,N_15088);
nand U15731 (N_15731,N_15408,N_15202);
or U15732 (N_15732,N_15030,N_15221);
xor U15733 (N_15733,N_15343,N_15083);
nor U15734 (N_15734,N_15442,N_15233);
nand U15735 (N_15735,N_15368,N_15193);
or U15736 (N_15736,N_15460,N_15024);
nand U15737 (N_15737,N_15256,N_15069);
and U15738 (N_15738,N_15378,N_15125);
or U15739 (N_15739,N_15419,N_15363);
or U15740 (N_15740,N_15375,N_15280);
and U15741 (N_15741,N_15198,N_15478);
nor U15742 (N_15742,N_15468,N_15167);
nor U15743 (N_15743,N_15356,N_15344);
and U15744 (N_15744,N_15298,N_15394);
nand U15745 (N_15745,N_15251,N_15067);
nor U15746 (N_15746,N_15124,N_15072);
or U15747 (N_15747,N_15431,N_15050);
nand U15748 (N_15748,N_15145,N_15351);
and U15749 (N_15749,N_15336,N_15409);
and U15750 (N_15750,N_15427,N_15356);
and U15751 (N_15751,N_15322,N_15304);
or U15752 (N_15752,N_15022,N_15035);
nor U15753 (N_15753,N_15350,N_15005);
and U15754 (N_15754,N_15263,N_15339);
xnor U15755 (N_15755,N_15235,N_15163);
or U15756 (N_15756,N_15474,N_15152);
and U15757 (N_15757,N_15235,N_15050);
xnor U15758 (N_15758,N_15252,N_15195);
nor U15759 (N_15759,N_15063,N_15429);
nor U15760 (N_15760,N_15242,N_15243);
nor U15761 (N_15761,N_15300,N_15431);
nand U15762 (N_15762,N_15084,N_15352);
or U15763 (N_15763,N_15469,N_15363);
nor U15764 (N_15764,N_15443,N_15287);
nand U15765 (N_15765,N_15356,N_15345);
or U15766 (N_15766,N_15319,N_15384);
nor U15767 (N_15767,N_15472,N_15032);
and U15768 (N_15768,N_15152,N_15280);
nor U15769 (N_15769,N_15132,N_15423);
nor U15770 (N_15770,N_15155,N_15212);
nor U15771 (N_15771,N_15115,N_15489);
nor U15772 (N_15772,N_15449,N_15053);
or U15773 (N_15773,N_15176,N_15101);
or U15774 (N_15774,N_15050,N_15361);
nor U15775 (N_15775,N_15494,N_15284);
nand U15776 (N_15776,N_15086,N_15137);
or U15777 (N_15777,N_15263,N_15270);
and U15778 (N_15778,N_15470,N_15134);
nand U15779 (N_15779,N_15082,N_15267);
and U15780 (N_15780,N_15050,N_15326);
nand U15781 (N_15781,N_15441,N_15095);
nor U15782 (N_15782,N_15183,N_15287);
and U15783 (N_15783,N_15087,N_15076);
xnor U15784 (N_15784,N_15119,N_15367);
nand U15785 (N_15785,N_15018,N_15113);
xnor U15786 (N_15786,N_15471,N_15105);
and U15787 (N_15787,N_15249,N_15246);
nor U15788 (N_15788,N_15317,N_15233);
nor U15789 (N_15789,N_15252,N_15209);
or U15790 (N_15790,N_15256,N_15377);
or U15791 (N_15791,N_15060,N_15279);
nand U15792 (N_15792,N_15090,N_15152);
nand U15793 (N_15793,N_15108,N_15026);
xnor U15794 (N_15794,N_15416,N_15082);
and U15795 (N_15795,N_15429,N_15133);
nor U15796 (N_15796,N_15038,N_15313);
nand U15797 (N_15797,N_15050,N_15184);
nor U15798 (N_15798,N_15015,N_15457);
nand U15799 (N_15799,N_15073,N_15165);
xnor U15800 (N_15800,N_15049,N_15203);
and U15801 (N_15801,N_15252,N_15038);
or U15802 (N_15802,N_15173,N_15005);
or U15803 (N_15803,N_15411,N_15446);
or U15804 (N_15804,N_15484,N_15258);
and U15805 (N_15805,N_15150,N_15364);
and U15806 (N_15806,N_15192,N_15274);
nand U15807 (N_15807,N_15089,N_15329);
nor U15808 (N_15808,N_15231,N_15041);
nor U15809 (N_15809,N_15091,N_15126);
nand U15810 (N_15810,N_15476,N_15347);
and U15811 (N_15811,N_15060,N_15105);
nor U15812 (N_15812,N_15244,N_15229);
nor U15813 (N_15813,N_15168,N_15435);
xor U15814 (N_15814,N_15412,N_15066);
nor U15815 (N_15815,N_15052,N_15312);
and U15816 (N_15816,N_15419,N_15413);
nor U15817 (N_15817,N_15252,N_15489);
nor U15818 (N_15818,N_15430,N_15470);
nor U15819 (N_15819,N_15172,N_15013);
xor U15820 (N_15820,N_15381,N_15486);
or U15821 (N_15821,N_15045,N_15420);
nor U15822 (N_15822,N_15339,N_15174);
nor U15823 (N_15823,N_15320,N_15160);
and U15824 (N_15824,N_15260,N_15451);
nand U15825 (N_15825,N_15167,N_15006);
nor U15826 (N_15826,N_15358,N_15308);
nand U15827 (N_15827,N_15331,N_15072);
xnor U15828 (N_15828,N_15168,N_15489);
nor U15829 (N_15829,N_15080,N_15046);
nor U15830 (N_15830,N_15334,N_15410);
or U15831 (N_15831,N_15097,N_15407);
or U15832 (N_15832,N_15197,N_15349);
and U15833 (N_15833,N_15405,N_15153);
and U15834 (N_15834,N_15262,N_15352);
nand U15835 (N_15835,N_15044,N_15066);
nor U15836 (N_15836,N_15304,N_15158);
nand U15837 (N_15837,N_15204,N_15096);
nand U15838 (N_15838,N_15137,N_15259);
or U15839 (N_15839,N_15097,N_15465);
nor U15840 (N_15840,N_15256,N_15099);
or U15841 (N_15841,N_15316,N_15348);
nand U15842 (N_15842,N_15146,N_15380);
nor U15843 (N_15843,N_15103,N_15118);
or U15844 (N_15844,N_15440,N_15130);
nand U15845 (N_15845,N_15410,N_15231);
and U15846 (N_15846,N_15351,N_15053);
or U15847 (N_15847,N_15237,N_15068);
nand U15848 (N_15848,N_15060,N_15433);
or U15849 (N_15849,N_15483,N_15068);
or U15850 (N_15850,N_15375,N_15435);
xor U15851 (N_15851,N_15218,N_15149);
nand U15852 (N_15852,N_15122,N_15389);
or U15853 (N_15853,N_15251,N_15090);
nor U15854 (N_15854,N_15136,N_15418);
and U15855 (N_15855,N_15255,N_15193);
or U15856 (N_15856,N_15370,N_15175);
or U15857 (N_15857,N_15054,N_15352);
and U15858 (N_15858,N_15226,N_15378);
and U15859 (N_15859,N_15022,N_15473);
and U15860 (N_15860,N_15371,N_15454);
nand U15861 (N_15861,N_15258,N_15407);
nor U15862 (N_15862,N_15144,N_15265);
xor U15863 (N_15863,N_15473,N_15064);
or U15864 (N_15864,N_15420,N_15349);
nand U15865 (N_15865,N_15119,N_15000);
nor U15866 (N_15866,N_15433,N_15296);
nand U15867 (N_15867,N_15434,N_15309);
or U15868 (N_15868,N_15122,N_15283);
xor U15869 (N_15869,N_15471,N_15192);
nand U15870 (N_15870,N_15435,N_15318);
or U15871 (N_15871,N_15006,N_15205);
or U15872 (N_15872,N_15385,N_15386);
nand U15873 (N_15873,N_15260,N_15278);
nor U15874 (N_15874,N_15133,N_15292);
and U15875 (N_15875,N_15307,N_15494);
or U15876 (N_15876,N_15176,N_15098);
and U15877 (N_15877,N_15365,N_15236);
nor U15878 (N_15878,N_15097,N_15305);
nand U15879 (N_15879,N_15216,N_15348);
nor U15880 (N_15880,N_15200,N_15001);
or U15881 (N_15881,N_15103,N_15230);
or U15882 (N_15882,N_15046,N_15389);
nor U15883 (N_15883,N_15278,N_15244);
and U15884 (N_15884,N_15341,N_15315);
and U15885 (N_15885,N_15067,N_15479);
nand U15886 (N_15886,N_15282,N_15468);
or U15887 (N_15887,N_15022,N_15449);
nor U15888 (N_15888,N_15023,N_15342);
nand U15889 (N_15889,N_15468,N_15381);
or U15890 (N_15890,N_15231,N_15252);
nor U15891 (N_15891,N_15149,N_15158);
nor U15892 (N_15892,N_15115,N_15213);
and U15893 (N_15893,N_15068,N_15264);
nand U15894 (N_15894,N_15345,N_15122);
nor U15895 (N_15895,N_15352,N_15327);
and U15896 (N_15896,N_15021,N_15479);
nor U15897 (N_15897,N_15439,N_15368);
nand U15898 (N_15898,N_15031,N_15180);
nand U15899 (N_15899,N_15060,N_15014);
and U15900 (N_15900,N_15115,N_15495);
and U15901 (N_15901,N_15142,N_15047);
or U15902 (N_15902,N_15187,N_15217);
nand U15903 (N_15903,N_15002,N_15115);
xnor U15904 (N_15904,N_15051,N_15126);
or U15905 (N_15905,N_15107,N_15069);
or U15906 (N_15906,N_15181,N_15203);
xor U15907 (N_15907,N_15487,N_15402);
nand U15908 (N_15908,N_15179,N_15366);
and U15909 (N_15909,N_15294,N_15031);
or U15910 (N_15910,N_15033,N_15073);
nand U15911 (N_15911,N_15237,N_15094);
and U15912 (N_15912,N_15228,N_15139);
and U15913 (N_15913,N_15055,N_15256);
and U15914 (N_15914,N_15312,N_15217);
nand U15915 (N_15915,N_15016,N_15266);
xnor U15916 (N_15916,N_15038,N_15400);
nand U15917 (N_15917,N_15055,N_15152);
xnor U15918 (N_15918,N_15258,N_15499);
nor U15919 (N_15919,N_15395,N_15498);
xnor U15920 (N_15920,N_15440,N_15298);
and U15921 (N_15921,N_15071,N_15445);
nor U15922 (N_15922,N_15311,N_15065);
nor U15923 (N_15923,N_15191,N_15158);
and U15924 (N_15924,N_15186,N_15372);
nand U15925 (N_15925,N_15289,N_15272);
or U15926 (N_15926,N_15259,N_15486);
nand U15927 (N_15927,N_15225,N_15102);
or U15928 (N_15928,N_15024,N_15483);
nand U15929 (N_15929,N_15198,N_15209);
and U15930 (N_15930,N_15158,N_15190);
or U15931 (N_15931,N_15088,N_15098);
nor U15932 (N_15932,N_15185,N_15260);
or U15933 (N_15933,N_15290,N_15413);
and U15934 (N_15934,N_15215,N_15112);
xor U15935 (N_15935,N_15429,N_15417);
nor U15936 (N_15936,N_15398,N_15023);
or U15937 (N_15937,N_15237,N_15242);
nand U15938 (N_15938,N_15322,N_15256);
xnor U15939 (N_15939,N_15030,N_15348);
nand U15940 (N_15940,N_15338,N_15065);
or U15941 (N_15941,N_15191,N_15256);
or U15942 (N_15942,N_15284,N_15384);
or U15943 (N_15943,N_15218,N_15301);
and U15944 (N_15944,N_15294,N_15338);
nand U15945 (N_15945,N_15432,N_15438);
or U15946 (N_15946,N_15276,N_15010);
nor U15947 (N_15947,N_15276,N_15252);
and U15948 (N_15948,N_15076,N_15114);
or U15949 (N_15949,N_15154,N_15446);
and U15950 (N_15950,N_15123,N_15316);
and U15951 (N_15951,N_15395,N_15380);
and U15952 (N_15952,N_15324,N_15057);
nor U15953 (N_15953,N_15296,N_15386);
nand U15954 (N_15954,N_15292,N_15399);
nor U15955 (N_15955,N_15100,N_15346);
nand U15956 (N_15956,N_15052,N_15275);
nor U15957 (N_15957,N_15082,N_15387);
or U15958 (N_15958,N_15031,N_15414);
and U15959 (N_15959,N_15294,N_15005);
and U15960 (N_15960,N_15419,N_15479);
nor U15961 (N_15961,N_15408,N_15384);
or U15962 (N_15962,N_15005,N_15453);
nor U15963 (N_15963,N_15268,N_15330);
nor U15964 (N_15964,N_15268,N_15138);
and U15965 (N_15965,N_15187,N_15201);
nand U15966 (N_15966,N_15277,N_15044);
and U15967 (N_15967,N_15066,N_15045);
nor U15968 (N_15968,N_15129,N_15046);
nor U15969 (N_15969,N_15077,N_15376);
or U15970 (N_15970,N_15143,N_15317);
and U15971 (N_15971,N_15471,N_15112);
or U15972 (N_15972,N_15288,N_15350);
or U15973 (N_15973,N_15061,N_15092);
nor U15974 (N_15974,N_15016,N_15427);
nor U15975 (N_15975,N_15006,N_15344);
and U15976 (N_15976,N_15125,N_15068);
and U15977 (N_15977,N_15244,N_15132);
nand U15978 (N_15978,N_15094,N_15379);
or U15979 (N_15979,N_15076,N_15469);
and U15980 (N_15980,N_15489,N_15444);
nand U15981 (N_15981,N_15410,N_15387);
and U15982 (N_15982,N_15369,N_15334);
nor U15983 (N_15983,N_15228,N_15484);
xnor U15984 (N_15984,N_15189,N_15279);
nor U15985 (N_15985,N_15494,N_15355);
or U15986 (N_15986,N_15347,N_15158);
or U15987 (N_15987,N_15294,N_15449);
nor U15988 (N_15988,N_15403,N_15127);
and U15989 (N_15989,N_15018,N_15042);
and U15990 (N_15990,N_15404,N_15073);
nor U15991 (N_15991,N_15493,N_15062);
nor U15992 (N_15992,N_15012,N_15175);
or U15993 (N_15993,N_15304,N_15266);
nand U15994 (N_15994,N_15149,N_15012);
or U15995 (N_15995,N_15054,N_15037);
nand U15996 (N_15996,N_15053,N_15488);
and U15997 (N_15997,N_15278,N_15407);
nor U15998 (N_15998,N_15266,N_15014);
or U15999 (N_15999,N_15127,N_15018);
nand U16000 (N_16000,N_15877,N_15789);
or U16001 (N_16001,N_15824,N_15729);
nand U16002 (N_16002,N_15583,N_15550);
nor U16003 (N_16003,N_15511,N_15698);
nand U16004 (N_16004,N_15983,N_15694);
and U16005 (N_16005,N_15816,N_15915);
or U16006 (N_16006,N_15620,N_15738);
or U16007 (N_16007,N_15935,N_15792);
and U16008 (N_16008,N_15897,N_15604);
nand U16009 (N_16009,N_15701,N_15732);
nand U16010 (N_16010,N_15829,N_15754);
or U16011 (N_16011,N_15838,N_15691);
nand U16012 (N_16012,N_15573,N_15516);
or U16013 (N_16013,N_15735,N_15861);
and U16014 (N_16014,N_15971,N_15921);
nor U16015 (N_16015,N_15966,N_15827);
and U16016 (N_16016,N_15723,N_15941);
xor U16017 (N_16017,N_15630,N_15908);
or U16018 (N_16018,N_15566,N_15993);
or U16019 (N_16019,N_15851,N_15543);
nor U16020 (N_16020,N_15678,N_15902);
nor U16021 (N_16021,N_15769,N_15687);
or U16022 (N_16022,N_15502,N_15844);
and U16023 (N_16023,N_15809,N_15777);
xnor U16024 (N_16024,N_15976,N_15812);
and U16025 (N_16025,N_15509,N_15540);
and U16026 (N_16026,N_15719,N_15549);
and U16027 (N_16027,N_15592,N_15696);
and U16028 (N_16028,N_15906,N_15710);
and U16029 (N_16029,N_15554,N_15841);
and U16030 (N_16030,N_15952,N_15986);
xnor U16031 (N_16031,N_15718,N_15544);
nor U16032 (N_16032,N_15677,N_15807);
nor U16033 (N_16033,N_15736,N_15940);
and U16034 (N_16034,N_15674,N_15531);
and U16035 (N_16035,N_15720,N_15582);
or U16036 (N_16036,N_15779,N_15783);
nor U16037 (N_16037,N_15639,N_15857);
and U16038 (N_16038,N_15995,N_15586);
or U16039 (N_16039,N_15740,N_15875);
and U16040 (N_16040,N_15895,N_15733);
and U16041 (N_16041,N_15842,N_15600);
xor U16042 (N_16042,N_15578,N_15521);
xor U16043 (N_16043,N_15506,N_15541);
nor U16044 (N_16044,N_15793,N_15645);
and U16045 (N_16045,N_15644,N_15852);
or U16046 (N_16046,N_15938,N_15896);
nor U16047 (N_16047,N_15788,N_15859);
nor U16048 (N_16048,N_15653,N_15761);
or U16049 (N_16049,N_15893,N_15886);
and U16050 (N_16050,N_15774,N_15819);
nand U16051 (N_16051,N_15560,N_15797);
nand U16052 (N_16052,N_15538,N_15529);
nand U16053 (N_16053,N_15956,N_15518);
or U16054 (N_16054,N_15655,N_15998);
nand U16055 (N_16055,N_15705,N_15669);
nand U16056 (N_16056,N_15756,N_15659);
nor U16057 (N_16057,N_15688,N_15985);
or U16058 (N_16058,N_15767,N_15929);
nor U16059 (N_16059,N_15730,N_15960);
or U16060 (N_16060,N_15519,N_15876);
or U16061 (N_16061,N_15551,N_15603);
nand U16062 (N_16062,N_15590,N_15682);
or U16063 (N_16063,N_15894,N_15672);
or U16064 (N_16064,N_15978,N_15642);
xor U16065 (N_16065,N_15855,N_15608);
or U16066 (N_16066,N_15662,N_15614);
nand U16067 (N_16067,N_15689,N_15647);
nor U16068 (N_16068,N_15634,N_15597);
xor U16069 (N_16069,N_15900,N_15850);
or U16070 (N_16070,N_15963,N_15778);
or U16071 (N_16071,N_15661,N_15822);
and U16072 (N_16072,N_15843,N_15871);
xor U16073 (N_16073,N_15628,N_15955);
nand U16074 (N_16074,N_15922,N_15626);
xnor U16075 (N_16075,N_15775,N_15625);
nor U16076 (N_16076,N_15890,N_15854);
nor U16077 (N_16077,N_15539,N_15664);
nor U16078 (N_16078,N_15892,N_15536);
or U16079 (N_16079,N_15984,N_15559);
and U16080 (N_16080,N_15982,N_15514);
and U16081 (N_16081,N_15651,N_15638);
or U16082 (N_16082,N_15602,N_15681);
xnor U16083 (N_16083,N_15517,N_15546);
and U16084 (N_16084,N_15680,N_15802);
and U16085 (N_16085,N_15524,N_15865);
nor U16086 (N_16086,N_15507,N_15588);
and U16087 (N_16087,N_15932,N_15618);
xor U16088 (N_16088,N_15530,N_15845);
or U16089 (N_16089,N_15558,N_15598);
or U16090 (N_16090,N_15770,N_15679);
nor U16091 (N_16091,N_15925,N_15716);
nor U16092 (N_16092,N_15866,N_15953);
or U16093 (N_16093,N_15621,N_15808);
nand U16094 (N_16094,N_15790,N_15753);
or U16095 (N_16095,N_15567,N_15747);
or U16096 (N_16096,N_15832,N_15833);
xor U16097 (N_16097,N_15795,N_15874);
nor U16098 (N_16098,N_15725,N_15570);
nand U16099 (N_16099,N_15878,N_15996);
nand U16100 (N_16100,N_15527,N_15772);
and U16101 (N_16101,N_15510,N_15919);
xor U16102 (N_16102,N_15826,N_15799);
and U16103 (N_16103,N_15967,N_15631);
or U16104 (N_16104,N_15746,N_15734);
and U16105 (N_16105,N_15656,N_15739);
nand U16106 (N_16106,N_15860,N_15836);
xor U16107 (N_16107,N_15555,N_15552);
and U16108 (N_16108,N_15849,N_15601);
nand U16109 (N_16109,N_15901,N_15846);
nor U16110 (N_16110,N_15992,N_15891);
nand U16111 (N_16111,N_15609,N_15727);
or U16112 (N_16112,N_15837,N_15883);
or U16113 (N_16113,N_15532,N_15596);
or U16114 (N_16114,N_15942,N_15685);
nand U16115 (N_16115,N_15933,N_15979);
nand U16116 (N_16116,N_15821,N_15830);
and U16117 (N_16117,N_15622,N_15786);
nand U16118 (N_16118,N_15828,N_15899);
and U16119 (N_16119,N_15773,N_15784);
nor U16120 (N_16120,N_15912,N_15806);
nand U16121 (N_16121,N_15646,N_15741);
and U16122 (N_16122,N_15684,N_15801);
and U16123 (N_16123,N_15749,N_15693);
nand U16124 (N_16124,N_15765,N_15632);
and U16125 (N_16125,N_15629,N_15743);
nand U16126 (N_16126,N_15962,N_15699);
xnor U16127 (N_16127,N_15523,N_15528);
or U16128 (N_16128,N_15948,N_15654);
nand U16129 (N_16129,N_15504,N_15839);
and U16130 (N_16130,N_15537,N_15577);
nand U16131 (N_16131,N_15904,N_15553);
and U16132 (N_16132,N_15853,N_15926);
or U16133 (N_16133,N_15800,N_15745);
nand U16134 (N_16134,N_15880,N_15615);
nand U16135 (N_16135,N_15752,N_15562);
xor U16136 (N_16136,N_15525,N_15649);
and U16137 (N_16137,N_15867,N_15804);
nor U16138 (N_16138,N_15835,N_15791);
and U16139 (N_16139,N_15593,N_15611);
nand U16140 (N_16140,N_15889,N_15568);
and U16141 (N_16141,N_15713,N_15755);
nand U16142 (N_16142,N_15671,N_15704);
xnor U16143 (N_16143,N_15556,N_15776);
or U16144 (N_16144,N_15690,N_15569);
and U16145 (N_16145,N_15605,N_15782);
nand U16146 (N_16146,N_15825,N_15658);
or U16147 (N_16147,N_15584,N_15565);
or U16148 (N_16148,N_15903,N_15794);
nand U16149 (N_16149,N_15939,N_15703);
nand U16150 (N_16150,N_15916,N_15771);
and U16151 (N_16151,N_15728,N_15726);
nand U16152 (N_16152,N_15599,N_15905);
nand U16153 (N_16153,N_15616,N_15545);
nand U16154 (N_16154,N_15928,N_15737);
nand U16155 (N_16155,N_15909,N_15633);
or U16156 (N_16156,N_15969,N_15574);
nand U16157 (N_16157,N_15652,N_15945);
nor U16158 (N_16158,N_15872,N_15997);
nor U16159 (N_16159,N_15968,N_15619);
and U16160 (N_16160,N_15760,N_15888);
nand U16161 (N_16161,N_15697,N_15815);
or U16162 (N_16162,N_15557,N_15974);
xnor U16163 (N_16163,N_15766,N_15810);
or U16164 (N_16164,N_15934,N_15627);
nor U16165 (N_16165,N_15898,N_15571);
nand U16166 (N_16166,N_15722,N_15930);
or U16167 (N_16167,N_15623,N_15548);
nor U16168 (N_16168,N_15526,N_15882);
nand U16169 (N_16169,N_15758,N_15561);
nor U16170 (N_16170,N_15575,N_15977);
nand U16171 (N_16171,N_15990,N_15964);
or U16172 (N_16172,N_15987,N_15650);
nor U16173 (N_16173,N_15706,N_15512);
xnor U16174 (N_16174,N_15643,N_15508);
and U16175 (N_16175,N_15763,N_15665);
xnor U16176 (N_16176,N_15831,N_15907);
and U16177 (N_16177,N_15613,N_15959);
or U16178 (N_16178,N_15721,N_15668);
xnor U16179 (N_16179,N_15607,N_15759);
xor U16180 (N_16180,N_15981,N_15803);
or U16181 (N_16181,N_15522,N_15748);
nand U16182 (N_16182,N_15811,N_15576);
nand U16183 (N_16183,N_15814,N_15980);
nand U16184 (N_16184,N_15589,N_15864);
nand U16185 (N_16185,N_15636,N_15666);
nand U16186 (N_16186,N_15683,N_15591);
nor U16187 (N_16187,N_15686,N_15887);
or U16188 (N_16188,N_15920,N_15660);
nand U16189 (N_16189,N_15870,N_15515);
and U16190 (N_16190,N_15823,N_15579);
xnor U16191 (N_16191,N_15834,N_15702);
or U16192 (N_16192,N_15798,N_15606);
nand U16193 (N_16193,N_15675,N_15595);
nor U16194 (N_16194,N_15975,N_15764);
nor U16195 (N_16195,N_15863,N_15780);
or U16196 (N_16196,N_15913,N_15988);
and U16197 (N_16197,N_15768,N_15572);
or U16198 (N_16198,N_15750,N_15881);
and U16199 (N_16199,N_15585,N_15648);
and U16200 (N_16200,N_15994,N_15635);
or U16201 (N_16201,N_15862,N_15717);
nand U16202 (N_16202,N_15762,N_15946);
and U16203 (N_16203,N_15885,N_15873);
xor U16204 (N_16204,N_15917,N_15944);
or U16205 (N_16205,N_15563,N_15847);
and U16206 (N_16206,N_15533,N_15751);
nand U16207 (N_16207,N_15501,N_15817);
nand U16208 (N_16208,N_15923,N_15637);
or U16209 (N_16209,N_15787,N_15840);
or U16210 (N_16210,N_15547,N_15961);
or U16211 (N_16211,N_15924,N_15503);
xnor U16212 (N_16212,N_15958,N_15587);
or U16213 (N_16213,N_15991,N_15520);
or U16214 (N_16214,N_15910,N_15667);
or U16215 (N_16215,N_15731,N_15911);
and U16216 (N_16216,N_15856,N_15973);
or U16217 (N_16217,N_15724,N_15715);
and U16218 (N_16218,N_15640,N_15692);
xnor U16219 (N_16219,N_15954,N_15785);
nand U16220 (N_16220,N_15972,N_15535);
or U16221 (N_16221,N_15868,N_15869);
nand U16222 (N_16222,N_15931,N_15927);
nor U16223 (N_16223,N_15610,N_15580);
nor U16224 (N_16224,N_15612,N_15884);
nand U16225 (N_16225,N_15542,N_15937);
and U16226 (N_16226,N_15500,N_15673);
nand U16227 (N_16227,N_15951,N_15709);
and U16228 (N_16228,N_15663,N_15936);
or U16229 (N_16229,N_15757,N_15564);
nor U16230 (N_16230,N_15848,N_15965);
xnor U16231 (N_16231,N_15714,N_15943);
xor U16232 (N_16232,N_15914,N_15957);
nor U16233 (N_16233,N_15918,N_15989);
or U16234 (N_16234,N_15594,N_15700);
nand U16235 (N_16235,N_15657,N_15947);
nand U16236 (N_16236,N_15970,N_15505);
xnor U16237 (N_16237,N_15879,N_15858);
nand U16238 (N_16238,N_15581,N_15670);
and U16239 (N_16239,N_15813,N_15742);
nand U16240 (N_16240,N_15796,N_15818);
nand U16241 (N_16241,N_15744,N_15999);
nand U16242 (N_16242,N_15676,N_15949);
or U16243 (N_16243,N_15711,N_15641);
and U16244 (N_16244,N_15712,N_15534);
and U16245 (N_16245,N_15513,N_15624);
and U16246 (N_16246,N_15781,N_15708);
or U16247 (N_16247,N_15820,N_15695);
or U16248 (N_16248,N_15707,N_15950);
nand U16249 (N_16249,N_15805,N_15617);
and U16250 (N_16250,N_15727,N_15566);
nand U16251 (N_16251,N_15931,N_15669);
and U16252 (N_16252,N_15858,N_15728);
or U16253 (N_16253,N_15817,N_15546);
and U16254 (N_16254,N_15670,N_15735);
or U16255 (N_16255,N_15824,N_15948);
or U16256 (N_16256,N_15632,N_15799);
nor U16257 (N_16257,N_15678,N_15886);
xnor U16258 (N_16258,N_15781,N_15954);
or U16259 (N_16259,N_15548,N_15848);
nand U16260 (N_16260,N_15529,N_15784);
and U16261 (N_16261,N_15893,N_15672);
or U16262 (N_16262,N_15664,N_15911);
and U16263 (N_16263,N_15571,N_15759);
nand U16264 (N_16264,N_15621,N_15751);
and U16265 (N_16265,N_15583,N_15715);
and U16266 (N_16266,N_15993,N_15755);
nand U16267 (N_16267,N_15759,N_15718);
xor U16268 (N_16268,N_15609,N_15683);
nor U16269 (N_16269,N_15991,N_15961);
or U16270 (N_16270,N_15880,N_15549);
nor U16271 (N_16271,N_15718,N_15751);
nor U16272 (N_16272,N_15855,N_15612);
nand U16273 (N_16273,N_15582,N_15910);
xnor U16274 (N_16274,N_15769,N_15997);
nor U16275 (N_16275,N_15999,N_15656);
nor U16276 (N_16276,N_15989,N_15531);
nor U16277 (N_16277,N_15757,N_15562);
nor U16278 (N_16278,N_15708,N_15754);
nor U16279 (N_16279,N_15695,N_15592);
nand U16280 (N_16280,N_15521,N_15897);
xnor U16281 (N_16281,N_15932,N_15896);
and U16282 (N_16282,N_15731,N_15571);
or U16283 (N_16283,N_15720,N_15608);
or U16284 (N_16284,N_15906,N_15703);
nand U16285 (N_16285,N_15880,N_15538);
or U16286 (N_16286,N_15693,N_15770);
or U16287 (N_16287,N_15989,N_15840);
nand U16288 (N_16288,N_15722,N_15638);
xor U16289 (N_16289,N_15805,N_15528);
or U16290 (N_16290,N_15644,N_15760);
or U16291 (N_16291,N_15736,N_15632);
nor U16292 (N_16292,N_15506,N_15892);
nand U16293 (N_16293,N_15833,N_15670);
and U16294 (N_16294,N_15666,N_15601);
and U16295 (N_16295,N_15846,N_15717);
or U16296 (N_16296,N_15673,N_15649);
nor U16297 (N_16297,N_15940,N_15841);
nor U16298 (N_16298,N_15525,N_15979);
xnor U16299 (N_16299,N_15665,N_15811);
or U16300 (N_16300,N_15675,N_15506);
nor U16301 (N_16301,N_15871,N_15522);
nor U16302 (N_16302,N_15681,N_15572);
nand U16303 (N_16303,N_15732,N_15580);
nand U16304 (N_16304,N_15721,N_15970);
nand U16305 (N_16305,N_15634,N_15908);
nand U16306 (N_16306,N_15694,N_15725);
nor U16307 (N_16307,N_15690,N_15874);
nor U16308 (N_16308,N_15813,N_15585);
nand U16309 (N_16309,N_15522,N_15760);
and U16310 (N_16310,N_15921,N_15861);
or U16311 (N_16311,N_15792,N_15975);
nand U16312 (N_16312,N_15712,N_15697);
nor U16313 (N_16313,N_15505,N_15718);
xor U16314 (N_16314,N_15921,N_15580);
nor U16315 (N_16315,N_15657,N_15506);
or U16316 (N_16316,N_15620,N_15743);
or U16317 (N_16317,N_15798,N_15651);
nor U16318 (N_16318,N_15877,N_15999);
nand U16319 (N_16319,N_15505,N_15827);
nor U16320 (N_16320,N_15846,N_15834);
nand U16321 (N_16321,N_15836,N_15982);
or U16322 (N_16322,N_15982,N_15718);
nor U16323 (N_16323,N_15968,N_15565);
nor U16324 (N_16324,N_15500,N_15519);
and U16325 (N_16325,N_15889,N_15577);
or U16326 (N_16326,N_15924,N_15570);
and U16327 (N_16327,N_15942,N_15834);
nand U16328 (N_16328,N_15586,N_15554);
xnor U16329 (N_16329,N_15528,N_15824);
nand U16330 (N_16330,N_15605,N_15557);
nand U16331 (N_16331,N_15864,N_15820);
nand U16332 (N_16332,N_15651,N_15668);
and U16333 (N_16333,N_15893,N_15816);
xnor U16334 (N_16334,N_15753,N_15729);
nor U16335 (N_16335,N_15640,N_15857);
xor U16336 (N_16336,N_15625,N_15708);
or U16337 (N_16337,N_15582,N_15954);
xnor U16338 (N_16338,N_15703,N_15640);
nand U16339 (N_16339,N_15713,N_15821);
nand U16340 (N_16340,N_15892,N_15914);
xnor U16341 (N_16341,N_15962,N_15961);
or U16342 (N_16342,N_15563,N_15925);
nand U16343 (N_16343,N_15623,N_15560);
and U16344 (N_16344,N_15599,N_15637);
nor U16345 (N_16345,N_15894,N_15849);
xnor U16346 (N_16346,N_15900,N_15677);
nand U16347 (N_16347,N_15624,N_15760);
xor U16348 (N_16348,N_15605,N_15964);
or U16349 (N_16349,N_15679,N_15621);
nand U16350 (N_16350,N_15647,N_15701);
and U16351 (N_16351,N_15875,N_15601);
or U16352 (N_16352,N_15571,N_15981);
xor U16353 (N_16353,N_15592,N_15664);
and U16354 (N_16354,N_15737,N_15832);
nor U16355 (N_16355,N_15989,N_15746);
nand U16356 (N_16356,N_15821,N_15805);
or U16357 (N_16357,N_15937,N_15721);
xnor U16358 (N_16358,N_15973,N_15661);
nor U16359 (N_16359,N_15570,N_15727);
and U16360 (N_16360,N_15638,N_15921);
xnor U16361 (N_16361,N_15552,N_15955);
nand U16362 (N_16362,N_15831,N_15701);
nor U16363 (N_16363,N_15793,N_15998);
and U16364 (N_16364,N_15595,N_15900);
nand U16365 (N_16365,N_15944,N_15737);
nand U16366 (N_16366,N_15910,N_15734);
nand U16367 (N_16367,N_15936,N_15650);
nor U16368 (N_16368,N_15782,N_15975);
and U16369 (N_16369,N_15669,N_15938);
nand U16370 (N_16370,N_15584,N_15889);
or U16371 (N_16371,N_15742,N_15637);
or U16372 (N_16372,N_15842,N_15622);
xor U16373 (N_16373,N_15512,N_15533);
nand U16374 (N_16374,N_15787,N_15581);
nand U16375 (N_16375,N_15992,N_15913);
and U16376 (N_16376,N_15541,N_15816);
nand U16377 (N_16377,N_15563,N_15595);
xnor U16378 (N_16378,N_15601,N_15587);
and U16379 (N_16379,N_15697,N_15853);
nand U16380 (N_16380,N_15675,N_15869);
and U16381 (N_16381,N_15656,N_15520);
and U16382 (N_16382,N_15567,N_15843);
nor U16383 (N_16383,N_15757,N_15532);
xnor U16384 (N_16384,N_15586,N_15521);
nand U16385 (N_16385,N_15682,N_15987);
and U16386 (N_16386,N_15549,N_15962);
and U16387 (N_16387,N_15731,N_15505);
nand U16388 (N_16388,N_15851,N_15790);
nor U16389 (N_16389,N_15894,N_15583);
nand U16390 (N_16390,N_15775,N_15782);
nor U16391 (N_16391,N_15557,N_15990);
and U16392 (N_16392,N_15816,N_15666);
nand U16393 (N_16393,N_15503,N_15529);
or U16394 (N_16394,N_15681,N_15895);
and U16395 (N_16395,N_15959,N_15758);
and U16396 (N_16396,N_15667,N_15577);
nand U16397 (N_16397,N_15928,N_15794);
or U16398 (N_16398,N_15764,N_15806);
nor U16399 (N_16399,N_15868,N_15803);
or U16400 (N_16400,N_15809,N_15801);
or U16401 (N_16401,N_15741,N_15638);
and U16402 (N_16402,N_15687,N_15970);
and U16403 (N_16403,N_15770,N_15617);
and U16404 (N_16404,N_15940,N_15633);
nor U16405 (N_16405,N_15676,N_15992);
or U16406 (N_16406,N_15535,N_15937);
xnor U16407 (N_16407,N_15977,N_15945);
or U16408 (N_16408,N_15673,N_15557);
or U16409 (N_16409,N_15592,N_15577);
nor U16410 (N_16410,N_15920,N_15688);
nand U16411 (N_16411,N_15827,N_15812);
nand U16412 (N_16412,N_15770,N_15726);
xor U16413 (N_16413,N_15540,N_15548);
nand U16414 (N_16414,N_15785,N_15533);
nand U16415 (N_16415,N_15713,N_15759);
and U16416 (N_16416,N_15557,N_15860);
nand U16417 (N_16417,N_15580,N_15814);
nor U16418 (N_16418,N_15809,N_15629);
and U16419 (N_16419,N_15976,N_15656);
or U16420 (N_16420,N_15604,N_15679);
or U16421 (N_16421,N_15630,N_15854);
nand U16422 (N_16422,N_15611,N_15759);
and U16423 (N_16423,N_15843,N_15669);
nand U16424 (N_16424,N_15686,N_15827);
and U16425 (N_16425,N_15708,N_15792);
nor U16426 (N_16426,N_15555,N_15875);
nor U16427 (N_16427,N_15818,N_15929);
nor U16428 (N_16428,N_15845,N_15844);
or U16429 (N_16429,N_15895,N_15534);
and U16430 (N_16430,N_15773,N_15751);
nor U16431 (N_16431,N_15990,N_15516);
and U16432 (N_16432,N_15914,N_15951);
or U16433 (N_16433,N_15732,N_15758);
nand U16434 (N_16434,N_15804,N_15671);
or U16435 (N_16435,N_15512,N_15869);
nor U16436 (N_16436,N_15963,N_15862);
nor U16437 (N_16437,N_15581,N_15543);
nand U16438 (N_16438,N_15678,N_15831);
or U16439 (N_16439,N_15578,N_15611);
nand U16440 (N_16440,N_15666,N_15801);
or U16441 (N_16441,N_15862,N_15677);
or U16442 (N_16442,N_15558,N_15619);
nor U16443 (N_16443,N_15668,N_15500);
xor U16444 (N_16444,N_15703,N_15678);
or U16445 (N_16445,N_15879,N_15807);
or U16446 (N_16446,N_15906,N_15657);
nand U16447 (N_16447,N_15675,N_15580);
nor U16448 (N_16448,N_15997,N_15848);
or U16449 (N_16449,N_15775,N_15596);
or U16450 (N_16450,N_15686,N_15785);
nor U16451 (N_16451,N_15988,N_15732);
and U16452 (N_16452,N_15884,N_15903);
and U16453 (N_16453,N_15751,N_15542);
and U16454 (N_16454,N_15632,N_15873);
nor U16455 (N_16455,N_15930,N_15762);
or U16456 (N_16456,N_15578,N_15522);
or U16457 (N_16457,N_15857,N_15902);
or U16458 (N_16458,N_15831,N_15633);
or U16459 (N_16459,N_15997,N_15903);
nor U16460 (N_16460,N_15708,N_15874);
and U16461 (N_16461,N_15594,N_15735);
and U16462 (N_16462,N_15883,N_15815);
and U16463 (N_16463,N_15860,N_15849);
or U16464 (N_16464,N_15796,N_15919);
nand U16465 (N_16465,N_15782,N_15754);
and U16466 (N_16466,N_15652,N_15747);
and U16467 (N_16467,N_15910,N_15604);
nor U16468 (N_16468,N_15537,N_15851);
xnor U16469 (N_16469,N_15968,N_15924);
xnor U16470 (N_16470,N_15693,N_15702);
and U16471 (N_16471,N_15760,N_15917);
and U16472 (N_16472,N_15973,N_15755);
and U16473 (N_16473,N_15698,N_15506);
nor U16474 (N_16474,N_15513,N_15521);
nor U16475 (N_16475,N_15649,N_15885);
xor U16476 (N_16476,N_15534,N_15739);
nor U16477 (N_16477,N_15568,N_15664);
nor U16478 (N_16478,N_15765,N_15952);
and U16479 (N_16479,N_15732,N_15929);
nand U16480 (N_16480,N_15699,N_15918);
and U16481 (N_16481,N_15823,N_15563);
nor U16482 (N_16482,N_15999,N_15884);
or U16483 (N_16483,N_15934,N_15970);
or U16484 (N_16484,N_15880,N_15535);
or U16485 (N_16485,N_15631,N_15902);
nand U16486 (N_16486,N_15877,N_15890);
nand U16487 (N_16487,N_15808,N_15656);
nand U16488 (N_16488,N_15578,N_15837);
nor U16489 (N_16489,N_15552,N_15572);
nand U16490 (N_16490,N_15831,N_15789);
nor U16491 (N_16491,N_15726,N_15731);
nor U16492 (N_16492,N_15714,N_15615);
nor U16493 (N_16493,N_15774,N_15672);
or U16494 (N_16494,N_15742,N_15588);
nand U16495 (N_16495,N_15650,N_15682);
nand U16496 (N_16496,N_15723,N_15599);
or U16497 (N_16497,N_15836,N_15560);
and U16498 (N_16498,N_15891,N_15686);
and U16499 (N_16499,N_15628,N_15621);
nor U16500 (N_16500,N_16442,N_16007);
or U16501 (N_16501,N_16106,N_16467);
or U16502 (N_16502,N_16371,N_16452);
or U16503 (N_16503,N_16014,N_16482);
and U16504 (N_16504,N_16187,N_16114);
nor U16505 (N_16505,N_16251,N_16330);
nor U16506 (N_16506,N_16107,N_16497);
or U16507 (N_16507,N_16468,N_16432);
or U16508 (N_16508,N_16080,N_16234);
and U16509 (N_16509,N_16450,N_16266);
nand U16510 (N_16510,N_16141,N_16319);
or U16511 (N_16511,N_16382,N_16196);
or U16512 (N_16512,N_16332,N_16439);
and U16513 (N_16513,N_16200,N_16479);
or U16514 (N_16514,N_16124,N_16282);
and U16515 (N_16515,N_16477,N_16147);
or U16516 (N_16516,N_16343,N_16095);
xnor U16517 (N_16517,N_16406,N_16093);
and U16518 (N_16518,N_16454,N_16444);
or U16519 (N_16519,N_16358,N_16088);
and U16520 (N_16520,N_16192,N_16369);
and U16521 (N_16521,N_16013,N_16478);
nor U16522 (N_16522,N_16404,N_16185);
nand U16523 (N_16523,N_16016,N_16020);
nor U16524 (N_16524,N_16203,N_16441);
nor U16525 (N_16525,N_16166,N_16264);
or U16526 (N_16526,N_16487,N_16328);
xnor U16527 (N_16527,N_16181,N_16065);
or U16528 (N_16528,N_16254,N_16492);
or U16529 (N_16529,N_16292,N_16183);
nor U16530 (N_16530,N_16082,N_16041);
and U16531 (N_16531,N_16436,N_16277);
and U16532 (N_16532,N_16311,N_16099);
and U16533 (N_16533,N_16098,N_16296);
nor U16534 (N_16534,N_16211,N_16257);
or U16535 (N_16535,N_16457,N_16462);
nor U16536 (N_16536,N_16310,N_16110);
or U16537 (N_16537,N_16290,N_16085);
xnor U16538 (N_16538,N_16475,N_16393);
and U16539 (N_16539,N_16250,N_16167);
nor U16540 (N_16540,N_16488,N_16092);
nor U16541 (N_16541,N_16179,N_16140);
xor U16542 (N_16542,N_16312,N_16394);
nor U16543 (N_16543,N_16164,N_16347);
and U16544 (N_16544,N_16419,N_16072);
nor U16545 (N_16545,N_16286,N_16491);
nor U16546 (N_16546,N_16224,N_16199);
or U16547 (N_16547,N_16342,N_16238);
or U16548 (N_16548,N_16461,N_16308);
nor U16549 (N_16549,N_16003,N_16142);
nand U16550 (N_16550,N_16077,N_16218);
and U16551 (N_16551,N_16026,N_16418);
nor U16552 (N_16552,N_16484,N_16109);
and U16553 (N_16553,N_16373,N_16175);
nand U16554 (N_16554,N_16425,N_16182);
nand U16555 (N_16555,N_16231,N_16485);
nor U16556 (N_16556,N_16120,N_16096);
nand U16557 (N_16557,N_16268,N_16322);
and U16558 (N_16558,N_16335,N_16431);
xor U16559 (N_16559,N_16407,N_16226);
or U16560 (N_16560,N_16243,N_16232);
or U16561 (N_16561,N_16314,N_16242);
nand U16562 (N_16562,N_16334,N_16102);
and U16563 (N_16563,N_16055,N_16036);
and U16564 (N_16564,N_16469,N_16091);
or U16565 (N_16565,N_16274,N_16409);
and U16566 (N_16566,N_16374,N_16113);
or U16567 (N_16567,N_16030,N_16078);
nand U16568 (N_16568,N_16193,N_16128);
nor U16569 (N_16569,N_16194,N_16202);
xor U16570 (N_16570,N_16354,N_16000);
or U16571 (N_16571,N_16390,N_16435);
or U16572 (N_16572,N_16136,N_16269);
or U16573 (N_16573,N_16453,N_16305);
nor U16574 (N_16574,N_16223,N_16320);
and U16575 (N_16575,N_16248,N_16121);
and U16576 (N_16576,N_16261,N_16051);
nand U16577 (N_16577,N_16372,N_16044);
nand U16578 (N_16578,N_16094,N_16410);
xnor U16579 (N_16579,N_16283,N_16050);
and U16580 (N_16580,N_16337,N_16229);
xnor U16581 (N_16581,N_16321,N_16376);
nor U16582 (N_16582,N_16236,N_16365);
and U16583 (N_16583,N_16151,N_16230);
nor U16584 (N_16584,N_16054,N_16087);
and U16585 (N_16585,N_16380,N_16481);
nor U16586 (N_16586,N_16246,N_16002);
nand U16587 (N_16587,N_16089,N_16493);
nor U16588 (N_16588,N_16081,N_16291);
nor U16589 (N_16589,N_16228,N_16195);
nand U16590 (N_16590,N_16428,N_16127);
or U16591 (N_16591,N_16021,N_16064);
and U16592 (N_16592,N_16103,N_16333);
nor U16593 (N_16593,N_16272,N_16402);
nand U16594 (N_16594,N_16169,N_16275);
or U16595 (N_16595,N_16152,N_16004);
and U16596 (N_16596,N_16253,N_16387);
nand U16597 (N_16597,N_16019,N_16355);
nand U16598 (N_16598,N_16213,N_16135);
and U16599 (N_16599,N_16401,N_16397);
or U16600 (N_16600,N_16008,N_16029);
nor U16601 (N_16601,N_16215,N_16460);
and U16602 (N_16602,N_16448,N_16326);
nand U16603 (N_16603,N_16219,N_16115);
nor U16604 (N_16604,N_16206,N_16160);
and U16605 (N_16605,N_16100,N_16172);
or U16606 (N_16606,N_16349,N_16367);
nand U16607 (N_16607,N_16212,N_16158);
nor U16608 (N_16608,N_16027,N_16023);
xor U16609 (N_16609,N_16139,N_16303);
nand U16610 (N_16610,N_16040,N_16170);
or U16611 (N_16611,N_16341,N_16412);
nand U16612 (N_16612,N_16163,N_16146);
nand U16613 (N_16613,N_16416,N_16244);
or U16614 (N_16614,N_16420,N_16344);
nand U16615 (N_16615,N_16233,N_16010);
nor U16616 (N_16616,N_16317,N_16357);
nand U16617 (N_16617,N_16227,N_16005);
and U16618 (N_16618,N_16383,N_16459);
or U16619 (N_16619,N_16368,N_16071);
nor U16620 (N_16620,N_16047,N_16345);
and U16621 (N_16621,N_16495,N_16309);
nor U16622 (N_16622,N_16255,N_16483);
nor U16623 (N_16623,N_16116,N_16148);
and U16624 (N_16624,N_16473,N_16067);
nor U16625 (N_16625,N_16384,N_16104);
nor U16626 (N_16626,N_16165,N_16249);
nand U16627 (N_16627,N_16413,N_16423);
nor U16628 (N_16628,N_16313,N_16119);
and U16629 (N_16629,N_16370,N_16038);
or U16630 (N_16630,N_16289,N_16417);
or U16631 (N_16631,N_16381,N_16024);
or U16632 (N_16632,N_16262,N_16396);
or U16633 (N_16633,N_16415,N_16329);
and U16634 (N_16634,N_16318,N_16480);
nor U16635 (N_16635,N_16018,N_16084);
nor U16636 (N_16636,N_16033,N_16247);
or U16637 (N_16637,N_16090,N_16034);
and U16638 (N_16638,N_16130,N_16405);
or U16639 (N_16639,N_16363,N_16252);
or U16640 (N_16640,N_16424,N_16063);
or U16641 (N_16641,N_16430,N_16391);
or U16642 (N_16642,N_16111,N_16009);
nand U16643 (N_16643,N_16399,N_16188);
nor U16644 (N_16644,N_16022,N_16466);
nand U16645 (N_16645,N_16346,N_16155);
and U16646 (N_16646,N_16201,N_16075);
nor U16647 (N_16647,N_16276,N_16361);
nor U16648 (N_16648,N_16304,N_16171);
or U16649 (N_16649,N_16101,N_16498);
nand U16650 (N_16650,N_16025,N_16489);
and U16651 (N_16651,N_16039,N_16348);
or U16652 (N_16652,N_16324,N_16364);
nor U16653 (N_16653,N_16267,N_16207);
or U16654 (N_16654,N_16126,N_16434);
nor U16655 (N_16655,N_16429,N_16221);
nor U16656 (N_16656,N_16204,N_16294);
and U16657 (N_16657,N_16131,N_16117);
and U16658 (N_16658,N_16043,N_16392);
nor U16659 (N_16659,N_16438,N_16316);
and U16660 (N_16660,N_16122,N_16145);
or U16661 (N_16661,N_16184,N_16057);
nand U16662 (N_16662,N_16208,N_16083);
nor U16663 (N_16663,N_16012,N_16076);
nand U16664 (N_16664,N_16327,N_16315);
and U16665 (N_16665,N_16217,N_16240);
and U16666 (N_16666,N_16451,N_16049);
nor U16667 (N_16667,N_16132,N_16470);
xnor U16668 (N_16668,N_16499,N_16331);
or U16669 (N_16669,N_16058,N_16225);
nor U16670 (N_16670,N_16061,N_16284);
nor U16671 (N_16671,N_16011,N_16301);
and U16672 (N_16672,N_16069,N_16123);
or U16673 (N_16673,N_16178,N_16377);
nor U16674 (N_16674,N_16271,N_16338);
nand U16675 (N_16675,N_16125,N_16045);
nor U16676 (N_16676,N_16414,N_16474);
nand U16677 (N_16677,N_16285,N_16388);
nand U16678 (N_16678,N_16340,N_16074);
nor U16679 (N_16679,N_16471,N_16028);
or U16680 (N_16680,N_16052,N_16150);
and U16681 (N_16681,N_16359,N_16306);
or U16682 (N_16682,N_16180,N_16398);
xor U16683 (N_16683,N_16437,N_16486);
and U16684 (N_16684,N_16302,N_16389);
nor U16685 (N_16685,N_16362,N_16307);
nand U16686 (N_16686,N_16189,N_16440);
xor U16687 (N_16687,N_16134,N_16385);
or U16688 (N_16688,N_16456,N_16157);
nand U16689 (N_16689,N_16445,N_16042);
xor U16690 (N_16690,N_16360,N_16149);
nand U16691 (N_16691,N_16153,N_16351);
xor U16692 (N_16692,N_16168,N_16053);
or U16693 (N_16693,N_16379,N_16258);
and U16694 (N_16694,N_16186,N_16220);
and U16695 (N_16695,N_16222,N_16006);
and U16696 (N_16696,N_16143,N_16325);
nor U16697 (N_16697,N_16162,N_16263);
and U16698 (N_16698,N_16447,N_16056);
nand U16699 (N_16699,N_16209,N_16298);
nand U16700 (N_16700,N_16032,N_16433);
nor U16701 (N_16701,N_16129,N_16449);
nor U16702 (N_16702,N_16472,N_16464);
nand U16703 (N_16703,N_16299,N_16070);
and U16704 (N_16704,N_16001,N_16017);
nand U16705 (N_16705,N_16494,N_16035);
or U16706 (N_16706,N_16210,N_16476);
nand U16707 (N_16707,N_16048,N_16353);
nor U16708 (N_16708,N_16403,N_16350);
and U16709 (N_16709,N_16118,N_16408);
or U16710 (N_16710,N_16270,N_16293);
nand U16711 (N_16711,N_16237,N_16336);
nand U16712 (N_16712,N_16112,N_16386);
nor U16713 (N_16713,N_16174,N_16133);
nor U16714 (N_16714,N_16059,N_16177);
or U16715 (N_16715,N_16176,N_16241);
and U16716 (N_16716,N_16144,N_16259);
nand U16717 (N_16717,N_16426,N_16281);
xor U16718 (N_16718,N_16490,N_16105);
and U16719 (N_16719,N_16260,N_16287);
nor U16720 (N_16720,N_16073,N_16245);
and U16721 (N_16721,N_16278,N_16356);
nor U16722 (N_16722,N_16173,N_16154);
nand U16723 (N_16723,N_16037,N_16463);
and U16724 (N_16724,N_16455,N_16060);
nand U16725 (N_16725,N_16265,N_16214);
nor U16726 (N_16726,N_16400,N_16079);
or U16727 (N_16727,N_16352,N_16411);
and U16728 (N_16728,N_16323,N_16297);
or U16729 (N_16729,N_16191,N_16239);
xnor U16730 (N_16730,N_16295,N_16279);
xnor U16731 (N_16731,N_16378,N_16097);
and U16732 (N_16732,N_16108,N_16086);
or U16733 (N_16733,N_16375,N_16216);
and U16734 (N_16734,N_16273,N_16339);
and U16735 (N_16735,N_16156,N_16205);
nand U16736 (N_16736,N_16138,N_16137);
nor U16737 (N_16737,N_16427,N_16046);
nor U16738 (N_16738,N_16422,N_16458);
nor U16739 (N_16739,N_16015,N_16395);
xnor U16740 (N_16740,N_16159,N_16280);
nand U16741 (N_16741,N_16198,N_16288);
nor U16742 (N_16742,N_16496,N_16465);
nand U16743 (N_16743,N_16256,N_16161);
nor U16744 (N_16744,N_16366,N_16068);
nor U16745 (N_16745,N_16300,N_16197);
nor U16746 (N_16746,N_16066,N_16062);
and U16747 (N_16747,N_16443,N_16421);
nor U16748 (N_16748,N_16446,N_16235);
and U16749 (N_16749,N_16190,N_16031);
nor U16750 (N_16750,N_16052,N_16139);
nor U16751 (N_16751,N_16073,N_16016);
and U16752 (N_16752,N_16175,N_16336);
and U16753 (N_16753,N_16308,N_16037);
and U16754 (N_16754,N_16284,N_16311);
nor U16755 (N_16755,N_16310,N_16335);
or U16756 (N_16756,N_16042,N_16210);
nor U16757 (N_16757,N_16319,N_16035);
xor U16758 (N_16758,N_16134,N_16497);
nor U16759 (N_16759,N_16308,N_16199);
and U16760 (N_16760,N_16174,N_16458);
nand U16761 (N_16761,N_16026,N_16397);
and U16762 (N_16762,N_16106,N_16249);
or U16763 (N_16763,N_16024,N_16308);
xnor U16764 (N_16764,N_16310,N_16468);
nand U16765 (N_16765,N_16294,N_16304);
or U16766 (N_16766,N_16118,N_16489);
and U16767 (N_16767,N_16014,N_16444);
nand U16768 (N_16768,N_16436,N_16235);
xnor U16769 (N_16769,N_16369,N_16161);
and U16770 (N_16770,N_16196,N_16415);
nor U16771 (N_16771,N_16196,N_16063);
and U16772 (N_16772,N_16143,N_16085);
or U16773 (N_16773,N_16044,N_16032);
nor U16774 (N_16774,N_16497,N_16125);
nor U16775 (N_16775,N_16137,N_16311);
nor U16776 (N_16776,N_16095,N_16306);
and U16777 (N_16777,N_16330,N_16279);
or U16778 (N_16778,N_16390,N_16088);
or U16779 (N_16779,N_16365,N_16129);
or U16780 (N_16780,N_16309,N_16275);
nand U16781 (N_16781,N_16393,N_16148);
or U16782 (N_16782,N_16006,N_16068);
nor U16783 (N_16783,N_16123,N_16124);
nor U16784 (N_16784,N_16151,N_16417);
nand U16785 (N_16785,N_16131,N_16480);
nand U16786 (N_16786,N_16148,N_16154);
nand U16787 (N_16787,N_16499,N_16400);
nor U16788 (N_16788,N_16196,N_16474);
and U16789 (N_16789,N_16180,N_16361);
or U16790 (N_16790,N_16046,N_16293);
nand U16791 (N_16791,N_16315,N_16153);
xor U16792 (N_16792,N_16240,N_16093);
and U16793 (N_16793,N_16332,N_16454);
or U16794 (N_16794,N_16132,N_16051);
and U16795 (N_16795,N_16313,N_16180);
or U16796 (N_16796,N_16419,N_16031);
nand U16797 (N_16797,N_16387,N_16038);
or U16798 (N_16798,N_16356,N_16483);
and U16799 (N_16799,N_16289,N_16249);
xnor U16800 (N_16800,N_16010,N_16408);
or U16801 (N_16801,N_16007,N_16478);
nor U16802 (N_16802,N_16483,N_16372);
or U16803 (N_16803,N_16122,N_16099);
nor U16804 (N_16804,N_16241,N_16122);
and U16805 (N_16805,N_16408,N_16394);
nor U16806 (N_16806,N_16243,N_16355);
or U16807 (N_16807,N_16490,N_16270);
or U16808 (N_16808,N_16473,N_16298);
xor U16809 (N_16809,N_16457,N_16193);
nor U16810 (N_16810,N_16244,N_16465);
nor U16811 (N_16811,N_16041,N_16300);
nand U16812 (N_16812,N_16272,N_16185);
nand U16813 (N_16813,N_16187,N_16117);
xnor U16814 (N_16814,N_16366,N_16309);
nand U16815 (N_16815,N_16414,N_16180);
or U16816 (N_16816,N_16060,N_16141);
nor U16817 (N_16817,N_16009,N_16413);
or U16818 (N_16818,N_16169,N_16010);
nand U16819 (N_16819,N_16458,N_16222);
nor U16820 (N_16820,N_16004,N_16084);
nor U16821 (N_16821,N_16074,N_16246);
and U16822 (N_16822,N_16125,N_16438);
xor U16823 (N_16823,N_16024,N_16117);
and U16824 (N_16824,N_16108,N_16089);
nor U16825 (N_16825,N_16219,N_16334);
nor U16826 (N_16826,N_16209,N_16121);
or U16827 (N_16827,N_16132,N_16337);
nor U16828 (N_16828,N_16174,N_16181);
nor U16829 (N_16829,N_16188,N_16299);
nand U16830 (N_16830,N_16335,N_16445);
nor U16831 (N_16831,N_16199,N_16036);
or U16832 (N_16832,N_16231,N_16472);
and U16833 (N_16833,N_16461,N_16159);
or U16834 (N_16834,N_16208,N_16495);
and U16835 (N_16835,N_16040,N_16222);
nand U16836 (N_16836,N_16282,N_16483);
nand U16837 (N_16837,N_16217,N_16409);
nand U16838 (N_16838,N_16412,N_16283);
nand U16839 (N_16839,N_16207,N_16112);
nor U16840 (N_16840,N_16421,N_16003);
nand U16841 (N_16841,N_16134,N_16123);
and U16842 (N_16842,N_16401,N_16343);
nand U16843 (N_16843,N_16466,N_16326);
nand U16844 (N_16844,N_16318,N_16068);
nand U16845 (N_16845,N_16344,N_16447);
nand U16846 (N_16846,N_16163,N_16342);
nand U16847 (N_16847,N_16094,N_16370);
or U16848 (N_16848,N_16384,N_16140);
or U16849 (N_16849,N_16126,N_16344);
nor U16850 (N_16850,N_16085,N_16434);
xor U16851 (N_16851,N_16279,N_16340);
or U16852 (N_16852,N_16177,N_16338);
nand U16853 (N_16853,N_16026,N_16069);
nor U16854 (N_16854,N_16395,N_16014);
and U16855 (N_16855,N_16067,N_16049);
or U16856 (N_16856,N_16183,N_16398);
and U16857 (N_16857,N_16015,N_16476);
nor U16858 (N_16858,N_16148,N_16433);
nand U16859 (N_16859,N_16260,N_16143);
and U16860 (N_16860,N_16247,N_16081);
nand U16861 (N_16861,N_16088,N_16378);
xnor U16862 (N_16862,N_16381,N_16061);
and U16863 (N_16863,N_16396,N_16328);
or U16864 (N_16864,N_16312,N_16246);
and U16865 (N_16865,N_16298,N_16270);
or U16866 (N_16866,N_16174,N_16382);
and U16867 (N_16867,N_16189,N_16340);
nor U16868 (N_16868,N_16162,N_16327);
and U16869 (N_16869,N_16322,N_16409);
xor U16870 (N_16870,N_16119,N_16341);
nand U16871 (N_16871,N_16213,N_16347);
nor U16872 (N_16872,N_16278,N_16188);
or U16873 (N_16873,N_16247,N_16041);
or U16874 (N_16874,N_16293,N_16331);
or U16875 (N_16875,N_16299,N_16118);
or U16876 (N_16876,N_16166,N_16239);
xnor U16877 (N_16877,N_16399,N_16387);
xor U16878 (N_16878,N_16265,N_16076);
xor U16879 (N_16879,N_16020,N_16209);
or U16880 (N_16880,N_16375,N_16159);
or U16881 (N_16881,N_16399,N_16481);
or U16882 (N_16882,N_16199,N_16413);
or U16883 (N_16883,N_16415,N_16099);
or U16884 (N_16884,N_16004,N_16160);
nand U16885 (N_16885,N_16056,N_16433);
or U16886 (N_16886,N_16251,N_16404);
and U16887 (N_16887,N_16286,N_16300);
or U16888 (N_16888,N_16045,N_16296);
and U16889 (N_16889,N_16408,N_16310);
and U16890 (N_16890,N_16172,N_16339);
and U16891 (N_16891,N_16428,N_16255);
nor U16892 (N_16892,N_16271,N_16076);
or U16893 (N_16893,N_16058,N_16140);
nor U16894 (N_16894,N_16487,N_16470);
or U16895 (N_16895,N_16129,N_16224);
and U16896 (N_16896,N_16275,N_16225);
or U16897 (N_16897,N_16195,N_16463);
nor U16898 (N_16898,N_16098,N_16003);
nand U16899 (N_16899,N_16452,N_16153);
or U16900 (N_16900,N_16432,N_16166);
nand U16901 (N_16901,N_16023,N_16145);
nand U16902 (N_16902,N_16024,N_16268);
and U16903 (N_16903,N_16490,N_16438);
and U16904 (N_16904,N_16238,N_16469);
nand U16905 (N_16905,N_16495,N_16302);
nor U16906 (N_16906,N_16163,N_16479);
and U16907 (N_16907,N_16469,N_16364);
xor U16908 (N_16908,N_16037,N_16400);
nor U16909 (N_16909,N_16259,N_16328);
and U16910 (N_16910,N_16356,N_16469);
and U16911 (N_16911,N_16392,N_16092);
nand U16912 (N_16912,N_16388,N_16295);
nand U16913 (N_16913,N_16288,N_16496);
nand U16914 (N_16914,N_16432,N_16062);
or U16915 (N_16915,N_16020,N_16421);
and U16916 (N_16916,N_16173,N_16191);
xor U16917 (N_16917,N_16106,N_16267);
and U16918 (N_16918,N_16444,N_16141);
nor U16919 (N_16919,N_16156,N_16088);
nand U16920 (N_16920,N_16082,N_16458);
xnor U16921 (N_16921,N_16058,N_16253);
nor U16922 (N_16922,N_16299,N_16090);
nor U16923 (N_16923,N_16402,N_16240);
and U16924 (N_16924,N_16462,N_16108);
nand U16925 (N_16925,N_16062,N_16276);
xnor U16926 (N_16926,N_16226,N_16036);
or U16927 (N_16927,N_16233,N_16329);
and U16928 (N_16928,N_16122,N_16360);
nor U16929 (N_16929,N_16193,N_16257);
xnor U16930 (N_16930,N_16249,N_16027);
or U16931 (N_16931,N_16083,N_16008);
or U16932 (N_16932,N_16328,N_16360);
nor U16933 (N_16933,N_16038,N_16125);
nand U16934 (N_16934,N_16268,N_16248);
or U16935 (N_16935,N_16421,N_16328);
and U16936 (N_16936,N_16102,N_16024);
or U16937 (N_16937,N_16376,N_16141);
nor U16938 (N_16938,N_16094,N_16363);
or U16939 (N_16939,N_16077,N_16351);
nor U16940 (N_16940,N_16040,N_16060);
nand U16941 (N_16941,N_16108,N_16192);
or U16942 (N_16942,N_16067,N_16465);
xor U16943 (N_16943,N_16260,N_16094);
nor U16944 (N_16944,N_16252,N_16056);
and U16945 (N_16945,N_16346,N_16016);
or U16946 (N_16946,N_16332,N_16079);
nor U16947 (N_16947,N_16373,N_16272);
xor U16948 (N_16948,N_16173,N_16461);
or U16949 (N_16949,N_16174,N_16470);
xor U16950 (N_16950,N_16438,N_16287);
nand U16951 (N_16951,N_16156,N_16475);
nor U16952 (N_16952,N_16192,N_16096);
nand U16953 (N_16953,N_16413,N_16483);
and U16954 (N_16954,N_16200,N_16070);
and U16955 (N_16955,N_16150,N_16198);
nor U16956 (N_16956,N_16215,N_16006);
xnor U16957 (N_16957,N_16335,N_16318);
nand U16958 (N_16958,N_16030,N_16000);
nor U16959 (N_16959,N_16252,N_16239);
nand U16960 (N_16960,N_16301,N_16475);
nor U16961 (N_16961,N_16013,N_16405);
and U16962 (N_16962,N_16080,N_16040);
or U16963 (N_16963,N_16469,N_16483);
nand U16964 (N_16964,N_16081,N_16231);
xor U16965 (N_16965,N_16132,N_16079);
nor U16966 (N_16966,N_16095,N_16036);
or U16967 (N_16967,N_16420,N_16105);
and U16968 (N_16968,N_16167,N_16141);
or U16969 (N_16969,N_16140,N_16459);
or U16970 (N_16970,N_16349,N_16342);
and U16971 (N_16971,N_16016,N_16103);
nand U16972 (N_16972,N_16392,N_16402);
and U16973 (N_16973,N_16212,N_16317);
nor U16974 (N_16974,N_16074,N_16195);
nand U16975 (N_16975,N_16039,N_16001);
and U16976 (N_16976,N_16002,N_16258);
and U16977 (N_16977,N_16122,N_16419);
and U16978 (N_16978,N_16474,N_16459);
or U16979 (N_16979,N_16388,N_16163);
and U16980 (N_16980,N_16299,N_16481);
or U16981 (N_16981,N_16212,N_16486);
xnor U16982 (N_16982,N_16458,N_16204);
nor U16983 (N_16983,N_16319,N_16137);
or U16984 (N_16984,N_16411,N_16378);
and U16985 (N_16985,N_16046,N_16000);
or U16986 (N_16986,N_16248,N_16210);
nor U16987 (N_16987,N_16124,N_16378);
or U16988 (N_16988,N_16383,N_16126);
xor U16989 (N_16989,N_16036,N_16086);
xnor U16990 (N_16990,N_16321,N_16218);
nand U16991 (N_16991,N_16220,N_16138);
or U16992 (N_16992,N_16198,N_16381);
and U16993 (N_16993,N_16081,N_16011);
and U16994 (N_16994,N_16121,N_16147);
nor U16995 (N_16995,N_16314,N_16295);
and U16996 (N_16996,N_16449,N_16190);
or U16997 (N_16997,N_16405,N_16471);
xor U16998 (N_16998,N_16433,N_16169);
or U16999 (N_16999,N_16355,N_16408);
nand U17000 (N_17000,N_16791,N_16645);
nand U17001 (N_17001,N_16832,N_16825);
nor U17002 (N_17002,N_16615,N_16844);
or U17003 (N_17003,N_16847,N_16540);
nand U17004 (N_17004,N_16931,N_16974);
nor U17005 (N_17005,N_16788,N_16530);
nor U17006 (N_17006,N_16767,N_16834);
or U17007 (N_17007,N_16848,N_16890);
nand U17008 (N_17008,N_16590,N_16623);
or U17009 (N_17009,N_16517,N_16628);
or U17010 (N_17010,N_16561,N_16732);
and U17011 (N_17011,N_16766,N_16954);
or U17012 (N_17012,N_16915,N_16925);
or U17013 (N_17013,N_16742,N_16529);
nor U17014 (N_17014,N_16755,N_16722);
nand U17015 (N_17015,N_16652,N_16984);
or U17016 (N_17016,N_16938,N_16760);
or U17017 (N_17017,N_16608,N_16700);
nand U17018 (N_17018,N_16690,N_16596);
nand U17019 (N_17019,N_16518,N_16990);
or U17020 (N_17020,N_16793,N_16637);
nor U17021 (N_17021,N_16758,N_16624);
xor U17022 (N_17022,N_16995,N_16924);
and U17023 (N_17023,N_16651,N_16829);
nand U17024 (N_17024,N_16694,N_16704);
nand U17025 (N_17025,N_16600,N_16705);
or U17026 (N_17026,N_16845,N_16908);
or U17027 (N_17027,N_16812,N_16846);
nand U17028 (N_17028,N_16750,N_16692);
and U17029 (N_17029,N_16661,N_16711);
nand U17030 (N_17030,N_16524,N_16911);
or U17031 (N_17031,N_16737,N_16878);
nor U17032 (N_17032,N_16718,N_16798);
or U17033 (N_17033,N_16960,N_16814);
nor U17034 (N_17034,N_16876,N_16958);
nor U17035 (N_17035,N_16653,N_16967);
nand U17036 (N_17036,N_16535,N_16935);
xor U17037 (N_17037,N_16778,N_16708);
and U17038 (N_17038,N_16866,N_16562);
or U17039 (N_17039,N_16827,N_16831);
or U17040 (N_17040,N_16559,N_16780);
nand U17041 (N_17041,N_16949,N_16959);
or U17042 (N_17042,N_16817,N_16862);
or U17043 (N_17043,N_16969,N_16527);
and U17044 (N_17044,N_16823,N_16724);
or U17045 (N_17045,N_16531,N_16882);
and U17046 (N_17046,N_16885,N_16551);
nor U17047 (N_17047,N_16856,N_16622);
and U17048 (N_17048,N_16973,N_16928);
and U17049 (N_17049,N_16859,N_16998);
and U17050 (N_17050,N_16514,N_16723);
nor U17051 (N_17051,N_16500,N_16887);
nor U17052 (N_17052,N_16671,N_16680);
nor U17053 (N_17053,N_16937,N_16821);
and U17054 (N_17054,N_16666,N_16644);
and U17055 (N_17055,N_16604,N_16640);
xor U17056 (N_17056,N_16710,N_16884);
and U17057 (N_17057,N_16765,N_16519);
and U17058 (N_17058,N_16956,N_16630);
nand U17059 (N_17059,N_16678,N_16769);
nand U17060 (N_17060,N_16675,N_16840);
nand U17061 (N_17061,N_16749,N_16759);
nor U17062 (N_17062,N_16532,N_16864);
nand U17063 (N_17063,N_16648,N_16903);
and U17064 (N_17064,N_16735,N_16617);
nor U17065 (N_17065,N_16719,N_16588);
nand U17066 (N_17066,N_16679,N_16507);
nor U17067 (N_17067,N_16695,N_16663);
and U17068 (N_17068,N_16612,N_16819);
nand U17069 (N_17069,N_16634,N_16701);
and U17070 (N_17070,N_16904,N_16923);
nor U17071 (N_17071,N_16883,N_16647);
and U17072 (N_17072,N_16568,N_16809);
nor U17073 (N_17073,N_16510,N_16785);
nand U17074 (N_17074,N_16886,N_16584);
nand U17075 (N_17075,N_16693,N_16968);
xor U17076 (N_17076,N_16738,N_16803);
nor U17077 (N_17077,N_16547,N_16768);
xnor U17078 (N_17078,N_16953,N_16513);
or U17079 (N_17079,N_16771,N_16592);
nor U17080 (N_17080,N_16966,N_16691);
nand U17081 (N_17081,N_16697,N_16997);
or U17082 (N_17082,N_16509,N_16774);
nand U17083 (N_17083,N_16613,N_16930);
xor U17084 (N_17084,N_16806,N_16939);
and U17085 (N_17085,N_16508,N_16669);
nor U17086 (N_17086,N_16786,N_16764);
nand U17087 (N_17087,N_16918,N_16957);
nand U17088 (N_17088,N_16744,N_16539);
nand U17089 (N_17089,N_16979,N_16972);
or U17090 (N_17090,N_16706,N_16970);
and U17091 (N_17091,N_16642,N_16578);
or U17092 (N_17092,N_16621,N_16583);
nand U17093 (N_17093,N_16865,N_16593);
xnor U17094 (N_17094,N_16556,N_16716);
xor U17095 (N_17095,N_16566,N_16567);
and U17096 (N_17096,N_16900,N_16837);
nor U17097 (N_17097,N_16897,N_16792);
and U17098 (N_17098,N_16790,N_16743);
and U17099 (N_17099,N_16901,N_16822);
and U17100 (N_17100,N_16763,N_16881);
nor U17101 (N_17101,N_16895,N_16689);
nor U17102 (N_17102,N_16734,N_16804);
and U17103 (N_17103,N_16504,N_16741);
xor U17104 (N_17104,N_16851,N_16523);
and U17105 (N_17105,N_16730,N_16521);
or U17106 (N_17106,N_16858,N_16824);
and U17107 (N_17107,N_16655,N_16892);
nand U17108 (N_17108,N_16565,N_16947);
or U17109 (N_17109,N_16586,N_16933);
nor U17110 (N_17110,N_16794,N_16975);
or U17111 (N_17111,N_16841,N_16502);
and U17112 (N_17112,N_16552,N_16673);
and U17113 (N_17113,N_16868,N_16989);
or U17114 (N_17114,N_16779,N_16811);
or U17115 (N_17115,N_16951,N_16677);
nand U17116 (N_17116,N_16554,N_16914);
and U17117 (N_17117,N_16601,N_16934);
nand U17118 (N_17118,N_16799,N_16999);
and U17119 (N_17119,N_16713,N_16861);
nand U17120 (N_17120,N_16842,N_16609);
xnor U17121 (N_17121,N_16849,N_16818);
nand U17122 (N_17122,N_16650,N_16776);
and U17123 (N_17123,N_16533,N_16542);
or U17124 (N_17124,N_16891,N_16912);
nor U17125 (N_17125,N_16796,N_16991);
and U17126 (N_17126,N_16838,N_16896);
nand U17127 (N_17127,N_16577,N_16942);
or U17128 (N_17128,N_16667,N_16726);
nor U17129 (N_17129,N_16581,N_16619);
or U17130 (N_17130,N_16994,N_16910);
xor U17131 (N_17131,N_16948,N_16982);
nand U17132 (N_17132,N_16987,N_16573);
xor U17133 (N_17133,N_16641,N_16707);
nor U17134 (N_17134,N_16570,N_16961);
nand U17135 (N_17135,N_16815,N_16550);
nand U17136 (N_17136,N_16620,N_16963);
xnor U17137 (N_17137,N_16952,N_16560);
or U17138 (N_17138,N_16585,N_16731);
or U17139 (N_17139,N_16875,N_16538);
nand U17140 (N_17140,N_16879,N_16522);
or U17141 (N_17141,N_16729,N_16919);
or U17142 (N_17142,N_16926,N_16907);
nor U17143 (N_17143,N_16537,N_16860);
and U17144 (N_17144,N_16712,N_16591);
nand U17145 (N_17145,N_16676,N_16605);
xor U17146 (N_17146,N_16668,N_16672);
or U17147 (N_17147,N_16899,N_16665);
xor U17148 (N_17148,N_16906,N_16872);
or U17149 (N_17149,N_16777,N_16546);
or U17150 (N_17150,N_16558,N_16874);
nor U17151 (N_17151,N_16870,N_16703);
or U17152 (N_17152,N_16674,N_16587);
nand U17153 (N_17153,N_16610,N_16913);
xor U17154 (N_17154,N_16603,N_16955);
or U17155 (N_17155,N_16921,N_16515);
nor U17156 (N_17156,N_16932,N_16501);
nand U17157 (N_17157,N_16770,N_16980);
or U17158 (N_17158,N_16635,N_16625);
xor U17159 (N_17159,N_16629,N_16800);
nor U17160 (N_17160,N_16506,N_16627);
or U17161 (N_17161,N_16852,N_16894);
or U17162 (N_17162,N_16606,N_16977);
and U17163 (N_17163,N_16557,N_16754);
or U17164 (N_17164,N_16761,N_16782);
or U17165 (N_17165,N_16863,N_16772);
nand U17166 (N_17166,N_16720,N_16725);
or U17167 (N_17167,N_16631,N_16922);
or U17168 (N_17168,N_16685,N_16783);
nand U17169 (N_17169,N_16850,N_16686);
and U17170 (N_17170,N_16962,N_16988);
and U17171 (N_17171,N_16830,N_16670);
nand U17172 (N_17172,N_16854,N_16563);
nor U17173 (N_17173,N_16787,N_16664);
and U17174 (N_17174,N_16736,N_16597);
xnor U17175 (N_17175,N_16826,N_16929);
and U17176 (N_17176,N_16503,N_16656);
nand U17177 (N_17177,N_16836,N_16688);
and U17178 (N_17178,N_16553,N_16857);
and U17179 (N_17179,N_16639,N_16867);
xor U17180 (N_17180,N_16985,N_16698);
and U17181 (N_17181,N_16598,N_16512);
nand U17182 (N_17182,N_16992,N_16549);
nor U17183 (N_17183,N_16916,N_16614);
or U17184 (N_17184,N_16602,N_16579);
and U17185 (N_17185,N_16657,N_16816);
or U17186 (N_17186,N_16888,N_16898);
nand U17187 (N_17187,N_16709,N_16589);
nor U17188 (N_17188,N_16681,N_16576);
nor U17189 (N_17189,N_16643,N_16871);
nor U17190 (N_17190,N_16905,N_16797);
nand U17191 (N_17191,N_16752,N_16795);
and U17192 (N_17192,N_16835,N_16802);
nand U17193 (N_17193,N_16715,N_16618);
nand U17194 (N_17194,N_16756,N_16505);
nand U17195 (N_17195,N_16748,N_16807);
and U17196 (N_17196,N_16936,N_16727);
or U17197 (N_17197,N_16682,N_16917);
and U17198 (N_17198,N_16654,N_16594);
nor U17199 (N_17199,N_16543,N_16636);
or U17200 (N_17200,N_16828,N_16976);
nand U17201 (N_17201,N_16784,N_16773);
nand U17202 (N_17202,N_16541,N_16940);
and U17203 (N_17203,N_16889,N_16745);
xor U17204 (N_17204,N_16662,N_16607);
and U17205 (N_17205,N_16632,N_16739);
or U17206 (N_17206,N_16595,N_16544);
nor U17207 (N_17207,N_16696,N_16660);
nor U17208 (N_17208,N_16950,N_16946);
or U17209 (N_17209,N_16611,N_16789);
and U17210 (N_17210,N_16775,N_16580);
or U17211 (N_17211,N_16920,N_16762);
and U17212 (N_17212,N_16909,N_16981);
xnor U17213 (N_17213,N_16927,N_16555);
and U17214 (N_17214,N_16684,N_16525);
nand U17215 (N_17215,N_16880,N_16626);
or U17216 (N_17216,N_16572,N_16893);
nor U17217 (N_17217,N_16575,N_16943);
nor U17218 (N_17218,N_16996,N_16702);
and U17219 (N_17219,N_16746,N_16813);
and U17220 (N_17220,N_16978,N_16599);
xnor U17221 (N_17221,N_16721,N_16569);
and U17222 (N_17222,N_16808,N_16714);
and U17223 (N_17223,N_16728,N_16516);
xor U17224 (N_17224,N_16659,N_16877);
nand U17225 (N_17225,N_16820,N_16964);
nand U17226 (N_17226,N_16717,N_16855);
or U17227 (N_17227,N_16781,N_16574);
nor U17228 (N_17228,N_16571,N_16520);
nand U17229 (N_17229,N_16983,N_16986);
xnor U17230 (N_17230,N_16528,N_16638);
or U17231 (N_17231,N_16941,N_16757);
nor U17232 (N_17232,N_16853,N_16833);
xor U17233 (N_17233,N_16753,N_16805);
nor U17234 (N_17234,N_16747,N_16646);
and U17235 (N_17235,N_16902,N_16740);
nand U17236 (N_17236,N_16873,N_16965);
or U17237 (N_17237,N_16843,N_16683);
or U17238 (N_17238,N_16801,N_16751);
and U17239 (N_17239,N_16548,N_16658);
nand U17240 (N_17240,N_16616,N_16733);
nor U17241 (N_17241,N_16649,N_16810);
and U17242 (N_17242,N_16839,N_16993);
nor U17243 (N_17243,N_16536,N_16511);
or U17244 (N_17244,N_16526,N_16971);
or U17245 (N_17245,N_16687,N_16633);
and U17246 (N_17246,N_16944,N_16545);
nor U17247 (N_17247,N_16699,N_16945);
nor U17248 (N_17248,N_16564,N_16534);
xor U17249 (N_17249,N_16869,N_16582);
nor U17250 (N_17250,N_16514,N_16799);
and U17251 (N_17251,N_16767,N_16657);
nand U17252 (N_17252,N_16947,N_16739);
and U17253 (N_17253,N_16522,N_16875);
nor U17254 (N_17254,N_16820,N_16500);
and U17255 (N_17255,N_16921,N_16778);
or U17256 (N_17256,N_16624,N_16636);
or U17257 (N_17257,N_16579,N_16924);
and U17258 (N_17258,N_16965,N_16833);
nand U17259 (N_17259,N_16993,N_16783);
and U17260 (N_17260,N_16727,N_16940);
xnor U17261 (N_17261,N_16828,N_16697);
nand U17262 (N_17262,N_16806,N_16899);
or U17263 (N_17263,N_16907,N_16832);
and U17264 (N_17264,N_16798,N_16980);
nor U17265 (N_17265,N_16720,N_16582);
nor U17266 (N_17266,N_16621,N_16541);
xnor U17267 (N_17267,N_16885,N_16931);
nand U17268 (N_17268,N_16551,N_16886);
nor U17269 (N_17269,N_16643,N_16717);
xnor U17270 (N_17270,N_16790,N_16853);
nor U17271 (N_17271,N_16718,N_16905);
xor U17272 (N_17272,N_16594,N_16832);
nand U17273 (N_17273,N_16667,N_16542);
and U17274 (N_17274,N_16865,N_16837);
or U17275 (N_17275,N_16620,N_16938);
or U17276 (N_17276,N_16828,N_16544);
nor U17277 (N_17277,N_16526,N_16556);
nor U17278 (N_17278,N_16767,N_16992);
or U17279 (N_17279,N_16525,N_16691);
nor U17280 (N_17280,N_16729,N_16799);
and U17281 (N_17281,N_16530,N_16553);
and U17282 (N_17282,N_16973,N_16652);
and U17283 (N_17283,N_16500,N_16987);
or U17284 (N_17284,N_16542,N_16543);
or U17285 (N_17285,N_16983,N_16534);
nor U17286 (N_17286,N_16579,N_16786);
and U17287 (N_17287,N_16831,N_16868);
and U17288 (N_17288,N_16652,N_16568);
nand U17289 (N_17289,N_16533,N_16951);
or U17290 (N_17290,N_16909,N_16927);
nand U17291 (N_17291,N_16834,N_16822);
nand U17292 (N_17292,N_16832,N_16925);
or U17293 (N_17293,N_16756,N_16946);
and U17294 (N_17294,N_16775,N_16801);
nor U17295 (N_17295,N_16613,N_16699);
nor U17296 (N_17296,N_16901,N_16508);
nand U17297 (N_17297,N_16931,N_16688);
nand U17298 (N_17298,N_16618,N_16985);
or U17299 (N_17299,N_16824,N_16717);
nor U17300 (N_17300,N_16866,N_16591);
nor U17301 (N_17301,N_16831,N_16722);
and U17302 (N_17302,N_16696,N_16599);
nand U17303 (N_17303,N_16837,N_16970);
nor U17304 (N_17304,N_16609,N_16973);
nor U17305 (N_17305,N_16631,N_16994);
xnor U17306 (N_17306,N_16543,N_16892);
nand U17307 (N_17307,N_16925,N_16607);
nor U17308 (N_17308,N_16689,N_16553);
or U17309 (N_17309,N_16720,N_16924);
nand U17310 (N_17310,N_16834,N_16686);
and U17311 (N_17311,N_16863,N_16651);
nor U17312 (N_17312,N_16701,N_16836);
nor U17313 (N_17313,N_16694,N_16636);
and U17314 (N_17314,N_16657,N_16945);
and U17315 (N_17315,N_16561,N_16899);
xor U17316 (N_17316,N_16755,N_16782);
xor U17317 (N_17317,N_16878,N_16512);
xor U17318 (N_17318,N_16977,N_16566);
and U17319 (N_17319,N_16580,N_16860);
nand U17320 (N_17320,N_16985,N_16504);
and U17321 (N_17321,N_16515,N_16887);
nand U17322 (N_17322,N_16994,N_16518);
or U17323 (N_17323,N_16635,N_16801);
and U17324 (N_17324,N_16928,N_16632);
and U17325 (N_17325,N_16640,N_16841);
xnor U17326 (N_17326,N_16850,N_16866);
nor U17327 (N_17327,N_16825,N_16698);
xor U17328 (N_17328,N_16957,N_16793);
nand U17329 (N_17329,N_16711,N_16557);
nand U17330 (N_17330,N_16929,N_16508);
nand U17331 (N_17331,N_16983,N_16816);
and U17332 (N_17332,N_16561,N_16769);
and U17333 (N_17333,N_16729,N_16718);
xor U17334 (N_17334,N_16854,N_16619);
and U17335 (N_17335,N_16605,N_16500);
nor U17336 (N_17336,N_16866,N_16528);
xnor U17337 (N_17337,N_16852,N_16810);
and U17338 (N_17338,N_16939,N_16995);
xnor U17339 (N_17339,N_16850,N_16707);
nor U17340 (N_17340,N_16866,N_16637);
nand U17341 (N_17341,N_16554,N_16959);
nor U17342 (N_17342,N_16978,N_16744);
nand U17343 (N_17343,N_16852,N_16836);
nor U17344 (N_17344,N_16635,N_16736);
nor U17345 (N_17345,N_16507,N_16903);
xor U17346 (N_17346,N_16700,N_16732);
or U17347 (N_17347,N_16990,N_16623);
xor U17348 (N_17348,N_16920,N_16742);
nand U17349 (N_17349,N_16901,N_16955);
nand U17350 (N_17350,N_16573,N_16569);
nor U17351 (N_17351,N_16608,N_16711);
nor U17352 (N_17352,N_16558,N_16580);
nand U17353 (N_17353,N_16659,N_16796);
nor U17354 (N_17354,N_16545,N_16886);
or U17355 (N_17355,N_16664,N_16790);
or U17356 (N_17356,N_16527,N_16561);
or U17357 (N_17357,N_16531,N_16620);
nand U17358 (N_17358,N_16965,N_16963);
xor U17359 (N_17359,N_16573,N_16806);
nor U17360 (N_17360,N_16785,N_16891);
xor U17361 (N_17361,N_16721,N_16983);
xnor U17362 (N_17362,N_16531,N_16750);
and U17363 (N_17363,N_16704,N_16956);
and U17364 (N_17364,N_16908,N_16629);
nor U17365 (N_17365,N_16639,N_16626);
nand U17366 (N_17366,N_16583,N_16728);
nand U17367 (N_17367,N_16560,N_16543);
nand U17368 (N_17368,N_16919,N_16629);
and U17369 (N_17369,N_16873,N_16844);
and U17370 (N_17370,N_16573,N_16872);
nor U17371 (N_17371,N_16503,N_16677);
nand U17372 (N_17372,N_16739,N_16594);
nand U17373 (N_17373,N_16522,N_16865);
xor U17374 (N_17374,N_16517,N_16849);
xor U17375 (N_17375,N_16832,N_16749);
or U17376 (N_17376,N_16820,N_16882);
xnor U17377 (N_17377,N_16871,N_16551);
or U17378 (N_17378,N_16952,N_16709);
and U17379 (N_17379,N_16723,N_16651);
and U17380 (N_17380,N_16823,N_16742);
and U17381 (N_17381,N_16772,N_16977);
nand U17382 (N_17382,N_16702,N_16988);
or U17383 (N_17383,N_16729,N_16856);
nor U17384 (N_17384,N_16771,N_16972);
or U17385 (N_17385,N_16781,N_16563);
or U17386 (N_17386,N_16509,N_16700);
nand U17387 (N_17387,N_16564,N_16945);
xnor U17388 (N_17388,N_16794,N_16647);
nand U17389 (N_17389,N_16785,N_16658);
nand U17390 (N_17390,N_16729,N_16813);
or U17391 (N_17391,N_16585,N_16639);
nor U17392 (N_17392,N_16823,N_16872);
nor U17393 (N_17393,N_16798,N_16702);
or U17394 (N_17394,N_16711,N_16796);
nand U17395 (N_17395,N_16989,N_16806);
and U17396 (N_17396,N_16735,N_16996);
or U17397 (N_17397,N_16933,N_16528);
nand U17398 (N_17398,N_16944,N_16558);
and U17399 (N_17399,N_16722,N_16823);
nand U17400 (N_17400,N_16976,N_16977);
and U17401 (N_17401,N_16958,N_16875);
or U17402 (N_17402,N_16980,N_16706);
nor U17403 (N_17403,N_16913,N_16695);
nand U17404 (N_17404,N_16766,N_16601);
or U17405 (N_17405,N_16795,N_16970);
or U17406 (N_17406,N_16836,N_16568);
nor U17407 (N_17407,N_16969,N_16614);
nand U17408 (N_17408,N_16829,N_16962);
or U17409 (N_17409,N_16910,N_16837);
or U17410 (N_17410,N_16612,N_16656);
xor U17411 (N_17411,N_16530,N_16574);
and U17412 (N_17412,N_16570,N_16993);
and U17413 (N_17413,N_16702,N_16712);
xor U17414 (N_17414,N_16717,N_16581);
or U17415 (N_17415,N_16810,N_16953);
nand U17416 (N_17416,N_16793,N_16913);
nand U17417 (N_17417,N_16645,N_16907);
or U17418 (N_17418,N_16768,N_16792);
nor U17419 (N_17419,N_16594,N_16572);
nor U17420 (N_17420,N_16938,N_16863);
nor U17421 (N_17421,N_16867,N_16792);
and U17422 (N_17422,N_16954,N_16682);
and U17423 (N_17423,N_16891,N_16946);
or U17424 (N_17424,N_16569,N_16611);
nor U17425 (N_17425,N_16563,N_16721);
nand U17426 (N_17426,N_16528,N_16500);
nor U17427 (N_17427,N_16587,N_16997);
nor U17428 (N_17428,N_16533,N_16502);
or U17429 (N_17429,N_16699,N_16859);
nand U17430 (N_17430,N_16966,N_16518);
and U17431 (N_17431,N_16502,N_16659);
or U17432 (N_17432,N_16912,N_16958);
and U17433 (N_17433,N_16551,N_16989);
nand U17434 (N_17434,N_16927,N_16781);
and U17435 (N_17435,N_16934,N_16931);
nand U17436 (N_17436,N_16804,N_16549);
nor U17437 (N_17437,N_16741,N_16732);
and U17438 (N_17438,N_16939,N_16954);
nand U17439 (N_17439,N_16990,N_16725);
nor U17440 (N_17440,N_16960,N_16931);
xor U17441 (N_17441,N_16926,N_16860);
xor U17442 (N_17442,N_16892,N_16730);
nor U17443 (N_17443,N_16910,N_16521);
nor U17444 (N_17444,N_16788,N_16991);
nand U17445 (N_17445,N_16908,N_16910);
nand U17446 (N_17446,N_16794,N_16532);
or U17447 (N_17447,N_16595,N_16760);
nand U17448 (N_17448,N_16777,N_16883);
nor U17449 (N_17449,N_16549,N_16955);
and U17450 (N_17450,N_16764,N_16816);
xor U17451 (N_17451,N_16630,N_16643);
nor U17452 (N_17452,N_16766,N_16938);
nand U17453 (N_17453,N_16676,N_16534);
and U17454 (N_17454,N_16632,N_16562);
and U17455 (N_17455,N_16686,N_16822);
nor U17456 (N_17456,N_16519,N_16923);
nor U17457 (N_17457,N_16988,N_16868);
nor U17458 (N_17458,N_16705,N_16620);
nand U17459 (N_17459,N_16849,N_16832);
nand U17460 (N_17460,N_16885,N_16986);
and U17461 (N_17461,N_16856,N_16847);
and U17462 (N_17462,N_16880,N_16684);
nand U17463 (N_17463,N_16763,N_16697);
and U17464 (N_17464,N_16613,N_16724);
and U17465 (N_17465,N_16794,N_16912);
nor U17466 (N_17466,N_16675,N_16849);
and U17467 (N_17467,N_16512,N_16998);
nor U17468 (N_17468,N_16724,N_16958);
and U17469 (N_17469,N_16548,N_16806);
or U17470 (N_17470,N_16699,N_16518);
or U17471 (N_17471,N_16526,N_16894);
and U17472 (N_17472,N_16710,N_16681);
nor U17473 (N_17473,N_16802,N_16624);
nand U17474 (N_17474,N_16989,N_16837);
nand U17475 (N_17475,N_16575,N_16949);
nor U17476 (N_17476,N_16715,N_16768);
or U17477 (N_17477,N_16568,N_16909);
nor U17478 (N_17478,N_16940,N_16559);
or U17479 (N_17479,N_16570,N_16879);
nand U17480 (N_17480,N_16582,N_16829);
and U17481 (N_17481,N_16771,N_16826);
or U17482 (N_17482,N_16946,N_16531);
nand U17483 (N_17483,N_16791,N_16855);
xnor U17484 (N_17484,N_16530,N_16785);
nor U17485 (N_17485,N_16613,N_16806);
and U17486 (N_17486,N_16638,N_16742);
nand U17487 (N_17487,N_16725,N_16782);
nor U17488 (N_17488,N_16544,N_16846);
nand U17489 (N_17489,N_16577,N_16667);
nand U17490 (N_17490,N_16795,N_16645);
nand U17491 (N_17491,N_16884,N_16673);
nand U17492 (N_17492,N_16588,N_16770);
nand U17493 (N_17493,N_16937,N_16878);
or U17494 (N_17494,N_16964,N_16924);
or U17495 (N_17495,N_16522,N_16514);
or U17496 (N_17496,N_16729,N_16581);
or U17497 (N_17497,N_16641,N_16590);
xnor U17498 (N_17498,N_16566,N_16721);
and U17499 (N_17499,N_16823,N_16515);
nor U17500 (N_17500,N_17256,N_17254);
nor U17501 (N_17501,N_17488,N_17266);
nand U17502 (N_17502,N_17248,N_17195);
nand U17503 (N_17503,N_17281,N_17468);
or U17504 (N_17504,N_17299,N_17024);
nand U17505 (N_17505,N_17217,N_17294);
or U17506 (N_17506,N_17194,N_17017);
nand U17507 (N_17507,N_17291,N_17493);
or U17508 (N_17508,N_17282,N_17404);
xnor U17509 (N_17509,N_17197,N_17381);
nor U17510 (N_17510,N_17022,N_17402);
nor U17511 (N_17511,N_17097,N_17384);
nor U17512 (N_17512,N_17130,N_17094);
nand U17513 (N_17513,N_17239,N_17487);
and U17514 (N_17514,N_17223,N_17079);
nand U17515 (N_17515,N_17001,N_17200);
nor U17516 (N_17516,N_17319,N_17111);
and U17517 (N_17517,N_17374,N_17028);
xnor U17518 (N_17518,N_17152,N_17457);
nand U17519 (N_17519,N_17161,N_17208);
or U17520 (N_17520,N_17421,N_17085);
nand U17521 (N_17521,N_17464,N_17241);
or U17522 (N_17522,N_17221,N_17049);
or U17523 (N_17523,N_17233,N_17175);
nor U17524 (N_17524,N_17155,N_17454);
or U17525 (N_17525,N_17082,N_17312);
nand U17526 (N_17526,N_17234,N_17396);
nand U17527 (N_17527,N_17344,N_17171);
nand U17528 (N_17528,N_17148,N_17490);
and U17529 (N_17529,N_17196,N_17000);
nand U17530 (N_17530,N_17474,N_17096);
nand U17531 (N_17531,N_17475,N_17057);
and U17532 (N_17532,N_17385,N_17352);
nor U17533 (N_17533,N_17495,N_17288);
or U17534 (N_17534,N_17335,N_17411);
nand U17535 (N_17535,N_17304,N_17320);
xor U17536 (N_17536,N_17461,N_17156);
and U17537 (N_17537,N_17446,N_17355);
and U17538 (N_17538,N_17040,N_17103);
or U17539 (N_17539,N_17382,N_17147);
nand U17540 (N_17540,N_17322,N_17203);
nand U17541 (N_17541,N_17192,N_17491);
and U17542 (N_17542,N_17286,N_17367);
xnor U17543 (N_17543,N_17230,N_17153);
nor U17544 (N_17544,N_17188,N_17422);
and U17545 (N_17545,N_17275,N_17357);
xnor U17546 (N_17546,N_17489,N_17013);
xnor U17547 (N_17547,N_17338,N_17328);
nor U17548 (N_17548,N_17370,N_17249);
nand U17549 (N_17549,N_17473,N_17176);
xnor U17550 (N_17550,N_17419,N_17347);
nand U17551 (N_17551,N_17225,N_17455);
nor U17552 (N_17552,N_17467,N_17071);
and U17553 (N_17553,N_17122,N_17073);
or U17554 (N_17554,N_17041,N_17383);
and U17555 (N_17555,N_17441,N_17497);
nor U17556 (N_17556,N_17339,N_17498);
xor U17557 (N_17557,N_17277,N_17180);
or U17558 (N_17558,N_17052,N_17010);
xor U17559 (N_17559,N_17062,N_17460);
xnor U17560 (N_17560,N_17260,N_17465);
or U17561 (N_17561,N_17100,N_17406);
or U17562 (N_17562,N_17169,N_17424);
nor U17563 (N_17563,N_17436,N_17163);
and U17564 (N_17564,N_17222,N_17093);
xnor U17565 (N_17565,N_17456,N_17128);
or U17566 (N_17566,N_17237,N_17226);
or U17567 (N_17567,N_17437,N_17451);
and U17568 (N_17568,N_17420,N_17345);
nor U17569 (N_17569,N_17127,N_17069);
or U17570 (N_17570,N_17269,N_17121);
or U17571 (N_17571,N_17227,N_17447);
or U17572 (N_17572,N_17137,N_17047);
nor U17573 (N_17573,N_17336,N_17481);
or U17574 (N_17574,N_17263,N_17056);
or U17575 (N_17575,N_17343,N_17327);
or U17576 (N_17576,N_17035,N_17334);
nor U17577 (N_17577,N_17238,N_17198);
or U17578 (N_17578,N_17048,N_17264);
nor U17579 (N_17579,N_17025,N_17020);
and U17580 (N_17580,N_17125,N_17141);
or U17581 (N_17581,N_17114,N_17004);
nor U17582 (N_17582,N_17009,N_17305);
nand U17583 (N_17583,N_17469,N_17251);
or U17584 (N_17584,N_17273,N_17438);
or U17585 (N_17585,N_17278,N_17314);
nand U17586 (N_17586,N_17365,N_17313);
nor U17587 (N_17587,N_17330,N_17287);
nor U17588 (N_17588,N_17038,N_17205);
xor U17589 (N_17589,N_17309,N_17340);
and U17590 (N_17590,N_17480,N_17002);
and U17591 (N_17591,N_17409,N_17432);
or U17592 (N_17592,N_17033,N_17204);
nand U17593 (N_17593,N_17311,N_17105);
or U17594 (N_17594,N_17247,N_17202);
or U17595 (N_17595,N_17075,N_17270);
nand U17596 (N_17596,N_17442,N_17417);
nor U17597 (N_17597,N_17037,N_17042);
nand U17598 (N_17598,N_17181,N_17191);
xnor U17599 (N_17599,N_17112,N_17139);
and U17600 (N_17600,N_17354,N_17389);
xnor U17601 (N_17601,N_17246,N_17435);
or U17602 (N_17602,N_17118,N_17290);
and U17603 (N_17603,N_17332,N_17390);
nand U17604 (N_17604,N_17350,N_17220);
or U17605 (N_17605,N_17440,N_17229);
nand U17606 (N_17606,N_17341,N_17280);
or U17607 (N_17607,N_17371,N_17496);
nor U17608 (N_17608,N_17250,N_17391);
xor U17609 (N_17609,N_17261,N_17064);
nand U17610 (N_17610,N_17272,N_17363);
nand U17611 (N_17611,N_17172,N_17008);
nand U17612 (N_17612,N_17209,N_17478);
and U17613 (N_17613,N_17124,N_17236);
or U17614 (N_17614,N_17159,N_17078);
and U17615 (N_17615,N_17329,N_17412);
or U17616 (N_17616,N_17110,N_17154);
or U17617 (N_17617,N_17206,N_17183);
and U17618 (N_17618,N_17072,N_17189);
and U17619 (N_17619,N_17258,N_17193);
or U17620 (N_17620,N_17218,N_17232);
or U17621 (N_17621,N_17321,N_17157);
nand U17622 (N_17622,N_17292,N_17484);
xor U17623 (N_17623,N_17164,N_17166);
xor U17624 (N_17624,N_17045,N_17162);
nand U17625 (N_17625,N_17060,N_17216);
or U17626 (N_17626,N_17207,N_17259);
nand U17627 (N_17627,N_17368,N_17353);
nand U17628 (N_17628,N_17149,N_17333);
and U17629 (N_17629,N_17058,N_17462);
and U17630 (N_17630,N_17360,N_17476);
or U17631 (N_17631,N_17120,N_17362);
and U17632 (N_17632,N_17426,N_17431);
and U17633 (N_17633,N_17021,N_17318);
and U17634 (N_17634,N_17351,N_17300);
and U17635 (N_17635,N_17415,N_17135);
xor U17636 (N_17636,N_17007,N_17032);
or U17637 (N_17637,N_17427,N_17499);
and U17638 (N_17638,N_17143,N_17129);
nor U17639 (N_17639,N_17317,N_17184);
nand U17640 (N_17640,N_17065,N_17265);
nand U17641 (N_17641,N_17190,N_17482);
xnor U17642 (N_17642,N_17109,N_17084);
or U17643 (N_17643,N_17090,N_17483);
and U17644 (N_17644,N_17301,N_17016);
and U17645 (N_17645,N_17276,N_17433);
nand U17646 (N_17646,N_17031,N_17324);
and U17647 (N_17647,N_17228,N_17131);
and U17648 (N_17648,N_17088,N_17036);
and U17649 (N_17649,N_17146,N_17279);
nor U17650 (N_17650,N_17253,N_17342);
and U17651 (N_17651,N_17133,N_17372);
nor U17652 (N_17652,N_17387,N_17182);
or U17653 (N_17653,N_17067,N_17295);
or U17654 (N_17654,N_17395,N_17053);
nand U17655 (N_17655,N_17136,N_17302);
and U17656 (N_17656,N_17403,N_17378);
or U17657 (N_17657,N_17174,N_17243);
and U17658 (N_17658,N_17026,N_17414);
xnor U17659 (N_17659,N_17380,N_17283);
nor U17660 (N_17660,N_17303,N_17293);
nor U17661 (N_17661,N_17087,N_17179);
and U17662 (N_17662,N_17034,N_17108);
and U17663 (N_17663,N_17472,N_17492);
and U17664 (N_17664,N_17224,N_17359);
and U17665 (N_17665,N_17019,N_17018);
nor U17666 (N_17666,N_17095,N_17061);
or U17667 (N_17667,N_17452,N_17219);
and U17668 (N_17668,N_17080,N_17126);
nand U17669 (N_17669,N_17450,N_17443);
and U17670 (N_17670,N_17214,N_17235);
nand U17671 (N_17671,N_17274,N_17086);
or U17672 (N_17672,N_17005,N_17337);
or U17673 (N_17673,N_17150,N_17310);
and U17674 (N_17674,N_17471,N_17083);
or U17675 (N_17675,N_17296,N_17211);
and U17676 (N_17676,N_17123,N_17101);
xor U17677 (N_17677,N_17459,N_17449);
nor U17678 (N_17678,N_17039,N_17413);
and U17679 (N_17679,N_17323,N_17494);
nor U17680 (N_17680,N_17011,N_17348);
and U17681 (N_17681,N_17160,N_17398);
xnor U17682 (N_17682,N_17029,N_17231);
and U17683 (N_17683,N_17187,N_17046);
and U17684 (N_17684,N_17358,N_17479);
and U17685 (N_17685,N_17470,N_17349);
and U17686 (N_17686,N_17307,N_17089);
nor U17687 (N_17687,N_17199,N_17074);
nor U17688 (N_17688,N_17325,N_17113);
or U17689 (N_17689,N_17014,N_17055);
nand U17690 (N_17690,N_17240,N_17375);
and U17691 (N_17691,N_17178,N_17298);
xnor U17692 (N_17692,N_17081,N_17331);
or U17693 (N_17693,N_17267,N_17027);
nand U17694 (N_17694,N_17144,N_17070);
xor U17695 (N_17695,N_17466,N_17405);
and U17696 (N_17696,N_17098,N_17167);
and U17697 (N_17697,N_17059,N_17364);
or U17698 (N_17698,N_17158,N_17444);
nor U17699 (N_17699,N_17284,N_17242);
nand U17700 (N_17700,N_17429,N_17428);
nor U17701 (N_17701,N_17458,N_17445);
or U17702 (N_17702,N_17142,N_17289);
nand U17703 (N_17703,N_17434,N_17271);
xor U17704 (N_17704,N_17115,N_17107);
nand U17705 (N_17705,N_17140,N_17023);
nand U17706 (N_17706,N_17379,N_17003);
or U17707 (N_17707,N_17106,N_17066);
nand U17708 (N_17708,N_17477,N_17377);
nor U17709 (N_17709,N_17346,N_17145);
and U17710 (N_17710,N_17134,N_17297);
nor U17711 (N_17711,N_17268,N_17376);
or U17712 (N_17712,N_17373,N_17186);
and U17713 (N_17713,N_17185,N_17050);
nand U17714 (N_17714,N_17392,N_17044);
or U17715 (N_17715,N_17006,N_17400);
or U17716 (N_17716,N_17117,N_17068);
nor U17717 (N_17717,N_17165,N_17423);
nor U17718 (N_17718,N_17245,N_17453);
nor U17719 (N_17719,N_17104,N_17116);
or U17720 (N_17720,N_17151,N_17244);
or U17721 (N_17721,N_17308,N_17076);
or U17722 (N_17722,N_17257,N_17215);
nor U17723 (N_17723,N_17369,N_17173);
or U17724 (N_17724,N_17397,N_17099);
nand U17725 (N_17725,N_17210,N_17091);
or U17726 (N_17726,N_17386,N_17168);
and U17727 (N_17727,N_17448,N_17485);
or U17728 (N_17728,N_17170,N_17012);
nand U17729 (N_17729,N_17356,N_17262);
xor U17730 (N_17730,N_17138,N_17486);
and U17731 (N_17731,N_17430,N_17054);
nor U17732 (N_17732,N_17407,N_17043);
nor U17733 (N_17733,N_17399,N_17252);
and U17734 (N_17734,N_17394,N_17439);
or U17735 (N_17735,N_17092,N_17361);
or U17736 (N_17736,N_17102,N_17051);
or U17737 (N_17737,N_17119,N_17285);
and U17738 (N_17738,N_17077,N_17326);
nor U17739 (N_17739,N_17408,N_17401);
or U17740 (N_17740,N_17015,N_17416);
nand U17741 (N_17741,N_17463,N_17366);
nand U17742 (N_17742,N_17177,N_17425);
or U17743 (N_17743,N_17410,N_17418);
xnor U17744 (N_17744,N_17393,N_17316);
or U17745 (N_17745,N_17306,N_17063);
xnor U17746 (N_17746,N_17201,N_17132);
nand U17747 (N_17747,N_17030,N_17388);
nand U17748 (N_17748,N_17255,N_17213);
or U17749 (N_17749,N_17212,N_17315);
nand U17750 (N_17750,N_17119,N_17211);
nor U17751 (N_17751,N_17415,N_17462);
xor U17752 (N_17752,N_17088,N_17010);
and U17753 (N_17753,N_17116,N_17138);
nor U17754 (N_17754,N_17160,N_17116);
nor U17755 (N_17755,N_17494,N_17190);
or U17756 (N_17756,N_17219,N_17384);
nor U17757 (N_17757,N_17378,N_17499);
xnor U17758 (N_17758,N_17416,N_17492);
xor U17759 (N_17759,N_17333,N_17339);
and U17760 (N_17760,N_17313,N_17487);
and U17761 (N_17761,N_17415,N_17307);
nand U17762 (N_17762,N_17491,N_17252);
and U17763 (N_17763,N_17218,N_17397);
or U17764 (N_17764,N_17196,N_17041);
nand U17765 (N_17765,N_17290,N_17396);
nor U17766 (N_17766,N_17099,N_17119);
nor U17767 (N_17767,N_17307,N_17424);
nor U17768 (N_17768,N_17016,N_17297);
or U17769 (N_17769,N_17322,N_17120);
nand U17770 (N_17770,N_17460,N_17497);
or U17771 (N_17771,N_17442,N_17293);
nand U17772 (N_17772,N_17270,N_17334);
or U17773 (N_17773,N_17418,N_17462);
and U17774 (N_17774,N_17432,N_17082);
and U17775 (N_17775,N_17426,N_17286);
or U17776 (N_17776,N_17235,N_17242);
nand U17777 (N_17777,N_17113,N_17153);
or U17778 (N_17778,N_17158,N_17455);
or U17779 (N_17779,N_17066,N_17434);
or U17780 (N_17780,N_17262,N_17207);
nand U17781 (N_17781,N_17208,N_17339);
nor U17782 (N_17782,N_17337,N_17368);
and U17783 (N_17783,N_17472,N_17329);
nand U17784 (N_17784,N_17028,N_17432);
and U17785 (N_17785,N_17233,N_17328);
nand U17786 (N_17786,N_17474,N_17495);
nand U17787 (N_17787,N_17436,N_17149);
and U17788 (N_17788,N_17121,N_17385);
nand U17789 (N_17789,N_17263,N_17331);
nand U17790 (N_17790,N_17131,N_17144);
nand U17791 (N_17791,N_17158,N_17124);
nand U17792 (N_17792,N_17410,N_17057);
and U17793 (N_17793,N_17404,N_17474);
nand U17794 (N_17794,N_17076,N_17345);
and U17795 (N_17795,N_17190,N_17131);
or U17796 (N_17796,N_17305,N_17235);
xnor U17797 (N_17797,N_17261,N_17257);
xor U17798 (N_17798,N_17236,N_17323);
nor U17799 (N_17799,N_17496,N_17316);
or U17800 (N_17800,N_17411,N_17367);
or U17801 (N_17801,N_17066,N_17017);
or U17802 (N_17802,N_17337,N_17421);
nand U17803 (N_17803,N_17436,N_17004);
nand U17804 (N_17804,N_17011,N_17490);
and U17805 (N_17805,N_17118,N_17356);
nand U17806 (N_17806,N_17012,N_17112);
nor U17807 (N_17807,N_17388,N_17386);
nor U17808 (N_17808,N_17071,N_17130);
nand U17809 (N_17809,N_17364,N_17164);
nor U17810 (N_17810,N_17235,N_17459);
nor U17811 (N_17811,N_17016,N_17319);
nor U17812 (N_17812,N_17149,N_17319);
or U17813 (N_17813,N_17037,N_17045);
xnor U17814 (N_17814,N_17377,N_17000);
and U17815 (N_17815,N_17026,N_17235);
and U17816 (N_17816,N_17367,N_17114);
or U17817 (N_17817,N_17473,N_17100);
and U17818 (N_17818,N_17170,N_17124);
and U17819 (N_17819,N_17351,N_17128);
nor U17820 (N_17820,N_17001,N_17242);
and U17821 (N_17821,N_17164,N_17222);
and U17822 (N_17822,N_17395,N_17249);
and U17823 (N_17823,N_17349,N_17496);
and U17824 (N_17824,N_17328,N_17356);
or U17825 (N_17825,N_17275,N_17181);
nand U17826 (N_17826,N_17157,N_17458);
or U17827 (N_17827,N_17392,N_17103);
and U17828 (N_17828,N_17137,N_17070);
and U17829 (N_17829,N_17387,N_17221);
nand U17830 (N_17830,N_17480,N_17166);
nand U17831 (N_17831,N_17038,N_17479);
or U17832 (N_17832,N_17276,N_17322);
nand U17833 (N_17833,N_17306,N_17443);
and U17834 (N_17834,N_17354,N_17323);
nand U17835 (N_17835,N_17137,N_17295);
nor U17836 (N_17836,N_17256,N_17224);
nor U17837 (N_17837,N_17487,N_17424);
nor U17838 (N_17838,N_17363,N_17336);
or U17839 (N_17839,N_17123,N_17086);
nor U17840 (N_17840,N_17302,N_17036);
xnor U17841 (N_17841,N_17114,N_17136);
and U17842 (N_17842,N_17041,N_17456);
nand U17843 (N_17843,N_17164,N_17463);
xnor U17844 (N_17844,N_17273,N_17267);
nor U17845 (N_17845,N_17278,N_17072);
or U17846 (N_17846,N_17015,N_17097);
and U17847 (N_17847,N_17457,N_17447);
or U17848 (N_17848,N_17170,N_17049);
and U17849 (N_17849,N_17359,N_17132);
nand U17850 (N_17850,N_17263,N_17497);
xor U17851 (N_17851,N_17471,N_17291);
and U17852 (N_17852,N_17171,N_17462);
or U17853 (N_17853,N_17139,N_17434);
and U17854 (N_17854,N_17401,N_17152);
nor U17855 (N_17855,N_17228,N_17203);
or U17856 (N_17856,N_17423,N_17249);
and U17857 (N_17857,N_17425,N_17158);
nand U17858 (N_17858,N_17179,N_17111);
nor U17859 (N_17859,N_17097,N_17374);
nor U17860 (N_17860,N_17296,N_17266);
or U17861 (N_17861,N_17439,N_17323);
or U17862 (N_17862,N_17009,N_17262);
nand U17863 (N_17863,N_17347,N_17376);
nor U17864 (N_17864,N_17158,N_17005);
nand U17865 (N_17865,N_17398,N_17256);
xnor U17866 (N_17866,N_17006,N_17249);
nor U17867 (N_17867,N_17014,N_17050);
nor U17868 (N_17868,N_17370,N_17017);
nand U17869 (N_17869,N_17329,N_17218);
xor U17870 (N_17870,N_17174,N_17131);
or U17871 (N_17871,N_17067,N_17203);
and U17872 (N_17872,N_17422,N_17465);
or U17873 (N_17873,N_17387,N_17426);
and U17874 (N_17874,N_17390,N_17320);
xnor U17875 (N_17875,N_17250,N_17338);
nand U17876 (N_17876,N_17209,N_17251);
and U17877 (N_17877,N_17088,N_17208);
xnor U17878 (N_17878,N_17287,N_17224);
nand U17879 (N_17879,N_17063,N_17205);
or U17880 (N_17880,N_17448,N_17413);
nor U17881 (N_17881,N_17250,N_17358);
or U17882 (N_17882,N_17441,N_17304);
xnor U17883 (N_17883,N_17468,N_17111);
and U17884 (N_17884,N_17101,N_17096);
nor U17885 (N_17885,N_17308,N_17494);
or U17886 (N_17886,N_17375,N_17106);
or U17887 (N_17887,N_17203,N_17104);
nor U17888 (N_17888,N_17349,N_17146);
nand U17889 (N_17889,N_17221,N_17279);
nand U17890 (N_17890,N_17225,N_17434);
or U17891 (N_17891,N_17106,N_17303);
and U17892 (N_17892,N_17268,N_17016);
and U17893 (N_17893,N_17317,N_17042);
nand U17894 (N_17894,N_17298,N_17305);
or U17895 (N_17895,N_17244,N_17478);
and U17896 (N_17896,N_17379,N_17183);
nor U17897 (N_17897,N_17048,N_17039);
nand U17898 (N_17898,N_17159,N_17342);
nand U17899 (N_17899,N_17217,N_17196);
nand U17900 (N_17900,N_17324,N_17435);
nand U17901 (N_17901,N_17220,N_17068);
or U17902 (N_17902,N_17367,N_17066);
nand U17903 (N_17903,N_17190,N_17485);
nor U17904 (N_17904,N_17204,N_17379);
nor U17905 (N_17905,N_17369,N_17335);
xor U17906 (N_17906,N_17008,N_17489);
nand U17907 (N_17907,N_17426,N_17284);
xnor U17908 (N_17908,N_17317,N_17301);
nand U17909 (N_17909,N_17397,N_17408);
nand U17910 (N_17910,N_17282,N_17024);
and U17911 (N_17911,N_17323,N_17198);
nor U17912 (N_17912,N_17319,N_17112);
nand U17913 (N_17913,N_17357,N_17465);
or U17914 (N_17914,N_17387,N_17068);
or U17915 (N_17915,N_17392,N_17411);
xor U17916 (N_17916,N_17184,N_17408);
nand U17917 (N_17917,N_17281,N_17368);
nor U17918 (N_17918,N_17222,N_17259);
and U17919 (N_17919,N_17099,N_17467);
or U17920 (N_17920,N_17095,N_17070);
or U17921 (N_17921,N_17285,N_17482);
nor U17922 (N_17922,N_17321,N_17480);
xnor U17923 (N_17923,N_17336,N_17392);
and U17924 (N_17924,N_17279,N_17234);
nor U17925 (N_17925,N_17044,N_17118);
nand U17926 (N_17926,N_17258,N_17168);
or U17927 (N_17927,N_17009,N_17278);
nor U17928 (N_17928,N_17008,N_17109);
nor U17929 (N_17929,N_17446,N_17070);
nor U17930 (N_17930,N_17202,N_17020);
and U17931 (N_17931,N_17151,N_17087);
nand U17932 (N_17932,N_17333,N_17355);
or U17933 (N_17933,N_17125,N_17108);
or U17934 (N_17934,N_17016,N_17442);
nand U17935 (N_17935,N_17295,N_17037);
nor U17936 (N_17936,N_17159,N_17291);
nor U17937 (N_17937,N_17157,N_17044);
nor U17938 (N_17938,N_17403,N_17315);
nand U17939 (N_17939,N_17136,N_17223);
or U17940 (N_17940,N_17088,N_17134);
nor U17941 (N_17941,N_17005,N_17025);
nand U17942 (N_17942,N_17165,N_17329);
or U17943 (N_17943,N_17095,N_17047);
xnor U17944 (N_17944,N_17394,N_17100);
nor U17945 (N_17945,N_17044,N_17184);
and U17946 (N_17946,N_17483,N_17277);
xnor U17947 (N_17947,N_17121,N_17216);
or U17948 (N_17948,N_17379,N_17193);
nand U17949 (N_17949,N_17218,N_17471);
xor U17950 (N_17950,N_17429,N_17234);
nand U17951 (N_17951,N_17227,N_17151);
or U17952 (N_17952,N_17486,N_17136);
and U17953 (N_17953,N_17316,N_17476);
or U17954 (N_17954,N_17054,N_17158);
nand U17955 (N_17955,N_17192,N_17372);
xnor U17956 (N_17956,N_17232,N_17272);
and U17957 (N_17957,N_17164,N_17024);
xnor U17958 (N_17958,N_17446,N_17023);
or U17959 (N_17959,N_17461,N_17028);
or U17960 (N_17960,N_17017,N_17011);
nor U17961 (N_17961,N_17290,N_17077);
xor U17962 (N_17962,N_17243,N_17067);
and U17963 (N_17963,N_17280,N_17298);
and U17964 (N_17964,N_17206,N_17471);
or U17965 (N_17965,N_17000,N_17074);
or U17966 (N_17966,N_17219,N_17256);
and U17967 (N_17967,N_17186,N_17047);
nor U17968 (N_17968,N_17308,N_17410);
nand U17969 (N_17969,N_17194,N_17282);
nor U17970 (N_17970,N_17264,N_17384);
nand U17971 (N_17971,N_17278,N_17320);
nand U17972 (N_17972,N_17086,N_17428);
xnor U17973 (N_17973,N_17390,N_17240);
nor U17974 (N_17974,N_17240,N_17144);
and U17975 (N_17975,N_17102,N_17403);
nand U17976 (N_17976,N_17195,N_17403);
and U17977 (N_17977,N_17099,N_17457);
or U17978 (N_17978,N_17381,N_17164);
nor U17979 (N_17979,N_17095,N_17075);
or U17980 (N_17980,N_17455,N_17051);
nand U17981 (N_17981,N_17221,N_17218);
or U17982 (N_17982,N_17137,N_17491);
and U17983 (N_17983,N_17125,N_17309);
and U17984 (N_17984,N_17284,N_17126);
and U17985 (N_17985,N_17093,N_17412);
nand U17986 (N_17986,N_17070,N_17380);
nand U17987 (N_17987,N_17393,N_17277);
nand U17988 (N_17988,N_17262,N_17410);
and U17989 (N_17989,N_17154,N_17025);
nor U17990 (N_17990,N_17498,N_17104);
and U17991 (N_17991,N_17132,N_17063);
nand U17992 (N_17992,N_17499,N_17219);
nand U17993 (N_17993,N_17367,N_17140);
nand U17994 (N_17994,N_17068,N_17190);
xnor U17995 (N_17995,N_17023,N_17345);
xnor U17996 (N_17996,N_17302,N_17492);
or U17997 (N_17997,N_17441,N_17309);
or U17998 (N_17998,N_17425,N_17298);
nand U17999 (N_17999,N_17039,N_17377);
and U18000 (N_18000,N_17625,N_17663);
nor U18001 (N_18001,N_17644,N_17590);
nand U18002 (N_18002,N_17820,N_17516);
or U18003 (N_18003,N_17555,N_17861);
nand U18004 (N_18004,N_17901,N_17731);
nor U18005 (N_18005,N_17802,N_17878);
nor U18006 (N_18006,N_17533,N_17744);
xor U18007 (N_18007,N_17924,N_17956);
nand U18008 (N_18008,N_17853,N_17967);
or U18009 (N_18009,N_17793,N_17636);
nor U18010 (N_18010,N_17952,N_17946);
or U18011 (N_18011,N_17943,N_17609);
xor U18012 (N_18012,N_17991,N_17859);
nand U18013 (N_18013,N_17714,N_17637);
nand U18014 (N_18014,N_17541,N_17762);
nor U18015 (N_18015,N_17912,N_17502);
and U18016 (N_18016,N_17993,N_17870);
xor U18017 (N_18017,N_17873,N_17900);
or U18018 (N_18018,N_17531,N_17990);
nor U18019 (N_18019,N_17825,N_17957);
nand U18020 (N_18020,N_17797,N_17908);
nor U18021 (N_18021,N_17680,N_17737);
and U18022 (N_18022,N_17725,N_17988);
and U18023 (N_18023,N_17501,N_17550);
nor U18024 (N_18024,N_17795,N_17638);
and U18025 (N_18025,N_17986,N_17572);
xnor U18026 (N_18026,N_17969,N_17530);
nor U18027 (N_18027,N_17998,N_17599);
nand U18028 (N_18028,N_17549,N_17951);
and U18029 (N_18029,N_17855,N_17769);
nor U18030 (N_18030,N_17950,N_17829);
or U18031 (N_18031,N_17862,N_17978);
nor U18032 (N_18032,N_17813,N_17819);
nand U18033 (N_18033,N_17573,N_17772);
xor U18034 (N_18034,N_17671,N_17657);
xor U18035 (N_18035,N_17740,N_17529);
nand U18036 (N_18036,N_17904,N_17992);
xnor U18037 (N_18037,N_17911,N_17936);
and U18038 (N_18038,N_17883,N_17561);
and U18039 (N_18039,N_17557,N_17712);
or U18040 (N_18040,N_17713,N_17526);
or U18041 (N_18041,N_17765,N_17849);
and U18042 (N_18042,N_17880,N_17848);
and U18043 (N_18043,N_17733,N_17606);
and U18044 (N_18044,N_17510,N_17705);
nand U18045 (N_18045,N_17521,N_17640);
or U18046 (N_18046,N_17701,N_17886);
or U18047 (N_18047,N_17589,N_17503);
nor U18048 (N_18048,N_17831,N_17796);
and U18049 (N_18049,N_17667,N_17566);
and U18050 (N_18050,N_17570,N_17664);
nor U18051 (N_18051,N_17708,N_17622);
and U18052 (N_18052,N_17665,N_17888);
and U18053 (N_18053,N_17920,N_17730);
or U18054 (N_18054,N_17587,N_17964);
or U18055 (N_18055,N_17546,N_17895);
nand U18056 (N_18056,N_17534,N_17923);
nor U18057 (N_18057,N_17783,N_17841);
and U18058 (N_18058,N_17710,N_17508);
or U18059 (N_18059,N_17605,N_17571);
xor U18060 (N_18060,N_17839,N_17939);
nand U18061 (N_18061,N_17728,N_17868);
nor U18062 (N_18062,N_17887,N_17741);
or U18063 (N_18063,N_17700,N_17683);
and U18064 (N_18064,N_17539,N_17834);
and U18065 (N_18065,N_17961,N_17679);
nand U18066 (N_18066,N_17812,N_17653);
nor U18067 (N_18067,N_17747,N_17630);
and U18068 (N_18068,N_17789,N_17689);
nand U18069 (N_18069,N_17615,N_17997);
or U18070 (N_18070,N_17514,N_17845);
nand U18071 (N_18071,N_17641,N_17832);
nand U18072 (N_18072,N_17734,N_17947);
and U18073 (N_18073,N_17914,N_17984);
nand U18074 (N_18074,N_17953,N_17519);
and U18075 (N_18075,N_17919,N_17786);
and U18076 (N_18076,N_17584,N_17836);
nor U18077 (N_18077,N_17600,N_17660);
and U18078 (N_18078,N_17909,N_17806);
xnor U18079 (N_18079,N_17542,N_17925);
or U18080 (N_18080,N_17575,N_17823);
and U18081 (N_18081,N_17535,N_17882);
and U18082 (N_18082,N_17977,N_17620);
nand U18083 (N_18083,N_17971,N_17751);
nand U18084 (N_18084,N_17881,N_17858);
nand U18085 (N_18085,N_17879,N_17717);
or U18086 (N_18086,N_17522,N_17523);
or U18087 (N_18087,N_17934,N_17596);
and U18088 (N_18088,N_17877,N_17965);
xnor U18089 (N_18089,N_17824,N_17724);
and U18090 (N_18090,N_17702,N_17856);
nand U18091 (N_18091,N_17822,N_17764);
nor U18092 (N_18092,N_17755,N_17774);
or U18093 (N_18093,N_17690,N_17742);
nand U18094 (N_18094,N_17661,N_17897);
nand U18095 (N_18095,N_17975,N_17811);
nand U18096 (N_18096,N_17576,N_17687);
nor U18097 (N_18097,N_17500,N_17669);
nand U18098 (N_18098,N_17757,N_17506);
nor U18099 (N_18099,N_17872,N_17935);
and U18100 (N_18100,N_17982,N_17787);
nor U18101 (N_18101,N_17885,N_17739);
xor U18102 (N_18102,N_17763,N_17659);
nor U18103 (N_18103,N_17838,N_17970);
or U18104 (N_18104,N_17624,N_17748);
nor U18105 (N_18105,N_17634,N_17803);
nor U18106 (N_18106,N_17632,N_17670);
and U18107 (N_18107,N_17685,N_17989);
or U18108 (N_18108,N_17963,N_17835);
nand U18109 (N_18109,N_17960,N_17564);
xor U18110 (N_18110,N_17828,N_17543);
nand U18111 (N_18111,N_17720,N_17581);
or U18112 (N_18112,N_17603,N_17628);
and U18113 (N_18113,N_17554,N_17583);
nand U18114 (N_18114,N_17906,N_17843);
or U18115 (N_18115,N_17654,N_17805);
and U18116 (N_18116,N_17722,N_17941);
or U18117 (N_18117,N_17944,N_17852);
nor U18118 (N_18118,N_17512,N_17794);
or U18119 (N_18119,N_17913,N_17703);
or U18120 (N_18120,N_17721,N_17545);
or U18121 (N_18121,N_17809,N_17651);
or U18122 (N_18122,N_17681,N_17626);
or U18123 (N_18123,N_17693,N_17611);
and U18124 (N_18124,N_17857,N_17821);
or U18125 (N_18125,N_17716,N_17623);
and U18126 (N_18126,N_17699,N_17719);
and U18127 (N_18127,N_17517,N_17610);
and U18128 (N_18128,N_17907,N_17694);
or U18129 (N_18129,N_17696,N_17955);
nand U18130 (N_18130,N_17894,N_17735);
nand U18131 (N_18131,N_17891,N_17771);
nor U18132 (N_18132,N_17921,N_17504);
nor U18133 (N_18133,N_17678,N_17642);
or U18134 (N_18134,N_17846,N_17738);
and U18135 (N_18135,N_17750,N_17954);
nor U18136 (N_18136,N_17892,N_17536);
and U18137 (N_18137,N_17926,N_17827);
or U18138 (N_18138,N_17792,N_17672);
or U18139 (N_18139,N_17760,N_17910);
nand U18140 (N_18140,N_17902,N_17509);
or U18141 (N_18141,N_17585,N_17903);
xnor U18142 (N_18142,N_17544,N_17949);
nor U18143 (N_18143,N_17758,N_17646);
nor U18144 (N_18144,N_17619,N_17867);
nor U18145 (N_18145,N_17966,N_17511);
nor U18146 (N_18146,N_17592,N_17562);
and U18147 (N_18147,N_17752,N_17974);
or U18148 (N_18148,N_17927,N_17602);
nor U18149 (N_18149,N_17692,N_17608);
nand U18150 (N_18150,N_17586,N_17840);
nor U18151 (N_18151,N_17648,N_17565);
or U18152 (N_18152,N_17707,N_17647);
or U18153 (N_18153,N_17513,N_17633);
nand U18154 (N_18154,N_17560,N_17790);
xnor U18155 (N_18155,N_17686,N_17736);
nand U18156 (N_18156,N_17756,N_17652);
or U18157 (N_18157,N_17781,N_17582);
and U18158 (N_18158,N_17767,N_17889);
nand U18159 (N_18159,N_17876,N_17948);
nor U18160 (N_18160,N_17621,N_17874);
nor U18161 (N_18161,N_17675,N_17842);
nand U18162 (N_18162,N_17761,N_17791);
and U18163 (N_18163,N_17658,N_17863);
nor U18164 (N_18164,N_17552,N_17732);
xor U18165 (N_18165,N_17674,N_17726);
nand U18166 (N_18166,N_17847,N_17780);
or U18167 (N_18167,N_17754,N_17649);
nor U18168 (N_18168,N_17807,N_17507);
nand U18169 (N_18169,N_17768,N_17580);
and U18170 (N_18170,N_17559,N_17778);
nand U18171 (N_18171,N_17898,N_17729);
nor U18172 (N_18172,N_17864,N_17505);
or U18173 (N_18173,N_17668,N_17650);
or U18174 (N_18174,N_17677,N_17551);
or U18175 (N_18175,N_17556,N_17817);
nand U18176 (N_18176,N_17577,N_17709);
or U18177 (N_18177,N_17727,N_17558);
or U18178 (N_18178,N_17918,N_17801);
or U18179 (N_18179,N_17759,N_17595);
nor U18180 (N_18180,N_17666,N_17698);
nand U18181 (N_18181,N_17745,N_17588);
and U18182 (N_18182,N_17601,N_17776);
nand U18183 (N_18183,N_17618,N_17704);
nand U18184 (N_18184,N_17553,N_17933);
or U18185 (N_18185,N_17784,N_17981);
or U18186 (N_18186,N_17869,N_17662);
nand U18187 (N_18187,N_17631,N_17833);
xnor U18188 (N_18188,N_17613,N_17890);
nor U18189 (N_18189,N_17958,N_17779);
nand U18190 (N_18190,N_17645,N_17865);
nand U18191 (N_18191,N_17567,N_17808);
nor U18192 (N_18192,N_17917,N_17785);
and U18193 (N_18193,N_17810,N_17749);
and U18194 (N_18194,N_17815,N_17568);
and U18195 (N_18195,N_17655,N_17985);
nor U18196 (N_18196,N_17973,N_17775);
nand U18197 (N_18197,N_17884,N_17816);
nand U18198 (N_18198,N_17799,N_17814);
or U18199 (N_18199,N_17673,N_17537);
nand U18200 (N_18200,N_17940,N_17569);
or U18201 (N_18201,N_17682,N_17715);
or U18202 (N_18202,N_17782,N_17777);
nor U18203 (N_18203,N_17854,N_17937);
and U18204 (N_18204,N_17614,N_17593);
and U18205 (N_18205,N_17612,N_17528);
or U18206 (N_18206,N_17656,N_17607);
nand U18207 (N_18207,N_17695,N_17639);
or U18208 (N_18208,N_17746,N_17540);
nor U18209 (N_18209,N_17627,N_17527);
or U18210 (N_18210,N_17643,N_17938);
and U18211 (N_18211,N_17979,N_17547);
nand U18212 (N_18212,N_17983,N_17987);
nand U18213 (N_18213,N_17995,N_17804);
nand U18214 (N_18214,N_17579,N_17525);
and U18215 (N_18215,N_17930,N_17697);
nand U18216 (N_18216,N_17574,N_17866);
nand U18217 (N_18217,N_17851,N_17893);
nor U18218 (N_18218,N_17837,N_17532);
or U18219 (N_18219,N_17830,N_17800);
xnor U18220 (N_18220,N_17563,N_17896);
nor U18221 (N_18221,N_17922,N_17968);
nand U18222 (N_18222,N_17932,N_17691);
and U18223 (N_18223,N_17711,N_17676);
nor U18224 (N_18224,N_17850,N_17598);
or U18225 (N_18225,N_17520,N_17875);
nand U18226 (N_18226,N_17591,N_17629);
and U18227 (N_18227,N_17548,N_17972);
or U18228 (N_18228,N_17788,N_17980);
nand U18229 (N_18229,N_17905,N_17723);
and U18230 (N_18230,N_17826,N_17616);
nand U18231 (N_18231,N_17798,N_17617);
and U18232 (N_18232,N_17635,N_17994);
or U18233 (N_18233,N_17996,N_17818);
xnor U18234 (N_18234,N_17860,N_17871);
nor U18235 (N_18235,N_17766,N_17844);
nand U18236 (N_18236,N_17597,N_17928);
nor U18237 (N_18237,N_17684,N_17718);
nor U18238 (N_18238,N_17773,N_17688);
nor U18239 (N_18239,N_17604,N_17538);
and U18240 (N_18240,N_17899,N_17976);
nor U18241 (N_18241,N_17594,N_17959);
or U18242 (N_18242,N_17518,N_17915);
nand U18243 (N_18243,N_17770,N_17962);
nand U18244 (N_18244,N_17999,N_17916);
nor U18245 (N_18245,N_17753,N_17515);
nor U18246 (N_18246,N_17931,N_17929);
and U18247 (N_18247,N_17578,N_17706);
nand U18248 (N_18248,N_17942,N_17524);
and U18249 (N_18249,N_17743,N_17945);
or U18250 (N_18250,N_17815,N_17503);
xnor U18251 (N_18251,N_17866,N_17981);
nor U18252 (N_18252,N_17651,N_17646);
nor U18253 (N_18253,N_17615,N_17900);
nor U18254 (N_18254,N_17812,N_17917);
and U18255 (N_18255,N_17781,N_17763);
or U18256 (N_18256,N_17874,N_17962);
xnor U18257 (N_18257,N_17620,N_17811);
or U18258 (N_18258,N_17541,N_17573);
or U18259 (N_18259,N_17566,N_17772);
nand U18260 (N_18260,N_17982,N_17952);
nand U18261 (N_18261,N_17897,N_17677);
and U18262 (N_18262,N_17685,N_17789);
and U18263 (N_18263,N_17574,N_17802);
or U18264 (N_18264,N_17639,N_17986);
nand U18265 (N_18265,N_17594,N_17767);
or U18266 (N_18266,N_17756,N_17903);
xnor U18267 (N_18267,N_17724,N_17673);
and U18268 (N_18268,N_17743,N_17781);
nor U18269 (N_18269,N_17611,N_17516);
or U18270 (N_18270,N_17850,N_17970);
nor U18271 (N_18271,N_17679,N_17925);
nand U18272 (N_18272,N_17862,N_17949);
nand U18273 (N_18273,N_17642,N_17975);
or U18274 (N_18274,N_17938,N_17616);
nor U18275 (N_18275,N_17853,N_17878);
or U18276 (N_18276,N_17576,N_17608);
or U18277 (N_18277,N_17633,N_17735);
nand U18278 (N_18278,N_17829,N_17617);
xnor U18279 (N_18279,N_17969,N_17747);
xnor U18280 (N_18280,N_17925,N_17719);
nand U18281 (N_18281,N_17628,N_17726);
or U18282 (N_18282,N_17571,N_17591);
and U18283 (N_18283,N_17943,N_17949);
xor U18284 (N_18284,N_17823,N_17950);
nand U18285 (N_18285,N_17866,N_17602);
and U18286 (N_18286,N_17853,N_17929);
nor U18287 (N_18287,N_17965,N_17959);
or U18288 (N_18288,N_17702,N_17529);
or U18289 (N_18289,N_17695,N_17791);
nand U18290 (N_18290,N_17656,N_17665);
nand U18291 (N_18291,N_17610,N_17900);
nor U18292 (N_18292,N_17789,N_17802);
and U18293 (N_18293,N_17655,N_17833);
nand U18294 (N_18294,N_17679,N_17602);
nor U18295 (N_18295,N_17643,N_17546);
nand U18296 (N_18296,N_17945,N_17754);
nor U18297 (N_18297,N_17949,N_17872);
or U18298 (N_18298,N_17797,N_17779);
nand U18299 (N_18299,N_17690,N_17922);
nand U18300 (N_18300,N_17791,N_17609);
and U18301 (N_18301,N_17718,N_17826);
and U18302 (N_18302,N_17873,N_17950);
and U18303 (N_18303,N_17615,N_17678);
nand U18304 (N_18304,N_17712,N_17758);
and U18305 (N_18305,N_17862,N_17786);
nor U18306 (N_18306,N_17819,N_17895);
nand U18307 (N_18307,N_17689,N_17919);
or U18308 (N_18308,N_17727,N_17658);
and U18309 (N_18309,N_17740,N_17539);
nor U18310 (N_18310,N_17522,N_17924);
nand U18311 (N_18311,N_17863,N_17898);
nor U18312 (N_18312,N_17533,N_17847);
nand U18313 (N_18313,N_17597,N_17584);
nor U18314 (N_18314,N_17812,N_17909);
nand U18315 (N_18315,N_17728,N_17980);
nand U18316 (N_18316,N_17624,N_17890);
and U18317 (N_18317,N_17793,N_17822);
or U18318 (N_18318,N_17997,N_17611);
and U18319 (N_18319,N_17777,N_17551);
or U18320 (N_18320,N_17794,N_17817);
and U18321 (N_18321,N_17626,N_17931);
nand U18322 (N_18322,N_17691,N_17919);
and U18323 (N_18323,N_17897,N_17911);
xor U18324 (N_18324,N_17524,N_17988);
or U18325 (N_18325,N_17727,N_17635);
xor U18326 (N_18326,N_17651,N_17788);
nand U18327 (N_18327,N_17523,N_17627);
or U18328 (N_18328,N_17511,N_17515);
or U18329 (N_18329,N_17838,N_17987);
or U18330 (N_18330,N_17785,N_17664);
nor U18331 (N_18331,N_17510,N_17953);
nor U18332 (N_18332,N_17584,N_17630);
nor U18333 (N_18333,N_17511,N_17555);
nand U18334 (N_18334,N_17520,N_17775);
and U18335 (N_18335,N_17626,N_17750);
nand U18336 (N_18336,N_17651,N_17767);
or U18337 (N_18337,N_17748,N_17559);
or U18338 (N_18338,N_17785,N_17657);
xnor U18339 (N_18339,N_17838,N_17582);
and U18340 (N_18340,N_17752,N_17785);
and U18341 (N_18341,N_17953,N_17501);
and U18342 (N_18342,N_17507,N_17528);
or U18343 (N_18343,N_17557,N_17732);
nand U18344 (N_18344,N_17961,N_17783);
or U18345 (N_18345,N_17565,N_17817);
or U18346 (N_18346,N_17706,N_17861);
and U18347 (N_18347,N_17984,N_17720);
nand U18348 (N_18348,N_17618,N_17627);
nor U18349 (N_18349,N_17667,N_17542);
and U18350 (N_18350,N_17718,N_17928);
or U18351 (N_18351,N_17764,N_17910);
nand U18352 (N_18352,N_17929,N_17604);
nand U18353 (N_18353,N_17716,N_17966);
or U18354 (N_18354,N_17858,N_17863);
nor U18355 (N_18355,N_17599,N_17891);
xor U18356 (N_18356,N_17579,N_17947);
nor U18357 (N_18357,N_17768,N_17973);
or U18358 (N_18358,N_17704,N_17886);
and U18359 (N_18359,N_17640,N_17883);
or U18360 (N_18360,N_17848,N_17881);
or U18361 (N_18361,N_17819,N_17761);
nand U18362 (N_18362,N_17646,N_17581);
or U18363 (N_18363,N_17735,N_17528);
or U18364 (N_18364,N_17603,N_17589);
and U18365 (N_18365,N_17918,N_17557);
and U18366 (N_18366,N_17539,N_17656);
nand U18367 (N_18367,N_17583,N_17543);
nand U18368 (N_18368,N_17524,N_17949);
or U18369 (N_18369,N_17710,N_17925);
nand U18370 (N_18370,N_17576,N_17948);
nor U18371 (N_18371,N_17812,N_17795);
nand U18372 (N_18372,N_17561,N_17869);
nand U18373 (N_18373,N_17889,N_17982);
and U18374 (N_18374,N_17776,N_17901);
nand U18375 (N_18375,N_17853,N_17579);
or U18376 (N_18376,N_17644,N_17722);
and U18377 (N_18377,N_17517,N_17510);
and U18378 (N_18378,N_17502,N_17678);
nor U18379 (N_18379,N_17814,N_17568);
or U18380 (N_18380,N_17643,N_17812);
nor U18381 (N_18381,N_17654,N_17663);
xnor U18382 (N_18382,N_17853,N_17569);
nor U18383 (N_18383,N_17853,N_17867);
nor U18384 (N_18384,N_17715,N_17790);
nor U18385 (N_18385,N_17549,N_17829);
or U18386 (N_18386,N_17712,N_17781);
and U18387 (N_18387,N_17674,N_17736);
or U18388 (N_18388,N_17827,N_17888);
or U18389 (N_18389,N_17596,N_17642);
or U18390 (N_18390,N_17736,N_17760);
or U18391 (N_18391,N_17589,N_17643);
xor U18392 (N_18392,N_17774,N_17599);
nand U18393 (N_18393,N_17723,N_17701);
and U18394 (N_18394,N_17817,N_17882);
nand U18395 (N_18395,N_17671,N_17855);
or U18396 (N_18396,N_17984,N_17721);
and U18397 (N_18397,N_17786,N_17882);
and U18398 (N_18398,N_17636,N_17876);
nand U18399 (N_18399,N_17933,N_17676);
nand U18400 (N_18400,N_17961,N_17537);
nand U18401 (N_18401,N_17933,N_17545);
or U18402 (N_18402,N_17950,N_17593);
or U18403 (N_18403,N_17860,N_17807);
nor U18404 (N_18404,N_17975,N_17910);
nand U18405 (N_18405,N_17509,N_17601);
xor U18406 (N_18406,N_17959,N_17847);
and U18407 (N_18407,N_17936,N_17957);
or U18408 (N_18408,N_17724,N_17979);
nand U18409 (N_18409,N_17665,N_17639);
nor U18410 (N_18410,N_17599,N_17851);
or U18411 (N_18411,N_17577,N_17604);
nor U18412 (N_18412,N_17968,N_17568);
nand U18413 (N_18413,N_17607,N_17722);
or U18414 (N_18414,N_17784,N_17975);
or U18415 (N_18415,N_17837,N_17829);
or U18416 (N_18416,N_17728,N_17897);
nor U18417 (N_18417,N_17596,N_17534);
or U18418 (N_18418,N_17645,N_17696);
nand U18419 (N_18419,N_17583,N_17882);
and U18420 (N_18420,N_17540,N_17617);
nand U18421 (N_18421,N_17661,N_17584);
xor U18422 (N_18422,N_17875,N_17844);
and U18423 (N_18423,N_17608,N_17728);
nor U18424 (N_18424,N_17752,N_17662);
or U18425 (N_18425,N_17576,N_17940);
and U18426 (N_18426,N_17902,N_17582);
xnor U18427 (N_18427,N_17559,N_17939);
and U18428 (N_18428,N_17585,N_17844);
or U18429 (N_18429,N_17773,N_17991);
and U18430 (N_18430,N_17625,N_17839);
xnor U18431 (N_18431,N_17808,N_17539);
or U18432 (N_18432,N_17702,N_17502);
nor U18433 (N_18433,N_17901,N_17583);
nor U18434 (N_18434,N_17533,N_17912);
or U18435 (N_18435,N_17847,N_17987);
and U18436 (N_18436,N_17704,N_17716);
nand U18437 (N_18437,N_17891,N_17924);
or U18438 (N_18438,N_17603,N_17502);
nand U18439 (N_18439,N_17649,N_17692);
nand U18440 (N_18440,N_17735,N_17846);
and U18441 (N_18441,N_17538,N_17702);
nand U18442 (N_18442,N_17677,N_17610);
xor U18443 (N_18443,N_17892,N_17899);
and U18444 (N_18444,N_17783,N_17906);
nand U18445 (N_18445,N_17691,N_17619);
nor U18446 (N_18446,N_17833,N_17730);
nand U18447 (N_18447,N_17712,N_17894);
nor U18448 (N_18448,N_17936,N_17706);
or U18449 (N_18449,N_17706,N_17994);
and U18450 (N_18450,N_17630,N_17691);
or U18451 (N_18451,N_17514,N_17848);
xor U18452 (N_18452,N_17832,N_17894);
nand U18453 (N_18453,N_17676,N_17632);
nand U18454 (N_18454,N_17758,N_17544);
xor U18455 (N_18455,N_17620,N_17948);
and U18456 (N_18456,N_17662,N_17998);
nand U18457 (N_18457,N_17505,N_17684);
nor U18458 (N_18458,N_17833,N_17819);
and U18459 (N_18459,N_17623,N_17879);
and U18460 (N_18460,N_17703,N_17742);
xor U18461 (N_18461,N_17853,N_17554);
nor U18462 (N_18462,N_17592,N_17742);
xnor U18463 (N_18463,N_17500,N_17830);
nor U18464 (N_18464,N_17902,N_17997);
and U18465 (N_18465,N_17821,N_17734);
nand U18466 (N_18466,N_17992,N_17605);
nor U18467 (N_18467,N_17897,N_17529);
nand U18468 (N_18468,N_17580,N_17520);
and U18469 (N_18469,N_17930,N_17521);
nand U18470 (N_18470,N_17735,N_17784);
or U18471 (N_18471,N_17698,N_17882);
and U18472 (N_18472,N_17863,N_17707);
or U18473 (N_18473,N_17629,N_17812);
or U18474 (N_18474,N_17919,N_17618);
and U18475 (N_18475,N_17550,N_17770);
and U18476 (N_18476,N_17612,N_17500);
or U18477 (N_18477,N_17589,N_17718);
or U18478 (N_18478,N_17919,N_17638);
or U18479 (N_18479,N_17543,N_17841);
or U18480 (N_18480,N_17985,N_17783);
nor U18481 (N_18481,N_17669,N_17934);
xnor U18482 (N_18482,N_17759,N_17807);
or U18483 (N_18483,N_17638,N_17673);
nand U18484 (N_18484,N_17890,N_17554);
nand U18485 (N_18485,N_17644,N_17973);
or U18486 (N_18486,N_17928,N_17793);
or U18487 (N_18487,N_17858,N_17601);
nand U18488 (N_18488,N_17640,N_17740);
or U18489 (N_18489,N_17943,N_17517);
or U18490 (N_18490,N_17585,N_17693);
nor U18491 (N_18491,N_17552,N_17988);
nor U18492 (N_18492,N_17746,N_17826);
or U18493 (N_18493,N_17926,N_17869);
or U18494 (N_18494,N_17954,N_17810);
and U18495 (N_18495,N_17901,N_17648);
nor U18496 (N_18496,N_17577,N_17737);
nor U18497 (N_18497,N_17521,N_17822);
nand U18498 (N_18498,N_17534,N_17511);
or U18499 (N_18499,N_17570,N_17700);
or U18500 (N_18500,N_18222,N_18077);
and U18501 (N_18501,N_18156,N_18125);
nand U18502 (N_18502,N_18417,N_18243);
and U18503 (N_18503,N_18007,N_18045);
or U18504 (N_18504,N_18386,N_18108);
nor U18505 (N_18505,N_18325,N_18395);
nand U18506 (N_18506,N_18389,N_18225);
xor U18507 (N_18507,N_18070,N_18409);
nor U18508 (N_18508,N_18307,N_18174);
nand U18509 (N_18509,N_18401,N_18122);
nand U18510 (N_18510,N_18457,N_18437);
nor U18511 (N_18511,N_18136,N_18178);
nor U18512 (N_18512,N_18373,N_18081);
nor U18513 (N_18513,N_18493,N_18140);
xnor U18514 (N_18514,N_18053,N_18367);
nor U18515 (N_18515,N_18481,N_18141);
nand U18516 (N_18516,N_18004,N_18072);
or U18517 (N_18517,N_18291,N_18458);
nand U18518 (N_18518,N_18476,N_18029);
nand U18519 (N_18519,N_18210,N_18244);
xnor U18520 (N_18520,N_18423,N_18215);
or U18521 (N_18521,N_18357,N_18134);
nor U18522 (N_18522,N_18094,N_18196);
and U18523 (N_18523,N_18245,N_18034);
and U18524 (N_18524,N_18005,N_18013);
nand U18525 (N_18525,N_18428,N_18133);
or U18526 (N_18526,N_18214,N_18202);
or U18527 (N_18527,N_18290,N_18316);
nand U18528 (N_18528,N_18184,N_18314);
and U18529 (N_18529,N_18119,N_18047);
and U18530 (N_18530,N_18265,N_18197);
and U18531 (N_18531,N_18015,N_18181);
nand U18532 (N_18532,N_18380,N_18361);
and U18533 (N_18533,N_18445,N_18486);
or U18534 (N_18534,N_18342,N_18092);
and U18535 (N_18535,N_18432,N_18326);
nand U18536 (N_18536,N_18293,N_18149);
nand U18537 (N_18537,N_18393,N_18399);
and U18538 (N_18538,N_18418,N_18376);
nand U18539 (N_18539,N_18180,N_18213);
nor U18540 (N_18540,N_18071,N_18339);
or U18541 (N_18541,N_18026,N_18407);
nor U18542 (N_18542,N_18038,N_18426);
nand U18543 (N_18543,N_18377,N_18456);
or U18544 (N_18544,N_18074,N_18043);
or U18545 (N_18545,N_18335,N_18260);
and U18546 (N_18546,N_18287,N_18429);
xor U18547 (N_18547,N_18443,N_18487);
nor U18548 (N_18548,N_18114,N_18374);
or U18549 (N_18549,N_18079,N_18421);
nor U18550 (N_18550,N_18115,N_18207);
nor U18551 (N_18551,N_18472,N_18468);
or U18552 (N_18552,N_18152,N_18471);
and U18553 (N_18553,N_18254,N_18451);
nand U18554 (N_18554,N_18059,N_18169);
nor U18555 (N_18555,N_18259,N_18246);
xnor U18556 (N_18556,N_18263,N_18262);
and U18557 (N_18557,N_18276,N_18075);
or U18558 (N_18558,N_18289,N_18479);
or U18559 (N_18559,N_18391,N_18102);
nor U18560 (N_18560,N_18192,N_18086);
nor U18561 (N_18561,N_18322,N_18396);
or U18562 (N_18562,N_18195,N_18057);
or U18563 (N_18563,N_18371,N_18462);
nand U18564 (N_18564,N_18039,N_18150);
and U18565 (N_18565,N_18235,N_18296);
nor U18566 (N_18566,N_18278,N_18261);
and U18567 (N_18567,N_18483,N_18121);
nor U18568 (N_18568,N_18362,N_18248);
nand U18569 (N_18569,N_18310,N_18475);
or U18570 (N_18570,N_18239,N_18069);
nand U18571 (N_18571,N_18292,N_18251);
and U18572 (N_18572,N_18336,N_18329);
nor U18573 (N_18573,N_18110,N_18242);
nor U18574 (N_18574,N_18284,N_18058);
nand U18575 (N_18575,N_18153,N_18040);
nand U18576 (N_18576,N_18282,N_18365);
nor U18577 (N_18577,N_18408,N_18320);
xnor U18578 (N_18578,N_18436,N_18406);
nand U18579 (N_18579,N_18008,N_18498);
and U18580 (N_18580,N_18105,N_18160);
nor U18581 (N_18581,N_18027,N_18341);
nor U18582 (N_18582,N_18454,N_18355);
nor U18583 (N_18583,N_18145,N_18104);
nor U18584 (N_18584,N_18354,N_18302);
nor U18585 (N_18585,N_18411,N_18098);
and U18586 (N_18586,N_18269,N_18494);
nor U18587 (N_18587,N_18394,N_18252);
nor U18588 (N_18588,N_18025,N_18020);
and U18589 (N_18589,N_18161,N_18188);
or U18590 (N_18590,N_18297,N_18450);
or U18591 (N_18591,N_18050,N_18489);
or U18592 (N_18592,N_18328,N_18400);
and U18593 (N_18593,N_18147,N_18019);
nand U18594 (N_18594,N_18440,N_18130);
nand U18595 (N_18595,N_18124,N_18324);
and U18596 (N_18596,N_18138,N_18205);
nor U18597 (N_18597,N_18186,N_18334);
nand U18598 (N_18598,N_18093,N_18203);
and U18599 (N_18599,N_18037,N_18496);
nand U18600 (N_18600,N_18378,N_18018);
nor U18601 (N_18601,N_18435,N_18273);
xnor U18602 (N_18602,N_18191,N_18023);
nand U18603 (N_18603,N_18173,N_18204);
nor U18604 (N_18604,N_18461,N_18158);
or U18605 (N_18605,N_18370,N_18000);
or U18606 (N_18606,N_18459,N_18277);
and U18607 (N_18607,N_18288,N_18414);
and U18608 (N_18608,N_18390,N_18463);
and U18609 (N_18609,N_18255,N_18103);
xor U18610 (N_18610,N_18484,N_18315);
nand U18611 (N_18611,N_18240,N_18460);
xnor U18612 (N_18612,N_18379,N_18311);
nand U18613 (N_18613,N_18340,N_18002);
and U18614 (N_18614,N_18280,N_18331);
or U18615 (N_18615,N_18030,N_18123);
and U18616 (N_18616,N_18490,N_18249);
or U18617 (N_18617,N_18247,N_18274);
or U18618 (N_18618,N_18358,N_18190);
nor U18619 (N_18619,N_18480,N_18258);
or U18620 (N_18620,N_18267,N_18430);
nor U18621 (N_18621,N_18351,N_18106);
and U18622 (N_18622,N_18434,N_18073);
xnor U18623 (N_18623,N_18182,N_18285);
and U18624 (N_18624,N_18343,N_18305);
or U18625 (N_18625,N_18356,N_18157);
nor U18626 (N_18626,N_18209,N_18323);
nor U18627 (N_18627,N_18368,N_18301);
or U18628 (N_18628,N_18091,N_18135);
nand U18629 (N_18629,N_18131,N_18142);
nor U18630 (N_18630,N_18206,N_18216);
and U18631 (N_18631,N_18308,N_18028);
nor U18632 (N_18632,N_18499,N_18303);
nor U18633 (N_18633,N_18228,N_18366);
nor U18634 (N_18634,N_18063,N_18067);
nor U18635 (N_18635,N_18482,N_18201);
and U18636 (N_18636,N_18198,N_18449);
xor U18637 (N_18637,N_18491,N_18080);
and U18638 (N_18638,N_18236,N_18473);
and U18639 (N_18639,N_18447,N_18384);
nand U18640 (N_18640,N_18497,N_18031);
and U18641 (N_18641,N_18346,N_18052);
nand U18642 (N_18642,N_18139,N_18372);
or U18643 (N_18643,N_18233,N_18185);
xor U18644 (N_18644,N_18097,N_18253);
nor U18645 (N_18645,N_18041,N_18272);
nand U18646 (N_18646,N_18218,N_18151);
or U18647 (N_18647,N_18381,N_18387);
or U18648 (N_18648,N_18083,N_18410);
nand U18649 (N_18649,N_18452,N_18194);
and U18650 (N_18650,N_18068,N_18232);
nor U18651 (N_18651,N_18076,N_18404);
nor U18652 (N_18652,N_18109,N_18444);
nor U18653 (N_18653,N_18003,N_18044);
nor U18654 (N_18654,N_18359,N_18264);
xor U18655 (N_18655,N_18229,N_18128);
or U18656 (N_18656,N_18046,N_18474);
nor U18657 (N_18657,N_18234,N_18446);
xor U18658 (N_18658,N_18238,N_18084);
nor U18659 (N_18659,N_18441,N_18318);
and U18660 (N_18660,N_18392,N_18159);
or U18661 (N_18661,N_18085,N_18143);
nor U18662 (N_18662,N_18369,N_18148);
and U18663 (N_18663,N_18189,N_18171);
xnor U18664 (N_18664,N_18100,N_18127);
nand U18665 (N_18665,N_18011,N_18398);
or U18666 (N_18666,N_18144,N_18212);
xor U18667 (N_18667,N_18382,N_18012);
and U18668 (N_18668,N_18137,N_18364);
and U18669 (N_18669,N_18363,N_18049);
nand U18670 (N_18670,N_18167,N_18065);
or U18671 (N_18671,N_18061,N_18425);
nand U18672 (N_18672,N_18337,N_18360);
nand U18673 (N_18673,N_18464,N_18485);
and U18674 (N_18674,N_18107,N_18146);
or U18675 (N_18675,N_18170,N_18298);
xnor U18676 (N_18676,N_18082,N_18162);
and U18677 (N_18677,N_18101,N_18448);
nor U18678 (N_18678,N_18442,N_18319);
or U18679 (N_18679,N_18056,N_18317);
nand U18680 (N_18680,N_18313,N_18295);
nor U18681 (N_18681,N_18266,N_18010);
and U18682 (N_18682,N_18397,N_18154);
and U18683 (N_18683,N_18090,N_18347);
or U18684 (N_18684,N_18415,N_18453);
nand U18685 (N_18685,N_18227,N_18226);
nand U18686 (N_18686,N_18022,N_18163);
and U18687 (N_18687,N_18433,N_18286);
nor U18688 (N_18688,N_18330,N_18168);
nand U18689 (N_18689,N_18111,N_18055);
and U18690 (N_18690,N_18164,N_18304);
nand U18691 (N_18691,N_18193,N_18348);
or U18692 (N_18692,N_18383,N_18279);
and U18693 (N_18693,N_18208,N_18021);
or U18694 (N_18694,N_18126,N_18118);
nand U18695 (N_18695,N_18035,N_18024);
xnor U18696 (N_18696,N_18385,N_18439);
and U18697 (N_18697,N_18350,N_18113);
nand U18698 (N_18698,N_18132,N_18062);
nand U18699 (N_18699,N_18175,N_18333);
nand U18700 (N_18700,N_18495,N_18353);
nand U18701 (N_18701,N_18223,N_18299);
nand U18702 (N_18702,N_18492,N_18467);
and U18703 (N_18703,N_18155,N_18177);
nor U18704 (N_18704,N_18051,N_18230);
and U18705 (N_18705,N_18017,N_18042);
nand U18706 (N_18706,N_18413,N_18183);
or U18707 (N_18707,N_18416,N_18419);
nand U18708 (N_18708,N_18089,N_18172);
or U18709 (N_18709,N_18231,N_18217);
nand U18710 (N_18710,N_18033,N_18469);
nor U18711 (N_18711,N_18117,N_18332);
nor U18712 (N_18712,N_18096,N_18219);
or U18713 (N_18713,N_18420,N_18345);
xor U18714 (N_18714,N_18422,N_18488);
and U18715 (N_18715,N_18087,N_18327);
or U18716 (N_18716,N_18250,N_18221);
and U18717 (N_18717,N_18006,N_18477);
and U18718 (N_18718,N_18116,N_18241);
nor U18719 (N_18719,N_18427,N_18283);
nand U18720 (N_18720,N_18300,N_18176);
and U18721 (N_18721,N_18375,N_18465);
and U18722 (N_18722,N_18112,N_18187);
and U18723 (N_18723,N_18352,N_18014);
nor U18724 (N_18724,N_18060,N_18211);
nand U18725 (N_18725,N_18179,N_18275);
or U18726 (N_18726,N_18470,N_18095);
and U18727 (N_18727,N_18294,N_18220);
nor U18728 (N_18728,N_18466,N_18088);
nor U18729 (N_18729,N_18455,N_18166);
nand U18730 (N_18730,N_18321,N_18099);
nand U18731 (N_18731,N_18165,N_18054);
or U18732 (N_18732,N_18309,N_18120);
nor U18733 (N_18733,N_18405,N_18403);
nand U18734 (N_18734,N_18478,N_18412);
or U18735 (N_18735,N_18344,N_18036);
nand U18736 (N_18736,N_18224,N_18200);
and U18737 (N_18737,N_18257,N_18001);
xnor U18738 (N_18738,N_18402,N_18237);
nand U18739 (N_18739,N_18349,N_18271);
and U18740 (N_18740,N_18424,N_18066);
nor U18741 (N_18741,N_18078,N_18281);
or U18742 (N_18742,N_18388,N_18048);
nor U18743 (N_18743,N_18438,N_18431);
and U18744 (N_18744,N_18129,N_18270);
and U18745 (N_18745,N_18338,N_18256);
nand U18746 (N_18746,N_18199,N_18306);
and U18747 (N_18747,N_18268,N_18032);
nand U18748 (N_18748,N_18009,N_18016);
or U18749 (N_18749,N_18312,N_18064);
and U18750 (N_18750,N_18177,N_18383);
and U18751 (N_18751,N_18382,N_18090);
and U18752 (N_18752,N_18182,N_18156);
or U18753 (N_18753,N_18299,N_18309);
and U18754 (N_18754,N_18207,N_18341);
or U18755 (N_18755,N_18411,N_18232);
and U18756 (N_18756,N_18295,N_18102);
or U18757 (N_18757,N_18302,N_18232);
and U18758 (N_18758,N_18006,N_18408);
xor U18759 (N_18759,N_18019,N_18279);
nand U18760 (N_18760,N_18022,N_18264);
nor U18761 (N_18761,N_18424,N_18146);
and U18762 (N_18762,N_18305,N_18271);
and U18763 (N_18763,N_18064,N_18104);
or U18764 (N_18764,N_18205,N_18437);
nor U18765 (N_18765,N_18262,N_18245);
nor U18766 (N_18766,N_18171,N_18410);
nor U18767 (N_18767,N_18180,N_18143);
nand U18768 (N_18768,N_18427,N_18254);
or U18769 (N_18769,N_18445,N_18040);
and U18770 (N_18770,N_18066,N_18434);
and U18771 (N_18771,N_18121,N_18480);
and U18772 (N_18772,N_18003,N_18464);
nand U18773 (N_18773,N_18004,N_18062);
nand U18774 (N_18774,N_18389,N_18344);
nand U18775 (N_18775,N_18263,N_18386);
nor U18776 (N_18776,N_18107,N_18176);
nand U18777 (N_18777,N_18384,N_18195);
nand U18778 (N_18778,N_18364,N_18152);
nand U18779 (N_18779,N_18380,N_18069);
nand U18780 (N_18780,N_18473,N_18278);
nand U18781 (N_18781,N_18498,N_18252);
nand U18782 (N_18782,N_18472,N_18300);
nor U18783 (N_18783,N_18451,N_18448);
xor U18784 (N_18784,N_18345,N_18249);
nor U18785 (N_18785,N_18387,N_18365);
nor U18786 (N_18786,N_18319,N_18034);
and U18787 (N_18787,N_18329,N_18009);
and U18788 (N_18788,N_18146,N_18112);
nand U18789 (N_18789,N_18243,N_18254);
nand U18790 (N_18790,N_18234,N_18466);
or U18791 (N_18791,N_18457,N_18245);
nand U18792 (N_18792,N_18168,N_18015);
and U18793 (N_18793,N_18052,N_18103);
and U18794 (N_18794,N_18294,N_18051);
or U18795 (N_18795,N_18133,N_18386);
and U18796 (N_18796,N_18281,N_18484);
nand U18797 (N_18797,N_18402,N_18230);
nor U18798 (N_18798,N_18267,N_18475);
nand U18799 (N_18799,N_18337,N_18419);
nor U18800 (N_18800,N_18236,N_18076);
nand U18801 (N_18801,N_18270,N_18132);
or U18802 (N_18802,N_18444,N_18373);
and U18803 (N_18803,N_18087,N_18456);
nor U18804 (N_18804,N_18103,N_18173);
nand U18805 (N_18805,N_18366,N_18009);
or U18806 (N_18806,N_18492,N_18469);
or U18807 (N_18807,N_18340,N_18280);
or U18808 (N_18808,N_18094,N_18078);
and U18809 (N_18809,N_18183,N_18059);
xnor U18810 (N_18810,N_18007,N_18235);
xnor U18811 (N_18811,N_18345,N_18302);
and U18812 (N_18812,N_18193,N_18033);
or U18813 (N_18813,N_18420,N_18063);
nor U18814 (N_18814,N_18261,N_18327);
nor U18815 (N_18815,N_18173,N_18293);
and U18816 (N_18816,N_18105,N_18336);
nand U18817 (N_18817,N_18086,N_18175);
and U18818 (N_18818,N_18187,N_18325);
nor U18819 (N_18819,N_18175,N_18198);
and U18820 (N_18820,N_18313,N_18066);
xor U18821 (N_18821,N_18385,N_18283);
nand U18822 (N_18822,N_18317,N_18081);
or U18823 (N_18823,N_18459,N_18241);
nand U18824 (N_18824,N_18438,N_18063);
xnor U18825 (N_18825,N_18257,N_18207);
and U18826 (N_18826,N_18482,N_18297);
xor U18827 (N_18827,N_18388,N_18098);
and U18828 (N_18828,N_18190,N_18107);
nor U18829 (N_18829,N_18476,N_18182);
nand U18830 (N_18830,N_18141,N_18477);
xor U18831 (N_18831,N_18467,N_18358);
nor U18832 (N_18832,N_18385,N_18473);
or U18833 (N_18833,N_18184,N_18299);
and U18834 (N_18834,N_18497,N_18401);
or U18835 (N_18835,N_18444,N_18395);
nor U18836 (N_18836,N_18232,N_18364);
and U18837 (N_18837,N_18452,N_18027);
nand U18838 (N_18838,N_18109,N_18084);
and U18839 (N_18839,N_18031,N_18479);
and U18840 (N_18840,N_18190,N_18218);
xnor U18841 (N_18841,N_18433,N_18144);
xnor U18842 (N_18842,N_18314,N_18082);
nand U18843 (N_18843,N_18031,N_18218);
nor U18844 (N_18844,N_18402,N_18083);
xor U18845 (N_18845,N_18038,N_18250);
nor U18846 (N_18846,N_18046,N_18069);
or U18847 (N_18847,N_18359,N_18195);
or U18848 (N_18848,N_18024,N_18240);
nor U18849 (N_18849,N_18062,N_18139);
and U18850 (N_18850,N_18352,N_18231);
nor U18851 (N_18851,N_18096,N_18137);
or U18852 (N_18852,N_18277,N_18382);
or U18853 (N_18853,N_18256,N_18483);
and U18854 (N_18854,N_18269,N_18457);
nor U18855 (N_18855,N_18465,N_18334);
nand U18856 (N_18856,N_18424,N_18389);
or U18857 (N_18857,N_18212,N_18428);
nand U18858 (N_18858,N_18438,N_18157);
and U18859 (N_18859,N_18131,N_18155);
xor U18860 (N_18860,N_18029,N_18420);
nor U18861 (N_18861,N_18474,N_18314);
nor U18862 (N_18862,N_18440,N_18457);
nor U18863 (N_18863,N_18155,N_18051);
nand U18864 (N_18864,N_18073,N_18014);
and U18865 (N_18865,N_18165,N_18107);
nand U18866 (N_18866,N_18153,N_18453);
or U18867 (N_18867,N_18237,N_18378);
and U18868 (N_18868,N_18431,N_18016);
and U18869 (N_18869,N_18108,N_18341);
nand U18870 (N_18870,N_18060,N_18176);
and U18871 (N_18871,N_18062,N_18388);
nor U18872 (N_18872,N_18107,N_18489);
nor U18873 (N_18873,N_18150,N_18497);
nor U18874 (N_18874,N_18490,N_18486);
nor U18875 (N_18875,N_18415,N_18148);
xor U18876 (N_18876,N_18202,N_18104);
nor U18877 (N_18877,N_18354,N_18496);
or U18878 (N_18878,N_18187,N_18470);
or U18879 (N_18879,N_18361,N_18157);
and U18880 (N_18880,N_18076,N_18014);
or U18881 (N_18881,N_18183,N_18260);
and U18882 (N_18882,N_18093,N_18152);
and U18883 (N_18883,N_18023,N_18137);
nor U18884 (N_18884,N_18391,N_18326);
nand U18885 (N_18885,N_18231,N_18370);
and U18886 (N_18886,N_18032,N_18178);
or U18887 (N_18887,N_18280,N_18394);
and U18888 (N_18888,N_18121,N_18420);
or U18889 (N_18889,N_18256,N_18223);
nand U18890 (N_18890,N_18027,N_18240);
or U18891 (N_18891,N_18172,N_18206);
nor U18892 (N_18892,N_18180,N_18053);
xnor U18893 (N_18893,N_18075,N_18343);
nand U18894 (N_18894,N_18168,N_18226);
or U18895 (N_18895,N_18246,N_18374);
nor U18896 (N_18896,N_18317,N_18319);
nand U18897 (N_18897,N_18160,N_18117);
and U18898 (N_18898,N_18357,N_18192);
and U18899 (N_18899,N_18436,N_18164);
or U18900 (N_18900,N_18497,N_18465);
nor U18901 (N_18901,N_18173,N_18247);
or U18902 (N_18902,N_18008,N_18249);
nand U18903 (N_18903,N_18308,N_18115);
xor U18904 (N_18904,N_18338,N_18472);
or U18905 (N_18905,N_18246,N_18125);
nand U18906 (N_18906,N_18001,N_18118);
and U18907 (N_18907,N_18164,N_18360);
nor U18908 (N_18908,N_18153,N_18246);
nor U18909 (N_18909,N_18121,N_18076);
nor U18910 (N_18910,N_18239,N_18183);
xor U18911 (N_18911,N_18398,N_18278);
nand U18912 (N_18912,N_18433,N_18285);
and U18913 (N_18913,N_18363,N_18104);
nand U18914 (N_18914,N_18073,N_18199);
nor U18915 (N_18915,N_18194,N_18459);
or U18916 (N_18916,N_18159,N_18476);
nand U18917 (N_18917,N_18405,N_18330);
and U18918 (N_18918,N_18143,N_18387);
and U18919 (N_18919,N_18168,N_18049);
nand U18920 (N_18920,N_18427,N_18321);
xnor U18921 (N_18921,N_18017,N_18176);
or U18922 (N_18922,N_18368,N_18477);
and U18923 (N_18923,N_18294,N_18483);
nor U18924 (N_18924,N_18326,N_18406);
and U18925 (N_18925,N_18497,N_18210);
nor U18926 (N_18926,N_18209,N_18092);
xnor U18927 (N_18927,N_18030,N_18264);
nor U18928 (N_18928,N_18227,N_18332);
and U18929 (N_18929,N_18429,N_18383);
nor U18930 (N_18930,N_18127,N_18462);
or U18931 (N_18931,N_18071,N_18201);
xnor U18932 (N_18932,N_18074,N_18237);
and U18933 (N_18933,N_18456,N_18342);
and U18934 (N_18934,N_18453,N_18146);
nand U18935 (N_18935,N_18116,N_18415);
xor U18936 (N_18936,N_18042,N_18127);
nor U18937 (N_18937,N_18320,N_18230);
nor U18938 (N_18938,N_18492,N_18459);
and U18939 (N_18939,N_18152,N_18140);
nor U18940 (N_18940,N_18059,N_18155);
nand U18941 (N_18941,N_18056,N_18079);
nor U18942 (N_18942,N_18162,N_18298);
nor U18943 (N_18943,N_18494,N_18149);
nor U18944 (N_18944,N_18345,N_18362);
nand U18945 (N_18945,N_18410,N_18209);
xor U18946 (N_18946,N_18308,N_18284);
and U18947 (N_18947,N_18178,N_18148);
nand U18948 (N_18948,N_18197,N_18281);
nor U18949 (N_18949,N_18162,N_18050);
and U18950 (N_18950,N_18306,N_18496);
nand U18951 (N_18951,N_18293,N_18063);
or U18952 (N_18952,N_18196,N_18288);
nand U18953 (N_18953,N_18144,N_18261);
nand U18954 (N_18954,N_18444,N_18267);
nand U18955 (N_18955,N_18206,N_18404);
and U18956 (N_18956,N_18175,N_18075);
nand U18957 (N_18957,N_18286,N_18003);
nand U18958 (N_18958,N_18426,N_18118);
xnor U18959 (N_18959,N_18215,N_18009);
and U18960 (N_18960,N_18232,N_18138);
or U18961 (N_18961,N_18262,N_18291);
xnor U18962 (N_18962,N_18155,N_18119);
nand U18963 (N_18963,N_18307,N_18283);
or U18964 (N_18964,N_18312,N_18011);
and U18965 (N_18965,N_18064,N_18132);
nor U18966 (N_18966,N_18292,N_18064);
nor U18967 (N_18967,N_18123,N_18117);
or U18968 (N_18968,N_18165,N_18296);
and U18969 (N_18969,N_18421,N_18184);
or U18970 (N_18970,N_18288,N_18303);
and U18971 (N_18971,N_18420,N_18471);
nor U18972 (N_18972,N_18493,N_18474);
nor U18973 (N_18973,N_18440,N_18439);
nand U18974 (N_18974,N_18346,N_18031);
xor U18975 (N_18975,N_18319,N_18386);
and U18976 (N_18976,N_18110,N_18015);
or U18977 (N_18977,N_18281,N_18420);
and U18978 (N_18978,N_18424,N_18095);
nor U18979 (N_18979,N_18397,N_18188);
nand U18980 (N_18980,N_18197,N_18240);
or U18981 (N_18981,N_18004,N_18393);
nor U18982 (N_18982,N_18252,N_18193);
and U18983 (N_18983,N_18098,N_18054);
nand U18984 (N_18984,N_18330,N_18404);
or U18985 (N_18985,N_18195,N_18322);
nand U18986 (N_18986,N_18247,N_18424);
nor U18987 (N_18987,N_18450,N_18129);
nor U18988 (N_18988,N_18112,N_18199);
or U18989 (N_18989,N_18484,N_18494);
and U18990 (N_18990,N_18467,N_18089);
and U18991 (N_18991,N_18433,N_18243);
and U18992 (N_18992,N_18389,N_18388);
and U18993 (N_18993,N_18162,N_18063);
xnor U18994 (N_18994,N_18312,N_18366);
nor U18995 (N_18995,N_18128,N_18368);
nor U18996 (N_18996,N_18004,N_18126);
and U18997 (N_18997,N_18314,N_18308);
or U18998 (N_18998,N_18069,N_18116);
nand U18999 (N_18999,N_18488,N_18026);
xor U19000 (N_19000,N_18708,N_18527);
and U19001 (N_19001,N_18524,N_18604);
xnor U19002 (N_19002,N_18645,N_18628);
and U19003 (N_19003,N_18822,N_18773);
nor U19004 (N_19004,N_18697,N_18817);
xnor U19005 (N_19005,N_18720,N_18737);
nand U19006 (N_19006,N_18622,N_18528);
nor U19007 (N_19007,N_18585,N_18784);
or U19008 (N_19008,N_18755,N_18651);
xor U19009 (N_19009,N_18928,N_18503);
nand U19010 (N_19010,N_18938,N_18787);
nor U19011 (N_19011,N_18756,N_18518);
and U19012 (N_19012,N_18570,N_18501);
nand U19013 (N_19013,N_18574,N_18836);
and U19014 (N_19014,N_18620,N_18843);
nor U19015 (N_19015,N_18985,N_18666);
and U19016 (N_19016,N_18839,N_18540);
nor U19017 (N_19017,N_18979,N_18742);
nor U19018 (N_19018,N_18543,N_18971);
nor U19019 (N_19019,N_18996,N_18754);
and U19020 (N_19020,N_18759,N_18687);
nor U19021 (N_19021,N_18724,N_18627);
and U19022 (N_19022,N_18532,N_18733);
and U19023 (N_19023,N_18740,N_18686);
nor U19024 (N_19024,N_18567,N_18646);
and U19025 (N_19025,N_18590,N_18576);
and U19026 (N_19026,N_18989,N_18901);
nand U19027 (N_19027,N_18725,N_18966);
and U19028 (N_19028,N_18772,N_18712);
nand U19029 (N_19029,N_18780,N_18571);
nand U19030 (N_19030,N_18991,N_18587);
nand U19031 (N_19031,N_18856,N_18658);
or U19032 (N_19032,N_18949,N_18738);
nor U19033 (N_19033,N_18509,N_18656);
nand U19034 (N_19034,N_18771,N_18888);
nand U19035 (N_19035,N_18704,N_18654);
and U19036 (N_19036,N_18522,N_18879);
nor U19037 (N_19037,N_18908,N_18769);
nand U19038 (N_19038,N_18547,N_18726);
and U19039 (N_19039,N_18977,N_18806);
nor U19040 (N_19040,N_18748,N_18601);
and U19041 (N_19041,N_18525,N_18707);
nand U19042 (N_19042,N_18828,N_18691);
and U19043 (N_19043,N_18659,N_18680);
or U19044 (N_19044,N_18618,N_18923);
nand U19045 (N_19045,N_18855,N_18785);
nor U19046 (N_19046,N_18500,N_18728);
nand U19047 (N_19047,N_18573,N_18519);
xnor U19048 (N_19048,N_18706,N_18980);
or U19049 (N_19049,N_18997,N_18983);
nor U19050 (N_19050,N_18745,N_18507);
or U19051 (N_19051,N_18894,N_18741);
or U19052 (N_19052,N_18671,N_18911);
and U19053 (N_19053,N_18982,N_18920);
and U19054 (N_19054,N_18994,N_18715);
and U19055 (N_19055,N_18538,N_18634);
or U19056 (N_19056,N_18936,N_18840);
or U19057 (N_19057,N_18611,N_18529);
nand U19058 (N_19058,N_18873,N_18998);
and U19059 (N_19059,N_18837,N_18557);
xor U19060 (N_19060,N_18695,N_18898);
nor U19061 (N_19061,N_18534,N_18871);
nor U19062 (N_19062,N_18692,N_18758);
nor U19063 (N_19063,N_18626,N_18762);
or U19064 (N_19064,N_18790,N_18963);
or U19065 (N_19065,N_18872,N_18635);
nor U19066 (N_19066,N_18841,N_18596);
and U19067 (N_19067,N_18517,N_18816);
and U19068 (N_19068,N_18743,N_18783);
and U19069 (N_19069,N_18801,N_18670);
nor U19070 (N_19070,N_18575,N_18905);
nand U19071 (N_19071,N_18577,N_18776);
nor U19072 (N_19072,N_18629,N_18513);
and U19073 (N_19073,N_18823,N_18912);
nand U19074 (N_19074,N_18674,N_18763);
nand U19075 (N_19075,N_18932,N_18609);
nor U19076 (N_19076,N_18781,N_18520);
nor U19077 (N_19077,N_18545,N_18885);
or U19078 (N_19078,N_18593,N_18633);
or U19079 (N_19079,N_18810,N_18892);
nand U19080 (N_19080,N_18655,N_18988);
nor U19081 (N_19081,N_18610,N_18744);
and U19082 (N_19082,N_18986,N_18650);
nand U19083 (N_19083,N_18564,N_18705);
nand U19084 (N_19084,N_18833,N_18751);
and U19085 (N_19085,N_18955,N_18887);
nand U19086 (N_19086,N_18603,N_18559);
and U19087 (N_19087,N_18796,N_18569);
or U19088 (N_19088,N_18915,N_18530);
nand U19089 (N_19089,N_18586,N_18962);
or U19090 (N_19090,N_18842,N_18964);
and U19091 (N_19091,N_18583,N_18795);
or U19092 (N_19092,N_18945,N_18684);
and U19093 (N_19093,N_18909,N_18794);
or U19094 (N_19094,N_18824,N_18811);
and U19095 (N_19095,N_18825,N_18652);
and U19096 (N_19096,N_18662,N_18753);
nor U19097 (N_19097,N_18690,N_18860);
xor U19098 (N_19098,N_18940,N_18959);
nor U19099 (N_19099,N_18749,N_18789);
and U19100 (N_19100,N_18821,N_18906);
nand U19101 (N_19101,N_18667,N_18891);
nor U19102 (N_19102,N_18799,N_18858);
nor U19103 (N_19103,N_18639,N_18599);
and U19104 (N_19104,N_18995,N_18578);
and U19105 (N_19105,N_18846,N_18808);
nand U19106 (N_19106,N_18869,N_18967);
and U19107 (N_19107,N_18689,N_18957);
and U19108 (N_19108,N_18850,N_18729);
xnor U19109 (N_19109,N_18791,N_18722);
xor U19110 (N_19110,N_18688,N_18660);
xor U19111 (N_19111,N_18902,N_18939);
nor U19112 (N_19112,N_18861,N_18812);
nor U19113 (N_19113,N_18876,N_18731);
or U19114 (N_19114,N_18975,N_18883);
or U19115 (N_19115,N_18640,N_18653);
and U19116 (N_19116,N_18782,N_18927);
and U19117 (N_19117,N_18913,N_18831);
or U19118 (N_19118,N_18919,N_18696);
nor U19119 (N_19119,N_18973,N_18638);
nand U19120 (N_19120,N_18851,N_18714);
nand U19121 (N_19121,N_18899,N_18732);
nor U19122 (N_19122,N_18661,N_18602);
nand U19123 (N_19123,N_18709,N_18968);
nand U19124 (N_19124,N_18711,N_18924);
or U19125 (N_19125,N_18561,N_18535);
xor U19126 (N_19126,N_18965,N_18550);
nor U19127 (N_19127,N_18765,N_18797);
nand U19128 (N_19128,N_18974,N_18558);
or U19129 (N_19129,N_18526,N_18948);
nand U19130 (N_19130,N_18566,N_18699);
nand U19131 (N_19131,N_18895,N_18641);
xnor U19132 (N_19132,N_18676,N_18533);
nand U19133 (N_19133,N_18778,N_18972);
xor U19134 (N_19134,N_18605,N_18969);
or U19135 (N_19135,N_18718,N_18844);
and U19136 (N_19136,N_18516,N_18907);
nand U19137 (N_19137,N_18890,N_18736);
and U19138 (N_19138,N_18954,N_18865);
or U19139 (N_19139,N_18878,N_18944);
and U19140 (N_19140,N_18556,N_18953);
nor U19141 (N_19141,N_18918,N_18942);
and U19142 (N_19142,N_18544,N_18829);
nand U19143 (N_19143,N_18904,N_18643);
nor U19144 (N_19144,N_18621,N_18681);
or U19145 (N_19145,N_18678,N_18752);
nor U19146 (N_19146,N_18929,N_18826);
and U19147 (N_19147,N_18713,N_18579);
nor U19148 (N_19148,N_18760,N_18882);
or U19149 (N_19149,N_18572,N_18900);
nor U19150 (N_19150,N_18508,N_18698);
nand U19151 (N_19151,N_18677,N_18701);
or U19152 (N_19152,N_18636,N_18672);
and U19153 (N_19153,N_18880,N_18875);
nand U19154 (N_19154,N_18694,N_18716);
nor U19155 (N_19155,N_18897,N_18931);
xnor U19156 (N_19156,N_18595,N_18774);
nor U19157 (N_19157,N_18703,N_18830);
and U19158 (N_19158,N_18584,N_18541);
or U19159 (N_19159,N_18625,N_18838);
or U19160 (N_19160,N_18608,N_18648);
nand U19161 (N_19161,N_18588,N_18960);
and U19162 (N_19162,N_18917,N_18592);
and U19163 (N_19163,N_18961,N_18649);
nand U19164 (N_19164,N_18637,N_18852);
or U19165 (N_19165,N_18798,N_18835);
nand U19166 (N_19166,N_18910,N_18976);
and U19167 (N_19167,N_18952,N_18515);
nand U19168 (N_19168,N_18613,N_18792);
nor U19169 (N_19169,N_18616,N_18673);
nand U19170 (N_19170,N_18683,N_18926);
nor U19171 (N_19171,N_18984,N_18597);
and U19172 (N_19172,N_18531,N_18663);
nand U19173 (N_19173,N_18647,N_18549);
nand U19174 (N_19174,N_18903,N_18624);
nand U19175 (N_19175,N_18548,N_18896);
nor U19176 (N_19176,N_18521,N_18542);
and U19177 (N_19177,N_18685,N_18893);
nand U19178 (N_19178,N_18868,N_18632);
or U19179 (N_19179,N_18614,N_18607);
nor U19180 (N_19180,N_18644,N_18886);
xor U19181 (N_19181,N_18615,N_18669);
or U19182 (N_19182,N_18819,N_18803);
or U19183 (N_19183,N_18807,N_18978);
nand U19184 (N_19184,N_18862,N_18657);
nor U19185 (N_19185,N_18770,N_18710);
nor U19186 (N_19186,N_18746,N_18664);
nor U19187 (N_19187,N_18777,N_18668);
nand U19188 (N_19188,N_18665,N_18933);
nor U19189 (N_19189,N_18606,N_18568);
or U19190 (N_19190,N_18943,N_18854);
nor U19191 (N_19191,N_18845,N_18700);
or U19192 (N_19192,N_18553,N_18630);
or U19193 (N_19193,N_18612,N_18813);
nor U19194 (N_19194,N_18934,N_18820);
nor U19195 (N_19195,N_18552,N_18512);
and U19196 (N_19196,N_18779,N_18867);
nand U19197 (N_19197,N_18832,N_18768);
nand U19198 (N_19198,N_18675,N_18565);
xnor U19199 (N_19199,N_18580,N_18546);
nor U19200 (N_19200,N_18992,N_18857);
nor U19201 (N_19201,N_18958,N_18788);
xnor U19202 (N_19202,N_18947,N_18619);
nand U19203 (N_19203,N_18950,N_18999);
or U19204 (N_19204,N_18551,N_18818);
and U19205 (N_19205,N_18510,N_18849);
nand U19206 (N_19206,N_18921,N_18719);
nand U19207 (N_19207,N_18881,N_18623);
or U19208 (N_19208,N_18735,N_18723);
nand U19209 (N_19209,N_18937,N_18600);
nor U19210 (N_19210,N_18589,N_18504);
or U19211 (N_19211,N_18859,N_18809);
or U19212 (N_19212,N_18591,N_18800);
and U19213 (N_19213,N_18946,N_18581);
nand U19214 (N_19214,N_18848,N_18563);
or U19215 (N_19215,N_18935,N_18537);
nand U19216 (N_19216,N_18562,N_18682);
and U19217 (N_19217,N_18930,N_18877);
nor U19218 (N_19218,N_18721,N_18702);
nor U19219 (N_19219,N_18536,N_18814);
and U19220 (N_19220,N_18827,N_18922);
or U19221 (N_19221,N_18617,N_18631);
nand U19222 (N_19222,N_18775,N_18505);
or U19223 (N_19223,N_18863,N_18853);
nor U19224 (N_19224,N_18511,N_18916);
and U19225 (N_19225,N_18764,N_18679);
xor U19226 (N_19226,N_18730,N_18956);
and U19227 (N_19227,N_18805,N_18747);
xnor U19228 (N_19228,N_18802,N_18642);
nor U19229 (N_19229,N_18925,N_18598);
and U19230 (N_19230,N_18757,N_18523);
nand U19231 (N_19231,N_18884,N_18874);
xnor U19232 (N_19232,N_18734,N_18951);
nor U19233 (N_19233,N_18717,N_18970);
nand U19234 (N_19234,N_18594,N_18914);
nor U19235 (N_19235,N_18864,N_18889);
nor U19236 (N_19236,N_18981,N_18761);
or U19237 (N_19237,N_18793,N_18554);
and U19238 (N_19238,N_18766,N_18560);
xnor U19239 (N_19239,N_18506,N_18582);
xnor U19240 (N_19240,N_18786,N_18750);
or U19241 (N_19241,N_18990,N_18987);
or U19242 (N_19242,N_18815,N_18804);
nor U19243 (N_19243,N_18555,N_18870);
nor U19244 (N_19244,N_18847,N_18739);
and U19245 (N_19245,N_18941,N_18866);
nand U19246 (N_19246,N_18693,N_18993);
nand U19247 (N_19247,N_18539,N_18727);
nor U19248 (N_19248,N_18834,N_18502);
nor U19249 (N_19249,N_18767,N_18514);
and U19250 (N_19250,N_18505,N_18583);
and U19251 (N_19251,N_18540,N_18929);
nor U19252 (N_19252,N_18968,N_18519);
or U19253 (N_19253,N_18977,N_18667);
nand U19254 (N_19254,N_18764,N_18676);
nor U19255 (N_19255,N_18934,N_18844);
nand U19256 (N_19256,N_18853,N_18822);
nand U19257 (N_19257,N_18568,N_18981);
nand U19258 (N_19258,N_18948,N_18694);
nor U19259 (N_19259,N_18537,N_18863);
or U19260 (N_19260,N_18914,N_18851);
or U19261 (N_19261,N_18542,N_18943);
nor U19262 (N_19262,N_18558,N_18881);
or U19263 (N_19263,N_18715,N_18576);
xor U19264 (N_19264,N_18854,N_18547);
nor U19265 (N_19265,N_18982,N_18804);
nor U19266 (N_19266,N_18826,N_18940);
xnor U19267 (N_19267,N_18686,N_18906);
nor U19268 (N_19268,N_18898,N_18702);
xor U19269 (N_19269,N_18657,N_18777);
nor U19270 (N_19270,N_18829,N_18672);
xor U19271 (N_19271,N_18854,N_18996);
nand U19272 (N_19272,N_18771,N_18640);
or U19273 (N_19273,N_18593,N_18557);
nor U19274 (N_19274,N_18942,N_18848);
nor U19275 (N_19275,N_18865,N_18794);
or U19276 (N_19276,N_18682,N_18553);
nor U19277 (N_19277,N_18664,N_18661);
nand U19278 (N_19278,N_18596,N_18849);
and U19279 (N_19279,N_18685,N_18819);
nand U19280 (N_19280,N_18935,N_18983);
and U19281 (N_19281,N_18835,N_18873);
nor U19282 (N_19282,N_18602,N_18738);
nor U19283 (N_19283,N_18874,N_18742);
nor U19284 (N_19284,N_18847,N_18914);
or U19285 (N_19285,N_18829,N_18557);
and U19286 (N_19286,N_18905,N_18984);
or U19287 (N_19287,N_18971,N_18825);
nand U19288 (N_19288,N_18996,N_18617);
xnor U19289 (N_19289,N_18819,N_18818);
xnor U19290 (N_19290,N_18616,N_18832);
nand U19291 (N_19291,N_18873,N_18858);
nor U19292 (N_19292,N_18617,N_18833);
nand U19293 (N_19293,N_18776,N_18921);
and U19294 (N_19294,N_18514,N_18853);
or U19295 (N_19295,N_18738,N_18762);
nand U19296 (N_19296,N_18721,N_18894);
nor U19297 (N_19297,N_18693,N_18535);
nand U19298 (N_19298,N_18586,N_18977);
and U19299 (N_19299,N_18739,N_18779);
nor U19300 (N_19300,N_18788,N_18873);
nor U19301 (N_19301,N_18743,N_18643);
xor U19302 (N_19302,N_18666,N_18850);
nand U19303 (N_19303,N_18543,N_18682);
or U19304 (N_19304,N_18866,N_18863);
or U19305 (N_19305,N_18894,N_18989);
xor U19306 (N_19306,N_18849,N_18559);
and U19307 (N_19307,N_18732,N_18866);
nor U19308 (N_19308,N_18800,N_18745);
or U19309 (N_19309,N_18605,N_18640);
nand U19310 (N_19310,N_18624,N_18834);
and U19311 (N_19311,N_18912,N_18788);
and U19312 (N_19312,N_18989,N_18671);
nand U19313 (N_19313,N_18838,N_18878);
nand U19314 (N_19314,N_18841,N_18695);
nand U19315 (N_19315,N_18800,N_18548);
xor U19316 (N_19316,N_18867,N_18852);
and U19317 (N_19317,N_18825,N_18626);
xor U19318 (N_19318,N_18568,N_18746);
nand U19319 (N_19319,N_18893,N_18817);
nor U19320 (N_19320,N_18567,N_18976);
or U19321 (N_19321,N_18584,N_18909);
nor U19322 (N_19322,N_18674,N_18660);
nand U19323 (N_19323,N_18564,N_18990);
nand U19324 (N_19324,N_18652,N_18600);
or U19325 (N_19325,N_18706,N_18690);
and U19326 (N_19326,N_18661,N_18828);
xnor U19327 (N_19327,N_18589,N_18540);
nor U19328 (N_19328,N_18883,N_18891);
nand U19329 (N_19329,N_18964,N_18638);
or U19330 (N_19330,N_18868,N_18837);
or U19331 (N_19331,N_18531,N_18790);
or U19332 (N_19332,N_18879,N_18560);
nor U19333 (N_19333,N_18735,N_18640);
or U19334 (N_19334,N_18918,N_18737);
nand U19335 (N_19335,N_18575,N_18845);
or U19336 (N_19336,N_18915,N_18726);
and U19337 (N_19337,N_18696,N_18619);
or U19338 (N_19338,N_18539,N_18782);
xnor U19339 (N_19339,N_18587,N_18589);
nand U19340 (N_19340,N_18771,N_18870);
and U19341 (N_19341,N_18876,N_18867);
nand U19342 (N_19342,N_18761,N_18667);
and U19343 (N_19343,N_18713,N_18883);
nand U19344 (N_19344,N_18614,N_18653);
xnor U19345 (N_19345,N_18674,N_18932);
or U19346 (N_19346,N_18926,N_18507);
xor U19347 (N_19347,N_18711,N_18892);
nand U19348 (N_19348,N_18719,N_18803);
or U19349 (N_19349,N_18654,N_18671);
or U19350 (N_19350,N_18679,N_18735);
xor U19351 (N_19351,N_18539,N_18627);
nor U19352 (N_19352,N_18695,N_18861);
or U19353 (N_19353,N_18708,N_18625);
nand U19354 (N_19354,N_18991,N_18958);
nor U19355 (N_19355,N_18898,N_18843);
or U19356 (N_19356,N_18641,N_18591);
and U19357 (N_19357,N_18656,N_18930);
xor U19358 (N_19358,N_18966,N_18866);
nand U19359 (N_19359,N_18829,N_18664);
or U19360 (N_19360,N_18703,N_18743);
and U19361 (N_19361,N_18855,N_18764);
and U19362 (N_19362,N_18593,N_18988);
nand U19363 (N_19363,N_18677,N_18621);
nand U19364 (N_19364,N_18914,N_18576);
and U19365 (N_19365,N_18995,N_18526);
nand U19366 (N_19366,N_18803,N_18746);
nand U19367 (N_19367,N_18764,N_18744);
and U19368 (N_19368,N_18512,N_18995);
nor U19369 (N_19369,N_18763,N_18908);
or U19370 (N_19370,N_18853,N_18760);
xnor U19371 (N_19371,N_18822,N_18607);
nand U19372 (N_19372,N_18560,N_18942);
or U19373 (N_19373,N_18729,N_18676);
nand U19374 (N_19374,N_18841,N_18977);
and U19375 (N_19375,N_18781,N_18658);
and U19376 (N_19376,N_18954,N_18631);
nor U19377 (N_19377,N_18939,N_18894);
nand U19378 (N_19378,N_18896,N_18891);
nand U19379 (N_19379,N_18872,N_18608);
nor U19380 (N_19380,N_18604,N_18624);
and U19381 (N_19381,N_18953,N_18601);
nor U19382 (N_19382,N_18801,N_18837);
xor U19383 (N_19383,N_18788,N_18906);
xnor U19384 (N_19384,N_18993,N_18777);
nand U19385 (N_19385,N_18792,N_18887);
or U19386 (N_19386,N_18799,N_18638);
nor U19387 (N_19387,N_18721,N_18963);
and U19388 (N_19388,N_18666,N_18786);
nand U19389 (N_19389,N_18874,N_18996);
nor U19390 (N_19390,N_18781,N_18659);
and U19391 (N_19391,N_18724,N_18516);
and U19392 (N_19392,N_18954,N_18712);
xnor U19393 (N_19393,N_18805,N_18929);
xor U19394 (N_19394,N_18984,N_18627);
and U19395 (N_19395,N_18901,N_18786);
nor U19396 (N_19396,N_18737,N_18744);
nand U19397 (N_19397,N_18897,N_18534);
and U19398 (N_19398,N_18951,N_18957);
or U19399 (N_19399,N_18757,N_18617);
nor U19400 (N_19400,N_18848,N_18906);
or U19401 (N_19401,N_18632,N_18729);
xor U19402 (N_19402,N_18833,N_18664);
nand U19403 (N_19403,N_18538,N_18792);
and U19404 (N_19404,N_18808,N_18653);
or U19405 (N_19405,N_18950,N_18881);
and U19406 (N_19406,N_18749,N_18819);
and U19407 (N_19407,N_18711,N_18867);
and U19408 (N_19408,N_18737,N_18919);
or U19409 (N_19409,N_18723,N_18917);
xor U19410 (N_19410,N_18945,N_18702);
xnor U19411 (N_19411,N_18988,N_18916);
nand U19412 (N_19412,N_18695,N_18596);
nand U19413 (N_19413,N_18600,N_18895);
or U19414 (N_19414,N_18556,N_18957);
and U19415 (N_19415,N_18579,N_18658);
nor U19416 (N_19416,N_18764,N_18746);
or U19417 (N_19417,N_18559,N_18785);
nor U19418 (N_19418,N_18526,N_18808);
nand U19419 (N_19419,N_18684,N_18542);
nand U19420 (N_19420,N_18793,N_18982);
nand U19421 (N_19421,N_18707,N_18703);
and U19422 (N_19422,N_18784,N_18552);
or U19423 (N_19423,N_18851,N_18999);
and U19424 (N_19424,N_18795,N_18931);
nand U19425 (N_19425,N_18712,N_18515);
or U19426 (N_19426,N_18525,N_18688);
and U19427 (N_19427,N_18846,N_18507);
or U19428 (N_19428,N_18572,N_18873);
nor U19429 (N_19429,N_18512,N_18786);
nor U19430 (N_19430,N_18867,N_18736);
and U19431 (N_19431,N_18943,N_18820);
and U19432 (N_19432,N_18736,N_18810);
nand U19433 (N_19433,N_18821,N_18546);
nor U19434 (N_19434,N_18999,N_18776);
or U19435 (N_19435,N_18914,N_18706);
and U19436 (N_19436,N_18940,N_18715);
nor U19437 (N_19437,N_18853,N_18983);
or U19438 (N_19438,N_18839,N_18862);
nor U19439 (N_19439,N_18930,N_18505);
nand U19440 (N_19440,N_18766,N_18787);
and U19441 (N_19441,N_18756,N_18535);
and U19442 (N_19442,N_18890,N_18771);
xnor U19443 (N_19443,N_18639,N_18969);
and U19444 (N_19444,N_18696,N_18537);
and U19445 (N_19445,N_18693,N_18911);
or U19446 (N_19446,N_18975,N_18971);
or U19447 (N_19447,N_18960,N_18833);
or U19448 (N_19448,N_18946,N_18639);
and U19449 (N_19449,N_18888,N_18729);
and U19450 (N_19450,N_18944,N_18643);
nor U19451 (N_19451,N_18915,N_18854);
and U19452 (N_19452,N_18808,N_18972);
and U19453 (N_19453,N_18946,N_18806);
and U19454 (N_19454,N_18935,N_18703);
nor U19455 (N_19455,N_18720,N_18898);
and U19456 (N_19456,N_18757,N_18662);
and U19457 (N_19457,N_18980,N_18553);
or U19458 (N_19458,N_18716,N_18511);
and U19459 (N_19459,N_18524,N_18561);
and U19460 (N_19460,N_18760,N_18732);
xor U19461 (N_19461,N_18601,N_18730);
or U19462 (N_19462,N_18858,N_18717);
nand U19463 (N_19463,N_18748,N_18538);
nor U19464 (N_19464,N_18802,N_18818);
nand U19465 (N_19465,N_18887,N_18505);
xnor U19466 (N_19466,N_18688,N_18627);
nand U19467 (N_19467,N_18688,N_18658);
nand U19468 (N_19468,N_18614,N_18726);
and U19469 (N_19469,N_18578,N_18799);
nor U19470 (N_19470,N_18702,N_18845);
nand U19471 (N_19471,N_18793,N_18622);
and U19472 (N_19472,N_18940,N_18614);
xor U19473 (N_19473,N_18710,N_18651);
and U19474 (N_19474,N_18562,N_18611);
xnor U19475 (N_19475,N_18712,N_18697);
xor U19476 (N_19476,N_18833,N_18514);
and U19477 (N_19477,N_18791,N_18530);
and U19478 (N_19478,N_18611,N_18538);
and U19479 (N_19479,N_18724,N_18788);
nand U19480 (N_19480,N_18597,N_18930);
nor U19481 (N_19481,N_18580,N_18764);
nor U19482 (N_19482,N_18658,N_18715);
nor U19483 (N_19483,N_18879,N_18741);
or U19484 (N_19484,N_18719,N_18951);
nand U19485 (N_19485,N_18671,N_18854);
nor U19486 (N_19486,N_18826,N_18994);
nor U19487 (N_19487,N_18761,N_18726);
and U19488 (N_19488,N_18506,N_18992);
or U19489 (N_19489,N_18761,N_18822);
or U19490 (N_19490,N_18735,N_18925);
nor U19491 (N_19491,N_18781,N_18822);
and U19492 (N_19492,N_18960,N_18618);
nand U19493 (N_19493,N_18680,N_18976);
xnor U19494 (N_19494,N_18816,N_18871);
and U19495 (N_19495,N_18993,N_18944);
nor U19496 (N_19496,N_18741,N_18580);
nand U19497 (N_19497,N_18843,N_18817);
or U19498 (N_19498,N_18999,N_18623);
or U19499 (N_19499,N_18849,N_18584);
nand U19500 (N_19500,N_19029,N_19084);
or U19501 (N_19501,N_19129,N_19406);
nor U19502 (N_19502,N_19237,N_19093);
nand U19503 (N_19503,N_19281,N_19303);
nor U19504 (N_19504,N_19257,N_19349);
nor U19505 (N_19505,N_19171,N_19321);
nor U19506 (N_19506,N_19099,N_19138);
and U19507 (N_19507,N_19497,N_19298);
xor U19508 (N_19508,N_19162,N_19293);
and U19509 (N_19509,N_19430,N_19197);
nor U19510 (N_19510,N_19477,N_19010);
nand U19511 (N_19511,N_19011,N_19377);
nand U19512 (N_19512,N_19492,N_19233);
or U19513 (N_19513,N_19285,N_19161);
and U19514 (N_19514,N_19498,N_19345);
or U19515 (N_19515,N_19135,N_19168);
nand U19516 (N_19516,N_19164,N_19317);
or U19517 (N_19517,N_19155,N_19122);
nand U19518 (N_19518,N_19152,N_19295);
or U19519 (N_19519,N_19254,N_19177);
xor U19520 (N_19520,N_19417,N_19100);
and U19521 (N_19521,N_19215,N_19310);
nor U19522 (N_19522,N_19314,N_19401);
and U19523 (N_19523,N_19399,N_19361);
and U19524 (N_19524,N_19114,N_19206);
nand U19525 (N_19525,N_19353,N_19278);
nor U19526 (N_19526,N_19242,N_19104);
nor U19527 (N_19527,N_19185,N_19072);
and U19528 (N_19528,N_19279,N_19284);
and U19529 (N_19529,N_19096,N_19064);
and U19530 (N_19530,N_19415,N_19355);
nor U19531 (N_19531,N_19336,N_19101);
xnor U19532 (N_19532,N_19250,N_19329);
and U19533 (N_19533,N_19360,N_19455);
xor U19534 (N_19534,N_19165,N_19069);
nor U19535 (N_19535,N_19202,N_19465);
or U19536 (N_19536,N_19179,N_19013);
nand U19537 (N_19537,N_19283,N_19265);
nand U19538 (N_19538,N_19367,N_19423);
nor U19539 (N_19539,N_19484,N_19103);
or U19540 (N_19540,N_19024,N_19395);
and U19541 (N_19541,N_19089,N_19343);
nand U19542 (N_19542,N_19494,N_19456);
xor U19543 (N_19543,N_19378,N_19228);
and U19544 (N_19544,N_19150,N_19174);
or U19545 (N_19545,N_19083,N_19366);
nor U19546 (N_19546,N_19264,N_19074);
nor U19547 (N_19547,N_19469,N_19490);
nand U19548 (N_19548,N_19212,N_19340);
and U19549 (N_19549,N_19200,N_19478);
or U19550 (N_19550,N_19239,N_19312);
nor U19551 (N_19551,N_19282,N_19144);
and U19552 (N_19552,N_19025,N_19141);
or U19553 (N_19553,N_19163,N_19274);
or U19554 (N_19554,N_19092,N_19365);
and U19555 (N_19555,N_19289,N_19180);
and U19556 (N_19556,N_19404,N_19139);
nor U19557 (N_19557,N_19449,N_19326);
and U19558 (N_19558,N_19117,N_19263);
or U19559 (N_19559,N_19389,N_19189);
nand U19560 (N_19560,N_19426,N_19061);
and U19561 (N_19561,N_19333,N_19454);
nor U19562 (N_19562,N_19322,N_19040);
nand U19563 (N_19563,N_19243,N_19451);
and U19564 (N_19564,N_19043,N_19082);
nand U19565 (N_19565,N_19255,N_19062);
and U19566 (N_19566,N_19119,N_19390);
and U19567 (N_19567,N_19223,N_19393);
and U19568 (N_19568,N_19194,N_19488);
nor U19569 (N_19569,N_19148,N_19300);
nor U19570 (N_19570,N_19009,N_19370);
nand U19571 (N_19571,N_19166,N_19066);
and U19572 (N_19572,N_19409,N_19432);
and U19573 (N_19573,N_19338,N_19457);
nand U19574 (N_19574,N_19435,N_19302);
nand U19575 (N_19575,N_19070,N_19363);
or U19576 (N_19576,N_19173,N_19036);
and U19577 (N_19577,N_19067,N_19416);
and U19578 (N_19578,N_19113,N_19203);
nand U19579 (N_19579,N_19238,N_19486);
xor U19580 (N_19580,N_19065,N_19109);
nor U19581 (N_19581,N_19499,N_19324);
and U19582 (N_19582,N_19211,N_19019);
nand U19583 (N_19583,N_19448,N_19294);
or U19584 (N_19584,N_19226,N_19419);
and U19585 (N_19585,N_19030,N_19334);
and U19586 (N_19586,N_19470,N_19346);
or U19587 (N_19587,N_19364,N_19268);
nor U19588 (N_19588,N_19485,N_19459);
nor U19589 (N_19589,N_19311,N_19436);
or U19590 (N_19590,N_19248,N_19088);
nor U19591 (N_19591,N_19269,N_19258);
nor U19592 (N_19592,N_19327,N_19115);
and U19593 (N_19593,N_19033,N_19041);
and U19594 (N_19594,N_19319,N_19146);
or U19595 (N_19595,N_19288,N_19397);
nor U19596 (N_19596,N_19190,N_19315);
nor U19597 (N_19597,N_19308,N_19304);
nand U19598 (N_19598,N_19352,N_19178);
nand U19599 (N_19599,N_19266,N_19480);
and U19600 (N_19600,N_19199,N_19079);
or U19601 (N_19601,N_19095,N_19388);
xor U19602 (N_19602,N_19332,N_19188);
or U19603 (N_19603,N_19493,N_19328);
and U19604 (N_19604,N_19128,N_19054);
nor U19605 (N_19605,N_19482,N_19374);
nor U19606 (N_19606,N_19342,N_19112);
and U19607 (N_19607,N_19496,N_19217);
nand U19608 (N_19608,N_19231,N_19331);
nand U19609 (N_19609,N_19198,N_19261);
and U19610 (N_19610,N_19309,N_19461);
or U19611 (N_19611,N_19458,N_19381);
or U19612 (N_19612,N_19136,N_19297);
or U19613 (N_19613,N_19132,N_19464);
nor U19614 (N_19614,N_19241,N_19276);
nor U19615 (N_19615,N_19330,N_19037);
or U19616 (N_19616,N_19042,N_19046);
nand U19617 (N_19617,N_19437,N_19421);
nand U19618 (N_19618,N_19251,N_19186);
and U19619 (N_19619,N_19442,N_19473);
nand U19620 (N_19620,N_19182,N_19240);
or U19621 (N_19621,N_19209,N_19472);
xor U19622 (N_19622,N_19181,N_19118);
and U19623 (N_19623,N_19051,N_19175);
nand U19624 (N_19624,N_19440,N_19005);
and U19625 (N_19625,N_19476,N_19354);
nor U19626 (N_19626,N_19433,N_19286);
nor U19627 (N_19627,N_19149,N_19154);
nor U19628 (N_19628,N_19375,N_19387);
xor U19629 (N_19629,N_19380,N_19467);
nand U19630 (N_19630,N_19259,N_19439);
nor U19631 (N_19631,N_19411,N_19272);
or U19632 (N_19632,N_19376,N_19438);
or U19633 (N_19633,N_19253,N_19147);
nand U19634 (N_19634,N_19450,N_19057);
nand U19635 (N_19635,N_19235,N_19016);
xnor U19636 (N_19636,N_19050,N_19191);
and U19637 (N_19637,N_19245,N_19134);
or U19638 (N_19638,N_19167,N_19140);
xor U19639 (N_19639,N_19244,N_19444);
nor U19640 (N_19640,N_19468,N_19462);
nand U19641 (N_19641,N_19106,N_19222);
and U19642 (N_19642,N_19172,N_19280);
nor U19643 (N_19643,N_19445,N_19313);
xor U19644 (N_19644,N_19169,N_19006);
xnor U19645 (N_19645,N_19252,N_19425);
nand U19646 (N_19646,N_19022,N_19205);
or U19647 (N_19647,N_19108,N_19145);
xor U19648 (N_19648,N_19369,N_19218);
and U19649 (N_19649,N_19463,N_19151);
or U19650 (N_19650,N_19133,N_19143);
xnor U19651 (N_19651,N_19098,N_19120);
or U19652 (N_19652,N_19073,N_19059);
and U19653 (N_19653,N_19058,N_19021);
or U19654 (N_19654,N_19213,N_19008);
and U19655 (N_19655,N_19225,N_19012);
nand U19656 (N_19656,N_19187,N_19420);
or U19657 (N_19657,N_19398,N_19039);
and U19658 (N_19658,N_19396,N_19474);
nand U19659 (N_19659,N_19017,N_19410);
xnor U19660 (N_19660,N_19344,N_19032);
xor U19661 (N_19661,N_19479,N_19111);
and U19662 (N_19662,N_19339,N_19236);
and U19663 (N_19663,N_19385,N_19495);
and U19664 (N_19664,N_19153,N_19158);
nor U19665 (N_19665,N_19193,N_19232);
and U19666 (N_19666,N_19210,N_19075);
nor U19667 (N_19667,N_19038,N_19481);
nor U19668 (N_19668,N_19031,N_19383);
nand U19669 (N_19669,N_19382,N_19219);
or U19670 (N_19670,N_19086,N_19077);
and U19671 (N_19671,N_19256,N_19045);
nor U19672 (N_19672,N_19359,N_19156);
and U19673 (N_19673,N_19224,N_19160);
or U19674 (N_19674,N_19471,N_19071);
xnor U19675 (N_19675,N_19137,N_19299);
nand U19676 (N_19676,N_19076,N_19348);
or U19677 (N_19677,N_19301,N_19052);
and U19678 (N_19678,N_19267,N_19405);
nor U19679 (N_19679,N_19443,N_19384);
nor U19680 (N_19680,N_19123,N_19105);
and U19681 (N_19681,N_19414,N_19216);
nor U19682 (N_19682,N_19028,N_19001);
xor U19683 (N_19683,N_19453,N_19371);
and U19684 (N_19684,N_19446,N_19452);
nand U19685 (N_19685,N_19434,N_19080);
nand U19686 (N_19686,N_19227,N_19356);
or U19687 (N_19687,N_19307,N_19026);
nor U19688 (N_19688,N_19287,N_19027);
and U19689 (N_19689,N_19131,N_19142);
nand U19690 (N_19690,N_19402,N_19192);
nand U19691 (N_19691,N_19130,N_19373);
and U19692 (N_19692,N_19273,N_19427);
and U19693 (N_19693,N_19403,N_19091);
nor U19694 (N_19694,N_19004,N_19418);
or U19695 (N_19695,N_19291,N_19170);
or U19696 (N_19696,N_19491,N_19277);
nor U19697 (N_19697,N_19475,N_19422);
nor U19698 (N_19698,N_19368,N_19483);
nand U19699 (N_19699,N_19335,N_19362);
xor U19700 (N_19700,N_19127,N_19220);
nor U19701 (N_19701,N_19275,N_19090);
and U19702 (N_19702,N_19081,N_19379);
or U19703 (N_19703,N_19372,N_19044);
nand U19704 (N_19704,N_19262,N_19053);
xor U19705 (N_19705,N_19247,N_19094);
xor U19706 (N_19706,N_19229,N_19157);
nor U19707 (N_19707,N_19015,N_19102);
xnor U19708 (N_19708,N_19358,N_19018);
or U19709 (N_19709,N_19020,N_19121);
xor U19710 (N_19710,N_19208,N_19408);
or U19711 (N_19711,N_19023,N_19320);
or U19712 (N_19712,N_19047,N_19110);
or U19713 (N_19713,N_19201,N_19176);
and U19714 (N_19714,N_19407,N_19400);
nor U19715 (N_19715,N_19068,N_19316);
nand U19716 (N_19716,N_19124,N_19195);
or U19717 (N_19717,N_19391,N_19296);
nand U19718 (N_19718,N_19428,N_19014);
and U19719 (N_19719,N_19429,N_19003);
nand U19720 (N_19720,N_19063,N_19196);
or U19721 (N_19721,N_19204,N_19035);
or U19722 (N_19722,N_19078,N_19126);
nor U19723 (N_19723,N_19323,N_19350);
nor U19724 (N_19724,N_19234,N_19392);
nand U19725 (N_19725,N_19159,N_19249);
nor U19726 (N_19726,N_19318,N_19447);
and U19727 (N_19727,N_19489,N_19048);
nand U19728 (N_19728,N_19056,N_19441);
and U19729 (N_19729,N_19325,N_19230);
nand U19730 (N_19730,N_19221,N_19183);
nor U19731 (N_19731,N_19413,N_19424);
and U19732 (N_19732,N_19116,N_19460);
nor U19733 (N_19733,N_19125,N_19431);
nor U19734 (N_19734,N_19246,N_19007);
nor U19735 (N_19735,N_19386,N_19184);
and U19736 (N_19736,N_19214,N_19055);
or U19737 (N_19737,N_19357,N_19049);
nor U19738 (N_19738,N_19270,N_19085);
xor U19739 (N_19739,N_19260,N_19060);
nand U19740 (N_19740,N_19347,N_19107);
nor U19741 (N_19741,N_19271,N_19207);
and U19742 (N_19742,N_19002,N_19034);
nand U19743 (N_19743,N_19290,N_19394);
xnor U19744 (N_19744,N_19466,N_19341);
nor U19745 (N_19745,N_19487,N_19351);
and U19746 (N_19746,N_19412,N_19292);
or U19747 (N_19747,N_19305,N_19000);
or U19748 (N_19748,N_19306,N_19337);
nor U19749 (N_19749,N_19087,N_19097);
nand U19750 (N_19750,N_19470,N_19069);
nor U19751 (N_19751,N_19280,N_19311);
or U19752 (N_19752,N_19101,N_19416);
or U19753 (N_19753,N_19154,N_19000);
nand U19754 (N_19754,N_19424,N_19446);
and U19755 (N_19755,N_19290,N_19191);
nor U19756 (N_19756,N_19149,N_19441);
nor U19757 (N_19757,N_19369,N_19098);
and U19758 (N_19758,N_19266,N_19441);
or U19759 (N_19759,N_19107,N_19187);
nor U19760 (N_19760,N_19360,N_19168);
nand U19761 (N_19761,N_19187,N_19437);
and U19762 (N_19762,N_19240,N_19474);
nand U19763 (N_19763,N_19011,N_19200);
nand U19764 (N_19764,N_19025,N_19084);
nor U19765 (N_19765,N_19311,N_19110);
and U19766 (N_19766,N_19050,N_19315);
nor U19767 (N_19767,N_19364,N_19335);
or U19768 (N_19768,N_19177,N_19247);
nor U19769 (N_19769,N_19209,N_19068);
nand U19770 (N_19770,N_19435,N_19083);
nand U19771 (N_19771,N_19388,N_19149);
xor U19772 (N_19772,N_19167,N_19194);
or U19773 (N_19773,N_19027,N_19315);
and U19774 (N_19774,N_19286,N_19135);
nor U19775 (N_19775,N_19242,N_19226);
or U19776 (N_19776,N_19178,N_19080);
and U19777 (N_19777,N_19491,N_19274);
nand U19778 (N_19778,N_19175,N_19449);
nor U19779 (N_19779,N_19033,N_19426);
and U19780 (N_19780,N_19472,N_19292);
and U19781 (N_19781,N_19456,N_19336);
nand U19782 (N_19782,N_19226,N_19195);
xnor U19783 (N_19783,N_19296,N_19174);
or U19784 (N_19784,N_19179,N_19163);
or U19785 (N_19785,N_19174,N_19204);
and U19786 (N_19786,N_19374,N_19026);
or U19787 (N_19787,N_19109,N_19441);
nand U19788 (N_19788,N_19489,N_19202);
or U19789 (N_19789,N_19172,N_19333);
xor U19790 (N_19790,N_19429,N_19382);
nand U19791 (N_19791,N_19493,N_19409);
or U19792 (N_19792,N_19115,N_19252);
and U19793 (N_19793,N_19316,N_19080);
and U19794 (N_19794,N_19280,N_19045);
nand U19795 (N_19795,N_19398,N_19109);
or U19796 (N_19796,N_19237,N_19080);
or U19797 (N_19797,N_19303,N_19123);
nor U19798 (N_19798,N_19077,N_19338);
and U19799 (N_19799,N_19355,N_19183);
xnor U19800 (N_19800,N_19385,N_19098);
nor U19801 (N_19801,N_19111,N_19143);
nor U19802 (N_19802,N_19342,N_19048);
or U19803 (N_19803,N_19003,N_19498);
nor U19804 (N_19804,N_19092,N_19103);
nor U19805 (N_19805,N_19377,N_19053);
nor U19806 (N_19806,N_19332,N_19148);
or U19807 (N_19807,N_19255,N_19317);
and U19808 (N_19808,N_19105,N_19323);
nand U19809 (N_19809,N_19419,N_19426);
nand U19810 (N_19810,N_19169,N_19257);
or U19811 (N_19811,N_19182,N_19183);
and U19812 (N_19812,N_19309,N_19304);
nor U19813 (N_19813,N_19460,N_19050);
or U19814 (N_19814,N_19362,N_19075);
nand U19815 (N_19815,N_19032,N_19274);
nand U19816 (N_19816,N_19212,N_19314);
xnor U19817 (N_19817,N_19158,N_19213);
nand U19818 (N_19818,N_19132,N_19382);
nor U19819 (N_19819,N_19434,N_19237);
nand U19820 (N_19820,N_19140,N_19353);
or U19821 (N_19821,N_19004,N_19220);
nand U19822 (N_19822,N_19305,N_19257);
nor U19823 (N_19823,N_19468,N_19047);
nor U19824 (N_19824,N_19123,N_19032);
or U19825 (N_19825,N_19326,N_19481);
nor U19826 (N_19826,N_19153,N_19187);
nor U19827 (N_19827,N_19199,N_19051);
nor U19828 (N_19828,N_19340,N_19497);
nand U19829 (N_19829,N_19126,N_19093);
or U19830 (N_19830,N_19376,N_19433);
and U19831 (N_19831,N_19292,N_19331);
or U19832 (N_19832,N_19278,N_19422);
nor U19833 (N_19833,N_19482,N_19227);
nand U19834 (N_19834,N_19326,N_19405);
or U19835 (N_19835,N_19225,N_19253);
xor U19836 (N_19836,N_19058,N_19254);
nor U19837 (N_19837,N_19126,N_19242);
and U19838 (N_19838,N_19102,N_19157);
nand U19839 (N_19839,N_19049,N_19466);
and U19840 (N_19840,N_19320,N_19378);
nand U19841 (N_19841,N_19474,N_19397);
nand U19842 (N_19842,N_19266,N_19135);
and U19843 (N_19843,N_19130,N_19279);
nor U19844 (N_19844,N_19467,N_19000);
or U19845 (N_19845,N_19235,N_19490);
nand U19846 (N_19846,N_19482,N_19213);
nor U19847 (N_19847,N_19197,N_19160);
nor U19848 (N_19848,N_19410,N_19060);
and U19849 (N_19849,N_19307,N_19037);
and U19850 (N_19850,N_19018,N_19441);
nor U19851 (N_19851,N_19481,N_19402);
nand U19852 (N_19852,N_19418,N_19151);
and U19853 (N_19853,N_19312,N_19184);
nor U19854 (N_19854,N_19265,N_19429);
nor U19855 (N_19855,N_19368,N_19025);
and U19856 (N_19856,N_19444,N_19247);
nor U19857 (N_19857,N_19456,N_19086);
nor U19858 (N_19858,N_19304,N_19239);
and U19859 (N_19859,N_19165,N_19375);
nor U19860 (N_19860,N_19276,N_19236);
and U19861 (N_19861,N_19057,N_19072);
xor U19862 (N_19862,N_19195,N_19364);
and U19863 (N_19863,N_19433,N_19068);
nor U19864 (N_19864,N_19336,N_19001);
or U19865 (N_19865,N_19018,N_19412);
nand U19866 (N_19866,N_19113,N_19485);
nor U19867 (N_19867,N_19032,N_19163);
xnor U19868 (N_19868,N_19452,N_19002);
nand U19869 (N_19869,N_19305,N_19114);
and U19870 (N_19870,N_19002,N_19132);
nand U19871 (N_19871,N_19256,N_19126);
nor U19872 (N_19872,N_19172,N_19008);
nand U19873 (N_19873,N_19084,N_19274);
nand U19874 (N_19874,N_19433,N_19084);
nor U19875 (N_19875,N_19392,N_19216);
xor U19876 (N_19876,N_19082,N_19050);
or U19877 (N_19877,N_19010,N_19491);
xor U19878 (N_19878,N_19484,N_19397);
nor U19879 (N_19879,N_19379,N_19459);
and U19880 (N_19880,N_19256,N_19326);
xnor U19881 (N_19881,N_19193,N_19468);
nor U19882 (N_19882,N_19334,N_19376);
and U19883 (N_19883,N_19498,N_19304);
nand U19884 (N_19884,N_19473,N_19430);
or U19885 (N_19885,N_19475,N_19362);
or U19886 (N_19886,N_19182,N_19374);
nand U19887 (N_19887,N_19256,N_19433);
nor U19888 (N_19888,N_19060,N_19277);
nand U19889 (N_19889,N_19297,N_19184);
nor U19890 (N_19890,N_19355,N_19299);
and U19891 (N_19891,N_19211,N_19088);
and U19892 (N_19892,N_19434,N_19311);
nor U19893 (N_19893,N_19454,N_19386);
or U19894 (N_19894,N_19193,N_19170);
nor U19895 (N_19895,N_19375,N_19053);
nor U19896 (N_19896,N_19197,N_19461);
and U19897 (N_19897,N_19152,N_19333);
and U19898 (N_19898,N_19039,N_19154);
nand U19899 (N_19899,N_19196,N_19312);
nand U19900 (N_19900,N_19401,N_19107);
nor U19901 (N_19901,N_19025,N_19035);
xor U19902 (N_19902,N_19197,N_19339);
and U19903 (N_19903,N_19381,N_19017);
nand U19904 (N_19904,N_19010,N_19276);
nand U19905 (N_19905,N_19261,N_19489);
or U19906 (N_19906,N_19035,N_19337);
or U19907 (N_19907,N_19016,N_19230);
nor U19908 (N_19908,N_19111,N_19053);
or U19909 (N_19909,N_19160,N_19019);
nand U19910 (N_19910,N_19058,N_19119);
nor U19911 (N_19911,N_19158,N_19256);
nand U19912 (N_19912,N_19436,N_19091);
and U19913 (N_19913,N_19444,N_19176);
or U19914 (N_19914,N_19493,N_19424);
xnor U19915 (N_19915,N_19118,N_19153);
nand U19916 (N_19916,N_19306,N_19113);
nand U19917 (N_19917,N_19230,N_19173);
nor U19918 (N_19918,N_19056,N_19263);
xnor U19919 (N_19919,N_19241,N_19132);
or U19920 (N_19920,N_19078,N_19000);
nor U19921 (N_19921,N_19392,N_19370);
nor U19922 (N_19922,N_19099,N_19291);
and U19923 (N_19923,N_19464,N_19056);
nor U19924 (N_19924,N_19291,N_19329);
nor U19925 (N_19925,N_19319,N_19191);
nor U19926 (N_19926,N_19257,N_19295);
and U19927 (N_19927,N_19243,N_19396);
and U19928 (N_19928,N_19055,N_19211);
nand U19929 (N_19929,N_19334,N_19433);
xnor U19930 (N_19930,N_19131,N_19305);
and U19931 (N_19931,N_19381,N_19399);
and U19932 (N_19932,N_19464,N_19447);
or U19933 (N_19933,N_19344,N_19000);
xor U19934 (N_19934,N_19016,N_19382);
nand U19935 (N_19935,N_19193,N_19283);
xnor U19936 (N_19936,N_19325,N_19473);
and U19937 (N_19937,N_19424,N_19228);
or U19938 (N_19938,N_19207,N_19308);
nand U19939 (N_19939,N_19263,N_19271);
or U19940 (N_19940,N_19341,N_19469);
nand U19941 (N_19941,N_19495,N_19410);
and U19942 (N_19942,N_19261,N_19185);
and U19943 (N_19943,N_19096,N_19332);
nand U19944 (N_19944,N_19185,N_19028);
nor U19945 (N_19945,N_19316,N_19041);
or U19946 (N_19946,N_19214,N_19283);
nand U19947 (N_19947,N_19392,N_19157);
or U19948 (N_19948,N_19236,N_19308);
or U19949 (N_19949,N_19344,N_19354);
or U19950 (N_19950,N_19310,N_19017);
and U19951 (N_19951,N_19494,N_19400);
nand U19952 (N_19952,N_19243,N_19347);
and U19953 (N_19953,N_19470,N_19178);
nor U19954 (N_19954,N_19337,N_19108);
nand U19955 (N_19955,N_19105,N_19361);
and U19956 (N_19956,N_19196,N_19022);
or U19957 (N_19957,N_19470,N_19357);
and U19958 (N_19958,N_19462,N_19145);
xnor U19959 (N_19959,N_19030,N_19321);
nand U19960 (N_19960,N_19282,N_19250);
and U19961 (N_19961,N_19140,N_19476);
and U19962 (N_19962,N_19397,N_19285);
nor U19963 (N_19963,N_19454,N_19055);
or U19964 (N_19964,N_19117,N_19438);
nor U19965 (N_19965,N_19223,N_19049);
or U19966 (N_19966,N_19265,N_19484);
and U19967 (N_19967,N_19335,N_19286);
nor U19968 (N_19968,N_19328,N_19174);
nor U19969 (N_19969,N_19047,N_19416);
nor U19970 (N_19970,N_19438,N_19351);
or U19971 (N_19971,N_19378,N_19336);
and U19972 (N_19972,N_19331,N_19160);
nor U19973 (N_19973,N_19060,N_19311);
or U19974 (N_19974,N_19012,N_19067);
nand U19975 (N_19975,N_19095,N_19039);
or U19976 (N_19976,N_19388,N_19473);
nor U19977 (N_19977,N_19112,N_19455);
nand U19978 (N_19978,N_19085,N_19010);
or U19979 (N_19979,N_19492,N_19454);
nand U19980 (N_19980,N_19362,N_19024);
nand U19981 (N_19981,N_19474,N_19076);
nor U19982 (N_19982,N_19011,N_19427);
nor U19983 (N_19983,N_19056,N_19162);
nor U19984 (N_19984,N_19008,N_19035);
nor U19985 (N_19985,N_19304,N_19047);
or U19986 (N_19986,N_19188,N_19416);
nand U19987 (N_19987,N_19454,N_19351);
nor U19988 (N_19988,N_19406,N_19474);
nor U19989 (N_19989,N_19241,N_19491);
or U19990 (N_19990,N_19465,N_19467);
nor U19991 (N_19991,N_19463,N_19266);
nand U19992 (N_19992,N_19333,N_19034);
nand U19993 (N_19993,N_19385,N_19071);
nand U19994 (N_19994,N_19006,N_19211);
nand U19995 (N_19995,N_19412,N_19066);
nor U19996 (N_19996,N_19202,N_19185);
or U19997 (N_19997,N_19325,N_19033);
nand U19998 (N_19998,N_19068,N_19055);
nor U19999 (N_19999,N_19140,N_19050);
nand U20000 (N_20000,N_19582,N_19788);
and U20001 (N_20001,N_19577,N_19791);
nand U20002 (N_20002,N_19803,N_19517);
and U20003 (N_20003,N_19916,N_19544);
nor U20004 (N_20004,N_19618,N_19507);
or U20005 (N_20005,N_19718,N_19684);
and U20006 (N_20006,N_19580,N_19824);
nor U20007 (N_20007,N_19797,N_19874);
xnor U20008 (N_20008,N_19663,N_19866);
or U20009 (N_20009,N_19912,N_19595);
nor U20010 (N_20010,N_19514,N_19652);
xor U20011 (N_20011,N_19815,N_19597);
nor U20012 (N_20012,N_19699,N_19850);
nor U20013 (N_20013,N_19871,N_19957);
nand U20014 (N_20014,N_19536,N_19929);
nand U20015 (N_20015,N_19708,N_19800);
and U20016 (N_20016,N_19933,N_19660);
and U20017 (N_20017,N_19570,N_19711);
nand U20018 (N_20018,N_19845,N_19943);
nand U20019 (N_20019,N_19758,N_19503);
or U20020 (N_20020,N_19651,N_19804);
and U20021 (N_20021,N_19567,N_19986);
nand U20022 (N_20022,N_19885,N_19978);
and U20023 (N_20023,N_19913,N_19695);
and U20024 (N_20024,N_19639,N_19636);
and U20025 (N_20025,N_19873,N_19553);
or U20026 (N_20026,N_19673,N_19564);
or U20027 (N_20027,N_19576,N_19691);
nor U20028 (N_20028,N_19801,N_19883);
xnor U20029 (N_20029,N_19900,N_19920);
and U20030 (N_20030,N_19585,N_19715);
nor U20031 (N_20031,N_19759,N_19568);
nand U20032 (N_20032,N_19907,N_19949);
and U20033 (N_20033,N_19887,N_19525);
nand U20034 (N_20034,N_19702,N_19808);
xnor U20035 (N_20035,N_19821,N_19643);
nand U20036 (N_20036,N_19970,N_19980);
nor U20037 (N_20037,N_19653,N_19918);
xor U20038 (N_20038,N_19852,N_19705);
and U20039 (N_20039,N_19965,N_19543);
nand U20040 (N_20040,N_19640,N_19868);
nand U20041 (N_20041,N_19766,N_19898);
xor U20042 (N_20042,N_19964,N_19942);
or U20043 (N_20043,N_19825,N_19589);
and U20044 (N_20044,N_19784,N_19648);
nand U20045 (N_20045,N_19510,N_19529);
nor U20046 (N_20046,N_19823,N_19538);
nand U20047 (N_20047,N_19515,N_19554);
nand U20048 (N_20048,N_19927,N_19977);
nand U20049 (N_20049,N_19692,N_19952);
nand U20050 (N_20050,N_19841,N_19789);
nor U20051 (N_20051,N_19712,N_19528);
and U20052 (N_20052,N_19592,N_19926);
and U20053 (N_20053,N_19537,N_19765);
nor U20054 (N_20054,N_19574,N_19521);
or U20055 (N_20055,N_19723,N_19886);
and U20056 (N_20056,N_19550,N_19747);
nand U20057 (N_20057,N_19737,N_19869);
nor U20058 (N_20058,N_19971,N_19674);
and U20059 (N_20059,N_19552,N_19627);
nand U20060 (N_20060,N_19729,N_19625);
or U20061 (N_20061,N_19844,N_19843);
or U20062 (N_20062,N_19509,N_19511);
or U20063 (N_20063,N_19617,N_19901);
nand U20064 (N_20064,N_19624,N_19855);
nand U20065 (N_20065,N_19632,N_19995);
xor U20066 (N_20066,N_19603,N_19777);
and U20067 (N_20067,N_19689,N_19809);
and U20068 (N_20068,N_19559,N_19984);
nor U20069 (N_20069,N_19516,N_19608);
nor U20070 (N_20070,N_19778,N_19865);
nand U20071 (N_20071,N_19752,N_19798);
nand U20072 (N_20072,N_19602,N_19902);
and U20073 (N_20073,N_19631,N_19593);
xor U20074 (N_20074,N_19762,N_19744);
or U20075 (N_20075,N_19944,N_19967);
nor U20076 (N_20076,N_19523,N_19742);
and U20077 (N_20077,N_19542,N_19993);
nand U20078 (N_20078,N_19879,N_19807);
nor U20079 (N_20079,N_19892,N_19781);
nand U20080 (N_20080,N_19930,N_19761);
or U20081 (N_20081,N_19741,N_19650);
nand U20082 (N_20082,N_19601,N_19560);
or U20083 (N_20083,N_19915,N_19906);
and U20084 (N_20084,N_19796,N_19848);
or U20085 (N_20085,N_19730,N_19688);
or U20086 (N_20086,N_19579,N_19793);
nor U20087 (N_20087,N_19780,N_19513);
nand U20088 (N_20088,N_19861,N_19731);
nand U20089 (N_20089,N_19569,N_19740);
or U20090 (N_20090,N_19749,N_19502);
nand U20091 (N_20091,N_19769,N_19508);
nor U20092 (N_20092,N_19614,N_19551);
or U20093 (N_20093,N_19735,N_19520);
nand U20094 (N_20094,N_19996,N_19954);
or U20095 (N_20095,N_19700,N_19630);
and U20096 (N_20096,N_19754,N_19764);
nand U20097 (N_20097,N_19587,N_19909);
nor U20098 (N_20098,N_19903,N_19704);
nor U20099 (N_20099,N_19757,N_19732);
nor U20100 (N_20100,N_19615,N_19782);
xnor U20101 (N_20101,N_19896,N_19555);
and U20102 (N_20102,N_19535,N_19816);
nand U20103 (N_20103,N_19549,N_19904);
or U20104 (N_20104,N_19987,N_19541);
or U20105 (N_20105,N_19836,N_19586);
and U20106 (N_20106,N_19534,N_19829);
or U20107 (N_20107,N_19572,N_19713);
nor U20108 (N_20108,N_19561,N_19575);
xnor U20109 (N_20109,N_19505,N_19839);
nand U20110 (N_20110,N_19858,N_19908);
and U20111 (N_20111,N_19774,N_19972);
and U20112 (N_20112,N_19607,N_19533);
xor U20113 (N_20113,N_19610,N_19812);
and U20114 (N_20114,N_19760,N_19799);
nor U20115 (N_20115,N_19733,N_19745);
nor U20116 (N_20116,N_19786,N_19881);
xnor U20117 (N_20117,N_19714,N_19897);
and U20118 (N_20118,N_19539,N_19696);
and U20119 (N_20119,N_19657,N_19795);
nor U20120 (N_20120,N_19566,N_19746);
nand U20121 (N_20121,N_19690,N_19991);
and U20122 (N_20122,N_19600,N_19983);
nor U20123 (N_20123,N_19773,N_19724);
xor U20124 (N_20124,N_19728,N_19750);
and U20125 (N_20125,N_19783,N_19981);
nand U20126 (N_20126,N_19994,N_19756);
and U20127 (N_20127,N_19725,N_19857);
and U20128 (N_20128,N_19654,N_19706);
and U20129 (N_20129,N_19500,N_19719);
nor U20130 (N_20130,N_19669,N_19922);
and U20131 (N_20131,N_19522,N_19670);
nand U20132 (N_20132,N_19672,N_19936);
xnor U20133 (N_20133,N_19847,N_19755);
and U20134 (N_20134,N_19598,N_19665);
and U20135 (N_20135,N_19717,N_19666);
nor U20136 (N_20136,N_19644,N_19583);
nor U20137 (N_20137,N_19935,N_19557);
and U20138 (N_20138,N_19787,N_19504);
or U20139 (N_20139,N_19872,N_19968);
nor U20140 (N_20140,N_19751,N_19888);
nor U20141 (N_20141,N_19776,N_19634);
nor U20142 (N_20142,N_19882,N_19818);
and U20143 (N_20143,N_19679,N_19726);
or U20144 (N_20144,N_19932,N_19524);
xnor U20145 (N_20145,N_19707,N_19853);
and U20146 (N_20146,N_19681,N_19743);
nor U20147 (N_20147,N_19736,N_19846);
xnor U20148 (N_20148,N_19939,N_19709);
nand U20149 (N_20149,N_19802,N_19512);
nor U20150 (N_20150,N_19641,N_19581);
xnor U20151 (N_20151,N_19680,N_19842);
nand U20152 (N_20152,N_19924,N_19938);
nand U20153 (N_20153,N_19979,N_19734);
or U20154 (N_20154,N_19792,N_19588);
or U20155 (N_20155,N_19662,N_19739);
nor U20156 (N_20156,N_19671,N_19623);
and U20157 (N_20157,N_19697,N_19998);
or U20158 (N_20158,N_19558,N_19895);
or U20159 (N_20159,N_19710,N_19947);
nor U20160 (N_20160,N_19698,N_19638);
nor U20161 (N_20161,N_19794,N_19934);
nor U20162 (N_20162,N_19628,N_19738);
or U20163 (N_20163,N_19545,N_19540);
nor U20164 (N_20164,N_19772,N_19547);
nor U20165 (N_20165,N_19518,N_19941);
nor U20166 (N_20166,N_19775,N_19790);
xor U20167 (N_20167,N_19911,N_19822);
nor U20168 (N_20168,N_19826,N_19677);
and U20169 (N_20169,N_19830,N_19611);
and U20170 (N_20170,N_19890,N_19937);
xor U20171 (N_20171,N_19685,N_19876);
or U20172 (N_20172,N_19893,N_19622);
and U20173 (N_20173,N_19925,N_19661);
nor U20174 (N_20174,N_19950,N_19501);
and U20175 (N_20175,N_19584,N_19889);
nor U20176 (N_20176,N_19649,N_19974);
nor U20177 (N_20177,N_19838,N_19856);
or U20178 (N_20178,N_19849,N_19837);
xnor U20179 (N_20179,N_19571,N_19976);
nor U20180 (N_20180,N_19999,N_19633);
or U20181 (N_20181,N_19867,N_19767);
xnor U20182 (N_20182,N_19556,N_19526);
xor U20183 (N_20183,N_19716,N_19519);
nand U20184 (N_20184,N_19530,N_19806);
nor U20185 (N_20185,N_19870,N_19946);
nor U20186 (N_20186,N_19811,N_19621);
nor U20187 (N_20187,N_19693,N_19810);
nor U20188 (N_20188,N_19779,N_19686);
nand U20189 (N_20189,N_19721,N_19854);
nor U20190 (N_20190,N_19834,N_19616);
or U20191 (N_20191,N_19785,N_19763);
and U20192 (N_20192,N_19635,N_19619);
or U20193 (N_20193,N_19905,N_19646);
and U20194 (N_20194,N_19864,N_19833);
xnor U20195 (N_20195,N_19532,N_19928);
and U20196 (N_20196,N_19923,N_19959);
and U20197 (N_20197,N_19527,N_19722);
nor U20198 (N_20198,N_19596,N_19963);
or U20199 (N_20199,N_19813,N_19960);
nand U20200 (N_20200,N_19955,N_19990);
xnor U20201 (N_20201,N_19682,N_19546);
nand U20202 (N_20202,N_19817,N_19748);
xor U20203 (N_20203,N_19753,N_19832);
nand U20204 (N_20204,N_19720,N_19961);
nor U20205 (N_20205,N_19859,N_19770);
or U20206 (N_20206,N_19835,N_19884);
nor U20207 (N_20207,N_19629,N_19613);
nand U20208 (N_20208,N_19891,N_19771);
xor U20209 (N_20209,N_19814,N_19620);
and U20210 (N_20210,N_19703,N_19658);
nand U20211 (N_20211,N_19548,N_19768);
xnor U20212 (N_20212,N_19940,N_19594);
nor U20213 (N_20213,N_19962,N_19694);
nand U20214 (N_20214,N_19878,N_19951);
or U20215 (N_20215,N_19988,N_19659);
nor U20216 (N_20216,N_19678,N_19805);
or U20217 (N_20217,N_19851,N_19563);
or U20218 (N_20218,N_19919,N_19969);
nor U20219 (N_20219,N_19863,N_19626);
nand U20220 (N_20220,N_19668,N_19921);
nor U20221 (N_20221,N_19676,N_19578);
and U20222 (N_20222,N_19637,N_19860);
xnor U20223 (N_20223,N_19910,N_19831);
and U20224 (N_20224,N_19820,N_19875);
and U20225 (N_20225,N_19573,N_19562);
or U20226 (N_20226,N_19675,N_19727);
nand U20227 (N_20227,N_19958,N_19687);
nor U20228 (N_20228,N_19827,N_19609);
nand U20229 (N_20229,N_19828,N_19612);
nand U20230 (N_20230,N_19931,N_19606);
or U20231 (N_20231,N_19975,N_19591);
xor U20232 (N_20232,N_19590,N_19945);
nand U20233 (N_20233,N_19565,N_19683);
nand U20234 (N_20234,N_19506,N_19948);
and U20235 (N_20235,N_19701,N_19664);
and U20236 (N_20236,N_19605,N_19985);
xor U20237 (N_20237,N_19840,N_19645);
or U20238 (N_20238,N_19992,N_19862);
xor U20239 (N_20239,N_19894,N_19604);
and U20240 (N_20240,N_19997,N_19647);
and U20241 (N_20241,N_19642,N_19953);
and U20242 (N_20242,N_19982,N_19655);
nor U20243 (N_20243,N_19914,N_19956);
nor U20244 (N_20244,N_19877,N_19989);
nor U20245 (N_20245,N_19899,N_19917);
and U20246 (N_20246,N_19667,N_19880);
nor U20247 (N_20247,N_19819,N_19531);
nor U20248 (N_20248,N_19599,N_19966);
nor U20249 (N_20249,N_19973,N_19656);
nor U20250 (N_20250,N_19684,N_19701);
or U20251 (N_20251,N_19648,N_19633);
or U20252 (N_20252,N_19536,N_19768);
nand U20253 (N_20253,N_19683,N_19564);
nor U20254 (N_20254,N_19513,N_19649);
or U20255 (N_20255,N_19683,N_19771);
xor U20256 (N_20256,N_19627,N_19547);
and U20257 (N_20257,N_19838,N_19849);
or U20258 (N_20258,N_19567,N_19883);
nor U20259 (N_20259,N_19925,N_19618);
nand U20260 (N_20260,N_19500,N_19873);
or U20261 (N_20261,N_19570,N_19875);
nor U20262 (N_20262,N_19618,N_19754);
nand U20263 (N_20263,N_19541,N_19595);
or U20264 (N_20264,N_19966,N_19810);
or U20265 (N_20265,N_19747,N_19650);
and U20266 (N_20266,N_19898,N_19972);
nand U20267 (N_20267,N_19725,N_19894);
or U20268 (N_20268,N_19591,N_19521);
or U20269 (N_20269,N_19949,N_19806);
nor U20270 (N_20270,N_19793,N_19909);
or U20271 (N_20271,N_19580,N_19985);
nor U20272 (N_20272,N_19699,N_19884);
xnor U20273 (N_20273,N_19726,N_19688);
nor U20274 (N_20274,N_19660,N_19733);
or U20275 (N_20275,N_19809,N_19990);
or U20276 (N_20276,N_19721,N_19820);
or U20277 (N_20277,N_19981,N_19900);
nand U20278 (N_20278,N_19936,N_19725);
or U20279 (N_20279,N_19560,N_19827);
and U20280 (N_20280,N_19643,N_19885);
nand U20281 (N_20281,N_19951,N_19710);
nand U20282 (N_20282,N_19919,N_19692);
xnor U20283 (N_20283,N_19846,N_19956);
nor U20284 (N_20284,N_19821,N_19581);
and U20285 (N_20285,N_19601,N_19838);
nor U20286 (N_20286,N_19763,N_19581);
and U20287 (N_20287,N_19713,N_19745);
and U20288 (N_20288,N_19632,N_19624);
xnor U20289 (N_20289,N_19678,N_19954);
and U20290 (N_20290,N_19556,N_19552);
nor U20291 (N_20291,N_19645,N_19934);
nor U20292 (N_20292,N_19859,N_19532);
nand U20293 (N_20293,N_19964,N_19842);
nor U20294 (N_20294,N_19686,N_19711);
or U20295 (N_20295,N_19579,N_19833);
nor U20296 (N_20296,N_19533,N_19887);
and U20297 (N_20297,N_19918,N_19628);
nand U20298 (N_20298,N_19669,N_19738);
or U20299 (N_20299,N_19729,N_19615);
or U20300 (N_20300,N_19601,N_19807);
nor U20301 (N_20301,N_19949,N_19947);
and U20302 (N_20302,N_19825,N_19889);
nand U20303 (N_20303,N_19920,N_19927);
and U20304 (N_20304,N_19503,N_19822);
nand U20305 (N_20305,N_19993,N_19817);
nor U20306 (N_20306,N_19920,N_19912);
or U20307 (N_20307,N_19878,N_19858);
nand U20308 (N_20308,N_19778,N_19797);
xnor U20309 (N_20309,N_19951,N_19520);
and U20310 (N_20310,N_19773,N_19728);
and U20311 (N_20311,N_19555,N_19969);
nand U20312 (N_20312,N_19841,N_19628);
nor U20313 (N_20313,N_19898,N_19792);
nand U20314 (N_20314,N_19707,N_19570);
and U20315 (N_20315,N_19641,N_19611);
or U20316 (N_20316,N_19961,N_19951);
nand U20317 (N_20317,N_19714,N_19604);
or U20318 (N_20318,N_19968,N_19917);
nand U20319 (N_20319,N_19632,N_19654);
or U20320 (N_20320,N_19888,N_19737);
nand U20321 (N_20321,N_19560,N_19619);
xnor U20322 (N_20322,N_19723,N_19633);
and U20323 (N_20323,N_19583,N_19833);
nor U20324 (N_20324,N_19763,N_19764);
nand U20325 (N_20325,N_19977,N_19759);
or U20326 (N_20326,N_19911,N_19999);
nand U20327 (N_20327,N_19799,N_19639);
and U20328 (N_20328,N_19721,N_19944);
and U20329 (N_20329,N_19628,N_19922);
and U20330 (N_20330,N_19501,N_19554);
or U20331 (N_20331,N_19592,N_19652);
nor U20332 (N_20332,N_19920,N_19803);
or U20333 (N_20333,N_19723,N_19715);
nand U20334 (N_20334,N_19910,N_19601);
nand U20335 (N_20335,N_19994,N_19563);
nand U20336 (N_20336,N_19557,N_19891);
or U20337 (N_20337,N_19786,N_19787);
nand U20338 (N_20338,N_19688,N_19773);
nor U20339 (N_20339,N_19917,N_19588);
or U20340 (N_20340,N_19913,N_19706);
or U20341 (N_20341,N_19543,N_19510);
nand U20342 (N_20342,N_19972,N_19648);
and U20343 (N_20343,N_19891,N_19816);
or U20344 (N_20344,N_19775,N_19523);
xnor U20345 (N_20345,N_19633,N_19541);
or U20346 (N_20346,N_19756,N_19638);
xnor U20347 (N_20347,N_19731,N_19728);
nor U20348 (N_20348,N_19771,N_19659);
nor U20349 (N_20349,N_19591,N_19982);
nor U20350 (N_20350,N_19672,N_19650);
or U20351 (N_20351,N_19595,N_19708);
nand U20352 (N_20352,N_19566,N_19838);
nor U20353 (N_20353,N_19816,N_19949);
or U20354 (N_20354,N_19987,N_19705);
and U20355 (N_20355,N_19612,N_19662);
nor U20356 (N_20356,N_19595,N_19582);
nand U20357 (N_20357,N_19721,N_19740);
or U20358 (N_20358,N_19639,N_19510);
xor U20359 (N_20359,N_19583,N_19762);
and U20360 (N_20360,N_19534,N_19806);
xor U20361 (N_20361,N_19583,N_19704);
nor U20362 (N_20362,N_19985,N_19701);
nor U20363 (N_20363,N_19603,N_19651);
xnor U20364 (N_20364,N_19608,N_19603);
and U20365 (N_20365,N_19858,N_19505);
nor U20366 (N_20366,N_19575,N_19560);
or U20367 (N_20367,N_19968,N_19992);
or U20368 (N_20368,N_19948,N_19988);
or U20369 (N_20369,N_19970,N_19969);
nand U20370 (N_20370,N_19668,N_19948);
and U20371 (N_20371,N_19838,N_19604);
or U20372 (N_20372,N_19887,N_19736);
nor U20373 (N_20373,N_19554,N_19758);
and U20374 (N_20374,N_19818,N_19536);
nor U20375 (N_20375,N_19925,N_19603);
nand U20376 (N_20376,N_19573,N_19502);
or U20377 (N_20377,N_19848,N_19787);
xor U20378 (N_20378,N_19558,N_19729);
nand U20379 (N_20379,N_19812,N_19622);
or U20380 (N_20380,N_19613,N_19897);
and U20381 (N_20381,N_19895,N_19938);
and U20382 (N_20382,N_19910,N_19797);
and U20383 (N_20383,N_19997,N_19648);
and U20384 (N_20384,N_19666,N_19889);
or U20385 (N_20385,N_19531,N_19558);
and U20386 (N_20386,N_19777,N_19650);
nand U20387 (N_20387,N_19681,N_19573);
and U20388 (N_20388,N_19803,N_19922);
or U20389 (N_20389,N_19965,N_19533);
nand U20390 (N_20390,N_19694,N_19625);
and U20391 (N_20391,N_19618,N_19667);
or U20392 (N_20392,N_19939,N_19877);
or U20393 (N_20393,N_19762,N_19592);
and U20394 (N_20394,N_19739,N_19957);
nor U20395 (N_20395,N_19988,N_19880);
nor U20396 (N_20396,N_19531,N_19721);
nor U20397 (N_20397,N_19657,N_19983);
or U20398 (N_20398,N_19852,N_19567);
nand U20399 (N_20399,N_19529,N_19936);
xor U20400 (N_20400,N_19965,N_19641);
and U20401 (N_20401,N_19685,N_19647);
nand U20402 (N_20402,N_19557,N_19744);
or U20403 (N_20403,N_19569,N_19731);
nor U20404 (N_20404,N_19587,N_19919);
nand U20405 (N_20405,N_19751,N_19826);
nor U20406 (N_20406,N_19729,N_19698);
xor U20407 (N_20407,N_19920,N_19517);
and U20408 (N_20408,N_19850,N_19511);
or U20409 (N_20409,N_19754,N_19969);
nor U20410 (N_20410,N_19993,N_19688);
nand U20411 (N_20411,N_19693,N_19644);
or U20412 (N_20412,N_19987,N_19998);
or U20413 (N_20413,N_19647,N_19696);
nor U20414 (N_20414,N_19729,N_19824);
nand U20415 (N_20415,N_19727,N_19538);
nor U20416 (N_20416,N_19574,N_19674);
nor U20417 (N_20417,N_19755,N_19818);
or U20418 (N_20418,N_19738,N_19773);
nor U20419 (N_20419,N_19842,N_19987);
and U20420 (N_20420,N_19695,N_19907);
nand U20421 (N_20421,N_19822,N_19930);
nor U20422 (N_20422,N_19878,N_19587);
or U20423 (N_20423,N_19964,N_19928);
or U20424 (N_20424,N_19755,N_19614);
and U20425 (N_20425,N_19933,N_19501);
or U20426 (N_20426,N_19777,N_19614);
or U20427 (N_20427,N_19854,N_19749);
and U20428 (N_20428,N_19644,N_19789);
and U20429 (N_20429,N_19688,N_19738);
nor U20430 (N_20430,N_19793,N_19808);
nor U20431 (N_20431,N_19828,N_19785);
xnor U20432 (N_20432,N_19585,N_19665);
nand U20433 (N_20433,N_19989,N_19592);
nand U20434 (N_20434,N_19781,N_19991);
or U20435 (N_20435,N_19995,N_19598);
nor U20436 (N_20436,N_19980,N_19558);
nand U20437 (N_20437,N_19511,N_19526);
or U20438 (N_20438,N_19760,N_19652);
or U20439 (N_20439,N_19518,N_19568);
xor U20440 (N_20440,N_19807,N_19912);
xnor U20441 (N_20441,N_19935,N_19881);
and U20442 (N_20442,N_19663,N_19737);
or U20443 (N_20443,N_19739,N_19524);
nor U20444 (N_20444,N_19600,N_19971);
and U20445 (N_20445,N_19663,N_19555);
or U20446 (N_20446,N_19962,N_19566);
and U20447 (N_20447,N_19687,N_19816);
nand U20448 (N_20448,N_19872,N_19610);
nand U20449 (N_20449,N_19921,N_19646);
or U20450 (N_20450,N_19590,N_19760);
nand U20451 (N_20451,N_19741,N_19546);
nand U20452 (N_20452,N_19926,N_19896);
nand U20453 (N_20453,N_19713,N_19621);
nand U20454 (N_20454,N_19941,N_19744);
or U20455 (N_20455,N_19835,N_19999);
and U20456 (N_20456,N_19977,N_19656);
or U20457 (N_20457,N_19791,N_19688);
and U20458 (N_20458,N_19618,N_19505);
nand U20459 (N_20459,N_19967,N_19549);
or U20460 (N_20460,N_19823,N_19793);
xor U20461 (N_20461,N_19661,N_19621);
xnor U20462 (N_20462,N_19648,N_19637);
nor U20463 (N_20463,N_19931,N_19867);
xnor U20464 (N_20464,N_19777,N_19651);
or U20465 (N_20465,N_19959,N_19577);
or U20466 (N_20466,N_19815,N_19779);
and U20467 (N_20467,N_19795,N_19968);
and U20468 (N_20468,N_19720,N_19797);
nor U20469 (N_20469,N_19561,N_19750);
nand U20470 (N_20470,N_19871,N_19573);
xor U20471 (N_20471,N_19924,N_19839);
nor U20472 (N_20472,N_19585,N_19743);
nor U20473 (N_20473,N_19909,N_19749);
nand U20474 (N_20474,N_19779,N_19871);
nand U20475 (N_20475,N_19506,N_19704);
nor U20476 (N_20476,N_19513,N_19800);
nand U20477 (N_20477,N_19635,N_19656);
xnor U20478 (N_20478,N_19706,N_19898);
and U20479 (N_20479,N_19840,N_19987);
and U20480 (N_20480,N_19746,N_19957);
or U20481 (N_20481,N_19740,N_19930);
and U20482 (N_20482,N_19842,N_19734);
nand U20483 (N_20483,N_19625,N_19990);
nor U20484 (N_20484,N_19535,N_19748);
nor U20485 (N_20485,N_19624,N_19808);
and U20486 (N_20486,N_19728,N_19991);
or U20487 (N_20487,N_19954,N_19581);
nand U20488 (N_20488,N_19971,N_19957);
and U20489 (N_20489,N_19678,N_19781);
nand U20490 (N_20490,N_19874,N_19628);
nor U20491 (N_20491,N_19656,N_19724);
xnor U20492 (N_20492,N_19793,N_19876);
and U20493 (N_20493,N_19558,N_19795);
and U20494 (N_20494,N_19544,N_19583);
or U20495 (N_20495,N_19885,N_19670);
and U20496 (N_20496,N_19538,N_19984);
or U20497 (N_20497,N_19579,N_19874);
nand U20498 (N_20498,N_19879,N_19752);
nand U20499 (N_20499,N_19527,N_19980);
nor U20500 (N_20500,N_20274,N_20097);
nor U20501 (N_20501,N_20071,N_20253);
nand U20502 (N_20502,N_20114,N_20178);
xor U20503 (N_20503,N_20399,N_20403);
or U20504 (N_20504,N_20009,N_20112);
and U20505 (N_20505,N_20383,N_20461);
xnor U20506 (N_20506,N_20139,N_20368);
or U20507 (N_20507,N_20470,N_20280);
and U20508 (N_20508,N_20268,N_20294);
nand U20509 (N_20509,N_20472,N_20485);
nand U20510 (N_20510,N_20207,N_20180);
nand U20511 (N_20511,N_20254,N_20035);
and U20512 (N_20512,N_20282,N_20323);
and U20513 (N_20513,N_20025,N_20275);
and U20514 (N_20514,N_20499,N_20435);
nand U20515 (N_20515,N_20482,N_20101);
and U20516 (N_20516,N_20169,N_20445);
or U20517 (N_20517,N_20456,N_20020);
and U20518 (N_20518,N_20128,N_20135);
or U20519 (N_20519,N_20251,N_20070);
nand U20520 (N_20520,N_20372,N_20428);
or U20521 (N_20521,N_20286,N_20444);
nand U20522 (N_20522,N_20492,N_20170);
nor U20523 (N_20523,N_20099,N_20134);
nand U20524 (N_20524,N_20050,N_20091);
and U20525 (N_20525,N_20053,N_20148);
and U20526 (N_20526,N_20182,N_20193);
nand U20527 (N_20527,N_20183,N_20033);
nand U20528 (N_20528,N_20156,N_20350);
xnor U20529 (N_20529,N_20455,N_20118);
xor U20530 (N_20530,N_20476,N_20332);
and U20531 (N_20531,N_20162,N_20015);
or U20532 (N_20532,N_20116,N_20073);
and U20533 (N_20533,N_20326,N_20493);
xor U20534 (N_20534,N_20259,N_20256);
nor U20535 (N_20535,N_20096,N_20481);
and U20536 (N_20536,N_20283,N_20122);
nand U20537 (N_20537,N_20154,N_20242);
and U20538 (N_20538,N_20055,N_20415);
and U20539 (N_20539,N_20315,N_20329);
or U20540 (N_20540,N_20152,N_20266);
nor U20541 (N_20541,N_20318,N_20407);
nand U20542 (N_20542,N_20382,N_20367);
nand U20543 (N_20543,N_20325,N_20001);
or U20544 (N_20544,N_20489,N_20413);
or U20545 (N_20545,N_20414,N_20230);
nand U20546 (N_20546,N_20363,N_20362);
nor U20547 (N_20547,N_20390,N_20306);
nand U20548 (N_20548,N_20014,N_20199);
nand U20549 (N_20549,N_20276,N_20153);
and U20550 (N_20550,N_20297,N_20337);
nor U20551 (N_20551,N_20453,N_20303);
nor U20552 (N_20552,N_20342,N_20007);
and U20553 (N_20553,N_20124,N_20218);
nor U20554 (N_20554,N_20331,N_20175);
nand U20555 (N_20555,N_20227,N_20384);
or U20556 (N_20556,N_20141,N_20249);
nor U20557 (N_20557,N_20443,N_20203);
nor U20558 (N_20558,N_20345,N_20349);
nor U20559 (N_20559,N_20458,N_20496);
xor U20560 (N_20560,N_20217,N_20334);
and U20561 (N_20561,N_20396,N_20225);
and U20562 (N_20562,N_20474,N_20408);
nor U20563 (N_20563,N_20074,N_20471);
nor U20564 (N_20564,N_20209,N_20067);
nor U20565 (N_20565,N_20094,N_20158);
and U20566 (N_20566,N_20263,N_20281);
nand U20567 (N_20567,N_20163,N_20298);
or U20568 (N_20568,N_20048,N_20467);
and U20569 (N_20569,N_20064,N_20108);
and U20570 (N_20570,N_20052,N_20075);
nand U20571 (N_20571,N_20495,N_20010);
or U20572 (N_20572,N_20236,N_20338);
nor U20573 (N_20573,N_20160,N_20082);
xor U20574 (N_20574,N_20023,N_20172);
nor U20575 (N_20575,N_20238,N_20400);
or U20576 (N_20576,N_20272,N_20173);
or U20577 (N_20577,N_20393,N_20340);
nor U20578 (N_20578,N_20054,N_20373);
nor U20579 (N_20579,N_20478,N_20296);
and U20580 (N_20580,N_20420,N_20189);
nand U20581 (N_20581,N_20464,N_20021);
and U20582 (N_20582,N_20061,N_20388);
or U20583 (N_20583,N_20235,N_20477);
and U20584 (N_20584,N_20410,N_20038);
nor U20585 (N_20585,N_20138,N_20398);
nor U20586 (N_20586,N_20127,N_20194);
nand U20587 (N_20587,N_20012,N_20140);
or U20588 (N_20588,N_20348,N_20098);
nand U20589 (N_20589,N_20335,N_20346);
and U20590 (N_20590,N_20125,N_20417);
xor U20591 (N_20591,N_20213,N_20198);
and U20592 (N_20592,N_20040,N_20279);
nand U20593 (N_20593,N_20111,N_20039);
or U20594 (N_20594,N_20095,N_20289);
or U20595 (N_20595,N_20299,N_20210);
nand U20596 (N_20596,N_20395,N_20191);
nor U20597 (N_20597,N_20089,N_20221);
or U20598 (N_20598,N_20231,N_20494);
nand U20599 (N_20599,N_20355,N_20257);
or U20600 (N_20600,N_20311,N_20484);
or U20601 (N_20601,N_20438,N_20295);
nand U20602 (N_20602,N_20437,N_20292);
nand U20603 (N_20603,N_20000,N_20186);
nor U20604 (N_20604,N_20145,N_20078);
and U20605 (N_20605,N_20404,N_20370);
nor U20606 (N_20606,N_20137,N_20196);
nor U20607 (N_20607,N_20214,N_20352);
nor U20608 (N_20608,N_20046,N_20327);
xnor U20609 (N_20609,N_20244,N_20265);
nand U20610 (N_20610,N_20245,N_20028);
and U20611 (N_20611,N_20416,N_20313);
nand U20612 (N_20612,N_20487,N_20226);
nor U20613 (N_20613,N_20387,N_20002);
nor U20614 (N_20614,N_20353,N_20376);
nand U20615 (N_20615,N_20460,N_20488);
nand U20616 (N_20616,N_20351,N_20117);
and U20617 (N_20617,N_20375,N_20320);
nand U20618 (N_20618,N_20463,N_20083);
nor U20619 (N_20619,N_20129,N_20284);
or U20620 (N_20620,N_20110,N_20239);
or U20621 (N_20621,N_20449,N_20109);
nand U20622 (N_20622,N_20465,N_20336);
or U20623 (N_20623,N_20392,N_20043);
nand U20624 (N_20624,N_20222,N_20219);
or U20625 (N_20625,N_20045,N_20439);
xnor U20626 (N_20626,N_20288,N_20146);
nor U20627 (N_20627,N_20149,N_20008);
or U20628 (N_20628,N_20309,N_20452);
nor U20629 (N_20629,N_20386,N_20079);
or U20630 (N_20630,N_20301,N_20005);
xor U20631 (N_20631,N_20041,N_20159);
or U20632 (N_20632,N_20243,N_20423);
nor U20633 (N_20633,N_20440,N_20076);
or U20634 (N_20634,N_20080,N_20252);
or U20635 (N_20635,N_20188,N_20308);
nand U20636 (N_20636,N_20013,N_20432);
or U20637 (N_20637,N_20267,N_20328);
nand U20638 (N_20638,N_20422,N_20291);
and U20639 (N_20639,N_20206,N_20365);
or U20640 (N_20640,N_20405,N_20446);
nor U20641 (N_20641,N_20434,N_20287);
nor U20642 (N_20642,N_20104,N_20229);
or U20643 (N_20643,N_20427,N_20107);
xnor U20644 (N_20644,N_20391,N_20459);
or U20645 (N_20645,N_20205,N_20237);
nand U20646 (N_20646,N_20174,N_20121);
nor U20647 (N_20647,N_20339,N_20072);
or U20648 (N_20648,N_20343,N_20319);
xor U20649 (N_20649,N_20269,N_20234);
and U20650 (N_20650,N_20171,N_20377);
and U20651 (N_20651,N_20321,N_20409);
xor U20652 (N_20652,N_20394,N_20441);
or U20653 (N_20653,N_20469,N_20113);
nor U20654 (N_20654,N_20360,N_20314);
or U20655 (N_20655,N_20442,N_20022);
or U20656 (N_20656,N_20077,N_20147);
and U20657 (N_20657,N_20016,N_20262);
nor U20658 (N_20658,N_20480,N_20497);
and U20659 (N_20659,N_20130,N_20034);
nor U20660 (N_20660,N_20371,N_20290);
nor U20661 (N_20661,N_20359,N_20255);
nor U20662 (N_20662,N_20019,N_20136);
nor U20663 (N_20663,N_20011,N_20240);
or U20664 (N_20664,N_20131,N_20086);
nand U20665 (N_20665,N_20277,N_20448);
nor U20666 (N_20666,N_20132,N_20241);
or U20667 (N_20667,N_20302,N_20233);
and U20668 (N_20668,N_20305,N_20151);
or U20669 (N_20669,N_20032,N_20462);
or U20670 (N_20670,N_20150,N_20026);
xnor U20671 (N_20671,N_20167,N_20030);
or U20672 (N_20672,N_20181,N_20491);
nor U20673 (N_20673,N_20119,N_20133);
and U20674 (N_20674,N_20100,N_20142);
or U20675 (N_20675,N_20184,N_20201);
and U20676 (N_20676,N_20300,N_20179);
nor U20677 (N_20677,N_20357,N_20278);
nor U20678 (N_20678,N_20258,N_20411);
and U20679 (N_20679,N_20081,N_20304);
nor U20680 (N_20680,N_20216,N_20211);
nand U20681 (N_20681,N_20450,N_20044);
nor U20682 (N_20682,N_20475,N_20168);
nand U20683 (N_20683,N_20029,N_20264);
and U20684 (N_20684,N_20115,N_20224);
and U20685 (N_20685,N_20483,N_20058);
nand U20686 (N_20686,N_20068,N_20424);
nand U20687 (N_20687,N_20195,N_20389);
or U20688 (N_20688,N_20215,N_20364);
nand U20689 (N_20689,N_20406,N_20164);
xnor U20690 (N_20690,N_20027,N_20322);
or U20691 (N_20691,N_20333,N_20358);
nor U20692 (N_20692,N_20024,N_20063);
nand U20693 (N_20693,N_20316,N_20317);
and U20694 (N_20694,N_20378,N_20347);
or U20695 (N_20695,N_20202,N_20473);
and U20696 (N_20696,N_20004,N_20246);
and U20697 (N_20697,N_20426,N_20085);
nand U20698 (N_20698,N_20385,N_20093);
or U20699 (N_20699,N_20451,N_20056);
nand U20700 (N_20700,N_20307,N_20155);
nor U20701 (N_20701,N_20069,N_20223);
nor U20702 (N_20702,N_20143,N_20466);
or U20703 (N_20703,N_20105,N_20436);
xor U20704 (N_20704,N_20042,N_20017);
nor U20705 (N_20705,N_20062,N_20192);
and U20706 (N_20706,N_20379,N_20165);
nor U20707 (N_20707,N_20006,N_20065);
xor U20708 (N_20708,N_20247,N_20312);
nand U20709 (N_20709,N_20176,N_20431);
and U20710 (N_20710,N_20421,N_20060);
nand U20711 (N_20711,N_20090,N_20418);
nand U20712 (N_20712,N_20273,N_20103);
xor U20713 (N_20713,N_20057,N_20447);
or U20714 (N_20714,N_20433,N_20228);
and U20715 (N_20715,N_20250,N_20261);
nor U20716 (N_20716,N_20106,N_20047);
nor U20717 (N_20717,N_20344,N_20324);
xnor U20718 (N_20718,N_20037,N_20285);
nand U20719 (N_20719,N_20049,N_20397);
and U20720 (N_20720,N_20157,N_20341);
or U20721 (N_20721,N_20208,N_20092);
nand U20722 (N_20722,N_20271,N_20051);
and U20723 (N_20723,N_20468,N_20479);
nor U20724 (N_20724,N_20380,N_20270);
nor U20725 (N_20725,N_20425,N_20486);
and U20726 (N_20726,N_20084,N_20361);
or U20727 (N_20727,N_20204,N_20356);
or U20728 (N_20728,N_20369,N_20454);
nand U20729 (N_20729,N_20457,N_20036);
and U20730 (N_20730,N_20087,N_20401);
nand U20731 (N_20731,N_20166,N_20366);
nand U20732 (N_20732,N_20429,N_20031);
and U20733 (N_20733,N_20066,N_20187);
and U20734 (N_20734,N_20260,N_20293);
nor U20735 (N_20735,N_20102,N_20381);
or U20736 (N_20736,N_20354,N_20212);
nor U20737 (N_20737,N_20220,N_20200);
or U20738 (N_20738,N_20185,N_20088);
nand U20739 (N_20739,N_20374,N_20232);
and U20740 (N_20740,N_20197,N_20490);
nand U20741 (N_20741,N_20144,N_20120);
xor U20742 (N_20742,N_20402,N_20190);
xnor U20743 (N_20743,N_20177,N_20126);
or U20744 (N_20744,N_20161,N_20310);
nand U20745 (N_20745,N_20018,N_20430);
nor U20746 (N_20746,N_20412,N_20003);
nand U20747 (N_20747,N_20248,N_20059);
and U20748 (N_20748,N_20419,N_20330);
nor U20749 (N_20749,N_20123,N_20498);
or U20750 (N_20750,N_20198,N_20376);
nand U20751 (N_20751,N_20124,N_20150);
or U20752 (N_20752,N_20065,N_20252);
or U20753 (N_20753,N_20097,N_20279);
and U20754 (N_20754,N_20051,N_20114);
nor U20755 (N_20755,N_20223,N_20428);
xnor U20756 (N_20756,N_20417,N_20197);
nand U20757 (N_20757,N_20112,N_20164);
xnor U20758 (N_20758,N_20105,N_20319);
nor U20759 (N_20759,N_20027,N_20252);
and U20760 (N_20760,N_20471,N_20344);
or U20761 (N_20761,N_20202,N_20137);
or U20762 (N_20762,N_20257,N_20466);
or U20763 (N_20763,N_20027,N_20324);
nor U20764 (N_20764,N_20220,N_20449);
or U20765 (N_20765,N_20424,N_20098);
nor U20766 (N_20766,N_20162,N_20157);
nor U20767 (N_20767,N_20452,N_20378);
or U20768 (N_20768,N_20299,N_20296);
nor U20769 (N_20769,N_20491,N_20054);
and U20770 (N_20770,N_20346,N_20487);
and U20771 (N_20771,N_20386,N_20365);
and U20772 (N_20772,N_20043,N_20449);
or U20773 (N_20773,N_20288,N_20339);
and U20774 (N_20774,N_20041,N_20382);
nand U20775 (N_20775,N_20008,N_20069);
nand U20776 (N_20776,N_20352,N_20205);
and U20777 (N_20777,N_20344,N_20251);
or U20778 (N_20778,N_20137,N_20004);
xor U20779 (N_20779,N_20474,N_20021);
and U20780 (N_20780,N_20267,N_20346);
and U20781 (N_20781,N_20494,N_20421);
nand U20782 (N_20782,N_20494,N_20430);
nor U20783 (N_20783,N_20034,N_20030);
nor U20784 (N_20784,N_20054,N_20343);
or U20785 (N_20785,N_20407,N_20169);
nand U20786 (N_20786,N_20212,N_20363);
or U20787 (N_20787,N_20133,N_20163);
nand U20788 (N_20788,N_20228,N_20245);
nor U20789 (N_20789,N_20345,N_20333);
nand U20790 (N_20790,N_20068,N_20273);
nand U20791 (N_20791,N_20251,N_20417);
nand U20792 (N_20792,N_20227,N_20201);
and U20793 (N_20793,N_20254,N_20328);
xnor U20794 (N_20794,N_20381,N_20084);
and U20795 (N_20795,N_20197,N_20481);
or U20796 (N_20796,N_20375,N_20154);
or U20797 (N_20797,N_20431,N_20257);
or U20798 (N_20798,N_20066,N_20475);
and U20799 (N_20799,N_20480,N_20142);
xnor U20800 (N_20800,N_20389,N_20308);
nor U20801 (N_20801,N_20360,N_20282);
or U20802 (N_20802,N_20463,N_20337);
or U20803 (N_20803,N_20321,N_20019);
and U20804 (N_20804,N_20251,N_20293);
nor U20805 (N_20805,N_20149,N_20330);
and U20806 (N_20806,N_20341,N_20227);
and U20807 (N_20807,N_20002,N_20364);
xnor U20808 (N_20808,N_20453,N_20022);
nand U20809 (N_20809,N_20344,N_20104);
or U20810 (N_20810,N_20462,N_20063);
and U20811 (N_20811,N_20456,N_20380);
nor U20812 (N_20812,N_20252,N_20160);
or U20813 (N_20813,N_20072,N_20325);
nor U20814 (N_20814,N_20350,N_20348);
and U20815 (N_20815,N_20248,N_20221);
or U20816 (N_20816,N_20347,N_20034);
nor U20817 (N_20817,N_20169,N_20082);
nand U20818 (N_20818,N_20349,N_20483);
and U20819 (N_20819,N_20196,N_20041);
or U20820 (N_20820,N_20421,N_20185);
and U20821 (N_20821,N_20498,N_20154);
nor U20822 (N_20822,N_20287,N_20205);
or U20823 (N_20823,N_20280,N_20482);
xnor U20824 (N_20824,N_20038,N_20402);
xnor U20825 (N_20825,N_20225,N_20480);
xnor U20826 (N_20826,N_20013,N_20093);
xnor U20827 (N_20827,N_20263,N_20109);
nor U20828 (N_20828,N_20022,N_20302);
or U20829 (N_20829,N_20080,N_20098);
nor U20830 (N_20830,N_20353,N_20181);
nand U20831 (N_20831,N_20478,N_20408);
nand U20832 (N_20832,N_20262,N_20188);
or U20833 (N_20833,N_20005,N_20303);
and U20834 (N_20834,N_20192,N_20346);
or U20835 (N_20835,N_20257,N_20472);
and U20836 (N_20836,N_20078,N_20012);
nand U20837 (N_20837,N_20277,N_20167);
xor U20838 (N_20838,N_20193,N_20253);
or U20839 (N_20839,N_20244,N_20474);
or U20840 (N_20840,N_20337,N_20128);
nor U20841 (N_20841,N_20178,N_20437);
and U20842 (N_20842,N_20302,N_20010);
nor U20843 (N_20843,N_20225,N_20403);
and U20844 (N_20844,N_20491,N_20084);
nand U20845 (N_20845,N_20052,N_20454);
and U20846 (N_20846,N_20378,N_20142);
nor U20847 (N_20847,N_20089,N_20127);
and U20848 (N_20848,N_20015,N_20274);
nand U20849 (N_20849,N_20486,N_20205);
or U20850 (N_20850,N_20260,N_20265);
or U20851 (N_20851,N_20004,N_20473);
or U20852 (N_20852,N_20040,N_20372);
nor U20853 (N_20853,N_20135,N_20102);
or U20854 (N_20854,N_20470,N_20373);
and U20855 (N_20855,N_20425,N_20277);
and U20856 (N_20856,N_20174,N_20468);
or U20857 (N_20857,N_20003,N_20273);
nand U20858 (N_20858,N_20394,N_20457);
xnor U20859 (N_20859,N_20456,N_20385);
nor U20860 (N_20860,N_20331,N_20309);
xor U20861 (N_20861,N_20477,N_20027);
nor U20862 (N_20862,N_20123,N_20031);
nand U20863 (N_20863,N_20390,N_20022);
nand U20864 (N_20864,N_20110,N_20296);
and U20865 (N_20865,N_20213,N_20062);
or U20866 (N_20866,N_20070,N_20174);
nor U20867 (N_20867,N_20419,N_20484);
and U20868 (N_20868,N_20182,N_20479);
nand U20869 (N_20869,N_20107,N_20358);
and U20870 (N_20870,N_20177,N_20123);
nand U20871 (N_20871,N_20404,N_20142);
nand U20872 (N_20872,N_20456,N_20137);
nor U20873 (N_20873,N_20356,N_20240);
and U20874 (N_20874,N_20398,N_20233);
or U20875 (N_20875,N_20047,N_20276);
and U20876 (N_20876,N_20171,N_20297);
nand U20877 (N_20877,N_20065,N_20472);
nor U20878 (N_20878,N_20378,N_20416);
or U20879 (N_20879,N_20108,N_20295);
or U20880 (N_20880,N_20439,N_20414);
nor U20881 (N_20881,N_20219,N_20189);
nand U20882 (N_20882,N_20496,N_20276);
nor U20883 (N_20883,N_20194,N_20313);
xor U20884 (N_20884,N_20443,N_20305);
or U20885 (N_20885,N_20319,N_20430);
and U20886 (N_20886,N_20312,N_20288);
nor U20887 (N_20887,N_20076,N_20390);
nand U20888 (N_20888,N_20441,N_20465);
nand U20889 (N_20889,N_20208,N_20094);
nand U20890 (N_20890,N_20462,N_20095);
and U20891 (N_20891,N_20090,N_20013);
nand U20892 (N_20892,N_20472,N_20197);
nor U20893 (N_20893,N_20393,N_20352);
nor U20894 (N_20894,N_20287,N_20029);
or U20895 (N_20895,N_20058,N_20321);
nand U20896 (N_20896,N_20056,N_20425);
xor U20897 (N_20897,N_20353,N_20324);
nor U20898 (N_20898,N_20223,N_20140);
and U20899 (N_20899,N_20257,N_20258);
and U20900 (N_20900,N_20130,N_20310);
nor U20901 (N_20901,N_20077,N_20257);
nor U20902 (N_20902,N_20031,N_20387);
and U20903 (N_20903,N_20208,N_20488);
nand U20904 (N_20904,N_20428,N_20014);
or U20905 (N_20905,N_20363,N_20488);
and U20906 (N_20906,N_20484,N_20061);
and U20907 (N_20907,N_20256,N_20239);
nand U20908 (N_20908,N_20088,N_20289);
or U20909 (N_20909,N_20450,N_20166);
or U20910 (N_20910,N_20070,N_20079);
nand U20911 (N_20911,N_20239,N_20397);
and U20912 (N_20912,N_20162,N_20371);
and U20913 (N_20913,N_20487,N_20097);
or U20914 (N_20914,N_20135,N_20409);
and U20915 (N_20915,N_20489,N_20377);
or U20916 (N_20916,N_20443,N_20299);
nand U20917 (N_20917,N_20238,N_20028);
and U20918 (N_20918,N_20367,N_20340);
or U20919 (N_20919,N_20389,N_20282);
or U20920 (N_20920,N_20350,N_20077);
and U20921 (N_20921,N_20449,N_20367);
nor U20922 (N_20922,N_20084,N_20118);
nand U20923 (N_20923,N_20087,N_20206);
or U20924 (N_20924,N_20193,N_20477);
nor U20925 (N_20925,N_20135,N_20468);
nor U20926 (N_20926,N_20386,N_20371);
nand U20927 (N_20927,N_20013,N_20278);
nor U20928 (N_20928,N_20071,N_20280);
or U20929 (N_20929,N_20089,N_20449);
nor U20930 (N_20930,N_20013,N_20055);
nand U20931 (N_20931,N_20450,N_20424);
nand U20932 (N_20932,N_20361,N_20370);
xor U20933 (N_20933,N_20442,N_20161);
or U20934 (N_20934,N_20035,N_20185);
nor U20935 (N_20935,N_20152,N_20491);
nor U20936 (N_20936,N_20171,N_20098);
or U20937 (N_20937,N_20225,N_20307);
and U20938 (N_20938,N_20062,N_20220);
or U20939 (N_20939,N_20105,N_20063);
nand U20940 (N_20940,N_20183,N_20462);
or U20941 (N_20941,N_20461,N_20376);
and U20942 (N_20942,N_20477,N_20119);
nor U20943 (N_20943,N_20014,N_20194);
nor U20944 (N_20944,N_20430,N_20104);
or U20945 (N_20945,N_20112,N_20111);
or U20946 (N_20946,N_20496,N_20232);
nor U20947 (N_20947,N_20347,N_20242);
nand U20948 (N_20948,N_20440,N_20130);
or U20949 (N_20949,N_20342,N_20319);
and U20950 (N_20950,N_20428,N_20397);
nor U20951 (N_20951,N_20138,N_20476);
or U20952 (N_20952,N_20145,N_20198);
and U20953 (N_20953,N_20108,N_20041);
and U20954 (N_20954,N_20499,N_20414);
nand U20955 (N_20955,N_20336,N_20004);
nand U20956 (N_20956,N_20214,N_20391);
and U20957 (N_20957,N_20123,N_20020);
nor U20958 (N_20958,N_20427,N_20452);
or U20959 (N_20959,N_20230,N_20309);
and U20960 (N_20960,N_20295,N_20144);
xnor U20961 (N_20961,N_20149,N_20351);
nand U20962 (N_20962,N_20343,N_20082);
or U20963 (N_20963,N_20323,N_20443);
nand U20964 (N_20964,N_20235,N_20042);
and U20965 (N_20965,N_20032,N_20202);
nand U20966 (N_20966,N_20214,N_20285);
nor U20967 (N_20967,N_20304,N_20025);
nand U20968 (N_20968,N_20465,N_20497);
nor U20969 (N_20969,N_20178,N_20452);
xor U20970 (N_20970,N_20349,N_20494);
nor U20971 (N_20971,N_20112,N_20385);
nand U20972 (N_20972,N_20472,N_20226);
and U20973 (N_20973,N_20201,N_20257);
nand U20974 (N_20974,N_20070,N_20493);
or U20975 (N_20975,N_20343,N_20435);
nand U20976 (N_20976,N_20296,N_20189);
nand U20977 (N_20977,N_20241,N_20384);
nand U20978 (N_20978,N_20272,N_20380);
and U20979 (N_20979,N_20088,N_20046);
and U20980 (N_20980,N_20469,N_20217);
nor U20981 (N_20981,N_20091,N_20270);
nand U20982 (N_20982,N_20252,N_20321);
nor U20983 (N_20983,N_20471,N_20297);
and U20984 (N_20984,N_20125,N_20171);
or U20985 (N_20985,N_20319,N_20405);
nand U20986 (N_20986,N_20440,N_20247);
nor U20987 (N_20987,N_20149,N_20217);
or U20988 (N_20988,N_20455,N_20157);
xor U20989 (N_20989,N_20057,N_20050);
nor U20990 (N_20990,N_20093,N_20154);
and U20991 (N_20991,N_20478,N_20041);
and U20992 (N_20992,N_20253,N_20314);
nor U20993 (N_20993,N_20272,N_20233);
or U20994 (N_20994,N_20010,N_20076);
nand U20995 (N_20995,N_20316,N_20239);
or U20996 (N_20996,N_20425,N_20120);
nand U20997 (N_20997,N_20146,N_20230);
nor U20998 (N_20998,N_20150,N_20022);
nor U20999 (N_20999,N_20217,N_20175);
and U21000 (N_21000,N_20715,N_20984);
nand U21001 (N_21001,N_20966,N_20864);
xor U21002 (N_21002,N_20595,N_20554);
and U21003 (N_21003,N_20996,N_20503);
or U21004 (N_21004,N_20939,N_20728);
and U21005 (N_21005,N_20985,N_20826);
nand U21006 (N_21006,N_20854,N_20981);
xnor U21007 (N_21007,N_20884,N_20776);
xor U21008 (N_21008,N_20899,N_20917);
or U21009 (N_21009,N_20798,N_20852);
or U21010 (N_21010,N_20875,N_20870);
or U21011 (N_21011,N_20581,N_20686);
nand U21012 (N_21012,N_20688,N_20518);
nor U21013 (N_21013,N_20646,N_20755);
and U21014 (N_21014,N_20820,N_20927);
nor U21015 (N_21015,N_20871,N_20703);
xor U21016 (N_21016,N_20598,N_20954);
nand U21017 (N_21017,N_20735,N_20658);
or U21018 (N_21018,N_20586,N_20922);
or U21019 (N_21019,N_20504,N_20987);
xor U21020 (N_21020,N_20788,N_20994);
or U21021 (N_21021,N_20670,N_20889);
and U21022 (N_21022,N_20748,N_20633);
and U21023 (N_21023,N_20969,N_20669);
and U21024 (N_21024,N_20746,N_20986);
nor U21025 (N_21025,N_20873,N_20695);
nor U21026 (N_21026,N_20578,N_20771);
nand U21027 (N_21027,N_20977,N_20766);
and U21028 (N_21028,N_20710,N_20804);
nand U21029 (N_21029,N_20759,N_20544);
nand U21030 (N_21030,N_20961,N_20550);
nor U21031 (N_21031,N_20713,N_20979);
or U21032 (N_21032,N_20543,N_20726);
or U21033 (N_21033,N_20835,N_20955);
nor U21034 (N_21034,N_20916,N_20747);
nor U21035 (N_21035,N_20973,N_20682);
or U21036 (N_21036,N_20823,N_20524);
xor U21037 (N_21037,N_20622,N_20529);
nor U21038 (N_21038,N_20563,N_20602);
nor U21039 (N_21039,N_20958,N_20806);
and U21040 (N_21040,N_20960,N_20509);
or U21041 (N_21041,N_20621,N_20729);
or U21042 (N_21042,N_20637,N_20991);
and U21043 (N_21043,N_20603,N_20894);
or U21044 (N_21044,N_20697,N_20600);
nor U21045 (N_21045,N_20962,N_20535);
nand U21046 (N_21046,N_20618,N_20664);
nand U21047 (N_21047,N_20877,N_20888);
nand U21048 (N_21048,N_20913,N_20858);
and U21049 (N_21049,N_20716,N_20723);
or U21050 (N_21050,N_20808,N_20549);
and U21051 (N_21051,N_20642,N_20860);
or U21052 (N_21052,N_20511,N_20721);
and U21053 (N_21053,N_20774,N_20878);
nand U21054 (N_21054,N_20588,N_20714);
nand U21055 (N_21055,N_20501,N_20972);
nand U21056 (N_21056,N_20677,N_20799);
nand U21057 (N_21057,N_20935,N_20886);
nor U21058 (N_21058,N_20515,N_20882);
nand U21059 (N_21059,N_20742,N_20575);
or U21060 (N_21060,N_20712,N_20900);
and U21061 (N_21061,N_20830,N_20690);
or U21062 (N_21062,N_20684,N_20946);
nor U21063 (N_21063,N_20626,N_20968);
and U21064 (N_21064,N_20532,N_20609);
nor U21065 (N_21065,N_20827,N_20567);
nor U21066 (N_21066,N_20767,N_20643);
xnor U21067 (N_21067,N_20657,N_20749);
nor U21068 (N_21068,N_20832,N_20615);
or U21069 (N_21069,N_20505,N_20665);
and U21070 (N_21070,N_20594,N_20980);
nor U21071 (N_21071,N_20560,N_20831);
or U21072 (N_21072,N_20592,N_20947);
and U21073 (N_21073,N_20660,N_20940);
nor U21074 (N_21074,N_20662,N_20542);
and U21075 (N_21075,N_20988,N_20949);
and U21076 (N_21076,N_20971,N_20925);
and U21077 (N_21077,N_20649,N_20627);
nand U21078 (N_21078,N_20739,N_20787);
nand U21079 (N_21079,N_20819,N_20537);
xor U21080 (N_21080,N_20920,N_20736);
nand U21081 (N_21081,N_20625,N_20890);
and U21082 (N_21082,N_20782,N_20693);
or U21083 (N_21083,N_20901,N_20601);
or U21084 (N_21084,N_20507,N_20815);
or U21085 (N_21085,N_20891,N_20751);
nor U21086 (N_21086,N_20704,N_20772);
nand U21087 (N_21087,N_20868,N_20573);
nor U21088 (N_21088,N_20585,N_20596);
nor U21089 (N_21089,N_20720,N_20841);
or U21090 (N_21090,N_20809,N_20647);
nand U21091 (N_21091,N_20789,N_20869);
and U21092 (N_21092,N_20803,N_20906);
or U21093 (N_21093,N_20508,N_20770);
and U21094 (N_21094,N_20895,N_20629);
xnor U21095 (N_21095,N_20692,N_20911);
or U21096 (N_21096,N_20941,N_20722);
nor U21097 (N_21097,N_20872,N_20967);
nor U21098 (N_21098,N_20502,N_20571);
and U21099 (N_21099,N_20879,N_20607);
and U21100 (N_21100,N_20671,N_20855);
or U21101 (N_21101,N_20593,N_20847);
nand U21102 (N_21102,N_20676,N_20956);
and U21103 (N_21103,N_20921,N_20564);
xor U21104 (N_21104,N_20517,N_20857);
and U21105 (N_21105,N_20661,N_20719);
nor U21106 (N_21106,N_20849,N_20597);
nand U21107 (N_21107,N_20942,N_20778);
and U21108 (N_21108,N_20853,N_20566);
nor U21109 (N_21109,N_20936,N_20863);
xor U21110 (N_21110,N_20689,N_20883);
or U21111 (N_21111,N_20975,N_20814);
nor U21112 (N_21112,N_20545,N_20839);
nor U21113 (N_21113,N_20699,N_20546);
or U21114 (N_21114,N_20978,N_20915);
nand U21115 (N_21115,N_20547,N_20737);
and U21116 (N_21116,N_20938,N_20659);
and U21117 (N_21117,N_20959,N_20928);
and U21118 (N_21118,N_20631,N_20711);
nor U21119 (N_21119,N_20738,N_20757);
nand U21120 (N_21120,N_20552,N_20848);
nor U21121 (N_21121,N_20687,N_20520);
and U21122 (N_21122,N_20612,N_20744);
and U21123 (N_21123,N_20796,N_20833);
nand U21124 (N_21124,N_20553,N_20800);
or U21125 (N_21125,N_20718,N_20702);
xnor U21126 (N_21126,N_20948,N_20812);
nand U21127 (N_21127,N_20707,N_20874);
nor U21128 (N_21128,N_20663,N_20666);
and U21129 (N_21129,N_20768,N_20574);
or U21130 (N_21130,N_20909,N_20732);
and U21131 (N_21131,N_20654,N_20912);
or U21132 (N_21132,N_20630,N_20565);
or U21133 (N_21133,N_20533,N_20865);
and U21134 (N_21134,N_20725,N_20953);
nand U21135 (N_21135,N_20807,N_20650);
nor U21136 (N_21136,N_20856,N_20569);
xnor U21137 (N_21137,N_20623,N_20777);
or U21138 (N_21138,N_20876,N_20580);
nor U21139 (N_21139,N_20816,N_20760);
nand U21140 (N_21140,N_20998,N_20965);
nand U21141 (N_21141,N_20606,N_20845);
nand U21142 (N_21142,N_20512,N_20608);
or U21143 (N_21143,N_20656,N_20951);
nand U21144 (N_21144,N_20634,N_20698);
and U21145 (N_21145,N_20817,N_20769);
nor U21146 (N_21146,N_20821,N_20577);
nor U21147 (N_21147,N_20842,N_20636);
or U21148 (N_21148,N_20616,N_20570);
nand U21149 (N_21149,N_20810,N_20793);
and U21150 (N_21150,N_20859,N_20558);
and U21151 (N_21151,N_20844,N_20785);
or U21152 (N_21152,N_20851,N_20582);
and U21153 (N_21153,N_20680,N_20651);
and U21154 (N_21154,N_20675,N_20648);
nor U21155 (N_21155,N_20526,N_20964);
and U21156 (N_21156,N_20786,N_20914);
nor U21157 (N_21157,N_20887,N_20758);
nand U21158 (N_21158,N_20624,N_20506);
nor U21159 (N_21159,N_20619,N_20898);
and U21160 (N_21160,N_20824,N_20705);
nor U21161 (N_21161,N_20668,N_20997);
or U21162 (N_21162,N_20773,N_20750);
xnor U21163 (N_21163,N_20933,N_20635);
nand U21164 (N_21164,N_20638,N_20620);
or U21165 (N_21165,N_20753,N_20811);
nand U21166 (N_21166,N_20640,N_20731);
xor U21167 (N_21167,N_20923,N_20893);
xor U21168 (N_21168,N_20937,N_20907);
nor U21169 (N_21169,N_20930,N_20797);
and U21170 (N_21170,N_20861,N_20926);
xnor U21171 (N_21171,N_20528,N_20934);
nand U21172 (N_21172,N_20822,N_20700);
and U21173 (N_21173,N_20963,N_20644);
and U21174 (N_21174,N_20613,N_20897);
and U21175 (N_21175,N_20999,N_20838);
nor U21176 (N_21176,N_20775,N_20694);
and U21177 (N_21177,N_20536,N_20673);
nand U21178 (N_21178,N_20674,N_20556);
and U21179 (N_21179,N_20557,N_20982);
nor U21180 (N_21180,N_20727,N_20599);
or U21181 (N_21181,N_20685,N_20896);
or U21182 (N_21182,N_20950,N_20611);
nor U21183 (N_21183,N_20783,N_20790);
nand U21184 (N_21184,N_20641,N_20829);
and U21185 (N_21185,N_20584,N_20579);
nor U21186 (N_21186,N_20763,N_20931);
nand U21187 (N_21187,N_20805,N_20678);
nand U21188 (N_21188,N_20919,N_20995);
and U21189 (N_21189,N_20840,N_20764);
nand U21190 (N_21190,N_20551,N_20706);
nor U21191 (N_21191,N_20681,N_20679);
nand U21192 (N_21192,N_20667,N_20880);
or U21193 (N_21193,N_20562,N_20541);
or U21194 (N_21194,N_20802,N_20780);
and U21195 (N_21195,N_20683,N_20514);
nor U21196 (N_21196,N_20743,N_20992);
nand U21197 (N_21197,N_20918,N_20614);
and U21198 (N_21198,N_20952,N_20867);
nor U21199 (N_21199,N_20583,N_20801);
nand U21200 (N_21200,N_20701,N_20752);
xor U21201 (N_21201,N_20741,N_20781);
xnor U21202 (N_21202,N_20945,N_20645);
and U21203 (N_21203,N_20510,N_20734);
nor U21204 (N_21204,N_20825,N_20795);
xnor U21205 (N_21205,N_20902,N_20572);
or U21206 (N_21206,N_20990,N_20850);
xor U21207 (N_21207,N_20655,N_20639);
nand U21208 (N_21208,N_20733,N_20730);
and U21209 (N_21209,N_20866,N_20500);
nand U21210 (N_21210,N_20754,N_20527);
nand U21211 (N_21211,N_20539,N_20970);
nor U21212 (N_21212,N_20779,N_20522);
nor U21213 (N_21213,N_20983,N_20904);
nor U21214 (N_21214,N_20837,N_20531);
nand U21215 (N_21215,N_20519,N_20653);
and U21216 (N_21216,N_20708,N_20910);
or U21217 (N_21217,N_20905,N_20709);
and U21218 (N_21218,N_20724,N_20836);
or U21219 (N_21219,N_20587,N_20559);
or U21220 (N_21220,N_20610,N_20993);
nand U21221 (N_21221,N_20604,N_20843);
or U21222 (N_21222,N_20976,N_20576);
or U21223 (N_21223,N_20892,N_20605);
nand U21224 (N_21224,N_20534,N_20765);
or U21225 (N_21225,N_20794,N_20828);
xnor U21226 (N_21226,N_20617,N_20791);
and U21227 (N_21227,N_20834,N_20513);
nor U21228 (N_21228,N_20944,N_20561);
nor U21229 (N_21229,N_20540,N_20974);
nor U21230 (N_21230,N_20523,N_20632);
and U21231 (N_21231,N_20908,N_20672);
nor U21232 (N_21232,N_20589,N_20516);
nand U21233 (N_21233,N_20792,N_20929);
and U21234 (N_21234,N_20521,N_20885);
or U21235 (N_21235,N_20548,N_20745);
and U21236 (N_21236,N_20740,N_20756);
and U21237 (N_21237,N_20696,N_20591);
and U21238 (N_21238,N_20761,N_20568);
nor U21239 (N_21239,N_20538,N_20932);
or U21240 (N_21240,N_20590,N_20846);
nand U21241 (N_21241,N_20943,N_20555);
and U21242 (N_21242,N_20530,N_20691);
nor U21243 (N_21243,N_20652,N_20762);
nor U21244 (N_21244,N_20862,N_20813);
and U21245 (N_21245,N_20525,N_20818);
nand U21246 (N_21246,N_20784,N_20989);
xnor U21247 (N_21247,N_20957,N_20881);
nand U21248 (N_21248,N_20924,N_20628);
nand U21249 (N_21249,N_20903,N_20717);
nand U21250 (N_21250,N_20790,N_20568);
and U21251 (N_21251,N_20982,N_20582);
and U21252 (N_21252,N_20880,N_20881);
or U21253 (N_21253,N_20593,N_20642);
or U21254 (N_21254,N_20555,N_20880);
or U21255 (N_21255,N_20920,N_20758);
and U21256 (N_21256,N_20637,N_20712);
and U21257 (N_21257,N_20765,N_20541);
nand U21258 (N_21258,N_20640,N_20810);
or U21259 (N_21259,N_20603,N_20553);
and U21260 (N_21260,N_20512,N_20649);
nor U21261 (N_21261,N_20969,N_20548);
nor U21262 (N_21262,N_20744,N_20992);
and U21263 (N_21263,N_20829,N_20807);
and U21264 (N_21264,N_20885,N_20674);
or U21265 (N_21265,N_20876,N_20649);
nand U21266 (N_21266,N_20600,N_20524);
nand U21267 (N_21267,N_20668,N_20694);
nor U21268 (N_21268,N_20810,N_20513);
nor U21269 (N_21269,N_20621,N_20951);
nand U21270 (N_21270,N_20832,N_20825);
xor U21271 (N_21271,N_20852,N_20546);
nor U21272 (N_21272,N_20959,N_20947);
xor U21273 (N_21273,N_20619,N_20636);
or U21274 (N_21274,N_20670,N_20676);
nand U21275 (N_21275,N_20556,N_20653);
and U21276 (N_21276,N_20954,N_20719);
and U21277 (N_21277,N_20872,N_20567);
nand U21278 (N_21278,N_20908,N_20716);
or U21279 (N_21279,N_20811,N_20953);
nand U21280 (N_21280,N_20885,N_20535);
xor U21281 (N_21281,N_20710,N_20744);
and U21282 (N_21282,N_20722,N_20868);
and U21283 (N_21283,N_20823,N_20869);
nor U21284 (N_21284,N_20783,N_20741);
and U21285 (N_21285,N_20617,N_20959);
nor U21286 (N_21286,N_20852,N_20907);
xor U21287 (N_21287,N_20668,N_20923);
or U21288 (N_21288,N_20986,N_20876);
and U21289 (N_21289,N_20617,N_20697);
nor U21290 (N_21290,N_20989,N_20583);
nor U21291 (N_21291,N_20668,N_20588);
nand U21292 (N_21292,N_20559,N_20729);
nand U21293 (N_21293,N_20985,N_20788);
xnor U21294 (N_21294,N_20740,N_20578);
xnor U21295 (N_21295,N_20630,N_20670);
and U21296 (N_21296,N_20629,N_20958);
and U21297 (N_21297,N_20939,N_20936);
nand U21298 (N_21298,N_20787,N_20720);
nand U21299 (N_21299,N_20785,N_20753);
and U21300 (N_21300,N_20643,N_20631);
and U21301 (N_21301,N_20844,N_20806);
nand U21302 (N_21302,N_20561,N_20885);
and U21303 (N_21303,N_20710,N_20827);
and U21304 (N_21304,N_20722,N_20802);
and U21305 (N_21305,N_20728,N_20827);
nand U21306 (N_21306,N_20983,N_20981);
nand U21307 (N_21307,N_20523,N_20504);
or U21308 (N_21308,N_20675,N_20525);
and U21309 (N_21309,N_20502,N_20554);
nor U21310 (N_21310,N_20859,N_20715);
or U21311 (N_21311,N_20738,N_20826);
nor U21312 (N_21312,N_20943,N_20907);
and U21313 (N_21313,N_20972,N_20885);
and U21314 (N_21314,N_20550,N_20574);
or U21315 (N_21315,N_20557,N_20552);
nand U21316 (N_21316,N_20921,N_20973);
nand U21317 (N_21317,N_20953,N_20847);
and U21318 (N_21318,N_20690,N_20982);
nand U21319 (N_21319,N_20904,N_20566);
and U21320 (N_21320,N_20625,N_20728);
nor U21321 (N_21321,N_20910,N_20977);
nand U21322 (N_21322,N_20668,N_20806);
xor U21323 (N_21323,N_20822,N_20857);
and U21324 (N_21324,N_20573,N_20529);
nor U21325 (N_21325,N_20624,N_20813);
nand U21326 (N_21326,N_20867,N_20832);
nand U21327 (N_21327,N_20971,N_20607);
and U21328 (N_21328,N_20840,N_20685);
nand U21329 (N_21329,N_20832,N_20914);
nand U21330 (N_21330,N_20845,N_20758);
nor U21331 (N_21331,N_20970,N_20675);
or U21332 (N_21332,N_20554,N_20988);
and U21333 (N_21333,N_20928,N_20807);
nand U21334 (N_21334,N_20677,N_20783);
and U21335 (N_21335,N_20607,N_20543);
or U21336 (N_21336,N_20504,N_20645);
nor U21337 (N_21337,N_20563,N_20780);
xnor U21338 (N_21338,N_20953,N_20786);
nand U21339 (N_21339,N_20812,N_20644);
nand U21340 (N_21340,N_20784,N_20938);
and U21341 (N_21341,N_20903,N_20972);
nor U21342 (N_21342,N_20933,N_20525);
nand U21343 (N_21343,N_20590,N_20749);
nand U21344 (N_21344,N_20581,N_20569);
nand U21345 (N_21345,N_20722,N_20959);
and U21346 (N_21346,N_20829,N_20792);
xor U21347 (N_21347,N_20666,N_20664);
or U21348 (N_21348,N_20571,N_20583);
and U21349 (N_21349,N_20613,N_20658);
or U21350 (N_21350,N_20840,N_20992);
nand U21351 (N_21351,N_20753,N_20770);
nor U21352 (N_21352,N_20501,N_20642);
nand U21353 (N_21353,N_20672,N_20707);
nor U21354 (N_21354,N_20924,N_20883);
and U21355 (N_21355,N_20819,N_20904);
xor U21356 (N_21356,N_20802,N_20879);
nor U21357 (N_21357,N_20652,N_20897);
nand U21358 (N_21358,N_20914,N_20522);
xor U21359 (N_21359,N_20805,N_20599);
nand U21360 (N_21360,N_20802,N_20936);
or U21361 (N_21361,N_20848,N_20948);
or U21362 (N_21362,N_20842,N_20993);
xor U21363 (N_21363,N_20769,N_20966);
xor U21364 (N_21364,N_20920,N_20591);
nor U21365 (N_21365,N_20998,N_20692);
nor U21366 (N_21366,N_20787,N_20600);
xnor U21367 (N_21367,N_20679,N_20944);
xnor U21368 (N_21368,N_20796,N_20995);
nor U21369 (N_21369,N_20518,N_20627);
nor U21370 (N_21370,N_20615,N_20627);
nor U21371 (N_21371,N_20725,N_20669);
nor U21372 (N_21372,N_20932,N_20930);
xor U21373 (N_21373,N_20711,N_20930);
and U21374 (N_21374,N_20585,N_20955);
or U21375 (N_21375,N_20863,N_20655);
and U21376 (N_21376,N_20566,N_20908);
xnor U21377 (N_21377,N_20840,N_20951);
nor U21378 (N_21378,N_20951,N_20871);
nand U21379 (N_21379,N_20640,N_20878);
nand U21380 (N_21380,N_20718,N_20529);
or U21381 (N_21381,N_20850,N_20799);
nor U21382 (N_21382,N_20529,N_20809);
nor U21383 (N_21383,N_20933,N_20992);
or U21384 (N_21384,N_20811,N_20747);
or U21385 (N_21385,N_20778,N_20584);
or U21386 (N_21386,N_20696,N_20861);
nor U21387 (N_21387,N_20510,N_20679);
and U21388 (N_21388,N_20959,N_20776);
nand U21389 (N_21389,N_20803,N_20866);
xor U21390 (N_21390,N_20545,N_20892);
nor U21391 (N_21391,N_20909,N_20601);
nor U21392 (N_21392,N_20860,N_20890);
or U21393 (N_21393,N_20814,N_20846);
or U21394 (N_21394,N_20710,N_20695);
xor U21395 (N_21395,N_20693,N_20667);
xnor U21396 (N_21396,N_20969,N_20938);
nor U21397 (N_21397,N_20603,N_20994);
and U21398 (N_21398,N_20690,N_20933);
or U21399 (N_21399,N_20648,N_20647);
or U21400 (N_21400,N_20940,N_20943);
nand U21401 (N_21401,N_20612,N_20644);
or U21402 (N_21402,N_20900,N_20561);
xnor U21403 (N_21403,N_20871,N_20859);
and U21404 (N_21404,N_20773,N_20736);
or U21405 (N_21405,N_20736,N_20769);
and U21406 (N_21406,N_20920,N_20522);
nor U21407 (N_21407,N_20973,N_20601);
and U21408 (N_21408,N_20916,N_20816);
and U21409 (N_21409,N_20577,N_20507);
and U21410 (N_21410,N_20747,N_20969);
nand U21411 (N_21411,N_20568,N_20562);
nand U21412 (N_21412,N_20784,N_20915);
or U21413 (N_21413,N_20710,N_20755);
or U21414 (N_21414,N_20916,N_20830);
or U21415 (N_21415,N_20568,N_20990);
or U21416 (N_21416,N_20878,N_20609);
or U21417 (N_21417,N_20504,N_20515);
nand U21418 (N_21418,N_20840,N_20758);
and U21419 (N_21419,N_20514,N_20551);
or U21420 (N_21420,N_20778,N_20599);
and U21421 (N_21421,N_20832,N_20945);
nor U21422 (N_21422,N_20799,N_20993);
nand U21423 (N_21423,N_20642,N_20768);
and U21424 (N_21424,N_20820,N_20765);
and U21425 (N_21425,N_20950,N_20747);
nand U21426 (N_21426,N_20812,N_20554);
and U21427 (N_21427,N_20695,N_20836);
xor U21428 (N_21428,N_20756,N_20786);
nor U21429 (N_21429,N_20668,N_20618);
and U21430 (N_21430,N_20761,N_20858);
and U21431 (N_21431,N_20734,N_20739);
and U21432 (N_21432,N_20752,N_20842);
nand U21433 (N_21433,N_20568,N_20658);
nand U21434 (N_21434,N_20851,N_20820);
nand U21435 (N_21435,N_20844,N_20838);
nand U21436 (N_21436,N_20911,N_20990);
or U21437 (N_21437,N_20986,N_20970);
and U21438 (N_21438,N_20881,N_20803);
nor U21439 (N_21439,N_20719,N_20521);
and U21440 (N_21440,N_20901,N_20736);
or U21441 (N_21441,N_20686,N_20548);
and U21442 (N_21442,N_20907,N_20918);
nand U21443 (N_21443,N_20732,N_20930);
nor U21444 (N_21444,N_20569,N_20685);
or U21445 (N_21445,N_20886,N_20982);
nand U21446 (N_21446,N_20545,N_20528);
and U21447 (N_21447,N_20597,N_20565);
nand U21448 (N_21448,N_20796,N_20609);
nor U21449 (N_21449,N_20921,N_20968);
nand U21450 (N_21450,N_20808,N_20592);
nand U21451 (N_21451,N_20749,N_20587);
and U21452 (N_21452,N_20688,N_20913);
and U21453 (N_21453,N_20728,N_20650);
nand U21454 (N_21454,N_20814,N_20727);
and U21455 (N_21455,N_20957,N_20967);
and U21456 (N_21456,N_20895,N_20548);
and U21457 (N_21457,N_20682,N_20803);
and U21458 (N_21458,N_20779,N_20916);
nor U21459 (N_21459,N_20695,N_20678);
nor U21460 (N_21460,N_20638,N_20564);
or U21461 (N_21461,N_20503,N_20897);
nor U21462 (N_21462,N_20722,N_20647);
nand U21463 (N_21463,N_20682,N_20503);
and U21464 (N_21464,N_20995,N_20779);
nand U21465 (N_21465,N_20740,N_20879);
and U21466 (N_21466,N_20719,N_20695);
nor U21467 (N_21467,N_20824,N_20539);
nand U21468 (N_21468,N_20800,N_20826);
nor U21469 (N_21469,N_20549,N_20746);
nor U21470 (N_21470,N_20824,N_20674);
nor U21471 (N_21471,N_20939,N_20681);
nand U21472 (N_21472,N_20604,N_20922);
or U21473 (N_21473,N_20732,N_20794);
xor U21474 (N_21474,N_20863,N_20609);
nand U21475 (N_21475,N_20858,N_20720);
or U21476 (N_21476,N_20956,N_20594);
and U21477 (N_21477,N_20974,N_20675);
or U21478 (N_21478,N_20807,N_20886);
xnor U21479 (N_21479,N_20609,N_20635);
nor U21480 (N_21480,N_20778,N_20729);
and U21481 (N_21481,N_20726,N_20989);
nand U21482 (N_21482,N_20862,N_20783);
xor U21483 (N_21483,N_20818,N_20672);
nor U21484 (N_21484,N_20550,N_20971);
or U21485 (N_21485,N_20586,N_20705);
nand U21486 (N_21486,N_20588,N_20934);
nand U21487 (N_21487,N_20585,N_20576);
nand U21488 (N_21488,N_20828,N_20969);
xor U21489 (N_21489,N_20758,N_20729);
nand U21490 (N_21490,N_20584,N_20780);
nor U21491 (N_21491,N_20765,N_20683);
nor U21492 (N_21492,N_20781,N_20519);
xor U21493 (N_21493,N_20798,N_20556);
or U21494 (N_21494,N_20615,N_20861);
or U21495 (N_21495,N_20937,N_20526);
nand U21496 (N_21496,N_20624,N_20557);
nand U21497 (N_21497,N_20970,N_20721);
or U21498 (N_21498,N_20570,N_20882);
and U21499 (N_21499,N_20913,N_20564);
nand U21500 (N_21500,N_21461,N_21212);
or U21501 (N_21501,N_21350,N_21166);
and U21502 (N_21502,N_21072,N_21439);
and U21503 (N_21503,N_21286,N_21027);
nand U21504 (N_21504,N_21100,N_21404);
nand U21505 (N_21505,N_21043,N_21265);
and U21506 (N_21506,N_21255,N_21460);
nand U21507 (N_21507,N_21332,N_21170);
nand U21508 (N_21508,N_21312,N_21297);
and U21509 (N_21509,N_21381,N_21154);
nor U21510 (N_21510,N_21472,N_21339);
and U21511 (N_21511,N_21457,N_21361);
and U21512 (N_21512,N_21483,N_21022);
nor U21513 (N_21513,N_21360,N_21225);
nand U21514 (N_21514,N_21038,N_21264);
nand U21515 (N_21515,N_21261,N_21064);
nor U21516 (N_21516,N_21096,N_21206);
xor U21517 (N_21517,N_21270,N_21198);
or U21518 (N_21518,N_21191,N_21383);
nand U21519 (N_21519,N_21498,N_21428);
nor U21520 (N_21520,N_21387,N_21474);
nand U21521 (N_21521,N_21056,N_21172);
or U21522 (N_21522,N_21378,N_21343);
nor U21523 (N_21523,N_21321,N_21389);
nand U21524 (N_21524,N_21213,N_21464);
xor U21525 (N_21525,N_21130,N_21340);
nand U21526 (N_21526,N_21160,N_21099);
or U21527 (N_21527,N_21303,N_21116);
nor U21528 (N_21528,N_21491,N_21415);
xnor U21529 (N_21529,N_21436,N_21456);
nor U21530 (N_21530,N_21115,N_21071);
nand U21531 (N_21531,N_21142,N_21251);
xnor U21532 (N_21532,N_21434,N_21399);
and U21533 (N_21533,N_21336,N_21246);
and U21534 (N_21534,N_21466,N_21290);
nor U21535 (N_21535,N_21074,N_21050);
nand U21536 (N_21536,N_21144,N_21053);
or U21537 (N_21537,N_21220,N_21242);
nand U21538 (N_21538,N_21318,N_21165);
nor U21539 (N_21539,N_21094,N_21259);
nand U21540 (N_21540,N_21224,N_21054);
nand U21541 (N_21541,N_21473,N_21407);
nand U21542 (N_21542,N_21450,N_21398);
and U21543 (N_21543,N_21396,N_21364);
or U21544 (N_21544,N_21269,N_21486);
xnor U21545 (N_21545,N_21310,N_21244);
and U21546 (N_21546,N_21218,N_21216);
xor U21547 (N_21547,N_21232,N_21017);
or U21548 (N_21548,N_21449,N_21186);
xnor U21549 (N_21549,N_21068,N_21189);
or U21550 (N_21550,N_21032,N_21114);
or U21551 (N_21551,N_21372,N_21499);
nor U21552 (N_21552,N_21233,N_21300);
nand U21553 (N_21553,N_21275,N_21370);
or U21554 (N_21554,N_21497,N_21322);
nor U21555 (N_21555,N_21397,N_21047);
xor U21556 (N_21556,N_21055,N_21247);
and U21557 (N_21557,N_21049,N_21257);
and U21558 (N_21558,N_21230,N_21204);
and U21559 (N_21559,N_21291,N_21459);
or U21560 (N_21560,N_21023,N_21152);
xor U21561 (N_21561,N_21347,N_21119);
and U21562 (N_21562,N_21059,N_21402);
or U21563 (N_21563,N_21042,N_21129);
and U21564 (N_21564,N_21195,N_21308);
xnor U21565 (N_21565,N_21177,N_21124);
or U21566 (N_21566,N_21319,N_21330);
nand U21567 (N_21567,N_21006,N_21423);
and U21568 (N_21568,N_21101,N_21469);
xnor U21569 (N_21569,N_21210,N_21240);
nor U21570 (N_21570,N_21093,N_21202);
or U21571 (N_21571,N_21097,N_21418);
nand U21572 (N_21572,N_21077,N_21446);
or U21573 (N_21573,N_21406,N_21482);
and U21574 (N_21574,N_21086,N_21488);
and U21575 (N_21575,N_21438,N_21139);
nor U21576 (N_21576,N_21203,N_21293);
nand U21577 (N_21577,N_21263,N_21117);
xor U21578 (N_21578,N_21085,N_21288);
xor U21579 (N_21579,N_21136,N_21409);
xor U21580 (N_21580,N_21181,N_21458);
nor U21581 (N_21581,N_21487,N_21348);
and U21582 (N_21582,N_21252,N_21476);
nand U21583 (N_21583,N_21173,N_21120);
nor U21584 (N_21584,N_21306,N_21284);
and U21585 (N_21585,N_21316,N_21337);
and U21586 (N_21586,N_21442,N_21024);
nand U21587 (N_21587,N_21333,N_21478);
nand U21588 (N_21588,N_21193,N_21048);
nand U21589 (N_21589,N_21278,N_21279);
nand U21590 (N_21590,N_21073,N_21123);
or U21591 (N_21591,N_21470,N_21179);
nand U21592 (N_21592,N_21107,N_21421);
nor U21593 (N_21593,N_21214,N_21400);
nor U21594 (N_21594,N_21234,N_21149);
or U21595 (N_21595,N_21271,N_21151);
xnor U21596 (N_21596,N_21126,N_21182);
or U21597 (N_21597,N_21125,N_21067);
nor U21598 (N_21598,N_21163,N_21062);
or U21599 (N_21599,N_21001,N_21040);
nand U21600 (N_21600,N_21237,N_21345);
or U21601 (N_21601,N_21135,N_21245);
nor U21602 (N_21602,N_21417,N_21395);
xnor U21603 (N_21603,N_21238,N_21133);
nor U21604 (N_21604,N_21044,N_21015);
or U21605 (N_21605,N_21307,N_21108);
or U21606 (N_21606,N_21034,N_21157);
and U21607 (N_21607,N_21137,N_21128);
nand U21608 (N_21608,N_21441,N_21065);
nand U21609 (N_21609,N_21187,N_21223);
nor U21610 (N_21610,N_21258,N_21298);
xnor U21611 (N_21611,N_21102,N_21036);
xor U21612 (N_21612,N_21164,N_21443);
nor U21613 (N_21613,N_21296,N_21021);
or U21614 (N_21614,N_21090,N_21080);
nand U21615 (N_21615,N_21197,N_21287);
nor U21616 (N_21616,N_21363,N_21026);
or U21617 (N_21617,N_21035,N_21283);
and U21618 (N_21618,N_21150,N_21490);
nor U21619 (N_21619,N_21411,N_21304);
nand U21620 (N_21620,N_21424,N_21243);
nand U21621 (N_21621,N_21200,N_21393);
nand U21622 (N_21622,N_21380,N_21430);
nor U21623 (N_21623,N_21352,N_21317);
nand U21624 (N_21624,N_21280,N_21127);
or U21625 (N_21625,N_21480,N_21199);
and U21626 (N_21626,N_21256,N_21250);
nand U21627 (N_21627,N_21103,N_21176);
nor U21628 (N_21628,N_21328,N_21394);
nor U21629 (N_21629,N_21121,N_21037);
or U21630 (N_21630,N_21433,N_21010);
nor U21631 (N_21631,N_21358,N_21109);
or U21632 (N_21632,N_21029,N_21002);
or U21633 (N_21633,N_21069,N_21083);
nor U21634 (N_21634,N_21344,N_21305);
nand U21635 (N_21635,N_21063,N_21081);
or U21636 (N_21636,N_21066,N_21341);
or U21637 (N_21637,N_21188,N_21386);
xor U21638 (N_21638,N_21159,N_21311);
xnor U21639 (N_21639,N_21095,N_21485);
xnor U21640 (N_21640,N_21475,N_21414);
nand U21641 (N_21641,N_21184,N_21468);
and U21642 (N_21642,N_21429,N_21426);
or U21643 (N_21643,N_21405,N_21260);
nand U21644 (N_21644,N_21357,N_21391);
and U21645 (N_21645,N_21329,N_21392);
nand U21646 (N_21646,N_21057,N_21228);
or U21647 (N_21647,N_21175,N_21005);
or U21648 (N_21648,N_21025,N_21289);
or U21649 (N_21649,N_21041,N_21326);
and U21650 (N_21650,N_21302,N_21362);
and U21651 (N_21651,N_21366,N_21236);
or U21652 (N_21652,N_21106,N_21020);
xnor U21653 (N_21653,N_21104,N_21373);
nor U21654 (N_21654,N_21138,N_21075);
xnor U21655 (N_21655,N_21309,N_21384);
nor U21656 (N_21656,N_21355,N_21431);
or U21657 (N_21657,N_21465,N_21285);
and U21658 (N_21658,N_21131,N_21167);
or U21659 (N_21659,N_21408,N_21008);
nand U21660 (N_21660,N_21454,N_21248);
or U21661 (N_21661,N_21004,N_21254);
nor U21662 (N_21662,N_21241,N_21379);
or U21663 (N_21663,N_21011,N_21003);
and U21664 (N_21664,N_21327,N_21219);
nand U21665 (N_21665,N_21158,N_21039);
xnor U21666 (N_21666,N_21292,N_21227);
nor U21667 (N_21667,N_21060,N_21194);
or U21668 (N_21668,N_21078,N_21013);
or U21669 (N_21669,N_21374,N_21016);
nor U21670 (N_21670,N_21413,N_21208);
or U21671 (N_21671,N_21432,N_21143);
or U21672 (N_21672,N_21422,N_21325);
or U21673 (N_21673,N_21425,N_21281);
nand U21674 (N_21674,N_21051,N_21496);
nor U21675 (N_21675,N_21058,N_21267);
nor U21676 (N_21676,N_21092,N_21435);
nor U21677 (N_21677,N_21141,N_21444);
nand U21678 (N_21678,N_21419,N_21087);
and U21679 (N_21679,N_21201,N_21205);
nor U21680 (N_21680,N_21410,N_21229);
nor U21681 (N_21681,N_21018,N_21376);
nor U21682 (N_21682,N_21192,N_21162);
or U21683 (N_21683,N_21353,N_21132);
xor U21684 (N_21684,N_21365,N_21088);
nand U21685 (N_21685,N_21009,N_21276);
nor U21686 (N_21686,N_21076,N_21105);
and U21687 (N_21687,N_21156,N_21161);
nor U21688 (N_21688,N_21437,N_21155);
or U21689 (N_21689,N_21226,N_21489);
nor U21690 (N_21690,N_21494,N_21014);
or U21691 (N_21691,N_21148,N_21215);
or U21692 (N_21692,N_21171,N_21122);
nor U21693 (N_21693,N_21084,N_21153);
and U21694 (N_21694,N_21046,N_21000);
nor U21695 (N_21695,N_21268,N_21481);
nand U21696 (N_21696,N_21338,N_21112);
or U21697 (N_21697,N_21221,N_21334);
and U21698 (N_21698,N_21349,N_21007);
or U21699 (N_21699,N_21385,N_21356);
or U21700 (N_21700,N_21113,N_21174);
nand U21701 (N_21701,N_21440,N_21335);
nand U21702 (N_21702,N_21253,N_21467);
nand U21703 (N_21703,N_21180,N_21448);
nand U21704 (N_21704,N_21030,N_21178);
or U21705 (N_21705,N_21479,N_21146);
xnor U21706 (N_21706,N_21211,N_21462);
and U21707 (N_21707,N_21196,N_21168);
nand U21708 (N_21708,N_21098,N_21299);
or U21709 (N_21709,N_21455,N_21209);
xor U21710 (N_21710,N_21061,N_21477);
nand U21711 (N_21711,N_21453,N_21012);
nor U21712 (N_21712,N_21323,N_21342);
or U21713 (N_21713,N_21346,N_21492);
xnor U21714 (N_21714,N_21375,N_21183);
xnor U21715 (N_21715,N_21207,N_21367);
nand U21716 (N_21716,N_21484,N_21382);
nor U21717 (N_21717,N_21273,N_21315);
and U21718 (N_21718,N_21351,N_21313);
or U21719 (N_21719,N_21028,N_21412);
nand U21720 (N_21720,N_21089,N_21277);
or U21721 (N_21721,N_21294,N_21359);
or U21722 (N_21722,N_21145,N_21320);
and U21723 (N_21723,N_21371,N_21274);
or U21724 (N_21724,N_21217,N_21354);
or U21725 (N_21725,N_21070,N_21445);
and U21726 (N_21726,N_21282,N_21471);
xor U21727 (N_21727,N_21388,N_21420);
nor U21728 (N_21728,N_21495,N_21324);
nor U21729 (N_21729,N_21401,N_21295);
nand U21730 (N_21730,N_21091,N_21239);
nor U21731 (N_21731,N_21262,N_21266);
xnor U21732 (N_21732,N_21222,N_21118);
xnor U21733 (N_21733,N_21140,N_21447);
and U21734 (N_21734,N_21301,N_21377);
nor U21735 (N_21735,N_21390,N_21045);
xor U21736 (N_21736,N_21079,N_21416);
nor U21737 (N_21737,N_21033,N_21452);
nor U21738 (N_21738,N_21272,N_21185);
or U21739 (N_21739,N_21368,N_21147);
and U21740 (N_21740,N_21314,N_21235);
nor U21741 (N_21741,N_21249,N_21052);
or U21742 (N_21742,N_21331,N_21019);
and U21743 (N_21743,N_21031,N_21403);
and U21744 (N_21744,N_21231,N_21463);
nor U21745 (N_21745,N_21493,N_21110);
and U21746 (N_21746,N_21190,N_21111);
nand U21747 (N_21747,N_21169,N_21451);
nor U21748 (N_21748,N_21369,N_21082);
and U21749 (N_21749,N_21134,N_21427);
nor U21750 (N_21750,N_21024,N_21077);
or U21751 (N_21751,N_21178,N_21124);
or U21752 (N_21752,N_21154,N_21275);
nand U21753 (N_21753,N_21000,N_21450);
nor U21754 (N_21754,N_21140,N_21469);
and U21755 (N_21755,N_21025,N_21180);
and U21756 (N_21756,N_21320,N_21066);
and U21757 (N_21757,N_21094,N_21391);
nand U21758 (N_21758,N_21048,N_21480);
nor U21759 (N_21759,N_21025,N_21000);
xor U21760 (N_21760,N_21397,N_21275);
nand U21761 (N_21761,N_21311,N_21035);
or U21762 (N_21762,N_21149,N_21279);
nand U21763 (N_21763,N_21434,N_21462);
and U21764 (N_21764,N_21012,N_21139);
and U21765 (N_21765,N_21015,N_21251);
or U21766 (N_21766,N_21041,N_21111);
nor U21767 (N_21767,N_21294,N_21163);
xor U21768 (N_21768,N_21365,N_21185);
or U21769 (N_21769,N_21302,N_21495);
and U21770 (N_21770,N_21200,N_21389);
nand U21771 (N_21771,N_21355,N_21017);
nand U21772 (N_21772,N_21367,N_21350);
nand U21773 (N_21773,N_21204,N_21339);
and U21774 (N_21774,N_21349,N_21223);
or U21775 (N_21775,N_21072,N_21065);
nand U21776 (N_21776,N_21110,N_21021);
nor U21777 (N_21777,N_21408,N_21290);
nand U21778 (N_21778,N_21473,N_21034);
and U21779 (N_21779,N_21453,N_21339);
nor U21780 (N_21780,N_21239,N_21458);
nor U21781 (N_21781,N_21316,N_21046);
nor U21782 (N_21782,N_21436,N_21308);
and U21783 (N_21783,N_21165,N_21490);
xnor U21784 (N_21784,N_21383,N_21400);
and U21785 (N_21785,N_21197,N_21202);
nand U21786 (N_21786,N_21376,N_21404);
and U21787 (N_21787,N_21212,N_21297);
or U21788 (N_21788,N_21243,N_21331);
and U21789 (N_21789,N_21453,N_21225);
nor U21790 (N_21790,N_21063,N_21403);
nand U21791 (N_21791,N_21125,N_21425);
xnor U21792 (N_21792,N_21469,N_21408);
and U21793 (N_21793,N_21243,N_21184);
nand U21794 (N_21794,N_21352,N_21216);
and U21795 (N_21795,N_21230,N_21449);
or U21796 (N_21796,N_21201,N_21322);
nor U21797 (N_21797,N_21019,N_21138);
xor U21798 (N_21798,N_21255,N_21093);
nor U21799 (N_21799,N_21251,N_21229);
or U21800 (N_21800,N_21380,N_21166);
or U21801 (N_21801,N_21161,N_21463);
xnor U21802 (N_21802,N_21234,N_21382);
or U21803 (N_21803,N_21352,N_21063);
and U21804 (N_21804,N_21245,N_21297);
nand U21805 (N_21805,N_21218,N_21278);
or U21806 (N_21806,N_21279,N_21421);
and U21807 (N_21807,N_21375,N_21069);
and U21808 (N_21808,N_21375,N_21271);
nor U21809 (N_21809,N_21370,N_21324);
and U21810 (N_21810,N_21063,N_21135);
or U21811 (N_21811,N_21485,N_21156);
nand U21812 (N_21812,N_21397,N_21118);
xnor U21813 (N_21813,N_21374,N_21132);
xnor U21814 (N_21814,N_21282,N_21017);
xnor U21815 (N_21815,N_21447,N_21204);
nor U21816 (N_21816,N_21489,N_21029);
or U21817 (N_21817,N_21195,N_21405);
nand U21818 (N_21818,N_21051,N_21014);
or U21819 (N_21819,N_21267,N_21171);
nand U21820 (N_21820,N_21369,N_21298);
nor U21821 (N_21821,N_21092,N_21407);
nor U21822 (N_21822,N_21152,N_21121);
or U21823 (N_21823,N_21004,N_21237);
and U21824 (N_21824,N_21166,N_21177);
or U21825 (N_21825,N_21093,N_21009);
and U21826 (N_21826,N_21219,N_21168);
or U21827 (N_21827,N_21050,N_21297);
and U21828 (N_21828,N_21102,N_21373);
or U21829 (N_21829,N_21073,N_21012);
and U21830 (N_21830,N_21489,N_21493);
nor U21831 (N_21831,N_21198,N_21187);
or U21832 (N_21832,N_21090,N_21233);
or U21833 (N_21833,N_21296,N_21398);
nor U21834 (N_21834,N_21146,N_21285);
nor U21835 (N_21835,N_21411,N_21212);
nand U21836 (N_21836,N_21385,N_21047);
nand U21837 (N_21837,N_21033,N_21416);
nand U21838 (N_21838,N_21334,N_21322);
nor U21839 (N_21839,N_21361,N_21302);
and U21840 (N_21840,N_21132,N_21042);
or U21841 (N_21841,N_21140,N_21049);
nand U21842 (N_21842,N_21082,N_21486);
and U21843 (N_21843,N_21194,N_21108);
xnor U21844 (N_21844,N_21189,N_21377);
or U21845 (N_21845,N_21399,N_21051);
and U21846 (N_21846,N_21484,N_21112);
nor U21847 (N_21847,N_21229,N_21136);
or U21848 (N_21848,N_21046,N_21348);
nor U21849 (N_21849,N_21170,N_21050);
or U21850 (N_21850,N_21071,N_21358);
xor U21851 (N_21851,N_21498,N_21231);
and U21852 (N_21852,N_21331,N_21288);
and U21853 (N_21853,N_21445,N_21346);
nand U21854 (N_21854,N_21386,N_21395);
or U21855 (N_21855,N_21027,N_21006);
or U21856 (N_21856,N_21390,N_21441);
xnor U21857 (N_21857,N_21088,N_21394);
nand U21858 (N_21858,N_21104,N_21099);
nor U21859 (N_21859,N_21075,N_21311);
nor U21860 (N_21860,N_21128,N_21179);
nand U21861 (N_21861,N_21214,N_21288);
nand U21862 (N_21862,N_21274,N_21403);
or U21863 (N_21863,N_21486,N_21175);
nand U21864 (N_21864,N_21441,N_21415);
and U21865 (N_21865,N_21442,N_21128);
nand U21866 (N_21866,N_21349,N_21299);
xnor U21867 (N_21867,N_21070,N_21411);
nor U21868 (N_21868,N_21408,N_21496);
nand U21869 (N_21869,N_21424,N_21138);
xor U21870 (N_21870,N_21367,N_21345);
nor U21871 (N_21871,N_21032,N_21350);
or U21872 (N_21872,N_21312,N_21076);
or U21873 (N_21873,N_21244,N_21066);
and U21874 (N_21874,N_21057,N_21287);
nor U21875 (N_21875,N_21297,N_21132);
nand U21876 (N_21876,N_21473,N_21071);
or U21877 (N_21877,N_21036,N_21447);
nor U21878 (N_21878,N_21256,N_21405);
nand U21879 (N_21879,N_21247,N_21260);
nor U21880 (N_21880,N_21157,N_21452);
and U21881 (N_21881,N_21276,N_21412);
nand U21882 (N_21882,N_21036,N_21122);
nor U21883 (N_21883,N_21376,N_21356);
and U21884 (N_21884,N_21469,N_21125);
nor U21885 (N_21885,N_21418,N_21186);
xor U21886 (N_21886,N_21467,N_21466);
nor U21887 (N_21887,N_21413,N_21376);
or U21888 (N_21888,N_21097,N_21096);
nor U21889 (N_21889,N_21458,N_21483);
xnor U21890 (N_21890,N_21019,N_21152);
nand U21891 (N_21891,N_21430,N_21273);
nor U21892 (N_21892,N_21403,N_21072);
nand U21893 (N_21893,N_21403,N_21171);
nand U21894 (N_21894,N_21127,N_21089);
nand U21895 (N_21895,N_21095,N_21170);
nor U21896 (N_21896,N_21206,N_21419);
nor U21897 (N_21897,N_21342,N_21416);
and U21898 (N_21898,N_21027,N_21119);
and U21899 (N_21899,N_21389,N_21005);
or U21900 (N_21900,N_21437,N_21211);
nor U21901 (N_21901,N_21436,N_21077);
and U21902 (N_21902,N_21190,N_21210);
nand U21903 (N_21903,N_21049,N_21167);
nor U21904 (N_21904,N_21160,N_21045);
and U21905 (N_21905,N_21489,N_21329);
nand U21906 (N_21906,N_21271,N_21461);
and U21907 (N_21907,N_21223,N_21486);
and U21908 (N_21908,N_21168,N_21403);
nand U21909 (N_21909,N_21232,N_21244);
nor U21910 (N_21910,N_21490,N_21464);
nand U21911 (N_21911,N_21031,N_21373);
nor U21912 (N_21912,N_21470,N_21417);
nand U21913 (N_21913,N_21400,N_21345);
nor U21914 (N_21914,N_21458,N_21111);
nand U21915 (N_21915,N_21359,N_21112);
nor U21916 (N_21916,N_21365,N_21430);
or U21917 (N_21917,N_21480,N_21176);
nand U21918 (N_21918,N_21356,N_21099);
xnor U21919 (N_21919,N_21086,N_21351);
nor U21920 (N_21920,N_21130,N_21073);
nand U21921 (N_21921,N_21343,N_21218);
nor U21922 (N_21922,N_21280,N_21154);
and U21923 (N_21923,N_21490,N_21383);
or U21924 (N_21924,N_21451,N_21001);
nand U21925 (N_21925,N_21177,N_21467);
and U21926 (N_21926,N_21332,N_21158);
nor U21927 (N_21927,N_21417,N_21231);
or U21928 (N_21928,N_21343,N_21088);
or U21929 (N_21929,N_21150,N_21488);
nor U21930 (N_21930,N_21082,N_21446);
nor U21931 (N_21931,N_21029,N_21423);
and U21932 (N_21932,N_21482,N_21136);
or U21933 (N_21933,N_21342,N_21413);
or U21934 (N_21934,N_21012,N_21154);
and U21935 (N_21935,N_21371,N_21181);
or U21936 (N_21936,N_21066,N_21467);
and U21937 (N_21937,N_21070,N_21058);
nor U21938 (N_21938,N_21274,N_21243);
nor U21939 (N_21939,N_21010,N_21450);
and U21940 (N_21940,N_21111,N_21338);
or U21941 (N_21941,N_21255,N_21479);
or U21942 (N_21942,N_21301,N_21072);
or U21943 (N_21943,N_21150,N_21182);
and U21944 (N_21944,N_21421,N_21267);
or U21945 (N_21945,N_21203,N_21097);
nand U21946 (N_21946,N_21452,N_21297);
or U21947 (N_21947,N_21330,N_21270);
xnor U21948 (N_21948,N_21479,N_21477);
nand U21949 (N_21949,N_21379,N_21095);
or U21950 (N_21950,N_21264,N_21006);
and U21951 (N_21951,N_21300,N_21136);
nor U21952 (N_21952,N_21401,N_21425);
nand U21953 (N_21953,N_21112,N_21365);
and U21954 (N_21954,N_21384,N_21282);
and U21955 (N_21955,N_21050,N_21006);
or U21956 (N_21956,N_21021,N_21133);
or U21957 (N_21957,N_21238,N_21230);
nand U21958 (N_21958,N_21251,N_21097);
xnor U21959 (N_21959,N_21134,N_21306);
nor U21960 (N_21960,N_21096,N_21094);
nand U21961 (N_21961,N_21228,N_21411);
and U21962 (N_21962,N_21336,N_21463);
and U21963 (N_21963,N_21272,N_21173);
xor U21964 (N_21964,N_21175,N_21273);
or U21965 (N_21965,N_21342,N_21489);
xor U21966 (N_21966,N_21418,N_21272);
or U21967 (N_21967,N_21140,N_21058);
nor U21968 (N_21968,N_21489,N_21144);
nand U21969 (N_21969,N_21205,N_21010);
nor U21970 (N_21970,N_21473,N_21162);
and U21971 (N_21971,N_21480,N_21182);
nor U21972 (N_21972,N_21044,N_21034);
and U21973 (N_21973,N_21088,N_21041);
nor U21974 (N_21974,N_21089,N_21364);
or U21975 (N_21975,N_21292,N_21162);
nor U21976 (N_21976,N_21127,N_21296);
nand U21977 (N_21977,N_21234,N_21369);
or U21978 (N_21978,N_21287,N_21393);
or U21979 (N_21979,N_21419,N_21288);
nand U21980 (N_21980,N_21200,N_21187);
and U21981 (N_21981,N_21397,N_21484);
nor U21982 (N_21982,N_21070,N_21436);
nand U21983 (N_21983,N_21367,N_21154);
nand U21984 (N_21984,N_21460,N_21380);
and U21985 (N_21985,N_21367,N_21432);
or U21986 (N_21986,N_21484,N_21415);
or U21987 (N_21987,N_21126,N_21249);
and U21988 (N_21988,N_21322,N_21338);
xor U21989 (N_21989,N_21220,N_21106);
nor U21990 (N_21990,N_21185,N_21088);
xor U21991 (N_21991,N_21376,N_21458);
nor U21992 (N_21992,N_21049,N_21002);
nand U21993 (N_21993,N_21006,N_21338);
nand U21994 (N_21994,N_21268,N_21062);
nand U21995 (N_21995,N_21130,N_21203);
nand U21996 (N_21996,N_21343,N_21174);
nor U21997 (N_21997,N_21071,N_21462);
nand U21998 (N_21998,N_21349,N_21202);
nand U21999 (N_21999,N_21404,N_21146);
and U22000 (N_22000,N_21732,N_21971);
nor U22001 (N_22001,N_21575,N_21852);
nor U22002 (N_22002,N_21976,N_21592);
nor U22003 (N_22003,N_21869,N_21996);
and U22004 (N_22004,N_21540,N_21777);
or U22005 (N_22005,N_21662,N_21628);
and U22006 (N_22006,N_21951,N_21938);
nand U22007 (N_22007,N_21847,N_21934);
or U22008 (N_22008,N_21990,N_21846);
nor U22009 (N_22009,N_21663,N_21578);
and U22010 (N_22010,N_21747,N_21969);
or U22011 (N_22011,N_21792,N_21964);
nand U22012 (N_22012,N_21854,N_21978);
and U22013 (N_22013,N_21911,N_21941);
nor U22014 (N_22014,N_21970,N_21625);
nor U22015 (N_22015,N_21639,N_21679);
nor U22016 (N_22016,N_21793,N_21764);
nand U22017 (N_22017,N_21811,N_21900);
nand U22018 (N_22018,N_21587,N_21708);
and U22019 (N_22019,N_21640,N_21877);
and U22020 (N_22020,N_21907,N_21956);
xnor U22021 (N_22021,N_21682,N_21830);
nor U22022 (N_22022,N_21913,N_21521);
and U22023 (N_22023,N_21901,N_21994);
and U22024 (N_22024,N_21714,N_21678);
nor U22025 (N_22025,N_21925,N_21706);
nand U22026 (N_22026,N_21801,N_21888);
or U22027 (N_22027,N_21776,N_21594);
xnor U22028 (N_22028,N_21790,N_21928);
nor U22029 (N_22029,N_21999,N_21556);
and U22030 (N_22030,N_21748,N_21885);
nand U22031 (N_22031,N_21853,N_21942);
or U22032 (N_22032,N_21570,N_21865);
or U22033 (N_22033,N_21689,N_21519);
or U22034 (N_22034,N_21543,N_21589);
nor U22035 (N_22035,N_21965,N_21805);
and U22036 (N_22036,N_21711,N_21960);
nand U22037 (N_22037,N_21810,N_21909);
nand U22038 (N_22038,N_21532,N_21768);
or U22039 (N_22039,N_21564,N_21986);
and U22040 (N_22040,N_21981,N_21939);
and U22041 (N_22041,N_21650,N_21765);
and U22042 (N_22042,N_21541,N_21850);
or U22043 (N_22043,N_21936,N_21522);
nand U22044 (N_22044,N_21574,N_21526);
nand U22045 (N_22045,N_21896,N_21596);
or U22046 (N_22046,N_21696,N_21755);
nand U22047 (N_22047,N_21812,N_21518);
nand U22048 (N_22048,N_21831,N_21547);
nand U22049 (N_22049,N_21557,N_21736);
and U22050 (N_22050,N_21549,N_21873);
nor U22051 (N_22051,N_21593,N_21733);
nor U22052 (N_22052,N_21641,N_21802);
and U22053 (N_22053,N_21757,N_21788);
nand U22054 (N_22054,N_21739,N_21848);
and U22055 (N_22055,N_21945,N_21535);
nor U22056 (N_22056,N_21503,N_21646);
nand U22057 (N_22057,N_21836,N_21983);
xnor U22058 (N_22058,N_21814,N_21858);
and U22059 (N_22059,N_21891,N_21502);
nor U22060 (N_22060,N_21955,N_21579);
nand U22061 (N_22061,N_21527,N_21681);
xnor U22062 (N_22062,N_21767,N_21712);
xor U22063 (N_22063,N_21989,N_21709);
or U22064 (N_22064,N_21600,N_21881);
or U22065 (N_22065,N_21742,N_21729);
or U22066 (N_22066,N_21829,N_21619);
or U22067 (N_22067,N_21963,N_21828);
xnor U22068 (N_22068,N_21694,N_21899);
or U22069 (N_22069,N_21751,N_21898);
nand U22070 (N_22070,N_21642,N_21720);
xor U22071 (N_22071,N_21966,N_21670);
nand U22072 (N_22072,N_21937,N_21538);
nor U22073 (N_22073,N_21508,N_21560);
and U22074 (N_22074,N_21948,N_21552);
or U22075 (N_22075,N_21837,N_21800);
or U22076 (N_22076,N_21878,N_21982);
and U22077 (N_22077,N_21779,N_21988);
and U22078 (N_22078,N_21601,N_21887);
or U22079 (N_22079,N_21664,N_21883);
xor U22080 (N_22080,N_21554,N_21632);
and U22081 (N_22081,N_21544,N_21821);
nor U22082 (N_22082,N_21571,N_21880);
xnor U22083 (N_22083,N_21809,N_21621);
nor U22084 (N_22084,N_21871,N_21895);
and U22085 (N_22085,N_21787,N_21804);
nor U22086 (N_22086,N_21954,N_21902);
nor U22087 (N_22087,N_21661,N_21676);
nor U22088 (N_22088,N_21692,N_21998);
nand U22089 (N_22089,N_21660,N_21760);
nor U22090 (N_22090,N_21824,N_21548);
or U22091 (N_22091,N_21944,N_21533);
and U22092 (N_22092,N_21607,N_21725);
nor U22093 (N_22093,N_21980,N_21700);
or U22094 (N_22094,N_21935,N_21961);
nand U22095 (N_22095,N_21746,N_21699);
nor U22096 (N_22096,N_21629,N_21603);
or U22097 (N_22097,N_21512,N_21856);
nand U22098 (N_22098,N_21940,N_21826);
nand U22099 (N_22099,N_21506,N_21823);
nand U22100 (N_22100,N_21542,N_21763);
nand U22101 (N_22101,N_21918,N_21919);
nor U22102 (N_22102,N_21819,N_21717);
nor U22103 (N_22103,N_21580,N_21611);
nand U22104 (N_22104,N_21946,N_21649);
nand U22105 (N_22105,N_21666,N_21766);
nor U22106 (N_22106,N_21816,N_21833);
and U22107 (N_22107,N_21703,N_21894);
or U22108 (N_22108,N_21573,N_21710);
or U22109 (N_22109,N_21673,N_21675);
or U22110 (N_22110,N_21950,N_21973);
and U22111 (N_22111,N_21588,N_21513);
nand U22112 (N_22112,N_21604,N_21558);
and U22113 (N_22113,N_21866,N_21618);
nor U22114 (N_22114,N_21778,N_21569);
nand U22115 (N_22115,N_21912,N_21683);
nand U22116 (N_22116,N_21627,N_21555);
or U22117 (N_22117,N_21862,N_21991);
and U22118 (N_22118,N_21718,N_21827);
xor U22119 (N_22119,N_21817,N_21545);
nand U22120 (N_22120,N_21652,N_21813);
and U22121 (N_22121,N_21845,N_21882);
nor U22122 (N_22122,N_21536,N_21968);
and U22123 (N_22123,N_21834,N_21616);
nand U22124 (N_22124,N_21537,N_21566);
or U22125 (N_22125,N_21731,N_21576);
nor U22126 (N_22126,N_21644,N_21719);
xor U22127 (N_22127,N_21977,N_21889);
and U22128 (N_22128,N_21745,N_21643);
or U22129 (N_22129,N_21550,N_21638);
xnor U22130 (N_22130,N_21608,N_21721);
or U22131 (N_22131,N_21959,N_21626);
nor U22132 (N_22132,N_21953,N_21553);
or U22133 (N_22133,N_21780,N_21943);
nand U22134 (N_22134,N_21920,N_21685);
and U22135 (N_22135,N_21926,N_21623);
nand U22136 (N_22136,N_21794,N_21688);
and U22137 (N_22137,N_21995,N_21658);
or U22138 (N_22138,N_21726,N_21539);
or U22139 (N_22139,N_21617,N_21500);
nand U22140 (N_22140,N_21752,N_21781);
and U22141 (N_22141,N_21645,N_21750);
xor U22142 (N_22142,N_21908,N_21864);
nor U22143 (N_22143,N_21905,N_21657);
and U22144 (N_22144,N_21947,N_21668);
or U22145 (N_22145,N_21724,N_21597);
or U22146 (N_22146,N_21528,N_21654);
and U22147 (N_22147,N_21789,N_21609);
or U22148 (N_22148,N_21842,N_21586);
nor U22149 (N_22149,N_21872,N_21761);
nor U22150 (N_22150,N_21504,N_21775);
nor U22151 (N_22151,N_21505,N_21738);
nand U22152 (N_22152,N_21653,N_21797);
and U22153 (N_22153,N_21677,N_21933);
xor U22154 (N_22154,N_21599,N_21843);
and U22155 (N_22155,N_21930,N_21822);
or U22156 (N_22156,N_21655,N_21507);
or U22157 (N_22157,N_21859,N_21516);
or U22158 (N_22158,N_21501,N_21784);
nand U22159 (N_22159,N_21511,N_21631);
or U22160 (N_22160,N_21952,N_21637);
nand U22161 (N_22161,N_21665,N_21927);
and U22162 (N_22162,N_21903,N_21734);
or U22163 (N_22163,N_21693,N_21838);
or U22164 (N_22164,N_21904,N_21774);
nor U22165 (N_22165,N_21922,N_21605);
nor U22166 (N_22166,N_21635,N_21713);
nand U22167 (N_22167,N_21754,N_21698);
xor U22168 (N_22168,N_21892,N_21667);
nand U22169 (N_22169,N_21572,N_21531);
and U22170 (N_22170,N_21598,N_21975);
xor U22171 (N_22171,N_21932,N_21705);
or U22172 (N_22172,N_21874,N_21671);
nand U22173 (N_22173,N_21987,N_21562);
xnor U22174 (N_22174,N_21860,N_21762);
nand U22175 (N_22175,N_21857,N_21759);
nand U22176 (N_22176,N_21770,N_21551);
xor U22177 (N_22177,N_21915,N_21840);
and U22178 (N_22178,N_21647,N_21741);
and U22179 (N_22179,N_21796,N_21844);
and U22180 (N_22180,N_21879,N_21884);
and U22181 (N_22181,N_21924,N_21876);
nor U22182 (N_22182,N_21515,N_21722);
nor U22183 (N_22183,N_21674,N_21523);
and U22184 (N_22184,N_21798,N_21806);
xor U22185 (N_22185,N_21851,N_21559);
and U22186 (N_22186,N_21634,N_21690);
or U22187 (N_22187,N_21656,N_21743);
nand U22188 (N_22188,N_21730,N_21735);
or U22189 (N_22189,N_21680,N_21737);
xor U22190 (N_22190,N_21565,N_21782);
nand U22191 (N_22191,N_21695,N_21524);
nand U22192 (N_22192,N_21613,N_21795);
nor U22193 (N_22193,N_21855,N_21577);
or U22194 (N_22194,N_21525,N_21839);
and U22195 (N_22195,N_21931,N_21591);
nor U22196 (N_22196,N_21808,N_21630);
nand U22197 (N_22197,N_21992,N_21756);
or U22198 (N_22198,N_21818,N_21534);
and U22199 (N_22199,N_21622,N_21957);
or U22200 (N_22200,N_21517,N_21893);
nor U22201 (N_22201,N_21697,N_21546);
xnor U22202 (N_22202,N_21758,N_21771);
nor U22203 (N_22203,N_21815,N_21584);
nor U22204 (N_22204,N_21672,N_21820);
and U22205 (N_22205,N_21993,N_21581);
nand U22206 (N_22206,N_21799,N_21595);
nor U22207 (N_22207,N_21509,N_21753);
nand U22208 (N_22208,N_21510,N_21979);
and U22209 (N_22209,N_21785,N_21568);
or U22210 (N_22210,N_21867,N_21561);
nand U22211 (N_22211,N_21728,N_21520);
nor U22212 (N_22212,N_21786,N_21659);
nand U22213 (N_22213,N_21783,N_21825);
nand U22214 (N_22214,N_21716,N_21702);
and U22215 (N_22215,N_21636,N_21958);
or U22216 (N_22216,N_21949,N_21917);
xnor U22217 (N_22217,N_21530,N_21749);
and U22218 (N_22218,N_21612,N_21651);
nor U22219 (N_22219,N_21684,N_21585);
xor U22220 (N_22220,N_21648,N_21727);
nand U22221 (N_22221,N_21985,N_21929);
nand U22222 (N_22222,N_21967,N_21567);
nand U22223 (N_22223,N_21886,N_21875);
nor U22224 (N_22224,N_21997,N_21772);
nand U22225 (N_22225,N_21583,N_21916);
or U22226 (N_22226,N_21868,N_21744);
and U22227 (N_22227,N_21707,N_21582);
nor U22228 (N_22228,N_21563,N_21602);
nand U22229 (N_22229,N_21807,N_21610);
nor U22230 (N_22230,N_21841,N_21723);
nand U22231 (N_22231,N_21514,N_21849);
nor U22232 (N_22232,N_21669,N_21910);
nand U22233 (N_22233,N_21906,N_21861);
nor U22234 (N_22234,N_21972,N_21835);
nor U22235 (N_22235,N_21606,N_21974);
nor U22236 (N_22236,N_21863,N_21633);
or U22237 (N_22237,N_21921,N_21529);
nor U22238 (N_22238,N_21687,N_21803);
or U22239 (N_22239,N_21897,N_21740);
and U22240 (N_22240,N_21962,N_21791);
nand U22241 (N_22241,N_21870,N_21624);
nor U22242 (N_22242,N_21614,N_21620);
xnor U22243 (N_22243,N_21832,N_21890);
nor U22244 (N_22244,N_21984,N_21704);
xor U22245 (N_22245,N_21691,N_21590);
nor U22246 (N_22246,N_21914,N_21615);
nor U22247 (N_22247,N_21715,N_21686);
nand U22248 (N_22248,N_21923,N_21769);
xor U22249 (N_22249,N_21701,N_21773);
and U22250 (N_22250,N_21763,N_21548);
xnor U22251 (N_22251,N_21981,N_21570);
and U22252 (N_22252,N_21921,N_21858);
and U22253 (N_22253,N_21968,N_21617);
nor U22254 (N_22254,N_21682,N_21988);
or U22255 (N_22255,N_21615,N_21543);
or U22256 (N_22256,N_21505,N_21843);
or U22257 (N_22257,N_21843,N_21826);
nor U22258 (N_22258,N_21908,N_21701);
or U22259 (N_22259,N_21559,N_21597);
and U22260 (N_22260,N_21698,N_21844);
or U22261 (N_22261,N_21890,N_21726);
nand U22262 (N_22262,N_21647,N_21884);
or U22263 (N_22263,N_21656,N_21995);
nand U22264 (N_22264,N_21853,N_21836);
or U22265 (N_22265,N_21769,N_21560);
xor U22266 (N_22266,N_21935,N_21912);
or U22267 (N_22267,N_21825,N_21859);
or U22268 (N_22268,N_21878,N_21578);
and U22269 (N_22269,N_21876,N_21821);
nor U22270 (N_22270,N_21945,N_21636);
nor U22271 (N_22271,N_21926,N_21815);
nand U22272 (N_22272,N_21703,N_21944);
and U22273 (N_22273,N_21784,N_21542);
nand U22274 (N_22274,N_21711,N_21918);
or U22275 (N_22275,N_21720,N_21899);
and U22276 (N_22276,N_21765,N_21730);
nand U22277 (N_22277,N_21752,N_21724);
nor U22278 (N_22278,N_21641,N_21739);
or U22279 (N_22279,N_21674,N_21619);
or U22280 (N_22280,N_21526,N_21692);
nand U22281 (N_22281,N_21881,N_21674);
or U22282 (N_22282,N_21936,N_21695);
nor U22283 (N_22283,N_21607,N_21829);
or U22284 (N_22284,N_21966,N_21508);
or U22285 (N_22285,N_21898,N_21765);
xor U22286 (N_22286,N_21813,N_21605);
nor U22287 (N_22287,N_21769,N_21524);
or U22288 (N_22288,N_21715,N_21994);
and U22289 (N_22289,N_21863,N_21947);
xnor U22290 (N_22290,N_21562,N_21978);
nor U22291 (N_22291,N_21566,N_21591);
nand U22292 (N_22292,N_21684,N_21740);
nand U22293 (N_22293,N_21852,N_21910);
or U22294 (N_22294,N_21892,N_21883);
nand U22295 (N_22295,N_21700,N_21599);
and U22296 (N_22296,N_21619,N_21540);
or U22297 (N_22297,N_21592,N_21726);
nand U22298 (N_22298,N_21722,N_21545);
xor U22299 (N_22299,N_21701,N_21652);
nand U22300 (N_22300,N_21781,N_21686);
or U22301 (N_22301,N_21982,N_21723);
or U22302 (N_22302,N_21734,N_21530);
and U22303 (N_22303,N_21769,N_21518);
and U22304 (N_22304,N_21994,N_21843);
and U22305 (N_22305,N_21512,N_21861);
and U22306 (N_22306,N_21660,N_21927);
xor U22307 (N_22307,N_21823,N_21716);
nand U22308 (N_22308,N_21574,N_21799);
nor U22309 (N_22309,N_21944,N_21785);
nand U22310 (N_22310,N_21869,N_21712);
and U22311 (N_22311,N_21559,N_21784);
and U22312 (N_22312,N_21821,N_21725);
or U22313 (N_22313,N_21943,N_21799);
nor U22314 (N_22314,N_21985,N_21713);
nand U22315 (N_22315,N_21635,N_21962);
or U22316 (N_22316,N_21882,N_21785);
or U22317 (N_22317,N_21847,N_21829);
nor U22318 (N_22318,N_21946,N_21739);
or U22319 (N_22319,N_21886,N_21665);
nor U22320 (N_22320,N_21755,N_21741);
and U22321 (N_22321,N_21996,N_21877);
nand U22322 (N_22322,N_21724,N_21857);
or U22323 (N_22323,N_21891,N_21975);
xnor U22324 (N_22324,N_21816,N_21976);
xnor U22325 (N_22325,N_21536,N_21626);
xor U22326 (N_22326,N_21845,N_21585);
or U22327 (N_22327,N_21761,N_21518);
or U22328 (N_22328,N_21723,N_21870);
nor U22329 (N_22329,N_21956,N_21528);
or U22330 (N_22330,N_21609,N_21531);
or U22331 (N_22331,N_21595,N_21896);
nor U22332 (N_22332,N_21864,N_21627);
or U22333 (N_22333,N_21640,N_21528);
and U22334 (N_22334,N_21809,N_21947);
nor U22335 (N_22335,N_21976,N_21744);
nand U22336 (N_22336,N_21843,N_21692);
nor U22337 (N_22337,N_21859,N_21910);
xnor U22338 (N_22338,N_21772,N_21586);
and U22339 (N_22339,N_21972,N_21978);
or U22340 (N_22340,N_21845,N_21843);
or U22341 (N_22341,N_21550,N_21980);
and U22342 (N_22342,N_21859,N_21786);
nand U22343 (N_22343,N_21540,N_21657);
nor U22344 (N_22344,N_21841,N_21691);
nor U22345 (N_22345,N_21844,N_21936);
and U22346 (N_22346,N_21690,N_21909);
or U22347 (N_22347,N_21849,N_21784);
nor U22348 (N_22348,N_21894,N_21768);
nor U22349 (N_22349,N_21825,N_21519);
nand U22350 (N_22350,N_21634,N_21587);
xor U22351 (N_22351,N_21684,N_21963);
nand U22352 (N_22352,N_21512,N_21532);
or U22353 (N_22353,N_21630,N_21659);
nand U22354 (N_22354,N_21685,N_21542);
nor U22355 (N_22355,N_21984,N_21645);
nor U22356 (N_22356,N_21666,N_21537);
or U22357 (N_22357,N_21743,N_21576);
nor U22358 (N_22358,N_21989,N_21697);
nand U22359 (N_22359,N_21887,N_21724);
or U22360 (N_22360,N_21900,N_21672);
and U22361 (N_22361,N_21744,N_21842);
nor U22362 (N_22362,N_21922,N_21576);
nand U22363 (N_22363,N_21730,N_21919);
or U22364 (N_22364,N_21689,N_21609);
nand U22365 (N_22365,N_21852,N_21897);
xnor U22366 (N_22366,N_21754,N_21837);
nor U22367 (N_22367,N_21823,N_21843);
or U22368 (N_22368,N_21960,N_21727);
and U22369 (N_22369,N_21724,N_21791);
nand U22370 (N_22370,N_21874,N_21702);
nand U22371 (N_22371,N_21554,N_21704);
and U22372 (N_22372,N_21711,N_21630);
nor U22373 (N_22373,N_21629,N_21906);
and U22374 (N_22374,N_21605,N_21777);
nor U22375 (N_22375,N_21863,N_21646);
nand U22376 (N_22376,N_21517,N_21673);
and U22377 (N_22377,N_21614,N_21738);
or U22378 (N_22378,N_21745,N_21744);
or U22379 (N_22379,N_21802,N_21845);
nor U22380 (N_22380,N_21555,N_21515);
nand U22381 (N_22381,N_21544,N_21959);
nor U22382 (N_22382,N_21559,N_21764);
nor U22383 (N_22383,N_21682,N_21581);
nand U22384 (N_22384,N_21740,N_21773);
nand U22385 (N_22385,N_21962,N_21727);
or U22386 (N_22386,N_21640,N_21704);
nand U22387 (N_22387,N_21674,N_21916);
and U22388 (N_22388,N_21985,N_21638);
nand U22389 (N_22389,N_21767,N_21845);
nand U22390 (N_22390,N_21677,N_21573);
nand U22391 (N_22391,N_21603,N_21617);
nor U22392 (N_22392,N_21877,N_21960);
and U22393 (N_22393,N_21999,N_21931);
nand U22394 (N_22394,N_21779,N_21807);
or U22395 (N_22395,N_21925,N_21853);
and U22396 (N_22396,N_21714,N_21965);
nand U22397 (N_22397,N_21673,N_21872);
xor U22398 (N_22398,N_21587,N_21549);
nor U22399 (N_22399,N_21508,N_21883);
xnor U22400 (N_22400,N_21516,N_21840);
or U22401 (N_22401,N_21500,N_21958);
nand U22402 (N_22402,N_21793,N_21909);
or U22403 (N_22403,N_21595,N_21519);
nand U22404 (N_22404,N_21891,N_21790);
nand U22405 (N_22405,N_21652,N_21790);
and U22406 (N_22406,N_21710,N_21893);
nand U22407 (N_22407,N_21556,N_21758);
and U22408 (N_22408,N_21727,N_21920);
nor U22409 (N_22409,N_21976,N_21827);
nor U22410 (N_22410,N_21642,N_21865);
nand U22411 (N_22411,N_21927,N_21662);
and U22412 (N_22412,N_21706,N_21828);
xnor U22413 (N_22413,N_21817,N_21970);
nand U22414 (N_22414,N_21910,N_21714);
nor U22415 (N_22415,N_21738,N_21576);
nor U22416 (N_22416,N_21942,N_21818);
and U22417 (N_22417,N_21971,N_21814);
nor U22418 (N_22418,N_21930,N_21747);
or U22419 (N_22419,N_21563,N_21953);
nand U22420 (N_22420,N_21553,N_21583);
nand U22421 (N_22421,N_21806,N_21534);
nand U22422 (N_22422,N_21632,N_21627);
nand U22423 (N_22423,N_21889,N_21773);
or U22424 (N_22424,N_21972,N_21954);
nor U22425 (N_22425,N_21681,N_21839);
nand U22426 (N_22426,N_21946,N_21638);
and U22427 (N_22427,N_21587,N_21644);
or U22428 (N_22428,N_21506,N_21764);
nor U22429 (N_22429,N_21631,N_21919);
or U22430 (N_22430,N_21770,N_21646);
nand U22431 (N_22431,N_21978,N_21938);
nand U22432 (N_22432,N_21693,N_21651);
and U22433 (N_22433,N_21667,N_21948);
xnor U22434 (N_22434,N_21644,N_21700);
nor U22435 (N_22435,N_21933,N_21729);
and U22436 (N_22436,N_21810,N_21936);
nor U22437 (N_22437,N_21795,N_21834);
and U22438 (N_22438,N_21931,N_21853);
nor U22439 (N_22439,N_21988,N_21860);
xnor U22440 (N_22440,N_21923,N_21510);
nand U22441 (N_22441,N_21894,N_21921);
or U22442 (N_22442,N_21593,N_21966);
or U22443 (N_22443,N_21800,N_21853);
xnor U22444 (N_22444,N_21668,N_21901);
nand U22445 (N_22445,N_21915,N_21743);
nand U22446 (N_22446,N_21959,N_21513);
nand U22447 (N_22447,N_21924,N_21950);
and U22448 (N_22448,N_21581,N_21555);
nor U22449 (N_22449,N_21563,N_21862);
nand U22450 (N_22450,N_21650,N_21537);
or U22451 (N_22451,N_21650,N_21846);
nand U22452 (N_22452,N_21969,N_21552);
nand U22453 (N_22453,N_21568,N_21663);
and U22454 (N_22454,N_21797,N_21873);
or U22455 (N_22455,N_21863,N_21735);
and U22456 (N_22456,N_21572,N_21978);
or U22457 (N_22457,N_21572,N_21520);
and U22458 (N_22458,N_21534,N_21673);
nand U22459 (N_22459,N_21682,N_21918);
nor U22460 (N_22460,N_21602,N_21787);
or U22461 (N_22461,N_21580,N_21820);
or U22462 (N_22462,N_21716,N_21607);
nor U22463 (N_22463,N_21588,N_21802);
nand U22464 (N_22464,N_21590,N_21729);
and U22465 (N_22465,N_21579,N_21620);
nand U22466 (N_22466,N_21778,N_21751);
nand U22467 (N_22467,N_21816,N_21533);
and U22468 (N_22468,N_21806,N_21657);
and U22469 (N_22469,N_21737,N_21793);
nor U22470 (N_22470,N_21959,N_21670);
nor U22471 (N_22471,N_21775,N_21635);
and U22472 (N_22472,N_21543,N_21577);
xor U22473 (N_22473,N_21650,N_21999);
nor U22474 (N_22474,N_21695,N_21923);
nor U22475 (N_22475,N_21809,N_21605);
nand U22476 (N_22476,N_21668,N_21973);
nand U22477 (N_22477,N_21692,N_21920);
or U22478 (N_22478,N_21827,N_21960);
and U22479 (N_22479,N_21627,N_21894);
xnor U22480 (N_22480,N_21721,N_21761);
and U22481 (N_22481,N_21840,N_21996);
nand U22482 (N_22482,N_21641,N_21828);
or U22483 (N_22483,N_21700,N_21666);
or U22484 (N_22484,N_21616,N_21703);
and U22485 (N_22485,N_21717,N_21803);
or U22486 (N_22486,N_21964,N_21877);
nor U22487 (N_22487,N_21837,N_21662);
or U22488 (N_22488,N_21636,N_21850);
and U22489 (N_22489,N_21589,N_21753);
xnor U22490 (N_22490,N_21950,N_21826);
nor U22491 (N_22491,N_21957,N_21795);
and U22492 (N_22492,N_21953,N_21551);
or U22493 (N_22493,N_21545,N_21937);
and U22494 (N_22494,N_21872,N_21928);
nand U22495 (N_22495,N_21978,N_21574);
nand U22496 (N_22496,N_21571,N_21889);
nand U22497 (N_22497,N_21693,N_21866);
or U22498 (N_22498,N_21633,N_21924);
nor U22499 (N_22499,N_21674,N_21733);
and U22500 (N_22500,N_22032,N_22085);
nor U22501 (N_22501,N_22102,N_22248);
or U22502 (N_22502,N_22250,N_22275);
and U22503 (N_22503,N_22489,N_22361);
or U22504 (N_22504,N_22016,N_22186);
or U22505 (N_22505,N_22445,N_22075);
or U22506 (N_22506,N_22055,N_22111);
nor U22507 (N_22507,N_22135,N_22197);
and U22508 (N_22508,N_22137,N_22217);
and U22509 (N_22509,N_22313,N_22004);
nor U22510 (N_22510,N_22292,N_22149);
and U22511 (N_22511,N_22079,N_22230);
and U22512 (N_22512,N_22009,N_22373);
or U22513 (N_22513,N_22067,N_22118);
nand U22514 (N_22514,N_22179,N_22383);
and U22515 (N_22515,N_22439,N_22254);
and U22516 (N_22516,N_22277,N_22065);
and U22517 (N_22517,N_22286,N_22060);
and U22518 (N_22518,N_22043,N_22478);
nand U22519 (N_22519,N_22435,N_22064);
or U22520 (N_22520,N_22037,N_22068);
and U22521 (N_22521,N_22307,N_22044);
and U22522 (N_22522,N_22334,N_22425);
nand U22523 (N_22523,N_22207,N_22433);
nand U22524 (N_22524,N_22295,N_22341);
nor U22525 (N_22525,N_22110,N_22348);
and U22526 (N_22526,N_22192,N_22430);
nand U22527 (N_22527,N_22368,N_22495);
nor U22528 (N_22528,N_22183,N_22443);
and U22529 (N_22529,N_22029,N_22306);
nor U22530 (N_22530,N_22208,N_22265);
nor U22531 (N_22531,N_22132,N_22237);
nor U22532 (N_22532,N_22235,N_22142);
or U22533 (N_22533,N_22491,N_22317);
and U22534 (N_22534,N_22176,N_22301);
nor U22535 (N_22535,N_22427,N_22473);
nand U22536 (N_22536,N_22063,N_22018);
nor U22537 (N_22537,N_22048,N_22402);
or U22538 (N_22538,N_22423,N_22136);
nand U22539 (N_22539,N_22087,N_22083);
nor U22540 (N_22540,N_22177,N_22471);
nor U22541 (N_22541,N_22028,N_22369);
or U22542 (N_22542,N_22020,N_22167);
nor U22543 (N_22543,N_22010,N_22349);
nand U22544 (N_22544,N_22239,N_22131);
nor U22545 (N_22545,N_22093,N_22145);
nor U22546 (N_22546,N_22338,N_22394);
nand U22547 (N_22547,N_22030,N_22271);
xor U22548 (N_22548,N_22357,N_22143);
and U22549 (N_22549,N_22127,N_22095);
nand U22550 (N_22550,N_22246,N_22360);
xor U22551 (N_22551,N_22469,N_22304);
and U22552 (N_22552,N_22314,N_22257);
nor U22553 (N_22553,N_22094,N_22023);
nor U22554 (N_22554,N_22448,N_22232);
and U22555 (N_22555,N_22310,N_22129);
and U22556 (N_22556,N_22008,N_22199);
nor U22557 (N_22557,N_22464,N_22399);
nor U22558 (N_22558,N_22178,N_22125);
xor U22559 (N_22559,N_22412,N_22276);
nand U22560 (N_22560,N_22355,N_22291);
or U22561 (N_22561,N_22293,N_22320);
and U22562 (N_22562,N_22024,N_22057);
nand U22563 (N_22563,N_22077,N_22461);
xor U22564 (N_22564,N_22409,N_22168);
or U22565 (N_22565,N_22336,N_22106);
and U22566 (N_22566,N_22185,N_22052);
and U22567 (N_22567,N_22269,N_22258);
or U22568 (N_22568,N_22418,N_22326);
and U22569 (N_22569,N_22196,N_22162);
nand U22570 (N_22570,N_22468,N_22283);
nand U22571 (N_22571,N_22463,N_22115);
and U22572 (N_22572,N_22014,N_22263);
and U22573 (N_22573,N_22034,N_22475);
nand U22574 (N_22574,N_22128,N_22352);
and U22575 (N_22575,N_22108,N_22488);
nand U22576 (N_22576,N_22410,N_22419);
and U22577 (N_22577,N_22172,N_22203);
or U22578 (N_22578,N_22157,N_22003);
or U22579 (N_22579,N_22450,N_22302);
nand U22580 (N_22580,N_22090,N_22000);
nand U22581 (N_22581,N_22353,N_22001);
nor U22582 (N_22582,N_22021,N_22156);
or U22583 (N_22583,N_22496,N_22038);
nor U22584 (N_22584,N_22025,N_22026);
and U22585 (N_22585,N_22432,N_22447);
and U22586 (N_22586,N_22340,N_22289);
and U22587 (N_22587,N_22190,N_22012);
nand U22588 (N_22588,N_22017,N_22103);
or U22589 (N_22589,N_22296,N_22243);
nor U22590 (N_22590,N_22411,N_22241);
and U22591 (N_22591,N_22392,N_22272);
and U22592 (N_22592,N_22315,N_22174);
nor U22593 (N_22593,N_22031,N_22238);
and U22594 (N_22594,N_22195,N_22245);
xnor U22595 (N_22595,N_22362,N_22184);
nor U22596 (N_22596,N_22456,N_22226);
or U22597 (N_22597,N_22138,N_22282);
nand U22598 (N_22598,N_22163,N_22462);
and U22599 (N_22599,N_22072,N_22221);
xor U22600 (N_22600,N_22170,N_22091);
nand U22601 (N_22601,N_22204,N_22007);
nand U22602 (N_22602,N_22354,N_22255);
xnor U22603 (N_22603,N_22401,N_22273);
or U22604 (N_22604,N_22122,N_22161);
or U22605 (N_22605,N_22387,N_22414);
nand U22606 (N_22606,N_22390,N_22346);
nor U22607 (N_22607,N_22405,N_22069);
or U22608 (N_22608,N_22180,N_22490);
and U22609 (N_22609,N_22049,N_22499);
and U22610 (N_22610,N_22147,N_22398);
nor U22611 (N_22611,N_22139,N_22242);
or U22612 (N_22612,N_22486,N_22374);
or U22613 (N_22613,N_22465,N_22449);
or U22614 (N_22614,N_22116,N_22487);
and U22615 (N_22615,N_22059,N_22454);
xor U22616 (N_22616,N_22153,N_22074);
xor U22617 (N_22617,N_22329,N_22251);
and U22618 (N_22618,N_22481,N_22019);
or U22619 (N_22619,N_22056,N_22497);
and U22620 (N_22620,N_22260,N_22287);
or U22621 (N_22621,N_22222,N_22218);
and U22622 (N_22622,N_22121,N_22047);
nor U22623 (N_22623,N_22407,N_22188);
and U22624 (N_22624,N_22482,N_22393);
or U22625 (N_22625,N_22078,N_22231);
or U22626 (N_22626,N_22321,N_22363);
nand U22627 (N_22627,N_22191,N_22022);
or U22628 (N_22628,N_22215,N_22460);
xnor U22629 (N_22629,N_22073,N_22385);
xnor U22630 (N_22630,N_22331,N_22485);
or U22631 (N_22631,N_22466,N_22080);
nand U22632 (N_22632,N_22367,N_22112);
and U22633 (N_22633,N_22396,N_22337);
and U22634 (N_22634,N_22268,N_22333);
and U22635 (N_22635,N_22324,N_22290);
or U22636 (N_22636,N_22384,N_22274);
xnor U22637 (N_22637,N_22437,N_22434);
nand U22638 (N_22638,N_22339,N_22366);
nor U22639 (N_22639,N_22446,N_22438);
and U22640 (N_22640,N_22327,N_22416);
or U22641 (N_22641,N_22299,N_22294);
and U22642 (N_22642,N_22388,N_22216);
and U22643 (N_22643,N_22041,N_22229);
nor U22644 (N_22644,N_22467,N_22259);
nand U22645 (N_22645,N_22046,N_22300);
or U22646 (N_22646,N_22279,N_22050);
and U22647 (N_22647,N_22494,N_22051);
or U22648 (N_22648,N_22380,N_22408);
and U22649 (N_22649,N_22479,N_22311);
nand U22650 (N_22650,N_22201,N_22126);
and U22651 (N_22651,N_22035,N_22422);
nor U22652 (N_22652,N_22305,N_22459);
nor U22653 (N_22653,N_22205,N_22330);
and U22654 (N_22654,N_22160,N_22428);
or U22655 (N_22655,N_22099,N_22148);
or U22656 (N_22656,N_22200,N_22270);
nor U22657 (N_22657,N_22084,N_22406);
nand U22658 (N_22658,N_22426,N_22236);
or U22659 (N_22659,N_22264,N_22134);
or U22660 (N_22660,N_22480,N_22011);
nand U22661 (N_22661,N_22391,N_22261);
and U22662 (N_22662,N_22097,N_22364);
or U22663 (N_22663,N_22061,N_22442);
and U22664 (N_22664,N_22140,N_22104);
or U22665 (N_22665,N_22284,N_22013);
or U22666 (N_22666,N_22451,N_22070);
and U22667 (N_22667,N_22206,N_22212);
nor U22668 (N_22668,N_22440,N_22002);
nor U22669 (N_22669,N_22303,N_22472);
nand U22670 (N_22670,N_22164,N_22249);
and U22671 (N_22671,N_22417,N_22123);
nand U22672 (N_22672,N_22114,N_22082);
xor U22673 (N_22673,N_22359,N_22493);
or U22674 (N_22674,N_22458,N_22244);
xnor U22675 (N_22675,N_22345,N_22171);
nor U22676 (N_22676,N_22088,N_22133);
nor U22677 (N_22677,N_22006,N_22308);
and U22678 (N_22678,N_22344,N_22223);
and U22679 (N_22679,N_22444,N_22150);
or U22680 (N_22680,N_22220,N_22389);
or U22681 (N_22681,N_22086,N_22198);
nand U22682 (N_22682,N_22247,N_22358);
nor U22683 (N_22683,N_22395,N_22042);
and U22684 (N_22684,N_22318,N_22397);
and U22685 (N_22685,N_22347,N_22159);
and U22686 (N_22686,N_22285,N_22240);
nor U22687 (N_22687,N_22076,N_22421);
nor U22688 (N_22688,N_22228,N_22413);
and U22689 (N_22689,N_22092,N_22202);
nor U22690 (N_22690,N_22098,N_22066);
and U22691 (N_22691,N_22288,N_22144);
and U22692 (N_22692,N_22370,N_22100);
nand U22693 (N_22693,N_22151,N_22256);
nor U22694 (N_22694,N_22312,N_22262);
nand U22695 (N_22695,N_22120,N_22350);
or U22696 (N_22696,N_22379,N_22053);
and U22697 (N_22697,N_22400,N_22278);
nand U22698 (N_22698,N_22483,N_22266);
nand U22699 (N_22699,N_22470,N_22209);
and U22700 (N_22700,N_22252,N_22477);
nand U22701 (N_22701,N_22130,N_22498);
or U22702 (N_22702,N_22297,N_22173);
nor U22703 (N_22703,N_22280,N_22429);
xor U22704 (N_22704,N_22081,N_22058);
and U22705 (N_22705,N_22211,N_22323);
nand U22706 (N_22706,N_22154,N_22219);
nand U22707 (N_22707,N_22381,N_22193);
xor U22708 (N_22708,N_22033,N_22182);
nor U22709 (N_22709,N_22351,N_22071);
nand U22710 (N_22710,N_22062,N_22403);
nor U22711 (N_22711,N_22169,N_22325);
nor U22712 (N_22712,N_22141,N_22453);
and U22713 (N_22713,N_22455,N_22005);
or U22714 (N_22714,N_22332,N_22015);
nor U22715 (N_22715,N_22328,N_22152);
and U22716 (N_22716,N_22227,N_22214);
or U22717 (N_22717,N_22124,N_22371);
nand U22718 (N_22718,N_22210,N_22105);
nor U22719 (N_22719,N_22036,N_22420);
nand U22720 (N_22720,N_22343,N_22234);
or U22721 (N_22721,N_22158,N_22378);
xnor U22722 (N_22722,N_22484,N_22372);
and U22723 (N_22723,N_22213,N_22404);
xor U22724 (N_22724,N_22054,N_22233);
or U22725 (N_22725,N_22424,N_22146);
nand U22726 (N_22726,N_22117,N_22319);
and U22727 (N_22727,N_22187,N_22101);
or U22728 (N_22728,N_22096,N_22027);
nor U22729 (N_22729,N_22492,N_22342);
nor U22730 (N_22730,N_22382,N_22166);
nor U22731 (N_22731,N_22253,N_22045);
xnor U22732 (N_22732,N_22457,N_22436);
xnor U22733 (N_22733,N_22441,N_22322);
nor U22734 (N_22734,N_22107,N_22431);
nor U22735 (N_22735,N_22298,N_22474);
nand U22736 (N_22736,N_22375,N_22089);
nor U22737 (N_22737,N_22039,N_22109);
nand U22738 (N_22738,N_22224,N_22267);
xnor U22739 (N_22739,N_22309,N_22165);
xnor U22740 (N_22740,N_22281,N_22175);
nor U22741 (N_22741,N_22189,N_22113);
nand U22742 (N_22742,N_22119,N_22181);
or U22743 (N_22743,N_22365,N_22476);
or U22744 (N_22744,N_22194,N_22356);
or U22745 (N_22745,N_22415,N_22335);
or U22746 (N_22746,N_22386,N_22316);
nand U22747 (N_22747,N_22040,N_22452);
xnor U22748 (N_22748,N_22225,N_22155);
nor U22749 (N_22749,N_22376,N_22377);
and U22750 (N_22750,N_22009,N_22197);
nor U22751 (N_22751,N_22000,N_22385);
nor U22752 (N_22752,N_22132,N_22344);
and U22753 (N_22753,N_22214,N_22298);
nand U22754 (N_22754,N_22384,N_22208);
nand U22755 (N_22755,N_22075,N_22265);
xor U22756 (N_22756,N_22267,N_22450);
or U22757 (N_22757,N_22207,N_22469);
xnor U22758 (N_22758,N_22405,N_22342);
and U22759 (N_22759,N_22011,N_22061);
nor U22760 (N_22760,N_22170,N_22317);
and U22761 (N_22761,N_22341,N_22466);
nand U22762 (N_22762,N_22115,N_22347);
or U22763 (N_22763,N_22390,N_22199);
and U22764 (N_22764,N_22364,N_22458);
nand U22765 (N_22765,N_22057,N_22027);
and U22766 (N_22766,N_22348,N_22463);
or U22767 (N_22767,N_22202,N_22420);
xor U22768 (N_22768,N_22491,N_22031);
nand U22769 (N_22769,N_22081,N_22034);
nand U22770 (N_22770,N_22482,N_22305);
xor U22771 (N_22771,N_22005,N_22113);
nor U22772 (N_22772,N_22486,N_22330);
nor U22773 (N_22773,N_22001,N_22160);
nor U22774 (N_22774,N_22281,N_22025);
nor U22775 (N_22775,N_22358,N_22086);
nand U22776 (N_22776,N_22041,N_22328);
nor U22777 (N_22777,N_22261,N_22395);
or U22778 (N_22778,N_22418,N_22091);
or U22779 (N_22779,N_22426,N_22167);
xnor U22780 (N_22780,N_22480,N_22363);
nor U22781 (N_22781,N_22175,N_22129);
or U22782 (N_22782,N_22235,N_22342);
nand U22783 (N_22783,N_22478,N_22227);
nand U22784 (N_22784,N_22266,N_22044);
nand U22785 (N_22785,N_22043,N_22454);
nor U22786 (N_22786,N_22099,N_22035);
nor U22787 (N_22787,N_22196,N_22198);
nor U22788 (N_22788,N_22432,N_22088);
nor U22789 (N_22789,N_22391,N_22216);
nor U22790 (N_22790,N_22312,N_22206);
or U22791 (N_22791,N_22273,N_22344);
or U22792 (N_22792,N_22443,N_22028);
nor U22793 (N_22793,N_22088,N_22360);
xnor U22794 (N_22794,N_22314,N_22413);
xnor U22795 (N_22795,N_22204,N_22060);
or U22796 (N_22796,N_22307,N_22259);
nand U22797 (N_22797,N_22359,N_22131);
nand U22798 (N_22798,N_22177,N_22008);
and U22799 (N_22799,N_22113,N_22307);
xor U22800 (N_22800,N_22380,N_22185);
nand U22801 (N_22801,N_22278,N_22367);
or U22802 (N_22802,N_22119,N_22312);
nor U22803 (N_22803,N_22426,N_22325);
and U22804 (N_22804,N_22211,N_22193);
nor U22805 (N_22805,N_22169,N_22434);
or U22806 (N_22806,N_22226,N_22098);
nand U22807 (N_22807,N_22254,N_22498);
and U22808 (N_22808,N_22191,N_22249);
nor U22809 (N_22809,N_22039,N_22328);
and U22810 (N_22810,N_22040,N_22189);
nand U22811 (N_22811,N_22487,N_22274);
xor U22812 (N_22812,N_22074,N_22180);
nor U22813 (N_22813,N_22063,N_22120);
or U22814 (N_22814,N_22352,N_22356);
xnor U22815 (N_22815,N_22231,N_22279);
nand U22816 (N_22816,N_22404,N_22349);
or U22817 (N_22817,N_22163,N_22347);
or U22818 (N_22818,N_22181,N_22458);
or U22819 (N_22819,N_22295,N_22021);
or U22820 (N_22820,N_22440,N_22221);
or U22821 (N_22821,N_22114,N_22052);
or U22822 (N_22822,N_22091,N_22089);
nand U22823 (N_22823,N_22228,N_22005);
and U22824 (N_22824,N_22285,N_22158);
nand U22825 (N_22825,N_22205,N_22274);
and U22826 (N_22826,N_22135,N_22055);
or U22827 (N_22827,N_22155,N_22493);
or U22828 (N_22828,N_22451,N_22073);
nor U22829 (N_22829,N_22434,N_22174);
nand U22830 (N_22830,N_22176,N_22048);
and U22831 (N_22831,N_22237,N_22124);
xor U22832 (N_22832,N_22074,N_22019);
or U22833 (N_22833,N_22404,N_22217);
nand U22834 (N_22834,N_22250,N_22134);
or U22835 (N_22835,N_22331,N_22147);
nand U22836 (N_22836,N_22450,N_22113);
nor U22837 (N_22837,N_22174,N_22024);
nand U22838 (N_22838,N_22430,N_22233);
and U22839 (N_22839,N_22331,N_22431);
and U22840 (N_22840,N_22420,N_22449);
or U22841 (N_22841,N_22482,N_22142);
nand U22842 (N_22842,N_22209,N_22116);
xnor U22843 (N_22843,N_22454,N_22211);
and U22844 (N_22844,N_22006,N_22485);
nor U22845 (N_22845,N_22030,N_22335);
nor U22846 (N_22846,N_22071,N_22098);
nor U22847 (N_22847,N_22145,N_22224);
nand U22848 (N_22848,N_22256,N_22279);
nand U22849 (N_22849,N_22126,N_22157);
xor U22850 (N_22850,N_22105,N_22073);
nand U22851 (N_22851,N_22091,N_22413);
xor U22852 (N_22852,N_22196,N_22452);
nor U22853 (N_22853,N_22110,N_22053);
xnor U22854 (N_22854,N_22388,N_22199);
nand U22855 (N_22855,N_22195,N_22227);
or U22856 (N_22856,N_22143,N_22354);
or U22857 (N_22857,N_22488,N_22297);
nor U22858 (N_22858,N_22365,N_22456);
and U22859 (N_22859,N_22258,N_22432);
or U22860 (N_22860,N_22459,N_22301);
nand U22861 (N_22861,N_22495,N_22231);
xnor U22862 (N_22862,N_22489,N_22469);
and U22863 (N_22863,N_22472,N_22481);
or U22864 (N_22864,N_22426,N_22332);
nand U22865 (N_22865,N_22378,N_22104);
nand U22866 (N_22866,N_22063,N_22203);
nand U22867 (N_22867,N_22487,N_22255);
nor U22868 (N_22868,N_22221,N_22069);
and U22869 (N_22869,N_22064,N_22170);
nand U22870 (N_22870,N_22219,N_22046);
and U22871 (N_22871,N_22207,N_22242);
or U22872 (N_22872,N_22249,N_22323);
nor U22873 (N_22873,N_22424,N_22475);
nand U22874 (N_22874,N_22435,N_22346);
nor U22875 (N_22875,N_22464,N_22435);
and U22876 (N_22876,N_22264,N_22433);
nand U22877 (N_22877,N_22279,N_22402);
and U22878 (N_22878,N_22041,N_22227);
nand U22879 (N_22879,N_22447,N_22254);
or U22880 (N_22880,N_22099,N_22492);
nor U22881 (N_22881,N_22184,N_22048);
and U22882 (N_22882,N_22082,N_22465);
nand U22883 (N_22883,N_22451,N_22329);
nor U22884 (N_22884,N_22170,N_22076);
or U22885 (N_22885,N_22252,N_22063);
nand U22886 (N_22886,N_22425,N_22025);
nor U22887 (N_22887,N_22291,N_22192);
nor U22888 (N_22888,N_22096,N_22246);
or U22889 (N_22889,N_22020,N_22302);
and U22890 (N_22890,N_22498,N_22313);
or U22891 (N_22891,N_22487,N_22459);
and U22892 (N_22892,N_22200,N_22466);
or U22893 (N_22893,N_22459,N_22447);
nor U22894 (N_22894,N_22360,N_22250);
and U22895 (N_22895,N_22323,N_22246);
and U22896 (N_22896,N_22339,N_22108);
nor U22897 (N_22897,N_22273,N_22319);
or U22898 (N_22898,N_22014,N_22462);
nand U22899 (N_22899,N_22445,N_22262);
and U22900 (N_22900,N_22025,N_22102);
nand U22901 (N_22901,N_22064,N_22153);
and U22902 (N_22902,N_22131,N_22253);
nand U22903 (N_22903,N_22184,N_22137);
or U22904 (N_22904,N_22466,N_22060);
or U22905 (N_22905,N_22060,N_22101);
xnor U22906 (N_22906,N_22012,N_22350);
or U22907 (N_22907,N_22175,N_22043);
nand U22908 (N_22908,N_22294,N_22475);
nand U22909 (N_22909,N_22380,N_22280);
nor U22910 (N_22910,N_22162,N_22475);
nor U22911 (N_22911,N_22437,N_22409);
and U22912 (N_22912,N_22073,N_22337);
or U22913 (N_22913,N_22392,N_22138);
nor U22914 (N_22914,N_22380,N_22445);
or U22915 (N_22915,N_22143,N_22458);
and U22916 (N_22916,N_22036,N_22424);
and U22917 (N_22917,N_22223,N_22260);
nand U22918 (N_22918,N_22432,N_22313);
and U22919 (N_22919,N_22026,N_22340);
nor U22920 (N_22920,N_22430,N_22107);
xnor U22921 (N_22921,N_22099,N_22322);
or U22922 (N_22922,N_22258,N_22434);
nor U22923 (N_22923,N_22158,N_22157);
nor U22924 (N_22924,N_22338,N_22156);
nor U22925 (N_22925,N_22457,N_22237);
nand U22926 (N_22926,N_22165,N_22142);
nor U22927 (N_22927,N_22179,N_22283);
and U22928 (N_22928,N_22367,N_22168);
or U22929 (N_22929,N_22478,N_22152);
nand U22930 (N_22930,N_22176,N_22453);
nand U22931 (N_22931,N_22366,N_22297);
nand U22932 (N_22932,N_22228,N_22326);
and U22933 (N_22933,N_22441,N_22485);
and U22934 (N_22934,N_22024,N_22195);
and U22935 (N_22935,N_22083,N_22171);
nand U22936 (N_22936,N_22260,N_22060);
nand U22937 (N_22937,N_22426,N_22045);
nor U22938 (N_22938,N_22077,N_22151);
xor U22939 (N_22939,N_22354,N_22274);
and U22940 (N_22940,N_22283,N_22214);
or U22941 (N_22941,N_22342,N_22372);
nand U22942 (N_22942,N_22492,N_22299);
or U22943 (N_22943,N_22435,N_22280);
or U22944 (N_22944,N_22257,N_22356);
nand U22945 (N_22945,N_22145,N_22436);
nand U22946 (N_22946,N_22325,N_22461);
nor U22947 (N_22947,N_22054,N_22274);
nor U22948 (N_22948,N_22454,N_22487);
or U22949 (N_22949,N_22289,N_22299);
nand U22950 (N_22950,N_22124,N_22395);
xor U22951 (N_22951,N_22366,N_22492);
nor U22952 (N_22952,N_22086,N_22304);
xnor U22953 (N_22953,N_22238,N_22077);
nor U22954 (N_22954,N_22171,N_22469);
and U22955 (N_22955,N_22496,N_22321);
or U22956 (N_22956,N_22219,N_22403);
xor U22957 (N_22957,N_22155,N_22202);
or U22958 (N_22958,N_22343,N_22247);
nand U22959 (N_22959,N_22437,N_22138);
or U22960 (N_22960,N_22324,N_22303);
nor U22961 (N_22961,N_22284,N_22021);
nor U22962 (N_22962,N_22490,N_22498);
or U22963 (N_22963,N_22306,N_22083);
or U22964 (N_22964,N_22442,N_22076);
nand U22965 (N_22965,N_22009,N_22450);
or U22966 (N_22966,N_22305,N_22168);
xor U22967 (N_22967,N_22380,N_22206);
nand U22968 (N_22968,N_22249,N_22204);
or U22969 (N_22969,N_22329,N_22272);
nor U22970 (N_22970,N_22152,N_22416);
xor U22971 (N_22971,N_22038,N_22392);
or U22972 (N_22972,N_22145,N_22208);
xnor U22973 (N_22973,N_22489,N_22270);
nand U22974 (N_22974,N_22106,N_22137);
nor U22975 (N_22975,N_22393,N_22165);
nand U22976 (N_22976,N_22014,N_22472);
nor U22977 (N_22977,N_22262,N_22313);
or U22978 (N_22978,N_22185,N_22440);
and U22979 (N_22979,N_22025,N_22115);
nand U22980 (N_22980,N_22147,N_22086);
and U22981 (N_22981,N_22031,N_22222);
nor U22982 (N_22982,N_22469,N_22404);
and U22983 (N_22983,N_22367,N_22105);
or U22984 (N_22984,N_22134,N_22431);
nand U22985 (N_22985,N_22144,N_22361);
xnor U22986 (N_22986,N_22222,N_22093);
nor U22987 (N_22987,N_22261,N_22272);
and U22988 (N_22988,N_22363,N_22413);
xor U22989 (N_22989,N_22147,N_22194);
nor U22990 (N_22990,N_22015,N_22195);
nand U22991 (N_22991,N_22441,N_22397);
nor U22992 (N_22992,N_22322,N_22186);
and U22993 (N_22993,N_22385,N_22466);
nor U22994 (N_22994,N_22473,N_22250);
nor U22995 (N_22995,N_22377,N_22385);
and U22996 (N_22996,N_22146,N_22292);
and U22997 (N_22997,N_22180,N_22471);
nand U22998 (N_22998,N_22078,N_22463);
nand U22999 (N_22999,N_22268,N_22276);
nand U23000 (N_23000,N_22697,N_22991);
and U23001 (N_23001,N_22717,N_22768);
nand U23002 (N_23002,N_22985,N_22605);
and U23003 (N_23003,N_22807,N_22892);
nor U23004 (N_23004,N_22908,N_22635);
nor U23005 (N_23005,N_22535,N_22804);
xor U23006 (N_23006,N_22563,N_22537);
nor U23007 (N_23007,N_22658,N_22874);
or U23008 (N_23008,N_22728,N_22968);
xor U23009 (N_23009,N_22770,N_22591);
and U23010 (N_23010,N_22707,N_22637);
and U23011 (N_23011,N_22611,N_22771);
and U23012 (N_23012,N_22622,N_22730);
and U23013 (N_23013,N_22789,N_22967);
or U23014 (N_23014,N_22671,N_22850);
and U23015 (N_23015,N_22833,N_22696);
or U23016 (N_23016,N_22872,N_22931);
xnor U23017 (N_23017,N_22932,N_22693);
or U23018 (N_23018,N_22513,N_22935);
and U23019 (N_23019,N_22746,N_22667);
and U23020 (N_23020,N_22787,N_22761);
nor U23021 (N_23021,N_22673,N_22737);
nor U23022 (N_23022,N_22661,N_22982);
nand U23023 (N_23023,N_22792,N_22900);
or U23024 (N_23024,N_22940,N_22589);
and U23025 (N_23025,N_22758,N_22674);
or U23026 (N_23026,N_22934,N_22799);
nand U23027 (N_23027,N_22554,N_22839);
and U23028 (N_23028,N_22654,N_22569);
xnor U23029 (N_23029,N_22953,N_22992);
nor U23030 (N_23030,N_22918,N_22690);
nor U23031 (N_23031,N_22677,N_22639);
or U23032 (N_23032,N_22902,N_22972);
or U23033 (N_23033,N_22765,N_22885);
nand U23034 (N_23034,N_22733,N_22561);
xor U23035 (N_23035,N_22757,N_22579);
nor U23036 (N_23036,N_22905,N_22855);
nand U23037 (N_23037,N_22689,N_22996);
nand U23038 (N_23038,N_22656,N_22847);
nand U23039 (N_23039,N_22676,N_22582);
nor U23040 (N_23040,N_22816,N_22861);
nor U23041 (N_23041,N_22539,N_22538);
nor U23042 (N_23042,N_22781,N_22973);
or U23043 (N_23043,N_22565,N_22809);
or U23044 (N_23044,N_22692,N_22526);
and U23045 (N_23045,N_22662,N_22887);
nor U23046 (N_23046,N_22923,N_22525);
nor U23047 (N_23047,N_22503,N_22597);
or U23048 (N_23048,N_22753,N_22927);
nor U23049 (N_23049,N_22558,N_22740);
nor U23050 (N_23050,N_22650,N_22655);
nand U23051 (N_23051,N_22783,N_22851);
nand U23052 (N_23052,N_22632,N_22718);
nand U23053 (N_23053,N_22846,N_22866);
xor U23054 (N_23054,N_22623,N_22977);
or U23055 (N_23055,N_22549,N_22803);
nand U23056 (N_23056,N_22610,N_22575);
xor U23057 (N_23057,N_22980,N_22741);
nand U23058 (N_23058,N_22506,N_22628);
and U23059 (N_23059,N_22911,N_22971);
or U23060 (N_23060,N_22772,N_22723);
nand U23061 (N_23061,N_22581,N_22750);
nand U23062 (N_23062,N_22536,N_22556);
nand U23063 (N_23063,N_22557,N_22668);
nand U23064 (N_23064,N_22684,N_22725);
nor U23065 (N_23065,N_22785,N_22821);
nand U23066 (N_23066,N_22744,N_22859);
nand U23067 (N_23067,N_22913,N_22864);
nor U23068 (N_23068,N_22815,N_22598);
or U23069 (N_23069,N_22638,N_22642);
nand U23070 (N_23070,N_22898,N_22606);
nor U23071 (N_23071,N_22801,N_22854);
or U23072 (N_23072,N_22921,N_22688);
and U23073 (N_23073,N_22865,N_22954);
nor U23074 (N_23074,N_22548,N_22641);
nand U23075 (N_23075,N_22883,N_22949);
nand U23076 (N_23076,N_22621,N_22564);
and U23077 (N_23077,N_22822,N_22834);
and U23078 (N_23078,N_22594,N_22670);
and U23079 (N_23079,N_22832,N_22615);
xnor U23080 (N_23080,N_22587,N_22876);
nor U23081 (N_23081,N_22517,N_22577);
nor U23082 (N_23082,N_22604,N_22736);
or U23083 (N_23083,N_22760,N_22508);
or U23084 (N_23084,N_22666,N_22708);
and U23085 (N_23085,N_22559,N_22997);
xnor U23086 (N_23086,N_22648,N_22889);
or U23087 (N_23087,N_22720,N_22919);
nor U23088 (N_23088,N_22995,N_22748);
nor U23089 (N_23089,N_22511,N_22906);
or U23090 (N_23090,N_22749,N_22586);
nand U23091 (N_23091,N_22867,N_22820);
nor U23092 (N_23092,N_22827,N_22555);
and U23093 (N_23093,N_22780,N_22626);
or U23094 (N_23094,N_22532,N_22520);
or U23095 (N_23095,N_22798,N_22607);
nor U23096 (N_23096,N_22726,N_22814);
or U23097 (N_23097,N_22766,N_22659);
nand U23098 (N_23098,N_22546,N_22672);
or U23099 (N_23099,N_22956,N_22849);
or U23100 (N_23100,N_22620,N_22764);
and U23101 (N_23101,N_22735,N_22826);
or U23102 (N_23102,N_22779,N_22875);
and U23103 (N_23103,N_22584,N_22619);
nand U23104 (N_23104,N_22522,N_22888);
or U23105 (N_23105,N_22544,N_22886);
and U23106 (N_23106,N_22570,N_22974);
and U23107 (N_23107,N_22975,N_22592);
nand U23108 (N_23108,N_22938,N_22928);
nor U23109 (N_23109,N_22710,N_22961);
nand U23110 (N_23110,N_22527,N_22574);
and U23111 (N_23111,N_22794,N_22682);
nor U23112 (N_23112,N_22614,N_22602);
nor U23113 (N_23113,N_22802,N_22942);
xnor U23114 (N_23114,N_22773,N_22685);
or U23115 (N_23115,N_22640,N_22657);
nand U23116 (N_23116,N_22683,N_22912);
and U23117 (N_23117,N_22817,N_22633);
xor U23118 (N_23118,N_22808,N_22578);
nand U23119 (N_23119,N_22848,N_22989);
nor U23120 (N_23120,N_22857,N_22862);
or U23121 (N_23121,N_22599,N_22796);
and U23122 (N_23122,N_22560,N_22810);
xnor U23123 (N_23123,N_22930,N_22836);
nor U23124 (N_23124,N_22825,N_22791);
nand U23125 (N_23125,N_22695,N_22660);
and U23126 (N_23126,N_22553,N_22743);
or U23127 (N_23127,N_22925,N_22722);
nand U23128 (N_23128,N_22944,N_22873);
and U23129 (N_23129,N_22813,N_22501);
nor U23130 (N_23130,N_22739,N_22646);
xor U23131 (N_23131,N_22812,N_22617);
and U23132 (N_23132,N_22616,N_22649);
nand U23133 (N_23133,N_22790,N_22533);
nand U23134 (N_23134,N_22981,N_22519);
and U23135 (N_23135,N_22751,N_22551);
nor U23136 (N_23136,N_22647,N_22528);
and U23137 (N_23137,N_22922,N_22829);
or U23138 (N_23138,N_22784,N_22521);
nor U23139 (N_23139,N_22881,N_22715);
nand U23140 (N_23140,N_22856,N_22515);
or U23141 (N_23141,N_22711,N_22776);
or U23142 (N_23142,N_22915,N_22531);
nor U23143 (N_23143,N_22745,N_22524);
nand U23144 (N_23144,N_22706,N_22727);
and U23145 (N_23145,N_22669,N_22734);
and U23146 (N_23146,N_22665,N_22907);
xor U23147 (N_23147,N_22600,N_22958);
nor U23148 (N_23148,N_22567,N_22845);
or U23149 (N_23149,N_22613,N_22651);
and U23150 (N_23150,N_22686,N_22568);
xnor U23151 (N_23151,N_22878,N_22762);
or U23152 (N_23152,N_22652,N_22719);
and U23153 (N_23153,N_22868,N_22699);
and U23154 (N_23154,N_22800,N_22767);
nor U23155 (N_23155,N_22920,N_22716);
and U23156 (N_23156,N_22926,N_22724);
or U23157 (N_23157,N_22644,N_22863);
nor U23158 (N_23158,N_22988,N_22998);
nand U23159 (N_23159,N_22609,N_22679);
nor U23160 (N_23160,N_22844,N_22562);
and U23161 (N_23161,N_22608,N_22512);
nand U23162 (N_23162,N_22732,N_22694);
nor U23163 (N_23163,N_22964,N_22755);
or U23164 (N_23164,N_22774,N_22712);
nand U23165 (N_23165,N_22534,N_22946);
nand U23166 (N_23166,N_22747,N_22583);
and U23167 (N_23167,N_22593,N_22970);
nand U23168 (N_23168,N_22899,N_22976);
xnor U23169 (N_23169,N_22952,N_22951);
nor U23170 (N_23170,N_22987,N_22993);
nand U23171 (N_23171,N_22763,N_22819);
nand U23172 (N_23172,N_22704,N_22675);
nand U23173 (N_23173,N_22653,N_22818);
nand U23174 (N_23174,N_22933,N_22843);
nor U23175 (N_23175,N_22738,N_22663);
or U23176 (N_23176,N_22978,N_22870);
xnor U23177 (N_23177,N_22937,N_22754);
nand U23178 (N_23178,N_22729,N_22838);
xnor U23179 (N_23179,N_22523,N_22957);
nor U23180 (N_23180,N_22590,N_22896);
nor U23181 (N_23181,N_22955,N_22778);
or U23182 (N_23182,N_22645,N_22909);
and U23183 (N_23183,N_22837,N_22631);
and U23184 (N_23184,N_22880,N_22860);
nand U23185 (N_23185,N_22786,N_22596);
xor U23186 (N_23186,N_22835,N_22500);
or U23187 (N_23187,N_22571,N_22945);
xor U23188 (N_23188,N_22936,N_22550);
and U23189 (N_23189,N_22756,N_22959);
nor U23190 (N_23190,N_22904,N_22731);
nor U23191 (N_23191,N_22601,N_22721);
or U23192 (N_23192,N_22687,N_22573);
nand U23193 (N_23193,N_22547,N_22680);
or U23194 (N_23194,N_22769,N_22929);
nand U23195 (N_23195,N_22540,N_22999);
nand U23196 (N_23196,N_22705,N_22782);
or U23197 (N_23197,N_22884,N_22947);
or U23198 (N_23198,N_22914,N_22831);
nor U23199 (N_23199,N_22624,N_22984);
nor U23200 (N_23200,N_22823,N_22924);
or U23201 (N_23201,N_22529,N_22806);
xor U23202 (N_23202,N_22797,N_22950);
and U23203 (N_23203,N_22903,N_22702);
xnor U23204 (N_23204,N_22618,N_22542);
nand U23205 (N_23205,N_22897,N_22939);
or U23206 (N_23206,N_22552,N_22703);
nand U23207 (N_23207,N_22795,N_22853);
nor U23208 (N_23208,N_22828,N_22509);
nand U23209 (N_23209,N_22681,N_22948);
nand U23210 (N_23210,N_22603,N_22983);
nor U23211 (N_23211,N_22830,N_22510);
or U23212 (N_23212,N_22858,N_22916);
nor U23213 (N_23213,N_22516,N_22709);
nand U23214 (N_23214,N_22910,N_22759);
or U23215 (N_23215,N_22879,N_22960);
or U23216 (N_23216,N_22585,N_22505);
or U23217 (N_23217,N_22901,N_22518);
xnor U23218 (N_23218,N_22698,N_22842);
and U23219 (N_23219,N_22541,N_22852);
or U23220 (N_23220,N_22700,N_22871);
and U23221 (N_23221,N_22788,N_22893);
or U23222 (N_23222,N_22580,N_22986);
xor U23223 (N_23223,N_22965,N_22514);
and U23224 (N_23224,N_22530,N_22576);
nand U23225 (N_23225,N_22941,N_22502);
nor U23226 (N_23226,N_22917,N_22625);
and U23227 (N_23227,N_22811,N_22627);
nand U23228 (N_23228,N_22636,N_22566);
nor U23229 (N_23229,N_22841,N_22994);
or U23230 (N_23230,N_22890,N_22877);
nand U23231 (N_23231,N_22691,N_22664);
nand U23232 (N_23232,N_22643,N_22840);
nor U23233 (N_23233,N_22894,N_22543);
nand U23234 (N_23234,N_22714,N_22629);
and U23235 (N_23235,N_22990,N_22742);
and U23236 (N_23236,N_22775,N_22824);
xnor U23237 (N_23237,N_22943,N_22966);
xor U23238 (N_23238,N_22630,N_22882);
xor U23239 (N_23239,N_22869,N_22963);
nor U23240 (N_23240,N_22805,N_22777);
and U23241 (N_23241,N_22678,N_22507);
or U23242 (N_23242,N_22545,N_22572);
and U23243 (N_23243,N_22969,N_22962);
nor U23244 (N_23244,N_22612,N_22634);
or U23245 (N_23245,N_22701,N_22595);
and U23246 (N_23246,N_22979,N_22752);
nor U23247 (N_23247,N_22713,N_22504);
or U23248 (N_23248,N_22793,N_22895);
or U23249 (N_23249,N_22891,N_22588);
nand U23250 (N_23250,N_22874,N_22635);
nor U23251 (N_23251,N_22640,N_22506);
nor U23252 (N_23252,N_22745,N_22800);
nand U23253 (N_23253,N_22842,N_22853);
and U23254 (N_23254,N_22678,N_22564);
or U23255 (N_23255,N_22894,N_22868);
or U23256 (N_23256,N_22579,N_22935);
and U23257 (N_23257,N_22639,N_22560);
nor U23258 (N_23258,N_22628,N_22968);
nand U23259 (N_23259,N_22816,N_22945);
nor U23260 (N_23260,N_22999,N_22779);
nor U23261 (N_23261,N_22817,N_22814);
nor U23262 (N_23262,N_22567,N_22944);
nor U23263 (N_23263,N_22573,N_22893);
nor U23264 (N_23264,N_22794,N_22613);
and U23265 (N_23265,N_22835,N_22658);
nor U23266 (N_23266,N_22588,N_22938);
nand U23267 (N_23267,N_22661,N_22515);
or U23268 (N_23268,N_22755,N_22987);
nor U23269 (N_23269,N_22960,N_22689);
xnor U23270 (N_23270,N_22898,N_22640);
and U23271 (N_23271,N_22651,N_22570);
nor U23272 (N_23272,N_22934,N_22798);
and U23273 (N_23273,N_22941,N_22660);
nand U23274 (N_23274,N_22763,N_22929);
or U23275 (N_23275,N_22539,N_22810);
and U23276 (N_23276,N_22996,N_22529);
nand U23277 (N_23277,N_22983,N_22991);
and U23278 (N_23278,N_22835,N_22884);
or U23279 (N_23279,N_22656,N_22919);
nand U23280 (N_23280,N_22799,N_22668);
nand U23281 (N_23281,N_22564,N_22697);
nor U23282 (N_23282,N_22979,N_22967);
nand U23283 (N_23283,N_22732,N_22852);
and U23284 (N_23284,N_22947,N_22558);
nor U23285 (N_23285,N_22766,N_22805);
and U23286 (N_23286,N_22845,N_22610);
nor U23287 (N_23287,N_22611,N_22913);
nand U23288 (N_23288,N_22763,N_22736);
and U23289 (N_23289,N_22968,N_22540);
or U23290 (N_23290,N_22883,N_22664);
xnor U23291 (N_23291,N_22922,N_22789);
nor U23292 (N_23292,N_22866,N_22742);
nor U23293 (N_23293,N_22774,N_22517);
nand U23294 (N_23294,N_22691,N_22591);
nand U23295 (N_23295,N_22511,N_22527);
or U23296 (N_23296,N_22858,N_22999);
or U23297 (N_23297,N_22853,N_22727);
or U23298 (N_23298,N_22832,N_22555);
nor U23299 (N_23299,N_22965,N_22799);
and U23300 (N_23300,N_22957,N_22654);
xnor U23301 (N_23301,N_22747,N_22546);
or U23302 (N_23302,N_22549,N_22700);
and U23303 (N_23303,N_22586,N_22838);
and U23304 (N_23304,N_22601,N_22618);
nor U23305 (N_23305,N_22799,N_22518);
nor U23306 (N_23306,N_22538,N_22691);
or U23307 (N_23307,N_22806,N_22664);
and U23308 (N_23308,N_22915,N_22938);
and U23309 (N_23309,N_22539,N_22812);
or U23310 (N_23310,N_22660,N_22743);
and U23311 (N_23311,N_22967,N_22570);
nor U23312 (N_23312,N_22830,N_22777);
and U23313 (N_23313,N_22594,N_22607);
xnor U23314 (N_23314,N_22627,N_22894);
xor U23315 (N_23315,N_22955,N_22794);
and U23316 (N_23316,N_22913,N_22886);
nand U23317 (N_23317,N_22766,N_22903);
nor U23318 (N_23318,N_22905,N_22718);
xor U23319 (N_23319,N_22999,N_22910);
and U23320 (N_23320,N_22536,N_22657);
and U23321 (N_23321,N_22830,N_22773);
and U23322 (N_23322,N_22802,N_22958);
and U23323 (N_23323,N_22855,N_22780);
nor U23324 (N_23324,N_22634,N_22907);
nor U23325 (N_23325,N_22816,N_22860);
nor U23326 (N_23326,N_22685,N_22646);
or U23327 (N_23327,N_22808,N_22932);
and U23328 (N_23328,N_22985,N_22850);
nand U23329 (N_23329,N_22699,N_22828);
or U23330 (N_23330,N_22533,N_22569);
or U23331 (N_23331,N_22862,N_22744);
nor U23332 (N_23332,N_22985,N_22736);
nor U23333 (N_23333,N_22575,N_22711);
or U23334 (N_23334,N_22595,N_22755);
and U23335 (N_23335,N_22788,N_22507);
xor U23336 (N_23336,N_22929,N_22517);
or U23337 (N_23337,N_22597,N_22978);
nand U23338 (N_23338,N_22837,N_22808);
nor U23339 (N_23339,N_22775,N_22888);
or U23340 (N_23340,N_22567,N_22728);
and U23341 (N_23341,N_22801,N_22618);
xnor U23342 (N_23342,N_22687,N_22912);
or U23343 (N_23343,N_22904,N_22863);
or U23344 (N_23344,N_22947,N_22581);
and U23345 (N_23345,N_22975,N_22823);
or U23346 (N_23346,N_22826,N_22878);
nand U23347 (N_23347,N_22951,N_22935);
nor U23348 (N_23348,N_22935,N_22786);
nor U23349 (N_23349,N_22555,N_22596);
and U23350 (N_23350,N_22813,N_22643);
or U23351 (N_23351,N_22752,N_22837);
or U23352 (N_23352,N_22584,N_22763);
nand U23353 (N_23353,N_22939,N_22895);
nand U23354 (N_23354,N_22772,N_22556);
nand U23355 (N_23355,N_22627,N_22645);
or U23356 (N_23356,N_22885,N_22942);
and U23357 (N_23357,N_22897,N_22698);
nand U23358 (N_23358,N_22889,N_22693);
nand U23359 (N_23359,N_22726,N_22651);
or U23360 (N_23360,N_22864,N_22665);
or U23361 (N_23361,N_22938,N_22981);
nand U23362 (N_23362,N_22645,N_22926);
nor U23363 (N_23363,N_22666,N_22931);
nand U23364 (N_23364,N_22585,N_22873);
and U23365 (N_23365,N_22955,N_22715);
and U23366 (N_23366,N_22739,N_22825);
nor U23367 (N_23367,N_22676,N_22701);
nand U23368 (N_23368,N_22931,N_22982);
and U23369 (N_23369,N_22542,N_22716);
xnor U23370 (N_23370,N_22800,N_22831);
and U23371 (N_23371,N_22871,N_22645);
or U23372 (N_23372,N_22525,N_22644);
or U23373 (N_23373,N_22571,N_22705);
nor U23374 (N_23374,N_22657,N_22704);
and U23375 (N_23375,N_22718,N_22696);
or U23376 (N_23376,N_22556,N_22929);
or U23377 (N_23377,N_22598,N_22972);
nand U23378 (N_23378,N_22587,N_22917);
nand U23379 (N_23379,N_22888,N_22946);
or U23380 (N_23380,N_22684,N_22687);
and U23381 (N_23381,N_22591,N_22853);
and U23382 (N_23382,N_22571,N_22917);
nor U23383 (N_23383,N_22734,N_22522);
and U23384 (N_23384,N_22683,N_22725);
nand U23385 (N_23385,N_22781,N_22920);
xnor U23386 (N_23386,N_22956,N_22633);
nor U23387 (N_23387,N_22535,N_22505);
or U23388 (N_23388,N_22550,N_22932);
nor U23389 (N_23389,N_22971,N_22892);
xor U23390 (N_23390,N_22803,N_22544);
nand U23391 (N_23391,N_22929,N_22649);
nor U23392 (N_23392,N_22566,N_22531);
and U23393 (N_23393,N_22739,N_22976);
nor U23394 (N_23394,N_22982,N_22751);
xnor U23395 (N_23395,N_22983,N_22523);
nand U23396 (N_23396,N_22888,N_22935);
and U23397 (N_23397,N_22811,N_22527);
nor U23398 (N_23398,N_22649,N_22638);
xor U23399 (N_23399,N_22737,N_22548);
nor U23400 (N_23400,N_22567,N_22871);
and U23401 (N_23401,N_22951,N_22941);
xnor U23402 (N_23402,N_22680,N_22697);
and U23403 (N_23403,N_22534,N_22984);
nand U23404 (N_23404,N_22794,N_22501);
nand U23405 (N_23405,N_22804,N_22787);
xnor U23406 (N_23406,N_22511,N_22982);
nor U23407 (N_23407,N_22534,N_22942);
and U23408 (N_23408,N_22716,N_22811);
or U23409 (N_23409,N_22628,N_22907);
xnor U23410 (N_23410,N_22528,N_22771);
nor U23411 (N_23411,N_22665,N_22791);
nand U23412 (N_23412,N_22924,N_22819);
xnor U23413 (N_23413,N_22818,N_22587);
nand U23414 (N_23414,N_22560,N_22617);
or U23415 (N_23415,N_22790,N_22631);
nor U23416 (N_23416,N_22943,N_22927);
nand U23417 (N_23417,N_22828,N_22893);
and U23418 (N_23418,N_22886,N_22683);
or U23419 (N_23419,N_22544,N_22696);
or U23420 (N_23420,N_22888,N_22994);
and U23421 (N_23421,N_22882,N_22707);
or U23422 (N_23422,N_22811,N_22636);
nor U23423 (N_23423,N_22583,N_22561);
nand U23424 (N_23424,N_22714,N_22776);
nor U23425 (N_23425,N_22633,N_22806);
nor U23426 (N_23426,N_22773,N_22612);
and U23427 (N_23427,N_22882,N_22568);
or U23428 (N_23428,N_22694,N_22582);
and U23429 (N_23429,N_22599,N_22941);
and U23430 (N_23430,N_22855,N_22505);
nor U23431 (N_23431,N_22778,N_22986);
and U23432 (N_23432,N_22605,N_22586);
nand U23433 (N_23433,N_22992,N_22750);
or U23434 (N_23434,N_22838,N_22818);
nand U23435 (N_23435,N_22942,N_22833);
and U23436 (N_23436,N_22707,N_22675);
or U23437 (N_23437,N_22641,N_22595);
and U23438 (N_23438,N_22613,N_22866);
or U23439 (N_23439,N_22661,N_22639);
nor U23440 (N_23440,N_22898,N_22619);
or U23441 (N_23441,N_22925,N_22682);
xor U23442 (N_23442,N_22814,N_22654);
and U23443 (N_23443,N_22977,N_22651);
nor U23444 (N_23444,N_22944,N_22508);
or U23445 (N_23445,N_22836,N_22748);
and U23446 (N_23446,N_22899,N_22792);
and U23447 (N_23447,N_22803,N_22852);
nand U23448 (N_23448,N_22804,N_22826);
nand U23449 (N_23449,N_22692,N_22819);
and U23450 (N_23450,N_22718,N_22791);
nor U23451 (N_23451,N_22630,N_22539);
nand U23452 (N_23452,N_22556,N_22859);
nor U23453 (N_23453,N_22664,N_22574);
xnor U23454 (N_23454,N_22688,N_22931);
or U23455 (N_23455,N_22836,N_22975);
nand U23456 (N_23456,N_22590,N_22895);
or U23457 (N_23457,N_22717,N_22512);
nor U23458 (N_23458,N_22770,N_22972);
nand U23459 (N_23459,N_22944,N_22829);
and U23460 (N_23460,N_22623,N_22737);
or U23461 (N_23461,N_22521,N_22737);
nand U23462 (N_23462,N_22507,N_22888);
nand U23463 (N_23463,N_22719,N_22852);
or U23464 (N_23464,N_22817,N_22958);
xnor U23465 (N_23465,N_22651,N_22740);
or U23466 (N_23466,N_22664,N_22735);
nor U23467 (N_23467,N_22623,N_22886);
nand U23468 (N_23468,N_22923,N_22898);
xor U23469 (N_23469,N_22725,N_22563);
and U23470 (N_23470,N_22735,N_22796);
and U23471 (N_23471,N_22640,N_22674);
nor U23472 (N_23472,N_22536,N_22990);
nor U23473 (N_23473,N_22893,N_22823);
or U23474 (N_23474,N_22792,N_22973);
nor U23475 (N_23475,N_22541,N_22773);
or U23476 (N_23476,N_22973,N_22937);
nand U23477 (N_23477,N_22526,N_22889);
and U23478 (N_23478,N_22933,N_22519);
nand U23479 (N_23479,N_22956,N_22585);
nand U23480 (N_23480,N_22781,N_22546);
nand U23481 (N_23481,N_22911,N_22661);
or U23482 (N_23482,N_22963,N_22723);
xor U23483 (N_23483,N_22986,N_22866);
or U23484 (N_23484,N_22978,N_22935);
or U23485 (N_23485,N_22770,N_22822);
or U23486 (N_23486,N_22748,N_22553);
or U23487 (N_23487,N_22956,N_22589);
or U23488 (N_23488,N_22913,N_22931);
and U23489 (N_23489,N_22519,N_22673);
or U23490 (N_23490,N_22998,N_22659);
and U23491 (N_23491,N_22701,N_22508);
or U23492 (N_23492,N_22606,N_22621);
nor U23493 (N_23493,N_22566,N_22743);
nand U23494 (N_23494,N_22662,N_22921);
nand U23495 (N_23495,N_22524,N_22677);
and U23496 (N_23496,N_22801,N_22883);
and U23497 (N_23497,N_22686,N_22514);
nor U23498 (N_23498,N_22697,N_22519);
and U23499 (N_23499,N_22889,N_22981);
nor U23500 (N_23500,N_23013,N_23303);
nor U23501 (N_23501,N_23166,N_23210);
and U23502 (N_23502,N_23353,N_23358);
nand U23503 (N_23503,N_23459,N_23361);
and U23504 (N_23504,N_23338,N_23054);
and U23505 (N_23505,N_23229,N_23474);
and U23506 (N_23506,N_23335,N_23016);
and U23507 (N_23507,N_23266,N_23235);
or U23508 (N_23508,N_23135,N_23379);
and U23509 (N_23509,N_23094,N_23035);
or U23510 (N_23510,N_23370,N_23351);
or U23511 (N_23511,N_23136,N_23195);
nor U23512 (N_23512,N_23364,N_23374);
and U23513 (N_23513,N_23243,N_23072);
or U23514 (N_23514,N_23423,N_23125);
or U23515 (N_23515,N_23393,N_23022);
xor U23516 (N_23516,N_23402,N_23213);
xor U23517 (N_23517,N_23205,N_23167);
nor U23518 (N_23518,N_23133,N_23148);
or U23519 (N_23519,N_23162,N_23071);
xor U23520 (N_23520,N_23105,N_23174);
xnor U23521 (N_23521,N_23040,N_23108);
or U23522 (N_23522,N_23089,N_23350);
or U23523 (N_23523,N_23065,N_23051);
and U23524 (N_23524,N_23420,N_23339);
or U23525 (N_23525,N_23170,N_23258);
nand U23526 (N_23526,N_23029,N_23319);
nor U23527 (N_23527,N_23486,N_23406);
nand U23528 (N_23528,N_23302,N_23285);
and U23529 (N_23529,N_23287,N_23346);
and U23530 (N_23530,N_23091,N_23134);
nand U23531 (N_23531,N_23396,N_23454);
or U23532 (N_23532,N_23099,N_23087);
nor U23533 (N_23533,N_23308,N_23069);
and U23534 (N_23534,N_23033,N_23063);
nor U23535 (N_23535,N_23100,N_23057);
and U23536 (N_23536,N_23360,N_23297);
nor U23537 (N_23537,N_23427,N_23276);
or U23538 (N_23538,N_23124,N_23356);
nand U23539 (N_23539,N_23321,N_23218);
nand U23540 (N_23540,N_23220,N_23048);
xor U23541 (N_23541,N_23467,N_23000);
nor U23542 (N_23542,N_23242,N_23192);
or U23543 (N_23543,N_23375,N_23263);
nor U23544 (N_23544,N_23155,N_23324);
and U23545 (N_23545,N_23096,N_23158);
nand U23546 (N_23546,N_23415,N_23140);
and U23547 (N_23547,N_23267,N_23281);
and U23548 (N_23548,N_23481,N_23095);
xor U23549 (N_23549,N_23203,N_23221);
or U23550 (N_23550,N_23104,N_23286);
and U23551 (N_23551,N_23132,N_23139);
and U23552 (N_23552,N_23190,N_23183);
nand U23553 (N_23553,N_23008,N_23495);
nor U23554 (N_23554,N_23288,N_23046);
and U23555 (N_23555,N_23426,N_23431);
nor U23556 (N_23556,N_23330,N_23097);
and U23557 (N_23557,N_23389,N_23270);
or U23558 (N_23558,N_23362,N_23386);
or U23559 (N_23559,N_23280,N_23015);
nor U23560 (N_23560,N_23007,N_23066);
and U23561 (N_23561,N_23416,N_23068);
nand U23562 (N_23562,N_23489,N_23122);
and U23563 (N_23563,N_23172,N_23202);
nand U23564 (N_23564,N_23469,N_23373);
xor U23565 (N_23565,N_23241,N_23143);
or U23566 (N_23566,N_23298,N_23391);
nand U23567 (N_23567,N_23200,N_23049);
nand U23568 (N_23568,N_23392,N_23471);
and U23569 (N_23569,N_23014,N_23106);
and U23570 (N_23570,N_23020,N_23043);
nand U23571 (N_23571,N_23357,N_23231);
nand U23572 (N_23572,N_23225,N_23333);
nor U23573 (N_23573,N_23309,N_23484);
or U23574 (N_23574,N_23145,N_23451);
nor U23575 (N_23575,N_23282,N_23291);
nor U23576 (N_23576,N_23304,N_23211);
nand U23577 (N_23577,N_23400,N_23146);
or U23578 (N_23578,N_23249,N_23073);
nor U23579 (N_23579,N_23448,N_23003);
nor U23580 (N_23580,N_23156,N_23337);
or U23581 (N_23581,N_23111,N_23058);
xor U23582 (N_23582,N_23317,N_23077);
and U23583 (N_23583,N_23409,N_23300);
and U23584 (N_23584,N_23296,N_23488);
nand U23585 (N_23585,N_23314,N_23163);
or U23586 (N_23586,N_23463,N_23318);
nor U23587 (N_23587,N_23452,N_23446);
nand U23588 (N_23588,N_23034,N_23215);
nand U23589 (N_23589,N_23045,N_23418);
nor U23590 (N_23590,N_23176,N_23305);
or U23591 (N_23591,N_23395,N_23376);
or U23592 (N_23592,N_23227,N_23354);
or U23593 (N_23593,N_23347,N_23457);
nor U23594 (N_23594,N_23327,N_23107);
nand U23595 (N_23595,N_23310,N_23271);
nor U23596 (N_23596,N_23175,N_23115);
and U23597 (N_23597,N_23284,N_23038);
and U23598 (N_23598,N_23342,N_23160);
or U23599 (N_23599,N_23414,N_23161);
nor U23600 (N_23600,N_23252,N_23432);
and U23601 (N_23601,N_23344,N_23447);
or U23602 (N_23602,N_23425,N_23422);
xor U23603 (N_23603,N_23178,N_23385);
xor U23604 (N_23604,N_23320,N_23401);
nand U23605 (N_23605,N_23259,N_23059);
or U23606 (N_23606,N_23397,N_23247);
nor U23607 (N_23607,N_23265,N_23329);
and U23608 (N_23608,N_23490,N_23365);
nor U23609 (N_23609,N_23199,N_23256);
and U23610 (N_23610,N_23430,N_23149);
nor U23611 (N_23611,N_23331,N_23336);
or U23612 (N_23612,N_23023,N_23042);
nand U23613 (N_23613,N_23212,N_23117);
nor U23614 (N_23614,N_23372,N_23261);
xnor U23615 (N_23615,N_23475,N_23387);
nand U23616 (N_23616,N_23173,N_23110);
nor U23617 (N_23617,N_23398,N_23348);
nand U23618 (N_23618,N_23466,N_23408);
nand U23619 (N_23619,N_23449,N_23165);
or U23620 (N_23620,N_23483,N_23237);
nor U23621 (N_23621,N_23157,N_23204);
and U23622 (N_23622,N_23381,N_23301);
or U23623 (N_23623,N_23223,N_23315);
nor U23624 (N_23624,N_23141,N_23487);
nor U23625 (N_23625,N_23001,N_23299);
or U23626 (N_23626,N_23456,N_23150);
and U23627 (N_23627,N_23368,N_23470);
or U23628 (N_23628,N_23179,N_23277);
and U23629 (N_23629,N_23080,N_23472);
nor U23630 (N_23630,N_23193,N_23168);
and U23631 (N_23631,N_23450,N_23292);
nand U23632 (N_23632,N_23030,N_23436);
xnor U23633 (N_23633,N_23419,N_23260);
nor U23634 (N_23634,N_23055,N_23206);
and U23635 (N_23635,N_23112,N_23369);
nand U23636 (N_23636,N_23118,N_23109);
nor U23637 (N_23637,N_23036,N_23222);
and U23638 (N_23638,N_23371,N_23061);
nor U23639 (N_23639,N_23274,N_23006);
nor U23640 (N_23640,N_23198,N_23289);
and U23641 (N_23641,N_23144,N_23005);
nor U23642 (N_23642,N_23191,N_23186);
nor U23643 (N_23643,N_23011,N_23151);
nor U23644 (N_23644,N_23154,N_23041);
nor U23645 (N_23645,N_23230,N_23208);
nor U23646 (N_23646,N_23088,N_23214);
or U23647 (N_23647,N_23120,N_23142);
nor U23648 (N_23648,N_23273,N_23429);
nor U23649 (N_23649,N_23209,N_23224);
nor U23650 (N_23650,N_23159,N_23238);
xnor U23651 (N_23651,N_23403,N_23216);
nand U23652 (N_23652,N_23445,N_23349);
nor U23653 (N_23653,N_23119,N_23332);
and U23654 (N_23654,N_23283,N_23064);
or U23655 (N_23655,N_23442,N_23384);
nand U23656 (N_23656,N_23441,N_23473);
or U23657 (N_23657,N_23184,N_23152);
or U23658 (N_23658,N_23207,N_23443);
or U23659 (N_23659,N_23239,N_23233);
nand U23660 (N_23660,N_23102,N_23017);
nand U23661 (N_23661,N_23078,N_23334);
and U23662 (N_23662,N_23312,N_23462);
nand U23663 (N_23663,N_23464,N_23056);
or U23664 (N_23664,N_23411,N_23126);
nor U23665 (N_23665,N_23367,N_23031);
and U23666 (N_23666,N_23116,N_23026);
xnor U23667 (N_23667,N_23460,N_23024);
nor U23668 (N_23668,N_23131,N_23421);
nand U23669 (N_23669,N_23485,N_23380);
nor U23670 (N_23670,N_23465,N_23121);
and U23671 (N_23671,N_23009,N_23081);
xnor U23672 (N_23672,N_23293,N_23188);
nor U23673 (N_23673,N_23458,N_23130);
or U23674 (N_23674,N_23478,N_23453);
and U23675 (N_23675,N_23477,N_23164);
or U23676 (N_23676,N_23295,N_23366);
nor U23677 (N_23677,N_23086,N_23412);
xor U23678 (N_23678,N_23187,N_23294);
nand U23679 (N_23679,N_23468,N_23434);
nand U23680 (N_23680,N_23169,N_23245);
nand U23681 (N_23681,N_23232,N_23062);
and U23682 (N_23682,N_23019,N_23083);
xnor U23683 (N_23683,N_23098,N_23196);
nand U23684 (N_23684,N_23246,N_23407);
or U23685 (N_23685,N_23345,N_23128);
nand U23686 (N_23686,N_23405,N_23383);
nor U23687 (N_23687,N_23359,N_23410);
nor U23688 (N_23688,N_23092,N_23114);
or U23689 (N_23689,N_23067,N_23404);
xnor U23690 (N_23690,N_23244,N_23388);
or U23691 (N_23691,N_23326,N_23461);
and U23692 (N_23692,N_23085,N_23090);
or U23693 (N_23693,N_23047,N_23240);
and U23694 (N_23694,N_23053,N_23343);
or U23695 (N_23695,N_23497,N_23076);
nor U23696 (N_23696,N_23363,N_23440);
nand U23697 (N_23697,N_23181,N_23306);
or U23698 (N_23698,N_23010,N_23194);
or U23699 (N_23699,N_23437,N_23093);
nor U23700 (N_23700,N_23251,N_23004);
or U23701 (N_23701,N_23328,N_23275);
and U23702 (N_23702,N_23262,N_23044);
nor U23703 (N_23703,N_23079,N_23253);
and U23704 (N_23704,N_23438,N_23248);
and U23705 (N_23705,N_23254,N_23236);
and U23706 (N_23706,N_23137,N_23413);
nor U23707 (N_23707,N_23268,N_23390);
and U23708 (N_23708,N_23226,N_23084);
nand U23709 (N_23709,N_23482,N_23075);
and U23710 (N_23710,N_23494,N_23219);
xor U23711 (N_23711,N_23060,N_23428);
and U23712 (N_23712,N_23018,N_23127);
nor U23713 (N_23713,N_23323,N_23234);
or U23714 (N_23714,N_23032,N_23250);
xnor U23715 (N_23715,N_23352,N_23340);
nor U23716 (N_23716,N_23129,N_23355);
nor U23717 (N_23717,N_23382,N_23480);
nand U23718 (N_23718,N_23037,N_23050);
and U23719 (N_23719,N_23439,N_23417);
and U23720 (N_23720,N_23307,N_23290);
nand U23721 (N_23721,N_23269,N_23185);
nand U23722 (N_23722,N_23378,N_23264);
or U23723 (N_23723,N_23272,N_23491);
or U23724 (N_23724,N_23498,N_23316);
or U23725 (N_23725,N_23123,N_23171);
nor U23726 (N_23726,N_23201,N_23025);
or U23727 (N_23727,N_23002,N_23492);
nand U23728 (N_23728,N_23435,N_23341);
xnor U23729 (N_23729,N_23228,N_23074);
or U23730 (N_23730,N_23279,N_23444);
or U23731 (N_23731,N_23082,N_23325);
nor U23732 (N_23732,N_23257,N_23496);
and U23733 (N_23733,N_23394,N_23153);
nand U23734 (N_23734,N_23455,N_23052);
and U23735 (N_23735,N_23433,N_23424);
nor U23736 (N_23736,N_23101,N_23476);
or U23737 (N_23737,N_23197,N_23499);
or U23738 (N_23738,N_23147,N_23313);
nor U23739 (N_23739,N_23377,N_23278);
or U23740 (N_23740,N_23322,N_23182);
nand U23741 (N_23741,N_23138,N_23103);
or U23742 (N_23742,N_23027,N_23189);
and U23743 (N_23743,N_23255,N_23028);
nor U23744 (N_23744,N_23012,N_23113);
nor U23745 (N_23745,N_23039,N_23070);
and U23746 (N_23746,N_23180,N_23493);
nor U23747 (N_23747,N_23177,N_23311);
or U23748 (N_23748,N_23217,N_23021);
nand U23749 (N_23749,N_23399,N_23479);
and U23750 (N_23750,N_23252,N_23196);
and U23751 (N_23751,N_23210,N_23306);
and U23752 (N_23752,N_23455,N_23299);
nand U23753 (N_23753,N_23102,N_23412);
xnor U23754 (N_23754,N_23424,N_23227);
nor U23755 (N_23755,N_23199,N_23369);
nor U23756 (N_23756,N_23303,N_23318);
nor U23757 (N_23757,N_23209,N_23269);
and U23758 (N_23758,N_23263,N_23276);
and U23759 (N_23759,N_23062,N_23233);
or U23760 (N_23760,N_23315,N_23073);
and U23761 (N_23761,N_23036,N_23289);
xor U23762 (N_23762,N_23139,N_23362);
or U23763 (N_23763,N_23439,N_23164);
and U23764 (N_23764,N_23460,N_23400);
nor U23765 (N_23765,N_23283,N_23305);
or U23766 (N_23766,N_23089,N_23065);
or U23767 (N_23767,N_23278,N_23339);
and U23768 (N_23768,N_23209,N_23148);
or U23769 (N_23769,N_23415,N_23463);
xnor U23770 (N_23770,N_23180,N_23436);
xor U23771 (N_23771,N_23439,N_23308);
xnor U23772 (N_23772,N_23491,N_23276);
nor U23773 (N_23773,N_23285,N_23310);
and U23774 (N_23774,N_23427,N_23203);
and U23775 (N_23775,N_23156,N_23068);
and U23776 (N_23776,N_23143,N_23081);
nand U23777 (N_23777,N_23355,N_23376);
xnor U23778 (N_23778,N_23107,N_23119);
nand U23779 (N_23779,N_23304,N_23149);
nor U23780 (N_23780,N_23014,N_23398);
nand U23781 (N_23781,N_23439,N_23051);
and U23782 (N_23782,N_23155,N_23086);
nand U23783 (N_23783,N_23349,N_23024);
nand U23784 (N_23784,N_23489,N_23328);
nand U23785 (N_23785,N_23251,N_23397);
or U23786 (N_23786,N_23431,N_23092);
and U23787 (N_23787,N_23319,N_23198);
or U23788 (N_23788,N_23080,N_23324);
nand U23789 (N_23789,N_23025,N_23194);
and U23790 (N_23790,N_23463,N_23091);
and U23791 (N_23791,N_23040,N_23198);
or U23792 (N_23792,N_23003,N_23145);
and U23793 (N_23793,N_23041,N_23034);
or U23794 (N_23794,N_23074,N_23335);
nand U23795 (N_23795,N_23143,N_23244);
and U23796 (N_23796,N_23283,N_23150);
xor U23797 (N_23797,N_23406,N_23412);
nand U23798 (N_23798,N_23455,N_23063);
or U23799 (N_23799,N_23266,N_23289);
xnor U23800 (N_23800,N_23310,N_23388);
or U23801 (N_23801,N_23221,N_23295);
and U23802 (N_23802,N_23443,N_23215);
or U23803 (N_23803,N_23444,N_23287);
and U23804 (N_23804,N_23215,N_23020);
or U23805 (N_23805,N_23038,N_23240);
nor U23806 (N_23806,N_23494,N_23349);
nor U23807 (N_23807,N_23329,N_23248);
and U23808 (N_23808,N_23178,N_23031);
or U23809 (N_23809,N_23168,N_23020);
nand U23810 (N_23810,N_23149,N_23104);
or U23811 (N_23811,N_23224,N_23259);
nor U23812 (N_23812,N_23324,N_23369);
and U23813 (N_23813,N_23303,N_23184);
nand U23814 (N_23814,N_23290,N_23014);
nand U23815 (N_23815,N_23103,N_23299);
or U23816 (N_23816,N_23041,N_23144);
nand U23817 (N_23817,N_23037,N_23167);
nor U23818 (N_23818,N_23018,N_23185);
nor U23819 (N_23819,N_23454,N_23102);
xnor U23820 (N_23820,N_23054,N_23162);
and U23821 (N_23821,N_23367,N_23480);
or U23822 (N_23822,N_23115,N_23456);
and U23823 (N_23823,N_23156,N_23100);
nor U23824 (N_23824,N_23115,N_23173);
or U23825 (N_23825,N_23260,N_23372);
nand U23826 (N_23826,N_23467,N_23027);
and U23827 (N_23827,N_23336,N_23230);
or U23828 (N_23828,N_23071,N_23447);
or U23829 (N_23829,N_23274,N_23321);
xor U23830 (N_23830,N_23180,N_23379);
nand U23831 (N_23831,N_23374,N_23083);
nand U23832 (N_23832,N_23244,N_23384);
or U23833 (N_23833,N_23436,N_23152);
and U23834 (N_23834,N_23144,N_23436);
xor U23835 (N_23835,N_23014,N_23368);
nand U23836 (N_23836,N_23216,N_23426);
or U23837 (N_23837,N_23468,N_23200);
or U23838 (N_23838,N_23077,N_23175);
and U23839 (N_23839,N_23430,N_23336);
and U23840 (N_23840,N_23164,N_23467);
nand U23841 (N_23841,N_23338,N_23248);
nor U23842 (N_23842,N_23116,N_23076);
or U23843 (N_23843,N_23345,N_23106);
and U23844 (N_23844,N_23170,N_23219);
and U23845 (N_23845,N_23354,N_23144);
and U23846 (N_23846,N_23101,N_23083);
nor U23847 (N_23847,N_23409,N_23141);
xnor U23848 (N_23848,N_23114,N_23455);
or U23849 (N_23849,N_23210,N_23182);
and U23850 (N_23850,N_23016,N_23209);
nand U23851 (N_23851,N_23303,N_23325);
nand U23852 (N_23852,N_23290,N_23170);
and U23853 (N_23853,N_23239,N_23391);
nor U23854 (N_23854,N_23382,N_23147);
nor U23855 (N_23855,N_23432,N_23020);
nor U23856 (N_23856,N_23496,N_23363);
and U23857 (N_23857,N_23036,N_23042);
and U23858 (N_23858,N_23366,N_23480);
nand U23859 (N_23859,N_23453,N_23082);
xor U23860 (N_23860,N_23264,N_23407);
or U23861 (N_23861,N_23490,N_23321);
or U23862 (N_23862,N_23291,N_23106);
and U23863 (N_23863,N_23331,N_23327);
and U23864 (N_23864,N_23085,N_23062);
nor U23865 (N_23865,N_23116,N_23079);
nor U23866 (N_23866,N_23065,N_23102);
and U23867 (N_23867,N_23486,N_23112);
and U23868 (N_23868,N_23264,N_23104);
nand U23869 (N_23869,N_23345,N_23188);
or U23870 (N_23870,N_23162,N_23288);
nor U23871 (N_23871,N_23390,N_23162);
nor U23872 (N_23872,N_23067,N_23351);
or U23873 (N_23873,N_23484,N_23362);
xor U23874 (N_23874,N_23335,N_23117);
or U23875 (N_23875,N_23350,N_23123);
or U23876 (N_23876,N_23210,N_23391);
nor U23877 (N_23877,N_23339,N_23020);
nor U23878 (N_23878,N_23100,N_23464);
xor U23879 (N_23879,N_23327,N_23138);
or U23880 (N_23880,N_23335,N_23364);
or U23881 (N_23881,N_23479,N_23130);
and U23882 (N_23882,N_23481,N_23387);
and U23883 (N_23883,N_23301,N_23084);
and U23884 (N_23884,N_23486,N_23420);
or U23885 (N_23885,N_23475,N_23287);
nor U23886 (N_23886,N_23177,N_23015);
nor U23887 (N_23887,N_23273,N_23359);
or U23888 (N_23888,N_23413,N_23184);
and U23889 (N_23889,N_23236,N_23279);
nor U23890 (N_23890,N_23143,N_23398);
nand U23891 (N_23891,N_23121,N_23268);
nand U23892 (N_23892,N_23299,N_23448);
or U23893 (N_23893,N_23365,N_23306);
xor U23894 (N_23894,N_23407,N_23300);
or U23895 (N_23895,N_23209,N_23420);
or U23896 (N_23896,N_23478,N_23444);
nand U23897 (N_23897,N_23471,N_23470);
and U23898 (N_23898,N_23337,N_23023);
or U23899 (N_23899,N_23389,N_23243);
and U23900 (N_23900,N_23364,N_23387);
or U23901 (N_23901,N_23231,N_23229);
nand U23902 (N_23902,N_23258,N_23123);
or U23903 (N_23903,N_23312,N_23084);
nand U23904 (N_23904,N_23394,N_23267);
nand U23905 (N_23905,N_23159,N_23490);
and U23906 (N_23906,N_23289,N_23225);
and U23907 (N_23907,N_23104,N_23127);
nor U23908 (N_23908,N_23031,N_23471);
or U23909 (N_23909,N_23226,N_23374);
nor U23910 (N_23910,N_23164,N_23234);
nand U23911 (N_23911,N_23242,N_23027);
and U23912 (N_23912,N_23117,N_23258);
nand U23913 (N_23913,N_23161,N_23363);
and U23914 (N_23914,N_23487,N_23074);
or U23915 (N_23915,N_23020,N_23423);
and U23916 (N_23916,N_23439,N_23238);
nand U23917 (N_23917,N_23396,N_23253);
nand U23918 (N_23918,N_23083,N_23205);
or U23919 (N_23919,N_23323,N_23009);
and U23920 (N_23920,N_23243,N_23141);
or U23921 (N_23921,N_23482,N_23211);
or U23922 (N_23922,N_23040,N_23493);
and U23923 (N_23923,N_23453,N_23248);
nand U23924 (N_23924,N_23168,N_23153);
nand U23925 (N_23925,N_23310,N_23158);
nand U23926 (N_23926,N_23304,N_23261);
and U23927 (N_23927,N_23378,N_23181);
or U23928 (N_23928,N_23381,N_23111);
nand U23929 (N_23929,N_23284,N_23386);
or U23930 (N_23930,N_23087,N_23115);
or U23931 (N_23931,N_23036,N_23028);
nor U23932 (N_23932,N_23224,N_23277);
and U23933 (N_23933,N_23282,N_23383);
xor U23934 (N_23934,N_23222,N_23430);
and U23935 (N_23935,N_23141,N_23470);
and U23936 (N_23936,N_23286,N_23385);
nand U23937 (N_23937,N_23363,N_23170);
or U23938 (N_23938,N_23289,N_23424);
and U23939 (N_23939,N_23489,N_23476);
nand U23940 (N_23940,N_23051,N_23002);
and U23941 (N_23941,N_23336,N_23116);
nand U23942 (N_23942,N_23177,N_23289);
nand U23943 (N_23943,N_23132,N_23332);
and U23944 (N_23944,N_23451,N_23108);
nor U23945 (N_23945,N_23043,N_23190);
nor U23946 (N_23946,N_23170,N_23185);
nor U23947 (N_23947,N_23188,N_23421);
xor U23948 (N_23948,N_23322,N_23085);
nor U23949 (N_23949,N_23094,N_23100);
nor U23950 (N_23950,N_23405,N_23300);
or U23951 (N_23951,N_23127,N_23440);
nand U23952 (N_23952,N_23030,N_23325);
and U23953 (N_23953,N_23300,N_23210);
and U23954 (N_23954,N_23168,N_23091);
nor U23955 (N_23955,N_23401,N_23470);
and U23956 (N_23956,N_23378,N_23359);
nand U23957 (N_23957,N_23151,N_23262);
nand U23958 (N_23958,N_23302,N_23067);
and U23959 (N_23959,N_23382,N_23458);
and U23960 (N_23960,N_23492,N_23132);
or U23961 (N_23961,N_23153,N_23440);
xor U23962 (N_23962,N_23373,N_23057);
nor U23963 (N_23963,N_23303,N_23020);
nand U23964 (N_23964,N_23030,N_23261);
xor U23965 (N_23965,N_23416,N_23288);
nand U23966 (N_23966,N_23302,N_23209);
nor U23967 (N_23967,N_23434,N_23250);
and U23968 (N_23968,N_23427,N_23321);
and U23969 (N_23969,N_23383,N_23444);
or U23970 (N_23970,N_23299,N_23437);
or U23971 (N_23971,N_23188,N_23371);
nand U23972 (N_23972,N_23047,N_23216);
nor U23973 (N_23973,N_23253,N_23068);
xnor U23974 (N_23974,N_23198,N_23293);
nor U23975 (N_23975,N_23290,N_23037);
nor U23976 (N_23976,N_23420,N_23083);
or U23977 (N_23977,N_23495,N_23066);
or U23978 (N_23978,N_23450,N_23085);
nor U23979 (N_23979,N_23058,N_23397);
nand U23980 (N_23980,N_23111,N_23144);
and U23981 (N_23981,N_23044,N_23461);
xnor U23982 (N_23982,N_23492,N_23383);
or U23983 (N_23983,N_23188,N_23050);
or U23984 (N_23984,N_23118,N_23053);
nand U23985 (N_23985,N_23485,N_23136);
nor U23986 (N_23986,N_23041,N_23460);
xnor U23987 (N_23987,N_23106,N_23066);
and U23988 (N_23988,N_23246,N_23313);
and U23989 (N_23989,N_23031,N_23069);
and U23990 (N_23990,N_23400,N_23147);
nand U23991 (N_23991,N_23368,N_23406);
or U23992 (N_23992,N_23480,N_23416);
nor U23993 (N_23993,N_23200,N_23365);
nand U23994 (N_23994,N_23362,N_23253);
and U23995 (N_23995,N_23374,N_23389);
xnor U23996 (N_23996,N_23144,N_23255);
or U23997 (N_23997,N_23409,N_23115);
and U23998 (N_23998,N_23307,N_23311);
or U23999 (N_23999,N_23411,N_23127);
and U24000 (N_24000,N_23902,N_23804);
or U24001 (N_24001,N_23581,N_23742);
and U24002 (N_24002,N_23850,N_23767);
nor U24003 (N_24003,N_23699,N_23951);
or U24004 (N_24004,N_23661,N_23664);
nand U24005 (N_24005,N_23504,N_23829);
nand U24006 (N_24006,N_23524,N_23554);
xnor U24007 (N_24007,N_23874,N_23971);
or U24008 (N_24008,N_23795,N_23866);
nor U24009 (N_24009,N_23539,N_23838);
and U24010 (N_24010,N_23522,N_23928);
nor U24011 (N_24011,N_23656,N_23514);
nand U24012 (N_24012,N_23662,N_23657);
or U24013 (N_24013,N_23594,N_23880);
xnor U24014 (N_24014,N_23520,N_23623);
or U24015 (N_24015,N_23527,N_23739);
nand U24016 (N_24016,N_23932,N_23984);
nor U24017 (N_24017,N_23882,N_23989);
or U24018 (N_24018,N_23863,N_23682);
nor U24019 (N_24019,N_23569,N_23813);
or U24020 (N_24020,N_23697,N_23564);
and U24021 (N_24021,N_23553,N_23714);
and U24022 (N_24022,N_23731,N_23884);
nand U24023 (N_24023,N_23784,N_23966);
nor U24024 (N_24024,N_23584,N_23870);
or U24025 (N_24025,N_23678,N_23961);
nor U24026 (N_24026,N_23647,N_23836);
and U24027 (N_24027,N_23865,N_23513);
nor U24028 (N_24028,N_23946,N_23531);
nor U24029 (N_24029,N_23687,N_23552);
xor U24030 (N_24030,N_23737,N_23544);
xnor U24031 (N_24031,N_23671,N_23568);
and U24032 (N_24032,N_23875,N_23782);
and U24033 (N_24033,N_23703,N_23645);
or U24034 (N_24034,N_23810,N_23638);
nand U24035 (N_24035,N_23503,N_23644);
xnor U24036 (N_24036,N_23943,N_23720);
nor U24037 (N_24037,N_23774,N_23941);
nand U24038 (N_24038,N_23740,N_23837);
nand U24039 (N_24039,N_23814,N_23815);
nor U24040 (N_24040,N_23582,N_23597);
or U24041 (N_24041,N_23912,N_23959);
nor U24042 (N_24042,N_23841,N_23999);
nand U24043 (N_24043,N_23631,N_23917);
xor U24044 (N_24044,N_23701,N_23608);
and U24045 (N_24045,N_23652,N_23603);
or U24046 (N_24046,N_23589,N_23995);
nor U24047 (N_24047,N_23980,N_23576);
nand U24048 (N_24048,N_23586,N_23695);
nand U24049 (N_24049,N_23864,N_23974);
nand U24050 (N_24050,N_23952,N_23844);
and U24051 (N_24051,N_23704,N_23533);
nand U24052 (N_24052,N_23909,N_23650);
nor U24053 (N_24053,N_23944,N_23925);
nor U24054 (N_24054,N_23537,N_23525);
nor U24055 (N_24055,N_23511,N_23571);
nor U24056 (N_24056,N_23660,N_23722);
and U24057 (N_24057,N_23688,N_23745);
nand U24058 (N_24058,N_23799,N_23842);
and U24059 (N_24059,N_23879,N_23939);
nor U24060 (N_24060,N_23759,N_23583);
nor U24061 (N_24061,N_23860,N_23857);
nor U24062 (N_24062,N_23518,N_23741);
xor U24063 (N_24063,N_23509,N_23715);
or U24064 (N_24064,N_23764,N_23729);
and U24065 (N_24065,N_23861,N_23903);
nand U24066 (N_24066,N_23901,N_23871);
and U24067 (N_24067,N_23913,N_23904);
nand U24068 (N_24068,N_23962,N_23878);
nor U24069 (N_24069,N_23614,N_23563);
nand U24070 (N_24070,N_23787,N_23725);
xnor U24071 (N_24071,N_23954,N_23821);
xnor U24072 (N_24072,N_23978,N_23790);
or U24073 (N_24073,N_23935,N_23967);
nand U24074 (N_24074,N_23910,N_23775);
and U24075 (N_24075,N_23970,N_23955);
and U24076 (N_24076,N_23834,N_23977);
nor U24077 (N_24077,N_23556,N_23599);
or U24078 (N_24078,N_23685,N_23711);
or U24079 (N_24079,N_23648,N_23762);
and U24080 (N_24080,N_23736,N_23947);
and U24081 (N_24081,N_23519,N_23986);
or U24082 (N_24082,N_23987,N_23748);
nand U24083 (N_24083,N_23642,N_23639);
and U24084 (N_24084,N_23786,N_23777);
nand U24085 (N_24085,N_23624,N_23749);
nand U24086 (N_24086,N_23953,N_23919);
nand U24087 (N_24087,N_23819,N_23532);
and U24088 (N_24088,N_23621,N_23684);
nand U24089 (N_24089,N_23921,N_23881);
or U24090 (N_24090,N_23508,N_23721);
or U24091 (N_24091,N_23789,N_23830);
and U24092 (N_24092,N_23856,N_23942);
nand U24093 (N_24093,N_23964,N_23724);
and U24094 (N_24094,N_23578,N_23773);
and U24095 (N_24095,N_23992,N_23716);
or U24096 (N_24096,N_23801,N_23757);
nand U24097 (N_24097,N_23752,N_23626);
nand U24098 (N_24098,N_23973,N_23765);
nor U24099 (N_24099,N_23700,N_23923);
and U24100 (N_24100,N_23848,N_23558);
or U24101 (N_24101,N_23896,N_23673);
nor U24102 (N_24102,N_23530,N_23976);
and U24103 (N_24103,N_23812,N_23965);
nor U24104 (N_24104,N_23694,N_23632);
nand U24105 (N_24105,N_23605,N_23689);
nand U24106 (N_24106,N_23797,N_23937);
or U24107 (N_24107,N_23933,N_23651);
or U24108 (N_24108,N_23845,N_23523);
nand U24109 (N_24109,N_23924,N_23717);
and U24110 (N_24110,N_23770,N_23990);
xor U24111 (N_24111,N_23920,N_23906);
nor U24112 (N_24112,N_23710,N_23505);
and U24113 (N_24113,N_23570,N_23963);
nor U24114 (N_24114,N_23911,N_23983);
or U24115 (N_24115,N_23824,N_23940);
nor U24116 (N_24116,N_23891,N_23634);
xor U24117 (N_24117,N_23596,N_23677);
nand U24118 (N_24118,N_23876,N_23618);
nor U24119 (N_24119,N_23549,N_23754);
or U24120 (N_24120,N_23674,N_23542);
nor U24121 (N_24121,N_23854,N_23681);
and U24122 (N_24122,N_23610,N_23600);
nand U24123 (N_24123,N_23654,N_23791);
xnor U24124 (N_24124,N_23506,N_23758);
xnor U24125 (N_24125,N_23931,N_23693);
nor U24126 (N_24126,N_23835,N_23653);
nand U24127 (N_24127,N_23692,N_23625);
xnor U24128 (N_24128,N_23772,N_23507);
and U24129 (N_24129,N_23659,N_23550);
and U24130 (N_24130,N_23823,N_23886);
nor U24131 (N_24131,N_23515,N_23580);
and U24132 (N_24132,N_23617,N_23991);
nor U24133 (N_24133,N_23869,N_23817);
or U24134 (N_24134,N_23590,N_23802);
or U24135 (N_24135,N_23769,N_23611);
or U24136 (N_24136,N_23691,N_23756);
and U24137 (N_24137,N_23766,N_23907);
nor U24138 (N_24138,N_23640,N_23683);
and U24139 (N_24139,N_23883,N_23635);
or U24140 (N_24140,N_23573,N_23646);
nand U24141 (N_24141,N_23822,N_23663);
and U24142 (N_24142,N_23619,N_23587);
nor U24143 (N_24143,N_23779,N_23627);
and U24144 (N_24144,N_23750,N_23892);
or U24145 (N_24145,N_23516,N_23858);
nor U24146 (N_24146,N_23852,N_23526);
xnor U24147 (N_24147,N_23807,N_23957);
and U24148 (N_24148,N_23719,N_23781);
nor U24149 (N_24149,N_23825,N_23843);
nor U24150 (N_24150,N_23805,N_23615);
nor U24151 (N_24151,N_23718,N_23649);
nor U24152 (N_24152,N_23686,N_23751);
or U24153 (N_24153,N_23551,N_23606);
xnor U24154 (N_24154,N_23643,N_23969);
or U24155 (N_24155,N_23985,N_23958);
and U24156 (N_24156,N_23847,N_23562);
or U24157 (N_24157,N_23534,N_23760);
xor U24158 (N_24158,N_23602,N_23818);
and U24159 (N_24159,N_23628,N_23894);
nor U24160 (N_24160,N_23755,N_23609);
or U24161 (N_24161,N_23872,N_23922);
nor U24162 (N_24162,N_23898,N_23555);
nor U24163 (N_24163,N_23577,N_23567);
or U24164 (N_24164,N_23560,N_23517);
nand U24165 (N_24165,N_23713,N_23900);
or U24166 (N_24166,N_23670,N_23579);
and U24167 (N_24167,N_23828,N_23612);
or U24168 (N_24168,N_23868,N_23604);
nand U24169 (N_24169,N_23798,N_23712);
nand U24170 (N_24170,N_23595,N_23897);
and U24171 (N_24171,N_23887,N_23601);
and U24172 (N_24172,N_23800,N_23929);
nand U24173 (N_24173,N_23633,N_23778);
nor U24174 (N_24174,N_23690,N_23734);
or U24175 (N_24175,N_23637,N_23588);
nor U24176 (N_24176,N_23949,N_23867);
and U24177 (N_24177,N_23809,N_23655);
nand U24178 (N_24178,N_23794,N_23675);
xnor U24179 (N_24179,N_23761,N_23981);
or U24180 (N_24180,N_23547,N_23806);
nand U24181 (N_24181,N_23780,N_23950);
nand U24182 (N_24182,N_23672,N_23945);
or U24183 (N_24183,N_23808,N_23540);
xor U24184 (N_24184,N_23744,N_23763);
or U24185 (N_24185,N_23667,N_23733);
and U24186 (N_24186,N_23616,N_23747);
and U24187 (N_24187,N_23669,N_23873);
nor U24188 (N_24188,N_23915,N_23908);
xor U24189 (N_24189,N_23575,N_23510);
or U24190 (N_24190,N_23541,N_23783);
nand U24191 (N_24191,N_23998,N_23574);
or U24192 (N_24192,N_23696,N_23811);
and U24193 (N_24193,N_23934,N_23679);
xnor U24194 (N_24194,N_23535,N_23888);
and U24195 (N_24195,N_23926,N_23839);
nor U24196 (N_24196,N_23668,N_23948);
nor U24197 (N_24197,N_23732,N_23592);
nand U24198 (N_24198,N_23796,N_23849);
nand U24199 (N_24199,N_23793,N_23676);
nor U24200 (N_24200,N_23855,N_23738);
nor U24201 (N_24201,N_23585,N_23994);
or U24202 (N_24202,N_23636,N_23607);
nor U24203 (N_24203,N_23622,N_23593);
and U24204 (N_24204,N_23831,N_23538);
nor U24205 (N_24205,N_23996,N_23895);
and U24206 (N_24206,N_23707,N_23833);
or U24207 (N_24207,N_23566,N_23545);
nor U24208 (N_24208,N_23521,N_23561);
and U24209 (N_24209,N_23972,N_23979);
or U24210 (N_24210,N_23768,N_23960);
and U24211 (N_24211,N_23853,N_23666);
nor U24212 (N_24212,N_23746,N_23727);
or U24213 (N_24213,N_23771,N_23877);
nor U24214 (N_24214,N_23753,N_23792);
nand U24215 (N_24215,N_23559,N_23698);
xor U24216 (N_24216,N_23680,N_23529);
and U24217 (N_24217,N_23927,N_23859);
xor U24218 (N_24218,N_23502,N_23816);
nand U24219 (N_24219,N_23899,N_23776);
nand U24220 (N_24220,N_23893,N_23889);
nor U24221 (N_24221,N_23705,N_23613);
nor U24222 (N_24222,N_23916,N_23820);
xnor U24223 (N_24223,N_23930,N_23572);
xnor U24224 (N_24224,N_23862,N_23846);
and U24225 (N_24225,N_23629,N_23730);
or U24226 (N_24226,N_23620,N_23803);
nor U24227 (N_24227,N_23543,N_23956);
or U24228 (N_24228,N_23827,N_23598);
and U24229 (N_24229,N_23936,N_23840);
nor U24230 (N_24230,N_23665,N_23702);
and U24231 (N_24231,N_23826,N_23591);
and U24232 (N_24232,N_23726,N_23630);
and U24233 (N_24233,N_23988,N_23728);
nor U24234 (N_24234,N_23832,N_23743);
and U24235 (N_24235,N_23918,N_23658);
nand U24236 (N_24236,N_23708,N_23641);
and U24237 (N_24237,N_23851,N_23528);
nor U24238 (N_24238,N_23706,N_23536);
or U24239 (N_24239,N_23723,N_23500);
xor U24240 (N_24240,N_23997,N_23548);
and U24241 (N_24241,N_23546,N_23788);
xor U24242 (N_24242,N_23785,N_23557);
nand U24243 (N_24243,N_23709,N_23501);
and U24244 (N_24244,N_23565,N_23982);
or U24245 (N_24245,N_23890,N_23968);
nand U24246 (N_24246,N_23993,N_23735);
nand U24247 (N_24247,N_23938,N_23914);
and U24248 (N_24248,N_23512,N_23885);
or U24249 (N_24249,N_23975,N_23905);
or U24250 (N_24250,N_23601,N_23906);
nand U24251 (N_24251,N_23720,N_23547);
or U24252 (N_24252,N_23780,N_23674);
and U24253 (N_24253,N_23601,N_23511);
nand U24254 (N_24254,N_23772,N_23902);
xor U24255 (N_24255,N_23957,N_23849);
or U24256 (N_24256,N_23973,N_23897);
nand U24257 (N_24257,N_23747,N_23513);
and U24258 (N_24258,N_23879,N_23669);
and U24259 (N_24259,N_23910,N_23526);
or U24260 (N_24260,N_23599,N_23995);
nor U24261 (N_24261,N_23638,N_23859);
and U24262 (N_24262,N_23553,N_23878);
and U24263 (N_24263,N_23805,N_23929);
nand U24264 (N_24264,N_23732,N_23555);
or U24265 (N_24265,N_23610,N_23719);
nor U24266 (N_24266,N_23998,N_23573);
nand U24267 (N_24267,N_23814,N_23921);
nand U24268 (N_24268,N_23588,N_23785);
nand U24269 (N_24269,N_23841,N_23765);
xor U24270 (N_24270,N_23871,N_23857);
nor U24271 (N_24271,N_23917,N_23613);
and U24272 (N_24272,N_23766,N_23687);
and U24273 (N_24273,N_23840,N_23549);
and U24274 (N_24274,N_23913,N_23694);
xnor U24275 (N_24275,N_23567,N_23755);
and U24276 (N_24276,N_23951,N_23684);
or U24277 (N_24277,N_23804,N_23859);
nor U24278 (N_24278,N_23782,N_23526);
xor U24279 (N_24279,N_23750,N_23742);
nand U24280 (N_24280,N_23546,N_23961);
and U24281 (N_24281,N_23638,N_23782);
and U24282 (N_24282,N_23697,N_23691);
nor U24283 (N_24283,N_23621,N_23971);
or U24284 (N_24284,N_23537,N_23607);
and U24285 (N_24285,N_23861,N_23538);
and U24286 (N_24286,N_23889,N_23977);
xnor U24287 (N_24287,N_23563,N_23893);
nand U24288 (N_24288,N_23952,N_23552);
and U24289 (N_24289,N_23804,N_23724);
nor U24290 (N_24290,N_23723,N_23941);
nand U24291 (N_24291,N_23765,N_23678);
nand U24292 (N_24292,N_23696,N_23649);
nand U24293 (N_24293,N_23818,N_23712);
nand U24294 (N_24294,N_23809,N_23994);
or U24295 (N_24295,N_23983,N_23652);
or U24296 (N_24296,N_23756,N_23541);
xor U24297 (N_24297,N_23665,N_23853);
or U24298 (N_24298,N_23763,N_23526);
nand U24299 (N_24299,N_23746,N_23965);
nor U24300 (N_24300,N_23787,N_23697);
or U24301 (N_24301,N_23580,N_23915);
nor U24302 (N_24302,N_23813,N_23585);
nor U24303 (N_24303,N_23812,N_23568);
and U24304 (N_24304,N_23724,N_23857);
nand U24305 (N_24305,N_23657,N_23766);
or U24306 (N_24306,N_23944,N_23517);
nor U24307 (N_24307,N_23670,N_23701);
nand U24308 (N_24308,N_23649,N_23805);
nand U24309 (N_24309,N_23853,N_23563);
or U24310 (N_24310,N_23685,N_23939);
nor U24311 (N_24311,N_23749,N_23977);
xnor U24312 (N_24312,N_23607,N_23811);
or U24313 (N_24313,N_23649,N_23777);
nor U24314 (N_24314,N_23886,N_23702);
nor U24315 (N_24315,N_23611,N_23554);
nor U24316 (N_24316,N_23760,N_23835);
and U24317 (N_24317,N_23530,N_23585);
nand U24318 (N_24318,N_23707,N_23914);
nor U24319 (N_24319,N_23538,N_23855);
xnor U24320 (N_24320,N_23616,N_23588);
or U24321 (N_24321,N_23788,N_23967);
and U24322 (N_24322,N_23949,N_23776);
nor U24323 (N_24323,N_23910,N_23875);
nor U24324 (N_24324,N_23556,N_23916);
nor U24325 (N_24325,N_23634,N_23508);
nand U24326 (N_24326,N_23894,N_23913);
nand U24327 (N_24327,N_23727,N_23575);
nand U24328 (N_24328,N_23807,N_23529);
and U24329 (N_24329,N_23544,N_23961);
or U24330 (N_24330,N_23785,N_23952);
xor U24331 (N_24331,N_23677,N_23907);
or U24332 (N_24332,N_23707,N_23743);
nor U24333 (N_24333,N_23597,N_23855);
or U24334 (N_24334,N_23540,N_23814);
nor U24335 (N_24335,N_23655,N_23791);
xnor U24336 (N_24336,N_23913,N_23753);
or U24337 (N_24337,N_23516,N_23649);
nor U24338 (N_24338,N_23796,N_23918);
nand U24339 (N_24339,N_23722,N_23717);
nand U24340 (N_24340,N_23992,N_23738);
or U24341 (N_24341,N_23771,N_23690);
and U24342 (N_24342,N_23594,N_23948);
xor U24343 (N_24343,N_23946,N_23737);
and U24344 (N_24344,N_23720,N_23682);
and U24345 (N_24345,N_23541,N_23820);
nor U24346 (N_24346,N_23879,N_23712);
and U24347 (N_24347,N_23682,N_23512);
xnor U24348 (N_24348,N_23526,N_23593);
nand U24349 (N_24349,N_23747,N_23986);
xnor U24350 (N_24350,N_23563,N_23551);
and U24351 (N_24351,N_23773,N_23709);
nor U24352 (N_24352,N_23536,N_23712);
nor U24353 (N_24353,N_23725,N_23576);
and U24354 (N_24354,N_23988,N_23725);
nor U24355 (N_24355,N_23865,N_23612);
nor U24356 (N_24356,N_23875,N_23851);
and U24357 (N_24357,N_23705,N_23982);
and U24358 (N_24358,N_23698,N_23750);
xnor U24359 (N_24359,N_23690,N_23938);
xor U24360 (N_24360,N_23516,N_23737);
or U24361 (N_24361,N_23642,N_23567);
nand U24362 (N_24362,N_23714,N_23796);
and U24363 (N_24363,N_23839,N_23641);
nor U24364 (N_24364,N_23952,N_23910);
nor U24365 (N_24365,N_23927,N_23909);
nor U24366 (N_24366,N_23864,N_23734);
nand U24367 (N_24367,N_23998,N_23794);
xor U24368 (N_24368,N_23889,N_23978);
and U24369 (N_24369,N_23854,N_23604);
or U24370 (N_24370,N_23897,N_23917);
or U24371 (N_24371,N_23903,N_23737);
or U24372 (N_24372,N_23627,N_23585);
or U24373 (N_24373,N_23994,N_23695);
nor U24374 (N_24374,N_23696,N_23636);
nand U24375 (N_24375,N_23892,N_23984);
nand U24376 (N_24376,N_23842,N_23780);
or U24377 (N_24377,N_23552,N_23801);
nor U24378 (N_24378,N_23891,N_23598);
nand U24379 (N_24379,N_23832,N_23749);
or U24380 (N_24380,N_23696,N_23592);
and U24381 (N_24381,N_23948,N_23822);
or U24382 (N_24382,N_23579,N_23519);
nand U24383 (N_24383,N_23526,N_23860);
or U24384 (N_24384,N_23952,N_23519);
nand U24385 (N_24385,N_23671,N_23757);
nor U24386 (N_24386,N_23647,N_23921);
nand U24387 (N_24387,N_23526,N_23877);
xnor U24388 (N_24388,N_23556,N_23550);
nor U24389 (N_24389,N_23890,N_23957);
and U24390 (N_24390,N_23957,N_23993);
xnor U24391 (N_24391,N_23762,N_23692);
or U24392 (N_24392,N_23548,N_23909);
and U24393 (N_24393,N_23858,N_23740);
nor U24394 (N_24394,N_23640,N_23539);
nor U24395 (N_24395,N_23754,N_23767);
or U24396 (N_24396,N_23864,N_23892);
and U24397 (N_24397,N_23564,N_23929);
nor U24398 (N_24398,N_23924,N_23919);
or U24399 (N_24399,N_23955,N_23578);
nand U24400 (N_24400,N_23573,N_23614);
nand U24401 (N_24401,N_23696,N_23921);
and U24402 (N_24402,N_23616,N_23822);
and U24403 (N_24403,N_23551,N_23815);
nand U24404 (N_24404,N_23682,N_23916);
nor U24405 (N_24405,N_23834,N_23842);
or U24406 (N_24406,N_23752,N_23513);
nor U24407 (N_24407,N_23848,N_23863);
and U24408 (N_24408,N_23706,N_23739);
and U24409 (N_24409,N_23529,N_23576);
nand U24410 (N_24410,N_23720,N_23635);
or U24411 (N_24411,N_23608,N_23739);
xor U24412 (N_24412,N_23821,N_23610);
xnor U24413 (N_24413,N_23997,N_23670);
nor U24414 (N_24414,N_23960,N_23851);
and U24415 (N_24415,N_23764,N_23601);
nor U24416 (N_24416,N_23783,N_23851);
nand U24417 (N_24417,N_23959,N_23754);
and U24418 (N_24418,N_23845,N_23935);
nand U24419 (N_24419,N_23771,N_23976);
and U24420 (N_24420,N_23970,N_23753);
or U24421 (N_24421,N_23889,N_23742);
and U24422 (N_24422,N_23720,N_23751);
nand U24423 (N_24423,N_23737,N_23846);
nand U24424 (N_24424,N_23724,N_23819);
nand U24425 (N_24425,N_23628,N_23735);
nor U24426 (N_24426,N_23596,N_23779);
or U24427 (N_24427,N_23656,N_23641);
xnor U24428 (N_24428,N_23769,N_23738);
nor U24429 (N_24429,N_23836,N_23547);
or U24430 (N_24430,N_23505,N_23567);
xnor U24431 (N_24431,N_23561,N_23958);
nand U24432 (N_24432,N_23976,N_23770);
or U24433 (N_24433,N_23730,N_23850);
or U24434 (N_24434,N_23582,N_23776);
and U24435 (N_24435,N_23880,N_23631);
nand U24436 (N_24436,N_23805,N_23638);
or U24437 (N_24437,N_23798,N_23699);
and U24438 (N_24438,N_23702,N_23562);
xnor U24439 (N_24439,N_23820,N_23774);
nor U24440 (N_24440,N_23767,N_23683);
xnor U24441 (N_24441,N_23787,N_23669);
xnor U24442 (N_24442,N_23784,N_23618);
xnor U24443 (N_24443,N_23538,N_23824);
and U24444 (N_24444,N_23805,N_23717);
or U24445 (N_24445,N_23974,N_23698);
or U24446 (N_24446,N_23614,N_23651);
nor U24447 (N_24447,N_23821,N_23797);
nor U24448 (N_24448,N_23823,N_23689);
or U24449 (N_24449,N_23897,N_23960);
nor U24450 (N_24450,N_23934,N_23513);
nor U24451 (N_24451,N_23624,N_23540);
or U24452 (N_24452,N_23955,N_23527);
or U24453 (N_24453,N_23647,N_23742);
nand U24454 (N_24454,N_23819,N_23677);
and U24455 (N_24455,N_23992,N_23828);
and U24456 (N_24456,N_23938,N_23751);
nand U24457 (N_24457,N_23959,N_23634);
nor U24458 (N_24458,N_23958,N_23963);
or U24459 (N_24459,N_23587,N_23868);
nor U24460 (N_24460,N_23641,N_23861);
nor U24461 (N_24461,N_23625,N_23617);
and U24462 (N_24462,N_23574,N_23891);
or U24463 (N_24463,N_23821,N_23921);
nor U24464 (N_24464,N_23756,N_23552);
nor U24465 (N_24465,N_23527,N_23622);
or U24466 (N_24466,N_23879,N_23882);
nand U24467 (N_24467,N_23620,N_23828);
nor U24468 (N_24468,N_23971,N_23605);
or U24469 (N_24469,N_23727,N_23878);
xor U24470 (N_24470,N_23719,N_23744);
xor U24471 (N_24471,N_23881,N_23578);
and U24472 (N_24472,N_23962,N_23886);
nor U24473 (N_24473,N_23844,N_23967);
or U24474 (N_24474,N_23811,N_23972);
nand U24475 (N_24475,N_23597,N_23594);
or U24476 (N_24476,N_23944,N_23661);
or U24477 (N_24477,N_23691,N_23695);
or U24478 (N_24478,N_23941,N_23642);
nand U24479 (N_24479,N_23718,N_23870);
nor U24480 (N_24480,N_23979,N_23627);
nor U24481 (N_24481,N_23836,N_23820);
nand U24482 (N_24482,N_23861,N_23964);
or U24483 (N_24483,N_23687,N_23661);
nand U24484 (N_24484,N_23511,N_23907);
and U24485 (N_24485,N_23508,N_23901);
nor U24486 (N_24486,N_23735,N_23615);
and U24487 (N_24487,N_23975,N_23588);
or U24488 (N_24488,N_23968,N_23714);
nand U24489 (N_24489,N_23784,N_23798);
nor U24490 (N_24490,N_23933,N_23902);
nor U24491 (N_24491,N_23701,N_23530);
and U24492 (N_24492,N_23643,N_23918);
or U24493 (N_24493,N_23850,N_23808);
xnor U24494 (N_24494,N_23780,N_23727);
nor U24495 (N_24495,N_23537,N_23727);
and U24496 (N_24496,N_23822,N_23937);
or U24497 (N_24497,N_23768,N_23979);
and U24498 (N_24498,N_23744,N_23884);
nand U24499 (N_24499,N_23890,N_23973);
or U24500 (N_24500,N_24481,N_24414);
nor U24501 (N_24501,N_24111,N_24030);
and U24502 (N_24502,N_24265,N_24338);
or U24503 (N_24503,N_24378,N_24350);
and U24504 (N_24504,N_24104,N_24389);
and U24505 (N_24505,N_24305,N_24297);
nor U24506 (N_24506,N_24263,N_24404);
and U24507 (N_24507,N_24408,N_24363);
xor U24508 (N_24508,N_24114,N_24425);
nor U24509 (N_24509,N_24276,N_24105);
nand U24510 (N_24510,N_24452,N_24087);
or U24511 (N_24511,N_24032,N_24061);
xnor U24512 (N_24512,N_24216,N_24482);
or U24513 (N_24513,N_24225,N_24280);
nand U24514 (N_24514,N_24018,N_24068);
nor U24515 (N_24515,N_24262,N_24247);
xor U24516 (N_24516,N_24093,N_24128);
or U24517 (N_24517,N_24116,N_24142);
or U24518 (N_24518,N_24147,N_24108);
and U24519 (N_24519,N_24190,N_24264);
nand U24520 (N_24520,N_24110,N_24460);
and U24521 (N_24521,N_24480,N_24468);
nand U24522 (N_24522,N_24293,N_24085);
and U24523 (N_24523,N_24437,N_24491);
nand U24524 (N_24524,N_24083,N_24155);
nand U24525 (N_24525,N_24149,N_24398);
or U24526 (N_24526,N_24181,N_24209);
nand U24527 (N_24527,N_24457,N_24047);
nand U24528 (N_24528,N_24086,N_24029);
and U24529 (N_24529,N_24072,N_24230);
nand U24530 (N_24530,N_24318,N_24429);
and U24531 (N_24531,N_24150,N_24129);
or U24532 (N_24532,N_24192,N_24436);
or U24533 (N_24533,N_24417,N_24455);
or U24534 (N_24534,N_24485,N_24394);
and U24535 (N_24535,N_24075,N_24431);
nor U24536 (N_24536,N_24490,N_24214);
and U24537 (N_24537,N_24148,N_24364);
xor U24538 (N_24538,N_24203,N_24245);
and U24539 (N_24539,N_24345,N_24058);
xnor U24540 (N_24540,N_24182,N_24407);
nand U24541 (N_24541,N_24416,N_24141);
nand U24542 (N_24542,N_24271,N_24441);
and U24543 (N_24543,N_24351,N_24326);
nor U24544 (N_24544,N_24220,N_24419);
or U24545 (N_24545,N_24342,N_24115);
xor U24546 (N_24546,N_24295,N_24454);
or U24547 (N_24547,N_24258,N_24023);
nor U24548 (N_24548,N_24473,N_24495);
nor U24549 (N_24549,N_24161,N_24004);
and U24550 (N_24550,N_24002,N_24470);
nand U24551 (N_24551,N_24212,N_24231);
and U24552 (N_24552,N_24423,N_24427);
and U24553 (N_24553,N_24021,N_24330);
nand U24554 (N_24554,N_24445,N_24022);
or U24555 (N_24555,N_24073,N_24173);
and U24556 (N_24556,N_24303,N_24366);
nand U24557 (N_24557,N_24362,N_24084);
or U24558 (N_24558,N_24145,N_24443);
nand U24559 (N_24559,N_24402,N_24463);
nand U24560 (N_24560,N_24444,N_24179);
nand U24561 (N_24561,N_24151,N_24406);
and U24562 (N_24562,N_24467,N_24356);
or U24563 (N_24563,N_24067,N_24180);
and U24564 (N_24564,N_24273,N_24392);
nor U24565 (N_24565,N_24285,N_24076);
or U24566 (N_24566,N_24438,N_24156);
and U24567 (N_24567,N_24449,N_24240);
nor U24568 (N_24568,N_24349,N_24287);
xnor U24569 (N_24569,N_24167,N_24456);
and U24570 (N_24570,N_24183,N_24331);
nor U24571 (N_24571,N_24393,N_24368);
xnor U24572 (N_24572,N_24301,N_24215);
nor U24573 (N_24573,N_24064,N_24211);
or U24574 (N_24574,N_24348,N_24282);
nor U24575 (N_24575,N_24132,N_24334);
and U24576 (N_24576,N_24246,N_24388);
xnor U24577 (N_24577,N_24405,N_24250);
nand U24578 (N_24578,N_24477,N_24113);
and U24579 (N_24579,N_24045,N_24090);
nand U24580 (N_24580,N_24284,N_24178);
nand U24581 (N_24581,N_24252,N_24077);
and U24582 (N_24582,N_24380,N_24381);
and U24583 (N_24583,N_24383,N_24377);
nand U24584 (N_24584,N_24496,N_24433);
nand U24585 (N_24585,N_24099,N_24315);
nand U24586 (N_24586,N_24081,N_24379);
and U24587 (N_24587,N_24261,N_24060);
nand U24588 (N_24588,N_24476,N_24223);
or U24589 (N_24589,N_24484,N_24307);
and U24590 (N_24590,N_24277,N_24109);
nor U24591 (N_24591,N_24100,N_24268);
nor U24592 (N_24592,N_24397,N_24292);
nor U24593 (N_24593,N_24453,N_24006);
xnor U24594 (N_24594,N_24234,N_24213);
nor U24595 (N_24595,N_24340,N_24298);
and U24596 (N_24596,N_24043,N_24079);
nand U24597 (N_24597,N_24497,N_24469);
xor U24598 (N_24598,N_24207,N_24387);
nand U24599 (N_24599,N_24311,N_24396);
nor U24600 (N_24600,N_24126,N_24369);
nor U24601 (N_24601,N_24028,N_24321);
nand U24602 (N_24602,N_24176,N_24420);
and U24603 (N_24603,N_24472,N_24102);
and U24604 (N_24604,N_24286,N_24010);
or U24605 (N_24605,N_24044,N_24434);
and U24606 (N_24606,N_24097,N_24353);
nor U24607 (N_24607,N_24488,N_24165);
nand U24608 (N_24608,N_24034,N_24143);
nand U24609 (N_24609,N_24154,N_24229);
or U24610 (N_24610,N_24187,N_24144);
and U24611 (N_24611,N_24251,N_24185);
nand U24612 (N_24612,N_24164,N_24300);
nor U24613 (N_24613,N_24347,N_24124);
xor U24614 (N_24614,N_24269,N_24189);
nor U24615 (N_24615,N_24162,N_24020);
and U24616 (N_24616,N_24281,N_24121);
and U24617 (N_24617,N_24123,N_24442);
nor U24618 (N_24618,N_24399,N_24304);
nor U24619 (N_24619,N_24339,N_24236);
or U24620 (N_24620,N_24249,N_24319);
nand U24621 (N_24621,N_24136,N_24198);
or U24622 (N_24622,N_24107,N_24248);
nor U24623 (N_24623,N_24447,N_24219);
nand U24624 (N_24624,N_24367,N_24375);
nand U24625 (N_24625,N_24233,N_24462);
and U24626 (N_24626,N_24283,N_24217);
and U24627 (N_24627,N_24157,N_24446);
nand U24628 (N_24628,N_24257,N_24094);
or U24629 (N_24629,N_24475,N_24486);
nand U24630 (N_24630,N_24421,N_24008);
nand U24631 (N_24631,N_24101,N_24054);
nor U24632 (N_24632,N_24140,N_24323);
nor U24633 (N_24633,N_24127,N_24357);
xor U24634 (N_24634,N_24479,N_24494);
nand U24635 (N_24635,N_24493,N_24222);
or U24636 (N_24636,N_24201,N_24137);
or U24637 (N_24637,N_24478,N_24066);
nor U24638 (N_24638,N_24074,N_24133);
nor U24639 (N_24639,N_24166,N_24053);
xnor U24640 (N_24640,N_24131,N_24314);
and U24641 (N_24641,N_24422,N_24412);
nand U24642 (N_24642,N_24027,N_24499);
or U24643 (N_24643,N_24009,N_24130);
nand U24644 (N_24644,N_24242,N_24270);
and U24645 (N_24645,N_24355,N_24371);
and U24646 (N_24646,N_24385,N_24036);
nand U24647 (N_24647,N_24051,N_24255);
and U24648 (N_24648,N_24193,N_24430);
nand U24649 (N_24649,N_24401,N_24428);
nor U24650 (N_24650,N_24317,N_24274);
nor U24651 (N_24651,N_24195,N_24384);
nor U24652 (N_24652,N_24333,N_24070);
or U24653 (N_24653,N_24341,N_24033);
nor U24654 (N_24654,N_24324,N_24310);
nand U24655 (N_24655,N_24120,N_24095);
nor U24656 (N_24656,N_24171,N_24418);
nor U24657 (N_24657,N_24177,N_24376);
nand U24658 (N_24658,N_24065,N_24117);
nor U24659 (N_24659,N_24259,N_24011);
nor U24660 (N_24660,N_24243,N_24218);
or U24661 (N_24661,N_24374,N_24163);
and U24662 (N_24662,N_24118,N_24146);
nand U24663 (N_24663,N_24253,N_24175);
and U24664 (N_24664,N_24237,N_24200);
xor U24665 (N_24665,N_24343,N_24103);
and U24666 (N_24666,N_24168,N_24410);
nand U24667 (N_24667,N_24400,N_24096);
nand U24668 (N_24668,N_24135,N_24386);
and U24669 (N_24669,N_24019,N_24139);
nand U24670 (N_24670,N_24160,N_24206);
and U24671 (N_24671,N_24365,N_24360);
nor U24672 (N_24672,N_24199,N_24332);
nor U24673 (N_24673,N_24153,N_24451);
and U24674 (N_24674,N_24188,N_24025);
nand U24675 (N_24675,N_24288,N_24091);
nand U24676 (N_24676,N_24046,N_24174);
or U24677 (N_24677,N_24291,N_24403);
nor U24678 (N_24678,N_24221,N_24228);
or U24679 (N_24679,N_24001,N_24224);
xor U24680 (N_24680,N_24336,N_24138);
and U24681 (N_24681,N_24050,N_24159);
or U24682 (N_24682,N_24191,N_24026);
or U24683 (N_24683,N_24069,N_24391);
nor U24684 (N_24684,N_24239,N_24395);
nor U24685 (N_24685,N_24306,N_24017);
and U24686 (N_24686,N_24092,N_24413);
or U24687 (N_24687,N_24309,N_24372);
nand U24688 (N_24688,N_24487,N_24275);
or U24689 (N_24689,N_24122,N_24040);
and U24690 (N_24690,N_24158,N_24256);
nand U24691 (N_24691,N_24489,N_24279);
and U24692 (N_24692,N_24059,N_24299);
and U24693 (N_24693,N_24204,N_24238);
nand U24694 (N_24694,N_24267,N_24232);
or U24695 (N_24695,N_24459,N_24056);
nand U24696 (N_24696,N_24170,N_24448);
nor U24697 (N_24697,N_24012,N_24450);
or U24698 (N_24698,N_24254,N_24031);
nand U24699 (N_24699,N_24226,N_24062);
nor U24700 (N_24700,N_24049,N_24202);
nand U24701 (N_24701,N_24435,N_24244);
and U24702 (N_24702,N_24227,N_24409);
nand U24703 (N_24703,N_24474,N_24057);
or U24704 (N_24704,N_24000,N_24492);
nand U24705 (N_24705,N_24346,N_24312);
or U24706 (N_24706,N_24039,N_24098);
nand U24707 (N_24707,N_24080,N_24194);
and U24708 (N_24708,N_24272,N_24007);
nand U24709 (N_24709,N_24052,N_24320);
or U24710 (N_24710,N_24037,N_24370);
or U24711 (N_24711,N_24390,N_24210);
nand U24712 (N_24712,N_24329,N_24205);
nor U24713 (N_24713,N_24041,N_24328);
and U24714 (N_24714,N_24461,N_24483);
nand U24715 (N_24715,N_24289,N_24241);
nand U24716 (N_24716,N_24260,N_24082);
nand U24717 (N_24717,N_24294,N_24184);
xnor U24718 (N_24718,N_24382,N_24440);
and U24719 (N_24719,N_24325,N_24302);
and U24720 (N_24720,N_24005,N_24042);
nor U24721 (N_24721,N_24266,N_24125);
nor U24722 (N_24722,N_24055,N_24327);
or U24723 (N_24723,N_24361,N_24411);
and U24724 (N_24724,N_24458,N_24119);
and U24725 (N_24725,N_24152,N_24063);
and U24726 (N_24726,N_24464,N_24038);
or U24727 (N_24727,N_24186,N_24296);
nand U24728 (N_24728,N_24112,N_24071);
nor U24729 (N_24729,N_24235,N_24354);
nand U24730 (N_24730,N_24089,N_24290);
or U24731 (N_24731,N_24322,N_24426);
and U24732 (N_24732,N_24003,N_24439);
and U24733 (N_24733,N_24498,N_24415);
nor U24734 (N_24734,N_24352,N_24308);
and U24735 (N_24735,N_24172,N_24466);
or U24736 (N_24736,N_24035,N_24373);
and U24737 (N_24737,N_24337,N_24358);
and U24738 (N_24738,N_24335,N_24278);
nor U24739 (N_24739,N_24344,N_24134);
nand U24740 (N_24740,N_24359,N_24197);
nand U24741 (N_24741,N_24313,N_24024);
and U24742 (N_24742,N_24078,N_24013);
and U24743 (N_24743,N_24316,N_24106);
or U24744 (N_24744,N_24465,N_24014);
and U24745 (N_24745,N_24196,N_24169);
nor U24746 (N_24746,N_24016,N_24432);
nor U24747 (N_24747,N_24424,N_24471);
nor U24748 (N_24748,N_24048,N_24015);
nor U24749 (N_24749,N_24088,N_24208);
and U24750 (N_24750,N_24090,N_24111);
or U24751 (N_24751,N_24067,N_24167);
nor U24752 (N_24752,N_24330,N_24383);
nor U24753 (N_24753,N_24333,N_24463);
nor U24754 (N_24754,N_24302,N_24238);
and U24755 (N_24755,N_24022,N_24161);
and U24756 (N_24756,N_24145,N_24442);
nor U24757 (N_24757,N_24009,N_24270);
or U24758 (N_24758,N_24159,N_24217);
nor U24759 (N_24759,N_24443,N_24483);
and U24760 (N_24760,N_24095,N_24398);
nor U24761 (N_24761,N_24295,N_24455);
nand U24762 (N_24762,N_24057,N_24028);
nand U24763 (N_24763,N_24264,N_24472);
nand U24764 (N_24764,N_24236,N_24031);
or U24765 (N_24765,N_24281,N_24111);
xor U24766 (N_24766,N_24469,N_24376);
nand U24767 (N_24767,N_24348,N_24395);
nand U24768 (N_24768,N_24010,N_24081);
nand U24769 (N_24769,N_24080,N_24004);
nor U24770 (N_24770,N_24020,N_24038);
nor U24771 (N_24771,N_24413,N_24075);
xor U24772 (N_24772,N_24151,N_24199);
and U24773 (N_24773,N_24370,N_24089);
and U24774 (N_24774,N_24272,N_24338);
and U24775 (N_24775,N_24453,N_24034);
nor U24776 (N_24776,N_24378,N_24472);
or U24777 (N_24777,N_24356,N_24292);
or U24778 (N_24778,N_24364,N_24169);
xor U24779 (N_24779,N_24420,N_24173);
nor U24780 (N_24780,N_24180,N_24338);
nand U24781 (N_24781,N_24335,N_24410);
nand U24782 (N_24782,N_24388,N_24068);
nand U24783 (N_24783,N_24352,N_24211);
nand U24784 (N_24784,N_24421,N_24155);
nand U24785 (N_24785,N_24342,N_24481);
or U24786 (N_24786,N_24219,N_24145);
xnor U24787 (N_24787,N_24446,N_24074);
and U24788 (N_24788,N_24060,N_24097);
nand U24789 (N_24789,N_24233,N_24043);
and U24790 (N_24790,N_24021,N_24196);
nor U24791 (N_24791,N_24342,N_24405);
nor U24792 (N_24792,N_24004,N_24233);
or U24793 (N_24793,N_24097,N_24177);
nand U24794 (N_24794,N_24326,N_24260);
nand U24795 (N_24795,N_24141,N_24252);
or U24796 (N_24796,N_24263,N_24308);
or U24797 (N_24797,N_24092,N_24398);
and U24798 (N_24798,N_24255,N_24371);
nand U24799 (N_24799,N_24029,N_24072);
and U24800 (N_24800,N_24401,N_24416);
xnor U24801 (N_24801,N_24360,N_24190);
nand U24802 (N_24802,N_24105,N_24399);
nor U24803 (N_24803,N_24250,N_24158);
or U24804 (N_24804,N_24320,N_24110);
nor U24805 (N_24805,N_24261,N_24199);
nand U24806 (N_24806,N_24225,N_24387);
and U24807 (N_24807,N_24446,N_24327);
nand U24808 (N_24808,N_24168,N_24154);
nor U24809 (N_24809,N_24136,N_24142);
nor U24810 (N_24810,N_24484,N_24040);
nor U24811 (N_24811,N_24170,N_24359);
nand U24812 (N_24812,N_24320,N_24183);
nor U24813 (N_24813,N_24118,N_24171);
xor U24814 (N_24814,N_24333,N_24106);
or U24815 (N_24815,N_24384,N_24393);
and U24816 (N_24816,N_24121,N_24469);
or U24817 (N_24817,N_24480,N_24181);
xnor U24818 (N_24818,N_24081,N_24216);
and U24819 (N_24819,N_24424,N_24480);
nor U24820 (N_24820,N_24334,N_24217);
or U24821 (N_24821,N_24304,N_24065);
nand U24822 (N_24822,N_24213,N_24399);
or U24823 (N_24823,N_24243,N_24375);
nand U24824 (N_24824,N_24125,N_24388);
and U24825 (N_24825,N_24258,N_24425);
nand U24826 (N_24826,N_24092,N_24098);
nand U24827 (N_24827,N_24115,N_24465);
nand U24828 (N_24828,N_24163,N_24335);
nand U24829 (N_24829,N_24457,N_24462);
nand U24830 (N_24830,N_24087,N_24193);
xor U24831 (N_24831,N_24398,N_24417);
or U24832 (N_24832,N_24044,N_24332);
nand U24833 (N_24833,N_24160,N_24446);
and U24834 (N_24834,N_24426,N_24323);
and U24835 (N_24835,N_24139,N_24307);
nand U24836 (N_24836,N_24326,N_24015);
nor U24837 (N_24837,N_24379,N_24012);
or U24838 (N_24838,N_24191,N_24301);
or U24839 (N_24839,N_24234,N_24172);
nand U24840 (N_24840,N_24328,N_24318);
and U24841 (N_24841,N_24003,N_24032);
nor U24842 (N_24842,N_24174,N_24446);
and U24843 (N_24843,N_24186,N_24012);
or U24844 (N_24844,N_24405,N_24404);
nand U24845 (N_24845,N_24060,N_24083);
xnor U24846 (N_24846,N_24047,N_24055);
xnor U24847 (N_24847,N_24274,N_24051);
xor U24848 (N_24848,N_24347,N_24451);
or U24849 (N_24849,N_24453,N_24215);
and U24850 (N_24850,N_24039,N_24457);
or U24851 (N_24851,N_24144,N_24116);
or U24852 (N_24852,N_24452,N_24022);
nand U24853 (N_24853,N_24096,N_24165);
nand U24854 (N_24854,N_24072,N_24336);
nand U24855 (N_24855,N_24117,N_24002);
or U24856 (N_24856,N_24185,N_24018);
nand U24857 (N_24857,N_24139,N_24100);
and U24858 (N_24858,N_24337,N_24414);
and U24859 (N_24859,N_24358,N_24022);
nor U24860 (N_24860,N_24154,N_24416);
or U24861 (N_24861,N_24453,N_24240);
or U24862 (N_24862,N_24453,N_24463);
or U24863 (N_24863,N_24050,N_24270);
or U24864 (N_24864,N_24325,N_24126);
or U24865 (N_24865,N_24495,N_24046);
nor U24866 (N_24866,N_24318,N_24329);
nor U24867 (N_24867,N_24095,N_24027);
nand U24868 (N_24868,N_24487,N_24117);
nand U24869 (N_24869,N_24473,N_24272);
nor U24870 (N_24870,N_24270,N_24462);
nand U24871 (N_24871,N_24287,N_24493);
nor U24872 (N_24872,N_24223,N_24047);
nor U24873 (N_24873,N_24244,N_24407);
nand U24874 (N_24874,N_24353,N_24283);
or U24875 (N_24875,N_24083,N_24402);
or U24876 (N_24876,N_24441,N_24015);
nor U24877 (N_24877,N_24132,N_24433);
nor U24878 (N_24878,N_24320,N_24496);
xnor U24879 (N_24879,N_24333,N_24163);
xnor U24880 (N_24880,N_24361,N_24249);
nand U24881 (N_24881,N_24295,N_24298);
nand U24882 (N_24882,N_24391,N_24421);
nor U24883 (N_24883,N_24177,N_24314);
or U24884 (N_24884,N_24192,N_24305);
or U24885 (N_24885,N_24100,N_24051);
or U24886 (N_24886,N_24282,N_24147);
or U24887 (N_24887,N_24071,N_24059);
and U24888 (N_24888,N_24082,N_24043);
or U24889 (N_24889,N_24291,N_24047);
or U24890 (N_24890,N_24487,N_24223);
nor U24891 (N_24891,N_24024,N_24497);
nand U24892 (N_24892,N_24373,N_24173);
xor U24893 (N_24893,N_24264,N_24415);
or U24894 (N_24894,N_24168,N_24314);
xor U24895 (N_24895,N_24059,N_24395);
and U24896 (N_24896,N_24465,N_24479);
or U24897 (N_24897,N_24411,N_24144);
or U24898 (N_24898,N_24388,N_24296);
or U24899 (N_24899,N_24326,N_24386);
nand U24900 (N_24900,N_24104,N_24246);
and U24901 (N_24901,N_24205,N_24018);
xor U24902 (N_24902,N_24379,N_24294);
nand U24903 (N_24903,N_24310,N_24099);
nand U24904 (N_24904,N_24382,N_24346);
nand U24905 (N_24905,N_24145,N_24298);
nand U24906 (N_24906,N_24296,N_24439);
nor U24907 (N_24907,N_24032,N_24361);
or U24908 (N_24908,N_24044,N_24475);
and U24909 (N_24909,N_24442,N_24127);
nand U24910 (N_24910,N_24206,N_24487);
and U24911 (N_24911,N_24487,N_24023);
nand U24912 (N_24912,N_24221,N_24007);
nand U24913 (N_24913,N_24177,N_24127);
nand U24914 (N_24914,N_24375,N_24283);
nor U24915 (N_24915,N_24251,N_24003);
and U24916 (N_24916,N_24373,N_24491);
nor U24917 (N_24917,N_24316,N_24139);
and U24918 (N_24918,N_24384,N_24319);
xor U24919 (N_24919,N_24282,N_24036);
or U24920 (N_24920,N_24390,N_24286);
nor U24921 (N_24921,N_24228,N_24276);
nand U24922 (N_24922,N_24002,N_24481);
or U24923 (N_24923,N_24432,N_24245);
or U24924 (N_24924,N_24219,N_24325);
nor U24925 (N_24925,N_24397,N_24346);
nor U24926 (N_24926,N_24113,N_24328);
nor U24927 (N_24927,N_24177,N_24111);
nor U24928 (N_24928,N_24098,N_24366);
nand U24929 (N_24929,N_24473,N_24285);
or U24930 (N_24930,N_24101,N_24303);
and U24931 (N_24931,N_24256,N_24055);
or U24932 (N_24932,N_24218,N_24027);
nor U24933 (N_24933,N_24069,N_24381);
nand U24934 (N_24934,N_24055,N_24338);
nand U24935 (N_24935,N_24256,N_24480);
nor U24936 (N_24936,N_24452,N_24401);
and U24937 (N_24937,N_24457,N_24243);
and U24938 (N_24938,N_24001,N_24474);
nand U24939 (N_24939,N_24399,N_24376);
and U24940 (N_24940,N_24387,N_24303);
or U24941 (N_24941,N_24088,N_24023);
xor U24942 (N_24942,N_24368,N_24414);
nor U24943 (N_24943,N_24412,N_24393);
nor U24944 (N_24944,N_24029,N_24415);
nor U24945 (N_24945,N_24365,N_24278);
or U24946 (N_24946,N_24344,N_24102);
xnor U24947 (N_24947,N_24271,N_24286);
and U24948 (N_24948,N_24398,N_24399);
and U24949 (N_24949,N_24184,N_24044);
or U24950 (N_24950,N_24323,N_24309);
nor U24951 (N_24951,N_24471,N_24037);
and U24952 (N_24952,N_24425,N_24185);
or U24953 (N_24953,N_24452,N_24235);
nor U24954 (N_24954,N_24337,N_24074);
or U24955 (N_24955,N_24293,N_24216);
nor U24956 (N_24956,N_24436,N_24255);
nor U24957 (N_24957,N_24484,N_24218);
nand U24958 (N_24958,N_24070,N_24394);
nor U24959 (N_24959,N_24441,N_24419);
nor U24960 (N_24960,N_24062,N_24191);
nor U24961 (N_24961,N_24284,N_24478);
nor U24962 (N_24962,N_24213,N_24428);
nor U24963 (N_24963,N_24421,N_24035);
nor U24964 (N_24964,N_24453,N_24183);
nand U24965 (N_24965,N_24338,N_24173);
and U24966 (N_24966,N_24117,N_24189);
and U24967 (N_24967,N_24063,N_24459);
and U24968 (N_24968,N_24261,N_24250);
and U24969 (N_24969,N_24356,N_24152);
xor U24970 (N_24970,N_24219,N_24393);
nand U24971 (N_24971,N_24015,N_24148);
nand U24972 (N_24972,N_24372,N_24370);
or U24973 (N_24973,N_24125,N_24264);
xnor U24974 (N_24974,N_24414,N_24037);
nand U24975 (N_24975,N_24188,N_24065);
nor U24976 (N_24976,N_24064,N_24275);
nand U24977 (N_24977,N_24020,N_24054);
or U24978 (N_24978,N_24148,N_24345);
and U24979 (N_24979,N_24251,N_24062);
nand U24980 (N_24980,N_24057,N_24282);
nor U24981 (N_24981,N_24355,N_24373);
and U24982 (N_24982,N_24208,N_24408);
nor U24983 (N_24983,N_24245,N_24412);
nor U24984 (N_24984,N_24139,N_24029);
or U24985 (N_24985,N_24123,N_24347);
and U24986 (N_24986,N_24114,N_24450);
nor U24987 (N_24987,N_24373,N_24180);
xor U24988 (N_24988,N_24362,N_24478);
nor U24989 (N_24989,N_24258,N_24370);
xnor U24990 (N_24990,N_24161,N_24202);
and U24991 (N_24991,N_24405,N_24417);
or U24992 (N_24992,N_24485,N_24374);
and U24993 (N_24993,N_24201,N_24414);
nor U24994 (N_24994,N_24179,N_24370);
and U24995 (N_24995,N_24339,N_24424);
nor U24996 (N_24996,N_24258,N_24304);
or U24997 (N_24997,N_24313,N_24216);
nor U24998 (N_24998,N_24416,N_24126);
or U24999 (N_24999,N_24136,N_24175);
nand U25000 (N_25000,N_24903,N_24871);
nand U25001 (N_25001,N_24588,N_24585);
nor U25002 (N_25002,N_24935,N_24560);
nor U25003 (N_25003,N_24881,N_24906);
and U25004 (N_25004,N_24739,N_24790);
and U25005 (N_25005,N_24643,N_24766);
nor U25006 (N_25006,N_24760,N_24944);
xnor U25007 (N_25007,N_24809,N_24964);
xnor U25008 (N_25008,N_24999,N_24831);
nor U25009 (N_25009,N_24783,N_24889);
or U25010 (N_25010,N_24583,N_24715);
and U25011 (N_25011,N_24846,N_24649);
nor U25012 (N_25012,N_24716,N_24695);
nand U25013 (N_25013,N_24866,N_24902);
nor U25014 (N_25014,N_24896,N_24669);
nand U25015 (N_25015,N_24650,N_24685);
nor U25016 (N_25016,N_24566,N_24569);
or U25017 (N_25017,N_24919,N_24860);
or U25018 (N_25018,N_24688,N_24573);
and U25019 (N_25019,N_24784,N_24642);
nand U25020 (N_25020,N_24820,N_24528);
nand U25021 (N_25021,N_24608,N_24771);
or U25022 (N_25022,N_24674,N_24923);
nor U25023 (N_25023,N_24795,N_24927);
nor U25024 (N_25024,N_24750,N_24587);
nand U25025 (N_25025,N_24780,N_24710);
nor U25026 (N_25026,N_24953,N_24930);
nor U25027 (N_25027,N_24668,N_24811);
and U25028 (N_25028,N_24533,N_24894);
or U25029 (N_25029,N_24842,N_24920);
or U25030 (N_25030,N_24598,N_24752);
or U25031 (N_25031,N_24539,N_24604);
nor U25032 (N_25032,N_24565,N_24523);
and U25033 (N_25033,N_24670,N_24756);
nor U25034 (N_25034,N_24929,N_24709);
or U25035 (N_25035,N_24839,N_24960);
or U25036 (N_25036,N_24757,N_24793);
xnor U25037 (N_25037,N_24991,N_24765);
nand U25038 (N_25038,N_24625,N_24891);
and U25039 (N_25039,N_24838,N_24821);
and U25040 (N_25040,N_24989,N_24720);
nor U25041 (N_25041,N_24713,N_24653);
or U25042 (N_25042,N_24869,N_24582);
xor U25043 (N_25043,N_24632,N_24753);
and U25044 (N_25044,N_24988,N_24961);
xnor U25045 (N_25045,N_24942,N_24531);
nor U25046 (N_25046,N_24652,N_24725);
or U25047 (N_25047,N_24778,N_24802);
or U25048 (N_25048,N_24622,N_24729);
xnor U25049 (N_25049,N_24648,N_24855);
nand U25050 (N_25050,N_24593,N_24629);
or U25051 (N_25051,N_24536,N_24967);
nor U25052 (N_25052,N_24799,N_24851);
and U25053 (N_25053,N_24703,N_24601);
and U25054 (N_25054,N_24665,N_24534);
or U25055 (N_25055,N_24529,N_24506);
nor U25056 (N_25056,N_24637,N_24873);
or U25057 (N_25057,N_24549,N_24812);
and U25058 (N_25058,N_24913,N_24594);
or U25059 (N_25059,N_24887,N_24907);
and U25060 (N_25060,N_24664,N_24511);
nor U25061 (N_25061,N_24574,N_24797);
and U25062 (N_25062,N_24614,N_24563);
and U25063 (N_25063,N_24973,N_24833);
and U25064 (N_25064,N_24879,N_24883);
nand U25065 (N_25065,N_24655,N_24639);
or U25066 (N_25066,N_24619,N_24740);
nor U25067 (N_25067,N_24509,N_24603);
and U25068 (N_25068,N_24801,N_24767);
xnor U25069 (N_25069,N_24521,N_24829);
nor U25070 (N_25070,N_24863,N_24749);
nand U25071 (N_25071,N_24792,N_24626);
and U25072 (N_25072,N_24949,N_24647);
nor U25073 (N_25073,N_24900,N_24575);
nor U25074 (N_25074,N_24915,N_24702);
or U25075 (N_25075,N_24644,N_24950);
and U25076 (N_25076,N_24692,N_24611);
nand U25077 (N_25077,N_24803,N_24963);
and U25078 (N_25078,N_24719,N_24865);
nand U25079 (N_25079,N_24623,N_24818);
and U25080 (N_25080,N_24607,N_24576);
or U25081 (N_25081,N_24736,N_24980);
and U25082 (N_25082,N_24718,N_24584);
nand U25083 (N_25083,N_24545,N_24578);
and U25084 (N_25084,N_24813,N_24504);
nand U25085 (N_25085,N_24946,N_24975);
xnor U25086 (N_25086,N_24662,N_24698);
nor U25087 (N_25087,N_24520,N_24852);
nand U25088 (N_25088,N_24597,N_24782);
nand U25089 (N_25089,N_24707,N_24502);
nor U25090 (N_25090,N_24675,N_24606);
or U25091 (N_25091,N_24610,N_24876);
xor U25092 (N_25092,N_24553,N_24505);
or U25093 (N_25093,N_24910,N_24895);
and U25094 (N_25094,N_24514,N_24556);
nand U25095 (N_25095,N_24878,N_24774);
nor U25096 (N_25096,N_24911,N_24945);
or U25097 (N_25097,N_24971,N_24554);
nand U25098 (N_25098,N_24886,N_24965);
and U25099 (N_25099,N_24954,N_24701);
nor U25100 (N_25100,N_24525,N_24691);
or U25101 (N_25101,N_24787,N_24741);
and U25102 (N_25102,N_24853,N_24618);
and U25103 (N_25103,N_24872,N_24806);
nand U25104 (N_25104,N_24624,N_24661);
nand U25105 (N_25105,N_24734,N_24515);
or U25106 (N_25106,N_24807,N_24956);
nand U25107 (N_25107,N_24850,N_24599);
xor U25108 (N_25108,N_24867,N_24969);
nand U25109 (N_25109,N_24837,N_24826);
nand U25110 (N_25110,N_24777,N_24737);
and U25111 (N_25111,N_24687,N_24640);
xnor U25112 (N_25112,N_24555,N_24762);
nand U25113 (N_25113,N_24841,N_24755);
or U25114 (N_25114,N_24526,N_24815);
or U25115 (N_25115,N_24579,N_24540);
xnor U25116 (N_25116,N_24538,N_24909);
nor U25117 (N_25117,N_24700,N_24816);
nand U25118 (N_25118,N_24830,N_24849);
or U25119 (N_25119,N_24683,N_24705);
nand U25120 (N_25120,N_24660,N_24800);
nor U25121 (N_25121,N_24985,N_24918);
nand U25122 (N_25122,N_24759,N_24602);
nand U25123 (N_25123,N_24684,N_24620);
and U25124 (N_25124,N_24877,N_24825);
and U25125 (N_25125,N_24532,N_24656);
or U25126 (N_25126,N_24596,N_24657);
nand U25127 (N_25127,N_24542,N_24951);
or U25128 (N_25128,N_24905,N_24933);
or U25129 (N_25129,N_24925,N_24912);
nand U25130 (N_25130,N_24834,N_24763);
nor U25131 (N_25131,N_24678,N_24559);
nor U25132 (N_25132,N_24519,N_24987);
or U25133 (N_25133,N_24547,N_24730);
xnor U25134 (N_25134,N_24970,N_24781);
nand U25135 (N_25135,N_24864,N_24690);
nand U25136 (N_25136,N_24546,N_24982);
or U25137 (N_25137,N_24998,N_24630);
nand U25138 (N_25138,N_24997,N_24748);
xor U25139 (N_25139,N_24577,N_24893);
nor U25140 (N_25140,N_24890,N_24580);
nand U25141 (N_25141,N_24571,N_24828);
and U25142 (N_25142,N_24609,N_24503);
nor U25143 (N_25143,N_24775,N_24827);
xnor U25144 (N_25144,N_24804,N_24861);
xor U25145 (N_25145,N_24731,N_24798);
nor U25146 (N_25146,N_24557,N_24938);
or U25147 (N_25147,N_24654,N_24810);
or U25148 (N_25148,N_24617,N_24732);
nor U25149 (N_25149,N_24727,N_24501);
and U25150 (N_25150,N_24844,N_24974);
and U25151 (N_25151,N_24758,N_24904);
nand U25152 (N_25152,N_24817,N_24516);
and U25153 (N_25153,N_24616,N_24633);
or U25154 (N_25154,N_24940,N_24544);
or U25155 (N_25155,N_24507,N_24641);
nor U25156 (N_25156,N_24561,N_24764);
nand U25157 (N_25157,N_24983,N_24972);
and U25158 (N_25158,N_24990,N_24882);
and U25159 (N_25159,N_24943,N_24550);
and U25160 (N_25160,N_24892,N_24543);
nor U25161 (N_25161,N_24722,N_24681);
nand U25162 (N_25162,N_24976,N_24667);
or U25163 (N_25163,N_24981,N_24885);
nor U25164 (N_25164,N_24677,N_24676);
nor U25165 (N_25165,N_24794,N_24570);
or U25166 (N_25166,N_24773,N_24984);
nand U25167 (N_25167,N_24897,N_24615);
nand U25168 (N_25168,N_24673,N_24992);
nand U25169 (N_25169,N_24856,N_24671);
nor U25170 (N_25170,N_24776,N_24635);
and U25171 (N_25171,N_24926,N_24843);
nand U25172 (N_25172,N_24779,N_24917);
nand U25173 (N_25173,N_24805,N_24789);
nor U25174 (N_25174,N_24979,N_24847);
or U25175 (N_25175,N_24510,N_24937);
or U25176 (N_25176,N_24589,N_24962);
nor U25177 (N_25177,N_24693,N_24880);
nor U25178 (N_25178,N_24738,N_24680);
nor U25179 (N_25179,N_24552,N_24939);
nand U25180 (N_25180,N_24541,N_24754);
or U25181 (N_25181,N_24899,N_24518);
or U25182 (N_25182,N_24530,N_24814);
and U25183 (N_25183,N_24697,N_24986);
or U25184 (N_25184,N_24977,N_24823);
nand U25185 (N_25185,N_24744,N_24572);
or U25186 (N_25186,N_24564,N_24706);
and U25187 (N_25187,N_24666,N_24735);
nor U25188 (N_25188,N_24908,N_24854);
nor U25189 (N_25189,N_24934,N_24862);
nand U25190 (N_25190,N_24936,N_24832);
nor U25191 (N_25191,N_24808,N_24634);
or U25192 (N_25192,N_24875,N_24708);
or U25193 (N_25193,N_24931,N_24835);
and U25194 (N_25194,N_24743,N_24558);
nor U25195 (N_25195,N_24955,N_24791);
or U25196 (N_25196,N_24612,N_24567);
and U25197 (N_25197,N_24659,N_24636);
and U25198 (N_25198,N_24724,N_24627);
nand U25199 (N_25199,N_24884,N_24796);
nor U25200 (N_25200,N_24848,N_24586);
nor U25201 (N_25201,N_24845,N_24605);
nand U25202 (N_25202,N_24682,N_24742);
xnor U25203 (N_25203,N_24524,N_24613);
nor U25204 (N_25204,N_24726,N_24958);
nor U25205 (N_25205,N_24996,N_24761);
xnor U25206 (N_25206,N_24568,N_24508);
nor U25207 (N_25207,N_24788,N_24840);
nand U25208 (N_25208,N_24527,N_24548);
nand U25209 (N_25209,N_24957,N_24948);
nor U25210 (N_25210,N_24858,N_24590);
and U25211 (N_25211,N_24914,N_24745);
or U25212 (N_25212,N_24645,N_24751);
and U25213 (N_25213,N_24786,N_24723);
nand U25214 (N_25214,N_24686,N_24966);
nand U25215 (N_25215,N_24733,N_24711);
nor U25216 (N_25216,N_24921,N_24898);
nand U25217 (N_25217,N_24663,N_24968);
and U25218 (N_25218,N_24699,N_24819);
nand U25219 (N_25219,N_24714,N_24631);
and U25220 (N_25220,N_24689,N_24746);
nand U25221 (N_25221,N_24646,N_24562);
nor U25222 (N_25222,N_24512,N_24901);
nand U25223 (N_25223,N_24628,N_24952);
nand U25224 (N_25224,N_24870,N_24704);
and U25225 (N_25225,N_24747,N_24772);
or U25226 (N_25226,N_24959,N_24836);
nand U25227 (N_25227,N_24947,N_24551);
xor U25228 (N_25228,N_24868,N_24822);
or U25229 (N_25229,N_24728,N_24717);
or U25230 (N_25230,N_24522,N_24672);
nand U25231 (N_25231,N_24994,N_24769);
nand U25232 (N_25232,N_24658,N_24785);
or U25233 (N_25233,N_24857,N_24537);
nand U25234 (N_25234,N_24621,N_24517);
or U25235 (N_25235,N_24638,N_24694);
nor U25236 (N_25236,N_24768,N_24824);
nor U25237 (N_25237,N_24595,N_24978);
nand U25238 (N_25238,N_24922,N_24928);
nor U25239 (N_25239,N_24770,N_24712);
nand U25240 (N_25240,N_24859,N_24535);
and U25241 (N_25241,N_24679,N_24592);
and U25242 (N_25242,N_24941,N_24916);
and U25243 (N_25243,N_24591,N_24696);
or U25244 (N_25244,N_24932,N_24874);
xor U25245 (N_25245,N_24651,N_24995);
xnor U25246 (N_25246,N_24888,N_24924);
or U25247 (N_25247,N_24721,N_24993);
nand U25248 (N_25248,N_24500,N_24600);
and U25249 (N_25249,N_24581,N_24513);
nor U25250 (N_25250,N_24846,N_24520);
xnor U25251 (N_25251,N_24654,N_24641);
and U25252 (N_25252,N_24558,N_24900);
nor U25253 (N_25253,N_24734,N_24969);
and U25254 (N_25254,N_24880,N_24924);
nor U25255 (N_25255,N_24551,N_24809);
or U25256 (N_25256,N_24628,N_24660);
nor U25257 (N_25257,N_24829,N_24737);
or U25258 (N_25258,N_24686,N_24605);
xnor U25259 (N_25259,N_24603,N_24974);
xnor U25260 (N_25260,N_24828,N_24976);
xnor U25261 (N_25261,N_24942,N_24566);
or U25262 (N_25262,N_24853,N_24921);
and U25263 (N_25263,N_24935,N_24578);
nand U25264 (N_25264,N_24898,N_24959);
and U25265 (N_25265,N_24811,N_24963);
and U25266 (N_25266,N_24526,N_24780);
and U25267 (N_25267,N_24690,N_24556);
and U25268 (N_25268,N_24525,N_24847);
and U25269 (N_25269,N_24750,N_24700);
nand U25270 (N_25270,N_24911,N_24508);
nand U25271 (N_25271,N_24571,N_24500);
or U25272 (N_25272,N_24825,N_24610);
and U25273 (N_25273,N_24926,N_24886);
nand U25274 (N_25274,N_24763,N_24822);
and U25275 (N_25275,N_24852,N_24817);
and U25276 (N_25276,N_24560,N_24586);
or U25277 (N_25277,N_24844,N_24515);
nand U25278 (N_25278,N_24866,N_24638);
or U25279 (N_25279,N_24797,N_24915);
and U25280 (N_25280,N_24538,N_24903);
and U25281 (N_25281,N_24841,N_24667);
nand U25282 (N_25282,N_24663,N_24592);
nor U25283 (N_25283,N_24647,N_24538);
and U25284 (N_25284,N_24615,N_24943);
nand U25285 (N_25285,N_24632,N_24754);
or U25286 (N_25286,N_24903,N_24588);
and U25287 (N_25287,N_24634,N_24639);
nor U25288 (N_25288,N_24653,N_24531);
or U25289 (N_25289,N_24631,N_24900);
and U25290 (N_25290,N_24649,N_24739);
nand U25291 (N_25291,N_24827,N_24829);
nor U25292 (N_25292,N_24999,N_24696);
nor U25293 (N_25293,N_24996,N_24759);
nand U25294 (N_25294,N_24792,N_24977);
or U25295 (N_25295,N_24758,N_24559);
and U25296 (N_25296,N_24873,N_24986);
nor U25297 (N_25297,N_24609,N_24551);
and U25298 (N_25298,N_24642,N_24695);
nor U25299 (N_25299,N_24815,N_24933);
nand U25300 (N_25300,N_24999,N_24974);
nand U25301 (N_25301,N_24708,N_24681);
xnor U25302 (N_25302,N_24938,N_24652);
or U25303 (N_25303,N_24659,N_24884);
and U25304 (N_25304,N_24682,N_24933);
nand U25305 (N_25305,N_24743,N_24644);
nor U25306 (N_25306,N_24961,N_24696);
xnor U25307 (N_25307,N_24725,N_24926);
or U25308 (N_25308,N_24902,N_24688);
and U25309 (N_25309,N_24823,N_24925);
nor U25310 (N_25310,N_24694,N_24914);
nand U25311 (N_25311,N_24526,N_24566);
xor U25312 (N_25312,N_24904,N_24883);
nor U25313 (N_25313,N_24771,N_24908);
and U25314 (N_25314,N_24611,N_24717);
nand U25315 (N_25315,N_24812,N_24548);
or U25316 (N_25316,N_24879,N_24598);
xor U25317 (N_25317,N_24567,N_24817);
or U25318 (N_25318,N_24864,N_24878);
nand U25319 (N_25319,N_24722,N_24789);
nor U25320 (N_25320,N_24658,N_24987);
nor U25321 (N_25321,N_24942,N_24877);
and U25322 (N_25322,N_24643,N_24702);
and U25323 (N_25323,N_24800,N_24690);
and U25324 (N_25324,N_24858,N_24518);
or U25325 (N_25325,N_24560,N_24739);
or U25326 (N_25326,N_24572,N_24546);
nand U25327 (N_25327,N_24623,N_24685);
and U25328 (N_25328,N_24547,N_24823);
nand U25329 (N_25329,N_24762,N_24862);
nor U25330 (N_25330,N_24892,N_24744);
or U25331 (N_25331,N_24713,N_24584);
nor U25332 (N_25332,N_24558,N_24681);
nor U25333 (N_25333,N_24685,N_24624);
nor U25334 (N_25334,N_24504,N_24510);
or U25335 (N_25335,N_24553,N_24968);
nor U25336 (N_25336,N_24845,N_24981);
or U25337 (N_25337,N_24528,N_24681);
and U25338 (N_25338,N_24834,N_24626);
and U25339 (N_25339,N_24931,N_24747);
and U25340 (N_25340,N_24543,N_24777);
nor U25341 (N_25341,N_24967,N_24717);
xnor U25342 (N_25342,N_24694,N_24762);
and U25343 (N_25343,N_24703,N_24568);
nand U25344 (N_25344,N_24661,N_24697);
nand U25345 (N_25345,N_24516,N_24791);
or U25346 (N_25346,N_24505,N_24535);
xor U25347 (N_25347,N_24822,N_24792);
nor U25348 (N_25348,N_24970,N_24512);
and U25349 (N_25349,N_24521,N_24863);
xnor U25350 (N_25350,N_24977,N_24903);
nand U25351 (N_25351,N_24931,N_24913);
nand U25352 (N_25352,N_24793,N_24854);
nand U25353 (N_25353,N_24709,N_24830);
or U25354 (N_25354,N_24816,N_24767);
nand U25355 (N_25355,N_24728,N_24790);
nor U25356 (N_25356,N_24594,N_24573);
nand U25357 (N_25357,N_24676,N_24914);
nor U25358 (N_25358,N_24897,N_24559);
and U25359 (N_25359,N_24671,N_24807);
or U25360 (N_25360,N_24850,N_24678);
nand U25361 (N_25361,N_24552,N_24952);
or U25362 (N_25362,N_24501,N_24568);
nor U25363 (N_25363,N_24709,N_24754);
nand U25364 (N_25364,N_24678,N_24556);
nand U25365 (N_25365,N_24788,N_24748);
nand U25366 (N_25366,N_24767,N_24540);
and U25367 (N_25367,N_24660,N_24850);
or U25368 (N_25368,N_24795,N_24708);
nor U25369 (N_25369,N_24773,N_24630);
and U25370 (N_25370,N_24730,N_24594);
and U25371 (N_25371,N_24910,N_24913);
and U25372 (N_25372,N_24813,N_24839);
and U25373 (N_25373,N_24868,N_24995);
or U25374 (N_25374,N_24655,N_24523);
and U25375 (N_25375,N_24635,N_24716);
or U25376 (N_25376,N_24729,N_24733);
nand U25377 (N_25377,N_24871,N_24582);
and U25378 (N_25378,N_24798,N_24592);
nand U25379 (N_25379,N_24951,N_24797);
nand U25380 (N_25380,N_24560,N_24675);
and U25381 (N_25381,N_24816,N_24694);
and U25382 (N_25382,N_24626,N_24934);
and U25383 (N_25383,N_24564,N_24584);
or U25384 (N_25384,N_24634,N_24797);
or U25385 (N_25385,N_24618,N_24977);
xor U25386 (N_25386,N_24503,N_24574);
nor U25387 (N_25387,N_24928,N_24835);
or U25388 (N_25388,N_24857,N_24614);
nor U25389 (N_25389,N_24665,N_24868);
nand U25390 (N_25390,N_24626,N_24549);
nand U25391 (N_25391,N_24865,N_24715);
nand U25392 (N_25392,N_24548,N_24784);
nor U25393 (N_25393,N_24642,N_24872);
and U25394 (N_25394,N_24820,N_24590);
nand U25395 (N_25395,N_24559,N_24535);
nor U25396 (N_25396,N_24565,N_24713);
or U25397 (N_25397,N_24585,N_24539);
nor U25398 (N_25398,N_24711,N_24963);
xor U25399 (N_25399,N_24841,N_24995);
xnor U25400 (N_25400,N_24972,N_24757);
or U25401 (N_25401,N_24651,N_24692);
or U25402 (N_25402,N_24515,N_24778);
nor U25403 (N_25403,N_24896,N_24522);
or U25404 (N_25404,N_24658,N_24891);
xor U25405 (N_25405,N_24787,N_24806);
and U25406 (N_25406,N_24573,N_24826);
and U25407 (N_25407,N_24669,N_24848);
nor U25408 (N_25408,N_24744,N_24589);
nand U25409 (N_25409,N_24509,N_24865);
and U25410 (N_25410,N_24828,N_24915);
or U25411 (N_25411,N_24939,N_24704);
xor U25412 (N_25412,N_24898,N_24739);
nor U25413 (N_25413,N_24590,N_24604);
or U25414 (N_25414,N_24814,N_24917);
and U25415 (N_25415,N_24699,N_24887);
nor U25416 (N_25416,N_24947,N_24530);
or U25417 (N_25417,N_24558,N_24895);
nand U25418 (N_25418,N_24532,N_24815);
or U25419 (N_25419,N_24676,N_24972);
nor U25420 (N_25420,N_24914,N_24657);
or U25421 (N_25421,N_24966,N_24797);
nor U25422 (N_25422,N_24875,N_24554);
xor U25423 (N_25423,N_24880,N_24646);
nand U25424 (N_25424,N_24964,N_24582);
or U25425 (N_25425,N_24751,N_24688);
nand U25426 (N_25426,N_24784,N_24811);
or U25427 (N_25427,N_24765,N_24803);
and U25428 (N_25428,N_24600,N_24794);
nand U25429 (N_25429,N_24619,N_24790);
or U25430 (N_25430,N_24995,N_24560);
and U25431 (N_25431,N_24538,N_24513);
nand U25432 (N_25432,N_24968,N_24940);
and U25433 (N_25433,N_24965,N_24535);
or U25434 (N_25434,N_24977,N_24775);
and U25435 (N_25435,N_24638,N_24639);
or U25436 (N_25436,N_24897,N_24592);
and U25437 (N_25437,N_24815,N_24547);
and U25438 (N_25438,N_24583,N_24699);
or U25439 (N_25439,N_24757,N_24665);
and U25440 (N_25440,N_24972,N_24943);
xor U25441 (N_25441,N_24805,N_24901);
or U25442 (N_25442,N_24648,N_24559);
and U25443 (N_25443,N_24823,N_24962);
and U25444 (N_25444,N_24570,N_24846);
or U25445 (N_25445,N_24681,N_24955);
nand U25446 (N_25446,N_24959,N_24634);
or U25447 (N_25447,N_24967,N_24599);
and U25448 (N_25448,N_24777,N_24962);
or U25449 (N_25449,N_24752,N_24537);
nor U25450 (N_25450,N_24677,N_24513);
or U25451 (N_25451,N_24599,N_24961);
nor U25452 (N_25452,N_24973,N_24893);
nand U25453 (N_25453,N_24801,N_24949);
nor U25454 (N_25454,N_24516,N_24779);
nor U25455 (N_25455,N_24673,N_24815);
xnor U25456 (N_25456,N_24902,N_24600);
nor U25457 (N_25457,N_24874,N_24744);
nor U25458 (N_25458,N_24640,N_24595);
or U25459 (N_25459,N_24562,N_24676);
nor U25460 (N_25460,N_24775,N_24859);
or U25461 (N_25461,N_24507,N_24666);
and U25462 (N_25462,N_24804,N_24994);
and U25463 (N_25463,N_24809,N_24606);
and U25464 (N_25464,N_24882,N_24509);
or U25465 (N_25465,N_24913,N_24752);
nand U25466 (N_25466,N_24737,N_24502);
xor U25467 (N_25467,N_24688,N_24960);
nand U25468 (N_25468,N_24931,N_24789);
or U25469 (N_25469,N_24792,N_24521);
nand U25470 (N_25470,N_24648,N_24857);
or U25471 (N_25471,N_24761,N_24918);
and U25472 (N_25472,N_24574,N_24941);
or U25473 (N_25473,N_24507,N_24674);
or U25474 (N_25474,N_24596,N_24527);
nand U25475 (N_25475,N_24970,N_24769);
nor U25476 (N_25476,N_24791,N_24696);
and U25477 (N_25477,N_24908,N_24757);
nor U25478 (N_25478,N_24852,N_24931);
or U25479 (N_25479,N_24596,N_24632);
xor U25480 (N_25480,N_24833,N_24757);
or U25481 (N_25481,N_24606,N_24713);
or U25482 (N_25482,N_24601,N_24850);
nand U25483 (N_25483,N_24574,N_24996);
or U25484 (N_25484,N_24769,N_24907);
xor U25485 (N_25485,N_24995,N_24763);
nor U25486 (N_25486,N_24698,N_24571);
nand U25487 (N_25487,N_24507,N_24993);
xnor U25488 (N_25488,N_24568,N_24727);
nor U25489 (N_25489,N_24904,N_24664);
nand U25490 (N_25490,N_24809,N_24957);
xor U25491 (N_25491,N_24701,N_24746);
nand U25492 (N_25492,N_24889,N_24620);
nor U25493 (N_25493,N_24762,N_24570);
nand U25494 (N_25494,N_24829,N_24905);
xnor U25495 (N_25495,N_24633,N_24594);
nor U25496 (N_25496,N_24712,N_24671);
and U25497 (N_25497,N_24950,N_24692);
nand U25498 (N_25498,N_24714,N_24518);
nand U25499 (N_25499,N_24871,N_24638);
and U25500 (N_25500,N_25398,N_25258);
nor U25501 (N_25501,N_25439,N_25355);
nand U25502 (N_25502,N_25382,N_25307);
nor U25503 (N_25503,N_25464,N_25026);
and U25504 (N_25504,N_25094,N_25342);
and U25505 (N_25505,N_25075,N_25227);
nand U25506 (N_25506,N_25270,N_25202);
nor U25507 (N_25507,N_25074,N_25318);
and U25508 (N_25508,N_25395,N_25169);
or U25509 (N_25509,N_25259,N_25172);
nor U25510 (N_25510,N_25397,N_25160);
nor U25511 (N_25511,N_25185,N_25337);
nor U25512 (N_25512,N_25155,N_25403);
nor U25513 (N_25513,N_25288,N_25377);
or U25514 (N_25514,N_25488,N_25257);
nor U25515 (N_25515,N_25113,N_25412);
nand U25516 (N_25516,N_25437,N_25388);
or U25517 (N_25517,N_25251,N_25289);
or U25518 (N_25518,N_25080,N_25046);
nor U25519 (N_25519,N_25170,N_25084);
nand U25520 (N_25520,N_25162,N_25021);
nor U25521 (N_25521,N_25306,N_25035);
nor U25522 (N_25522,N_25285,N_25315);
xnor U25523 (N_25523,N_25472,N_25276);
xor U25524 (N_25524,N_25128,N_25373);
xor U25525 (N_25525,N_25062,N_25233);
or U25526 (N_25526,N_25129,N_25201);
nand U25527 (N_25527,N_25441,N_25436);
nand U25528 (N_25528,N_25340,N_25376);
and U25529 (N_25529,N_25279,N_25192);
xor U25530 (N_25530,N_25426,N_25438);
nor U25531 (N_25531,N_25256,N_25011);
nand U25532 (N_25532,N_25103,N_25245);
nor U25533 (N_25533,N_25061,N_25043);
nor U25534 (N_25534,N_25098,N_25089);
nor U25535 (N_25535,N_25273,N_25165);
nand U25536 (N_25536,N_25252,N_25299);
and U25537 (N_25537,N_25283,N_25174);
and U25538 (N_25538,N_25459,N_25339);
nor U25539 (N_25539,N_25360,N_25331);
and U25540 (N_25540,N_25460,N_25215);
nor U25541 (N_25541,N_25321,N_25404);
and U25542 (N_25542,N_25137,N_25349);
nand U25543 (N_25543,N_25292,N_25456);
or U25544 (N_25544,N_25275,N_25146);
or U25545 (N_25545,N_25230,N_25486);
or U25546 (N_25546,N_25371,N_25317);
nand U25547 (N_25547,N_25153,N_25301);
and U25548 (N_25548,N_25217,N_25281);
nand U25549 (N_25549,N_25417,N_25478);
nor U25550 (N_25550,N_25343,N_25222);
and U25551 (N_25551,N_25225,N_25498);
or U25552 (N_25552,N_25189,N_25408);
or U25553 (N_25553,N_25370,N_25167);
nand U25554 (N_25554,N_25381,N_25243);
or U25555 (N_25555,N_25302,N_25467);
nor U25556 (N_25556,N_25314,N_25250);
and U25557 (N_25557,N_25284,N_25271);
nor U25558 (N_25558,N_25014,N_25124);
nand U25559 (N_25559,N_25244,N_25042);
or U25560 (N_25560,N_25158,N_25198);
nand U25561 (N_25561,N_25248,N_25034);
or U25562 (N_25562,N_25325,N_25450);
or U25563 (N_25563,N_25296,N_25221);
nand U25564 (N_25564,N_25290,N_25096);
nor U25565 (N_25565,N_25088,N_25131);
or U25566 (N_25566,N_25140,N_25375);
nand U25567 (N_25567,N_25183,N_25237);
nor U25568 (N_25568,N_25380,N_25324);
or U25569 (N_25569,N_25440,N_25040);
nor U25570 (N_25570,N_25102,N_25383);
nor U25571 (N_25571,N_25235,N_25418);
and U25572 (N_25572,N_25175,N_25009);
and U25573 (N_25573,N_25423,N_25070);
nand U25574 (N_25574,N_25204,N_25414);
and U25575 (N_25575,N_25017,N_25186);
and U25576 (N_25576,N_25006,N_25372);
nand U25577 (N_25577,N_25309,N_25038);
or U25578 (N_25578,N_25166,N_25127);
or U25579 (N_25579,N_25462,N_25051);
and U25580 (N_25580,N_25210,N_25039);
and U25581 (N_25581,N_25219,N_25308);
nand U25582 (N_25582,N_25120,N_25249);
and U25583 (N_25583,N_25067,N_25126);
and U25584 (N_25584,N_25068,N_25135);
nor U25585 (N_25585,N_25147,N_25143);
nor U25586 (N_25586,N_25367,N_25463);
nor U25587 (N_25587,N_25311,N_25136);
or U25588 (N_25588,N_25013,N_25001);
and U25589 (N_25589,N_25291,N_25150);
and U25590 (N_25590,N_25180,N_25260);
nor U25591 (N_25591,N_25176,N_25108);
and U25592 (N_25592,N_25416,N_25332);
and U25593 (N_25593,N_25117,N_25037);
nand U25594 (N_25594,N_25393,N_25220);
and U25595 (N_25595,N_25479,N_25020);
nand U25596 (N_25596,N_25442,N_25238);
nand U25597 (N_25597,N_25207,N_25200);
nand U25598 (N_25598,N_25358,N_25141);
nor U25599 (N_25599,N_25066,N_25179);
or U25600 (N_25600,N_25104,N_25214);
nor U25601 (N_25601,N_25193,N_25163);
and U25602 (N_25602,N_25000,N_25338);
nor U25603 (N_25603,N_25254,N_25224);
nand U25604 (N_25604,N_25287,N_25030);
or U25605 (N_25605,N_25407,N_25057);
nand U25606 (N_25606,N_25101,N_25389);
or U25607 (N_25607,N_25424,N_25125);
nor U25608 (N_25608,N_25234,N_25316);
nand U25609 (N_25609,N_25494,N_25100);
nor U25610 (N_25610,N_25240,N_25282);
nor U25611 (N_25611,N_25497,N_25277);
nand U25612 (N_25612,N_25263,N_25022);
and U25613 (N_25613,N_25199,N_25151);
nor U25614 (N_25614,N_25490,N_25181);
xnor U25615 (N_25615,N_25378,N_25480);
or U25616 (N_25616,N_25032,N_25392);
xor U25617 (N_25617,N_25365,N_25431);
and U25618 (N_25618,N_25148,N_25123);
nand U25619 (N_25619,N_25298,N_25267);
or U25620 (N_25620,N_25093,N_25313);
xnor U25621 (N_25621,N_25402,N_25405);
nand U25622 (N_25622,N_25171,N_25081);
or U25623 (N_25623,N_25229,N_25159);
nand U25624 (N_25624,N_25194,N_25491);
or U25625 (N_25625,N_25465,N_25453);
nand U25626 (N_25626,N_25029,N_25008);
nand U25627 (N_25627,N_25203,N_25354);
and U25628 (N_25628,N_25114,N_25335);
nor U25629 (N_25629,N_25269,N_25266);
and U25630 (N_25630,N_25481,N_25005);
nand U25631 (N_25631,N_25149,N_25322);
and U25632 (N_25632,N_25419,N_25087);
xor U25633 (N_25633,N_25468,N_25359);
xnor U25634 (N_25634,N_25107,N_25063);
and U25635 (N_25635,N_25330,N_25073);
and U25636 (N_25636,N_25195,N_25487);
nand U25637 (N_25637,N_25293,N_25178);
and U25638 (N_25638,N_25188,N_25430);
xor U25639 (N_25639,N_25305,N_25482);
and U25640 (N_25640,N_25329,N_25493);
nor U25641 (N_25641,N_25484,N_25461);
nand U25642 (N_25642,N_25246,N_25091);
nand U25643 (N_25643,N_25010,N_25433);
and U25644 (N_25644,N_25023,N_25223);
nor U25645 (N_25645,N_25134,N_25092);
and U25646 (N_25646,N_25396,N_25344);
nand U25647 (N_25647,N_25420,N_25077);
or U25648 (N_25648,N_25352,N_25242);
xor U25649 (N_25649,N_25489,N_25320);
nand U25650 (N_25650,N_25390,N_25004);
or U25651 (N_25651,N_25144,N_25012);
nand U25652 (N_25652,N_25212,N_25054);
or U25653 (N_25653,N_25142,N_25112);
nand U25654 (N_25654,N_25157,N_25110);
or U25655 (N_25655,N_25427,N_25268);
or U25656 (N_25656,N_25394,N_25278);
nand U25657 (N_25657,N_25095,N_25016);
xnor U25658 (N_25658,N_25492,N_25466);
or U25659 (N_25659,N_25319,N_25025);
or U25660 (N_25660,N_25297,N_25205);
or U25661 (N_25661,N_25083,N_25072);
nor U25662 (N_25662,N_25323,N_25122);
nand U25663 (N_25663,N_25121,N_25443);
or U25664 (N_25664,N_25105,N_25085);
xnor U25665 (N_25665,N_25056,N_25184);
nand U25666 (N_25666,N_25346,N_25231);
nor U25667 (N_25667,N_25152,N_25187);
nor U25668 (N_25668,N_25018,N_25048);
and U25669 (N_25669,N_25304,N_25274);
nor U25670 (N_25670,N_25253,N_25024);
nor U25671 (N_25671,N_25280,N_25471);
and U25672 (N_25672,N_25448,N_25347);
and U25673 (N_25673,N_25469,N_25138);
nor U25674 (N_25674,N_25064,N_25476);
and U25675 (N_25675,N_25435,N_25044);
and U25676 (N_25676,N_25033,N_25058);
nor U25677 (N_25677,N_25115,N_25421);
nand U25678 (N_25678,N_25050,N_25272);
nand U25679 (N_25679,N_25399,N_25161);
or U25680 (N_25680,N_25387,N_25164);
or U25681 (N_25681,N_25239,N_25019);
xnor U25682 (N_25682,N_25116,N_25356);
or U25683 (N_25683,N_25090,N_25391);
nor U25684 (N_25684,N_25078,N_25097);
nor U25685 (N_25685,N_25213,N_25052);
or U25686 (N_25686,N_25379,N_25082);
nand U25687 (N_25687,N_25197,N_25357);
or U25688 (N_25688,N_25353,N_25428);
nor U25689 (N_25689,N_25099,N_25053);
or U25690 (N_25690,N_25341,N_25328);
and U25691 (N_25691,N_25401,N_25232);
or U25692 (N_25692,N_25031,N_25457);
nor U25693 (N_25693,N_25363,N_25485);
or U25694 (N_25694,N_25060,N_25310);
and U25695 (N_25695,N_25139,N_25059);
and U25696 (N_25696,N_25345,N_25434);
or U25697 (N_25697,N_25015,N_25133);
and U25698 (N_25698,N_25470,N_25451);
or U25699 (N_25699,N_25429,N_25262);
and U25700 (N_25700,N_25445,N_25411);
and U25701 (N_25701,N_25236,N_25473);
nor U25702 (N_25702,N_25362,N_25496);
and U25703 (N_25703,N_25196,N_25351);
nand U25704 (N_25704,N_25079,N_25300);
xnor U25705 (N_25705,N_25047,N_25190);
nor U25706 (N_25706,N_25182,N_25368);
xor U25707 (N_25707,N_25173,N_25415);
and U25708 (N_25708,N_25111,N_25495);
and U25709 (N_25709,N_25264,N_25336);
nand U25710 (N_25710,N_25286,N_25261);
and U25711 (N_25711,N_25409,N_25002);
nand U25712 (N_25712,N_25369,N_25425);
nor U25713 (N_25713,N_25130,N_25410);
nand U25714 (N_25714,N_25477,N_25265);
nor U25715 (N_25715,N_25191,N_25446);
nor U25716 (N_25716,N_25168,N_25086);
nor U25717 (N_25717,N_25449,N_25350);
or U25718 (N_25718,N_25109,N_25474);
nand U25719 (N_25719,N_25326,N_25400);
nor U25720 (N_25720,N_25228,N_25003);
or U25721 (N_25721,N_25294,N_25364);
nand U25722 (N_25722,N_25444,N_25154);
xnor U25723 (N_25723,N_25384,N_25361);
nand U25724 (N_25724,N_25156,N_25385);
nor U25725 (N_25725,N_25366,N_25071);
nor U25726 (N_25726,N_25247,N_25455);
nor U25727 (N_25727,N_25255,N_25007);
nand U25728 (N_25728,N_25447,N_25374);
and U25729 (N_25729,N_25119,N_25432);
nand U25730 (N_25730,N_25312,N_25483);
xor U25731 (N_25731,N_25208,N_25177);
or U25732 (N_25732,N_25295,N_25027);
xor U25733 (N_25733,N_25036,N_25218);
nor U25734 (N_25734,N_25303,N_25386);
nand U25735 (N_25735,N_25216,N_25413);
or U25736 (N_25736,N_25334,N_25452);
nand U25737 (N_25737,N_25226,N_25065);
and U25738 (N_25738,N_25132,N_25076);
nor U25739 (N_25739,N_25209,N_25069);
nand U25740 (N_25740,N_25333,N_25206);
and U25741 (N_25741,N_25211,N_25045);
nor U25742 (N_25742,N_25475,N_25118);
nor U25743 (N_25743,N_25055,N_25348);
nor U25744 (N_25744,N_25499,N_25327);
nor U25745 (N_25745,N_25406,N_25454);
nand U25746 (N_25746,N_25028,N_25422);
or U25747 (N_25747,N_25458,N_25145);
nor U25748 (N_25748,N_25106,N_25241);
nor U25749 (N_25749,N_25041,N_25049);
nor U25750 (N_25750,N_25174,N_25038);
or U25751 (N_25751,N_25398,N_25298);
or U25752 (N_25752,N_25274,N_25288);
nand U25753 (N_25753,N_25386,N_25068);
nor U25754 (N_25754,N_25336,N_25224);
and U25755 (N_25755,N_25272,N_25280);
or U25756 (N_25756,N_25119,N_25486);
or U25757 (N_25757,N_25366,N_25259);
and U25758 (N_25758,N_25479,N_25135);
or U25759 (N_25759,N_25409,N_25319);
and U25760 (N_25760,N_25415,N_25182);
and U25761 (N_25761,N_25083,N_25062);
or U25762 (N_25762,N_25007,N_25165);
nor U25763 (N_25763,N_25308,N_25180);
nor U25764 (N_25764,N_25055,N_25107);
nor U25765 (N_25765,N_25138,N_25273);
xor U25766 (N_25766,N_25295,N_25347);
nor U25767 (N_25767,N_25409,N_25091);
nor U25768 (N_25768,N_25344,N_25108);
or U25769 (N_25769,N_25367,N_25288);
or U25770 (N_25770,N_25441,N_25243);
or U25771 (N_25771,N_25084,N_25190);
and U25772 (N_25772,N_25051,N_25420);
nand U25773 (N_25773,N_25197,N_25386);
nor U25774 (N_25774,N_25279,N_25479);
or U25775 (N_25775,N_25319,N_25395);
nor U25776 (N_25776,N_25437,N_25220);
nor U25777 (N_25777,N_25281,N_25250);
nand U25778 (N_25778,N_25328,N_25090);
and U25779 (N_25779,N_25194,N_25390);
and U25780 (N_25780,N_25413,N_25058);
xnor U25781 (N_25781,N_25408,N_25318);
nand U25782 (N_25782,N_25046,N_25132);
nor U25783 (N_25783,N_25496,N_25146);
xnor U25784 (N_25784,N_25219,N_25485);
nor U25785 (N_25785,N_25406,N_25299);
and U25786 (N_25786,N_25497,N_25225);
and U25787 (N_25787,N_25218,N_25368);
nor U25788 (N_25788,N_25257,N_25064);
nand U25789 (N_25789,N_25088,N_25474);
xor U25790 (N_25790,N_25023,N_25229);
nor U25791 (N_25791,N_25414,N_25427);
or U25792 (N_25792,N_25056,N_25316);
or U25793 (N_25793,N_25237,N_25261);
nand U25794 (N_25794,N_25052,N_25028);
nand U25795 (N_25795,N_25360,N_25299);
nor U25796 (N_25796,N_25420,N_25091);
or U25797 (N_25797,N_25348,N_25134);
and U25798 (N_25798,N_25333,N_25411);
nor U25799 (N_25799,N_25067,N_25286);
nor U25800 (N_25800,N_25232,N_25436);
or U25801 (N_25801,N_25394,N_25387);
or U25802 (N_25802,N_25452,N_25006);
and U25803 (N_25803,N_25364,N_25008);
nand U25804 (N_25804,N_25171,N_25368);
nand U25805 (N_25805,N_25444,N_25371);
nand U25806 (N_25806,N_25010,N_25163);
or U25807 (N_25807,N_25307,N_25381);
nor U25808 (N_25808,N_25065,N_25062);
and U25809 (N_25809,N_25195,N_25125);
or U25810 (N_25810,N_25244,N_25480);
nor U25811 (N_25811,N_25058,N_25207);
nor U25812 (N_25812,N_25006,N_25054);
and U25813 (N_25813,N_25266,N_25299);
or U25814 (N_25814,N_25392,N_25396);
nor U25815 (N_25815,N_25013,N_25360);
and U25816 (N_25816,N_25257,N_25297);
nand U25817 (N_25817,N_25366,N_25292);
and U25818 (N_25818,N_25007,N_25231);
or U25819 (N_25819,N_25333,N_25176);
nand U25820 (N_25820,N_25249,N_25124);
and U25821 (N_25821,N_25326,N_25072);
nor U25822 (N_25822,N_25231,N_25432);
nor U25823 (N_25823,N_25306,N_25339);
nor U25824 (N_25824,N_25153,N_25342);
and U25825 (N_25825,N_25333,N_25227);
nor U25826 (N_25826,N_25464,N_25358);
nand U25827 (N_25827,N_25378,N_25485);
nor U25828 (N_25828,N_25448,N_25477);
and U25829 (N_25829,N_25335,N_25407);
and U25830 (N_25830,N_25214,N_25187);
xor U25831 (N_25831,N_25118,N_25113);
xnor U25832 (N_25832,N_25332,N_25318);
and U25833 (N_25833,N_25286,N_25272);
and U25834 (N_25834,N_25325,N_25036);
nand U25835 (N_25835,N_25076,N_25484);
nor U25836 (N_25836,N_25237,N_25063);
and U25837 (N_25837,N_25476,N_25342);
nand U25838 (N_25838,N_25302,N_25092);
nand U25839 (N_25839,N_25124,N_25105);
nor U25840 (N_25840,N_25063,N_25219);
xnor U25841 (N_25841,N_25007,N_25113);
or U25842 (N_25842,N_25109,N_25342);
nand U25843 (N_25843,N_25402,N_25198);
and U25844 (N_25844,N_25493,N_25202);
nand U25845 (N_25845,N_25162,N_25048);
nand U25846 (N_25846,N_25118,N_25447);
or U25847 (N_25847,N_25372,N_25398);
or U25848 (N_25848,N_25447,N_25078);
xnor U25849 (N_25849,N_25331,N_25489);
nor U25850 (N_25850,N_25032,N_25425);
and U25851 (N_25851,N_25282,N_25497);
nor U25852 (N_25852,N_25443,N_25034);
nor U25853 (N_25853,N_25446,N_25483);
xor U25854 (N_25854,N_25288,N_25013);
and U25855 (N_25855,N_25405,N_25472);
and U25856 (N_25856,N_25093,N_25452);
or U25857 (N_25857,N_25380,N_25376);
nand U25858 (N_25858,N_25431,N_25326);
or U25859 (N_25859,N_25000,N_25265);
nand U25860 (N_25860,N_25111,N_25415);
nor U25861 (N_25861,N_25349,N_25484);
and U25862 (N_25862,N_25282,N_25072);
and U25863 (N_25863,N_25370,N_25005);
nor U25864 (N_25864,N_25031,N_25365);
nor U25865 (N_25865,N_25206,N_25357);
and U25866 (N_25866,N_25494,N_25215);
and U25867 (N_25867,N_25056,N_25146);
and U25868 (N_25868,N_25422,N_25246);
nor U25869 (N_25869,N_25348,N_25156);
and U25870 (N_25870,N_25229,N_25413);
and U25871 (N_25871,N_25399,N_25480);
nand U25872 (N_25872,N_25059,N_25191);
nand U25873 (N_25873,N_25027,N_25101);
or U25874 (N_25874,N_25129,N_25083);
nor U25875 (N_25875,N_25374,N_25415);
nand U25876 (N_25876,N_25434,N_25269);
or U25877 (N_25877,N_25105,N_25157);
nor U25878 (N_25878,N_25343,N_25225);
nor U25879 (N_25879,N_25036,N_25472);
or U25880 (N_25880,N_25002,N_25407);
nor U25881 (N_25881,N_25316,N_25034);
nor U25882 (N_25882,N_25335,N_25290);
and U25883 (N_25883,N_25027,N_25463);
nand U25884 (N_25884,N_25474,N_25330);
and U25885 (N_25885,N_25401,N_25442);
nand U25886 (N_25886,N_25002,N_25272);
and U25887 (N_25887,N_25132,N_25451);
xor U25888 (N_25888,N_25431,N_25135);
and U25889 (N_25889,N_25438,N_25497);
xor U25890 (N_25890,N_25165,N_25259);
xnor U25891 (N_25891,N_25021,N_25444);
xnor U25892 (N_25892,N_25160,N_25422);
nor U25893 (N_25893,N_25007,N_25344);
and U25894 (N_25894,N_25297,N_25387);
or U25895 (N_25895,N_25137,N_25038);
nor U25896 (N_25896,N_25318,N_25228);
and U25897 (N_25897,N_25331,N_25101);
nand U25898 (N_25898,N_25450,N_25212);
and U25899 (N_25899,N_25126,N_25486);
nand U25900 (N_25900,N_25067,N_25298);
and U25901 (N_25901,N_25451,N_25163);
or U25902 (N_25902,N_25353,N_25263);
nand U25903 (N_25903,N_25459,N_25087);
nor U25904 (N_25904,N_25267,N_25295);
nor U25905 (N_25905,N_25393,N_25055);
xor U25906 (N_25906,N_25200,N_25462);
or U25907 (N_25907,N_25470,N_25362);
nand U25908 (N_25908,N_25403,N_25441);
nor U25909 (N_25909,N_25497,N_25044);
nor U25910 (N_25910,N_25014,N_25024);
and U25911 (N_25911,N_25023,N_25417);
or U25912 (N_25912,N_25200,N_25195);
or U25913 (N_25913,N_25237,N_25071);
nand U25914 (N_25914,N_25371,N_25476);
nand U25915 (N_25915,N_25342,N_25403);
nor U25916 (N_25916,N_25120,N_25245);
and U25917 (N_25917,N_25003,N_25447);
xor U25918 (N_25918,N_25330,N_25381);
and U25919 (N_25919,N_25167,N_25060);
nand U25920 (N_25920,N_25108,N_25232);
nor U25921 (N_25921,N_25282,N_25404);
nand U25922 (N_25922,N_25126,N_25010);
nor U25923 (N_25923,N_25232,N_25276);
xor U25924 (N_25924,N_25076,N_25464);
xnor U25925 (N_25925,N_25482,N_25384);
nor U25926 (N_25926,N_25409,N_25064);
or U25927 (N_25927,N_25315,N_25019);
or U25928 (N_25928,N_25446,N_25423);
xnor U25929 (N_25929,N_25376,N_25373);
nor U25930 (N_25930,N_25182,N_25129);
nand U25931 (N_25931,N_25479,N_25111);
nand U25932 (N_25932,N_25285,N_25046);
nor U25933 (N_25933,N_25156,N_25060);
or U25934 (N_25934,N_25479,N_25454);
nand U25935 (N_25935,N_25384,N_25490);
xor U25936 (N_25936,N_25381,N_25003);
and U25937 (N_25937,N_25432,N_25227);
or U25938 (N_25938,N_25428,N_25297);
nor U25939 (N_25939,N_25190,N_25153);
nor U25940 (N_25940,N_25372,N_25281);
xnor U25941 (N_25941,N_25046,N_25186);
or U25942 (N_25942,N_25319,N_25213);
nor U25943 (N_25943,N_25082,N_25335);
xor U25944 (N_25944,N_25126,N_25089);
or U25945 (N_25945,N_25241,N_25150);
nor U25946 (N_25946,N_25278,N_25317);
nand U25947 (N_25947,N_25361,N_25321);
or U25948 (N_25948,N_25386,N_25351);
nand U25949 (N_25949,N_25472,N_25039);
nand U25950 (N_25950,N_25359,N_25177);
xor U25951 (N_25951,N_25406,N_25466);
nor U25952 (N_25952,N_25223,N_25397);
nand U25953 (N_25953,N_25232,N_25105);
and U25954 (N_25954,N_25255,N_25139);
xor U25955 (N_25955,N_25120,N_25449);
xor U25956 (N_25956,N_25287,N_25033);
nand U25957 (N_25957,N_25336,N_25341);
or U25958 (N_25958,N_25442,N_25293);
nor U25959 (N_25959,N_25152,N_25294);
xnor U25960 (N_25960,N_25127,N_25425);
xor U25961 (N_25961,N_25445,N_25409);
and U25962 (N_25962,N_25155,N_25408);
or U25963 (N_25963,N_25215,N_25225);
nand U25964 (N_25964,N_25014,N_25418);
or U25965 (N_25965,N_25111,N_25468);
nor U25966 (N_25966,N_25010,N_25255);
or U25967 (N_25967,N_25108,N_25450);
or U25968 (N_25968,N_25014,N_25169);
nor U25969 (N_25969,N_25079,N_25005);
and U25970 (N_25970,N_25227,N_25204);
nand U25971 (N_25971,N_25026,N_25482);
nand U25972 (N_25972,N_25092,N_25448);
nand U25973 (N_25973,N_25154,N_25448);
nand U25974 (N_25974,N_25277,N_25025);
nand U25975 (N_25975,N_25202,N_25278);
or U25976 (N_25976,N_25379,N_25319);
or U25977 (N_25977,N_25202,N_25096);
or U25978 (N_25978,N_25356,N_25385);
nor U25979 (N_25979,N_25408,N_25131);
nor U25980 (N_25980,N_25168,N_25294);
nand U25981 (N_25981,N_25201,N_25052);
and U25982 (N_25982,N_25324,N_25131);
nor U25983 (N_25983,N_25370,N_25037);
and U25984 (N_25984,N_25084,N_25253);
and U25985 (N_25985,N_25206,N_25417);
nor U25986 (N_25986,N_25434,N_25327);
and U25987 (N_25987,N_25407,N_25079);
nor U25988 (N_25988,N_25020,N_25304);
and U25989 (N_25989,N_25311,N_25357);
or U25990 (N_25990,N_25052,N_25249);
or U25991 (N_25991,N_25485,N_25280);
nor U25992 (N_25992,N_25012,N_25186);
xor U25993 (N_25993,N_25281,N_25072);
nor U25994 (N_25994,N_25220,N_25004);
or U25995 (N_25995,N_25462,N_25019);
or U25996 (N_25996,N_25449,N_25417);
nor U25997 (N_25997,N_25245,N_25210);
nand U25998 (N_25998,N_25246,N_25050);
and U25999 (N_25999,N_25421,N_25478);
xor U26000 (N_26000,N_25950,N_25601);
and U26001 (N_26001,N_25704,N_25757);
nor U26002 (N_26002,N_25807,N_25958);
and U26003 (N_26003,N_25594,N_25901);
and U26004 (N_26004,N_25572,N_25888);
xor U26005 (N_26005,N_25504,N_25837);
xnor U26006 (N_26006,N_25624,N_25514);
and U26007 (N_26007,N_25649,N_25522);
nand U26008 (N_26008,N_25937,N_25894);
xor U26009 (N_26009,N_25538,N_25783);
nor U26010 (N_26010,N_25832,N_25710);
or U26011 (N_26011,N_25812,N_25596);
nand U26012 (N_26012,N_25665,N_25571);
and U26013 (N_26013,N_25718,N_25906);
or U26014 (N_26014,N_25819,N_25887);
xnor U26015 (N_26015,N_25520,N_25912);
nor U26016 (N_26016,N_25735,N_25761);
nor U26017 (N_26017,N_25661,N_25513);
or U26018 (N_26018,N_25968,N_25873);
or U26019 (N_26019,N_25676,N_25566);
nor U26020 (N_26020,N_25989,N_25565);
and U26021 (N_26021,N_25825,N_25568);
nor U26022 (N_26022,N_25729,N_25781);
nand U26023 (N_26023,N_25830,N_25821);
nor U26024 (N_26024,N_25780,N_25838);
nor U26025 (N_26025,N_25550,N_25778);
nor U26026 (N_26026,N_25715,N_25552);
and U26027 (N_26027,N_25553,N_25760);
or U26028 (N_26028,N_25848,N_25836);
nand U26029 (N_26029,N_25831,N_25699);
nand U26030 (N_26030,N_25633,N_25864);
nor U26031 (N_26031,N_25965,N_25856);
nor U26032 (N_26032,N_25608,N_25849);
and U26033 (N_26033,N_25586,N_25507);
or U26034 (N_26034,N_25839,N_25687);
or U26035 (N_26035,N_25771,N_25744);
nand U26036 (N_26036,N_25991,N_25853);
and U26037 (N_26037,N_25655,N_25891);
or U26038 (N_26038,N_25660,N_25510);
nand U26039 (N_26039,N_25820,N_25843);
or U26040 (N_26040,N_25647,N_25946);
nand U26041 (N_26041,N_25555,N_25706);
nor U26042 (N_26042,N_25897,N_25930);
nor U26043 (N_26043,N_25598,N_25896);
nand U26044 (N_26044,N_25716,N_25614);
nor U26045 (N_26045,N_25658,N_25548);
or U26046 (N_26046,N_25755,N_25707);
nor U26047 (N_26047,N_25768,N_25788);
and U26048 (N_26048,N_25573,N_25623);
nor U26049 (N_26049,N_25517,N_25993);
nand U26050 (N_26050,N_25717,N_25956);
and U26051 (N_26051,N_25728,N_25943);
or U26052 (N_26052,N_25875,N_25845);
nand U26053 (N_26053,N_25712,N_25521);
or U26054 (N_26054,N_25949,N_25703);
nand U26055 (N_26055,N_25722,N_25861);
and U26056 (N_26056,N_25952,N_25854);
or U26057 (N_26057,N_25595,N_25570);
xnor U26058 (N_26058,N_25635,N_25743);
xnor U26059 (N_26059,N_25732,N_25785);
and U26060 (N_26060,N_25876,N_25580);
nor U26061 (N_26061,N_25673,N_25597);
nand U26062 (N_26062,N_25809,N_25619);
and U26063 (N_26063,N_25721,N_25698);
nor U26064 (N_26064,N_25988,N_25840);
and U26065 (N_26065,N_25682,N_25858);
or U26066 (N_26066,N_25805,N_25563);
nor U26067 (N_26067,N_25525,N_25745);
nor U26068 (N_26068,N_25713,N_25724);
and U26069 (N_26069,N_25589,N_25671);
and U26070 (N_26070,N_25694,N_25680);
nand U26071 (N_26071,N_25947,N_25827);
and U26072 (N_26072,N_25777,N_25625);
nor U26073 (N_26073,N_25506,N_25651);
nand U26074 (N_26074,N_25791,N_25942);
and U26075 (N_26075,N_25591,N_25662);
and U26076 (N_26076,N_25786,N_25561);
nand U26077 (N_26077,N_25674,N_25762);
and U26078 (N_26078,N_25979,N_25905);
nand U26079 (N_26079,N_25871,N_25892);
nor U26080 (N_26080,N_25530,N_25746);
and U26081 (N_26081,N_25643,N_25650);
or U26082 (N_26082,N_25810,N_25515);
nor U26083 (N_26083,N_25971,N_25683);
or U26084 (N_26084,N_25939,N_25789);
nor U26085 (N_26085,N_25659,N_25535);
and U26086 (N_26086,N_25984,N_25799);
nand U26087 (N_26087,N_25636,N_25867);
or U26088 (N_26088,N_25857,N_25811);
nand U26089 (N_26089,N_25657,N_25737);
or U26090 (N_26090,N_25969,N_25907);
nand U26091 (N_26091,N_25954,N_25590);
nand U26092 (N_26092,N_25526,N_25924);
nor U26093 (N_26093,N_25641,N_25842);
and U26094 (N_26094,N_25536,N_25990);
and U26095 (N_26095,N_25938,N_25529);
and U26096 (N_26096,N_25828,N_25618);
nor U26097 (N_26097,N_25995,N_25932);
or U26098 (N_26098,N_25973,N_25759);
nand U26099 (N_26099,N_25739,N_25604);
nand U26100 (N_26100,N_25727,N_25544);
nor U26101 (N_26101,N_25584,N_25774);
nor U26102 (N_26102,N_25880,N_25941);
and U26103 (N_26103,N_25534,N_25927);
nand U26104 (N_26104,N_25546,N_25523);
nor U26105 (N_26105,N_25630,N_25962);
nor U26106 (N_26106,N_25773,N_25961);
or U26107 (N_26107,N_25846,N_25637);
or U26108 (N_26108,N_25667,N_25879);
nor U26109 (N_26109,N_25539,N_25669);
nand U26110 (N_26110,N_25602,N_25929);
nand U26111 (N_26111,N_25914,N_25654);
nor U26112 (N_26112,N_25626,N_25502);
nor U26113 (N_26113,N_25560,N_25516);
nor U26114 (N_26114,N_25859,N_25508);
xor U26115 (N_26115,N_25797,N_25889);
and U26116 (N_26116,N_25692,N_25668);
nor U26117 (N_26117,N_25751,N_25622);
and U26118 (N_26118,N_25653,N_25588);
xor U26119 (N_26119,N_25974,N_25642);
nand U26120 (N_26120,N_25690,N_25533);
nand U26121 (N_26121,N_25611,N_25801);
or U26122 (N_26122,N_25599,N_25558);
or U26123 (N_26123,N_25613,N_25579);
nor U26124 (N_26124,N_25562,N_25869);
or U26125 (N_26125,N_25955,N_25957);
nand U26126 (N_26126,N_25631,N_25987);
nand U26127 (N_26127,N_25933,N_25615);
and U26128 (N_26128,N_25612,N_25754);
nand U26129 (N_26129,N_25764,N_25640);
and U26130 (N_26130,N_25822,N_25769);
xor U26131 (N_26131,N_25996,N_25936);
nor U26132 (N_26132,N_25787,N_25926);
or U26133 (N_26133,N_25582,N_25977);
nor U26134 (N_26134,N_25567,N_25554);
or U26135 (N_26135,N_25531,N_25500);
and U26136 (N_26136,N_25731,N_25793);
or U26137 (N_26137,N_25679,N_25714);
and U26138 (N_26138,N_25920,N_25756);
nor U26139 (N_26139,N_25592,N_25511);
nor U26140 (N_26140,N_25855,N_25616);
nand U26141 (N_26141,N_25980,N_25577);
or U26142 (N_26142,N_25862,N_25772);
or U26143 (N_26143,N_25519,N_25639);
or U26144 (N_26144,N_25695,N_25620);
xor U26145 (N_26145,N_25986,N_25865);
and U26146 (N_26146,N_25847,N_25823);
and U26147 (N_26147,N_25833,N_25931);
nand U26148 (N_26148,N_25528,N_25734);
or U26149 (N_26149,N_25863,N_25542);
and U26150 (N_26150,N_25505,N_25678);
nor U26151 (N_26151,N_25998,N_25804);
and U26152 (N_26152,N_25899,N_25557);
xor U26153 (N_26153,N_25796,N_25709);
xnor U26154 (N_26154,N_25841,N_25587);
nand U26155 (N_26155,N_25644,N_25564);
nand U26156 (N_26156,N_25798,N_25617);
nand U26157 (N_26157,N_25559,N_25792);
or U26158 (N_26158,N_25917,N_25720);
and U26159 (N_26159,N_25909,N_25999);
nand U26160 (N_26160,N_25908,N_25736);
nor U26161 (N_26161,N_25829,N_25632);
and U26162 (N_26162,N_25697,N_25882);
nand U26163 (N_26163,N_25850,N_25681);
and U26164 (N_26164,N_25960,N_25688);
xor U26165 (N_26165,N_25913,N_25978);
nor U26166 (N_26166,N_25923,N_25878);
nor U26167 (N_26167,N_25868,N_25527);
xor U26168 (N_26168,N_25675,N_25652);
and U26169 (N_26169,N_25775,N_25748);
nand U26170 (N_26170,N_25782,N_25541);
or U26171 (N_26171,N_25994,N_25621);
nand U26172 (N_26172,N_25606,N_25663);
and U26173 (N_26173,N_25902,N_25686);
or U26174 (N_26174,N_25818,N_25648);
or U26175 (N_26175,N_25672,N_25767);
nor U26176 (N_26176,N_25593,N_25922);
nor U26177 (N_26177,N_25666,N_25967);
nand U26178 (N_26178,N_25696,N_25940);
and U26179 (N_26179,N_25629,N_25750);
or U26180 (N_26180,N_25609,N_25972);
or U26181 (N_26181,N_25963,N_25890);
and U26182 (N_26182,N_25503,N_25753);
or U26183 (N_26183,N_25951,N_25740);
nand U26184 (N_26184,N_25997,N_25711);
xnor U26185 (N_26185,N_25870,N_25705);
nor U26186 (N_26186,N_25701,N_25603);
or U26187 (N_26187,N_25860,N_25900);
or U26188 (N_26188,N_25928,N_25547);
nand U26189 (N_26189,N_25708,N_25685);
nor U26190 (N_26190,N_25851,N_25985);
or U26191 (N_26191,N_25852,N_25747);
or U26192 (N_26192,N_25816,N_25749);
xnor U26193 (N_26193,N_25815,N_25540);
xor U26194 (N_26194,N_25945,N_25719);
and U26195 (N_26195,N_25784,N_25903);
and U26196 (N_26196,N_25512,N_25970);
nand U26197 (N_26197,N_25600,N_25866);
or U26198 (N_26198,N_25574,N_25742);
nor U26199 (N_26199,N_25733,N_25808);
nor U26200 (N_26200,N_25532,N_25645);
or U26201 (N_26201,N_25585,N_25738);
xnor U26202 (N_26202,N_25677,N_25803);
xor U26203 (N_26203,N_25959,N_25814);
nor U26204 (N_26204,N_25779,N_25966);
and U26205 (N_26205,N_25537,N_25992);
nand U26206 (N_26206,N_25578,N_25964);
and U26207 (N_26207,N_25693,N_25730);
nor U26208 (N_26208,N_25607,N_25634);
nand U26209 (N_26209,N_25638,N_25551);
nor U26210 (N_26210,N_25885,N_25794);
nand U26211 (N_26211,N_25911,N_25915);
nand U26212 (N_26212,N_25543,N_25898);
and U26213 (N_26213,N_25881,N_25983);
nand U26214 (N_26214,N_25834,N_25509);
nor U26215 (N_26215,N_25916,N_25575);
or U26216 (N_26216,N_25576,N_25524);
or U26217 (N_26217,N_25776,N_25795);
nor U26218 (N_26218,N_25806,N_25884);
and U26219 (N_26219,N_25953,N_25723);
or U26220 (N_26220,N_25910,N_25790);
and U26221 (N_26221,N_25725,N_25765);
nor U26222 (N_26222,N_25689,N_25691);
nand U26223 (N_26223,N_25934,N_25944);
or U26224 (N_26224,N_25741,N_25770);
nor U26225 (N_26225,N_25918,N_25895);
nand U26226 (N_26226,N_25844,N_25904);
or U26227 (N_26227,N_25872,N_25817);
nor U26228 (N_26228,N_25700,N_25981);
nor U26229 (N_26229,N_25893,N_25569);
or U26230 (N_26230,N_25919,N_25766);
or U26231 (N_26231,N_25948,N_25501);
nor U26232 (N_26232,N_25763,N_25646);
or U26233 (N_26233,N_25752,N_25581);
or U26234 (N_26234,N_25583,N_25670);
or U26235 (N_26235,N_25556,N_25976);
nor U26236 (N_26236,N_25835,N_25684);
nand U26237 (N_26237,N_25726,N_25874);
and U26238 (N_26238,N_25925,N_25610);
nand U26239 (N_26239,N_25545,N_25656);
nor U26240 (N_26240,N_25877,N_25826);
nand U26241 (N_26241,N_25982,N_25627);
or U26242 (N_26242,N_25935,N_25802);
or U26243 (N_26243,N_25921,N_25702);
and U26244 (N_26244,N_25813,N_25628);
nor U26245 (N_26245,N_25518,N_25886);
nand U26246 (N_26246,N_25549,N_25800);
nor U26247 (N_26247,N_25664,N_25824);
nor U26248 (N_26248,N_25883,N_25605);
or U26249 (N_26249,N_25758,N_25975);
and U26250 (N_26250,N_25556,N_25660);
or U26251 (N_26251,N_25865,N_25813);
and U26252 (N_26252,N_25569,N_25571);
nand U26253 (N_26253,N_25850,N_25987);
xor U26254 (N_26254,N_25644,N_25562);
and U26255 (N_26255,N_25595,N_25545);
xor U26256 (N_26256,N_25510,N_25857);
nor U26257 (N_26257,N_25777,N_25964);
nor U26258 (N_26258,N_25887,N_25767);
nor U26259 (N_26259,N_25588,N_25629);
nor U26260 (N_26260,N_25665,N_25765);
nor U26261 (N_26261,N_25951,N_25881);
or U26262 (N_26262,N_25993,N_25678);
nor U26263 (N_26263,N_25992,N_25588);
nand U26264 (N_26264,N_25652,N_25934);
nand U26265 (N_26265,N_25631,N_25625);
and U26266 (N_26266,N_25861,N_25854);
and U26267 (N_26267,N_25550,N_25597);
or U26268 (N_26268,N_25875,N_25607);
or U26269 (N_26269,N_25945,N_25578);
and U26270 (N_26270,N_25880,N_25804);
or U26271 (N_26271,N_25603,N_25924);
and U26272 (N_26272,N_25526,N_25879);
or U26273 (N_26273,N_25998,N_25799);
or U26274 (N_26274,N_25998,N_25952);
and U26275 (N_26275,N_25565,N_25977);
xor U26276 (N_26276,N_25703,N_25622);
nand U26277 (N_26277,N_25560,N_25673);
or U26278 (N_26278,N_25709,N_25841);
nor U26279 (N_26279,N_25644,N_25748);
nor U26280 (N_26280,N_25644,N_25939);
or U26281 (N_26281,N_25740,N_25627);
or U26282 (N_26282,N_25711,N_25720);
nand U26283 (N_26283,N_25840,N_25850);
nor U26284 (N_26284,N_25823,N_25580);
and U26285 (N_26285,N_25712,N_25918);
nand U26286 (N_26286,N_25658,N_25759);
nand U26287 (N_26287,N_25955,N_25852);
or U26288 (N_26288,N_25735,N_25895);
and U26289 (N_26289,N_25579,N_25954);
nor U26290 (N_26290,N_25565,N_25870);
nor U26291 (N_26291,N_25798,N_25821);
nand U26292 (N_26292,N_25899,N_25838);
and U26293 (N_26293,N_25640,N_25784);
xor U26294 (N_26294,N_25532,N_25899);
nand U26295 (N_26295,N_25619,N_25932);
nor U26296 (N_26296,N_25624,N_25526);
nand U26297 (N_26297,N_25585,N_25659);
nand U26298 (N_26298,N_25852,N_25553);
nand U26299 (N_26299,N_25549,N_25780);
xor U26300 (N_26300,N_25928,N_25715);
nor U26301 (N_26301,N_25796,N_25525);
nor U26302 (N_26302,N_25565,N_25832);
nand U26303 (N_26303,N_25755,N_25997);
or U26304 (N_26304,N_25964,N_25539);
nor U26305 (N_26305,N_25880,N_25841);
or U26306 (N_26306,N_25816,N_25878);
xor U26307 (N_26307,N_25725,N_25561);
nand U26308 (N_26308,N_25876,N_25754);
or U26309 (N_26309,N_25956,N_25963);
and U26310 (N_26310,N_25799,N_25965);
or U26311 (N_26311,N_25884,N_25957);
xor U26312 (N_26312,N_25617,N_25500);
or U26313 (N_26313,N_25723,N_25839);
nand U26314 (N_26314,N_25686,N_25556);
nor U26315 (N_26315,N_25867,N_25970);
or U26316 (N_26316,N_25651,N_25971);
nor U26317 (N_26317,N_25580,N_25886);
nor U26318 (N_26318,N_25902,N_25674);
nor U26319 (N_26319,N_25889,N_25971);
or U26320 (N_26320,N_25749,N_25904);
nand U26321 (N_26321,N_25618,N_25598);
nand U26322 (N_26322,N_25619,N_25945);
or U26323 (N_26323,N_25777,N_25776);
and U26324 (N_26324,N_25753,N_25641);
nor U26325 (N_26325,N_25673,N_25508);
and U26326 (N_26326,N_25762,N_25689);
nand U26327 (N_26327,N_25897,N_25739);
and U26328 (N_26328,N_25961,N_25694);
nor U26329 (N_26329,N_25580,N_25724);
nand U26330 (N_26330,N_25596,N_25737);
nand U26331 (N_26331,N_25798,N_25551);
and U26332 (N_26332,N_25909,N_25822);
or U26333 (N_26333,N_25929,N_25893);
nor U26334 (N_26334,N_25894,N_25531);
xor U26335 (N_26335,N_25670,N_25986);
or U26336 (N_26336,N_25630,N_25515);
and U26337 (N_26337,N_25732,N_25789);
or U26338 (N_26338,N_25576,N_25694);
or U26339 (N_26339,N_25999,N_25527);
nand U26340 (N_26340,N_25689,N_25776);
nor U26341 (N_26341,N_25698,N_25526);
nor U26342 (N_26342,N_25894,N_25500);
nor U26343 (N_26343,N_25970,N_25728);
or U26344 (N_26344,N_25739,N_25699);
nor U26345 (N_26345,N_25719,N_25810);
nand U26346 (N_26346,N_25901,N_25726);
xor U26347 (N_26347,N_25576,N_25592);
nand U26348 (N_26348,N_25589,N_25718);
nor U26349 (N_26349,N_25650,N_25596);
and U26350 (N_26350,N_25960,N_25671);
and U26351 (N_26351,N_25932,N_25788);
xnor U26352 (N_26352,N_25646,N_25716);
nor U26353 (N_26353,N_25755,N_25958);
xor U26354 (N_26354,N_25556,N_25771);
nand U26355 (N_26355,N_25741,N_25979);
and U26356 (N_26356,N_25911,N_25872);
nor U26357 (N_26357,N_25846,N_25769);
nor U26358 (N_26358,N_25524,N_25756);
xnor U26359 (N_26359,N_25756,N_25638);
nand U26360 (N_26360,N_25635,N_25894);
nor U26361 (N_26361,N_25768,N_25914);
xor U26362 (N_26362,N_25923,N_25709);
and U26363 (N_26363,N_25555,N_25866);
or U26364 (N_26364,N_25924,N_25836);
nand U26365 (N_26365,N_25842,N_25618);
or U26366 (N_26366,N_25620,N_25595);
and U26367 (N_26367,N_25829,N_25861);
nand U26368 (N_26368,N_25686,N_25719);
nand U26369 (N_26369,N_25954,N_25690);
and U26370 (N_26370,N_25542,N_25664);
or U26371 (N_26371,N_25662,N_25949);
or U26372 (N_26372,N_25505,N_25823);
nor U26373 (N_26373,N_25755,N_25637);
nand U26374 (N_26374,N_25533,N_25604);
or U26375 (N_26375,N_25746,N_25659);
and U26376 (N_26376,N_25641,N_25988);
or U26377 (N_26377,N_25818,N_25761);
nand U26378 (N_26378,N_25516,N_25538);
nor U26379 (N_26379,N_25826,N_25674);
nor U26380 (N_26380,N_25821,N_25547);
nand U26381 (N_26381,N_25972,N_25735);
or U26382 (N_26382,N_25658,N_25983);
or U26383 (N_26383,N_25650,N_25667);
or U26384 (N_26384,N_25563,N_25554);
nand U26385 (N_26385,N_25902,N_25756);
nand U26386 (N_26386,N_25767,N_25859);
and U26387 (N_26387,N_25772,N_25689);
and U26388 (N_26388,N_25963,N_25806);
and U26389 (N_26389,N_25614,N_25521);
xnor U26390 (N_26390,N_25952,N_25631);
nand U26391 (N_26391,N_25544,N_25664);
or U26392 (N_26392,N_25697,N_25959);
nand U26393 (N_26393,N_25728,N_25924);
nor U26394 (N_26394,N_25758,N_25676);
nor U26395 (N_26395,N_25616,N_25868);
nand U26396 (N_26396,N_25750,N_25877);
nor U26397 (N_26397,N_25798,N_25714);
or U26398 (N_26398,N_25579,N_25698);
and U26399 (N_26399,N_25729,N_25861);
nand U26400 (N_26400,N_25762,N_25961);
and U26401 (N_26401,N_25596,N_25604);
or U26402 (N_26402,N_25825,N_25940);
nor U26403 (N_26403,N_25667,N_25516);
nand U26404 (N_26404,N_25639,N_25638);
or U26405 (N_26405,N_25983,N_25542);
and U26406 (N_26406,N_25587,N_25885);
and U26407 (N_26407,N_25937,N_25658);
nand U26408 (N_26408,N_25919,N_25768);
and U26409 (N_26409,N_25673,N_25810);
nor U26410 (N_26410,N_25787,N_25577);
nor U26411 (N_26411,N_25633,N_25609);
nand U26412 (N_26412,N_25654,N_25750);
xor U26413 (N_26413,N_25575,N_25735);
or U26414 (N_26414,N_25712,N_25628);
xor U26415 (N_26415,N_25584,N_25687);
nor U26416 (N_26416,N_25856,N_25559);
xor U26417 (N_26417,N_25775,N_25989);
xor U26418 (N_26418,N_25955,N_25630);
nand U26419 (N_26419,N_25738,N_25535);
nand U26420 (N_26420,N_25765,N_25987);
nor U26421 (N_26421,N_25829,N_25824);
xor U26422 (N_26422,N_25579,N_25743);
nor U26423 (N_26423,N_25736,N_25900);
or U26424 (N_26424,N_25794,N_25511);
nor U26425 (N_26425,N_25554,N_25600);
and U26426 (N_26426,N_25940,N_25911);
nand U26427 (N_26427,N_25880,N_25548);
and U26428 (N_26428,N_25526,N_25911);
nand U26429 (N_26429,N_25979,N_25587);
and U26430 (N_26430,N_25854,N_25608);
nand U26431 (N_26431,N_25826,N_25800);
nor U26432 (N_26432,N_25716,N_25872);
and U26433 (N_26433,N_25652,N_25709);
nor U26434 (N_26434,N_25615,N_25717);
nor U26435 (N_26435,N_25943,N_25989);
xor U26436 (N_26436,N_25813,N_25994);
nand U26437 (N_26437,N_25506,N_25698);
nand U26438 (N_26438,N_25892,N_25941);
nand U26439 (N_26439,N_25828,N_25670);
nor U26440 (N_26440,N_25616,N_25728);
nor U26441 (N_26441,N_25525,N_25921);
and U26442 (N_26442,N_25702,N_25904);
or U26443 (N_26443,N_25865,N_25529);
nand U26444 (N_26444,N_25704,N_25666);
xor U26445 (N_26445,N_25899,N_25661);
nor U26446 (N_26446,N_25976,N_25620);
nor U26447 (N_26447,N_25667,N_25570);
or U26448 (N_26448,N_25818,N_25763);
and U26449 (N_26449,N_25847,N_25738);
xnor U26450 (N_26450,N_25788,N_25786);
nor U26451 (N_26451,N_25938,N_25620);
xor U26452 (N_26452,N_25744,N_25665);
xor U26453 (N_26453,N_25566,N_25614);
nand U26454 (N_26454,N_25755,N_25539);
and U26455 (N_26455,N_25922,N_25664);
nor U26456 (N_26456,N_25575,N_25645);
nor U26457 (N_26457,N_25905,N_25725);
or U26458 (N_26458,N_25585,N_25993);
nand U26459 (N_26459,N_25607,N_25891);
and U26460 (N_26460,N_25743,N_25659);
and U26461 (N_26461,N_25507,N_25650);
and U26462 (N_26462,N_25633,N_25825);
nand U26463 (N_26463,N_25838,N_25776);
nand U26464 (N_26464,N_25626,N_25547);
xnor U26465 (N_26465,N_25663,N_25956);
nor U26466 (N_26466,N_25571,N_25559);
or U26467 (N_26467,N_25578,N_25705);
nand U26468 (N_26468,N_25994,N_25761);
or U26469 (N_26469,N_25871,N_25579);
and U26470 (N_26470,N_25559,N_25619);
or U26471 (N_26471,N_25531,N_25795);
and U26472 (N_26472,N_25850,N_25814);
xor U26473 (N_26473,N_25727,N_25704);
and U26474 (N_26474,N_25765,N_25914);
and U26475 (N_26475,N_25753,N_25565);
or U26476 (N_26476,N_25687,N_25887);
and U26477 (N_26477,N_25509,N_25634);
nor U26478 (N_26478,N_25756,N_25583);
nand U26479 (N_26479,N_25917,N_25999);
and U26480 (N_26480,N_25796,N_25613);
or U26481 (N_26481,N_25898,N_25696);
nor U26482 (N_26482,N_25655,N_25574);
or U26483 (N_26483,N_25800,N_25512);
and U26484 (N_26484,N_25502,N_25852);
nor U26485 (N_26485,N_25698,N_25754);
or U26486 (N_26486,N_25788,N_25836);
nand U26487 (N_26487,N_25889,N_25781);
nand U26488 (N_26488,N_25705,N_25846);
or U26489 (N_26489,N_25647,N_25863);
nand U26490 (N_26490,N_25886,N_25857);
nand U26491 (N_26491,N_25959,N_25896);
nor U26492 (N_26492,N_25693,N_25970);
and U26493 (N_26493,N_25555,N_25558);
and U26494 (N_26494,N_25797,N_25591);
and U26495 (N_26495,N_25611,N_25871);
nand U26496 (N_26496,N_25891,N_25976);
nand U26497 (N_26497,N_25723,N_25594);
or U26498 (N_26498,N_25847,N_25599);
or U26499 (N_26499,N_25748,N_25736);
nand U26500 (N_26500,N_26438,N_26381);
or U26501 (N_26501,N_26152,N_26209);
nor U26502 (N_26502,N_26356,N_26490);
and U26503 (N_26503,N_26178,N_26095);
xor U26504 (N_26504,N_26293,N_26359);
nand U26505 (N_26505,N_26116,N_26074);
xor U26506 (N_26506,N_26051,N_26472);
nor U26507 (N_26507,N_26377,N_26428);
and U26508 (N_26508,N_26370,N_26418);
nand U26509 (N_26509,N_26189,N_26460);
nand U26510 (N_26510,N_26055,N_26140);
and U26511 (N_26511,N_26279,N_26271);
xor U26512 (N_26512,N_26027,N_26410);
nor U26513 (N_26513,N_26196,N_26379);
and U26514 (N_26514,N_26324,N_26194);
nand U26515 (N_26515,N_26469,N_26394);
nand U26516 (N_26516,N_26232,N_26492);
or U26517 (N_26517,N_26338,N_26243);
nor U26518 (N_26518,N_26372,N_26415);
nand U26519 (N_26519,N_26302,N_26175);
nor U26520 (N_26520,N_26070,N_26367);
nor U26521 (N_26521,N_26488,N_26192);
and U26522 (N_26522,N_26396,N_26177);
and U26523 (N_26523,N_26364,N_26383);
nand U26524 (N_26524,N_26464,N_26273);
xor U26525 (N_26525,N_26165,N_26064);
or U26526 (N_26526,N_26053,N_26373);
xor U26527 (N_26527,N_26242,N_26229);
nand U26528 (N_26528,N_26183,N_26404);
nor U26529 (N_26529,N_26130,N_26000);
xnor U26530 (N_26530,N_26199,N_26421);
or U26531 (N_26531,N_26061,N_26172);
or U26532 (N_26532,N_26223,N_26049);
nand U26533 (N_26533,N_26202,N_26007);
nor U26534 (N_26534,N_26237,N_26250);
or U26535 (N_26535,N_26352,N_26230);
nor U26536 (N_26536,N_26327,N_26354);
and U26537 (N_26537,N_26092,N_26119);
nand U26538 (N_26538,N_26045,N_26337);
or U26539 (N_26539,N_26440,N_26283);
or U26540 (N_26540,N_26125,N_26066);
nand U26541 (N_26541,N_26282,N_26032);
nand U26542 (N_26542,N_26360,N_26059);
and U26543 (N_26543,N_26076,N_26176);
xnor U26544 (N_26544,N_26269,N_26082);
nand U26545 (N_26545,N_26117,N_26395);
xnor U26546 (N_26546,N_26482,N_26047);
nand U26547 (N_26547,N_26301,N_26445);
and U26548 (N_26548,N_26328,N_26320);
nor U26549 (N_26549,N_26434,N_26067);
nor U26550 (N_26550,N_26086,N_26365);
nand U26551 (N_26551,N_26128,N_26406);
and U26552 (N_26552,N_26288,N_26080);
or U26553 (N_26553,N_26499,N_26110);
and U26554 (N_26554,N_26233,N_26161);
xor U26555 (N_26555,N_26310,N_26275);
nand U26556 (N_26556,N_26257,N_26323);
nor U26557 (N_26557,N_26446,N_26393);
xnor U26558 (N_26558,N_26171,N_26050);
or U26559 (N_26559,N_26039,N_26433);
nor U26560 (N_26560,N_26432,N_26091);
or U26561 (N_26561,N_26435,N_26498);
nor U26562 (N_26562,N_26309,N_26225);
nor U26563 (N_26563,N_26124,N_26217);
xnor U26564 (N_26564,N_26109,N_26481);
nor U26565 (N_26565,N_26495,N_26292);
or U26566 (N_26566,N_26258,N_26284);
xor U26567 (N_26567,N_26035,N_26038);
and U26568 (N_26568,N_26376,N_26078);
or U26569 (N_26569,N_26397,N_26113);
or U26570 (N_26570,N_26062,N_26439);
xor U26571 (N_26571,N_26190,N_26368);
or U26572 (N_26572,N_26238,N_26017);
xor U26573 (N_26573,N_26147,N_26148);
and U26574 (N_26574,N_26494,N_26090);
or U26575 (N_26575,N_26259,N_26249);
and U26576 (N_26576,N_26387,N_26380);
nor U26577 (N_26577,N_26025,N_26414);
and U26578 (N_26578,N_26371,N_26105);
or U26579 (N_26579,N_26036,N_26164);
and U26580 (N_26580,N_26193,N_26458);
or U26581 (N_26581,N_26350,N_26306);
nand U26582 (N_26582,N_26332,N_26448);
nand U26583 (N_26583,N_26334,N_26197);
nand U26584 (N_26584,N_26023,N_26089);
and U26585 (N_26585,N_26112,N_26386);
or U26586 (N_26586,N_26083,N_26281);
or U26587 (N_26587,N_26041,N_26043);
or U26588 (N_26588,N_26211,N_26142);
xnor U26589 (N_26589,N_26162,N_26447);
nand U26590 (N_26590,N_26305,N_26361);
or U26591 (N_26591,N_26134,N_26491);
xor U26592 (N_26592,N_26444,N_26342);
nand U26593 (N_26593,N_26436,N_26056);
or U26594 (N_26594,N_26253,N_26442);
xor U26595 (N_26595,N_26160,N_26493);
nand U26596 (N_26596,N_26236,N_26026);
or U26597 (N_26597,N_26069,N_26318);
or U26598 (N_26598,N_26263,N_26475);
nor U26599 (N_26599,N_26001,N_26188);
xnor U26600 (N_26600,N_26011,N_26181);
nor U26601 (N_26601,N_26419,N_26412);
and U26602 (N_26602,N_26473,N_26215);
xnor U26603 (N_26603,N_26075,N_26248);
or U26604 (N_26604,N_26405,N_26042);
nand U26605 (N_26605,N_26022,N_26052);
xor U26606 (N_26606,N_26030,N_26009);
and U26607 (N_26607,N_26099,N_26144);
and U26608 (N_26608,N_26173,N_26307);
or U26609 (N_26609,N_26348,N_26463);
nand U26610 (N_26610,N_26311,N_26330);
xnor U26611 (N_26611,N_26487,N_26417);
and U26612 (N_26612,N_26468,N_26382);
and U26613 (N_26613,N_26201,N_26212);
xor U26614 (N_26614,N_26431,N_26347);
nor U26615 (N_26615,N_26168,N_26443);
nand U26616 (N_26616,N_26261,N_26103);
nand U26617 (N_26617,N_26020,N_26040);
xnor U26618 (N_26618,N_26264,N_26118);
nand U26619 (N_26619,N_26024,N_26300);
nand U26620 (N_26620,N_26422,N_26384);
or U26621 (N_26621,N_26018,N_26340);
or U26622 (N_26622,N_26329,N_26298);
nand U26623 (N_26623,N_26010,N_26313);
nand U26624 (N_26624,N_26466,N_26156);
nand U26625 (N_26625,N_26085,N_26423);
or U26626 (N_26626,N_26150,N_26013);
and U26627 (N_26627,N_26451,N_26133);
nor U26628 (N_26628,N_26402,N_26325);
or U26629 (N_26629,N_26467,N_26299);
xor U26630 (N_26630,N_26274,N_26399);
and U26631 (N_26631,N_26121,N_26063);
nand U26632 (N_26632,N_26002,N_26449);
nor U26633 (N_26633,N_26339,N_26483);
nand U26634 (N_26634,N_26278,N_26268);
or U26635 (N_26635,N_26145,N_26304);
or U26636 (N_26636,N_26478,N_26403);
xor U26637 (N_26637,N_26138,N_26077);
nor U26638 (N_26638,N_26094,N_26108);
nand U26639 (N_26639,N_26441,N_26005);
nor U26640 (N_26640,N_26126,N_26480);
and U26641 (N_26641,N_26459,N_26272);
or U26642 (N_26642,N_26413,N_26155);
or U26643 (N_26643,N_26252,N_26336);
nand U26644 (N_26644,N_26097,N_26220);
and U26645 (N_26645,N_26004,N_26407);
or U26646 (N_26646,N_26425,N_26398);
nand U26647 (N_26647,N_26191,N_26222);
nand U26648 (N_26648,N_26270,N_26186);
or U26649 (N_26649,N_26411,N_26021);
nor U26650 (N_26650,N_26245,N_26149);
nor U26651 (N_26651,N_26401,N_26450);
nand U26652 (N_26652,N_26187,N_26241);
nor U26653 (N_26653,N_26048,N_26213);
xor U26654 (N_26654,N_26346,N_26184);
and U26655 (N_26655,N_26331,N_26060);
or U26656 (N_26656,N_26366,N_26294);
or U26657 (N_26657,N_26219,N_26426);
or U26658 (N_26658,N_26221,N_26104);
or U26659 (N_26659,N_26014,N_26317);
nand U26660 (N_26660,N_26079,N_26054);
or U26661 (N_26661,N_26476,N_26461);
nor U26662 (N_26662,N_26295,N_26343);
or U26663 (N_26663,N_26102,N_26456);
xor U26664 (N_26664,N_26256,N_26058);
or U26665 (N_26665,N_26037,N_26231);
or U26666 (N_26666,N_26391,N_26003);
and U26667 (N_26667,N_26319,N_26132);
or U26668 (N_26668,N_26345,N_26267);
nand U26669 (N_26669,N_26170,N_26424);
nor U26670 (N_26670,N_26206,N_26087);
nor U26671 (N_26671,N_26057,N_26321);
nor U26672 (N_26672,N_26214,N_26088);
xor U26673 (N_26673,N_26137,N_26335);
nor U26674 (N_26674,N_26163,N_26470);
and U26675 (N_26675,N_26107,N_26008);
or U26676 (N_26676,N_26120,N_26114);
or U26677 (N_26677,N_26374,N_26157);
or U26678 (N_26678,N_26166,N_26277);
or U26679 (N_26679,N_26357,N_26111);
nand U26680 (N_26680,N_26247,N_26068);
and U26681 (N_26681,N_26169,N_26135);
nor U26682 (N_26682,N_26228,N_26390);
and U26683 (N_26683,N_26081,N_26158);
and U26684 (N_26684,N_26378,N_26203);
or U26685 (N_26685,N_26489,N_26098);
xnor U26686 (N_26686,N_26392,N_26101);
or U26687 (N_26687,N_26455,N_26484);
nand U26688 (N_26688,N_26012,N_26028);
and U26689 (N_26689,N_26180,N_26251);
nor U26690 (N_26690,N_26362,N_26216);
nand U26691 (N_26691,N_26084,N_26474);
nor U26692 (N_26692,N_26006,N_26314);
xor U26693 (N_26693,N_26122,N_26333);
or U26694 (N_26694,N_26266,N_26308);
nand U26695 (N_26695,N_26131,N_26303);
nor U26696 (N_26696,N_26254,N_26200);
and U26697 (N_26697,N_26019,N_26453);
nor U26698 (N_26698,N_26287,N_26141);
nand U26699 (N_26699,N_26355,N_26143);
or U26700 (N_26700,N_26351,N_26179);
or U26701 (N_26701,N_26388,N_26286);
nand U26702 (N_26702,N_26234,N_26115);
nand U26703 (N_26703,N_26218,N_26239);
or U26704 (N_26704,N_26205,N_26073);
and U26705 (N_26705,N_26151,N_26016);
and U26706 (N_26706,N_26358,N_26198);
and U26707 (N_26707,N_26457,N_26235);
or U26708 (N_26708,N_26315,N_26265);
nand U26709 (N_26709,N_26207,N_26290);
or U26710 (N_26710,N_26465,N_26071);
or U26711 (N_26711,N_26430,N_26400);
or U26712 (N_26712,N_26437,N_26363);
and U26713 (N_26713,N_26389,N_26224);
nor U26714 (N_26714,N_26153,N_26262);
and U26715 (N_26715,N_26260,N_26296);
nor U26716 (N_26716,N_26497,N_26429);
nor U26717 (N_26717,N_26033,N_26195);
nor U26718 (N_26718,N_26154,N_26454);
nor U26719 (N_26719,N_26322,N_26353);
or U26720 (N_26720,N_26065,N_26280);
or U26721 (N_26721,N_26167,N_26129);
nand U26722 (N_26722,N_26244,N_26486);
nor U26723 (N_26723,N_26208,N_26093);
or U26724 (N_26724,N_26369,N_26204);
xnor U26725 (N_26725,N_26246,N_26072);
nand U26726 (N_26726,N_26159,N_26210);
or U26727 (N_26727,N_26136,N_26471);
nor U26728 (N_26728,N_26015,N_26185);
nor U26729 (N_26729,N_26349,N_26316);
nand U26730 (N_26730,N_26291,N_26485);
nor U26731 (N_26731,N_26375,N_26255);
nor U26732 (N_26732,N_26409,N_26139);
and U26733 (N_26733,N_26408,N_26416);
or U26734 (N_26734,N_26031,N_26127);
xnor U26735 (N_26735,N_26044,N_26462);
nand U26736 (N_26736,N_26452,N_26289);
nand U26737 (N_26737,N_26427,N_26496);
nor U26738 (N_26738,N_26326,N_26100);
and U26739 (N_26739,N_26034,N_26312);
nor U26740 (N_26740,N_26146,N_26341);
nand U26741 (N_26741,N_26227,N_26477);
nor U26742 (N_26742,N_26297,N_26106);
and U26743 (N_26743,N_26479,N_26096);
or U26744 (N_26744,N_26182,N_26123);
nor U26745 (N_26745,N_26385,N_26029);
nor U26746 (N_26746,N_26420,N_26240);
xnor U26747 (N_26747,N_26046,N_26174);
and U26748 (N_26748,N_26285,N_26276);
nand U26749 (N_26749,N_26344,N_26226);
and U26750 (N_26750,N_26274,N_26160);
or U26751 (N_26751,N_26156,N_26062);
xor U26752 (N_26752,N_26282,N_26382);
nand U26753 (N_26753,N_26120,N_26002);
nand U26754 (N_26754,N_26337,N_26283);
or U26755 (N_26755,N_26289,N_26366);
nor U26756 (N_26756,N_26190,N_26211);
nand U26757 (N_26757,N_26014,N_26374);
nor U26758 (N_26758,N_26251,N_26182);
and U26759 (N_26759,N_26258,N_26042);
or U26760 (N_26760,N_26439,N_26107);
and U26761 (N_26761,N_26003,N_26345);
nor U26762 (N_26762,N_26029,N_26051);
and U26763 (N_26763,N_26037,N_26286);
and U26764 (N_26764,N_26473,N_26272);
nor U26765 (N_26765,N_26142,N_26168);
xnor U26766 (N_26766,N_26083,N_26300);
xnor U26767 (N_26767,N_26105,N_26223);
xnor U26768 (N_26768,N_26488,N_26072);
nand U26769 (N_26769,N_26143,N_26412);
nor U26770 (N_26770,N_26280,N_26117);
or U26771 (N_26771,N_26078,N_26217);
and U26772 (N_26772,N_26253,N_26469);
nand U26773 (N_26773,N_26343,N_26271);
nor U26774 (N_26774,N_26016,N_26076);
nand U26775 (N_26775,N_26392,N_26439);
nand U26776 (N_26776,N_26003,N_26362);
or U26777 (N_26777,N_26078,N_26008);
nor U26778 (N_26778,N_26239,N_26412);
and U26779 (N_26779,N_26052,N_26254);
or U26780 (N_26780,N_26220,N_26223);
nor U26781 (N_26781,N_26260,N_26367);
nand U26782 (N_26782,N_26144,N_26020);
nor U26783 (N_26783,N_26160,N_26286);
or U26784 (N_26784,N_26423,N_26153);
and U26785 (N_26785,N_26303,N_26302);
nand U26786 (N_26786,N_26251,N_26216);
nand U26787 (N_26787,N_26175,N_26345);
nor U26788 (N_26788,N_26017,N_26079);
or U26789 (N_26789,N_26114,N_26487);
or U26790 (N_26790,N_26137,N_26383);
or U26791 (N_26791,N_26245,N_26126);
nor U26792 (N_26792,N_26111,N_26478);
nor U26793 (N_26793,N_26128,N_26125);
nand U26794 (N_26794,N_26056,N_26026);
or U26795 (N_26795,N_26111,N_26459);
nor U26796 (N_26796,N_26465,N_26167);
or U26797 (N_26797,N_26153,N_26394);
xnor U26798 (N_26798,N_26482,N_26196);
and U26799 (N_26799,N_26088,N_26377);
nor U26800 (N_26800,N_26238,N_26413);
nand U26801 (N_26801,N_26450,N_26370);
or U26802 (N_26802,N_26164,N_26279);
or U26803 (N_26803,N_26479,N_26157);
nand U26804 (N_26804,N_26240,N_26245);
or U26805 (N_26805,N_26033,N_26285);
nand U26806 (N_26806,N_26395,N_26196);
or U26807 (N_26807,N_26402,N_26366);
and U26808 (N_26808,N_26439,N_26153);
nor U26809 (N_26809,N_26274,N_26191);
or U26810 (N_26810,N_26161,N_26166);
nor U26811 (N_26811,N_26381,N_26133);
and U26812 (N_26812,N_26405,N_26039);
xnor U26813 (N_26813,N_26399,N_26454);
nor U26814 (N_26814,N_26183,N_26153);
and U26815 (N_26815,N_26472,N_26429);
nand U26816 (N_26816,N_26049,N_26150);
or U26817 (N_26817,N_26497,N_26111);
and U26818 (N_26818,N_26442,N_26004);
nand U26819 (N_26819,N_26490,N_26075);
and U26820 (N_26820,N_26119,N_26445);
and U26821 (N_26821,N_26075,N_26346);
nor U26822 (N_26822,N_26450,N_26458);
or U26823 (N_26823,N_26078,N_26106);
nor U26824 (N_26824,N_26259,N_26484);
nand U26825 (N_26825,N_26161,N_26110);
xnor U26826 (N_26826,N_26026,N_26085);
xor U26827 (N_26827,N_26300,N_26234);
nand U26828 (N_26828,N_26064,N_26040);
nor U26829 (N_26829,N_26431,N_26174);
and U26830 (N_26830,N_26487,N_26415);
nand U26831 (N_26831,N_26091,N_26273);
and U26832 (N_26832,N_26037,N_26297);
nor U26833 (N_26833,N_26187,N_26087);
nor U26834 (N_26834,N_26388,N_26438);
xor U26835 (N_26835,N_26357,N_26360);
nand U26836 (N_26836,N_26361,N_26067);
or U26837 (N_26837,N_26337,N_26404);
and U26838 (N_26838,N_26401,N_26150);
nor U26839 (N_26839,N_26137,N_26450);
or U26840 (N_26840,N_26231,N_26476);
or U26841 (N_26841,N_26442,N_26002);
nand U26842 (N_26842,N_26061,N_26427);
or U26843 (N_26843,N_26369,N_26043);
or U26844 (N_26844,N_26491,N_26208);
xnor U26845 (N_26845,N_26062,N_26354);
and U26846 (N_26846,N_26317,N_26304);
nor U26847 (N_26847,N_26432,N_26177);
nor U26848 (N_26848,N_26448,N_26214);
nor U26849 (N_26849,N_26108,N_26277);
or U26850 (N_26850,N_26010,N_26150);
xnor U26851 (N_26851,N_26123,N_26030);
nand U26852 (N_26852,N_26013,N_26035);
nand U26853 (N_26853,N_26486,N_26324);
or U26854 (N_26854,N_26292,N_26483);
and U26855 (N_26855,N_26033,N_26342);
or U26856 (N_26856,N_26414,N_26008);
or U26857 (N_26857,N_26053,N_26107);
or U26858 (N_26858,N_26454,N_26278);
or U26859 (N_26859,N_26097,N_26172);
and U26860 (N_26860,N_26395,N_26097);
and U26861 (N_26861,N_26415,N_26208);
or U26862 (N_26862,N_26196,N_26107);
or U26863 (N_26863,N_26470,N_26246);
xor U26864 (N_26864,N_26088,N_26023);
nand U26865 (N_26865,N_26340,N_26182);
nand U26866 (N_26866,N_26306,N_26347);
or U26867 (N_26867,N_26213,N_26185);
nand U26868 (N_26868,N_26276,N_26242);
nand U26869 (N_26869,N_26162,N_26337);
nor U26870 (N_26870,N_26427,N_26497);
nor U26871 (N_26871,N_26266,N_26439);
and U26872 (N_26872,N_26105,N_26006);
nor U26873 (N_26873,N_26223,N_26110);
xor U26874 (N_26874,N_26081,N_26041);
nor U26875 (N_26875,N_26455,N_26155);
or U26876 (N_26876,N_26106,N_26308);
and U26877 (N_26877,N_26143,N_26469);
nor U26878 (N_26878,N_26386,N_26117);
and U26879 (N_26879,N_26378,N_26491);
nand U26880 (N_26880,N_26213,N_26178);
nor U26881 (N_26881,N_26320,N_26071);
and U26882 (N_26882,N_26266,N_26132);
nor U26883 (N_26883,N_26084,N_26368);
nor U26884 (N_26884,N_26179,N_26054);
nand U26885 (N_26885,N_26310,N_26182);
nor U26886 (N_26886,N_26071,N_26208);
nor U26887 (N_26887,N_26216,N_26458);
or U26888 (N_26888,N_26115,N_26421);
nor U26889 (N_26889,N_26358,N_26417);
or U26890 (N_26890,N_26326,N_26243);
or U26891 (N_26891,N_26325,N_26433);
xnor U26892 (N_26892,N_26072,N_26384);
or U26893 (N_26893,N_26317,N_26160);
nand U26894 (N_26894,N_26442,N_26224);
and U26895 (N_26895,N_26380,N_26081);
nor U26896 (N_26896,N_26346,N_26073);
nor U26897 (N_26897,N_26124,N_26130);
nand U26898 (N_26898,N_26363,N_26399);
nor U26899 (N_26899,N_26039,N_26078);
nand U26900 (N_26900,N_26428,N_26307);
and U26901 (N_26901,N_26331,N_26100);
or U26902 (N_26902,N_26086,N_26091);
and U26903 (N_26903,N_26499,N_26282);
or U26904 (N_26904,N_26278,N_26361);
or U26905 (N_26905,N_26203,N_26388);
nand U26906 (N_26906,N_26186,N_26311);
nand U26907 (N_26907,N_26176,N_26300);
or U26908 (N_26908,N_26134,N_26117);
nand U26909 (N_26909,N_26002,N_26249);
and U26910 (N_26910,N_26157,N_26139);
or U26911 (N_26911,N_26491,N_26273);
nand U26912 (N_26912,N_26053,N_26012);
xor U26913 (N_26913,N_26044,N_26435);
nand U26914 (N_26914,N_26051,N_26073);
nand U26915 (N_26915,N_26169,N_26424);
nor U26916 (N_26916,N_26460,N_26391);
or U26917 (N_26917,N_26478,N_26194);
or U26918 (N_26918,N_26496,N_26399);
nor U26919 (N_26919,N_26114,N_26149);
xor U26920 (N_26920,N_26322,N_26015);
or U26921 (N_26921,N_26392,N_26038);
nor U26922 (N_26922,N_26390,N_26167);
nand U26923 (N_26923,N_26006,N_26019);
nor U26924 (N_26924,N_26281,N_26323);
nand U26925 (N_26925,N_26410,N_26439);
nand U26926 (N_26926,N_26144,N_26286);
nand U26927 (N_26927,N_26007,N_26219);
nor U26928 (N_26928,N_26158,N_26113);
nor U26929 (N_26929,N_26167,N_26162);
and U26930 (N_26930,N_26397,N_26053);
nor U26931 (N_26931,N_26450,N_26274);
nand U26932 (N_26932,N_26077,N_26335);
nand U26933 (N_26933,N_26297,N_26381);
xor U26934 (N_26934,N_26014,N_26230);
nor U26935 (N_26935,N_26308,N_26136);
and U26936 (N_26936,N_26093,N_26173);
nand U26937 (N_26937,N_26488,N_26325);
and U26938 (N_26938,N_26001,N_26021);
nand U26939 (N_26939,N_26354,N_26060);
or U26940 (N_26940,N_26253,N_26214);
xnor U26941 (N_26941,N_26138,N_26143);
nand U26942 (N_26942,N_26129,N_26060);
and U26943 (N_26943,N_26146,N_26070);
or U26944 (N_26944,N_26174,N_26410);
xnor U26945 (N_26945,N_26156,N_26234);
or U26946 (N_26946,N_26480,N_26288);
nand U26947 (N_26947,N_26191,N_26195);
nor U26948 (N_26948,N_26240,N_26255);
nand U26949 (N_26949,N_26401,N_26030);
and U26950 (N_26950,N_26272,N_26339);
nor U26951 (N_26951,N_26007,N_26308);
xor U26952 (N_26952,N_26389,N_26268);
or U26953 (N_26953,N_26237,N_26267);
and U26954 (N_26954,N_26329,N_26049);
nor U26955 (N_26955,N_26403,N_26241);
and U26956 (N_26956,N_26171,N_26045);
nor U26957 (N_26957,N_26182,N_26164);
nand U26958 (N_26958,N_26240,N_26338);
xor U26959 (N_26959,N_26308,N_26043);
and U26960 (N_26960,N_26393,N_26100);
or U26961 (N_26961,N_26406,N_26356);
nand U26962 (N_26962,N_26424,N_26078);
xnor U26963 (N_26963,N_26107,N_26057);
nor U26964 (N_26964,N_26000,N_26010);
xor U26965 (N_26965,N_26168,N_26401);
and U26966 (N_26966,N_26179,N_26237);
and U26967 (N_26967,N_26351,N_26461);
nor U26968 (N_26968,N_26310,N_26286);
xnor U26969 (N_26969,N_26399,N_26413);
xnor U26970 (N_26970,N_26203,N_26312);
nand U26971 (N_26971,N_26047,N_26233);
nor U26972 (N_26972,N_26324,N_26350);
or U26973 (N_26973,N_26343,N_26218);
nor U26974 (N_26974,N_26048,N_26429);
nor U26975 (N_26975,N_26495,N_26255);
and U26976 (N_26976,N_26386,N_26340);
or U26977 (N_26977,N_26272,N_26033);
or U26978 (N_26978,N_26182,N_26255);
nand U26979 (N_26979,N_26029,N_26174);
or U26980 (N_26980,N_26154,N_26115);
or U26981 (N_26981,N_26486,N_26110);
and U26982 (N_26982,N_26209,N_26168);
or U26983 (N_26983,N_26243,N_26400);
or U26984 (N_26984,N_26250,N_26494);
xor U26985 (N_26985,N_26151,N_26118);
nand U26986 (N_26986,N_26288,N_26304);
xor U26987 (N_26987,N_26196,N_26218);
nor U26988 (N_26988,N_26251,N_26250);
xnor U26989 (N_26989,N_26457,N_26091);
nor U26990 (N_26990,N_26487,N_26399);
nand U26991 (N_26991,N_26471,N_26190);
and U26992 (N_26992,N_26414,N_26006);
nand U26993 (N_26993,N_26165,N_26497);
and U26994 (N_26994,N_26367,N_26442);
xor U26995 (N_26995,N_26335,N_26340);
nor U26996 (N_26996,N_26261,N_26109);
nor U26997 (N_26997,N_26247,N_26037);
or U26998 (N_26998,N_26438,N_26049);
nand U26999 (N_26999,N_26014,N_26292);
nor U27000 (N_27000,N_26650,N_26817);
and U27001 (N_27001,N_26883,N_26680);
nand U27002 (N_27002,N_26536,N_26830);
or U27003 (N_27003,N_26842,N_26845);
nor U27004 (N_27004,N_26749,N_26862);
xor U27005 (N_27005,N_26695,N_26756);
xnor U27006 (N_27006,N_26596,N_26517);
or U27007 (N_27007,N_26739,N_26580);
xor U27008 (N_27008,N_26878,N_26638);
nor U27009 (N_27009,N_26909,N_26884);
nor U27010 (N_27010,N_26791,N_26581);
or U27011 (N_27011,N_26934,N_26915);
and U27012 (N_27012,N_26571,N_26569);
and U27013 (N_27013,N_26718,N_26534);
nor U27014 (N_27014,N_26560,N_26958);
and U27015 (N_27015,N_26577,N_26998);
and U27016 (N_27016,N_26832,N_26824);
nor U27017 (N_27017,N_26576,N_26941);
nand U27018 (N_27018,N_26773,N_26837);
nor U27019 (N_27019,N_26765,N_26659);
nand U27020 (N_27020,N_26582,N_26699);
nor U27021 (N_27021,N_26991,N_26953);
and U27022 (N_27022,N_26808,N_26822);
nor U27023 (N_27023,N_26811,N_26965);
nand U27024 (N_27024,N_26508,N_26573);
or U27025 (N_27025,N_26886,N_26538);
or U27026 (N_27026,N_26684,N_26974);
nand U27027 (N_27027,N_26768,N_26733);
and U27028 (N_27028,N_26711,N_26697);
and U27029 (N_27029,N_26653,N_26829);
nand U27030 (N_27030,N_26605,N_26907);
nor U27031 (N_27031,N_26891,N_26633);
nand U27032 (N_27032,N_26637,N_26640);
and U27033 (N_27033,N_26703,N_26621);
nand U27034 (N_27034,N_26944,N_26724);
nor U27035 (N_27035,N_26720,N_26895);
or U27036 (N_27036,N_26980,N_26685);
nor U27037 (N_27037,N_26964,N_26570);
nor U27038 (N_27038,N_26537,N_26892);
nand U27039 (N_27039,N_26868,N_26696);
xnor U27040 (N_27040,N_26632,N_26962);
and U27041 (N_27041,N_26533,N_26528);
and U27042 (N_27042,N_26910,N_26922);
nor U27043 (N_27043,N_26849,N_26579);
and U27044 (N_27044,N_26505,N_26858);
or U27045 (N_27045,N_26729,N_26841);
or U27046 (N_27046,N_26549,N_26693);
nand U27047 (N_27047,N_26672,N_26903);
and U27048 (N_27048,N_26762,N_26625);
nand U27049 (N_27049,N_26595,N_26926);
and U27050 (N_27050,N_26651,N_26995);
xor U27051 (N_27051,N_26669,N_26876);
xor U27052 (N_27052,N_26561,N_26890);
and U27053 (N_27053,N_26750,N_26987);
xnor U27054 (N_27054,N_26532,N_26678);
nand U27055 (N_27055,N_26935,N_26609);
nand U27056 (N_27056,N_26742,N_26504);
or U27057 (N_27057,N_26911,N_26531);
or U27058 (N_27058,N_26847,N_26558);
nand U27059 (N_27059,N_26732,N_26951);
nand U27060 (N_27060,N_26787,N_26687);
nand U27061 (N_27061,N_26646,N_26942);
or U27062 (N_27062,N_26818,N_26740);
xor U27063 (N_27063,N_26779,N_26700);
nor U27064 (N_27064,N_26893,N_26983);
nor U27065 (N_27065,N_26937,N_26857);
and U27066 (N_27066,N_26624,N_26555);
and U27067 (N_27067,N_26919,N_26527);
or U27068 (N_27068,N_26949,N_26611);
xnor U27069 (N_27069,N_26745,N_26928);
nand U27070 (N_27070,N_26511,N_26513);
or U27071 (N_27071,N_26815,N_26856);
xor U27072 (N_27072,N_26820,N_26821);
nor U27073 (N_27073,N_26812,N_26978);
nand U27074 (N_27074,N_26599,N_26827);
nand U27075 (N_27075,N_26683,N_26789);
nand U27076 (N_27076,N_26620,N_26501);
xor U27077 (N_27077,N_26667,N_26657);
nand U27078 (N_27078,N_26925,N_26639);
and U27079 (N_27079,N_26786,N_26645);
and U27080 (N_27080,N_26722,N_26715);
and U27081 (N_27081,N_26996,N_26559);
or U27082 (N_27082,N_26810,N_26723);
xor U27083 (N_27083,N_26838,N_26590);
or U27084 (N_27084,N_26634,N_26591);
nand U27085 (N_27085,N_26675,N_26719);
nor U27086 (N_27086,N_26516,N_26557);
nand U27087 (N_27087,N_26647,N_26714);
xnor U27088 (N_27088,N_26997,N_26930);
xnor U27089 (N_27089,N_26933,N_26506);
nand U27090 (N_27090,N_26906,N_26946);
or U27091 (N_27091,N_26593,N_26548);
nand U27092 (N_27092,N_26967,N_26668);
nand U27093 (N_27093,N_26709,N_26575);
xor U27094 (N_27094,N_26870,N_26888);
nor U27095 (N_27095,N_26585,N_26831);
or U27096 (N_27096,N_26957,N_26968);
nand U27097 (N_27097,N_26807,N_26682);
nor U27098 (N_27098,N_26594,N_26689);
or U27099 (N_27099,N_26916,N_26835);
xor U27100 (N_27100,N_26660,N_26871);
nand U27101 (N_27101,N_26801,N_26502);
or U27102 (N_27102,N_26948,N_26661);
or U27103 (N_27103,N_26936,N_26523);
or U27104 (N_27104,N_26799,N_26836);
and U27105 (N_27105,N_26999,N_26840);
or U27106 (N_27106,N_26726,N_26588);
xor U27107 (N_27107,N_26704,N_26777);
nand U27108 (N_27108,N_26984,N_26526);
and U27109 (N_27109,N_26601,N_26769);
nor U27110 (N_27110,N_26943,N_26778);
or U27111 (N_27111,N_26587,N_26900);
nand U27112 (N_27112,N_26763,N_26529);
xor U27113 (N_27113,N_26955,N_26612);
nand U27114 (N_27114,N_26521,N_26618);
nor U27115 (N_27115,N_26859,N_26814);
and U27116 (N_27116,N_26986,N_26867);
and U27117 (N_27117,N_26607,N_26568);
nand U27118 (N_27118,N_26602,N_26563);
and U27119 (N_27119,N_26880,N_26960);
nand U27120 (N_27120,N_26619,N_26664);
nor U27121 (N_27121,N_26674,N_26735);
nor U27122 (N_27122,N_26804,N_26852);
or U27123 (N_27123,N_26813,N_26794);
nor U27124 (N_27124,N_26947,N_26809);
and U27125 (N_27125,N_26544,N_26597);
nand U27126 (N_27126,N_26782,N_26929);
nor U27127 (N_27127,N_26616,N_26507);
nand U27128 (N_27128,N_26872,N_26701);
and U27129 (N_27129,N_26793,N_26774);
xnor U27130 (N_27130,N_26894,N_26780);
or U27131 (N_27131,N_26716,N_26889);
and U27132 (N_27132,N_26728,N_26753);
nand U27133 (N_27133,N_26881,N_26692);
or U27134 (N_27134,N_26988,N_26717);
and U27135 (N_27135,N_26913,N_26551);
and U27136 (N_27136,N_26979,N_26865);
and U27137 (N_27137,N_26912,N_26754);
nor U27138 (N_27138,N_26673,N_26567);
nor U27139 (N_27139,N_26931,N_26874);
or U27140 (N_27140,N_26954,N_26713);
or U27141 (N_27141,N_26956,N_26795);
nand U27142 (N_27142,N_26725,N_26643);
nor U27143 (N_27143,N_26901,N_26707);
and U27144 (N_27144,N_26741,N_26604);
or U27145 (N_27145,N_26676,N_26691);
or U27146 (N_27146,N_26819,N_26710);
xnor U27147 (N_27147,N_26826,N_26792);
xnor U27148 (N_27148,N_26530,N_26851);
nand U27149 (N_27149,N_26515,N_26785);
or U27150 (N_27150,N_26738,N_26712);
nor U27151 (N_27151,N_26781,N_26545);
or U27152 (N_27152,N_26721,N_26823);
or U27153 (N_27153,N_26863,N_26914);
and U27154 (N_27154,N_26525,N_26622);
and U27155 (N_27155,N_26615,N_26921);
or U27156 (N_27156,N_26783,N_26854);
or U27157 (N_27157,N_26614,N_26552);
or U27158 (N_27158,N_26644,N_26636);
nor U27159 (N_27159,N_26514,N_26802);
nor U27160 (N_27160,N_26975,N_26706);
and U27161 (N_27161,N_26839,N_26642);
and U27162 (N_27162,N_26864,N_26879);
nand U27163 (N_27163,N_26510,N_26751);
nand U27164 (N_27164,N_26666,N_26989);
nor U27165 (N_27165,N_26629,N_26990);
nand U27166 (N_27166,N_26663,N_26603);
and U27167 (N_27167,N_26945,N_26797);
nand U27168 (N_27168,N_26952,N_26757);
nand U27169 (N_27169,N_26677,N_26737);
nor U27170 (N_27170,N_26656,N_26994);
xor U27171 (N_27171,N_26731,N_26519);
and U27172 (N_27172,N_26939,N_26985);
and U27173 (N_27173,N_26776,N_26973);
nand U27174 (N_27174,N_26679,N_26758);
nand U27175 (N_27175,N_26586,N_26578);
xor U27176 (N_27176,N_26631,N_26755);
and U27177 (N_27177,N_26882,N_26743);
and U27178 (N_27178,N_26898,N_26961);
and U27179 (N_27179,N_26690,N_26565);
nand U27180 (N_27180,N_26924,N_26566);
or U27181 (N_27181,N_26708,N_26908);
and U27182 (N_27182,N_26698,N_26736);
and U27183 (N_27183,N_26652,N_26512);
nor U27184 (N_27184,N_26535,N_26539);
nand U27185 (N_27185,N_26583,N_26784);
nand U27186 (N_27186,N_26855,N_26542);
nor U27187 (N_27187,N_26959,N_26746);
or U27188 (N_27188,N_26550,N_26972);
and U27189 (N_27189,N_26630,N_26592);
or U27190 (N_27190,N_26606,N_26613);
or U27191 (N_27191,N_26556,N_26843);
nand U27192 (N_27192,N_26627,N_26608);
nand U27193 (N_27193,N_26727,N_26553);
nor U27194 (N_27194,N_26918,N_26798);
nor U27195 (N_27195,N_26917,N_26543);
or U27196 (N_27196,N_26681,N_26833);
nor U27197 (N_27197,N_26899,N_26805);
xnor U27198 (N_27198,N_26686,N_26747);
and U27199 (N_27199,N_26770,N_26861);
or U27200 (N_27200,N_26982,N_26800);
nor U27201 (N_27201,N_26897,N_26705);
or U27202 (N_27202,N_26617,N_26626);
and U27203 (N_27203,N_26844,N_26920);
nand U27204 (N_27204,N_26966,N_26748);
xor U27205 (N_27205,N_26759,N_26963);
nor U27206 (N_27206,N_26992,N_26938);
and U27207 (N_27207,N_26702,N_26834);
or U27208 (N_27208,N_26775,N_26655);
and U27209 (N_27209,N_26860,N_26971);
xnor U27210 (N_27210,N_26658,N_26600);
nand U27211 (N_27211,N_26764,N_26546);
or U27212 (N_27212,N_26584,N_26554);
nand U27213 (N_27213,N_26628,N_26873);
nand U27214 (N_27214,N_26744,N_26500);
nand U27215 (N_27215,N_26509,N_26932);
or U27216 (N_27216,N_26766,N_26503);
and U27217 (N_27217,N_26641,N_26562);
or U27218 (N_27218,N_26665,N_26788);
nor U27219 (N_27219,N_26541,N_26752);
nor U27220 (N_27220,N_26904,N_26940);
nor U27221 (N_27221,N_26790,N_26970);
nand U27222 (N_27222,N_26734,N_26572);
and U27223 (N_27223,N_26885,N_26796);
and U27224 (N_27224,N_26887,N_26969);
and U27225 (N_27225,N_26520,N_26648);
nor U27226 (N_27226,N_26850,N_26649);
or U27227 (N_27227,N_26866,N_26671);
and U27228 (N_27228,N_26760,N_26761);
and U27229 (N_27229,N_26877,N_26977);
nand U27230 (N_27230,N_26976,N_26522);
and U27231 (N_27231,N_26670,N_26803);
and U27232 (N_27232,N_26598,N_26771);
or U27233 (N_27233,N_26905,N_26993);
nor U27234 (N_27234,N_26547,N_26896);
and U27235 (N_27235,N_26869,N_26610);
or U27236 (N_27236,N_26950,N_26518);
or U27237 (N_27237,N_26816,N_26902);
nor U27238 (N_27238,N_26853,N_26688);
xor U27239 (N_27239,N_26923,N_26623);
nor U27240 (N_27240,N_26564,N_26767);
nor U27241 (N_27241,N_26806,N_26730);
or U27242 (N_27242,N_26875,N_26540);
nor U27243 (N_27243,N_26846,N_26662);
nand U27244 (N_27244,N_26772,N_26981);
nand U27245 (N_27245,N_26848,N_26927);
xnor U27246 (N_27246,N_26635,N_26589);
nand U27247 (N_27247,N_26654,N_26524);
nand U27248 (N_27248,N_26828,N_26694);
nand U27249 (N_27249,N_26825,N_26574);
nand U27250 (N_27250,N_26677,N_26578);
or U27251 (N_27251,N_26608,N_26618);
nor U27252 (N_27252,N_26740,N_26822);
nor U27253 (N_27253,N_26900,N_26674);
or U27254 (N_27254,N_26989,N_26664);
nand U27255 (N_27255,N_26527,N_26753);
or U27256 (N_27256,N_26579,N_26946);
or U27257 (N_27257,N_26656,N_26889);
and U27258 (N_27258,N_26857,N_26594);
xor U27259 (N_27259,N_26875,N_26589);
nor U27260 (N_27260,N_26585,N_26872);
nand U27261 (N_27261,N_26540,N_26651);
nand U27262 (N_27262,N_26801,N_26869);
or U27263 (N_27263,N_26939,N_26515);
nand U27264 (N_27264,N_26510,N_26794);
and U27265 (N_27265,N_26941,N_26677);
and U27266 (N_27266,N_26716,N_26555);
or U27267 (N_27267,N_26865,N_26936);
nor U27268 (N_27268,N_26913,N_26568);
xor U27269 (N_27269,N_26616,N_26703);
nand U27270 (N_27270,N_26660,N_26693);
nor U27271 (N_27271,N_26505,N_26846);
and U27272 (N_27272,N_26978,N_26788);
or U27273 (N_27273,N_26758,N_26940);
nor U27274 (N_27274,N_26878,N_26644);
nand U27275 (N_27275,N_26666,N_26913);
and U27276 (N_27276,N_26809,N_26690);
nand U27277 (N_27277,N_26993,N_26898);
and U27278 (N_27278,N_26515,N_26604);
nor U27279 (N_27279,N_26586,N_26817);
nor U27280 (N_27280,N_26654,N_26672);
or U27281 (N_27281,N_26900,N_26626);
nor U27282 (N_27282,N_26842,N_26897);
nand U27283 (N_27283,N_26909,N_26727);
or U27284 (N_27284,N_26790,N_26776);
xor U27285 (N_27285,N_26978,N_26521);
nand U27286 (N_27286,N_26540,N_26930);
or U27287 (N_27287,N_26937,N_26643);
or U27288 (N_27288,N_26614,N_26568);
nand U27289 (N_27289,N_26746,N_26643);
nand U27290 (N_27290,N_26902,N_26561);
nor U27291 (N_27291,N_26926,N_26898);
and U27292 (N_27292,N_26678,N_26970);
and U27293 (N_27293,N_26835,N_26843);
and U27294 (N_27294,N_26540,N_26929);
nor U27295 (N_27295,N_26864,N_26597);
and U27296 (N_27296,N_26735,N_26924);
nand U27297 (N_27297,N_26950,N_26629);
nor U27298 (N_27298,N_26812,N_26992);
xor U27299 (N_27299,N_26890,N_26619);
nand U27300 (N_27300,N_26811,N_26558);
and U27301 (N_27301,N_26892,N_26801);
and U27302 (N_27302,N_26791,N_26880);
and U27303 (N_27303,N_26525,N_26918);
nor U27304 (N_27304,N_26953,N_26814);
and U27305 (N_27305,N_26973,N_26982);
nand U27306 (N_27306,N_26883,N_26698);
nand U27307 (N_27307,N_26990,N_26787);
nand U27308 (N_27308,N_26949,N_26774);
nand U27309 (N_27309,N_26840,N_26907);
nand U27310 (N_27310,N_26593,N_26536);
and U27311 (N_27311,N_26978,N_26846);
xnor U27312 (N_27312,N_26651,N_26627);
and U27313 (N_27313,N_26650,N_26761);
nor U27314 (N_27314,N_26896,N_26664);
nand U27315 (N_27315,N_26509,N_26580);
or U27316 (N_27316,N_26759,N_26593);
or U27317 (N_27317,N_26520,N_26573);
and U27318 (N_27318,N_26889,N_26645);
nor U27319 (N_27319,N_26535,N_26553);
nand U27320 (N_27320,N_26602,N_26880);
or U27321 (N_27321,N_26551,N_26701);
or U27322 (N_27322,N_26829,N_26847);
nor U27323 (N_27323,N_26907,N_26500);
or U27324 (N_27324,N_26614,N_26527);
or U27325 (N_27325,N_26784,N_26788);
nand U27326 (N_27326,N_26847,N_26846);
and U27327 (N_27327,N_26793,N_26962);
nand U27328 (N_27328,N_26508,N_26614);
and U27329 (N_27329,N_26818,N_26927);
and U27330 (N_27330,N_26566,N_26688);
and U27331 (N_27331,N_26844,N_26871);
or U27332 (N_27332,N_26783,N_26612);
or U27333 (N_27333,N_26573,N_26602);
nand U27334 (N_27334,N_26880,N_26936);
nor U27335 (N_27335,N_26722,N_26558);
and U27336 (N_27336,N_26505,N_26800);
and U27337 (N_27337,N_26699,N_26786);
xor U27338 (N_27338,N_26889,N_26647);
nand U27339 (N_27339,N_26517,N_26844);
nand U27340 (N_27340,N_26500,N_26502);
nor U27341 (N_27341,N_26686,N_26873);
xnor U27342 (N_27342,N_26615,N_26651);
nand U27343 (N_27343,N_26878,N_26653);
or U27344 (N_27344,N_26936,N_26553);
and U27345 (N_27345,N_26973,N_26679);
nand U27346 (N_27346,N_26855,N_26826);
and U27347 (N_27347,N_26918,N_26896);
or U27348 (N_27348,N_26713,N_26756);
xor U27349 (N_27349,N_26885,N_26522);
and U27350 (N_27350,N_26820,N_26664);
and U27351 (N_27351,N_26910,N_26873);
nor U27352 (N_27352,N_26692,N_26981);
nand U27353 (N_27353,N_26981,N_26785);
and U27354 (N_27354,N_26590,N_26835);
nor U27355 (N_27355,N_26830,N_26544);
and U27356 (N_27356,N_26740,N_26782);
nand U27357 (N_27357,N_26967,N_26809);
or U27358 (N_27358,N_26754,N_26722);
xnor U27359 (N_27359,N_26556,N_26876);
and U27360 (N_27360,N_26880,N_26870);
nand U27361 (N_27361,N_26629,N_26612);
nor U27362 (N_27362,N_26595,N_26504);
nand U27363 (N_27363,N_26565,N_26731);
nand U27364 (N_27364,N_26791,N_26631);
nor U27365 (N_27365,N_26886,N_26588);
and U27366 (N_27366,N_26953,N_26995);
or U27367 (N_27367,N_26937,N_26664);
nand U27368 (N_27368,N_26587,N_26940);
xnor U27369 (N_27369,N_26889,N_26830);
nand U27370 (N_27370,N_26678,N_26835);
nor U27371 (N_27371,N_26891,N_26524);
nor U27372 (N_27372,N_26804,N_26999);
nand U27373 (N_27373,N_26532,N_26617);
or U27374 (N_27374,N_26719,N_26808);
xnor U27375 (N_27375,N_26669,N_26676);
nor U27376 (N_27376,N_26883,N_26541);
nand U27377 (N_27377,N_26575,N_26682);
nor U27378 (N_27378,N_26780,N_26923);
and U27379 (N_27379,N_26591,N_26723);
or U27380 (N_27380,N_26666,N_26595);
nor U27381 (N_27381,N_26667,N_26769);
xor U27382 (N_27382,N_26679,N_26616);
or U27383 (N_27383,N_26962,N_26825);
and U27384 (N_27384,N_26807,N_26532);
nand U27385 (N_27385,N_26871,N_26582);
nand U27386 (N_27386,N_26550,N_26988);
or U27387 (N_27387,N_26767,N_26697);
nand U27388 (N_27388,N_26719,N_26735);
nand U27389 (N_27389,N_26806,N_26932);
and U27390 (N_27390,N_26682,N_26979);
or U27391 (N_27391,N_26764,N_26745);
nor U27392 (N_27392,N_26951,N_26561);
and U27393 (N_27393,N_26862,N_26832);
nand U27394 (N_27394,N_26510,N_26528);
or U27395 (N_27395,N_26602,N_26954);
and U27396 (N_27396,N_26983,N_26695);
and U27397 (N_27397,N_26975,N_26718);
nand U27398 (N_27398,N_26783,N_26604);
and U27399 (N_27399,N_26812,N_26605);
nand U27400 (N_27400,N_26548,N_26679);
nor U27401 (N_27401,N_26643,N_26822);
and U27402 (N_27402,N_26766,N_26957);
or U27403 (N_27403,N_26902,N_26717);
or U27404 (N_27404,N_26788,N_26625);
or U27405 (N_27405,N_26889,N_26704);
nand U27406 (N_27406,N_26812,N_26828);
nor U27407 (N_27407,N_26661,N_26619);
or U27408 (N_27408,N_26955,N_26831);
and U27409 (N_27409,N_26645,N_26673);
nand U27410 (N_27410,N_26891,N_26725);
nand U27411 (N_27411,N_26878,N_26852);
xnor U27412 (N_27412,N_26558,N_26816);
and U27413 (N_27413,N_26639,N_26857);
nand U27414 (N_27414,N_26631,N_26928);
and U27415 (N_27415,N_26917,N_26666);
nand U27416 (N_27416,N_26763,N_26839);
nand U27417 (N_27417,N_26679,N_26528);
nor U27418 (N_27418,N_26895,N_26819);
and U27419 (N_27419,N_26988,N_26959);
or U27420 (N_27420,N_26716,N_26758);
nand U27421 (N_27421,N_26986,N_26602);
nand U27422 (N_27422,N_26521,N_26981);
xnor U27423 (N_27423,N_26869,N_26663);
or U27424 (N_27424,N_26887,N_26797);
nand U27425 (N_27425,N_26799,N_26569);
nand U27426 (N_27426,N_26793,N_26617);
nor U27427 (N_27427,N_26987,N_26836);
nand U27428 (N_27428,N_26712,N_26618);
nor U27429 (N_27429,N_26619,N_26787);
and U27430 (N_27430,N_26714,N_26827);
or U27431 (N_27431,N_26971,N_26783);
nand U27432 (N_27432,N_26963,N_26727);
nand U27433 (N_27433,N_26528,N_26762);
xor U27434 (N_27434,N_26822,N_26604);
xor U27435 (N_27435,N_26992,N_26785);
xnor U27436 (N_27436,N_26566,N_26525);
nand U27437 (N_27437,N_26904,N_26695);
nand U27438 (N_27438,N_26535,N_26597);
nor U27439 (N_27439,N_26602,N_26513);
nor U27440 (N_27440,N_26799,N_26812);
or U27441 (N_27441,N_26863,N_26692);
nor U27442 (N_27442,N_26510,N_26756);
or U27443 (N_27443,N_26924,N_26851);
or U27444 (N_27444,N_26871,N_26540);
or U27445 (N_27445,N_26787,N_26755);
nand U27446 (N_27446,N_26596,N_26901);
nand U27447 (N_27447,N_26734,N_26806);
nor U27448 (N_27448,N_26602,N_26709);
nand U27449 (N_27449,N_26740,N_26717);
or U27450 (N_27450,N_26751,N_26913);
and U27451 (N_27451,N_26876,N_26887);
nand U27452 (N_27452,N_26996,N_26983);
xor U27453 (N_27453,N_26620,N_26522);
or U27454 (N_27454,N_26672,N_26571);
or U27455 (N_27455,N_26624,N_26669);
nand U27456 (N_27456,N_26561,N_26930);
and U27457 (N_27457,N_26774,N_26968);
and U27458 (N_27458,N_26567,N_26655);
or U27459 (N_27459,N_26838,N_26907);
and U27460 (N_27460,N_26735,N_26937);
nand U27461 (N_27461,N_26989,N_26563);
and U27462 (N_27462,N_26920,N_26784);
nand U27463 (N_27463,N_26549,N_26642);
xnor U27464 (N_27464,N_26545,N_26833);
nand U27465 (N_27465,N_26860,N_26761);
nand U27466 (N_27466,N_26779,N_26638);
xor U27467 (N_27467,N_26828,N_26838);
and U27468 (N_27468,N_26780,N_26702);
nor U27469 (N_27469,N_26913,N_26620);
and U27470 (N_27470,N_26730,N_26634);
nand U27471 (N_27471,N_26693,N_26803);
nor U27472 (N_27472,N_26509,N_26794);
and U27473 (N_27473,N_26681,N_26794);
nand U27474 (N_27474,N_26722,N_26961);
nand U27475 (N_27475,N_26637,N_26739);
nor U27476 (N_27476,N_26667,N_26818);
nand U27477 (N_27477,N_26846,N_26820);
and U27478 (N_27478,N_26680,N_26691);
nand U27479 (N_27479,N_26823,N_26646);
nand U27480 (N_27480,N_26801,N_26542);
xnor U27481 (N_27481,N_26555,N_26616);
and U27482 (N_27482,N_26979,N_26546);
xnor U27483 (N_27483,N_26590,N_26858);
and U27484 (N_27484,N_26745,N_26529);
or U27485 (N_27485,N_26591,N_26712);
xnor U27486 (N_27486,N_26593,N_26774);
nand U27487 (N_27487,N_26536,N_26723);
nand U27488 (N_27488,N_26688,N_26536);
xor U27489 (N_27489,N_26837,N_26672);
and U27490 (N_27490,N_26560,N_26547);
xor U27491 (N_27491,N_26617,N_26582);
nor U27492 (N_27492,N_26560,N_26599);
and U27493 (N_27493,N_26610,N_26984);
and U27494 (N_27494,N_26538,N_26707);
nand U27495 (N_27495,N_26560,N_26937);
nor U27496 (N_27496,N_26582,N_26575);
xor U27497 (N_27497,N_26535,N_26505);
nor U27498 (N_27498,N_26929,N_26631);
and U27499 (N_27499,N_26988,N_26801);
nand U27500 (N_27500,N_27308,N_27204);
nor U27501 (N_27501,N_27357,N_27222);
nor U27502 (N_27502,N_27274,N_27095);
nand U27503 (N_27503,N_27226,N_27118);
and U27504 (N_27504,N_27399,N_27296);
and U27505 (N_27505,N_27041,N_27255);
nor U27506 (N_27506,N_27326,N_27049);
or U27507 (N_27507,N_27024,N_27079);
nor U27508 (N_27508,N_27054,N_27432);
and U27509 (N_27509,N_27100,N_27203);
nor U27510 (N_27510,N_27172,N_27408);
xnor U27511 (N_27511,N_27253,N_27328);
nor U27512 (N_27512,N_27365,N_27461);
or U27513 (N_27513,N_27477,N_27021);
nor U27514 (N_27514,N_27367,N_27020);
and U27515 (N_27515,N_27097,N_27352);
nor U27516 (N_27516,N_27320,N_27453);
and U27517 (N_27517,N_27363,N_27149);
or U27518 (N_27518,N_27498,N_27317);
or U27519 (N_27519,N_27252,N_27474);
xor U27520 (N_27520,N_27034,N_27346);
or U27521 (N_27521,N_27398,N_27211);
nor U27522 (N_27522,N_27392,N_27212);
nor U27523 (N_27523,N_27166,N_27364);
nand U27524 (N_27524,N_27048,N_27366);
nand U27525 (N_27525,N_27455,N_27194);
nand U27526 (N_27526,N_27153,N_27450);
or U27527 (N_27527,N_27496,N_27445);
xor U27528 (N_27528,N_27428,N_27487);
nand U27529 (N_27529,N_27281,N_27161);
or U27530 (N_27530,N_27080,N_27176);
nand U27531 (N_27531,N_27259,N_27099);
and U27532 (N_27532,N_27311,N_27451);
and U27533 (N_27533,N_27094,N_27427);
and U27534 (N_27534,N_27234,N_27199);
or U27535 (N_27535,N_27307,N_27171);
or U27536 (N_27536,N_27385,N_27288);
and U27537 (N_27537,N_27125,N_27232);
and U27538 (N_27538,N_27287,N_27179);
xor U27539 (N_27539,N_27060,N_27042);
nand U27540 (N_27540,N_27243,N_27278);
nand U27541 (N_27541,N_27121,N_27272);
and U27542 (N_27542,N_27207,N_27492);
and U27543 (N_27543,N_27426,N_27009);
xor U27544 (N_27544,N_27425,N_27472);
nand U27545 (N_27545,N_27490,N_27050);
nand U27546 (N_27546,N_27333,N_27303);
nand U27547 (N_27547,N_27456,N_27025);
nand U27548 (N_27548,N_27197,N_27148);
and U27549 (N_27549,N_27129,N_27460);
and U27550 (N_27550,N_27375,N_27033);
or U27551 (N_27551,N_27292,N_27324);
or U27552 (N_27552,N_27098,N_27202);
or U27553 (N_27553,N_27184,N_27290);
xnor U27554 (N_27554,N_27400,N_27383);
or U27555 (N_27555,N_27002,N_27151);
and U27556 (N_27556,N_27348,N_27231);
nor U27557 (N_27557,N_27051,N_27217);
and U27558 (N_27558,N_27423,N_27407);
nand U27559 (N_27559,N_27209,N_27242);
nand U27560 (N_27560,N_27101,N_27028);
nand U27561 (N_27561,N_27391,N_27146);
nor U27562 (N_27562,N_27168,N_27145);
nand U27563 (N_27563,N_27323,N_27486);
nor U27564 (N_27564,N_27201,N_27373);
nand U27565 (N_27565,N_27330,N_27036);
and U27566 (N_27566,N_27260,N_27052);
or U27567 (N_27567,N_27283,N_27340);
nor U27568 (N_27568,N_27044,N_27047);
nor U27569 (N_27569,N_27318,N_27435);
or U27570 (N_27570,N_27132,N_27314);
and U27571 (N_27571,N_27447,N_27462);
nand U27572 (N_27572,N_27141,N_27069);
nor U27573 (N_27573,N_27291,N_27017);
xnor U27574 (N_27574,N_27264,N_27062);
or U27575 (N_27575,N_27342,N_27188);
xor U27576 (N_27576,N_27268,N_27421);
nand U27577 (N_27577,N_27302,N_27227);
nand U27578 (N_27578,N_27313,N_27003);
nand U27579 (N_27579,N_27196,N_27219);
and U27580 (N_27580,N_27241,N_27183);
nor U27581 (N_27581,N_27481,N_27466);
xnor U27582 (N_27582,N_27422,N_27465);
nand U27583 (N_27583,N_27412,N_27133);
or U27584 (N_27584,N_27381,N_27256);
nand U27585 (N_27585,N_27390,N_27355);
xor U27586 (N_27586,N_27289,N_27103);
and U27587 (N_27587,N_27198,N_27306);
nor U27588 (N_27588,N_27075,N_27066);
xor U27589 (N_27589,N_27248,N_27473);
xnor U27590 (N_27590,N_27011,N_27218);
xor U27591 (N_27591,N_27470,N_27074);
or U27592 (N_27592,N_27345,N_27378);
nor U27593 (N_27593,N_27005,N_27065);
nand U27594 (N_27594,N_27039,N_27404);
and U27595 (N_27595,N_27464,N_27082);
and U27596 (N_27596,N_27413,N_27055);
xnor U27597 (N_27597,N_27495,N_27104);
nor U27598 (N_27598,N_27270,N_27371);
nor U27599 (N_27599,N_27022,N_27078);
and U27600 (N_27600,N_27059,N_27216);
and U27601 (N_27601,N_27434,N_27221);
nor U27602 (N_27602,N_27395,N_27163);
nor U27603 (N_27603,N_27489,N_27170);
or U27604 (N_27604,N_27027,N_27416);
or U27605 (N_27605,N_27494,N_27117);
and U27606 (N_27606,N_27147,N_27092);
nor U27607 (N_27607,N_27093,N_27205);
nand U27608 (N_27608,N_27338,N_27158);
or U27609 (N_27609,N_27137,N_27483);
nand U27610 (N_27610,N_27354,N_27106);
or U27611 (N_27611,N_27388,N_27006);
or U27612 (N_27612,N_27443,N_27126);
nor U27613 (N_27613,N_27056,N_27479);
nor U27614 (N_27614,N_27294,N_27436);
nand U27615 (N_27615,N_27418,N_27402);
nor U27616 (N_27616,N_27411,N_27332);
xnor U27617 (N_27617,N_27076,N_27361);
nand U27618 (N_27618,N_27123,N_27085);
or U27619 (N_27619,N_27190,N_27305);
or U27620 (N_27620,N_27182,N_27316);
nor U27621 (N_27621,N_27206,N_27409);
nand U27622 (N_27622,N_27279,N_27084);
nor U27623 (N_27623,N_27077,N_27269);
and U27624 (N_27624,N_27417,N_27458);
or U27625 (N_27625,N_27112,N_27230);
nor U27626 (N_27626,N_27459,N_27349);
or U27627 (N_27627,N_27178,N_27235);
or U27628 (N_27628,N_27224,N_27249);
and U27629 (N_27629,N_27467,N_27040);
and U27630 (N_27630,N_27007,N_27030);
nand U27631 (N_27631,N_27322,N_27299);
xor U27632 (N_27632,N_27236,N_27159);
xor U27633 (N_27633,N_27446,N_27251);
or U27634 (N_27634,N_27499,N_27189);
nand U27635 (N_27635,N_27008,N_27061);
or U27636 (N_27636,N_27312,N_27156);
nand U27637 (N_27637,N_27067,N_27396);
nor U27638 (N_27638,N_27140,N_27327);
xor U27639 (N_27639,N_27334,N_27239);
nor U27640 (N_27640,N_27120,N_27439);
or U27641 (N_27641,N_27444,N_27023);
nand U27642 (N_27642,N_27257,N_27379);
xnor U27643 (N_27643,N_27468,N_27452);
xnor U27644 (N_27644,N_27154,N_27053);
and U27645 (N_27645,N_27142,N_27362);
nor U27646 (N_27646,N_27174,N_27448);
nand U27647 (N_27647,N_27130,N_27293);
nor U27648 (N_27648,N_27360,N_27480);
or U27649 (N_27649,N_27081,N_27454);
nor U27650 (N_27650,N_27070,N_27261);
and U27651 (N_27651,N_27277,N_27115);
or U27652 (N_27652,N_27116,N_27353);
or U27653 (N_27653,N_27043,N_27245);
nand U27654 (N_27654,N_27157,N_27128);
and U27655 (N_27655,N_27233,N_27215);
nand U27656 (N_27656,N_27406,N_27238);
nor U27657 (N_27657,N_27343,N_27484);
nand U27658 (N_27658,N_27437,N_27463);
and U27659 (N_27659,N_27032,N_27150);
or U27660 (N_27660,N_27029,N_27136);
and U27661 (N_27661,N_27482,N_27026);
nand U27662 (N_27662,N_27135,N_27329);
or U27663 (N_27663,N_27018,N_27152);
or U27664 (N_27664,N_27393,N_27262);
and U27665 (N_27665,N_27380,N_27193);
or U27666 (N_27666,N_27019,N_27250);
nand U27667 (N_27667,N_27058,N_27280);
nor U27668 (N_27668,N_27321,N_27109);
and U27669 (N_27669,N_27223,N_27089);
nor U27670 (N_27670,N_27341,N_27297);
and U27671 (N_27671,N_27471,N_27405);
nor U27672 (N_27672,N_27073,N_27335);
and U27673 (N_27673,N_27001,N_27394);
or U27674 (N_27674,N_27382,N_27139);
or U27675 (N_27675,N_27491,N_27195);
and U27676 (N_27676,N_27387,N_27497);
nand U27677 (N_27677,N_27310,N_27347);
xor U27678 (N_27678,N_27038,N_27068);
or U27679 (N_27679,N_27108,N_27441);
nor U27680 (N_27680,N_27397,N_27298);
or U27681 (N_27681,N_27185,N_27493);
nor U27682 (N_27682,N_27114,N_27225);
nor U27683 (N_27683,N_27370,N_27263);
nand U27684 (N_27684,N_27071,N_27440);
nor U27685 (N_27685,N_27384,N_27300);
and U27686 (N_27686,N_27469,N_27275);
nand U27687 (N_27687,N_27015,N_27372);
nand U27688 (N_27688,N_27265,N_27045);
or U27689 (N_27689,N_27107,N_27415);
nand U27690 (N_27690,N_27119,N_27358);
nor U27691 (N_27691,N_27127,N_27475);
or U27692 (N_27692,N_27111,N_27144);
and U27693 (N_27693,N_27177,N_27000);
nor U27694 (N_27694,N_27319,N_27401);
nand U27695 (N_27695,N_27337,N_27210);
or U27696 (N_27696,N_27339,N_27386);
nand U27697 (N_27697,N_27431,N_27229);
and U27698 (N_27698,N_27162,N_27273);
nand U27699 (N_27699,N_27488,N_27301);
nand U27700 (N_27700,N_27012,N_27403);
or U27701 (N_27701,N_27110,N_27134);
nand U27702 (N_27702,N_27004,N_27186);
nand U27703 (N_27703,N_27072,N_27155);
xnor U27704 (N_27704,N_27258,N_27377);
nand U27705 (N_27705,N_27331,N_27429);
or U27706 (N_27706,N_27284,N_27063);
nor U27707 (N_27707,N_27336,N_27304);
nand U27708 (N_27708,N_27187,N_27088);
nand U27709 (N_27709,N_27181,N_27037);
nand U27710 (N_27710,N_27192,N_27457);
nor U27711 (N_27711,N_27143,N_27369);
nor U27712 (N_27712,N_27351,N_27350);
and U27713 (N_27713,N_27105,N_27374);
and U27714 (N_27714,N_27282,N_27035);
nand U27715 (N_27715,N_27124,N_27169);
and U27716 (N_27716,N_27131,N_27414);
nand U27717 (N_27717,N_27449,N_27276);
nor U27718 (N_27718,N_27213,N_27285);
xor U27719 (N_27719,N_27064,N_27090);
and U27720 (N_27720,N_27376,N_27368);
and U27721 (N_27721,N_27359,N_27016);
nor U27722 (N_27722,N_27086,N_27246);
and U27723 (N_27723,N_27325,N_27267);
nor U27724 (N_27724,N_27228,N_27102);
nand U27725 (N_27725,N_27442,N_27485);
xor U27726 (N_27726,N_27167,N_27244);
nand U27727 (N_27727,N_27430,N_27014);
xor U27728 (N_27728,N_27010,N_27410);
nor U27729 (N_27729,N_27254,N_27122);
or U27730 (N_27730,N_27091,N_27113);
or U27731 (N_27731,N_27344,N_27164);
nand U27732 (N_27732,N_27476,N_27295);
nor U27733 (N_27733,N_27057,N_27478);
nand U27734 (N_27734,N_27165,N_27424);
or U27735 (N_27735,N_27083,N_27087);
or U27736 (N_27736,N_27271,N_27046);
or U27737 (N_27737,N_27266,N_27356);
nand U27738 (N_27738,N_27309,N_27175);
or U27739 (N_27739,N_27173,N_27180);
nor U27740 (N_27740,N_27096,N_27208);
nor U27741 (N_27741,N_27220,N_27389);
and U27742 (N_27742,N_27433,N_27315);
and U27743 (N_27743,N_27286,N_27031);
nor U27744 (N_27744,N_27191,N_27438);
nor U27745 (N_27745,N_27420,N_27214);
nor U27746 (N_27746,N_27200,N_27160);
or U27747 (N_27747,N_27419,N_27138);
nand U27748 (N_27748,N_27247,N_27237);
or U27749 (N_27749,N_27013,N_27240);
and U27750 (N_27750,N_27276,N_27249);
xnor U27751 (N_27751,N_27485,N_27492);
and U27752 (N_27752,N_27007,N_27134);
or U27753 (N_27753,N_27355,N_27325);
nand U27754 (N_27754,N_27492,N_27071);
and U27755 (N_27755,N_27417,N_27467);
or U27756 (N_27756,N_27281,N_27094);
or U27757 (N_27757,N_27302,N_27150);
nand U27758 (N_27758,N_27302,N_27435);
and U27759 (N_27759,N_27321,N_27315);
nor U27760 (N_27760,N_27499,N_27236);
nand U27761 (N_27761,N_27045,N_27163);
and U27762 (N_27762,N_27132,N_27190);
or U27763 (N_27763,N_27427,N_27241);
and U27764 (N_27764,N_27225,N_27195);
nor U27765 (N_27765,N_27083,N_27187);
xor U27766 (N_27766,N_27305,N_27344);
and U27767 (N_27767,N_27173,N_27178);
nor U27768 (N_27768,N_27006,N_27103);
and U27769 (N_27769,N_27387,N_27482);
xor U27770 (N_27770,N_27015,N_27462);
xor U27771 (N_27771,N_27126,N_27230);
nor U27772 (N_27772,N_27015,N_27298);
xor U27773 (N_27773,N_27263,N_27498);
xnor U27774 (N_27774,N_27233,N_27316);
nor U27775 (N_27775,N_27106,N_27398);
nand U27776 (N_27776,N_27441,N_27329);
or U27777 (N_27777,N_27275,N_27149);
or U27778 (N_27778,N_27410,N_27485);
nand U27779 (N_27779,N_27002,N_27403);
nor U27780 (N_27780,N_27246,N_27416);
nor U27781 (N_27781,N_27258,N_27133);
nand U27782 (N_27782,N_27037,N_27224);
and U27783 (N_27783,N_27262,N_27107);
nor U27784 (N_27784,N_27378,N_27398);
or U27785 (N_27785,N_27061,N_27094);
nor U27786 (N_27786,N_27461,N_27348);
or U27787 (N_27787,N_27318,N_27083);
nand U27788 (N_27788,N_27032,N_27057);
xnor U27789 (N_27789,N_27468,N_27327);
or U27790 (N_27790,N_27218,N_27342);
nor U27791 (N_27791,N_27398,N_27035);
or U27792 (N_27792,N_27062,N_27430);
nor U27793 (N_27793,N_27209,N_27461);
nor U27794 (N_27794,N_27192,N_27338);
nand U27795 (N_27795,N_27318,N_27352);
nand U27796 (N_27796,N_27352,N_27110);
xnor U27797 (N_27797,N_27030,N_27065);
nor U27798 (N_27798,N_27215,N_27313);
nor U27799 (N_27799,N_27229,N_27111);
nor U27800 (N_27800,N_27138,N_27049);
nor U27801 (N_27801,N_27313,N_27017);
nand U27802 (N_27802,N_27081,N_27166);
nor U27803 (N_27803,N_27082,N_27306);
and U27804 (N_27804,N_27207,N_27173);
and U27805 (N_27805,N_27343,N_27165);
nand U27806 (N_27806,N_27095,N_27424);
and U27807 (N_27807,N_27075,N_27383);
and U27808 (N_27808,N_27332,N_27360);
or U27809 (N_27809,N_27001,N_27332);
nand U27810 (N_27810,N_27101,N_27209);
nor U27811 (N_27811,N_27396,N_27377);
and U27812 (N_27812,N_27381,N_27200);
nand U27813 (N_27813,N_27003,N_27173);
nor U27814 (N_27814,N_27057,N_27413);
nand U27815 (N_27815,N_27249,N_27288);
nand U27816 (N_27816,N_27429,N_27222);
nor U27817 (N_27817,N_27156,N_27372);
nor U27818 (N_27818,N_27125,N_27461);
nor U27819 (N_27819,N_27120,N_27237);
or U27820 (N_27820,N_27183,N_27390);
nand U27821 (N_27821,N_27280,N_27368);
or U27822 (N_27822,N_27114,N_27213);
or U27823 (N_27823,N_27174,N_27042);
and U27824 (N_27824,N_27261,N_27172);
xor U27825 (N_27825,N_27295,N_27025);
and U27826 (N_27826,N_27406,N_27016);
nand U27827 (N_27827,N_27036,N_27008);
nor U27828 (N_27828,N_27164,N_27127);
nand U27829 (N_27829,N_27127,N_27278);
and U27830 (N_27830,N_27286,N_27307);
nor U27831 (N_27831,N_27414,N_27267);
nor U27832 (N_27832,N_27081,N_27193);
or U27833 (N_27833,N_27099,N_27288);
nand U27834 (N_27834,N_27164,N_27117);
or U27835 (N_27835,N_27330,N_27283);
or U27836 (N_27836,N_27443,N_27142);
nand U27837 (N_27837,N_27398,N_27052);
nor U27838 (N_27838,N_27032,N_27400);
or U27839 (N_27839,N_27268,N_27300);
nand U27840 (N_27840,N_27083,N_27431);
nor U27841 (N_27841,N_27206,N_27482);
xor U27842 (N_27842,N_27267,N_27389);
nor U27843 (N_27843,N_27477,N_27111);
and U27844 (N_27844,N_27160,N_27104);
nor U27845 (N_27845,N_27065,N_27054);
or U27846 (N_27846,N_27161,N_27235);
nand U27847 (N_27847,N_27194,N_27135);
or U27848 (N_27848,N_27280,N_27303);
or U27849 (N_27849,N_27428,N_27159);
xnor U27850 (N_27850,N_27029,N_27202);
xor U27851 (N_27851,N_27385,N_27188);
or U27852 (N_27852,N_27368,N_27382);
nand U27853 (N_27853,N_27208,N_27020);
nand U27854 (N_27854,N_27413,N_27498);
and U27855 (N_27855,N_27139,N_27101);
nand U27856 (N_27856,N_27130,N_27434);
nor U27857 (N_27857,N_27479,N_27434);
or U27858 (N_27858,N_27328,N_27125);
xnor U27859 (N_27859,N_27020,N_27124);
or U27860 (N_27860,N_27095,N_27186);
or U27861 (N_27861,N_27478,N_27066);
nor U27862 (N_27862,N_27344,N_27034);
nand U27863 (N_27863,N_27110,N_27049);
and U27864 (N_27864,N_27361,N_27354);
or U27865 (N_27865,N_27377,N_27163);
or U27866 (N_27866,N_27096,N_27443);
nand U27867 (N_27867,N_27216,N_27370);
and U27868 (N_27868,N_27089,N_27382);
and U27869 (N_27869,N_27125,N_27343);
nor U27870 (N_27870,N_27420,N_27044);
xor U27871 (N_27871,N_27134,N_27060);
nand U27872 (N_27872,N_27094,N_27039);
or U27873 (N_27873,N_27212,N_27390);
and U27874 (N_27874,N_27356,N_27430);
and U27875 (N_27875,N_27045,N_27390);
nand U27876 (N_27876,N_27435,N_27352);
nand U27877 (N_27877,N_27129,N_27004);
and U27878 (N_27878,N_27193,N_27106);
and U27879 (N_27879,N_27264,N_27495);
nor U27880 (N_27880,N_27412,N_27242);
xor U27881 (N_27881,N_27100,N_27300);
nand U27882 (N_27882,N_27262,N_27494);
or U27883 (N_27883,N_27484,N_27095);
or U27884 (N_27884,N_27414,N_27047);
nand U27885 (N_27885,N_27280,N_27255);
nor U27886 (N_27886,N_27462,N_27166);
xor U27887 (N_27887,N_27311,N_27250);
nor U27888 (N_27888,N_27052,N_27000);
and U27889 (N_27889,N_27060,N_27238);
nand U27890 (N_27890,N_27358,N_27209);
and U27891 (N_27891,N_27479,N_27381);
nand U27892 (N_27892,N_27283,N_27160);
nand U27893 (N_27893,N_27194,N_27233);
nand U27894 (N_27894,N_27346,N_27020);
and U27895 (N_27895,N_27477,N_27001);
and U27896 (N_27896,N_27259,N_27417);
and U27897 (N_27897,N_27414,N_27466);
nor U27898 (N_27898,N_27282,N_27328);
nand U27899 (N_27899,N_27480,N_27129);
nor U27900 (N_27900,N_27330,N_27138);
nor U27901 (N_27901,N_27278,N_27094);
nor U27902 (N_27902,N_27415,N_27445);
nand U27903 (N_27903,N_27310,N_27246);
and U27904 (N_27904,N_27392,N_27263);
nor U27905 (N_27905,N_27497,N_27128);
nand U27906 (N_27906,N_27125,N_27433);
or U27907 (N_27907,N_27275,N_27097);
xnor U27908 (N_27908,N_27192,N_27160);
or U27909 (N_27909,N_27084,N_27290);
or U27910 (N_27910,N_27479,N_27498);
or U27911 (N_27911,N_27111,N_27489);
nor U27912 (N_27912,N_27198,N_27378);
or U27913 (N_27913,N_27138,N_27073);
and U27914 (N_27914,N_27018,N_27022);
nor U27915 (N_27915,N_27119,N_27227);
or U27916 (N_27916,N_27279,N_27146);
or U27917 (N_27917,N_27080,N_27114);
nand U27918 (N_27918,N_27437,N_27188);
nand U27919 (N_27919,N_27381,N_27399);
nand U27920 (N_27920,N_27354,N_27054);
nand U27921 (N_27921,N_27084,N_27167);
and U27922 (N_27922,N_27275,N_27388);
nor U27923 (N_27923,N_27006,N_27424);
and U27924 (N_27924,N_27481,N_27090);
nand U27925 (N_27925,N_27232,N_27488);
and U27926 (N_27926,N_27208,N_27032);
or U27927 (N_27927,N_27240,N_27148);
nor U27928 (N_27928,N_27451,N_27033);
nand U27929 (N_27929,N_27096,N_27102);
and U27930 (N_27930,N_27255,N_27217);
and U27931 (N_27931,N_27034,N_27179);
or U27932 (N_27932,N_27326,N_27342);
and U27933 (N_27933,N_27152,N_27272);
or U27934 (N_27934,N_27224,N_27244);
xnor U27935 (N_27935,N_27181,N_27028);
nor U27936 (N_27936,N_27097,N_27258);
and U27937 (N_27937,N_27105,N_27229);
nor U27938 (N_27938,N_27030,N_27134);
or U27939 (N_27939,N_27015,N_27363);
nor U27940 (N_27940,N_27268,N_27143);
nand U27941 (N_27941,N_27008,N_27130);
and U27942 (N_27942,N_27136,N_27269);
nand U27943 (N_27943,N_27495,N_27022);
nor U27944 (N_27944,N_27179,N_27352);
nand U27945 (N_27945,N_27150,N_27303);
xor U27946 (N_27946,N_27067,N_27317);
xor U27947 (N_27947,N_27335,N_27129);
or U27948 (N_27948,N_27090,N_27311);
nor U27949 (N_27949,N_27304,N_27424);
nand U27950 (N_27950,N_27394,N_27070);
nor U27951 (N_27951,N_27242,N_27218);
nor U27952 (N_27952,N_27442,N_27065);
nor U27953 (N_27953,N_27127,N_27139);
and U27954 (N_27954,N_27101,N_27163);
nor U27955 (N_27955,N_27242,N_27283);
or U27956 (N_27956,N_27392,N_27165);
or U27957 (N_27957,N_27128,N_27237);
nor U27958 (N_27958,N_27034,N_27184);
nand U27959 (N_27959,N_27073,N_27244);
and U27960 (N_27960,N_27053,N_27125);
nor U27961 (N_27961,N_27318,N_27188);
nand U27962 (N_27962,N_27356,N_27009);
and U27963 (N_27963,N_27202,N_27158);
or U27964 (N_27964,N_27116,N_27242);
nand U27965 (N_27965,N_27147,N_27139);
and U27966 (N_27966,N_27374,N_27343);
nor U27967 (N_27967,N_27271,N_27275);
nand U27968 (N_27968,N_27131,N_27393);
and U27969 (N_27969,N_27287,N_27062);
or U27970 (N_27970,N_27433,N_27133);
and U27971 (N_27971,N_27071,N_27060);
or U27972 (N_27972,N_27462,N_27480);
nand U27973 (N_27973,N_27342,N_27048);
nor U27974 (N_27974,N_27340,N_27499);
or U27975 (N_27975,N_27226,N_27004);
nand U27976 (N_27976,N_27470,N_27319);
and U27977 (N_27977,N_27053,N_27039);
nor U27978 (N_27978,N_27365,N_27262);
nand U27979 (N_27979,N_27425,N_27088);
nand U27980 (N_27980,N_27269,N_27383);
nor U27981 (N_27981,N_27201,N_27077);
or U27982 (N_27982,N_27327,N_27092);
xnor U27983 (N_27983,N_27040,N_27059);
and U27984 (N_27984,N_27257,N_27011);
nor U27985 (N_27985,N_27125,N_27318);
or U27986 (N_27986,N_27230,N_27240);
nor U27987 (N_27987,N_27251,N_27265);
or U27988 (N_27988,N_27084,N_27493);
or U27989 (N_27989,N_27166,N_27455);
xor U27990 (N_27990,N_27306,N_27469);
and U27991 (N_27991,N_27276,N_27230);
xnor U27992 (N_27992,N_27000,N_27056);
or U27993 (N_27993,N_27048,N_27170);
nand U27994 (N_27994,N_27233,N_27164);
nand U27995 (N_27995,N_27160,N_27100);
or U27996 (N_27996,N_27372,N_27121);
or U27997 (N_27997,N_27376,N_27284);
nand U27998 (N_27998,N_27083,N_27277);
and U27999 (N_27999,N_27187,N_27271);
xor U28000 (N_28000,N_27976,N_27558);
nor U28001 (N_28001,N_27817,N_27864);
nand U28002 (N_28002,N_27823,N_27839);
and U28003 (N_28003,N_27614,N_27527);
and U28004 (N_28004,N_27835,N_27623);
and U28005 (N_28005,N_27871,N_27962);
nand U28006 (N_28006,N_27844,N_27500);
nor U28007 (N_28007,N_27521,N_27607);
xnor U28008 (N_28008,N_27855,N_27984);
nor U28009 (N_28009,N_27541,N_27951);
or U28010 (N_28010,N_27783,N_27529);
nor U28011 (N_28011,N_27751,N_27767);
nand U28012 (N_28012,N_27795,N_27760);
or U28013 (N_28013,N_27909,N_27849);
and U28014 (N_28014,N_27780,N_27757);
xor U28015 (N_28015,N_27724,N_27756);
or U28016 (N_28016,N_27803,N_27603);
nand U28017 (N_28017,N_27716,N_27714);
and U28018 (N_28018,N_27519,N_27938);
nand U28019 (N_28019,N_27690,N_27738);
or U28020 (N_28020,N_27890,N_27931);
nor U28021 (N_28021,N_27547,N_27761);
or U28022 (N_28022,N_27967,N_27704);
or U28023 (N_28023,N_27677,N_27619);
xnor U28024 (N_28024,N_27867,N_27902);
xor U28025 (N_28025,N_27509,N_27635);
or U28026 (N_28026,N_27634,N_27748);
nor U28027 (N_28027,N_27678,N_27566);
nor U28028 (N_28028,N_27671,N_27622);
or U28029 (N_28029,N_27964,N_27605);
nor U28030 (N_28030,N_27950,N_27514);
and U28031 (N_28031,N_27977,N_27667);
nand U28032 (N_28032,N_27752,N_27824);
or U28033 (N_28033,N_27560,N_27779);
nand U28034 (N_28034,N_27926,N_27991);
xor U28035 (N_28035,N_27801,N_27765);
and U28036 (N_28036,N_27569,N_27762);
and U28037 (N_28037,N_27654,N_27978);
nor U28038 (N_28038,N_27775,N_27531);
nand U28039 (N_28039,N_27524,N_27778);
or U28040 (N_28040,N_27729,N_27737);
nor U28041 (N_28041,N_27682,N_27829);
and U28042 (N_28042,N_27787,N_27980);
and U28043 (N_28043,N_27518,N_27968);
xor U28044 (N_28044,N_27631,N_27916);
xor U28045 (N_28045,N_27670,N_27853);
and U28046 (N_28046,N_27505,N_27847);
or U28047 (N_28047,N_27565,N_27639);
xor U28048 (N_28048,N_27673,N_27656);
nor U28049 (N_28049,N_27741,N_27895);
nand U28050 (N_28050,N_27593,N_27579);
nor U28051 (N_28051,N_27574,N_27810);
or U28052 (N_28052,N_27963,N_27989);
or U28053 (N_28053,N_27905,N_27731);
and U28054 (N_28054,N_27982,N_27646);
or U28055 (N_28055,N_27537,N_27929);
and U28056 (N_28056,N_27675,N_27845);
nand U28057 (N_28057,N_27821,N_27684);
or U28058 (N_28058,N_27986,N_27502);
nor U28059 (N_28059,N_27702,N_27655);
and U28060 (N_28060,N_27552,N_27814);
or U28061 (N_28061,N_27893,N_27770);
or U28062 (N_28062,N_27686,N_27640);
nor U28063 (N_28063,N_27557,N_27597);
and U28064 (N_28064,N_27504,N_27973);
xnor U28065 (N_28065,N_27936,N_27674);
nor U28066 (N_28066,N_27696,N_27993);
nand U28067 (N_28067,N_27570,N_27587);
or U28068 (N_28068,N_27854,N_27862);
nor U28069 (N_28069,N_27934,N_27992);
or U28070 (N_28070,N_27930,N_27754);
or U28071 (N_28071,N_27617,N_27694);
and U28072 (N_28072,N_27651,N_27881);
and U28073 (N_28073,N_27961,N_27740);
nand U28074 (N_28074,N_27918,N_27739);
or U28075 (N_28075,N_27753,N_27959);
nor U28076 (N_28076,N_27663,N_27523);
nor U28077 (N_28077,N_27685,N_27517);
and U28078 (N_28078,N_27556,N_27712);
or U28079 (N_28079,N_27925,N_27653);
and U28080 (N_28080,N_27588,N_27589);
and U28081 (N_28081,N_27596,N_27990);
nand U28082 (N_28082,N_27979,N_27723);
and U28083 (N_28083,N_27793,N_27915);
or U28084 (N_28084,N_27911,N_27535);
nor U28085 (N_28085,N_27609,N_27534);
or U28086 (N_28086,N_27940,N_27553);
nand U28087 (N_28087,N_27530,N_27710);
nand U28088 (N_28088,N_27953,N_27896);
nor U28089 (N_28089,N_27841,N_27863);
nand U28090 (N_28090,N_27742,N_27550);
nand U28091 (N_28091,N_27734,N_27618);
nor U28092 (N_28092,N_27861,N_27647);
and U28093 (N_28093,N_27781,N_27797);
nor U28094 (N_28094,N_27875,N_27981);
nand U28095 (N_28095,N_27876,N_27826);
nor U28096 (N_28096,N_27573,N_27620);
or U28097 (N_28097,N_27818,N_27580);
xnor U28098 (N_28098,N_27621,N_27600);
or U28099 (N_28099,N_27644,N_27768);
nor U28100 (N_28100,N_27727,N_27726);
or U28101 (N_28101,N_27827,N_27695);
nor U28102 (N_28102,N_27660,N_27626);
or U28103 (N_28103,N_27718,N_27539);
nor U28104 (N_28104,N_27608,N_27822);
nor U28105 (N_28105,N_27939,N_27616);
nand U28106 (N_28106,N_27949,N_27882);
nor U28107 (N_28107,N_27825,N_27544);
and U28108 (N_28108,N_27944,N_27883);
or U28109 (N_28109,N_27503,N_27657);
nor U28110 (N_28110,N_27528,N_27860);
nor U28111 (N_28111,N_27516,N_27869);
and U28112 (N_28112,N_27561,N_27628);
xor U28113 (N_28113,N_27804,N_27679);
and U28114 (N_28114,N_27791,N_27585);
xnor U28115 (N_28115,N_27652,N_27711);
or U28116 (N_28116,N_27586,N_27919);
nand U28117 (N_28117,N_27549,N_27923);
nand U28118 (N_28118,N_27928,N_27763);
nand U28119 (N_28119,N_27636,N_27637);
and U28120 (N_28120,N_27615,N_27820);
nand U28121 (N_28121,N_27999,N_27955);
nand U28122 (N_28122,N_27747,N_27945);
or U28123 (N_28123,N_27515,N_27551);
or U28124 (N_28124,N_27785,N_27725);
nand U28125 (N_28125,N_27813,N_27758);
or U28126 (N_28126,N_27645,N_27717);
nor U28127 (N_28127,N_27733,N_27922);
and U28128 (N_28128,N_27613,N_27567);
or U28129 (N_28129,N_27513,N_27611);
nor U28130 (N_28130,N_27970,N_27848);
nor U28131 (N_28131,N_27691,N_27800);
nand U28132 (N_28132,N_27538,N_27601);
or U28133 (N_28133,N_27598,N_27831);
nand U28134 (N_28134,N_27536,N_27836);
nand U28135 (N_28135,N_27721,N_27746);
and U28136 (N_28136,N_27811,N_27735);
nand U28137 (N_28137,N_27946,N_27624);
nor U28138 (N_28138,N_27599,N_27759);
nand U28139 (N_28139,N_27815,N_27892);
or U28140 (N_28140,N_27947,N_27577);
nand U28141 (N_28141,N_27998,N_27769);
nor U28142 (N_28142,N_27957,N_27920);
and U28143 (N_28143,N_27901,N_27857);
xor U28144 (N_28144,N_27546,N_27590);
nor U28145 (N_28145,N_27559,N_27943);
or U28146 (N_28146,N_27545,N_27886);
or U28147 (N_28147,N_27865,N_27856);
or U28148 (N_28148,N_27850,N_27720);
and U28149 (N_28149,N_27766,N_27809);
and U28150 (N_28150,N_27958,N_27948);
and U28151 (N_28151,N_27868,N_27879);
nor U28152 (N_28152,N_27969,N_27563);
or U28153 (N_28153,N_27507,N_27576);
and U28154 (N_28154,N_27708,N_27927);
and U28155 (N_28155,N_27894,N_27917);
or U28156 (N_28156,N_27555,N_27744);
or U28157 (N_28157,N_27807,N_27533);
or U28158 (N_28158,N_27907,N_27707);
nor U28159 (N_28159,N_27812,N_27884);
and U28160 (N_28160,N_27838,N_27806);
nor U28161 (N_28161,N_27833,N_27642);
nand U28162 (N_28162,N_27680,N_27832);
or U28163 (N_28163,N_27952,N_27932);
and U28164 (N_28164,N_27776,N_27912);
or U28165 (N_28165,N_27796,N_27974);
and U28166 (N_28166,N_27575,N_27885);
and U28167 (N_28167,N_27942,N_27520);
and U28168 (N_28168,N_27699,N_27782);
or U28169 (N_28169,N_27698,N_27828);
nor U28170 (N_28170,N_27543,N_27641);
nor U28171 (N_28171,N_27996,N_27542);
or U28172 (N_28172,N_27995,N_27910);
nor U28173 (N_28173,N_27512,N_27819);
or U28174 (N_28174,N_27786,N_27564);
nor U28175 (N_28175,N_27629,N_27956);
and U28176 (N_28176,N_27852,N_27899);
nand U28177 (N_28177,N_27887,N_27914);
or U28178 (N_28178,N_27594,N_27501);
or U28179 (N_28179,N_27802,N_27692);
or U28180 (N_28180,N_27706,N_27562);
or U28181 (N_28181,N_27681,N_27526);
nor U28182 (N_28182,N_27921,N_27506);
nor U28183 (N_28183,N_27591,N_27701);
nand U28184 (N_28184,N_27532,N_27630);
and U28185 (N_28185,N_27592,N_27571);
and U28186 (N_28186,N_27960,N_27997);
or U28187 (N_28187,N_27777,N_27870);
nand U28188 (N_28188,N_27935,N_27662);
xor U28189 (N_28189,N_27830,N_27703);
or U28190 (N_28190,N_27966,N_27937);
xor U28191 (N_28191,N_27625,N_27846);
nand U28192 (N_28192,N_27985,N_27627);
or U28193 (N_28193,N_27908,N_27578);
xnor U28194 (N_28194,N_27750,N_27858);
nor U28195 (N_28195,N_27941,N_27843);
or U28196 (N_28196,N_27730,N_27683);
and U28197 (N_28197,N_27602,N_27799);
nor U28198 (N_28198,N_27650,N_27745);
nand U28199 (N_28199,N_27665,N_27595);
and U28200 (N_28200,N_27643,N_27773);
or U28201 (N_28201,N_27715,N_27668);
nand U28202 (N_28202,N_27792,N_27888);
nor U28203 (N_28203,N_27584,N_27971);
or U28204 (N_28204,N_27900,N_27736);
nand U28205 (N_28205,N_27872,N_27612);
or U28206 (N_28206,N_27764,N_27722);
nor U28207 (N_28207,N_27851,N_27664);
or U28208 (N_28208,N_27994,N_27661);
and U28209 (N_28209,N_27889,N_27859);
or U28210 (N_28210,N_27913,N_27891);
or U28211 (N_28211,N_27583,N_27878);
or U28212 (N_28212,N_27897,N_27713);
and U28213 (N_28213,N_27700,N_27784);
nor U28214 (N_28214,N_27688,N_27522);
nor U28215 (N_28215,N_27693,N_27808);
nor U28216 (N_28216,N_27749,N_27508);
nand U28217 (N_28217,N_27772,N_27816);
and U28218 (N_28218,N_27604,N_27898);
or U28219 (N_28219,N_27610,N_27511);
and U28220 (N_28220,N_27548,N_27774);
or U28221 (N_28221,N_27648,N_27697);
and U28222 (N_28222,N_27771,N_27790);
or U28223 (N_28223,N_27906,N_27719);
nor U28224 (N_28224,N_27842,N_27873);
or U28225 (N_28225,N_27705,N_27554);
nand U28226 (N_28226,N_27988,N_27743);
nand U28227 (N_28227,N_27877,N_27638);
nor U28228 (N_28228,N_27649,N_27568);
nor U28229 (N_28229,N_27666,N_27633);
or U28230 (N_28230,N_27972,N_27904);
and U28231 (N_28231,N_27755,N_27709);
nor U28232 (N_28232,N_27965,N_27606);
nor U28233 (N_28233,N_27880,N_27903);
nor U28234 (N_28234,N_27954,N_27728);
and U28235 (N_28235,N_27987,N_27510);
nand U28236 (N_28236,N_27676,N_27540);
nor U28237 (N_28237,N_27789,N_27659);
nor U28238 (N_28238,N_27732,N_27689);
xor U28239 (N_28239,N_27983,N_27874);
nand U28240 (N_28240,N_27866,N_27581);
or U28241 (N_28241,N_27798,N_27840);
nand U28242 (N_28242,N_27788,N_27632);
nand U28243 (N_28243,N_27658,N_27924);
nand U28244 (N_28244,N_27669,N_27834);
nand U28245 (N_28245,N_27933,N_27572);
or U28246 (N_28246,N_27687,N_27975);
nor U28247 (N_28247,N_27672,N_27837);
xor U28248 (N_28248,N_27794,N_27525);
or U28249 (N_28249,N_27582,N_27805);
nand U28250 (N_28250,N_27942,N_27771);
nand U28251 (N_28251,N_27897,N_27736);
and U28252 (N_28252,N_27915,N_27739);
nor U28253 (N_28253,N_27920,N_27686);
and U28254 (N_28254,N_27516,N_27865);
or U28255 (N_28255,N_27984,N_27679);
and U28256 (N_28256,N_27743,N_27538);
nor U28257 (N_28257,N_27613,N_27651);
and U28258 (N_28258,N_27777,N_27771);
nand U28259 (N_28259,N_27615,N_27945);
and U28260 (N_28260,N_27623,N_27979);
nor U28261 (N_28261,N_27955,N_27549);
or U28262 (N_28262,N_27606,N_27962);
nor U28263 (N_28263,N_27779,N_27889);
nor U28264 (N_28264,N_27502,N_27845);
or U28265 (N_28265,N_27952,N_27769);
or U28266 (N_28266,N_27516,N_27569);
nand U28267 (N_28267,N_27772,N_27567);
or U28268 (N_28268,N_27571,N_27757);
or U28269 (N_28269,N_27626,N_27896);
nand U28270 (N_28270,N_27620,N_27537);
nand U28271 (N_28271,N_27536,N_27784);
nor U28272 (N_28272,N_27756,N_27581);
or U28273 (N_28273,N_27959,N_27775);
or U28274 (N_28274,N_27790,N_27882);
or U28275 (N_28275,N_27936,N_27726);
nand U28276 (N_28276,N_27532,N_27599);
or U28277 (N_28277,N_27766,N_27660);
or U28278 (N_28278,N_27733,N_27818);
nor U28279 (N_28279,N_27805,N_27594);
nor U28280 (N_28280,N_27790,N_27508);
nor U28281 (N_28281,N_27658,N_27586);
nor U28282 (N_28282,N_27733,N_27638);
nand U28283 (N_28283,N_27659,N_27861);
nand U28284 (N_28284,N_27779,N_27628);
or U28285 (N_28285,N_27999,N_27508);
or U28286 (N_28286,N_27954,N_27630);
or U28287 (N_28287,N_27834,N_27611);
and U28288 (N_28288,N_27717,N_27840);
nor U28289 (N_28289,N_27861,N_27968);
or U28290 (N_28290,N_27801,N_27610);
or U28291 (N_28291,N_27813,N_27566);
nor U28292 (N_28292,N_27653,N_27619);
or U28293 (N_28293,N_27544,N_27827);
nor U28294 (N_28294,N_27637,N_27784);
or U28295 (N_28295,N_27742,N_27881);
nand U28296 (N_28296,N_27839,N_27534);
or U28297 (N_28297,N_27685,N_27670);
nor U28298 (N_28298,N_27800,N_27876);
nand U28299 (N_28299,N_27510,N_27591);
nand U28300 (N_28300,N_27852,N_27627);
or U28301 (N_28301,N_27616,N_27822);
and U28302 (N_28302,N_27579,N_27762);
or U28303 (N_28303,N_27700,N_27959);
nor U28304 (N_28304,N_27875,N_27988);
xnor U28305 (N_28305,N_27571,N_27840);
or U28306 (N_28306,N_27866,N_27655);
and U28307 (N_28307,N_27902,N_27535);
and U28308 (N_28308,N_27510,N_27913);
nand U28309 (N_28309,N_27579,N_27587);
nand U28310 (N_28310,N_27774,N_27891);
nand U28311 (N_28311,N_27701,N_27587);
nand U28312 (N_28312,N_27544,N_27501);
xor U28313 (N_28313,N_27536,N_27890);
nor U28314 (N_28314,N_27920,N_27628);
xnor U28315 (N_28315,N_27591,N_27670);
or U28316 (N_28316,N_27633,N_27848);
nand U28317 (N_28317,N_27554,N_27746);
xor U28318 (N_28318,N_27641,N_27581);
and U28319 (N_28319,N_27649,N_27910);
nand U28320 (N_28320,N_27825,N_27526);
nor U28321 (N_28321,N_27931,N_27667);
nor U28322 (N_28322,N_27552,N_27679);
nand U28323 (N_28323,N_27569,N_27680);
nand U28324 (N_28324,N_27858,N_27556);
nand U28325 (N_28325,N_27912,N_27933);
nor U28326 (N_28326,N_27742,N_27807);
or U28327 (N_28327,N_27716,N_27596);
or U28328 (N_28328,N_27509,N_27768);
or U28329 (N_28329,N_27978,N_27872);
and U28330 (N_28330,N_27874,N_27817);
nand U28331 (N_28331,N_27736,N_27725);
and U28332 (N_28332,N_27854,N_27703);
nand U28333 (N_28333,N_27604,N_27636);
or U28334 (N_28334,N_27910,N_27563);
and U28335 (N_28335,N_27963,N_27616);
nor U28336 (N_28336,N_27796,N_27903);
nor U28337 (N_28337,N_27501,N_27636);
and U28338 (N_28338,N_27768,N_27569);
or U28339 (N_28339,N_27686,N_27930);
or U28340 (N_28340,N_27732,N_27616);
nand U28341 (N_28341,N_27940,N_27734);
xnor U28342 (N_28342,N_27510,N_27511);
nor U28343 (N_28343,N_27734,N_27939);
or U28344 (N_28344,N_27913,N_27529);
or U28345 (N_28345,N_27860,N_27588);
nor U28346 (N_28346,N_27886,N_27555);
nor U28347 (N_28347,N_27863,N_27806);
nor U28348 (N_28348,N_27697,N_27643);
and U28349 (N_28349,N_27947,N_27855);
and U28350 (N_28350,N_27850,N_27938);
xor U28351 (N_28351,N_27825,N_27954);
or U28352 (N_28352,N_27844,N_27768);
and U28353 (N_28353,N_27875,N_27952);
nand U28354 (N_28354,N_27815,N_27645);
xor U28355 (N_28355,N_27751,N_27868);
or U28356 (N_28356,N_27766,N_27593);
xor U28357 (N_28357,N_27892,N_27501);
or U28358 (N_28358,N_27661,N_27938);
nand U28359 (N_28359,N_27594,N_27616);
nand U28360 (N_28360,N_27676,N_27634);
nand U28361 (N_28361,N_27773,N_27977);
or U28362 (N_28362,N_27863,N_27939);
xnor U28363 (N_28363,N_27596,N_27962);
nand U28364 (N_28364,N_27559,N_27862);
nand U28365 (N_28365,N_27548,N_27585);
and U28366 (N_28366,N_27942,N_27698);
nor U28367 (N_28367,N_27902,N_27690);
nor U28368 (N_28368,N_27731,N_27885);
xor U28369 (N_28369,N_27891,N_27927);
or U28370 (N_28370,N_27562,N_27737);
xor U28371 (N_28371,N_27765,N_27684);
nand U28372 (N_28372,N_27702,N_27507);
nor U28373 (N_28373,N_27879,N_27884);
nor U28374 (N_28374,N_27876,N_27676);
nand U28375 (N_28375,N_27836,N_27568);
and U28376 (N_28376,N_27728,N_27612);
nor U28377 (N_28377,N_27673,N_27682);
and U28378 (N_28378,N_27752,N_27732);
nor U28379 (N_28379,N_27933,N_27923);
or U28380 (N_28380,N_27908,N_27599);
nor U28381 (N_28381,N_27932,N_27556);
nand U28382 (N_28382,N_27530,N_27954);
nor U28383 (N_28383,N_27972,N_27583);
xnor U28384 (N_28384,N_27629,N_27895);
or U28385 (N_28385,N_27880,N_27942);
and U28386 (N_28386,N_27980,N_27763);
xor U28387 (N_28387,N_27535,N_27687);
nand U28388 (N_28388,N_27873,N_27619);
nor U28389 (N_28389,N_27795,N_27989);
and U28390 (N_28390,N_27589,N_27950);
nand U28391 (N_28391,N_27578,N_27966);
xnor U28392 (N_28392,N_27644,N_27706);
and U28393 (N_28393,N_27754,N_27849);
and U28394 (N_28394,N_27553,N_27895);
nand U28395 (N_28395,N_27785,N_27933);
nor U28396 (N_28396,N_27535,N_27996);
nor U28397 (N_28397,N_27540,N_27955);
nand U28398 (N_28398,N_27643,N_27692);
and U28399 (N_28399,N_27901,N_27609);
xor U28400 (N_28400,N_27521,N_27760);
nor U28401 (N_28401,N_27574,N_27611);
xor U28402 (N_28402,N_27798,N_27647);
and U28403 (N_28403,N_27907,N_27725);
xnor U28404 (N_28404,N_27780,N_27812);
nand U28405 (N_28405,N_27780,N_27789);
nand U28406 (N_28406,N_27962,N_27935);
nor U28407 (N_28407,N_27584,N_27986);
nand U28408 (N_28408,N_27998,N_27784);
nand U28409 (N_28409,N_27689,N_27518);
or U28410 (N_28410,N_27792,N_27683);
nand U28411 (N_28411,N_27875,N_27612);
or U28412 (N_28412,N_27509,N_27837);
nor U28413 (N_28413,N_27917,N_27790);
nor U28414 (N_28414,N_27562,N_27623);
or U28415 (N_28415,N_27908,N_27992);
or U28416 (N_28416,N_27960,N_27810);
or U28417 (N_28417,N_27733,N_27612);
nor U28418 (N_28418,N_27776,N_27640);
and U28419 (N_28419,N_27956,N_27841);
nor U28420 (N_28420,N_27678,N_27897);
and U28421 (N_28421,N_27837,N_27612);
or U28422 (N_28422,N_27893,N_27806);
nor U28423 (N_28423,N_27614,N_27572);
nor U28424 (N_28424,N_27625,N_27728);
or U28425 (N_28425,N_27642,N_27608);
nand U28426 (N_28426,N_27934,N_27733);
and U28427 (N_28427,N_27754,N_27590);
nand U28428 (N_28428,N_27774,N_27814);
nand U28429 (N_28429,N_27805,N_27967);
xor U28430 (N_28430,N_27899,N_27888);
and U28431 (N_28431,N_27953,N_27779);
and U28432 (N_28432,N_27856,N_27832);
or U28433 (N_28433,N_27628,N_27830);
and U28434 (N_28434,N_27700,N_27695);
and U28435 (N_28435,N_27524,N_27690);
and U28436 (N_28436,N_27723,N_27779);
nor U28437 (N_28437,N_27651,N_27513);
xor U28438 (N_28438,N_27533,N_27603);
nor U28439 (N_28439,N_27587,N_27591);
nand U28440 (N_28440,N_27984,N_27838);
nor U28441 (N_28441,N_27584,N_27793);
and U28442 (N_28442,N_27609,N_27886);
and U28443 (N_28443,N_27939,N_27930);
or U28444 (N_28444,N_27975,N_27972);
nor U28445 (N_28445,N_27589,N_27518);
nor U28446 (N_28446,N_27650,N_27736);
nand U28447 (N_28447,N_27598,N_27520);
or U28448 (N_28448,N_27846,N_27575);
xnor U28449 (N_28449,N_27750,N_27669);
and U28450 (N_28450,N_27719,N_27978);
or U28451 (N_28451,N_27935,N_27606);
or U28452 (N_28452,N_27530,N_27619);
nor U28453 (N_28453,N_27968,N_27952);
or U28454 (N_28454,N_27718,N_27729);
or U28455 (N_28455,N_27850,N_27825);
and U28456 (N_28456,N_27834,N_27623);
and U28457 (N_28457,N_27760,N_27715);
nor U28458 (N_28458,N_27806,N_27999);
and U28459 (N_28459,N_27534,N_27828);
or U28460 (N_28460,N_27803,N_27697);
and U28461 (N_28461,N_27558,N_27752);
and U28462 (N_28462,N_27597,N_27763);
or U28463 (N_28463,N_27826,N_27601);
or U28464 (N_28464,N_27561,N_27853);
and U28465 (N_28465,N_27851,N_27523);
or U28466 (N_28466,N_27544,N_27618);
and U28467 (N_28467,N_27983,N_27608);
nor U28468 (N_28468,N_27912,N_27881);
and U28469 (N_28469,N_27859,N_27671);
and U28470 (N_28470,N_27824,N_27997);
and U28471 (N_28471,N_27596,N_27819);
or U28472 (N_28472,N_27559,N_27663);
or U28473 (N_28473,N_27878,N_27818);
and U28474 (N_28474,N_27824,N_27678);
nand U28475 (N_28475,N_27617,N_27560);
nor U28476 (N_28476,N_27901,N_27929);
and U28477 (N_28477,N_27991,N_27884);
xor U28478 (N_28478,N_27642,N_27721);
nand U28479 (N_28479,N_27848,N_27727);
nand U28480 (N_28480,N_27845,N_27745);
nand U28481 (N_28481,N_27579,N_27975);
nor U28482 (N_28482,N_27827,N_27664);
nand U28483 (N_28483,N_27790,N_27763);
nor U28484 (N_28484,N_27861,N_27579);
nor U28485 (N_28485,N_27911,N_27898);
and U28486 (N_28486,N_27980,N_27666);
and U28487 (N_28487,N_27566,N_27510);
and U28488 (N_28488,N_27856,N_27516);
nor U28489 (N_28489,N_27693,N_27870);
nor U28490 (N_28490,N_27962,N_27902);
nor U28491 (N_28491,N_27506,N_27969);
xor U28492 (N_28492,N_27632,N_27982);
and U28493 (N_28493,N_27744,N_27530);
and U28494 (N_28494,N_27739,N_27623);
nand U28495 (N_28495,N_27643,N_27802);
nand U28496 (N_28496,N_27910,N_27534);
or U28497 (N_28497,N_27508,N_27563);
nand U28498 (N_28498,N_27894,N_27815);
nand U28499 (N_28499,N_27572,N_27528);
or U28500 (N_28500,N_28492,N_28285);
nand U28501 (N_28501,N_28410,N_28240);
or U28502 (N_28502,N_28489,N_28397);
nand U28503 (N_28503,N_28278,N_28050);
and U28504 (N_28504,N_28399,N_28252);
or U28505 (N_28505,N_28407,N_28173);
nor U28506 (N_28506,N_28193,N_28010);
and U28507 (N_28507,N_28080,N_28154);
nor U28508 (N_28508,N_28257,N_28148);
or U28509 (N_28509,N_28333,N_28431);
or U28510 (N_28510,N_28265,N_28079);
or U28511 (N_28511,N_28022,N_28027);
xnor U28512 (N_28512,N_28018,N_28174);
nand U28513 (N_28513,N_28189,N_28415);
or U28514 (N_28514,N_28029,N_28023);
or U28515 (N_28515,N_28056,N_28307);
or U28516 (N_28516,N_28336,N_28344);
xor U28517 (N_28517,N_28479,N_28171);
xnor U28518 (N_28518,N_28038,N_28209);
nand U28519 (N_28519,N_28380,N_28368);
nand U28520 (N_28520,N_28314,N_28065);
and U28521 (N_28521,N_28256,N_28087);
or U28522 (N_28522,N_28076,N_28367);
nor U28523 (N_28523,N_28444,N_28082);
and U28524 (N_28524,N_28453,N_28205);
nor U28525 (N_28525,N_28284,N_28261);
and U28526 (N_28526,N_28213,N_28101);
or U28527 (N_28527,N_28329,N_28192);
nor U28528 (N_28528,N_28390,N_28150);
xor U28529 (N_28529,N_28125,N_28127);
and U28530 (N_28530,N_28179,N_28136);
and U28531 (N_28531,N_28411,N_28019);
nor U28532 (N_28532,N_28001,N_28139);
nor U28533 (N_28533,N_28498,N_28325);
nor U28534 (N_28534,N_28129,N_28300);
or U28535 (N_28535,N_28230,N_28147);
and U28536 (N_28536,N_28194,N_28096);
nand U28537 (N_28537,N_28327,N_28398);
xor U28538 (N_28538,N_28042,N_28310);
or U28539 (N_28539,N_28451,N_28374);
nand U28540 (N_28540,N_28334,N_28035);
nor U28541 (N_28541,N_28346,N_28468);
or U28542 (N_28542,N_28402,N_28359);
or U28543 (N_28543,N_28475,N_28033);
and U28544 (N_28544,N_28476,N_28248);
nand U28545 (N_28545,N_28465,N_28236);
nand U28546 (N_28546,N_28447,N_28370);
nand U28547 (N_28547,N_28461,N_28424);
and U28548 (N_28548,N_28088,N_28323);
nor U28549 (N_28549,N_28316,N_28083);
nor U28550 (N_28550,N_28055,N_28481);
or U28551 (N_28551,N_28024,N_28073);
nor U28552 (N_28552,N_28051,N_28124);
and U28553 (N_28553,N_28181,N_28164);
and U28554 (N_28554,N_28190,N_28132);
or U28555 (N_28555,N_28490,N_28384);
and U28556 (N_28556,N_28483,N_28058);
xor U28557 (N_28557,N_28199,N_28007);
and U28558 (N_28558,N_28090,N_28470);
nor U28559 (N_28559,N_28028,N_28456);
or U28560 (N_28560,N_28195,N_28393);
nand U28561 (N_28561,N_28288,N_28432);
nor U28562 (N_28562,N_28341,N_28255);
or U28563 (N_28563,N_28435,N_28228);
or U28564 (N_28564,N_28302,N_28304);
nand U28565 (N_28565,N_28178,N_28214);
xor U28566 (N_28566,N_28419,N_28141);
nand U28567 (N_28567,N_28246,N_28176);
nor U28568 (N_28568,N_28168,N_28363);
or U28569 (N_28569,N_28482,N_28471);
and U28570 (N_28570,N_28420,N_28259);
nor U28571 (N_28571,N_28108,N_28006);
and U28572 (N_28572,N_28045,N_28268);
nor U28573 (N_28573,N_28440,N_28392);
nor U28574 (N_28574,N_28070,N_28005);
nand U28575 (N_28575,N_28446,N_28123);
nor U28576 (N_28576,N_28182,N_28460);
xnor U28577 (N_28577,N_28169,N_28060);
nand U28578 (N_28578,N_28091,N_28237);
or U28579 (N_28579,N_28075,N_28478);
or U28580 (N_28580,N_28339,N_28250);
nand U28581 (N_28581,N_28383,N_28115);
or U28582 (N_28582,N_28499,N_28217);
and U28583 (N_28583,N_28021,N_28280);
nand U28584 (N_28584,N_28494,N_28200);
nand U28585 (N_28585,N_28202,N_28296);
nand U28586 (N_28586,N_28305,N_28436);
and U28587 (N_28587,N_28328,N_28251);
and U28588 (N_28588,N_28098,N_28198);
nor U28589 (N_28589,N_28409,N_28442);
and U28590 (N_28590,N_28289,N_28238);
or U28591 (N_28591,N_28116,N_28121);
xnor U28592 (N_28592,N_28216,N_28002);
or U28593 (N_28593,N_28474,N_28464);
nand U28594 (N_28594,N_28000,N_28275);
or U28595 (N_28595,N_28269,N_28286);
and U28596 (N_28596,N_28496,N_28351);
xor U28597 (N_28597,N_28375,N_28331);
and U28598 (N_28598,N_28040,N_28340);
nand U28599 (N_28599,N_28235,N_28381);
nand U28600 (N_28600,N_28247,N_28163);
and U28601 (N_28601,N_28077,N_28074);
xnor U28602 (N_28602,N_28473,N_28356);
xor U28603 (N_28603,N_28271,N_28158);
and U28604 (N_28604,N_28321,N_28072);
nand U28605 (N_28605,N_28320,N_28396);
xor U28606 (N_28606,N_28308,N_28379);
and U28607 (N_28607,N_28239,N_28353);
nor U28608 (N_28608,N_28231,N_28264);
nand U28609 (N_28609,N_28137,N_28354);
and U28610 (N_28610,N_28242,N_28153);
or U28611 (N_28611,N_28241,N_28488);
or U28612 (N_28612,N_28061,N_28089);
and U28613 (N_28613,N_28343,N_28317);
and U28614 (N_28614,N_28282,N_28012);
and U28615 (N_28615,N_28034,N_28400);
and U28616 (N_28616,N_28497,N_28130);
nand U28617 (N_28617,N_28480,N_28207);
nor U28618 (N_28618,N_28262,N_28416);
nor U28619 (N_28619,N_28225,N_28011);
nand U28620 (N_28620,N_28218,N_28454);
nor U28621 (N_28621,N_28263,N_28360);
or U28622 (N_28622,N_28401,N_28149);
nor U28623 (N_28623,N_28313,N_28113);
nand U28624 (N_28624,N_28388,N_28165);
nand U28625 (N_28625,N_28175,N_28043);
and U28626 (N_28626,N_28326,N_28430);
or U28627 (N_28627,N_28106,N_28233);
nand U28628 (N_28628,N_28063,N_28303);
or U28629 (N_28629,N_28365,N_28413);
nor U28630 (N_28630,N_28078,N_28185);
or U28631 (N_28631,N_28391,N_28142);
and U28632 (N_28632,N_28421,N_28276);
xnor U28633 (N_28633,N_28166,N_28159);
or U28634 (N_28634,N_28274,N_28290);
and U28635 (N_28635,N_28270,N_28345);
nor U28636 (N_28636,N_28441,N_28099);
nor U28637 (N_28637,N_28445,N_28428);
nor U28638 (N_28638,N_28036,N_28120);
xor U28639 (N_28639,N_28016,N_28203);
and U28640 (N_28640,N_28459,N_28423);
and U28641 (N_28641,N_28003,N_28462);
nor U28642 (N_28642,N_28057,N_28352);
nor U28643 (N_28643,N_28162,N_28466);
and U28644 (N_28644,N_28103,N_28092);
nor U28645 (N_28645,N_28467,N_28366);
nand U28646 (N_28646,N_28220,N_28067);
nand U28647 (N_28647,N_28348,N_28105);
or U28648 (N_28648,N_28052,N_28102);
and U28649 (N_28649,N_28094,N_28350);
nor U28650 (N_28650,N_28046,N_28114);
and U28651 (N_28651,N_28201,N_28439);
nor U28652 (N_28652,N_28491,N_28287);
nand U28653 (N_28653,N_28244,N_28186);
or U28654 (N_28654,N_28143,N_28294);
nor U28655 (N_28655,N_28319,N_28293);
nand U28656 (N_28656,N_28039,N_28206);
and U28657 (N_28657,N_28311,N_28484);
nand U28658 (N_28658,N_28272,N_28020);
nor U28659 (N_28659,N_28188,N_28364);
and U28660 (N_28660,N_28455,N_28306);
nor U28661 (N_28661,N_28109,N_28229);
and U28662 (N_28662,N_28062,N_28371);
nand U28663 (N_28663,N_28254,N_28477);
nand U28664 (N_28664,N_28155,N_28232);
and U28665 (N_28665,N_28291,N_28133);
nor U28666 (N_28666,N_28463,N_28112);
nor U28667 (N_28667,N_28004,N_28032);
and U28668 (N_28668,N_28180,N_28427);
or U28669 (N_28669,N_28357,N_28119);
and U28670 (N_28670,N_28298,N_28361);
nor U28671 (N_28671,N_28406,N_28458);
nor U28672 (N_28672,N_28008,N_28448);
xor U28673 (N_28673,N_28118,N_28170);
nor U28674 (N_28674,N_28387,N_28197);
or U28675 (N_28675,N_28315,N_28223);
and U28676 (N_28676,N_28295,N_28131);
nor U28677 (N_28677,N_28085,N_28041);
or U28678 (N_28678,N_28013,N_28338);
nor U28679 (N_28679,N_28064,N_28349);
and U28680 (N_28680,N_28086,N_28243);
xor U28681 (N_28681,N_28335,N_28224);
nand U28682 (N_28682,N_28100,N_28157);
xor U28683 (N_28683,N_28245,N_28048);
nand U28684 (N_28684,N_28373,N_28324);
nand U28685 (N_28685,N_28187,N_28140);
nand U28686 (N_28686,N_28204,N_28309);
and U28687 (N_28687,N_28408,N_28412);
or U28688 (N_28688,N_28030,N_28128);
or U28689 (N_28689,N_28234,N_28267);
nor U28690 (N_28690,N_28025,N_28457);
or U28691 (N_28691,N_28281,N_28084);
nand U28692 (N_28692,N_28443,N_28208);
and U28693 (N_28693,N_28277,N_28044);
or U28694 (N_28694,N_28212,N_28167);
xnor U28695 (N_28695,N_28434,N_28226);
or U28696 (N_28696,N_28342,N_28219);
nand U28697 (N_28697,N_28081,N_28362);
nand U28698 (N_28698,N_28279,N_28015);
nand U28699 (N_28699,N_28332,N_28386);
and U28700 (N_28700,N_28196,N_28414);
or U28701 (N_28701,N_28376,N_28068);
xor U28702 (N_28702,N_28372,N_28172);
nand U28703 (N_28703,N_28297,N_28438);
nor U28704 (N_28704,N_28418,N_28404);
nor U28705 (N_28705,N_28151,N_28450);
xor U28706 (N_28706,N_28135,N_28227);
nor U28707 (N_28707,N_28210,N_28469);
xnor U28708 (N_28708,N_28292,N_28183);
nand U28709 (N_28709,N_28134,N_28395);
nor U28710 (N_28710,N_28066,N_28394);
and U28711 (N_28711,N_28337,N_28312);
nand U28712 (N_28712,N_28382,N_28385);
nor U28713 (N_28713,N_28184,N_28266);
nand U28714 (N_28714,N_28249,N_28253);
nor U28715 (N_28715,N_28433,N_28377);
and U28716 (N_28716,N_28258,N_28485);
nand U28717 (N_28717,N_28449,N_28322);
xnor U28718 (N_28718,N_28299,N_28495);
or U28719 (N_28719,N_28437,N_28152);
and U28720 (N_28720,N_28389,N_28425);
xor U28721 (N_28721,N_28037,N_28493);
xnor U28722 (N_28722,N_28472,N_28097);
and U28723 (N_28723,N_28378,N_28049);
nor U28724 (N_28724,N_28069,N_28059);
nand U28725 (N_28725,N_28177,N_28145);
nand U28726 (N_28726,N_28107,N_28031);
or U28727 (N_28727,N_28358,N_28487);
and U28728 (N_28728,N_28160,N_28009);
or U28729 (N_28729,N_28191,N_28221);
and U28730 (N_28730,N_28117,N_28126);
xor U28731 (N_28731,N_28095,N_28138);
nand U28732 (N_28732,N_28215,N_28403);
nor U28733 (N_28733,N_28047,N_28369);
and U28734 (N_28734,N_28054,N_28017);
nand U28735 (N_28735,N_28014,N_28452);
nor U28736 (N_28736,N_28417,N_28429);
or U28737 (N_28737,N_28405,N_28156);
or U28738 (N_28738,N_28161,N_28071);
nand U28739 (N_28739,N_28330,N_28110);
and U28740 (N_28740,N_28026,N_28422);
nand U28741 (N_28741,N_28273,N_28283);
and U28742 (N_28742,N_28211,N_28301);
nor U28743 (N_28743,N_28122,N_28260);
or U28744 (N_28744,N_28355,N_28144);
nand U28745 (N_28745,N_28222,N_28347);
nor U28746 (N_28746,N_28486,N_28318);
nand U28747 (N_28747,N_28426,N_28104);
nor U28748 (N_28748,N_28093,N_28053);
or U28749 (N_28749,N_28146,N_28111);
and U28750 (N_28750,N_28119,N_28218);
and U28751 (N_28751,N_28207,N_28431);
nor U28752 (N_28752,N_28195,N_28489);
and U28753 (N_28753,N_28471,N_28296);
or U28754 (N_28754,N_28328,N_28064);
and U28755 (N_28755,N_28031,N_28293);
and U28756 (N_28756,N_28462,N_28468);
and U28757 (N_28757,N_28344,N_28478);
xnor U28758 (N_28758,N_28168,N_28498);
or U28759 (N_28759,N_28049,N_28066);
nor U28760 (N_28760,N_28425,N_28326);
nand U28761 (N_28761,N_28336,N_28086);
nor U28762 (N_28762,N_28241,N_28229);
and U28763 (N_28763,N_28097,N_28468);
nor U28764 (N_28764,N_28181,N_28013);
and U28765 (N_28765,N_28228,N_28381);
and U28766 (N_28766,N_28496,N_28287);
xnor U28767 (N_28767,N_28153,N_28340);
nand U28768 (N_28768,N_28409,N_28089);
nor U28769 (N_28769,N_28277,N_28003);
or U28770 (N_28770,N_28294,N_28408);
and U28771 (N_28771,N_28342,N_28315);
or U28772 (N_28772,N_28286,N_28261);
nor U28773 (N_28773,N_28098,N_28112);
xnor U28774 (N_28774,N_28122,N_28231);
nor U28775 (N_28775,N_28379,N_28110);
and U28776 (N_28776,N_28285,N_28121);
or U28777 (N_28777,N_28222,N_28306);
xnor U28778 (N_28778,N_28312,N_28094);
and U28779 (N_28779,N_28010,N_28166);
nor U28780 (N_28780,N_28325,N_28190);
or U28781 (N_28781,N_28336,N_28493);
and U28782 (N_28782,N_28226,N_28218);
nor U28783 (N_28783,N_28452,N_28413);
nor U28784 (N_28784,N_28471,N_28019);
nor U28785 (N_28785,N_28132,N_28439);
and U28786 (N_28786,N_28054,N_28280);
and U28787 (N_28787,N_28469,N_28305);
nor U28788 (N_28788,N_28232,N_28319);
nand U28789 (N_28789,N_28162,N_28377);
or U28790 (N_28790,N_28079,N_28139);
nand U28791 (N_28791,N_28172,N_28151);
nand U28792 (N_28792,N_28104,N_28110);
xnor U28793 (N_28793,N_28320,N_28390);
nand U28794 (N_28794,N_28450,N_28396);
and U28795 (N_28795,N_28220,N_28009);
nor U28796 (N_28796,N_28343,N_28334);
nand U28797 (N_28797,N_28298,N_28273);
nand U28798 (N_28798,N_28170,N_28484);
or U28799 (N_28799,N_28307,N_28459);
nand U28800 (N_28800,N_28195,N_28378);
nor U28801 (N_28801,N_28280,N_28268);
nor U28802 (N_28802,N_28030,N_28404);
nand U28803 (N_28803,N_28387,N_28247);
nor U28804 (N_28804,N_28385,N_28271);
or U28805 (N_28805,N_28083,N_28085);
and U28806 (N_28806,N_28341,N_28006);
and U28807 (N_28807,N_28435,N_28346);
or U28808 (N_28808,N_28117,N_28439);
or U28809 (N_28809,N_28295,N_28189);
nand U28810 (N_28810,N_28345,N_28199);
nand U28811 (N_28811,N_28035,N_28276);
or U28812 (N_28812,N_28013,N_28193);
or U28813 (N_28813,N_28035,N_28099);
nor U28814 (N_28814,N_28476,N_28002);
or U28815 (N_28815,N_28473,N_28277);
nor U28816 (N_28816,N_28037,N_28151);
and U28817 (N_28817,N_28474,N_28429);
nand U28818 (N_28818,N_28099,N_28340);
nand U28819 (N_28819,N_28120,N_28102);
or U28820 (N_28820,N_28423,N_28341);
nand U28821 (N_28821,N_28282,N_28383);
or U28822 (N_28822,N_28255,N_28337);
or U28823 (N_28823,N_28035,N_28126);
nand U28824 (N_28824,N_28180,N_28408);
and U28825 (N_28825,N_28196,N_28355);
nor U28826 (N_28826,N_28046,N_28454);
and U28827 (N_28827,N_28141,N_28316);
or U28828 (N_28828,N_28291,N_28160);
nand U28829 (N_28829,N_28111,N_28272);
nor U28830 (N_28830,N_28403,N_28295);
and U28831 (N_28831,N_28170,N_28374);
xnor U28832 (N_28832,N_28072,N_28147);
nand U28833 (N_28833,N_28243,N_28370);
or U28834 (N_28834,N_28305,N_28346);
nor U28835 (N_28835,N_28260,N_28285);
nor U28836 (N_28836,N_28283,N_28084);
nor U28837 (N_28837,N_28406,N_28064);
or U28838 (N_28838,N_28074,N_28399);
nand U28839 (N_28839,N_28277,N_28406);
or U28840 (N_28840,N_28475,N_28435);
nand U28841 (N_28841,N_28351,N_28277);
nand U28842 (N_28842,N_28376,N_28423);
nand U28843 (N_28843,N_28468,N_28082);
nor U28844 (N_28844,N_28096,N_28180);
nand U28845 (N_28845,N_28059,N_28068);
or U28846 (N_28846,N_28447,N_28040);
and U28847 (N_28847,N_28403,N_28275);
nand U28848 (N_28848,N_28301,N_28010);
or U28849 (N_28849,N_28194,N_28499);
or U28850 (N_28850,N_28179,N_28455);
and U28851 (N_28851,N_28198,N_28410);
nand U28852 (N_28852,N_28334,N_28480);
and U28853 (N_28853,N_28344,N_28003);
nand U28854 (N_28854,N_28308,N_28051);
nor U28855 (N_28855,N_28350,N_28264);
nand U28856 (N_28856,N_28126,N_28313);
xor U28857 (N_28857,N_28495,N_28489);
or U28858 (N_28858,N_28202,N_28022);
nor U28859 (N_28859,N_28115,N_28461);
and U28860 (N_28860,N_28425,N_28113);
nor U28861 (N_28861,N_28167,N_28479);
or U28862 (N_28862,N_28121,N_28115);
or U28863 (N_28863,N_28487,N_28307);
and U28864 (N_28864,N_28030,N_28206);
or U28865 (N_28865,N_28412,N_28291);
and U28866 (N_28866,N_28302,N_28444);
nor U28867 (N_28867,N_28141,N_28457);
or U28868 (N_28868,N_28295,N_28306);
nand U28869 (N_28869,N_28435,N_28404);
nand U28870 (N_28870,N_28208,N_28027);
nand U28871 (N_28871,N_28472,N_28194);
nor U28872 (N_28872,N_28046,N_28302);
nand U28873 (N_28873,N_28499,N_28185);
nand U28874 (N_28874,N_28316,N_28340);
and U28875 (N_28875,N_28113,N_28385);
xor U28876 (N_28876,N_28028,N_28160);
nor U28877 (N_28877,N_28022,N_28250);
nor U28878 (N_28878,N_28276,N_28482);
nand U28879 (N_28879,N_28201,N_28210);
or U28880 (N_28880,N_28308,N_28120);
or U28881 (N_28881,N_28466,N_28040);
nand U28882 (N_28882,N_28038,N_28150);
nand U28883 (N_28883,N_28345,N_28317);
xor U28884 (N_28884,N_28222,N_28002);
or U28885 (N_28885,N_28259,N_28263);
or U28886 (N_28886,N_28372,N_28026);
or U28887 (N_28887,N_28172,N_28435);
and U28888 (N_28888,N_28309,N_28359);
or U28889 (N_28889,N_28220,N_28165);
and U28890 (N_28890,N_28414,N_28097);
nand U28891 (N_28891,N_28453,N_28328);
nand U28892 (N_28892,N_28375,N_28264);
and U28893 (N_28893,N_28420,N_28200);
and U28894 (N_28894,N_28237,N_28313);
or U28895 (N_28895,N_28291,N_28408);
or U28896 (N_28896,N_28129,N_28418);
or U28897 (N_28897,N_28493,N_28188);
xor U28898 (N_28898,N_28275,N_28351);
nand U28899 (N_28899,N_28464,N_28222);
and U28900 (N_28900,N_28097,N_28227);
nand U28901 (N_28901,N_28269,N_28017);
nor U28902 (N_28902,N_28083,N_28070);
nand U28903 (N_28903,N_28002,N_28483);
or U28904 (N_28904,N_28381,N_28447);
and U28905 (N_28905,N_28217,N_28448);
nand U28906 (N_28906,N_28278,N_28393);
or U28907 (N_28907,N_28330,N_28340);
and U28908 (N_28908,N_28394,N_28480);
or U28909 (N_28909,N_28355,N_28333);
nor U28910 (N_28910,N_28202,N_28191);
or U28911 (N_28911,N_28487,N_28186);
nor U28912 (N_28912,N_28185,N_28157);
and U28913 (N_28913,N_28001,N_28116);
or U28914 (N_28914,N_28043,N_28427);
and U28915 (N_28915,N_28263,N_28475);
xnor U28916 (N_28916,N_28191,N_28039);
nor U28917 (N_28917,N_28014,N_28107);
and U28918 (N_28918,N_28147,N_28082);
xor U28919 (N_28919,N_28006,N_28473);
or U28920 (N_28920,N_28229,N_28224);
nand U28921 (N_28921,N_28408,N_28277);
nand U28922 (N_28922,N_28177,N_28170);
and U28923 (N_28923,N_28229,N_28282);
or U28924 (N_28924,N_28101,N_28239);
and U28925 (N_28925,N_28266,N_28019);
nand U28926 (N_28926,N_28202,N_28067);
nor U28927 (N_28927,N_28280,N_28349);
nor U28928 (N_28928,N_28358,N_28117);
nor U28929 (N_28929,N_28466,N_28005);
xnor U28930 (N_28930,N_28350,N_28269);
and U28931 (N_28931,N_28447,N_28402);
xor U28932 (N_28932,N_28300,N_28459);
or U28933 (N_28933,N_28173,N_28187);
nor U28934 (N_28934,N_28354,N_28128);
and U28935 (N_28935,N_28244,N_28028);
or U28936 (N_28936,N_28194,N_28358);
and U28937 (N_28937,N_28485,N_28210);
nor U28938 (N_28938,N_28256,N_28364);
xnor U28939 (N_28939,N_28486,N_28048);
and U28940 (N_28940,N_28093,N_28158);
or U28941 (N_28941,N_28158,N_28405);
and U28942 (N_28942,N_28192,N_28343);
nor U28943 (N_28943,N_28261,N_28290);
or U28944 (N_28944,N_28313,N_28229);
xor U28945 (N_28945,N_28306,N_28037);
nand U28946 (N_28946,N_28104,N_28343);
nor U28947 (N_28947,N_28231,N_28260);
nor U28948 (N_28948,N_28001,N_28219);
and U28949 (N_28949,N_28450,N_28104);
or U28950 (N_28950,N_28079,N_28117);
and U28951 (N_28951,N_28482,N_28409);
nand U28952 (N_28952,N_28123,N_28140);
and U28953 (N_28953,N_28078,N_28012);
nand U28954 (N_28954,N_28011,N_28386);
nand U28955 (N_28955,N_28479,N_28130);
nor U28956 (N_28956,N_28227,N_28426);
nor U28957 (N_28957,N_28249,N_28416);
xor U28958 (N_28958,N_28398,N_28324);
nand U28959 (N_28959,N_28032,N_28031);
and U28960 (N_28960,N_28066,N_28112);
nor U28961 (N_28961,N_28012,N_28310);
nand U28962 (N_28962,N_28346,N_28448);
nor U28963 (N_28963,N_28121,N_28303);
nand U28964 (N_28964,N_28023,N_28049);
or U28965 (N_28965,N_28100,N_28370);
or U28966 (N_28966,N_28063,N_28292);
xnor U28967 (N_28967,N_28099,N_28292);
nor U28968 (N_28968,N_28395,N_28241);
and U28969 (N_28969,N_28081,N_28163);
and U28970 (N_28970,N_28034,N_28339);
xor U28971 (N_28971,N_28169,N_28450);
and U28972 (N_28972,N_28018,N_28371);
or U28973 (N_28973,N_28322,N_28343);
nand U28974 (N_28974,N_28293,N_28461);
xnor U28975 (N_28975,N_28296,N_28007);
nor U28976 (N_28976,N_28428,N_28314);
xor U28977 (N_28977,N_28283,N_28131);
xnor U28978 (N_28978,N_28422,N_28020);
nand U28979 (N_28979,N_28117,N_28069);
nand U28980 (N_28980,N_28459,N_28340);
nor U28981 (N_28981,N_28244,N_28267);
xor U28982 (N_28982,N_28090,N_28343);
or U28983 (N_28983,N_28138,N_28075);
xnor U28984 (N_28984,N_28004,N_28190);
nand U28985 (N_28985,N_28075,N_28078);
and U28986 (N_28986,N_28258,N_28432);
and U28987 (N_28987,N_28234,N_28108);
xnor U28988 (N_28988,N_28460,N_28015);
or U28989 (N_28989,N_28370,N_28292);
and U28990 (N_28990,N_28397,N_28113);
or U28991 (N_28991,N_28002,N_28180);
nor U28992 (N_28992,N_28329,N_28184);
or U28993 (N_28993,N_28127,N_28395);
and U28994 (N_28994,N_28093,N_28068);
nor U28995 (N_28995,N_28210,N_28065);
nor U28996 (N_28996,N_28062,N_28098);
nor U28997 (N_28997,N_28397,N_28129);
and U28998 (N_28998,N_28079,N_28085);
nor U28999 (N_28999,N_28314,N_28308);
or U29000 (N_29000,N_28999,N_28714);
xor U29001 (N_29001,N_28882,N_28892);
xor U29002 (N_29002,N_28806,N_28644);
nand U29003 (N_29003,N_28510,N_28589);
nor U29004 (N_29004,N_28720,N_28549);
xnor U29005 (N_29005,N_28989,N_28725);
xnor U29006 (N_29006,N_28960,N_28835);
nor U29007 (N_29007,N_28581,N_28755);
and U29008 (N_29008,N_28854,N_28823);
nor U29009 (N_29009,N_28862,N_28524);
nand U29010 (N_29010,N_28937,N_28632);
xnor U29011 (N_29011,N_28596,N_28583);
nand U29012 (N_29012,N_28958,N_28630);
or U29013 (N_29013,N_28711,N_28848);
nor U29014 (N_29014,N_28907,N_28622);
nor U29015 (N_29015,N_28784,N_28606);
nand U29016 (N_29016,N_28821,N_28810);
and U29017 (N_29017,N_28788,N_28785);
nor U29018 (N_29018,N_28517,N_28790);
nand U29019 (N_29019,N_28814,N_28528);
nor U29020 (N_29020,N_28991,N_28750);
xnor U29021 (N_29021,N_28833,N_28932);
nand U29022 (N_29022,N_28543,N_28856);
or U29023 (N_29023,N_28713,N_28998);
nand U29024 (N_29024,N_28552,N_28874);
nand U29025 (N_29025,N_28863,N_28676);
nor U29026 (N_29026,N_28929,N_28565);
nor U29027 (N_29027,N_28610,N_28769);
or U29028 (N_29028,N_28759,N_28888);
or U29029 (N_29029,N_28727,N_28945);
nand U29030 (N_29030,N_28926,N_28608);
nand U29031 (N_29031,N_28811,N_28896);
nand U29032 (N_29032,N_28600,N_28972);
nand U29033 (N_29033,N_28846,N_28681);
or U29034 (N_29034,N_28566,N_28982);
nor U29035 (N_29035,N_28602,N_28903);
nand U29036 (N_29036,N_28574,N_28919);
and U29037 (N_29037,N_28917,N_28872);
nor U29038 (N_29038,N_28590,N_28700);
xor U29039 (N_29039,N_28656,N_28747);
xor U29040 (N_29040,N_28936,N_28749);
nand U29041 (N_29041,N_28950,N_28618);
nor U29042 (N_29042,N_28651,N_28577);
and U29043 (N_29043,N_28959,N_28890);
xor U29044 (N_29044,N_28557,N_28962);
nand U29045 (N_29045,N_28969,N_28516);
or U29046 (N_29046,N_28551,N_28956);
nor U29047 (N_29047,N_28812,N_28721);
xor U29048 (N_29048,N_28520,N_28740);
xnor U29049 (N_29049,N_28643,N_28922);
and U29050 (N_29050,N_28766,N_28900);
or U29051 (N_29051,N_28935,N_28704);
or U29052 (N_29052,N_28976,N_28573);
nor U29053 (N_29053,N_28792,N_28579);
nand U29054 (N_29054,N_28985,N_28760);
nand U29055 (N_29055,N_28787,N_28842);
xnor U29056 (N_29056,N_28830,N_28580);
nand U29057 (N_29057,N_28658,N_28564);
or U29058 (N_29058,N_28660,N_28518);
or U29059 (N_29059,N_28712,N_28587);
or U29060 (N_29060,N_28649,N_28592);
or U29061 (N_29061,N_28911,N_28883);
and U29062 (N_29062,N_28975,N_28659);
or U29063 (N_29063,N_28930,N_28594);
xor U29064 (N_29064,N_28916,N_28559);
nand U29065 (N_29065,N_28619,N_28815);
nand U29066 (N_29066,N_28561,N_28623);
xor U29067 (N_29067,N_28902,N_28662);
or U29068 (N_29068,N_28536,N_28921);
nor U29069 (N_29069,N_28736,N_28523);
nor U29070 (N_29070,N_28885,N_28940);
nand U29071 (N_29071,N_28988,N_28665);
or U29072 (N_29072,N_28764,N_28604);
or U29073 (N_29073,N_28970,N_28692);
and U29074 (N_29074,N_28794,N_28550);
xnor U29075 (N_29075,N_28677,N_28624);
xnor U29076 (N_29076,N_28555,N_28529);
nand U29077 (N_29077,N_28904,N_28819);
or U29078 (N_29078,N_28642,N_28763);
or U29079 (N_29079,N_28756,N_28718);
and U29080 (N_29080,N_28527,N_28703);
nor U29081 (N_29081,N_28974,N_28847);
nor U29082 (N_29082,N_28813,N_28947);
nor U29083 (N_29083,N_28734,N_28938);
or U29084 (N_29084,N_28715,N_28723);
or U29085 (N_29085,N_28758,N_28831);
or U29086 (N_29086,N_28901,N_28620);
or U29087 (N_29087,N_28946,N_28695);
or U29088 (N_29088,N_28893,N_28939);
nor U29089 (N_29089,N_28684,N_28648);
xor U29090 (N_29090,N_28776,N_28864);
or U29091 (N_29091,N_28669,N_28575);
nor U29092 (N_29092,N_28647,N_28914);
nand U29093 (N_29093,N_28650,N_28729);
nor U29094 (N_29094,N_28514,N_28507);
or U29095 (N_29095,N_28997,N_28558);
and U29096 (N_29096,N_28732,N_28722);
and U29097 (N_29097,N_28957,N_28913);
or U29098 (N_29098,N_28672,N_28840);
nand U29099 (N_29099,N_28568,N_28951);
or U29100 (N_29100,N_28817,N_28591);
or U29101 (N_29101,N_28653,N_28641);
and U29102 (N_29102,N_28702,N_28891);
xor U29103 (N_29103,N_28639,N_28730);
xor U29104 (N_29104,N_28513,N_28675);
nand U29105 (N_29105,N_28538,N_28889);
nand U29106 (N_29106,N_28934,N_28801);
and U29107 (N_29107,N_28906,N_28967);
and U29108 (N_29108,N_28563,N_28636);
nand U29109 (N_29109,N_28719,N_28705);
nand U29110 (N_29110,N_28880,N_28841);
or U29111 (N_29111,N_28767,N_28865);
or U29112 (N_29112,N_28953,N_28878);
and U29113 (N_29113,N_28990,N_28912);
xnor U29114 (N_29114,N_28818,N_28508);
and U29115 (N_29115,N_28678,N_28645);
and U29116 (N_29116,N_28824,N_28915);
nor U29117 (N_29117,N_28526,N_28731);
and U29118 (N_29118,N_28502,N_28857);
xnor U29119 (N_29119,N_28775,N_28586);
or U29120 (N_29120,N_28544,N_28768);
or U29121 (N_29121,N_28687,N_28634);
nor U29122 (N_29122,N_28805,N_28515);
nor U29123 (N_29123,N_28569,N_28927);
or U29124 (N_29124,N_28688,N_28609);
xor U29125 (N_29125,N_28782,N_28797);
or U29126 (N_29126,N_28631,N_28652);
and U29127 (N_29127,N_28978,N_28986);
or U29128 (N_29128,N_28942,N_28837);
nor U29129 (N_29129,N_28850,N_28627);
or U29130 (N_29130,N_28739,N_28598);
nand U29131 (N_29131,N_28534,N_28964);
or U29132 (N_29132,N_28667,N_28873);
and U29133 (N_29133,N_28548,N_28859);
and U29134 (N_29134,N_28709,N_28503);
nor U29135 (N_29135,N_28984,N_28680);
nand U29136 (N_29136,N_28640,N_28708);
or U29137 (N_29137,N_28612,N_28757);
xnor U29138 (N_29138,N_28992,N_28697);
nor U29139 (N_29139,N_28673,N_28663);
and U29140 (N_29140,N_28522,N_28773);
or U29141 (N_29141,N_28851,N_28511);
nor U29142 (N_29142,N_28500,N_28621);
or U29143 (N_29143,N_28617,N_28679);
and U29144 (N_29144,N_28875,N_28855);
and U29145 (N_29145,N_28876,N_28807);
xor U29146 (N_29146,N_28877,N_28949);
nand U29147 (N_29147,N_28699,N_28898);
xnor U29148 (N_29148,N_28966,N_28633);
nand U29149 (N_29149,N_28869,N_28793);
and U29150 (N_29150,N_28710,N_28924);
xnor U29151 (N_29151,N_28770,N_28887);
nor U29152 (N_29152,N_28836,N_28961);
nand U29153 (N_29153,N_28778,N_28707);
nand U29154 (N_29154,N_28560,N_28765);
nand U29155 (N_29155,N_28802,N_28777);
xnor U29156 (N_29156,N_28716,N_28562);
and U29157 (N_29157,N_28535,N_28597);
nor U29158 (N_29158,N_28762,N_28868);
and U29159 (N_29159,N_28706,N_28605);
or U29160 (N_29160,N_28822,N_28931);
nor U29161 (N_29161,N_28585,N_28541);
xor U29162 (N_29162,N_28744,N_28748);
xor U29163 (N_29163,N_28571,N_28803);
or U29164 (N_29164,N_28996,N_28741);
nand U29165 (N_29165,N_28601,N_28682);
nand U29166 (N_29166,N_28944,N_28728);
nand U29167 (N_29167,N_28908,N_28895);
nor U29168 (N_29168,N_28671,N_28858);
nor U29169 (N_29169,N_28745,N_28800);
or U29170 (N_29170,N_28533,N_28780);
or U29171 (N_29171,N_28973,N_28983);
or U29172 (N_29172,N_28826,N_28691);
nand U29173 (N_29173,N_28698,N_28531);
or U29174 (N_29174,N_28894,N_28584);
nand U29175 (N_29175,N_28761,N_28979);
and U29176 (N_29176,N_28920,N_28981);
nand U29177 (N_29177,N_28799,N_28897);
and U29178 (N_29178,N_28816,N_28735);
nor U29179 (N_29179,N_28832,N_28545);
xnor U29180 (N_29180,N_28952,N_28532);
or U29181 (N_29181,N_28603,N_28607);
nor U29182 (N_29182,N_28726,N_28742);
nand U29183 (N_29183,N_28779,N_28582);
or U29184 (N_29184,N_28724,N_28685);
or U29185 (N_29185,N_28521,N_28933);
and U29186 (N_29186,N_28870,N_28925);
nand U29187 (N_29187,N_28839,N_28899);
nor U29188 (N_29188,N_28808,N_28753);
nand U29189 (N_29189,N_28751,N_28843);
nand U29190 (N_29190,N_28501,N_28553);
and U29191 (N_29191,N_28852,N_28664);
and U29192 (N_29192,N_28572,N_28690);
and U29193 (N_29193,N_28537,N_28905);
xnor U29194 (N_29194,N_28578,N_28657);
nor U29195 (N_29195,N_28879,N_28928);
or U29196 (N_29196,N_28737,N_28546);
or U29197 (N_29197,N_28849,N_28834);
xor U29198 (N_29198,N_28625,N_28752);
or U29199 (N_29199,N_28506,N_28955);
and U29200 (N_29200,N_28820,N_28540);
nor U29201 (N_29201,N_28804,N_28881);
and U29202 (N_29202,N_28654,N_28772);
nand U29203 (N_29203,N_28971,N_28683);
and U29204 (N_29204,N_28588,N_28626);
nor U29205 (N_29205,N_28791,N_28827);
or U29206 (N_29206,N_28884,N_28798);
or U29207 (N_29207,N_28615,N_28995);
or U29208 (N_29208,N_28613,N_28993);
nor U29209 (N_29209,N_28666,N_28783);
nand U29210 (N_29210,N_28556,N_28542);
xor U29211 (N_29211,N_28871,N_28923);
nor U29212 (N_29212,N_28733,N_28638);
nor U29213 (N_29213,N_28505,N_28509);
or U29214 (N_29214,N_28668,N_28686);
or U29215 (N_29215,N_28693,N_28629);
nor U29216 (N_29216,N_28599,N_28829);
nor U29217 (N_29217,N_28570,N_28963);
and U29218 (N_29218,N_28954,N_28789);
or U29219 (N_29219,N_28977,N_28786);
or U29220 (N_29220,N_28593,N_28948);
nand U29221 (N_29221,N_28525,N_28635);
xor U29222 (N_29222,N_28628,N_28861);
or U29223 (N_29223,N_28994,N_28909);
nand U29224 (N_29224,N_28828,N_28918);
and U29225 (N_29225,N_28853,N_28867);
and U29226 (N_29226,N_28674,N_28689);
and U29227 (N_29227,N_28701,N_28530);
nand U29228 (N_29228,N_28576,N_28965);
and U29229 (N_29229,N_28694,N_28754);
and U29230 (N_29230,N_28825,N_28504);
and U29231 (N_29231,N_28838,N_28845);
xor U29232 (N_29232,N_28539,N_28844);
xnor U29233 (N_29233,N_28866,N_28795);
nor U29234 (N_29234,N_28743,N_28860);
nand U29235 (N_29235,N_28567,N_28968);
or U29236 (N_29236,N_28595,N_28987);
nor U29237 (N_29237,N_28941,N_28771);
or U29238 (N_29238,N_28512,N_28910);
and U29239 (N_29239,N_28655,N_28781);
or U29240 (N_29240,N_28696,N_28661);
nor U29241 (N_29241,N_28886,N_28616);
nand U29242 (N_29242,N_28980,N_28554);
or U29243 (N_29243,N_28746,N_28738);
or U29244 (N_29244,N_28809,N_28717);
nand U29245 (N_29245,N_28774,N_28611);
or U29246 (N_29246,N_28519,N_28646);
nor U29247 (N_29247,N_28614,N_28670);
nor U29248 (N_29248,N_28943,N_28796);
and U29249 (N_29249,N_28547,N_28637);
nand U29250 (N_29250,N_28708,N_28886);
nor U29251 (N_29251,N_28539,N_28905);
nor U29252 (N_29252,N_28673,N_28714);
nand U29253 (N_29253,N_28739,N_28652);
and U29254 (N_29254,N_28738,N_28654);
nand U29255 (N_29255,N_28667,N_28547);
or U29256 (N_29256,N_28806,N_28600);
or U29257 (N_29257,N_28719,N_28704);
and U29258 (N_29258,N_28892,N_28648);
nand U29259 (N_29259,N_28605,N_28544);
or U29260 (N_29260,N_28553,N_28780);
nand U29261 (N_29261,N_28924,N_28980);
xnor U29262 (N_29262,N_28570,N_28972);
or U29263 (N_29263,N_28892,N_28942);
nor U29264 (N_29264,N_28919,N_28577);
nand U29265 (N_29265,N_28798,N_28760);
nand U29266 (N_29266,N_28831,N_28804);
and U29267 (N_29267,N_28868,N_28700);
nor U29268 (N_29268,N_28626,N_28685);
nand U29269 (N_29269,N_28626,N_28835);
nand U29270 (N_29270,N_28964,N_28969);
nor U29271 (N_29271,N_28862,N_28675);
nand U29272 (N_29272,N_28922,N_28669);
or U29273 (N_29273,N_28591,N_28748);
nor U29274 (N_29274,N_28510,N_28965);
nor U29275 (N_29275,N_28717,N_28564);
nand U29276 (N_29276,N_28589,N_28938);
nand U29277 (N_29277,N_28993,N_28938);
nand U29278 (N_29278,N_28806,N_28864);
xor U29279 (N_29279,N_28659,N_28503);
nor U29280 (N_29280,N_28733,N_28952);
nor U29281 (N_29281,N_28652,N_28677);
nor U29282 (N_29282,N_28837,N_28522);
nor U29283 (N_29283,N_28787,N_28575);
xor U29284 (N_29284,N_28944,N_28649);
nor U29285 (N_29285,N_28526,N_28518);
and U29286 (N_29286,N_28687,N_28822);
nand U29287 (N_29287,N_28841,N_28871);
or U29288 (N_29288,N_28562,N_28932);
nor U29289 (N_29289,N_28985,N_28994);
and U29290 (N_29290,N_28719,N_28715);
and U29291 (N_29291,N_28822,N_28978);
and U29292 (N_29292,N_28898,N_28516);
nor U29293 (N_29293,N_28891,N_28810);
or U29294 (N_29294,N_28581,N_28693);
and U29295 (N_29295,N_28911,N_28858);
and U29296 (N_29296,N_28557,N_28712);
nand U29297 (N_29297,N_28551,N_28572);
or U29298 (N_29298,N_28700,N_28675);
nand U29299 (N_29299,N_28825,N_28827);
nor U29300 (N_29300,N_28872,N_28855);
and U29301 (N_29301,N_28987,N_28643);
nand U29302 (N_29302,N_28771,N_28963);
or U29303 (N_29303,N_28671,N_28506);
or U29304 (N_29304,N_28878,N_28646);
nand U29305 (N_29305,N_28873,N_28931);
nor U29306 (N_29306,N_28745,N_28628);
nand U29307 (N_29307,N_28866,N_28575);
nand U29308 (N_29308,N_28693,N_28889);
and U29309 (N_29309,N_28564,N_28686);
nor U29310 (N_29310,N_28928,N_28534);
xnor U29311 (N_29311,N_28629,N_28776);
nor U29312 (N_29312,N_28709,N_28949);
nand U29313 (N_29313,N_28550,N_28533);
nor U29314 (N_29314,N_28525,N_28862);
nand U29315 (N_29315,N_28823,N_28650);
and U29316 (N_29316,N_28976,N_28612);
nor U29317 (N_29317,N_28547,N_28716);
nand U29318 (N_29318,N_28854,N_28566);
nand U29319 (N_29319,N_28643,N_28647);
xnor U29320 (N_29320,N_28837,N_28847);
and U29321 (N_29321,N_28861,N_28595);
nand U29322 (N_29322,N_28883,N_28530);
nor U29323 (N_29323,N_28962,N_28928);
nor U29324 (N_29324,N_28899,N_28946);
nor U29325 (N_29325,N_28590,N_28647);
and U29326 (N_29326,N_28596,N_28890);
xor U29327 (N_29327,N_28614,N_28972);
and U29328 (N_29328,N_28889,N_28614);
and U29329 (N_29329,N_28849,N_28515);
xnor U29330 (N_29330,N_28890,N_28716);
and U29331 (N_29331,N_28689,N_28870);
or U29332 (N_29332,N_28824,N_28994);
nand U29333 (N_29333,N_28863,N_28563);
or U29334 (N_29334,N_28690,N_28712);
xnor U29335 (N_29335,N_28613,N_28919);
and U29336 (N_29336,N_28883,N_28620);
nor U29337 (N_29337,N_28606,N_28571);
xor U29338 (N_29338,N_28991,N_28837);
nand U29339 (N_29339,N_28911,N_28524);
nand U29340 (N_29340,N_28831,N_28539);
and U29341 (N_29341,N_28838,N_28571);
nor U29342 (N_29342,N_28640,N_28774);
nor U29343 (N_29343,N_28832,N_28635);
nand U29344 (N_29344,N_28708,N_28762);
nand U29345 (N_29345,N_28504,N_28645);
nand U29346 (N_29346,N_28640,N_28641);
nor U29347 (N_29347,N_28714,N_28504);
and U29348 (N_29348,N_28614,N_28763);
or U29349 (N_29349,N_28516,N_28672);
nand U29350 (N_29350,N_28861,N_28616);
nand U29351 (N_29351,N_28777,N_28776);
and U29352 (N_29352,N_28615,N_28608);
nand U29353 (N_29353,N_28845,N_28850);
or U29354 (N_29354,N_28653,N_28736);
nand U29355 (N_29355,N_28652,N_28763);
nor U29356 (N_29356,N_28736,N_28565);
nor U29357 (N_29357,N_28808,N_28629);
or U29358 (N_29358,N_28833,N_28912);
and U29359 (N_29359,N_28674,N_28932);
nor U29360 (N_29360,N_28971,N_28854);
and U29361 (N_29361,N_28604,N_28573);
and U29362 (N_29362,N_28530,N_28775);
nand U29363 (N_29363,N_28976,N_28555);
nand U29364 (N_29364,N_28740,N_28965);
nor U29365 (N_29365,N_28950,N_28770);
xor U29366 (N_29366,N_28877,N_28725);
nor U29367 (N_29367,N_28923,N_28888);
or U29368 (N_29368,N_28573,N_28847);
xor U29369 (N_29369,N_28648,N_28553);
or U29370 (N_29370,N_28863,N_28994);
nor U29371 (N_29371,N_28536,N_28511);
nand U29372 (N_29372,N_28992,N_28691);
and U29373 (N_29373,N_28863,N_28845);
and U29374 (N_29374,N_28532,N_28606);
or U29375 (N_29375,N_28943,N_28964);
nor U29376 (N_29376,N_28716,N_28503);
nand U29377 (N_29377,N_28714,N_28687);
xnor U29378 (N_29378,N_28837,N_28795);
nor U29379 (N_29379,N_28732,N_28762);
nand U29380 (N_29380,N_28589,N_28799);
nor U29381 (N_29381,N_28825,N_28754);
and U29382 (N_29382,N_28896,N_28964);
and U29383 (N_29383,N_28680,N_28997);
xnor U29384 (N_29384,N_28639,N_28668);
or U29385 (N_29385,N_28938,N_28567);
nand U29386 (N_29386,N_28732,N_28636);
nand U29387 (N_29387,N_28839,N_28614);
nor U29388 (N_29388,N_28724,N_28910);
nor U29389 (N_29389,N_28724,N_28982);
or U29390 (N_29390,N_28939,N_28833);
nor U29391 (N_29391,N_28915,N_28911);
or U29392 (N_29392,N_28827,N_28866);
nand U29393 (N_29393,N_28538,N_28810);
and U29394 (N_29394,N_28705,N_28720);
nand U29395 (N_29395,N_28511,N_28925);
or U29396 (N_29396,N_28539,N_28583);
nand U29397 (N_29397,N_28563,N_28853);
nand U29398 (N_29398,N_28682,N_28630);
or U29399 (N_29399,N_28582,N_28617);
xor U29400 (N_29400,N_28720,N_28749);
and U29401 (N_29401,N_28723,N_28542);
or U29402 (N_29402,N_28828,N_28626);
nor U29403 (N_29403,N_28812,N_28601);
nor U29404 (N_29404,N_28677,N_28648);
or U29405 (N_29405,N_28697,N_28732);
or U29406 (N_29406,N_28519,N_28937);
and U29407 (N_29407,N_28646,N_28927);
nor U29408 (N_29408,N_28989,N_28514);
or U29409 (N_29409,N_28621,N_28554);
or U29410 (N_29410,N_28527,N_28777);
or U29411 (N_29411,N_28954,N_28605);
and U29412 (N_29412,N_28528,N_28906);
or U29413 (N_29413,N_28996,N_28539);
nand U29414 (N_29414,N_28951,N_28540);
nand U29415 (N_29415,N_28629,N_28682);
nor U29416 (N_29416,N_28891,N_28613);
nand U29417 (N_29417,N_28877,N_28631);
xor U29418 (N_29418,N_28542,N_28916);
nor U29419 (N_29419,N_28893,N_28948);
nand U29420 (N_29420,N_28733,N_28593);
nand U29421 (N_29421,N_28865,N_28730);
or U29422 (N_29422,N_28870,N_28933);
or U29423 (N_29423,N_28748,N_28679);
nand U29424 (N_29424,N_28574,N_28546);
nor U29425 (N_29425,N_28933,N_28846);
nand U29426 (N_29426,N_28504,N_28976);
nor U29427 (N_29427,N_28992,N_28830);
nor U29428 (N_29428,N_28727,N_28792);
and U29429 (N_29429,N_28978,N_28709);
nand U29430 (N_29430,N_28919,N_28585);
or U29431 (N_29431,N_28510,N_28595);
xor U29432 (N_29432,N_28542,N_28802);
nor U29433 (N_29433,N_28981,N_28578);
xnor U29434 (N_29434,N_28595,N_28691);
and U29435 (N_29435,N_28600,N_28919);
and U29436 (N_29436,N_28781,N_28640);
nand U29437 (N_29437,N_28918,N_28868);
or U29438 (N_29438,N_28640,N_28779);
or U29439 (N_29439,N_28594,N_28581);
nor U29440 (N_29440,N_28751,N_28899);
or U29441 (N_29441,N_28906,N_28700);
and U29442 (N_29442,N_28917,N_28521);
nand U29443 (N_29443,N_28579,N_28811);
and U29444 (N_29444,N_28781,N_28883);
and U29445 (N_29445,N_28917,N_28939);
nand U29446 (N_29446,N_28846,N_28815);
xor U29447 (N_29447,N_28857,N_28911);
nand U29448 (N_29448,N_28621,N_28601);
nand U29449 (N_29449,N_28742,N_28924);
nand U29450 (N_29450,N_28946,N_28906);
nand U29451 (N_29451,N_28924,N_28802);
nor U29452 (N_29452,N_28572,N_28979);
and U29453 (N_29453,N_28918,N_28623);
nand U29454 (N_29454,N_28880,N_28637);
nor U29455 (N_29455,N_28714,N_28536);
and U29456 (N_29456,N_28549,N_28818);
and U29457 (N_29457,N_28976,N_28671);
or U29458 (N_29458,N_28697,N_28544);
nand U29459 (N_29459,N_28829,N_28958);
nor U29460 (N_29460,N_28810,N_28674);
nand U29461 (N_29461,N_28604,N_28862);
nor U29462 (N_29462,N_28518,N_28673);
nor U29463 (N_29463,N_28884,N_28503);
nor U29464 (N_29464,N_28693,N_28679);
and U29465 (N_29465,N_28887,N_28935);
or U29466 (N_29466,N_28612,N_28800);
or U29467 (N_29467,N_28919,N_28752);
or U29468 (N_29468,N_28839,N_28695);
nand U29469 (N_29469,N_28897,N_28719);
and U29470 (N_29470,N_28796,N_28826);
nor U29471 (N_29471,N_28648,N_28683);
or U29472 (N_29472,N_28713,N_28694);
or U29473 (N_29473,N_28710,N_28562);
nand U29474 (N_29474,N_28557,N_28844);
and U29475 (N_29475,N_28748,N_28823);
or U29476 (N_29476,N_28954,N_28973);
and U29477 (N_29477,N_28791,N_28515);
nor U29478 (N_29478,N_28573,N_28609);
and U29479 (N_29479,N_28787,N_28679);
nor U29480 (N_29480,N_28636,N_28683);
nor U29481 (N_29481,N_28537,N_28768);
nand U29482 (N_29482,N_28659,N_28978);
nand U29483 (N_29483,N_28803,N_28838);
nor U29484 (N_29484,N_28591,N_28774);
nor U29485 (N_29485,N_28612,N_28584);
and U29486 (N_29486,N_28785,N_28744);
nand U29487 (N_29487,N_28509,N_28730);
and U29488 (N_29488,N_28708,N_28945);
and U29489 (N_29489,N_28648,N_28996);
and U29490 (N_29490,N_28763,N_28500);
and U29491 (N_29491,N_28669,N_28951);
nand U29492 (N_29492,N_28670,N_28785);
nand U29493 (N_29493,N_28737,N_28593);
nor U29494 (N_29494,N_28521,N_28758);
nand U29495 (N_29495,N_28755,N_28541);
or U29496 (N_29496,N_28628,N_28770);
or U29497 (N_29497,N_28853,N_28715);
nand U29498 (N_29498,N_28659,N_28741);
or U29499 (N_29499,N_28999,N_28735);
and U29500 (N_29500,N_29113,N_29394);
or U29501 (N_29501,N_29473,N_29237);
nor U29502 (N_29502,N_29356,N_29442);
and U29503 (N_29503,N_29483,N_29277);
or U29504 (N_29504,N_29374,N_29360);
or U29505 (N_29505,N_29139,N_29013);
nor U29506 (N_29506,N_29003,N_29372);
nand U29507 (N_29507,N_29050,N_29097);
and U29508 (N_29508,N_29281,N_29399);
and U29509 (N_29509,N_29248,N_29011);
and U29510 (N_29510,N_29099,N_29334);
and U29511 (N_29511,N_29202,N_29088);
xnor U29512 (N_29512,N_29347,N_29370);
xor U29513 (N_29513,N_29185,N_29467);
or U29514 (N_29514,N_29335,N_29104);
nor U29515 (N_29515,N_29386,N_29366);
nor U29516 (N_29516,N_29406,N_29087);
or U29517 (N_29517,N_29269,N_29349);
nor U29518 (N_29518,N_29175,N_29379);
and U29519 (N_29519,N_29101,N_29034);
nand U29520 (N_29520,N_29393,N_29261);
nand U29521 (N_29521,N_29130,N_29491);
and U29522 (N_29522,N_29172,N_29472);
or U29523 (N_29523,N_29299,N_29353);
or U29524 (N_29524,N_29476,N_29159);
nor U29525 (N_29525,N_29188,N_29322);
nand U29526 (N_29526,N_29471,N_29425);
nand U29527 (N_29527,N_29316,N_29153);
and U29528 (N_29528,N_29085,N_29403);
nor U29529 (N_29529,N_29214,N_29218);
and U29530 (N_29530,N_29337,N_29060);
nor U29531 (N_29531,N_29441,N_29273);
nand U29532 (N_29532,N_29246,N_29027);
nand U29533 (N_29533,N_29300,N_29332);
and U29534 (N_29534,N_29245,N_29090);
and U29535 (N_29535,N_29220,N_29047);
or U29536 (N_29536,N_29482,N_29200);
or U29537 (N_29537,N_29124,N_29186);
or U29538 (N_29538,N_29169,N_29145);
nor U29539 (N_29539,N_29233,N_29391);
and U29540 (N_29540,N_29057,N_29475);
and U29541 (N_29541,N_29267,N_29021);
nor U29542 (N_29542,N_29401,N_29466);
and U29543 (N_29543,N_29424,N_29496);
and U29544 (N_29544,N_29304,N_29439);
or U29545 (N_29545,N_29301,N_29479);
nor U29546 (N_29546,N_29089,N_29162);
and U29547 (N_29547,N_29008,N_29210);
nand U29548 (N_29548,N_29385,N_29446);
nor U29549 (N_29549,N_29161,N_29224);
or U29550 (N_29550,N_29096,N_29131);
nand U29551 (N_29551,N_29453,N_29211);
and U29552 (N_29552,N_29118,N_29413);
xnor U29553 (N_29553,N_29309,N_29028);
nor U29554 (N_29554,N_29249,N_29076);
nor U29555 (N_29555,N_29286,N_29375);
and U29556 (N_29556,N_29265,N_29495);
and U29557 (N_29557,N_29389,N_29216);
or U29558 (N_29558,N_29138,N_29344);
or U29559 (N_29559,N_29177,N_29255);
and U29560 (N_29560,N_29461,N_29387);
nor U29561 (N_29561,N_29449,N_29244);
nor U29562 (N_29562,N_29056,N_29423);
xor U29563 (N_29563,N_29095,N_29014);
or U29564 (N_29564,N_29080,N_29031);
or U29565 (N_29565,N_29236,N_29459);
or U29566 (N_29566,N_29054,N_29263);
or U29567 (N_29567,N_29287,N_29359);
xor U29568 (N_29568,N_29317,N_29376);
xnor U29569 (N_29569,N_29230,N_29416);
nor U29570 (N_29570,N_29331,N_29070);
nand U29571 (N_29571,N_29121,N_29445);
or U29572 (N_29572,N_29208,N_29284);
or U29573 (N_29573,N_29452,N_29081);
and U29574 (N_29574,N_29123,N_29402);
nand U29575 (N_29575,N_29274,N_29498);
and U29576 (N_29576,N_29152,N_29320);
nand U29577 (N_29577,N_29390,N_29410);
or U29578 (N_29578,N_29183,N_29132);
nand U29579 (N_29579,N_29158,N_29392);
nor U29580 (N_29580,N_29134,N_29078);
or U29581 (N_29581,N_29381,N_29321);
or U29582 (N_29582,N_29181,N_29045);
and U29583 (N_29583,N_29155,N_29324);
xor U29584 (N_29584,N_29067,N_29336);
xor U29585 (N_29585,N_29010,N_29174);
nand U29586 (N_29586,N_29485,N_29039);
and U29587 (N_29587,N_29166,N_29136);
or U29588 (N_29588,N_29122,N_29357);
nand U29589 (N_29589,N_29457,N_29296);
or U29590 (N_29590,N_29411,N_29384);
nand U29591 (N_29591,N_29084,N_29346);
xor U29592 (N_29592,N_29035,N_29041);
nor U29593 (N_29593,N_29016,N_29448);
and U29594 (N_29594,N_29422,N_29253);
or U29595 (N_29595,N_29001,N_29213);
nand U29596 (N_29596,N_29456,N_29007);
nand U29597 (N_29597,N_29142,N_29022);
and U29598 (N_29598,N_29062,N_29256);
nor U29599 (N_29599,N_29319,N_29182);
or U29600 (N_29600,N_29365,N_29173);
or U29601 (N_29601,N_29023,N_29083);
or U29602 (N_29602,N_29077,N_29156);
xor U29603 (N_29603,N_29484,N_29373);
and U29604 (N_29604,N_29487,N_29184);
or U29605 (N_29605,N_29493,N_29240);
and U29606 (N_29606,N_29030,N_29092);
and U29607 (N_29607,N_29292,N_29378);
xor U29608 (N_29608,N_29140,N_29431);
nor U29609 (N_29609,N_29432,N_29454);
and U29610 (N_29610,N_29180,N_29205);
nor U29611 (N_29611,N_29222,N_29228);
and U29612 (N_29612,N_29380,N_29111);
nor U29613 (N_29613,N_29225,N_29051);
nand U29614 (N_29614,N_29190,N_29151);
and U29615 (N_29615,N_29458,N_29364);
nor U29616 (N_29616,N_29264,N_29234);
xnor U29617 (N_29617,N_29009,N_29368);
or U29618 (N_29618,N_29407,N_29477);
or U29619 (N_29619,N_29193,N_29000);
and U29620 (N_29620,N_29105,N_29404);
nor U29621 (N_29621,N_29318,N_29271);
and U29622 (N_29622,N_29146,N_29178);
nand U29623 (N_29623,N_29437,N_29191);
nand U29624 (N_29624,N_29443,N_29143);
nor U29625 (N_29625,N_29154,N_29341);
nand U29626 (N_29626,N_29073,N_29192);
xor U29627 (N_29627,N_29053,N_29419);
nor U29628 (N_29628,N_29086,N_29427);
xor U29629 (N_29629,N_29114,N_29283);
nand U29630 (N_29630,N_29306,N_29017);
nor U29631 (N_29631,N_29302,N_29494);
or U29632 (N_29632,N_29232,N_29323);
or U29633 (N_29633,N_29415,N_29266);
nand U29634 (N_29634,N_29223,N_29204);
and U29635 (N_29635,N_29098,N_29470);
nor U29636 (N_29636,N_29260,N_29075);
and U29637 (N_29637,N_29215,N_29106);
or U29638 (N_29638,N_29037,N_29135);
nand U29639 (N_29639,N_29032,N_29438);
and U29640 (N_29640,N_29094,N_29072);
and U29641 (N_29641,N_29462,N_29069);
nor U29642 (N_29642,N_29270,N_29128);
nand U29643 (N_29643,N_29018,N_29147);
or U29644 (N_29644,N_29235,N_29110);
or U29645 (N_29645,N_29327,N_29238);
and U29646 (N_29646,N_29354,N_29486);
nor U29647 (N_29647,N_29333,N_29282);
and U29648 (N_29648,N_29217,N_29229);
nor U29649 (N_29649,N_29285,N_29463);
nor U29650 (N_29650,N_29071,N_29382);
and U29651 (N_29651,N_29395,N_29250);
and U29652 (N_29652,N_29068,N_29164);
nor U29653 (N_29653,N_29465,N_29171);
nand U29654 (N_29654,N_29257,N_29421);
or U29655 (N_29655,N_29297,N_29046);
nand U29656 (N_29656,N_29428,N_29004);
nor U29657 (N_29657,N_29025,N_29189);
and U29658 (N_29658,N_29420,N_29444);
nand U29659 (N_29659,N_29355,N_29430);
xor U29660 (N_29660,N_29129,N_29052);
or U29661 (N_29661,N_29489,N_29065);
and U29662 (N_29662,N_29126,N_29199);
nor U29663 (N_29663,N_29313,N_29388);
nor U29664 (N_29664,N_29195,N_29371);
nand U29665 (N_29665,N_29338,N_29490);
nand U29666 (N_29666,N_29207,N_29455);
nor U29667 (N_29667,N_29329,N_29109);
or U29668 (N_29668,N_29339,N_29362);
nor U29669 (N_29669,N_29196,N_29012);
nor U29670 (N_29670,N_29157,N_29417);
nand U29671 (N_29671,N_29328,N_29451);
and U29672 (N_29672,N_29043,N_29042);
and U29673 (N_29673,N_29170,N_29061);
or U29674 (N_29674,N_29272,N_29377);
nor U29675 (N_29675,N_29117,N_29279);
nor U29676 (N_29676,N_29242,N_29221);
nand U29677 (N_29677,N_29127,N_29289);
or U29678 (N_29678,N_29450,N_29160);
nor U29679 (N_29679,N_29044,N_29194);
nor U29680 (N_29680,N_29468,N_29150);
xor U29681 (N_29681,N_29049,N_29414);
nand U29682 (N_29682,N_29033,N_29116);
nand U29683 (N_29683,N_29029,N_29315);
xor U29684 (N_29684,N_29298,N_29325);
xnor U29685 (N_29685,N_29103,N_29440);
and U29686 (N_29686,N_29115,N_29201);
or U29687 (N_29687,N_29040,N_29093);
nand U29688 (N_29688,N_29262,N_29102);
nor U29689 (N_29689,N_29167,N_29227);
nor U29690 (N_29690,N_29293,N_29342);
and U29691 (N_29691,N_29412,N_29383);
nand U29692 (N_29692,N_29064,N_29002);
nor U29693 (N_29693,N_29006,N_29429);
and U29694 (N_29694,N_29165,N_29247);
and U29695 (N_29695,N_29308,N_29361);
nand U29696 (N_29696,N_29268,N_29091);
nor U29697 (N_29697,N_29259,N_29082);
and U29698 (N_29698,N_29005,N_29241);
and U29699 (N_29699,N_29363,N_29251);
nor U29700 (N_29700,N_29469,N_29447);
and U29701 (N_29701,N_29149,N_29100);
nor U29702 (N_29702,N_29163,N_29499);
xor U29703 (N_29703,N_29055,N_29187);
nand U29704 (N_29704,N_29397,N_29464);
or U29705 (N_29705,N_29294,N_29203);
xnor U29706 (N_29706,N_29400,N_29079);
nand U29707 (N_29707,N_29433,N_29426);
or U29708 (N_29708,N_29340,N_29275);
nor U29709 (N_29709,N_29295,N_29254);
nand U29710 (N_29710,N_29176,N_29144);
xor U29711 (N_29711,N_29303,N_29480);
nand U29712 (N_29712,N_29133,N_29398);
nor U29713 (N_29713,N_29481,N_29020);
nor U29714 (N_29714,N_29280,N_29409);
xnor U29715 (N_29715,N_29258,N_29492);
and U29716 (N_29716,N_29408,N_29345);
and U29717 (N_29717,N_29436,N_29058);
or U29718 (N_29718,N_29141,N_29059);
nor U29719 (N_29719,N_29418,N_29307);
nand U29720 (N_29720,N_29243,N_29405);
and U29721 (N_29721,N_29311,N_29305);
or U29722 (N_29722,N_29206,N_29343);
nor U29723 (N_29723,N_29478,N_29066);
or U29724 (N_29724,N_29063,N_29367);
nand U29725 (N_29725,N_29026,N_29107);
or U29726 (N_29726,N_29231,N_29209);
nand U29727 (N_29727,N_29120,N_29435);
and U29728 (N_29728,N_29239,N_29314);
or U29729 (N_29729,N_29310,N_29197);
or U29730 (N_29730,N_29119,N_29278);
nor U29731 (N_29731,N_29148,N_29024);
or U29732 (N_29732,N_29460,N_29351);
xor U29733 (N_29733,N_29048,N_29252);
or U29734 (N_29734,N_29036,N_29015);
nand U29735 (N_29735,N_29352,N_29369);
xor U29736 (N_29736,N_29291,N_29074);
nor U29737 (N_29737,N_29137,N_29108);
or U29738 (N_29738,N_29348,N_29434);
nand U29739 (N_29739,N_29198,N_29330);
and U29740 (N_29740,N_29112,N_29019);
and U29741 (N_29741,N_29219,N_29276);
and U29742 (N_29742,N_29350,N_29290);
nand U29743 (N_29743,N_29326,N_29179);
and U29744 (N_29744,N_29168,N_29312);
and U29745 (N_29745,N_29288,N_29226);
nand U29746 (N_29746,N_29212,N_29038);
nand U29747 (N_29747,N_29358,N_29474);
and U29748 (N_29748,N_29125,N_29497);
and U29749 (N_29749,N_29488,N_29396);
and U29750 (N_29750,N_29084,N_29071);
or U29751 (N_29751,N_29051,N_29490);
and U29752 (N_29752,N_29411,N_29421);
or U29753 (N_29753,N_29464,N_29197);
nor U29754 (N_29754,N_29250,N_29196);
nand U29755 (N_29755,N_29422,N_29218);
and U29756 (N_29756,N_29092,N_29124);
nor U29757 (N_29757,N_29104,N_29046);
nand U29758 (N_29758,N_29435,N_29215);
xnor U29759 (N_29759,N_29011,N_29443);
nand U29760 (N_29760,N_29316,N_29205);
and U29761 (N_29761,N_29100,N_29269);
nor U29762 (N_29762,N_29393,N_29309);
and U29763 (N_29763,N_29293,N_29339);
xor U29764 (N_29764,N_29316,N_29391);
xnor U29765 (N_29765,N_29360,N_29134);
xnor U29766 (N_29766,N_29157,N_29495);
and U29767 (N_29767,N_29381,N_29318);
or U29768 (N_29768,N_29123,N_29192);
and U29769 (N_29769,N_29463,N_29250);
nand U29770 (N_29770,N_29488,N_29225);
and U29771 (N_29771,N_29055,N_29001);
or U29772 (N_29772,N_29440,N_29172);
xnor U29773 (N_29773,N_29367,N_29385);
nor U29774 (N_29774,N_29030,N_29000);
or U29775 (N_29775,N_29323,N_29302);
nand U29776 (N_29776,N_29315,N_29156);
nand U29777 (N_29777,N_29466,N_29454);
and U29778 (N_29778,N_29491,N_29074);
nor U29779 (N_29779,N_29391,N_29343);
nor U29780 (N_29780,N_29358,N_29146);
or U29781 (N_29781,N_29347,N_29456);
xor U29782 (N_29782,N_29367,N_29378);
or U29783 (N_29783,N_29221,N_29008);
or U29784 (N_29784,N_29372,N_29048);
or U29785 (N_29785,N_29404,N_29209);
nand U29786 (N_29786,N_29004,N_29076);
nand U29787 (N_29787,N_29193,N_29154);
or U29788 (N_29788,N_29456,N_29031);
nor U29789 (N_29789,N_29472,N_29043);
and U29790 (N_29790,N_29442,N_29296);
and U29791 (N_29791,N_29219,N_29372);
and U29792 (N_29792,N_29292,N_29156);
or U29793 (N_29793,N_29411,N_29007);
and U29794 (N_29794,N_29007,N_29356);
or U29795 (N_29795,N_29146,N_29360);
nand U29796 (N_29796,N_29431,N_29213);
xnor U29797 (N_29797,N_29149,N_29347);
nor U29798 (N_29798,N_29353,N_29075);
nor U29799 (N_29799,N_29367,N_29431);
and U29800 (N_29800,N_29212,N_29368);
and U29801 (N_29801,N_29304,N_29153);
or U29802 (N_29802,N_29318,N_29086);
nand U29803 (N_29803,N_29224,N_29228);
nor U29804 (N_29804,N_29178,N_29158);
or U29805 (N_29805,N_29400,N_29217);
nand U29806 (N_29806,N_29462,N_29232);
xor U29807 (N_29807,N_29294,N_29355);
and U29808 (N_29808,N_29449,N_29103);
and U29809 (N_29809,N_29479,N_29494);
and U29810 (N_29810,N_29082,N_29203);
xnor U29811 (N_29811,N_29337,N_29262);
nor U29812 (N_29812,N_29139,N_29300);
and U29813 (N_29813,N_29334,N_29137);
xor U29814 (N_29814,N_29490,N_29488);
xor U29815 (N_29815,N_29065,N_29050);
nor U29816 (N_29816,N_29411,N_29398);
or U29817 (N_29817,N_29323,N_29471);
or U29818 (N_29818,N_29457,N_29492);
nor U29819 (N_29819,N_29380,N_29010);
and U29820 (N_29820,N_29115,N_29265);
nor U29821 (N_29821,N_29003,N_29156);
nand U29822 (N_29822,N_29365,N_29148);
nor U29823 (N_29823,N_29207,N_29401);
and U29824 (N_29824,N_29324,N_29140);
and U29825 (N_29825,N_29089,N_29285);
nor U29826 (N_29826,N_29214,N_29058);
or U29827 (N_29827,N_29111,N_29214);
or U29828 (N_29828,N_29266,N_29107);
and U29829 (N_29829,N_29116,N_29071);
or U29830 (N_29830,N_29452,N_29045);
nor U29831 (N_29831,N_29463,N_29064);
or U29832 (N_29832,N_29186,N_29126);
nand U29833 (N_29833,N_29143,N_29498);
nand U29834 (N_29834,N_29398,N_29140);
and U29835 (N_29835,N_29378,N_29457);
xnor U29836 (N_29836,N_29432,N_29246);
or U29837 (N_29837,N_29449,N_29374);
nor U29838 (N_29838,N_29058,N_29243);
nor U29839 (N_29839,N_29319,N_29381);
nand U29840 (N_29840,N_29227,N_29346);
xor U29841 (N_29841,N_29457,N_29337);
nor U29842 (N_29842,N_29315,N_29041);
or U29843 (N_29843,N_29211,N_29423);
nor U29844 (N_29844,N_29108,N_29140);
nand U29845 (N_29845,N_29385,N_29342);
nand U29846 (N_29846,N_29143,N_29063);
and U29847 (N_29847,N_29292,N_29071);
or U29848 (N_29848,N_29162,N_29381);
or U29849 (N_29849,N_29374,N_29336);
or U29850 (N_29850,N_29186,N_29315);
nand U29851 (N_29851,N_29309,N_29218);
and U29852 (N_29852,N_29398,N_29173);
and U29853 (N_29853,N_29467,N_29054);
nand U29854 (N_29854,N_29254,N_29341);
and U29855 (N_29855,N_29460,N_29348);
or U29856 (N_29856,N_29265,N_29106);
nor U29857 (N_29857,N_29250,N_29319);
and U29858 (N_29858,N_29139,N_29290);
nor U29859 (N_29859,N_29185,N_29308);
and U29860 (N_29860,N_29445,N_29468);
nor U29861 (N_29861,N_29030,N_29038);
or U29862 (N_29862,N_29262,N_29276);
and U29863 (N_29863,N_29050,N_29257);
and U29864 (N_29864,N_29426,N_29384);
nor U29865 (N_29865,N_29351,N_29380);
or U29866 (N_29866,N_29253,N_29291);
nor U29867 (N_29867,N_29085,N_29477);
xor U29868 (N_29868,N_29219,N_29486);
or U29869 (N_29869,N_29476,N_29362);
or U29870 (N_29870,N_29261,N_29113);
nor U29871 (N_29871,N_29040,N_29387);
nor U29872 (N_29872,N_29058,N_29340);
and U29873 (N_29873,N_29164,N_29163);
nor U29874 (N_29874,N_29204,N_29363);
nor U29875 (N_29875,N_29479,N_29019);
nand U29876 (N_29876,N_29468,N_29095);
and U29877 (N_29877,N_29138,N_29043);
or U29878 (N_29878,N_29433,N_29373);
or U29879 (N_29879,N_29149,N_29152);
xnor U29880 (N_29880,N_29127,N_29457);
nor U29881 (N_29881,N_29295,N_29200);
nand U29882 (N_29882,N_29231,N_29063);
and U29883 (N_29883,N_29000,N_29012);
or U29884 (N_29884,N_29211,N_29168);
nand U29885 (N_29885,N_29160,N_29050);
nor U29886 (N_29886,N_29300,N_29391);
and U29887 (N_29887,N_29303,N_29486);
nand U29888 (N_29888,N_29469,N_29078);
nand U29889 (N_29889,N_29130,N_29396);
and U29890 (N_29890,N_29040,N_29376);
nor U29891 (N_29891,N_29383,N_29318);
or U29892 (N_29892,N_29330,N_29482);
nand U29893 (N_29893,N_29432,N_29375);
and U29894 (N_29894,N_29110,N_29035);
nor U29895 (N_29895,N_29346,N_29427);
or U29896 (N_29896,N_29367,N_29434);
nor U29897 (N_29897,N_29323,N_29074);
nand U29898 (N_29898,N_29131,N_29275);
nor U29899 (N_29899,N_29381,N_29327);
nor U29900 (N_29900,N_29496,N_29358);
nand U29901 (N_29901,N_29215,N_29087);
and U29902 (N_29902,N_29396,N_29226);
xnor U29903 (N_29903,N_29233,N_29294);
or U29904 (N_29904,N_29251,N_29451);
or U29905 (N_29905,N_29162,N_29269);
xor U29906 (N_29906,N_29116,N_29146);
nand U29907 (N_29907,N_29300,N_29268);
nor U29908 (N_29908,N_29148,N_29413);
xnor U29909 (N_29909,N_29152,N_29426);
and U29910 (N_29910,N_29428,N_29301);
nor U29911 (N_29911,N_29313,N_29081);
nand U29912 (N_29912,N_29446,N_29345);
or U29913 (N_29913,N_29201,N_29456);
and U29914 (N_29914,N_29274,N_29426);
and U29915 (N_29915,N_29214,N_29341);
and U29916 (N_29916,N_29169,N_29062);
nor U29917 (N_29917,N_29481,N_29298);
nand U29918 (N_29918,N_29357,N_29329);
or U29919 (N_29919,N_29150,N_29045);
nand U29920 (N_29920,N_29477,N_29281);
nand U29921 (N_29921,N_29035,N_29071);
and U29922 (N_29922,N_29043,N_29372);
nor U29923 (N_29923,N_29009,N_29010);
or U29924 (N_29924,N_29251,N_29163);
nor U29925 (N_29925,N_29304,N_29121);
nand U29926 (N_29926,N_29227,N_29041);
and U29927 (N_29927,N_29383,N_29071);
or U29928 (N_29928,N_29351,N_29363);
nor U29929 (N_29929,N_29214,N_29416);
and U29930 (N_29930,N_29001,N_29306);
nand U29931 (N_29931,N_29499,N_29009);
and U29932 (N_29932,N_29069,N_29441);
or U29933 (N_29933,N_29178,N_29347);
nand U29934 (N_29934,N_29218,N_29467);
and U29935 (N_29935,N_29156,N_29045);
or U29936 (N_29936,N_29216,N_29296);
and U29937 (N_29937,N_29135,N_29067);
or U29938 (N_29938,N_29263,N_29477);
and U29939 (N_29939,N_29340,N_29067);
and U29940 (N_29940,N_29313,N_29378);
or U29941 (N_29941,N_29303,N_29344);
nand U29942 (N_29942,N_29308,N_29139);
nand U29943 (N_29943,N_29087,N_29139);
xor U29944 (N_29944,N_29138,N_29135);
nand U29945 (N_29945,N_29030,N_29371);
xor U29946 (N_29946,N_29442,N_29345);
nor U29947 (N_29947,N_29220,N_29368);
or U29948 (N_29948,N_29264,N_29307);
nor U29949 (N_29949,N_29118,N_29345);
and U29950 (N_29950,N_29225,N_29011);
and U29951 (N_29951,N_29322,N_29242);
nor U29952 (N_29952,N_29383,N_29001);
nor U29953 (N_29953,N_29341,N_29100);
and U29954 (N_29954,N_29253,N_29045);
or U29955 (N_29955,N_29291,N_29002);
and U29956 (N_29956,N_29304,N_29254);
xor U29957 (N_29957,N_29277,N_29269);
and U29958 (N_29958,N_29479,N_29249);
and U29959 (N_29959,N_29200,N_29474);
and U29960 (N_29960,N_29140,N_29049);
xnor U29961 (N_29961,N_29377,N_29286);
or U29962 (N_29962,N_29025,N_29362);
nor U29963 (N_29963,N_29127,N_29168);
nor U29964 (N_29964,N_29213,N_29203);
xor U29965 (N_29965,N_29114,N_29284);
xnor U29966 (N_29966,N_29330,N_29176);
nand U29967 (N_29967,N_29467,N_29423);
nor U29968 (N_29968,N_29056,N_29322);
nor U29969 (N_29969,N_29221,N_29421);
xor U29970 (N_29970,N_29061,N_29312);
nor U29971 (N_29971,N_29210,N_29425);
xor U29972 (N_29972,N_29282,N_29095);
nor U29973 (N_29973,N_29473,N_29047);
or U29974 (N_29974,N_29407,N_29231);
nor U29975 (N_29975,N_29290,N_29225);
and U29976 (N_29976,N_29425,N_29211);
xnor U29977 (N_29977,N_29033,N_29090);
and U29978 (N_29978,N_29315,N_29030);
and U29979 (N_29979,N_29162,N_29253);
or U29980 (N_29980,N_29218,N_29406);
nor U29981 (N_29981,N_29055,N_29143);
and U29982 (N_29982,N_29158,N_29465);
and U29983 (N_29983,N_29203,N_29128);
nand U29984 (N_29984,N_29236,N_29124);
and U29985 (N_29985,N_29165,N_29127);
and U29986 (N_29986,N_29216,N_29452);
nand U29987 (N_29987,N_29033,N_29161);
xnor U29988 (N_29988,N_29284,N_29191);
nand U29989 (N_29989,N_29318,N_29300);
nand U29990 (N_29990,N_29391,N_29412);
and U29991 (N_29991,N_29098,N_29127);
and U29992 (N_29992,N_29239,N_29065);
nor U29993 (N_29993,N_29255,N_29119);
nand U29994 (N_29994,N_29454,N_29096);
or U29995 (N_29995,N_29355,N_29081);
or U29996 (N_29996,N_29213,N_29360);
xor U29997 (N_29997,N_29160,N_29118);
nor U29998 (N_29998,N_29303,N_29301);
nor U29999 (N_29999,N_29049,N_29153);
nor U30000 (N_30000,N_29793,N_29615);
or U30001 (N_30001,N_29604,N_29570);
and U30002 (N_30002,N_29571,N_29751);
xnor U30003 (N_30003,N_29979,N_29501);
or U30004 (N_30004,N_29671,N_29623);
nand U30005 (N_30005,N_29773,N_29957);
nand U30006 (N_30006,N_29714,N_29962);
nand U30007 (N_30007,N_29936,N_29802);
nor U30008 (N_30008,N_29889,N_29865);
or U30009 (N_30009,N_29996,N_29645);
nor U30010 (N_30010,N_29814,N_29992);
xor U30011 (N_30011,N_29965,N_29854);
or U30012 (N_30012,N_29937,N_29838);
nor U30013 (N_30013,N_29929,N_29703);
nor U30014 (N_30014,N_29797,N_29526);
or U30015 (N_30015,N_29672,N_29517);
or U30016 (N_30016,N_29502,N_29626);
xnor U30017 (N_30017,N_29805,N_29588);
or U30018 (N_30018,N_29920,N_29956);
nand U30019 (N_30019,N_29777,N_29737);
xnor U30020 (N_30020,N_29946,N_29606);
and U30021 (N_30021,N_29682,N_29534);
nor U30022 (N_30022,N_29758,N_29701);
xor U30023 (N_30023,N_29594,N_29704);
and U30024 (N_30024,N_29766,N_29527);
nor U30025 (N_30025,N_29646,N_29537);
or U30026 (N_30026,N_29665,N_29923);
and U30027 (N_30027,N_29644,N_29762);
and U30028 (N_30028,N_29840,N_29613);
nand U30029 (N_30029,N_29640,N_29643);
or U30030 (N_30030,N_29636,N_29991);
and U30031 (N_30031,N_29964,N_29503);
xnor U30032 (N_30032,N_29883,N_29817);
and U30033 (N_30033,N_29719,N_29598);
or U30034 (N_30034,N_29545,N_29507);
and U30035 (N_30035,N_29811,N_29715);
nand U30036 (N_30036,N_29879,N_29585);
or U30037 (N_30037,N_29949,N_29930);
nor U30038 (N_30038,N_29548,N_29736);
and U30039 (N_30039,N_29721,N_29668);
or U30040 (N_30040,N_29911,N_29738);
or U30041 (N_30041,N_29987,N_29584);
and U30042 (N_30042,N_29832,N_29898);
nand U30043 (N_30043,N_29972,N_29899);
nand U30044 (N_30044,N_29712,N_29576);
and U30045 (N_30045,N_29560,N_29620);
xnor U30046 (N_30046,N_29885,N_29639);
nor U30047 (N_30047,N_29687,N_29755);
nand U30048 (N_30048,N_29870,N_29711);
or U30049 (N_30049,N_29670,N_29819);
or U30050 (N_30050,N_29628,N_29593);
nand U30051 (N_30051,N_29667,N_29908);
or U30052 (N_30052,N_29546,N_29746);
nor U30053 (N_30053,N_29788,N_29562);
nand U30054 (N_30054,N_29863,N_29520);
and U30055 (N_30055,N_29980,N_29945);
nand U30056 (N_30056,N_29845,N_29589);
or U30057 (N_30057,N_29891,N_29839);
or U30058 (N_30058,N_29754,N_29932);
nand U30059 (N_30059,N_29795,N_29647);
and U30060 (N_30060,N_29504,N_29824);
or U30061 (N_30061,N_29694,N_29761);
nor U30062 (N_30062,N_29709,N_29774);
nand U30063 (N_30063,N_29919,N_29505);
and U30064 (N_30064,N_29515,N_29592);
nand U30065 (N_30065,N_29798,N_29903);
and U30066 (N_30066,N_29988,N_29688);
and U30067 (N_30067,N_29747,N_29901);
nor U30068 (N_30068,N_29720,N_29599);
or U30069 (N_30069,N_29816,N_29535);
and U30070 (N_30070,N_29629,N_29782);
or U30071 (N_30071,N_29904,N_29935);
and U30072 (N_30072,N_29781,N_29931);
or U30073 (N_30073,N_29986,N_29506);
or U30074 (N_30074,N_29952,N_29834);
and U30075 (N_30075,N_29861,N_29740);
or U30076 (N_30076,N_29950,N_29918);
and U30077 (N_30077,N_29691,N_29806);
or U30078 (N_30078,N_29605,N_29561);
nand U30079 (N_30079,N_29897,N_29828);
nand U30080 (N_30080,N_29698,N_29942);
nand U30081 (N_30081,N_29511,N_29739);
nand U30082 (N_30082,N_29808,N_29539);
or U30083 (N_30083,N_29666,N_29540);
and U30084 (N_30084,N_29678,N_29752);
or U30085 (N_30085,N_29522,N_29621);
nand U30086 (N_30086,N_29985,N_29702);
nor U30087 (N_30087,N_29884,N_29696);
nand U30088 (N_30088,N_29882,N_29780);
and U30089 (N_30089,N_29513,N_29710);
and U30090 (N_30090,N_29743,N_29982);
nand U30091 (N_30091,N_29547,N_29812);
or U30092 (N_30092,N_29800,N_29954);
nor U30093 (N_30093,N_29959,N_29757);
nand U30094 (N_30094,N_29809,N_29858);
and U30095 (N_30095,N_29581,N_29971);
or U30096 (N_30096,N_29917,N_29566);
nor U30097 (N_30097,N_29693,N_29940);
nand U30098 (N_30098,N_29902,N_29748);
nor U30099 (N_30099,N_29896,N_29794);
nand U30100 (N_30100,N_29852,N_29669);
xnor U30101 (N_30101,N_29567,N_29681);
and U30102 (N_30102,N_29587,N_29841);
nand U30103 (N_30103,N_29772,N_29705);
and U30104 (N_30104,N_29549,N_29765);
nand U30105 (N_30105,N_29998,N_29555);
or U30106 (N_30106,N_29791,N_29827);
nand U30107 (N_30107,N_29608,N_29776);
nand U30108 (N_30108,N_29699,N_29722);
and U30109 (N_30109,N_29862,N_29610);
and U30110 (N_30110,N_29536,N_29831);
nand U30111 (N_30111,N_29759,N_29966);
nor U30112 (N_30112,N_29893,N_29915);
xor U30113 (N_30113,N_29600,N_29627);
nand U30114 (N_30114,N_29944,N_29663);
xnor U30115 (N_30115,N_29963,N_29654);
or U30116 (N_30116,N_29813,N_29994);
nor U30117 (N_30117,N_29895,N_29662);
or U30118 (N_30118,N_29708,N_29951);
or U30119 (N_30119,N_29619,N_29529);
and U30120 (N_30120,N_29857,N_29771);
and U30121 (N_30121,N_29881,N_29750);
and U30122 (N_30122,N_29922,N_29789);
and U30123 (N_30123,N_29677,N_29652);
and U30124 (N_30124,N_29509,N_29717);
and U30125 (N_30125,N_29855,N_29579);
nor U30126 (N_30126,N_29916,N_29564);
and U30127 (N_30127,N_29925,N_29744);
or U30128 (N_30128,N_29790,N_29799);
or U30129 (N_30129,N_29989,N_29968);
xor U30130 (N_30130,N_29878,N_29869);
or U30131 (N_30131,N_29638,N_29616);
nand U30132 (N_30132,N_29836,N_29853);
nor U30133 (N_30133,N_29970,N_29846);
or U30134 (N_30134,N_29573,N_29538);
nand U30135 (N_30135,N_29770,N_29591);
nand U30136 (N_30136,N_29907,N_29675);
nand U30137 (N_30137,N_29533,N_29912);
or U30138 (N_30138,N_29601,N_29820);
nor U30139 (N_30139,N_29871,N_29732);
nand U30140 (N_30140,N_29928,N_29848);
or U30141 (N_30141,N_29731,N_29974);
and U30142 (N_30142,N_29574,N_29769);
nor U30143 (N_30143,N_29822,N_29778);
nor U30144 (N_30144,N_29847,N_29657);
nand U30145 (N_30145,N_29713,N_29837);
and U30146 (N_30146,N_29978,N_29597);
nand U30147 (N_30147,N_29528,N_29921);
nand U30148 (N_30148,N_29784,N_29868);
nor U30149 (N_30149,N_29558,N_29559);
nor U30150 (N_30150,N_29697,N_29826);
nor U30151 (N_30151,N_29723,N_29787);
xnor U30152 (N_30152,N_29660,N_29933);
xor U30153 (N_30153,N_29661,N_29823);
and U30154 (N_30154,N_29725,N_29872);
and U30155 (N_30155,N_29727,N_29867);
and U30156 (N_30156,N_29909,N_29641);
nor U30157 (N_30157,N_29984,N_29842);
and U30158 (N_30158,N_29553,N_29999);
nor U30159 (N_30159,N_29947,N_29653);
nand U30160 (N_30160,N_29541,N_29960);
nor U30161 (N_30161,N_29900,N_29637);
and U30162 (N_30162,N_29631,N_29851);
nand U30163 (N_30163,N_29939,N_29718);
nor U30164 (N_30164,N_29583,N_29582);
or U30165 (N_30165,N_29676,N_29821);
or U30166 (N_30166,N_29531,N_29633);
and U30167 (N_30167,N_29810,N_29807);
and U30168 (N_30168,N_29658,N_29686);
nor U30169 (N_30169,N_29888,N_29734);
or U30170 (N_30170,N_29792,N_29651);
or U30171 (N_30171,N_29568,N_29938);
xnor U30172 (N_30172,N_29887,N_29892);
nor U30173 (N_30173,N_29679,N_29655);
or U30174 (N_30174,N_29707,N_29550);
or U30175 (N_30175,N_29625,N_29642);
or U30176 (N_30176,N_29634,N_29864);
xnor U30177 (N_30177,N_29523,N_29607);
or U30178 (N_30178,N_29519,N_29815);
nand U30179 (N_30179,N_29521,N_29981);
nand U30180 (N_30180,N_29779,N_29542);
or U30181 (N_30181,N_29603,N_29659);
nand U30182 (N_30182,N_29516,N_29804);
nor U30183 (N_30183,N_29913,N_29756);
nor U30184 (N_30184,N_29941,N_29783);
and U30185 (N_30185,N_29849,N_29544);
nor U30186 (N_30186,N_29674,N_29976);
xnor U30187 (N_30187,N_29575,N_29524);
nor U30188 (N_30188,N_29635,N_29927);
nor U30189 (N_30189,N_29983,N_29914);
nor U30190 (N_30190,N_29695,N_29510);
and U30191 (N_30191,N_29866,N_29844);
or U30192 (N_30192,N_29609,N_29801);
and U30193 (N_30193,N_29572,N_29632);
or U30194 (N_30194,N_29993,N_29512);
and U30195 (N_30195,N_29997,N_29680);
nor U30196 (N_30196,N_29690,N_29689);
and U30197 (N_30197,N_29733,N_29786);
nor U30198 (N_30198,N_29578,N_29934);
nor U30199 (N_30199,N_29990,N_29875);
nor U30200 (N_30200,N_29890,N_29877);
nor U30201 (N_30201,N_29730,N_29684);
or U30202 (N_30202,N_29775,N_29551);
and U30203 (N_30203,N_29835,N_29905);
xnor U30204 (N_30204,N_29729,N_29948);
and U30205 (N_30205,N_29818,N_29728);
nor U30206 (N_30206,N_29543,N_29995);
nand U30207 (N_30207,N_29767,N_29830);
nand U30208 (N_30208,N_29552,N_29630);
xnor U30209 (N_30209,N_29880,N_29716);
nor U30210 (N_30210,N_29833,N_29596);
and U30211 (N_30211,N_29859,N_29745);
nor U30212 (N_30212,N_29656,N_29742);
xnor U30213 (N_30213,N_29967,N_29876);
nand U30214 (N_30214,N_29958,N_29924);
or U30215 (N_30215,N_29973,N_29650);
xor U30216 (N_30216,N_29700,N_29649);
and U30217 (N_30217,N_29768,N_29843);
xor U30218 (N_30218,N_29977,N_29554);
nor U30219 (N_30219,N_29614,N_29943);
nor U30220 (N_30220,N_29685,N_29514);
or U30221 (N_30221,N_29673,N_29563);
or U30222 (N_30222,N_29741,N_29532);
and U30223 (N_30223,N_29530,N_29590);
nand U30224 (N_30224,N_29969,N_29618);
nor U30225 (N_30225,N_29508,N_29886);
nand U30226 (N_30226,N_29975,N_29763);
or U30227 (N_30227,N_29622,N_29910);
and U30228 (N_30228,N_29953,N_29749);
xnor U30229 (N_30229,N_29955,N_29586);
nor U30230 (N_30230,N_29518,N_29873);
and U30231 (N_30231,N_29500,N_29664);
nor U30232 (N_30232,N_29602,N_29785);
nand U30233 (N_30233,N_29557,N_29874);
or U30234 (N_30234,N_29556,N_29611);
and U30235 (N_30235,N_29706,N_29803);
or U30236 (N_30236,N_29764,N_29612);
xnor U30237 (N_30237,N_29906,N_29724);
nand U30238 (N_30238,N_29692,N_29760);
and U30239 (N_30239,N_29595,N_29753);
xor U30240 (N_30240,N_29856,N_29926);
nor U30241 (N_30241,N_29525,N_29683);
or U30242 (N_30242,N_29726,N_29735);
nand U30243 (N_30243,N_29565,N_29894);
nand U30244 (N_30244,N_29624,N_29961);
nand U30245 (N_30245,N_29850,N_29860);
and U30246 (N_30246,N_29825,N_29569);
nand U30247 (N_30247,N_29617,N_29648);
nand U30248 (N_30248,N_29796,N_29580);
and U30249 (N_30249,N_29577,N_29829);
xnor U30250 (N_30250,N_29785,N_29965);
nor U30251 (N_30251,N_29822,N_29552);
nand U30252 (N_30252,N_29532,N_29661);
nand U30253 (N_30253,N_29681,N_29569);
xor U30254 (N_30254,N_29763,N_29701);
nand U30255 (N_30255,N_29686,N_29980);
nand U30256 (N_30256,N_29746,N_29707);
and U30257 (N_30257,N_29861,N_29886);
or U30258 (N_30258,N_29541,N_29754);
nor U30259 (N_30259,N_29903,N_29827);
and U30260 (N_30260,N_29653,N_29714);
nor U30261 (N_30261,N_29902,N_29721);
and U30262 (N_30262,N_29974,N_29510);
xor U30263 (N_30263,N_29522,N_29943);
or U30264 (N_30264,N_29723,N_29685);
nand U30265 (N_30265,N_29638,N_29682);
nor U30266 (N_30266,N_29550,N_29824);
or U30267 (N_30267,N_29757,N_29845);
xor U30268 (N_30268,N_29851,N_29840);
nor U30269 (N_30269,N_29763,N_29812);
nand U30270 (N_30270,N_29655,N_29546);
and U30271 (N_30271,N_29884,N_29997);
nand U30272 (N_30272,N_29885,N_29882);
nor U30273 (N_30273,N_29873,N_29760);
and U30274 (N_30274,N_29664,N_29886);
and U30275 (N_30275,N_29987,N_29808);
nand U30276 (N_30276,N_29562,N_29790);
nor U30277 (N_30277,N_29638,N_29684);
and U30278 (N_30278,N_29826,N_29682);
nor U30279 (N_30279,N_29855,N_29885);
and U30280 (N_30280,N_29794,N_29563);
nor U30281 (N_30281,N_29845,N_29985);
or U30282 (N_30282,N_29918,N_29873);
or U30283 (N_30283,N_29701,N_29804);
nand U30284 (N_30284,N_29866,N_29826);
xor U30285 (N_30285,N_29560,N_29879);
and U30286 (N_30286,N_29882,N_29968);
and U30287 (N_30287,N_29985,N_29888);
nand U30288 (N_30288,N_29900,N_29880);
or U30289 (N_30289,N_29621,N_29742);
nand U30290 (N_30290,N_29936,N_29949);
and U30291 (N_30291,N_29695,N_29990);
and U30292 (N_30292,N_29588,N_29611);
and U30293 (N_30293,N_29657,N_29663);
nand U30294 (N_30294,N_29959,N_29727);
and U30295 (N_30295,N_29508,N_29658);
nor U30296 (N_30296,N_29939,N_29716);
nor U30297 (N_30297,N_29993,N_29558);
or U30298 (N_30298,N_29661,N_29764);
nand U30299 (N_30299,N_29541,N_29940);
and U30300 (N_30300,N_29664,N_29972);
or U30301 (N_30301,N_29786,N_29663);
and U30302 (N_30302,N_29762,N_29993);
nor U30303 (N_30303,N_29632,N_29629);
and U30304 (N_30304,N_29882,N_29646);
and U30305 (N_30305,N_29533,N_29974);
nand U30306 (N_30306,N_29816,N_29633);
nand U30307 (N_30307,N_29703,N_29976);
and U30308 (N_30308,N_29672,N_29955);
nor U30309 (N_30309,N_29993,N_29505);
nor U30310 (N_30310,N_29666,N_29866);
xor U30311 (N_30311,N_29776,N_29892);
nor U30312 (N_30312,N_29911,N_29770);
or U30313 (N_30313,N_29520,N_29517);
nand U30314 (N_30314,N_29645,N_29941);
or U30315 (N_30315,N_29654,N_29713);
nand U30316 (N_30316,N_29581,N_29896);
and U30317 (N_30317,N_29709,N_29878);
xnor U30318 (N_30318,N_29730,N_29791);
or U30319 (N_30319,N_29835,N_29689);
and U30320 (N_30320,N_29693,N_29820);
nor U30321 (N_30321,N_29523,N_29925);
nor U30322 (N_30322,N_29959,N_29799);
and U30323 (N_30323,N_29634,N_29852);
nand U30324 (N_30324,N_29774,N_29669);
nor U30325 (N_30325,N_29983,N_29521);
or U30326 (N_30326,N_29689,N_29966);
nor U30327 (N_30327,N_29795,N_29566);
nand U30328 (N_30328,N_29541,N_29830);
or U30329 (N_30329,N_29649,N_29739);
xor U30330 (N_30330,N_29966,N_29753);
and U30331 (N_30331,N_29634,N_29529);
nand U30332 (N_30332,N_29955,N_29595);
nor U30333 (N_30333,N_29855,N_29752);
or U30334 (N_30334,N_29672,N_29590);
or U30335 (N_30335,N_29768,N_29535);
nand U30336 (N_30336,N_29606,N_29838);
nor U30337 (N_30337,N_29783,N_29652);
xnor U30338 (N_30338,N_29741,N_29884);
nor U30339 (N_30339,N_29552,N_29609);
nor U30340 (N_30340,N_29732,N_29543);
nor U30341 (N_30341,N_29750,N_29927);
or U30342 (N_30342,N_29672,N_29519);
nor U30343 (N_30343,N_29562,N_29526);
and U30344 (N_30344,N_29546,N_29576);
and U30345 (N_30345,N_29567,N_29845);
nand U30346 (N_30346,N_29725,N_29907);
nor U30347 (N_30347,N_29704,N_29808);
nor U30348 (N_30348,N_29913,N_29876);
nand U30349 (N_30349,N_29774,N_29658);
nand U30350 (N_30350,N_29917,N_29905);
nand U30351 (N_30351,N_29803,N_29509);
nand U30352 (N_30352,N_29991,N_29526);
nand U30353 (N_30353,N_29633,N_29878);
nand U30354 (N_30354,N_29787,N_29505);
nor U30355 (N_30355,N_29974,N_29732);
nor U30356 (N_30356,N_29716,N_29500);
or U30357 (N_30357,N_29967,N_29579);
nand U30358 (N_30358,N_29893,N_29922);
nor U30359 (N_30359,N_29682,N_29750);
and U30360 (N_30360,N_29689,N_29593);
nand U30361 (N_30361,N_29575,N_29636);
and U30362 (N_30362,N_29840,N_29570);
or U30363 (N_30363,N_29860,N_29764);
nor U30364 (N_30364,N_29976,N_29773);
nor U30365 (N_30365,N_29845,N_29647);
and U30366 (N_30366,N_29503,N_29880);
nor U30367 (N_30367,N_29554,N_29879);
xor U30368 (N_30368,N_29530,N_29787);
or U30369 (N_30369,N_29762,N_29709);
and U30370 (N_30370,N_29904,N_29554);
nand U30371 (N_30371,N_29885,N_29813);
nand U30372 (N_30372,N_29792,N_29522);
or U30373 (N_30373,N_29967,N_29762);
nand U30374 (N_30374,N_29846,N_29969);
nand U30375 (N_30375,N_29506,N_29560);
nand U30376 (N_30376,N_29937,N_29571);
nand U30377 (N_30377,N_29795,N_29710);
or U30378 (N_30378,N_29746,N_29754);
nor U30379 (N_30379,N_29969,N_29523);
xor U30380 (N_30380,N_29921,N_29929);
nor U30381 (N_30381,N_29971,N_29755);
nor U30382 (N_30382,N_29654,N_29904);
xor U30383 (N_30383,N_29721,N_29527);
or U30384 (N_30384,N_29667,N_29769);
nand U30385 (N_30385,N_29750,N_29619);
nor U30386 (N_30386,N_29668,N_29618);
nand U30387 (N_30387,N_29671,N_29746);
xor U30388 (N_30388,N_29717,N_29713);
xnor U30389 (N_30389,N_29670,N_29887);
xor U30390 (N_30390,N_29861,N_29994);
xor U30391 (N_30391,N_29882,N_29652);
or U30392 (N_30392,N_29566,N_29525);
nand U30393 (N_30393,N_29780,N_29661);
or U30394 (N_30394,N_29604,N_29762);
nand U30395 (N_30395,N_29751,N_29553);
nand U30396 (N_30396,N_29982,N_29930);
nor U30397 (N_30397,N_29773,N_29592);
nand U30398 (N_30398,N_29663,N_29990);
nand U30399 (N_30399,N_29697,N_29850);
nor U30400 (N_30400,N_29597,N_29513);
and U30401 (N_30401,N_29585,N_29623);
and U30402 (N_30402,N_29654,N_29888);
xnor U30403 (N_30403,N_29991,N_29905);
nor U30404 (N_30404,N_29953,N_29819);
or U30405 (N_30405,N_29636,N_29647);
and U30406 (N_30406,N_29837,N_29854);
and U30407 (N_30407,N_29955,N_29563);
nor U30408 (N_30408,N_29724,N_29765);
and U30409 (N_30409,N_29717,N_29914);
xor U30410 (N_30410,N_29644,N_29838);
and U30411 (N_30411,N_29582,N_29555);
or U30412 (N_30412,N_29501,N_29911);
nand U30413 (N_30413,N_29799,N_29712);
nand U30414 (N_30414,N_29987,N_29887);
nand U30415 (N_30415,N_29767,N_29969);
nand U30416 (N_30416,N_29766,N_29710);
nand U30417 (N_30417,N_29561,N_29529);
and U30418 (N_30418,N_29953,N_29519);
nor U30419 (N_30419,N_29652,N_29951);
xor U30420 (N_30420,N_29520,N_29779);
xnor U30421 (N_30421,N_29918,N_29647);
nor U30422 (N_30422,N_29804,N_29782);
and U30423 (N_30423,N_29688,N_29821);
nor U30424 (N_30424,N_29995,N_29666);
or U30425 (N_30425,N_29727,N_29601);
xnor U30426 (N_30426,N_29858,N_29678);
and U30427 (N_30427,N_29730,N_29921);
nor U30428 (N_30428,N_29646,N_29553);
nor U30429 (N_30429,N_29809,N_29585);
nor U30430 (N_30430,N_29895,N_29825);
nand U30431 (N_30431,N_29784,N_29597);
and U30432 (N_30432,N_29584,N_29917);
nor U30433 (N_30433,N_29996,N_29751);
nand U30434 (N_30434,N_29861,N_29628);
or U30435 (N_30435,N_29979,N_29654);
nand U30436 (N_30436,N_29948,N_29927);
nor U30437 (N_30437,N_29798,N_29719);
nand U30438 (N_30438,N_29707,N_29840);
xnor U30439 (N_30439,N_29534,N_29966);
nand U30440 (N_30440,N_29944,N_29683);
nand U30441 (N_30441,N_29576,N_29688);
and U30442 (N_30442,N_29810,N_29743);
xor U30443 (N_30443,N_29831,N_29783);
and U30444 (N_30444,N_29880,N_29847);
and U30445 (N_30445,N_29507,N_29794);
nor U30446 (N_30446,N_29932,N_29548);
or U30447 (N_30447,N_29875,N_29702);
nor U30448 (N_30448,N_29985,N_29700);
and U30449 (N_30449,N_29760,N_29522);
or U30450 (N_30450,N_29687,N_29971);
nand U30451 (N_30451,N_29998,N_29658);
xnor U30452 (N_30452,N_29740,N_29642);
and U30453 (N_30453,N_29770,N_29768);
or U30454 (N_30454,N_29545,N_29660);
xor U30455 (N_30455,N_29561,N_29955);
or U30456 (N_30456,N_29638,N_29888);
xnor U30457 (N_30457,N_29716,N_29944);
nand U30458 (N_30458,N_29988,N_29969);
or U30459 (N_30459,N_29547,N_29850);
or U30460 (N_30460,N_29908,N_29583);
or U30461 (N_30461,N_29748,N_29829);
or U30462 (N_30462,N_29568,N_29895);
nor U30463 (N_30463,N_29548,N_29994);
xnor U30464 (N_30464,N_29592,N_29838);
nand U30465 (N_30465,N_29786,N_29822);
nand U30466 (N_30466,N_29911,N_29802);
or U30467 (N_30467,N_29816,N_29812);
or U30468 (N_30468,N_29732,N_29953);
or U30469 (N_30469,N_29977,N_29892);
nand U30470 (N_30470,N_29704,N_29668);
or U30471 (N_30471,N_29883,N_29548);
and U30472 (N_30472,N_29881,N_29733);
nand U30473 (N_30473,N_29653,N_29759);
nand U30474 (N_30474,N_29585,N_29672);
xor U30475 (N_30475,N_29500,N_29762);
or U30476 (N_30476,N_29535,N_29686);
and U30477 (N_30477,N_29637,N_29701);
nand U30478 (N_30478,N_29956,N_29641);
and U30479 (N_30479,N_29501,N_29582);
or U30480 (N_30480,N_29595,N_29743);
nand U30481 (N_30481,N_29611,N_29999);
or U30482 (N_30482,N_29837,N_29510);
or U30483 (N_30483,N_29855,N_29695);
xnor U30484 (N_30484,N_29914,N_29975);
and U30485 (N_30485,N_29859,N_29730);
or U30486 (N_30486,N_29861,N_29578);
and U30487 (N_30487,N_29504,N_29700);
or U30488 (N_30488,N_29914,N_29672);
and U30489 (N_30489,N_29817,N_29625);
and U30490 (N_30490,N_29512,N_29541);
and U30491 (N_30491,N_29714,N_29931);
or U30492 (N_30492,N_29545,N_29750);
or U30493 (N_30493,N_29551,N_29892);
nor U30494 (N_30494,N_29926,N_29940);
nand U30495 (N_30495,N_29548,N_29501);
nand U30496 (N_30496,N_29547,N_29924);
nor U30497 (N_30497,N_29632,N_29944);
and U30498 (N_30498,N_29908,N_29787);
xor U30499 (N_30499,N_29697,N_29686);
nand U30500 (N_30500,N_30072,N_30338);
or U30501 (N_30501,N_30140,N_30025);
nand U30502 (N_30502,N_30288,N_30131);
or U30503 (N_30503,N_30396,N_30371);
xnor U30504 (N_30504,N_30239,N_30382);
nor U30505 (N_30505,N_30180,N_30185);
nor U30506 (N_30506,N_30093,N_30473);
nand U30507 (N_30507,N_30437,N_30449);
or U30508 (N_30508,N_30499,N_30399);
and U30509 (N_30509,N_30061,N_30033);
xor U30510 (N_30510,N_30422,N_30106);
xnor U30511 (N_30511,N_30290,N_30209);
and U30512 (N_30512,N_30087,N_30038);
or U30513 (N_30513,N_30293,N_30126);
or U30514 (N_30514,N_30109,N_30323);
nor U30515 (N_30515,N_30245,N_30156);
nand U30516 (N_30516,N_30212,N_30194);
nor U30517 (N_30517,N_30283,N_30363);
nor U30518 (N_30518,N_30259,N_30280);
xor U30519 (N_30519,N_30099,N_30011);
and U30520 (N_30520,N_30378,N_30297);
or U30521 (N_30521,N_30240,N_30308);
nor U30522 (N_30522,N_30215,N_30276);
nand U30523 (N_30523,N_30368,N_30309);
nand U30524 (N_30524,N_30429,N_30151);
nor U30525 (N_30525,N_30157,N_30265);
nor U30526 (N_30526,N_30301,N_30486);
nor U30527 (N_30527,N_30487,N_30386);
nand U30528 (N_30528,N_30128,N_30319);
xor U30529 (N_30529,N_30235,N_30342);
nand U30530 (N_30530,N_30497,N_30067);
nor U30531 (N_30531,N_30136,N_30475);
and U30532 (N_30532,N_30381,N_30451);
nand U30533 (N_30533,N_30158,N_30398);
or U30534 (N_30534,N_30271,N_30188);
nor U30535 (N_30535,N_30218,N_30171);
or U30536 (N_30536,N_30431,N_30257);
nor U30537 (N_30537,N_30272,N_30270);
or U30538 (N_30538,N_30095,N_30494);
xnor U30539 (N_30539,N_30457,N_30329);
nand U30540 (N_30540,N_30123,N_30455);
nand U30541 (N_30541,N_30263,N_30222);
nor U30542 (N_30542,N_30146,N_30178);
and U30543 (N_30543,N_30223,N_30278);
nand U30544 (N_30544,N_30167,N_30445);
and U30545 (N_30545,N_30474,N_30419);
nor U30546 (N_30546,N_30277,N_30393);
and U30547 (N_30547,N_30054,N_30037);
xnor U30548 (N_30548,N_30010,N_30485);
or U30549 (N_30549,N_30339,N_30217);
nand U30550 (N_30550,N_30410,N_30361);
and U30551 (N_30551,N_30441,N_30048);
nor U30552 (N_30552,N_30482,N_30089);
or U30553 (N_30553,N_30456,N_30112);
nor U30554 (N_30554,N_30160,N_30478);
nor U30555 (N_30555,N_30143,N_30114);
and U30556 (N_30556,N_30241,N_30039);
nor U30557 (N_30557,N_30227,N_30274);
nand U30558 (N_30558,N_30450,N_30207);
nor U30559 (N_30559,N_30104,N_30284);
nand U30560 (N_30560,N_30029,N_30017);
or U30561 (N_30561,N_30059,N_30150);
nor U30562 (N_30562,N_30032,N_30056);
nand U30563 (N_30563,N_30145,N_30229);
or U30564 (N_30564,N_30460,N_30330);
or U30565 (N_30565,N_30233,N_30074);
or U30566 (N_30566,N_30020,N_30395);
or U30567 (N_30567,N_30190,N_30357);
nor U30568 (N_30568,N_30332,N_30163);
nor U30569 (N_30569,N_30124,N_30314);
or U30570 (N_30570,N_30362,N_30458);
nand U30571 (N_30571,N_30287,N_30211);
or U30572 (N_30572,N_30387,N_30289);
and U30573 (N_30573,N_30453,N_30462);
or U30574 (N_30574,N_30351,N_30137);
or U30575 (N_30575,N_30465,N_30484);
and U30576 (N_30576,N_30367,N_30385);
and U30577 (N_30577,N_30333,N_30310);
and U30578 (N_30578,N_30053,N_30463);
and U30579 (N_30579,N_30366,N_30414);
or U30580 (N_30580,N_30097,N_30083);
or U30581 (N_30581,N_30466,N_30344);
and U30582 (N_30582,N_30448,N_30258);
nor U30583 (N_30583,N_30173,N_30108);
nand U30584 (N_30584,N_30380,N_30237);
xor U30585 (N_30585,N_30063,N_30049);
or U30586 (N_30586,N_30320,N_30423);
or U30587 (N_30587,N_30243,N_30015);
nor U30588 (N_30588,N_30321,N_30070);
nand U30589 (N_30589,N_30082,N_30267);
nor U30590 (N_30590,N_30428,N_30088);
nand U30591 (N_30591,N_30420,N_30296);
and U30592 (N_30592,N_30328,N_30447);
or U30593 (N_30593,N_30213,N_30129);
and U30594 (N_30594,N_30149,N_30075);
and U30595 (N_30595,N_30078,N_30165);
nor U30596 (N_30596,N_30182,N_30230);
xor U30597 (N_30597,N_30370,N_30418);
nand U30598 (N_30598,N_30306,N_30169);
xor U30599 (N_30599,N_30477,N_30302);
and U30600 (N_30600,N_30000,N_30312);
or U30601 (N_30601,N_30242,N_30216);
and U30602 (N_30602,N_30350,N_30353);
and U30603 (N_30603,N_30291,N_30413);
nor U30604 (N_30604,N_30231,N_30042);
nand U30605 (N_30605,N_30476,N_30341);
or U30606 (N_30606,N_30246,N_30379);
or U30607 (N_30607,N_30408,N_30050);
or U30608 (N_30608,N_30102,N_30299);
nand U30609 (N_30609,N_30044,N_30345);
nand U30610 (N_30610,N_30421,N_30135);
or U30611 (N_30611,N_30094,N_30286);
nor U30612 (N_30612,N_30252,N_30498);
or U30613 (N_30613,N_30427,N_30161);
nor U30614 (N_30614,N_30077,N_30004);
or U30615 (N_30615,N_30183,N_30406);
and U30616 (N_30616,N_30111,N_30226);
and U30617 (N_30617,N_30193,N_30110);
or U30618 (N_30618,N_30266,N_30355);
nand U30619 (N_30619,N_30006,N_30069);
nor U30620 (N_30620,N_30384,N_30253);
nand U30621 (N_30621,N_30142,N_30304);
nand U30622 (N_30622,N_30496,N_30426);
or U30623 (N_30623,N_30365,N_30411);
and U30624 (N_30624,N_30347,N_30214);
and U30625 (N_30625,N_30247,N_30184);
nand U30626 (N_30626,N_30046,N_30176);
xnor U30627 (N_30627,N_30018,N_30402);
nor U30628 (N_30628,N_30096,N_30373);
xnor U30629 (N_30629,N_30461,N_30022);
or U30630 (N_30630,N_30250,N_30221);
nor U30631 (N_30631,N_30005,N_30442);
nor U30632 (N_30632,N_30260,N_30115);
xnor U30633 (N_30633,N_30138,N_30224);
and U30634 (N_30634,N_30051,N_30202);
and U30635 (N_30635,N_30407,N_30043);
nand U30636 (N_30636,N_30040,N_30027);
nor U30637 (N_30637,N_30269,N_30187);
nor U30638 (N_30638,N_30489,N_30443);
or U30639 (N_30639,N_30275,N_30092);
and U30640 (N_30640,N_30228,N_30264);
nand U30641 (N_30641,N_30196,N_30117);
and U30642 (N_30642,N_30469,N_30392);
nor U30643 (N_30643,N_30295,N_30483);
nand U30644 (N_30644,N_30348,N_30454);
or U30645 (N_30645,N_30085,N_30389);
nand U30646 (N_30646,N_30132,N_30472);
and U30647 (N_30647,N_30175,N_30107);
nand U30648 (N_30648,N_30101,N_30424);
and U30649 (N_30649,N_30444,N_30086);
xnor U30650 (N_30650,N_30007,N_30438);
xnor U30651 (N_30651,N_30327,N_30134);
and U30652 (N_30652,N_30377,N_30208);
and U30653 (N_30653,N_30139,N_30415);
and U30654 (N_30654,N_30446,N_30023);
and U30655 (N_30655,N_30273,N_30019);
or U30656 (N_30656,N_30383,N_30325);
or U30657 (N_30657,N_30113,N_30204);
nand U30658 (N_30658,N_30153,N_30219);
or U30659 (N_30659,N_30249,N_30390);
and U30660 (N_30660,N_30491,N_30152);
or U30661 (N_30661,N_30232,N_30292);
xnor U30662 (N_30662,N_30154,N_30008);
nor U30663 (N_30663,N_30002,N_30026);
xnor U30664 (N_30664,N_30354,N_30014);
and U30665 (N_30665,N_30116,N_30452);
nor U30666 (N_30666,N_30303,N_30065);
nor U30667 (N_30667,N_30311,N_30066);
nand U30668 (N_30668,N_30166,N_30047);
nand U30669 (N_30669,N_30103,N_30073);
nand U30670 (N_30670,N_30409,N_30125);
and U30671 (N_30671,N_30028,N_30021);
and U30672 (N_30672,N_30034,N_30013);
and U30673 (N_30673,N_30220,N_30331);
nand U30674 (N_30674,N_30493,N_30261);
nor U30675 (N_30675,N_30076,N_30360);
nor U30676 (N_30676,N_30440,N_30436);
and U30677 (N_30677,N_30236,N_30324);
nor U30678 (N_30678,N_30343,N_30003);
nand U30679 (N_30679,N_30201,N_30159);
nand U30680 (N_30680,N_30467,N_30009);
nand U30681 (N_30681,N_30434,N_30198);
nand U30682 (N_30682,N_30045,N_30100);
or U30683 (N_30683,N_30471,N_30412);
xor U30684 (N_30684,N_30244,N_30254);
xnor U30685 (N_30685,N_30459,N_30359);
or U30686 (N_30686,N_30133,N_30481);
nor U30687 (N_30687,N_30480,N_30401);
nor U30688 (N_30688,N_30064,N_30326);
nand U30689 (N_30689,N_30144,N_30234);
and U30690 (N_30690,N_30118,N_30195);
and U30691 (N_30691,N_30369,N_30335);
and U30692 (N_30692,N_30001,N_30349);
or U30693 (N_30693,N_30430,N_30425);
nor U30694 (N_30694,N_30294,N_30179);
or U30695 (N_30695,N_30305,N_30432);
nand U30696 (N_30696,N_30417,N_30256);
or U30697 (N_30697,N_30238,N_30318);
nand U30698 (N_30698,N_30041,N_30439);
nand U30699 (N_30699,N_30285,N_30334);
or U30700 (N_30700,N_30036,N_30192);
and U30701 (N_30701,N_30358,N_30174);
or U30702 (N_30702,N_30336,N_30162);
nand U30703 (N_30703,N_30388,N_30376);
or U30704 (N_30704,N_30281,N_30079);
and U30705 (N_30705,N_30322,N_30168);
xnor U30706 (N_30706,N_30164,N_30203);
or U30707 (N_30707,N_30375,N_30121);
nand U30708 (N_30708,N_30364,N_30081);
nand U30709 (N_30709,N_30391,N_30404);
and U30710 (N_30710,N_30197,N_30090);
or U30711 (N_30711,N_30468,N_30313);
or U30712 (N_30712,N_30105,N_30057);
xnor U30713 (N_30713,N_30120,N_30170);
nand U30714 (N_30714,N_30300,N_30058);
and U30715 (N_30715,N_30433,N_30127);
xor U30716 (N_30716,N_30394,N_30372);
nor U30717 (N_30717,N_30262,N_30470);
nand U30718 (N_30718,N_30405,N_30298);
or U30719 (N_30719,N_30282,N_30397);
xnor U30720 (N_30720,N_30030,N_30122);
xor U30721 (N_30721,N_30316,N_30416);
nor U30722 (N_30722,N_30479,N_30248);
and U30723 (N_30723,N_30490,N_30181);
or U30724 (N_30724,N_30210,N_30403);
nand U30725 (N_30725,N_30464,N_30186);
nand U30726 (N_30726,N_30225,N_30346);
nor U30727 (N_30727,N_30307,N_30031);
xnor U30728 (N_30728,N_30012,N_30172);
nand U30729 (N_30729,N_30148,N_30119);
and U30730 (N_30730,N_30060,N_30199);
or U30731 (N_30731,N_30024,N_30098);
and U30732 (N_30732,N_30062,N_30255);
and U30733 (N_30733,N_30141,N_30279);
or U30734 (N_30734,N_30205,N_30130);
xor U30735 (N_30735,N_30071,N_30435);
and U30736 (N_30736,N_30356,N_30315);
nor U30737 (N_30737,N_30317,N_30147);
or U30738 (N_30738,N_30080,N_30400);
nor U30739 (N_30739,N_30268,N_30177);
nor U30740 (N_30740,N_30337,N_30488);
nor U30741 (N_30741,N_30084,N_30206);
and U30742 (N_30742,N_30016,N_30191);
or U30743 (N_30743,N_30055,N_30155);
or U30744 (N_30744,N_30052,N_30374);
nor U30745 (N_30745,N_30495,N_30200);
nor U30746 (N_30746,N_30189,N_30251);
and U30747 (N_30747,N_30035,N_30068);
and U30748 (N_30748,N_30091,N_30340);
nor U30749 (N_30749,N_30352,N_30492);
nand U30750 (N_30750,N_30299,N_30304);
nand U30751 (N_30751,N_30164,N_30303);
or U30752 (N_30752,N_30485,N_30017);
nor U30753 (N_30753,N_30402,N_30395);
nand U30754 (N_30754,N_30042,N_30072);
nor U30755 (N_30755,N_30111,N_30307);
or U30756 (N_30756,N_30235,N_30201);
nor U30757 (N_30757,N_30102,N_30118);
nand U30758 (N_30758,N_30231,N_30215);
nand U30759 (N_30759,N_30477,N_30171);
and U30760 (N_30760,N_30077,N_30310);
nand U30761 (N_30761,N_30449,N_30439);
or U30762 (N_30762,N_30312,N_30111);
and U30763 (N_30763,N_30261,N_30378);
nand U30764 (N_30764,N_30448,N_30405);
nand U30765 (N_30765,N_30238,N_30357);
nor U30766 (N_30766,N_30117,N_30338);
and U30767 (N_30767,N_30415,N_30160);
or U30768 (N_30768,N_30483,N_30493);
or U30769 (N_30769,N_30019,N_30428);
nor U30770 (N_30770,N_30129,N_30145);
or U30771 (N_30771,N_30125,N_30444);
nand U30772 (N_30772,N_30243,N_30440);
and U30773 (N_30773,N_30023,N_30184);
nand U30774 (N_30774,N_30392,N_30190);
nor U30775 (N_30775,N_30269,N_30413);
or U30776 (N_30776,N_30357,N_30179);
and U30777 (N_30777,N_30489,N_30226);
xor U30778 (N_30778,N_30120,N_30369);
or U30779 (N_30779,N_30066,N_30262);
nor U30780 (N_30780,N_30294,N_30118);
and U30781 (N_30781,N_30269,N_30346);
or U30782 (N_30782,N_30293,N_30070);
nor U30783 (N_30783,N_30016,N_30070);
xor U30784 (N_30784,N_30499,N_30411);
or U30785 (N_30785,N_30284,N_30216);
and U30786 (N_30786,N_30485,N_30344);
nand U30787 (N_30787,N_30403,N_30302);
and U30788 (N_30788,N_30344,N_30056);
nor U30789 (N_30789,N_30497,N_30223);
nand U30790 (N_30790,N_30058,N_30395);
nor U30791 (N_30791,N_30355,N_30443);
xor U30792 (N_30792,N_30061,N_30020);
and U30793 (N_30793,N_30016,N_30312);
and U30794 (N_30794,N_30028,N_30325);
and U30795 (N_30795,N_30267,N_30435);
xor U30796 (N_30796,N_30043,N_30476);
nand U30797 (N_30797,N_30095,N_30433);
nand U30798 (N_30798,N_30311,N_30069);
nor U30799 (N_30799,N_30140,N_30001);
nor U30800 (N_30800,N_30254,N_30255);
nand U30801 (N_30801,N_30014,N_30374);
nand U30802 (N_30802,N_30076,N_30496);
or U30803 (N_30803,N_30049,N_30012);
nor U30804 (N_30804,N_30341,N_30009);
nand U30805 (N_30805,N_30476,N_30321);
nand U30806 (N_30806,N_30316,N_30093);
and U30807 (N_30807,N_30200,N_30215);
and U30808 (N_30808,N_30041,N_30434);
nor U30809 (N_30809,N_30279,N_30153);
nand U30810 (N_30810,N_30082,N_30123);
and U30811 (N_30811,N_30429,N_30026);
nand U30812 (N_30812,N_30109,N_30063);
nand U30813 (N_30813,N_30162,N_30002);
nor U30814 (N_30814,N_30474,N_30478);
nor U30815 (N_30815,N_30340,N_30108);
nor U30816 (N_30816,N_30089,N_30267);
or U30817 (N_30817,N_30419,N_30242);
nand U30818 (N_30818,N_30018,N_30472);
or U30819 (N_30819,N_30188,N_30419);
or U30820 (N_30820,N_30349,N_30031);
or U30821 (N_30821,N_30418,N_30347);
xnor U30822 (N_30822,N_30113,N_30091);
and U30823 (N_30823,N_30460,N_30245);
and U30824 (N_30824,N_30121,N_30245);
or U30825 (N_30825,N_30134,N_30264);
nand U30826 (N_30826,N_30064,N_30389);
nor U30827 (N_30827,N_30341,N_30008);
and U30828 (N_30828,N_30034,N_30086);
and U30829 (N_30829,N_30317,N_30415);
nand U30830 (N_30830,N_30127,N_30184);
nor U30831 (N_30831,N_30498,N_30259);
nor U30832 (N_30832,N_30102,N_30233);
nor U30833 (N_30833,N_30407,N_30373);
or U30834 (N_30834,N_30093,N_30192);
nor U30835 (N_30835,N_30050,N_30119);
and U30836 (N_30836,N_30450,N_30081);
xor U30837 (N_30837,N_30074,N_30094);
or U30838 (N_30838,N_30394,N_30347);
or U30839 (N_30839,N_30333,N_30117);
xnor U30840 (N_30840,N_30498,N_30378);
nor U30841 (N_30841,N_30175,N_30486);
and U30842 (N_30842,N_30010,N_30138);
nor U30843 (N_30843,N_30000,N_30486);
and U30844 (N_30844,N_30367,N_30280);
nand U30845 (N_30845,N_30300,N_30375);
and U30846 (N_30846,N_30214,N_30389);
nor U30847 (N_30847,N_30180,N_30353);
and U30848 (N_30848,N_30288,N_30336);
xnor U30849 (N_30849,N_30156,N_30005);
nor U30850 (N_30850,N_30279,N_30329);
xor U30851 (N_30851,N_30400,N_30410);
nand U30852 (N_30852,N_30075,N_30435);
and U30853 (N_30853,N_30497,N_30088);
nor U30854 (N_30854,N_30100,N_30290);
nand U30855 (N_30855,N_30425,N_30410);
or U30856 (N_30856,N_30114,N_30164);
and U30857 (N_30857,N_30416,N_30129);
nand U30858 (N_30858,N_30481,N_30192);
nand U30859 (N_30859,N_30462,N_30232);
and U30860 (N_30860,N_30079,N_30065);
nor U30861 (N_30861,N_30256,N_30259);
nor U30862 (N_30862,N_30489,N_30129);
and U30863 (N_30863,N_30071,N_30049);
and U30864 (N_30864,N_30352,N_30390);
or U30865 (N_30865,N_30336,N_30003);
nor U30866 (N_30866,N_30173,N_30184);
nand U30867 (N_30867,N_30263,N_30409);
nand U30868 (N_30868,N_30184,N_30338);
or U30869 (N_30869,N_30184,N_30492);
or U30870 (N_30870,N_30028,N_30210);
nor U30871 (N_30871,N_30163,N_30349);
or U30872 (N_30872,N_30320,N_30177);
nand U30873 (N_30873,N_30438,N_30087);
nand U30874 (N_30874,N_30486,N_30443);
nor U30875 (N_30875,N_30018,N_30322);
and U30876 (N_30876,N_30281,N_30090);
nand U30877 (N_30877,N_30218,N_30370);
nand U30878 (N_30878,N_30241,N_30124);
xor U30879 (N_30879,N_30162,N_30385);
nand U30880 (N_30880,N_30047,N_30183);
or U30881 (N_30881,N_30297,N_30126);
nand U30882 (N_30882,N_30375,N_30457);
xor U30883 (N_30883,N_30045,N_30464);
xnor U30884 (N_30884,N_30480,N_30042);
and U30885 (N_30885,N_30089,N_30477);
or U30886 (N_30886,N_30486,N_30225);
and U30887 (N_30887,N_30206,N_30202);
nor U30888 (N_30888,N_30152,N_30202);
and U30889 (N_30889,N_30299,N_30143);
nand U30890 (N_30890,N_30070,N_30083);
nor U30891 (N_30891,N_30435,N_30486);
nor U30892 (N_30892,N_30115,N_30355);
and U30893 (N_30893,N_30492,N_30474);
or U30894 (N_30894,N_30488,N_30019);
nor U30895 (N_30895,N_30485,N_30333);
xor U30896 (N_30896,N_30414,N_30024);
nor U30897 (N_30897,N_30452,N_30126);
or U30898 (N_30898,N_30032,N_30171);
and U30899 (N_30899,N_30165,N_30350);
or U30900 (N_30900,N_30365,N_30454);
nor U30901 (N_30901,N_30017,N_30165);
and U30902 (N_30902,N_30044,N_30157);
nand U30903 (N_30903,N_30420,N_30162);
and U30904 (N_30904,N_30175,N_30326);
or U30905 (N_30905,N_30329,N_30267);
and U30906 (N_30906,N_30006,N_30397);
and U30907 (N_30907,N_30101,N_30350);
or U30908 (N_30908,N_30149,N_30240);
and U30909 (N_30909,N_30425,N_30023);
and U30910 (N_30910,N_30164,N_30127);
and U30911 (N_30911,N_30393,N_30144);
xor U30912 (N_30912,N_30327,N_30157);
or U30913 (N_30913,N_30037,N_30267);
nand U30914 (N_30914,N_30416,N_30232);
nor U30915 (N_30915,N_30259,N_30001);
xnor U30916 (N_30916,N_30301,N_30312);
xor U30917 (N_30917,N_30135,N_30465);
and U30918 (N_30918,N_30150,N_30186);
and U30919 (N_30919,N_30060,N_30018);
nand U30920 (N_30920,N_30454,N_30245);
nor U30921 (N_30921,N_30297,N_30302);
nand U30922 (N_30922,N_30251,N_30058);
nand U30923 (N_30923,N_30345,N_30301);
nand U30924 (N_30924,N_30094,N_30431);
nor U30925 (N_30925,N_30426,N_30247);
nand U30926 (N_30926,N_30186,N_30036);
nand U30927 (N_30927,N_30091,N_30372);
nand U30928 (N_30928,N_30399,N_30345);
and U30929 (N_30929,N_30108,N_30429);
nand U30930 (N_30930,N_30251,N_30481);
nand U30931 (N_30931,N_30049,N_30100);
or U30932 (N_30932,N_30435,N_30112);
nand U30933 (N_30933,N_30440,N_30206);
nor U30934 (N_30934,N_30301,N_30241);
and U30935 (N_30935,N_30230,N_30251);
or U30936 (N_30936,N_30129,N_30411);
or U30937 (N_30937,N_30271,N_30418);
and U30938 (N_30938,N_30131,N_30458);
and U30939 (N_30939,N_30369,N_30405);
nand U30940 (N_30940,N_30224,N_30049);
xor U30941 (N_30941,N_30495,N_30317);
nor U30942 (N_30942,N_30141,N_30225);
and U30943 (N_30943,N_30273,N_30454);
or U30944 (N_30944,N_30353,N_30204);
or U30945 (N_30945,N_30266,N_30302);
and U30946 (N_30946,N_30350,N_30045);
xor U30947 (N_30947,N_30274,N_30354);
and U30948 (N_30948,N_30289,N_30284);
and U30949 (N_30949,N_30393,N_30387);
nand U30950 (N_30950,N_30065,N_30339);
or U30951 (N_30951,N_30020,N_30216);
nor U30952 (N_30952,N_30194,N_30148);
or U30953 (N_30953,N_30385,N_30412);
nand U30954 (N_30954,N_30333,N_30299);
nor U30955 (N_30955,N_30102,N_30264);
nand U30956 (N_30956,N_30268,N_30015);
and U30957 (N_30957,N_30134,N_30295);
nor U30958 (N_30958,N_30417,N_30135);
nor U30959 (N_30959,N_30470,N_30055);
xor U30960 (N_30960,N_30268,N_30215);
and U30961 (N_30961,N_30303,N_30107);
nor U30962 (N_30962,N_30267,N_30187);
and U30963 (N_30963,N_30149,N_30391);
nand U30964 (N_30964,N_30035,N_30093);
nor U30965 (N_30965,N_30335,N_30358);
or U30966 (N_30966,N_30358,N_30244);
nand U30967 (N_30967,N_30422,N_30054);
nor U30968 (N_30968,N_30076,N_30315);
nor U30969 (N_30969,N_30430,N_30258);
nor U30970 (N_30970,N_30265,N_30171);
or U30971 (N_30971,N_30351,N_30352);
nand U30972 (N_30972,N_30422,N_30250);
nand U30973 (N_30973,N_30139,N_30322);
or U30974 (N_30974,N_30001,N_30316);
and U30975 (N_30975,N_30131,N_30462);
and U30976 (N_30976,N_30193,N_30425);
and U30977 (N_30977,N_30007,N_30266);
or U30978 (N_30978,N_30385,N_30422);
xor U30979 (N_30979,N_30344,N_30283);
nor U30980 (N_30980,N_30350,N_30335);
or U30981 (N_30981,N_30151,N_30183);
nor U30982 (N_30982,N_30423,N_30231);
nand U30983 (N_30983,N_30480,N_30143);
nor U30984 (N_30984,N_30447,N_30056);
nand U30985 (N_30985,N_30245,N_30320);
nor U30986 (N_30986,N_30313,N_30303);
or U30987 (N_30987,N_30013,N_30460);
nand U30988 (N_30988,N_30487,N_30285);
nor U30989 (N_30989,N_30219,N_30192);
or U30990 (N_30990,N_30382,N_30249);
nand U30991 (N_30991,N_30448,N_30385);
nand U30992 (N_30992,N_30152,N_30337);
or U30993 (N_30993,N_30412,N_30495);
or U30994 (N_30994,N_30296,N_30314);
and U30995 (N_30995,N_30377,N_30035);
and U30996 (N_30996,N_30106,N_30201);
nor U30997 (N_30997,N_30083,N_30066);
xnor U30998 (N_30998,N_30150,N_30432);
nor U30999 (N_30999,N_30382,N_30457);
nor U31000 (N_31000,N_30771,N_30602);
nor U31001 (N_31001,N_30671,N_30815);
nor U31002 (N_31002,N_30797,N_30726);
nor U31003 (N_31003,N_30621,N_30606);
nand U31004 (N_31004,N_30552,N_30502);
nand U31005 (N_31005,N_30698,N_30584);
and U31006 (N_31006,N_30988,N_30569);
or U31007 (N_31007,N_30512,N_30919);
and U31008 (N_31008,N_30648,N_30731);
or U31009 (N_31009,N_30717,N_30948);
nand U31010 (N_31010,N_30761,N_30898);
and U31011 (N_31011,N_30923,N_30622);
and U31012 (N_31012,N_30715,N_30549);
and U31013 (N_31013,N_30810,N_30800);
nand U31014 (N_31014,N_30645,N_30708);
nor U31015 (N_31015,N_30792,N_30906);
nor U31016 (N_31016,N_30767,N_30755);
nor U31017 (N_31017,N_30694,N_30647);
nor U31018 (N_31018,N_30505,N_30588);
nand U31019 (N_31019,N_30951,N_30786);
xnor U31020 (N_31020,N_30553,N_30848);
nand U31021 (N_31021,N_30641,N_30738);
nor U31022 (N_31022,N_30974,N_30835);
or U31023 (N_31023,N_30904,N_30889);
nand U31024 (N_31024,N_30610,N_30633);
or U31025 (N_31025,N_30653,N_30691);
xnor U31026 (N_31026,N_30913,N_30750);
or U31027 (N_31027,N_30659,N_30541);
or U31028 (N_31028,N_30873,N_30916);
and U31029 (N_31029,N_30944,N_30687);
or U31030 (N_31030,N_30928,N_30530);
nand U31031 (N_31031,N_30837,N_30893);
nor U31032 (N_31032,N_30561,N_30508);
nand U31033 (N_31033,N_30853,N_30805);
nand U31034 (N_31034,N_30884,N_30878);
or U31035 (N_31035,N_30589,N_30583);
nor U31036 (N_31036,N_30918,N_30892);
nor U31037 (N_31037,N_30776,N_30763);
or U31038 (N_31038,N_30794,N_30960);
xor U31039 (N_31039,N_30592,N_30959);
or U31040 (N_31040,N_30877,N_30866);
nor U31041 (N_31041,N_30733,N_30790);
and U31042 (N_31042,N_30981,N_30526);
nand U31043 (N_31043,N_30768,N_30683);
nor U31044 (N_31044,N_30799,N_30545);
nor U31045 (N_31045,N_30780,N_30670);
nor U31046 (N_31046,N_30891,N_30743);
or U31047 (N_31047,N_30539,N_30876);
nor U31048 (N_31048,N_30858,N_30964);
nor U31049 (N_31049,N_30772,N_30535);
or U31050 (N_31050,N_30787,N_30663);
nor U31051 (N_31051,N_30826,N_30968);
nor U31052 (N_31052,N_30934,N_30806);
or U31053 (N_31053,N_30961,N_30516);
nor U31054 (N_31054,N_30735,N_30966);
nand U31055 (N_31055,N_30555,N_30989);
nor U31056 (N_31056,N_30596,N_30542);
and U31057 (N_31057,N_30572,N_30783);
nor U31058 (N_31058,N_30684,N_30534);
and U31059 (N_31059,N_30723,N_30804);
nand U31060 (N_31060,N_30649,N_30574);
and U31061 (N_31061,N_30947,N_30888);
and U31062 (N_31062,N_30700,N_30576);
nand U31063 (N_31063,N_30567,N_30887);
or U31064 (N_31064,N_30568,N_30655);
nor U31065 (N_31065,N_30896,N_30582);
and U31066 (N_31066,N_30527,N_30643);
nor U31067 (N_31067,N_30688,N_30886);
nor U31068 (N_31068,N_30519,N_30751);
nand U31069 (N_31069,N_30618,N_30611);
nor U31070 (N_31070,N_30920,N_30812);
and U31071 (N_31071,N_30737,N_30608);
or U31072 (N_31072,N_30669,N_30500);
nor U31073 (N_31073,N_30802,N_30970);
nor U31074 (N_31074,N_30976,N_30680);
nor U31075 (N_31075,N_30722,N_30521);
and U31076 (N_31076,N_30860,N_30556);
or U31077 (N_31077,N_30749,N_30693);
nor U31078 (N_31078,N_30739,N_30942);
xor U31079 (N_31079,N_30581,N_30836);
nor U31080 (N_31080,N_30808,N_30701);
nor U31081 (N_31081,N_30990,N_30511);
xnor U31082 (N_31082,N_30862,N_30779);
or U31083 (N_31083,N_30536,N_30875);
xor U31084 (N_31084,N_30965,N_30651);
or U31085 (N_31085,N_30832,N_30769);
nor U31086 (N_31086,N_30656,N_30632);
nor U31087 (N_31087,N_30562,N_30957);
or U31088 (N_31088,N_30544,N_30666);
nor U31089 (N_31089,N_30855,N_30984);
and U31090 (N_31090,N_30522,N_30793);
and U31091 (N_31091,N_30980,N_30996);
and U31092 (N_31092,N_30593,N_30977);
xnor U31093 (N_31093,N_30841,N_30969);
nor U31094 (N_31094,N_30658,N_30880);
or U31095 (N_31095,N_30842,N_30746);
or U31096 (N_31096,N_30897,N_30646);
nand U31097 (N_31097,N_30933,N_30624);
and U31098 (N_31098,N_30986,N_30564);
nand U31099 (N_31099,N_30774,N_30927);
xnor U31100 (N_31100,N_30570,N_30931);
and U31101 (N_31101,N_30538,N_30598);
and U31102 (N_31102,N_30932,N_30650);
xnor U31103 (N_31103,N_30908,N_30854);
xnor U31104 (N_31104,N_30910,N_30742);
nand U31105 (N_31105,N_30825,N_30798);
nand U31106 (N_31106,N_30637,N_30952);
nor U31107 (N_31107,N_30859,N_30506);
nor U31108 (N_31108,N_30631,N_30902);
or U31109 (N_31109,N_30660,N_30785);
and U31110 (N_31110,N_30662,N_30962);
nand U31111 (N_31111,N_30803,N_30504);
and U31112 (N_31112,N_30585,N_30849);
and U31113 (N_31113,N_30547,N_30953);
and U31114 (N_31114,N_30674,N_30972);
nor U31115 (N_31115,N_30741,N_30850);
or U31116 (N_31116,N_30635,N_30675);
or U31117 (N_31117,N_30559,N_30885);
xor U31118 (N_31118,N_30921,N_30525);
nand U31119 (N_31119,N_30946,N_30727);
and U31120 (N_31120,N_30725,N_30677);
nor U31121 (N_31121,N_30834,N_30955);
xnor U31122 (N_31122,N_30702,N_30587);
and U31123 (N_31123,N_30999,N_30846);
nor U31124 (N_31124,N_30938,N_30811);
and U31125 (N_31125,N_30578,N_30503);
nand U31126 (N_31126,N_30560,N_30668);
nand U31127 (N_31127,N_30550,N_30629);
and U31128 (N_31128,N_30992,N_30630);
nand U31129 (N_31129,N_30925,N_30626);
nand U31130 (N_31130,N_30609,N_30724);
and U31131 (N_31131,N_30642,N_30565);
and U31132 (N_31132,N_30987,N_30847);
and U31133 (N_31133,N_30732,N_30828);
nor U31134 (N_31134,N_30707,N_30807);
nand U31135 (N_31135,N_30801,N_30533);
nor U31136 (N_31136,N_30628,N_30730);
xnor U31137 (N_31137,N_30900,N_30905);
and U31138 (N_31138,N_30819,N_30845);
nand U31139 (N_31139,N_30672,N_30557);
nand U31140 (N_31140,N_30518,N_30685);
and U31141 (N_31141,N_30765,N_30781);
and U31142 (N_31142,N_30995,N_30940);
and U31143 (N_31143,N_30840,N_30580);
nand U31144 (N_31144,N_30958,N_30829);
or U31145 (N_31145,N_30571,N_30721);
xor U31146 (N_31146,N_30983,N_30788);
nor U31147 (N_31147,N_30754,N_30861);
nand U31148 (N_31148,N_30869,N_30759);
nand U31149 (N_31149,N_30736,N_30704);
xnor U31150 (N_31150,N_30782,N_30907);
or U31151 (N_31151,N_30915,N_30871);
or U31152 (N_31152,N_30554,N_30509);
and U31153 (N_31153,N_30757,N_30982);
or U31154 (N_31154,N_30752,N_30507);
xor U31155 (N_31155,N_30956,N_30716);
nand U31156 (N_31156,N_30856,N_30706);
or U31157 (N_31157,N_30558,N_30949);
and U31158 (N_31158,N_30531,N_30524);
or U31159 (N_31159,N_30978,N_30773);
nor U31160 (N_31160,N_30857,N_30625);
nor U31161 (N_31161,N_30528,N_30501);
nand U31162 (N_31162,N_30679,N_30764);
and U31163 (N_31163,N_30579,N_30546);
nand U31164 (N_31164,N_30822,N_30863);
or U31165 (N_31165,N_30520,N_30747);
nand U31166 (N_31166,N_30667,N_30634);
or U31167 (N_31167,N_30600,N_30657);
nand U31168 (N_31168,N_30939,N_30613);
nand U31169 (N_31169,N_30758,N_30770);
nand U31170 (N_31170,N_30686,N_30912);
and U31171 (N_31171,N_30678,N_30573);
nand U31172 (N_31172,N_30994,N_30895);
or U31173 (N_31173,N_30664,N_30720);
or U31174 (N_31174,N_30638,N_30831);
xnor U31175 (N_31175,N_30879,N_30605);
or U31176 (N_31176,N_30548,N_30639);
xnor U31177 (N_31177,N_30870,N_30813);
nor U31178 (N_31178,N_30963,N_30543);
xor U31179 (N_31179,N_30874,N_30839);
or U31180 (N_31180,N_30599,N_30523);
or U31181 (N_31181,N_30930,N_30917);
and U31182 (N_31182,N_30760,N_30690);
nor U31183 (N_31183,N_30971,N_30745);
nand U31184 (N_31184,N_30681,N_30899);
nor U31185 (N_31185,N_30601,N_30586);
nor U31186 (N_31186,N_30537,N_30775);
nor U31187 (N_31187,N_30766,N_30778);
nand U31188 (N_31188,N_30851,N_30838);
xnor U31189 (N_31189,N_30740,N_30914);
or U31190 (N_31190,N_30865,N_30619);
or U31191 (N_31191,N_30867,N_30709);
xor U31192 (N_31192,N_30777,N_30872);
and U31193 (N_31193,N_30513,N_30517);
and U31194 (N_31194,N_30591,N_30689);
nand U31195 (N_31195,N_30665,N_30590);
and U31196 (N_31196,N_30607,N_30644);
nand U31197 (N_31197,N_30551,N_30843);
or U31198 (N_31198,N_30936,N_30753);
or U31199 (N_31199,N_30729,N_30756);
nand U31200 (N_31200,N_30719,N_30911);
and U31201 (N_31201,N_30699,N_30926);
nand U31202 (N_31202,N_30950,N_30617);
nor U31203 (N_31203,N_30993,N_30814);
nand U31204 (N_31204,N_30827,N_30816);
nand U31205 (N_31205,N_30563,N_30823);
and U31206 (N_31206,N_30673,N_30935);
or U31207 (N_31207,N_30762,N_30575);
xnor U31208 (N_31208,N_30692,N_30973);
nor U31209 (N_31209,N_30954,N_30945);
xnor U31210 (N_31210,N_30728,N_30529);
and U31211 (N_31211,N_30710,N_30791);
nor U31212 (N_31212,N_30703,N_30909);
or U31213 (N_31213,N_30975,N_30795);
or U31214 (N_31214,N_30695,N_30682);
and U31215 (N_31215,N_30784,N_30929);
nand U31216 (N_31216,N_30614,N_30718);
and U31217 (N_31217,N_30943,N_30796);
and U31218 (N_31218,N_30821,N_30713);
nor U31219 (N_31219,N_30824,N_30937);
nand U31220 (N_31220,N_30833,N_30903);
and U31221 (N_31221,N_30820,N_30623);
nand U31222 (N_31222,N_30612,N_30510);
nand U31223 (N_31223,N_30744,N_30852);
xor U31224 (N_31224,N_30924,N_30881);
nand U31225 (N_31225,N_30636,N_30515);
and U31226 (N_31226,N_30577,N_30985);
nor U31227 (N_31227,N_30789,N_30640);
nor U31228 (N_31228,N_30661,N_30597);
nor U31229 (N_31229,N_30696,N_30818);
nand U31230 (N_31230,N_30540,N_30532);
and U31231 (N_31231,N_30979,N_30967);
nor U31232 (N_31232,N_30654,N_30616);
and U31233 (N_31233,N_30566,N_30595);
nor U31234 (N_31234,N_30603,N_30620);
or U31235 (N_31235,N_30890,N_30830);
xor U31236 (N_31236,N_30922,N_30734);
nor U31237 (N_31237,N_30604,N_30712);
or U31238 (N_31238,N_30894,N_30817);
nand U31239 (N_31239,N_30864,N_30991);
or U31240 (N_31240,N_30844,N_30697);
nand U31241 (N_31241,N_30809,N_30998);
nor U31242 (N_31242,N_30676,N_30882);
or U31243 (N_31243,N_30714,N_30594);
and U31244 (N_31244,N_30748,N_30615);
nand U31245 (N_31245,N_30652,N_30941);
and U31246 (N_31246,N_30883,N_30711);
or U31247 (N_31247,N_30627,N_30901);
and U31248 (N_31248,N_30514,N_30868);
nand U31249 (N_31249,N_30705,N_30997);
and U31250 (N_31250,N_30824,N_30888);
and U31251 (N_31251,N_30517,N_30657);
nand U31252 (N_31252,N_30684,N_30919);
nor U31253 (N_31253,N_30621,N_30569);
nor U31254 (N_31254,N_30601,N_30815);
nand U31255 (N_31255,N_30801,N_30989);
and U31256 (N_31256,N_30952,N_30806);
nand U31257 (N_31257,N_30906,N_30805);
or U31258 (N_31258,N_30710,N_30566);
or U31259 (N_31259,N_30737,N_30864);
nor U31260 (N_31260,N_30517,N_30530);
nor U31261 (N_31261,N_30529,N_30921);
or U31262 (N_31262,N_30660,N_30644);
and U31263 (N_31263,N_30821,N_30823);
nand U31264 (N_31264,N_30975,N_30518);
and U31265 (N_31265,N_30796,N_30804);
or U31266 (N_31266,N_30724,N_30568);
and U31267 (N_31267,N_30857,N_30995);
nand U31268 (N_31268,N_30600,N_30727);
xor U31269 (N_31269,N_30795,N_30760);
or U31270 (N_31270,N_30601,N_30759);
nand U31271 (N_31271,N_30734,N_30771);
nor U31272 (N_31272,N_30713,N_30536);
xor U31273 (N_31273,N_30576,N_30693);
and U31274 (N_31274,N_30743,N_30572);
nand U31275 (N_31275,N_30822,N_30716);
nand U31276 (N_31276,N_30745,N_30676);
nor U31277 (N_31277,N_30738,N_30736);
nand U31278 (N_31278,N_30878,N_30783);
xnor U31279 (N_31279,N_30791,N_30529);
xnor U31280 (N_31280,N_30536,N_30725);
and U31281 (N_31281,N_30643,N_30817);
and U31282 (N_31282,N_30723,N_30908);
and U31283 (N_31283,N_30505,N_30927);
nand U31284 (N_31284,N_30994,N_30896);
or U31285 (N_31285,N_30999,N_30874);
nand U31286 (N_31286,N_30530,N_30888);
nand U31287 (N_31287,N_30887,N_30575);
and U31288 (N_31288,N_30900,N_30707);
and U31289 (N_31289,N_30686,N_30861);
and U31290 (N_31290,N_30568,N_30833);
and U31291 (N_31291,N_30753,N_30679);
nand U31292 (N_31292,N_30676,N_30636);
nand U31293 (N_31293,N_30525,N_30998);
or U31294 (N_31294,N_30803,N_30584);
or U31295 (N_31295,N_30993,N_30868);
nand U31296 (N_31296,N_30604,N_30793);
nor U31297 (N_31297,N_30674,N_30918);
and U31298 (N_31298,N_30695,N_30548);
xnor U31299 (N_31299,N_30704,N_30949);
and U31300 (N_31300,N_30605,N_30688);
or U31301 (N_31301,N_30698,N_30601);
nand U31302 (N_31302,N_30617,N_30666);
nor U31303 (N_31303,N_30700,N_30867);
or U31304 (N_31304,N_30638,N_30773);
or U31305 (N_31305,N_30638,N_30765);
nor U31306 (N_31306,N_30931,N_30649);
or U31307 (N_31307,N_30541,N_30605);
or U31308 (N_31308,N_30675,N_30572);
nor U31309 (N_31309,N_30517,N_30567);
xor U31310 (N_31310,N_30969,N_30554);
and U31311 (N_31311,N_30527,N_30579);
and U31312 (N_31312,N_30972,N_30977);
xnor U31313 (N_31313,N_30812,N_30676);
or U31314 (N_31314,N_30907,N_30647);
nor U31315 (N_31315,N_30942,N_30752);
nor U31316 (N_31316,N_30865,N_30796);
nand U31317 (N_31317,N_30622,N_30975);
xor U31318 (N_31318,N_30672,N_30934);
and U31319 (N_31319,N_30771,N_30567);
and U31320 (N_31320,N_30561,N_30673);
nor U31321 (N_31321,N_30951,N_30514);
or U31322 (N_31322,N_30896,N_30557);
or U31323 (N_31323,N_30791,N_30555);
nand U31324 (N_31324,N_30635,N_30731);
xor U31325 (N_31325,N_30903,N_30814);
and U31326 (N_31326,N_30836,N_30692);
xnor U31327 (N_31327,N_30775,N_30654);
or U31328 (N_31328,N_30656,N_30835);
or U31329 (N_31329,N_30754,N_30590);
nand U31330 (N_31330,N_30944,N_30731);
nor U31331 (N_31331,N_30956,N_30878);
xor U31332 (N_31332,N_30732,N_30620);
nor U31333 (N_31333,N_30904,N_30569);
or U31334 (N_31334,N_30956,N_30757);
nor U31335 (N_31335,N_30951,N_30839);
and U31336 (N_31336,N_30598,N_30636);
nor U31337 (N_31337,N_30570,N_30514);
xnor U31338 (N_31338,N_30947,N_30703);
xor U31339 (N_31339,N_30585,N_30724);
or U31340 (N_31340,N_30625,N_30717);
nand U31341 (N_31341,N_30841,N_30871);
nand U31342 (N_31342,N_30671,N_30589);
nor U31343 (N_31343,N_30716,N_30586);
nand U31344 (N_31344,N_30664,N_30854);
and U31345 (N_31345,N_30919,N_30866);
nor U31346 (N_31346,N_30830,N_30823);
or U31347 (N_31347,N_30635,N_30528);
nor U31348 (N_31348,N_30667,N_30830);
nor U31349 (N_31349,N_30886,N_30522);
nand U31350 (N_31350,N_30784,N_30993);
nand U31351 (N_31351,N_30976,N_30651);
nor U31352 (N_31352,N_30873,N_30826);
nand U31353 (N_31353,N_30515,N_30840);
nor U31354 (N_31354,N_30854,N_30833);
nand U31355 (N_31355,N_30868,N_30509);
nor U31356 (N_31356,N_30534,N_30788);
and U31357 (N_31357,N_30688,N_30518);
nor U31358 (N_31358,N_30723,N_30978);
or U31359 (N_31359,N_30818,N_30985);
nor U31360 (N_31360,N_30815,N_30557);
or U31361 (N_31361,N_30528,N_30840);
and U31362 (N_31362,N_30522,N_30865);
nand U31363 (N_31363,N_30567,N_30664);
or U31364 (N_31364,N_30865,N_30694);
and U31365 (N_31365,N_30937,N_30729);
or U31366 (N_31366,N_30679,N_30520);
xnor U31367 (N_31367,N_30895,N_30508);
nor U31368 (N_31368,N_30975,N_30909);
or U31369 (N_31369,N_30693,N_30810);
nand U31370 (N_31370,N_30846,N_30610);
or U31371 (N_31371,N_30840,N_30745);
and U31372 (N_31372,N_30533,N_30581);
nand U31373 (N_31373,N_30725,N_30637);
and U31374 (N_31374,N_30926,N_30872);
nor U31375 (N_31375,N_30651,N_30601);
and U31376 (N_31376,N_30871,N_30606);
or U31377 (N_31377,N_30867,N_30771);
or U31378 (N_31378,N_30994,N_30998);
and U31379 (N_31379,N_30825,N_30792);
or U31380 (N_31380,N_30684,N_30839);
or U31381 (N_31381,N_30628,N_30980);
nor U31382 (N_31382,N_30811,N_30653);
and U31383 (N_31383,N_30521,N_30620);
or U31384 (N_31384,N_30797,N_30821);
and U31385 (N_31385,N_30786,N_30913);
or U31386 (N_31386,N_30665,N_30877);
or U31387 (N_31387,N_30590,N_30846);
or U31388 (N_31388,N_30568,N_30922);
nand U31389 (N_31389,N_30857,N_30504);
nand U31390 (N_31390,N_30656,N_30948);
or U31391 (N_31391,N_30636,N_30684);
or U31392 (N_31392,N_30677,N_30544);
and U31393 (N_31393,N_30545,N_30782);
or U31394 (N_31394,N_30712,N_30621);
and U31395 (N_31395,N_30613,N_30702);
and U31396 (N_31396,N_30715,N_30975);
nand U31397 (N_31397,N_30791,N_30708);
and U31398 (N_31398,N_30789,N_30783);
nor U31399 (N_31399,N_30563,N_30995);
or U31400 (N_31400,N_30667,N_30784);
nor U31401 (N_31401,N_30614,N_30864);
nor U31402 (N_31402,N_30531,N_30541);
nand U31403 (N_31403,N_30722,N_30862);
and U31404 (N_31404,N_30738,N_30825);
nor U31405 (N_31405,N_30686,N_30866);
nor U31406 (N_31406,N_30996,N_30760);
or U31407 (N_31407,N_30633,N_30565);
or U31408 (N_31408,N_30914,N_30762);
xor U31409 (N_31409,N_30868,N_30690);
or U31410 (N_31410,N_30793,N_30774);
nand U31411 (N_31411,N_30767,N_30816);
nor U31412 (N_31412,N_30582,N_30826);
nor U31413 (N_31413,N_30538,N_30733);
nand U31414 (N_31414,N_30660,N_30664);
nand U31415 (N_31415,N_30589,N_30651);
nand U31416 (N_31416,N_30519,N_30710);
xor U31417 (N_31417,N_30674,N_30934);
nor U31418 (N_31418,N_30671,N_30943);
nand U31419 (N_31419,N_30616,N_30594);
or U31420 (N_31420,N_30838,N_30936);
nor U31421 (N_31421,N_30732,N_30981);
nand U31422 (N_31422,N_30705,N_30994);
or U31423 (N_31423,N_30773,N_30729);
or U31424 (N_31424,N_30681,N_30580);
nand U31425 (N_31425,N_30784,N_30970);
nor U31426 (N_31426,N_30544,N_30855);
or U31427 (N_31427,N_30694,N_30656);
nor U31428 (N_31428,N_30781,N_30545);
nor U31429 (N_31429,N_30752,N_30671);
and U31430 (N_31430,N_30989,N_30537);
nand U31431 (N_31431,N_30744,N_30524);
nor U31432 (N_31432,N_30696,N_30911);
xor U31433 (N_31433,N_30781,N_30987);
nor U31434 (N_31434,N_30647,N_30716);
xor U31435 (N_31435,N_30998,N_30517);
nor U31436 (N_31436,N_30614,N_30930);
nand U31437 (N_31437,N_30771,N_30817);
nand U31438 (N_31438,N_30820,N_30645);
nand U31439 (N_31439,N_30624,N_30517);
and U31440 (N_31440,N_30798,N_30857);
nand U31441 (N_31441,N_30770,N_30635);
xnor U31442 (N_31442,N_30984,N_30592);
or U31443 (N_31443,N_30809,N_30815);
nand U31444 (N_31444,N_30866,N_30667);
xnor U31445 (N_31445,N_30860,N_30548);
or U31446 (N_31446,N_30667,N_30615);
and U31447 (N_31447,N_30886,N_30524);
nand U31448 (N_31448,N_30915,N_30949);
and U31449 (N_31449,N_30598,N_30945);
and U31450 (N_31450,N_30580,N_30714);
and U31451 (N_31451,N_30752,N_30850);
and U31452 (N_31452,N_30904,N_30667);
nor U31453 (N_31453,N_30597,N_30626);
and U31454 (N_31454,N_30960,N_30651);
nor U31455 (N_31455,N_30971,N_30935);
or U31456 (N_31456,N_30985,N_30708);
nand U31457 (N_31457,N_30625,N_30735);
nand U31458 (N_31458,N_30562,N_30988);
or U31459 (N_31459,N_30508,N_30837);
nor U31460 (N_31460,N_30914,N_30546);
nand U31461 (N_31461,N_30629,N_30878);
and U31462 (N_31462,N_30788,N_30674);
or U31463 (N_31463,N_30871,N_30705);
nor U31464 (N_31464,N_30619,N_30899);
or U31465 (N_31465,N_30912,N_30963);
and U31466 (N_31466,N_30569,N_30991);
and U31467 (N_31467,N_30846,N_30807);
xor U31468 (N_31468,N_30949,N_30636);
or U31469 (N_31469,N_30843,N_30511);
xor U31470 (N_31470,N_30980,N_30746);
nand U31471 (N_31471,N_30660,N_30603);
or U31472 (N_31472,N_30889,N_30928);
nor U31473 (N_31473,N_30658,N_30629);
and U31474 (N_31474,N_30778,N_30592);
or U31475 (N_31475,N_30661,N_30556);
nand U31476 (N_31476,N_30945,N_30697);
nand U31477 (N_31477,N_30604,N_30555);
and U31478 (N_31478,N_30790,N_30501);
nand U31479 (N_31479,N_30706,N_30850);
xnor U31480 (N_31480,N_30906,N_30984);
nor U31481 (N_31481,N_30844,N_30698);
or U31482 (N_31482,N_30772,N_30760);
nor U31483 (N_31483,N_30774,N_30590);
xor U31484 (N_31484,N_30998,N_30613);
or U31485 (N_31485,N_30566,N_30525);
or U31486 (N_31486,N_30974,N_30506);
xor U31487 (N_31487,N_30923,N_30869);
nor U31488 (N_31488,N_30832,N_30778);
or U31489 (N_31489,N_30582,N_30848);
and U31490 (N_31490,N_30997,N_30514);
nand U31491 (N_31491,N_30826,N_30651);
or U31492 (N_31492,N_30878,N_30727);
or U31493 (N_31493,N_30532,N_30802);
and U31494 (N_31494,N_30859,N_30770);
nand U31495 (N_31495,N_30628,N_30834);
xnor U31496 (N_31496,N_30729,N_30855);
nor U31497 (N_31497,N_30748,N_30625);
and U31498 (N_31498,N_30997,N_30547);
and U31499 (N_31499,N_30980,N_30948);
nand U31500 (N_31500,N_31413,N_31168);
nand U31501 (N_31501,N_31482,N_31111);
nor U31502 (N_31502,N_31348,N_31495);
and U31503 (N_31503,N_31016,N_31308);
and U31504 (N_31504,N_31396,N_31044);
or U31505 (N_31505,N_31331,N_31174);
or U31506 (N_31506,N_31198,N_31231);
nand U31507 (N_31507,N_31234,N_31257);
or U31508 (N_31508,N_31136,N_31059);
or U31509 (N_31509,N_31210,N_31486);
and U31510 (N_31510,N_31477,N_31155);
nor U31511 (N_31511,N_31449,N_31065);
xnor U31512 (N_31512,N_31214,N_31432);
or U31513 (N_31513,N_31106,N_31200);
nand U31514 (N_31514,N_31406,N_31349);
nor U31515 (N_31515,N_31218,N_31304);
nand U31516 (N_31516,N_31430,N_31368);
nand U31517 (N_31517,N_31407,N_31139);
nor U31518 (N_31518,N_31404,N_31239);
and U31519 (N_31519,N_31305,N_31343);
and U31520 (N_31520,N_31110,N_31202);
nand U31521 (N_31521,N_31251,N_31058);
nand U31522 (N_31522,N_31116,N_31276);
or U31523 (N_31523,N_31060,N_31385);
or U31524 (N_31524,N_31439,N_31123);
nand U31525 (N_31525,N_31473,N_31340);
nor U31526 (N_31526,N_31100,N_31487);
xor U31527 (N_31527,N_31144,N_31209);
nand U31528 (N_31528,N_31480,N_31279);
xor U31529 (N_31529,N_31208,N_31127);
xnor U31530 (N_31530,N_31086,N_31325);
or U31531 (N_31531,N_31120,N_31441);
or U31532 (N_31532,N_31133,N_31095);
or U31533 (N_31533,N_31048,N_31266);
nor U31534 (N_31534,N_31498,N_31020);
or U31535 (N_31535,N_31091,N_31244);
or U31536 (N_31536,N_31103,N_31367);
nand U31537 (N_31537,N_31177,N_31280);
and U31538 (N_31538,N_31314,N_31289);
nor U31539 (N_31539,N_31435,N_31221);
and U31540 (N_31540,N_31466,N_31328);
and U31541 (N_31541,N_31295,N_31452);
nor U31542 (N_31542,N_31063,N_31363);
nand U31543 (N_31543,N_31274,N_31445);
and U31544 (N_31544,N_31339,N_31252);
or U31545 (N_31545,N_31131,N_31219);
nand U31546 (N_31546,N_31410,N_31113);
and U31547 (N_31547,N_31423,N_31137);
xor U31548 (N_31548,N_31094,N_31447);
nor U31549 (N_31549,N_31357,N_31153);
nor U31550 (N_31550,N_31281,N_31062);
and U31551 (N_31551,N_31278,N_31260);
nor U31552 (N_31552,N_31199,N_31000);
nor U31553 (N_31553,N_31135,N_31076);
and U31554 (N_31554,N_31027,N_31483);
nand U31555 (N_31555,N_31286,N_31351);
nor U31556 (N_31556,N_31415,N_31246);
and U31557 (N_31557,N_31190,N_31356);
nand U31558 (N_31558,N_31457,N_31322);
or U31559 (N_31559,N_31227,N_31247);
nor U31560 (N_31560,N_31292,N_31241);
or U31561 (N_31561,N_31284,N_31017);
or U31562 (N_31562,N_31419,N_31165);
and U31563 (N_31563,N_31022,N_31262);
nor U31564 (N_31564,N_31023,N_31372);
nand U31565 (N_31565,N_31118,N_31312);
nand U31566 (N_31566,N_31005,N_31185);
and U31567 (N_31567,N_31364,N_31474);
nor U31568 (N_31568,N_31162,N_31342);
nor U31569 (N_31569,N_31374,N_31034);
or U31570 (N_31570,N_31269,N_31053);
or U31571 (N_31571,N_31186,N_31398);
nor U31572 (N_31572,N_31159,N_31150);
and U31573 (N_31573,N_31256,N_31238);
nand U31574 (N_31574,N_31187,N_31327);
nor U31575 (N_31575,N_31476,N_31080);
nor U31576 (N_31576,N_31164,N_31326);
or U31577 (N_31577,N_31294,N_31300);
or U31578 (N_31578,N_31307,N_31104);
and U31579 (N_31579,N_31365,N_31132);
nand U31580 (N_31580,N_31037,N_31147);
or U31581 (N_31581,N_31283,N_31298);
and U31582 (N_31582,N_31124,N_31157);
and U31583 (N_31583,N_31296,N_31389);
xor U31584 (N_31584,N_31097,N_31018);
nand U31585 (N_31585,N_31277,N_31098);
and U31586 (N_31586,N_31196,N_31206);
and U31587 (N_31587,N_31032,N_31010);
nand U31588 (N_31588,N_31195,N_31318);
or U31589 (N_31589,N_31149,N_31068);
and U31590 (N_31590,N_31382,N_31213);
or U31591 (N_31591,N_31056,N_31122);
nor U31592 (N_31592,N_31377,N_31460);
or U31593 (N_31593,N_31184,N_31216);
nor U31594 (N_31594,N_31454,N_31496);
xnor U31595 (N_31595,N_31288,N_31161);
xor U31596 (N_31596,N_31145,N_31141);
or U31597 (N_31597,N_31003,N_31041);
and U31598 (N_31598,N_31259,N_31101);
nor U31599 (N_31599,N_31222,N_31030);
nand U31600 (N_31600,N_31061,N_31067);
nand U31601 (N_31601,N_31417,N_31489);
xor U31602 (N_31602,N_31464,N_31261);
and U31603 (N_31603,N_31493,N_31180);
or U31604 (N_31604,N_31049,N_31455);
nand U31605 (N_31605,N_31172,N_31393);
nor U31606 (N_31606,N_31315,N_31412);
nand U31607 (N_31607,N_31258,N_31178);
or U31608 (N_31608,N_31448,N_31009);
nand U31609 (N_31609,N_31171,N_31337);
xnor U31610 (N_31610,N_31004,N_31057);
nand U31611 (N_31611,N_31485,N_31170);
nand U31612 (N_31612,N_31007,N_31084);
nand U31613 (N_31613,N_31429,N_31310);
nor U31614 (N_31614,N_31181,N_31399);
nand U31615 (N_31615,N_31243,N_31384);
or U31616 (N_31616,N_31176,N_31070);
or U31617 (N_31617,N_31245,N_31418);
or U31618 (N_31618,N_31203,N_31047);
and U31619 (N_31619,N_31054,N_31105);
and U31620 (N_31620,N_31484,N_31442);
nor U31621 (N_31621,N_31275,N_31248);
nand U31622 (N_31622,N_31375,N_31237);
xnor U31623 (N_31623,N_31211,N_31428);
nand U31624 (N_31624,N_31425,N_31414);
or U31625 (N_31625,N_31033,N_31468);
nor U31626 (N_31626,N_31263,N_31072);
and U31627 (N_31627,N_31008,N_31424);
nor U31628 (N_31628,N_31205,N_31040);
and U31629 (N_31629,N_31463,N_31319);
nand U31630 (N_31630,N_31042,N_31458);
xnor U31631 (N_31631,N_31142,N_31360);
or U31632 (N_31632,N_31163,N_31117);
or U31633 (N_31633,N_31055,N_31401);
and U31634 (N_31634,N_31250,N_31012);
xnor U31635 (N_31635,N_31287,N_31015);
and U31636 (N_31636,N_31311,N_31402);
and U31637 (N_31637,N_31450,N_31183);
and U31638 (N_31638,N_31108,N_31240);
xor U31639 (N_31639,N_31353,N_31193);
and U31640 (N_31640,N_31082,N_31126);
xnor U31641 (N_31641,N_31273,N_31488);
or U31642 (N_31642,N_31066,N_31235);
xor U31643 (N_31643,N_31217,N_31052);
nor U31644 (N_31644,N_31189,N_31045);
nand U31645 (N_31645,N_31138,N_31443);
xnor U31646 (N_31646,N_31151,N_31090);
and U31647 (N_31647,N_31359,N_31242);
or U31648 (N_31648,N_31395,N_31471);
and U31649 (N_31649,N_31341,N_31229);
nor U31650 (N_31650,N_31352,N_31011);
nor U31651 (N_31651,N_31285,N_31387);
nand U31652 (N_31652,N_31249,N_31381);
and U31653 (N_31653,N_31083,N_31469);
or U31654 (N_31654,N_31306,N_31014);
nand U31655 (N_31655,N_31021,N_31461);
or U31656 (N_31656,N_31336,N_31254);
or U31657 (N_31657,N_31265,N_31369);
nor U31658 (N_31658,N_31370,N_31267);
nor U31659 (N_31659,N_31081,N_31099);
and U31660 (N_31660,N_31107,N_31119);
and U31661 (N_31661,N_31400,N_31029);
and U31662 (N_31662,N_31475,N_31437);
nand U31663 (N_31663,N_31102,N_31109);
nand U31664 (N_31664,N_31050,N_31332);
nor U31665 (N_31665,N_31478,N_31143);
nor U31666 (N_31666,N_31397,N_31226);
or U31667 (N_31667,N_31223,N_31167);
xor U31668 (N_31668,N_31074,N_31197);
and U31669 (N_31669,N_31433,N_31492);
and U31670 (N_31670,N_31264,N_31255);
nor U31671 (N_31671,N_31130,N_31301);
and U31672 (N_31672,N_31467,N_31272);
or U31673 (N_31673,N_31329,N_31236);
nand U31674 (N_31674,N_31313,N_31134);
nor U31675 (N_31675,N_31392,N_31494);
and U31676 (N_31676,N_31499,N_31253);
or U31677 (N_31677,N_31085,N_31391);
nor U31678 (N_31678,N_31324,N_31152);
or U31679 (N_31679,N_31019,N_31230);
nand U31680 (N_31680,N_31179,N_31465);
nand U31681 (N_31681,N_31051,N_31380);
and U31682 (N_31682,N_31358,N_31491);
or U31683 (N_31683,N_31320,N_31232);
nor U31684 (N_31684,N_31146,N_31470);
xnor U31685 (N_31685,N_31077,N_31379);
and U31686 (N_31686,N_31355,N_31173);
and U31687 (N_31687,N_31096,N_31166);
and U31688 (N_31688,N_31148,N_31490);
and U31689 (N_31689,N_31421,N_31212);
nor U31690 (N_31690,N_31079,N_31129);
nor U31691 (N_31691,N_31225,N_31362);
nand U31692 (N_31692,N_31479,N_31128);
and U31693 (N_31693,N_31125,N_31481);
and U31694 (N_31694,N_31290,N_31182);
or U31695 (N_31695,N_31409,N_31201);
or U31696 (N_31696,N_31440,N_31036);
and U31697 (N_31697,N_31291,N_31092);
or U31698 (N_31698,N_31175,N_31031);
or U31699 (N_31699,N_31446,N_31071);
xnor U31700 (N_31700,N_31158,N_31366);
nor U31701 (N_31701,N_31330,N_31140);
nor U31702 (N_31702,N_31188,N_31089);
nor U31703 (N_31703,N_31302,N_31388);
xnor U31704 (N_31704,N_31282,N_31233);
and U31705 (N_31705,N_31344,N_31075);
nand U31706 (N_31706,N_31347,N_31078);
and U31707 (N_31707,N_31431,N_31299);
xnor U31708 (N_31708,N_31025,N_31204);
nor U31709 (N_31709,N_31444,N_31228);
nor U31710 (N_31710,N_31069,N_31043);
nand U31711 (N_31711,N_31378,N_31038);
nand U31712 (N_31712,N_31001,N_31024);
nand U31713 (N_31713,N_31064,N_31191);
nand U31714 (N_31714,N_31346,N_31115);
nand U31715 (N_31715,N_31154,N_31028);
or U31716 (N_31716,N_31408,N_31093);
nand U31717 (N_31717,N_31039,N_31416);
nand U31718 (N_31718,N_31427,N_31386);
and U31719 (N_31719,N_31156,N_31321);
and U31720 (N_31720,N_31333,N_31121);
or U31721 (N_31721,N_31220,N_31422);
xnor U31722 (N_31722,N_31114,N_31317);
or U31723 (N_31723,N_31026,N_31192);
nand U31724 (N_31724,N_31373,N_31451);
or U31725 (N_31725,N_31472,N_31350);
nor U31726 (N_31726,N_31268,N_31293);
or U31727 (N_31727,N_31405,N_31160);
or U31728 (N_31728,N_31194,N_31371);
and U31729 (N_31729,N_31335,N_31394);
and U31730 (N_31730,N_31013,N_31169);
nor U31731 (N_31731,N_31215,N_31497);
nor U31732 (N_31732,N_31035,N_31224);
nor U31733 (N_31733,N_31453,N_31006);
nand U31734 (N_31734,N_31434,N_31361);
nand U31735 (N_31735,N_31426,N_31420);
xor U31736 (N_31736,N_31087,N_31270);
nand U31737 (N_31737,N_31390,N_31112);
or U31738 (N_31738,N_31459,N_31207);
or U31739 (N_31739,N_31303,N_31316);
or U31740 (N_31740,N_31345,N_31338);
and U31741 (N_31741,N_31046,N_31376);
or U31742 (N_31742,N_31403,N_31297);
or U31743 (N_31743,N_31438,N_31073);
and U31744 (N_31744,N_31088,N_31002);
nor U31745 (N_31745,N_31323,N_31383);
or U31746 (N_31746,N_31411,N_31462);
nand U31747 (N_31747,N_31456,N_31436);
xnor U31748 (N_31748,N_31271,N_31354);
nor U31749 (N_31749,N_31334,N_31309);
nor U31750 (N_31750,N_31227,N_31362);
nand U31751 (N_31751,N_31117,N_31441);
or U31752 (N_31752,N_31315,N_31080);
nand U31753 (N_31753,N_31428,N_31120);
xor U31754 (N_31754,N_31497,N_31024);
nand U31755 (N_31755,N_31303,N_31013);
nand U31756 (N_31756,N_31313,N_31363);
nand U31757 (N_31757,N_31397,N_31151);
and U31758 (N_31758,N_31101,N_31377);
xor U31759 (N_31759,N_31481,N_31160);
nand U31760 (N_31760,N_31494,N_31087);
nand U31761 (N_31761,N_31063,N_31313);
nand U31762 (N_31762,N_31050,N_31265);
or U31763 (N_31763,N_31338,N_31247);
nor U31764 (N_31764,N_31337,N_31057);
nand U31765 (N_31765,N_31050,N_31157);
and U31766 (N_31766,N_31118,N_31394);
nand U31767 (N_31767,N_31294,N_31068);
nor U31768 (N_31768,N_31364,N_31258);
nand U31769 (N_31769,N_31425,N_31491);
nand U31770 (N_31770,N_31220,N_31253);
nor U31771 (N_31771,N_31476,N_31274);
or U31772 (N_31772,N_31275,N_31415);
nor U31773 (N_31773,N_31325,N_31415);
nand U31774 (N_31774,N_31347,N_31369);
or U31775 (N_31775,N_31318,N_31230);
or U31776 (N_31776,N_31023,N_31440);
nor U31777 (N_31777,N_31424,N_31253);
and U31778 (N_31778,N_31048,N_31308);
xor U31779 (N_31779,N_31133,N_31415);
nand U31780 (N_31780,N_31045,N_31294);
nor U31781 (N_31781,N_31446,N_31390);
and U31782 (N_31782,N_31100,N_31286);
or U31783 (N_31783,N_31450,N_31266);
nor U31784 (N_31784,N_31381,N_31407);
or U31785 (N_31785,N_31368,N_31014);
xor U31786 (N_31786,N_31250,N_31280);
nor U31787 (N_31787,N_31081,N_31008);
nor U31788 (N_31788,N_31316,N_31042);
or U31789 (N_31789,N_31351,N_31100);
or U31790 (N_31790,N_31006,N_31227);
or U31791 (N_31791,N_31376,N_31357);
and U31792 (N_31792,N_31439,N_31299);
or U31793 (N_31793,N_31375,N_31494);
nor U31794 (N_31794,N_31280,N_31245);
nand U31795 (N_31795,N_31312,N_31320);
or U31796 (N_31796,N_31457,N_31356);
xor U31797 (N_31797,N_31067,N_31424);
and U31798 (N_31798,N_31056,N_31171);
and U31799 (N_31799,N_31113,N_31056);
nand U31800 (N_31800,N_31124,N_31159);
nand U31801 (N_31801,N_31358,N_31230);
nor U31802 (N_31802,N_31164,N_31363);
or U31803 (N_31803,N_31134,N_31467);
nor U31804 (N_31804,N_31476,N_31495);
or U31805 (N_31805,N_31083,N_31233);
and U31806 (N_31806,N_31336,N_31047);
nor U31807 (N_31807,N_31253,N_31111);
nand U31808 (N_31808,N_31107,N_31365);
and U31809 (N_31809,N_31397,N_31154);
nor U31810 (N_31810,N_31337,N_31061);
or U31811 (N_31811,N_31008,N_31220);
or U31812 (N_31812,N_31485,N_31220);
xor U31813 (N_31813,N_31283,N_31342);
and U31814 (N_31814,N_31323,N_31282);
and U31815 (N_31815,N_31011,N_31421);
nand U31816 (N_31816,N_31047,N_31270);
xnor U31817 (N_31817,N_31256,N_31411);
or U31818 (N_31818,N_31121,N_31082);
nor U31819 (N_31819,N_31113,N_31479);
xor U31820 (N_31820,N_31222,N_31190);
and U31821 (N_31821,N_31241,N_31301);
or U31822 (N_31822,N_31180,N_31031);
nor U31823 (N_31823,N_31160,N_31428);
nor U31824 (N_31824,N_31005,N_31253);
xor U31825 (N_31825,N_31012,N_31358);
nand U31826 (N_31826,N_31250,N_31482);
and U31827 (N_31827,N_31496,N_31233);
nand U31828 (N_31828,N_31486,N_31347);
or U31829 (N_31829,N_31310,N_31035);
or U31830 (N_31830,N_31336,N_31003);
nand U31831 (N_31831,N_31405,N_31211);
nand U31832 (N_31832,N_31070,N_31317);
nor U31833 (N_31833,N_31322,N_31117);
xnor U31834 (N_31834,N_31311,N_31396);
nand U31835 (N_31835,N_31366,N_31065);
and U31836 (N_31836,N_31296,N_31266);
or U31837 (N_31837,N_31492,N_31181);
nand U31838 (N_31838,N_31356,N_31309);
nand U31839 (N_31839,N_31055,N_31105);
nand U31840 (N_31840,N_31482,N_31478);
xor U31841 (N_31841,N_31242,N_31336);
nor U31842 (N_31842,N_31175,N_31003);
or U31843 (N_31843,N_31464,N_31222);
or U31844 (N_31844,N_31341,N_31056);
nand U31845 (N_31845,N_31180,N_31495);
and U31846 (N_31846,N_31423,N_31103);
or U31847 (N_31847,N_31239,N_31341);
nand U31848 (N_31848,N_31137,N_31473);
xor U31849 (N_31849,N_31147,N_31445);
xnor U31850 (N_31850,N_31406,N_31279);
or U31851 (N_31851,N_31326,N_31163);
and U31852 (N_31852,N_31477,N_31160);
nor U31853 (N_31853,N_31273,N_31239);
nor U31854 (N_31854,N_31444,N_31352);
and U31855 (N_31855,N_31173,N_31470);
nor U31856 (N_31856,N_31420,N_31051);
or U31857 (N_31857,N_31435,N_31144);
or U31858 (N_31858,N_31017,N_31205);
nand U31859 (N_31859,N_31078,N_31170);
and U31860 (N_31860,N_31310,N_31322);
or U31861 (N_31861,N_31125,N_31400);
and U31862 (N_31862,N_31087,N_31023);
or U31863 (N_31863,N_31143,N_31052);
nor U31864 (N_31864,N_31188,N_31475);
and U31865 (N_31865,N_31261,N_31036);
nor U31866 (N_31866,N_31309,N_31184);
nor U31867 (N_31867,N_31073,N_31127);
nor U31868 (N_31868,N_31197,N_31018);
nand U31869 (N_31869,N_31235,N_31239);
nand U31870 (N_31870,N_31018,N_31226);
nand U31871 (N_31871,N_31087,N_31400);
nand U31872 (N_31872,N_31260,N_31094);
nand U31873 (N_31873,N_31036,N_31299);
and U31874 (N_31874,N_31272,N_31393);
and U31875 (N_31875,N_31240,N_31292);
xor U31876 (N_31876,N_31059,N_31470);
nand U31877 (N_31877,N_31485,N_31172);
or U31878 (N_31878,N_31445,N_31418);
or U31879 (N_31879,N_31390,N_31036);
nand U31880 (N_31880,N_31129,N_31412);
or U31881 (N_31881,N_31165,N_31351);
or U31882 (N_31882,N_31033,N_31028);
or U31883 (N_31883,N_31279,N_31434);
and U31884 (N_31884,N_31371,N_31256);
nor U31885 (N_31885,N_31348,N_31277);
and U31886 (N_31886,N_31444,N_31389);
nor U31887 (N_31887,N_31049,N_31062);
or U31888 (N_31888,N_31075,N_31121);
xnor U31889 (N_31889,N_31390,N_31371);
nor U31890 (N_31890,N_31265,N_31366);
nor U31891 (N_31891,N_31111,N_31458);
nor U31892 (N_31892,N_31073,N_31265);
and U31893 (N_31893,N_31169,N_31282);
or U31894 (N_31894,N_31070,N_31084);
xnor U31895 (N_31895,N_31212,N_31343);
and U31896 (N_31896,N_31005,N_31358);
nor U31897 (N_31897,N_31417,N_31089);
or U31898 (N_31898,N_31470,N_31383);
and U31899 (N_31899,N_31158,N_31350);
nand U31900 (N_31900,N_31400,N_31477);
nor U31901 (N_31901,N_31011,N_31488);
and U31902 (N_31902,N_31334,N_31131);
nand U31903 (N_31903,N_31230,N_31048);
or U31904 (N_31904,N_31084,N_31303);
nand U31905 (N_31905,N_31179,N_31416);
nor U31906 (N_31906,N_31212,N_31498);
nor U31907 (N_31907,N_31127,N_31175);
or U31908 (N_31908,N_31077,N_31088);
xnor U31909 (N_31909,N_31137,N_31249);
nand U31910 (N_31910,N_31327,N_31064);
and U31911 (N_31911,N_31153,N_31228);
nand U31912 (N_31912,N_31103,N_31122);
or U31913 (N_31913,N_31339,N_31299);
and U31914 (N_31914,N_31205,N_31486);
nor U31915 (N_31915,N_31032,N_31290);
nand U31916 (N_31916,N_31224,N_31407);
or U31917 (N_31917,N_31129,N_31426);
or U31918 (N_31918,N_31318,N_31476);
or U31919 (N_31919,N_31475,N_31351);
nor U31920 (N_31920,N_31226,N_31363);
and U31921 (N_31921,N_31027,N_31129);
and U31922 (N_31922,N_31292,N_31130);
nor U31923 (N_31923,N_31180,N_31274);
or U31924 (N_31924,N_31346,N_31317);
and U31925 (N_31925,N_31410,N_31255);
nand U31926 (N_31926,N_31442,N_31062);
or U31927 (N_31927,N_31188,N_31028);
nor U31928 (N_31928,N_31406,N_31395);
nor U31929 (N_31929,N_31383,N_31292);
nor U31930 (N_31930,N_31152,N_31302);
or U31931 (N_31931,N_31097,N_31111);
xnor U31932 (N_31932,N_31377,N_31414);
nand U31933 (N_31933,N_31348,N_31384);
or U31934 (N_31934,N_31137,N_31389);
or U31935 (N_31935,N_31409,N_31040);
nand U31936 (N_31936,N_31377,N_31162);
and U31937 (N_31937,N_31391,N_31098);
nand U31938 (N_31938,N_31168,N_31176);
nor U31939 (N_31939,N_31263,N_31427);
and U31940 (N_31940,N_31086,N_31293);
and U31941 (N_31941,N_31160,N_31030);
and U31942 (N_31942,N_31112,N_31046);
and U31943 (N_31943,N_31198,N_31217);
nor U31944 (N_31944,N_31156,N_31074);
xnor U31945 (N_31945,N_31212,N_31458);
nand U31946 (N_31946,N_31458,N_31166);
nor U31947 (N_31947,N_31353,N_31258);
xor U31948 (N_31948,N_31401,N_31149);
or U31949 (N_31949,N_31119,N_31016);
nand U31950 (N_31950,N_31256,N_31143);
nor U31951 (N_31951,N_31228,N_31451);
nor U31952 (N_31952,N_31231,N_31354);
nor U31953 (N_31953,N_31406,N_31461);
nand U31954 (N_31954,N_31193,N_31352);
xnor U31955 (N_31955,N_31434,N_31368);
nand U31956 (N_31956,N_31087,N_31119);
and U31957 (N_31957,N_31261,N_31170);
and U31958 (N_31958,N_31340,N_31406);
nor U31959 (N_31959,N_31008,N_31411);
or U31960 (N_31960,N_31298,N_31226);
nor U31961 (N_31961,N_31058,N_31474);
nor U31962 (N_31962,N_31221,N_31047);
xnor U31963 (N_31963,N_31489,N_31187);
and U31964 (N_31964,N_31325,N_31305);
nor U31965 (N_31965,N_31290,N_31020);
nor U31966 (N_31966,N_31202,N_31161);
nor U31967 (N_31967,N_31054,N_31099);
nor U31968 (N_31968,N_31142,N_31068);
nand U31969 (N_31969,N_31059,N_31494);
nand U31970 (N_31970,N_31314,N_31270);
or U31971 (N_31971,N_31011,N_31411);
or U31972 (N_31972,N_31453,N_31282);
nand U31973 (N_31973,N_31396,N_31065);
or U31974 (N_31974,N_31389,N_31365);
and U31975 (N_31975,N_31013,N_31277);
nor U31976 (N_31976,N_31470,N_31234);
nand U31977 (N_31977,N_31096,N_31117);
nand U31978 (N_31978,N_31388,N_31030);
nor U31979 (N_31979,N_31232,N_31275);
or U31980 (N_31980,N_31165,N_31413);
nand U31981 (N_31981,N_31123,N_31113);
xor U31982 (N_31982,N_31347,N_31425);
xnor U31983 (N_31983,N_31349,N_31033);
or U31984 (N_31984,N_31246,N_31279);
nor U31985 (N_31985,N_31164,N_31398);
nand U31986 (N_31986,N_31484,N_31092);
nor U31987 (N_31987,N_31213,N_31133);
nor U31988 (N_31988,N_31477,N_31286);
and U31989 (N_31989,N_31389,N_31452);
and U31990 (N_31990,N_31080,N_31173);
nor U31991 (N_31991,N_31193,N_31432);
and U31992 (N_31992,N_31424,N_31115);
and U31993 (N_31993,N_31320,N_31394);
nand U31994 (N_31994,N_31443,N_31261);
nor U31995 (N_31995,N_31205,N_31302);
and U31996 (N_31996,N_31401,N_31464);
nand U31997 (N_31997,N_31335,N_31417);
xor U31998 (N_31998,N_31050,N_31141);
or U31999 (N_31999,N_31323,N_31189);
xor U32000 (N_32000,N_31787,N_31769);
nor U32001 (N_32001,N_31875,N_31685);
nand U32002 (N_32002,N_31957,N_31573);
nor U32003 (N_32003,N_31906,N_31966);
or U32004 (N_32004,N_31645,N_31507);
xnor U32005 (N_32005,N_31965,N_31979);
and U32006 (N_32006,N_31525,N_31680);
nor U32007 (N_32007,N_31803,N_31516);
nand U32008 (N_32008,N_31641,N_31701);
or U32009 (N_32009,N_31816,N_31929);
nand U32010 (N_32010,N_31721,N_31667);
nand U32011 (N_32011,N_31873,N_31559);
xnor U32012 (N_32012,N_31774,N_31713);
and U32013 (N_32013,N_31669,N_31886);
or U32014 (N_32014,N_31688,N_31682);
nand U32015 (N_32015,N_31830,N_31663);
nor U32016 (N_32016,N_31594,N_31659);
nor U32017 (N_32017,N_31959,N_31722);
and U32018 (N_32018,N_31916,N_31623);
and U32019 (N_32019,N_31547,N_31674);
and U32020 (N_32020,N_31628,N_31927);
xor U32021 (N_32021,N_31613,N_31924);
nor U32022 (N_32022,N_31677,N_31513);
nor U32023 (N_32023,N_31562,N_31897);
nand U32024 (N_32024,N_31726,N_31735);
or U32025 (N_32025,N_31901,N_31828);
xnor U32026 (N_32026,N_31502,N_31838);
xor U32027 (N_32027,N_31601,N_31619);
and U32028 (N_32028,N_31978,N_31988);
or U32029 (N_32029,N_31938,N_31676);
or U32030 (N_32030,N_31653,N_31611);
nor U32031 (N_32031,N_31687,N_31541);
nand U32032 (N_32032,N_31555,N_31603);
nand U32033 (N_32033,N_31753,N_31931);
or U32034 (N_32034,N_31574,N_31567);
and U32035 (N_32035,N_31770,N_31958);
or U32036 (N_32036,N_31968,N_31622);
nand U32037 (N_32037,N_31666,N_31987);
nand U32038 (N_32038,N_31941,N_31766);
nand U32039 (N_32039,N_31524,N_31584);
nor U32040 (N_32040,N_31575,N_31986);
nand U32041 (N_32041,N_31934,N_31727);
nor U32042 (N_32042,N_31718,N_31748);
or U32043 (N_32043,N_31790,N_31570);
or U32044 (N_32044,N_31734,N_31856);
nor U32045 (N_32045,N_31964,N_31837);
xor U32046 (N_32046,N_31702,N_31984);
and U32047 (N_32047,N_31944,N_31843);
nor U32048 (N_32048,N_31907,N_31913);
and U32049 (N_32049,N_31894,N_31665);
nor U32050 (N_32050,N_31861,N_31751);
nor U32051 (N_32051,N_31813,N_31733);
nand U32052 (N_32052,N_31605,N_31930);
or U32053 (N_32053,N_31689,N_31851);
or U32054 (N_32054,N_31536,N_31880);
nand U32055 (N_32055,N_31607,N_31834);
xnor U32056 (N_32056,N_31662,N_31954);
nor U32057 (N_32057,N_31951,N_31678);
or U32058 (N_32058,N_31824,N_31928);
nor U32059 (N_32059,N_31657,N_31848);
and U32060 (N_32060,N_31707,N_31962);
or U32061 (N_32061,N_31878,N_31889);
nor U32062 (N_32062,N_31757,N_31716);
nand U32063 (N_32063,N_31548,N_31719);
nand U32064 (N_32064,N_31528,N_31936);
nor U32065 (N_32065,N_31772,N_31963);
nor U32066 (N_32066,N_31630,N_31960);
or U32067 (N_32067,N_31569,N_31729);
or U32068 (N_32068,N_31893,N_31832);
xor U32069 (N_32069,N_31910,N_31629);
nor U32070 (N_32070,N_31699,N_31723);
nor U32071 (N_32071,N_31937,N_31802);
nand U32072 (N_32072,N_31637,N_31724);
and U32073 (N_32073,N_31614,N_31577);
or U32074 (N_32074,N_31595,N_31867);
nor U32075 (N_32075,N_31836,N_31887);
nor U32076 (N_32076,N_31847,N_31974);
or U32077 (N_32077,N_31994,N_31804);
nor U32078 (N_32078,N_31668,N_31796);
xnor U32079 (N_32079,N_31535,N_31534);
and U32080 (N_32080,N_31797,N_31952);
or U32081 (N_32081,N_31649,N_31658);
xor U32082 (N_32082,N_31743,N_31985);
nand U32083 (N_32083,N_31530,N_31865);
or U32084 (N_32084,N_31864,N_31806);
or U32085 (N_32085,N_31884,N_31531);
xor U32086 (N_32086,N_31932,N_31872);
and U32087 (N_32087,N_31800,N_31681);
or U32088 (N_32088,N_31869,N_31514);
or U32089 (N_32089,N_31749,N_31839);
and U32090 (N_32090,N_31909,N_31679);
and U32091 (N_32091,N_31717,N_31792);
xor U32092 (N_32092,N_31660,N_31620);
or U32093 (N_32093,N_31538,N_31550);
nor U32094 (N_32094,N_31709,N_31754);
and U32095 (N_32095,N_31639,N_31608);
and U32096 (N_32096,N_31644,N_31624);
nor U32097 (N_32097,N_31672,N_31744);
nor U32098 (N_32098,N_31921,N_31908);
and U32099 (N_32099,N_31715,N_31610);
and U32100 (N_32100,N_31755,N_31593);
and U32101 (N_32101,N_31915,N_31731);
and U32102 (N_32102,N_31829,N_31596);
nand U32103 (N_32103,N_31784,N_31788);
xor U32104 (N_32104,N_31549,N_31862);
nor U32105 (N_32105,N_31609,N_31691);
nand U32106 (N_32106,N_31583,N_31825);
or U32107 (N_32107,N_31551,N_31858);
and U32108 (N_32108,N_31747,N_31526);
nor U32109 (N_32109,N_31982,N_31693);
or U32110 (N_32110,N_31768,N_31565);
or U32111 (N_32111,N_31556,N_31798);
and U32112 (N_32112,N_31779,N_31617);
or U32113 (N_32113,N_31750,N_31956);
and U32114 (N_32114,N_31859,N_31640);
xor U32115 (N_32115,N_31521,N_31794);
and U32116 (N_32116,N_31590,N_31741);
or U32117 (N_32117,N_31914,N_31580);
or U32118 (N_32118,N_31592,N_31627);
and U32119 (N_32119,N_31566,N_31578);
nand U32120 (N_32120,N_31799,N_31997);
nand U32121 (N_32121,N_31523,N_31553);
or U32122 (N_32122,N_31650,N_31876);
nand U32123 (N_32123,N_31899,N_31903);
or U32124 (N_32124,N_31920,N_31683);
and U32125 (N_32125,N_31852,N_31849);
or U32126 (N_32126,N_31891,N_31585);
nand U32127 (N_32127,N_31781,N_31892);
or U32128 (N_32128,N_31615,N_31654);
xnor U32129 (N_32129,N_31883,N_31618);
or U32130 (N_32130,N_31673,N_31568);
or U32131 (N_32131,N_31517,N_31780);
nor U32132 (N_32132,N_31764,N_31571);
nand U32133 (N_32133,N_31992,N_31874);
nor U32134 (N_32134,N_31948,N_31826);
or U32135 (N_32135,N_31684,N_31821);
or U32136 (N_32136,N_31902,N_31708);
nor U32137 (N_32137,N_31651,N_31777);
nor U32138 (N_32138,N_31817,N_31519);
or U32139 (N_32139,N_31625,N_31977);
or U32140 (N_32140,N_31763,N_31833);
xor U32141 (N_32141,N_31969,N_31647);
xor U32142 (N_32142,N_31926,N_31540);
nor U32143 (N_32143,N_31587,N_31515);
or U32144 (N_32144,N_31612,N_31697);
or U32145 (N_32145,N_31560,N_31706);
and U32146 (N_32146,N_31890,N_31812);
and U32147 (N_32147,N_31818,N_31670);
nor U32148 (N_32148,N_31738,N_31632);
or U32149 (N_32149,N_31918,N_31631);
xnor U32150 (N_32150,N_31822,N_31840);
nor U32151 (N_32151,N_31881,N_31845);
or U32152 (N_32152,N_31767,N_31501);
and U32153 (N_32153,N_31616,N_31773);
nor U32154 (N_32154,N_31919,N_31989);
nor U32155 (N_32155,N_31819,N_31942);
and U32156 (N_32156,N_31537,N_31863);
or U32157 (N_32157,N_31815,N_31505);
and U32158 (N_32158,N_31811,N_31967);
or U32159 (N_32159,N_31529,N_31564);
xnor U32160 (N_32160,N_31879,N_31835);
and U32161 (N_32161,N_31973,N_31980);
nor U32162 (N_32162,N_31643,N_31945);
nor U32163 (N_32163,N_31563,N_31971);
or U32164 (N_32164,N_31546,N_31694);
nand U32165 (N_32165,N_31939,N_31572);
nand U32166 (N_32166,N_31905,N_31656);
nor U32167 (N_32167,N_31991,N_31506);
and U32168 (N_32168,N_31740,N_31807);
xnor U32169 (N_32169,N_31855,N_31972);
nor U32170 (N_32170,N_31761,N_31882);
nor U32171 (N_32171,N_31911,N_31725);
or U32172 (N_32172,N_31655,N_31844);
nor U32173 (N_32173,N_31898,N_31503);
and U32174 (N_32174,N_31935,N_31756);
nand U32175 (N_32175,N_31604,N_31542);
or U32176 (N_32176,N_31976,N_31805);
nand U32177 (N_32177,N_31652,N_31695);
or U32178 (N_32178,N_31664,N_31808);
nand U32179 (N_32179,N_31917,N_31850);
xor U32180 (N_32180,N_31510,N_31646);
and U32181 (N_32181,N_31539,N_31745);
nor U32182 (N_32182,N_31675,N_31504);
xor U32183 (N_32183,N_31760,N_31633);
nor U32184 (N_32184,N_31714,N_31728);
nand U32185 (N_32185,N_31842,N_31561);
nor U32186 (N_32186,N_31955,N_31775);
xnor U32187 (N_32187,N_31885,N_31661);
and U32188 (N_32188,N_31557,N_31933);
nor U32189 (N_32189,N_31552,N_31636);
and U32190 (N_32190,N_31710,N_31739);
or U32191 (N_32191,N_31500,N_31581);
nand U32192 (N_32192,N_31512,N_31854);
nand U32193 (N_32193,N_31999,N_31746);
and U32194 (N_32194,N_31696,N_31995);
and U32195 (N_32195,N_31544,N_31947);
xnor U32196 (N_32196,N_31801,N_31888);
nor U32197 (N_32197,N_31522,N_31904);
and U32198 (N_32198,N_31970,N_31518);
nand U32199 (N_32199,N_31690,N_31543);
and U32200 (N_32200,N_31634,N_31949);
or U32201 (N_32201,N_31759,N_31532);
and U32202 (N_32202,N_31900,N_31589);
and U32203 (N_32203,N_31732,N_31606);
nor U32204 (N_32204,N_31950,N_31635);
xnor U32205 (N_32205,N_31730,N_31712);
and U32206 (N_32206,N_31704,N_31698);
and U32207 (N_32207,N_31576,N_31602);
nor U32208 (N_32208,N_31692,N_31598);
nand U32209 (N_32209,N_31975,N_31827);
and U32210 (N_32210,N_31554,N_31791);
nand U32211 (N_32211,N_31940,N_31720);
or U32212 (N_32212,N_31686,N_31520);
or U32213 (N_32213,N_31993,N_31857);
nor U32214 (N_32214,N_31545,N_31765);
nor U32215 (N_32215,N_31591,N_31814);
xnor U32216 (N_32216,N_31786,N_31752);
and U32217 (N_32217,N_31923,N_31533);
and U32218 (N_32218,N_31793,N_31946);
xnor U32219 (N_32219,N_31912,N_31961);
nand U32220 (N_32220,N_31642,N_31711);
and U32221 (N_32221,N_31558,N_31866);
nand U32222 (N_32222,N_31925,N_31586);
nand U32223 (N_32223,N_31853,N_31626);
or U32224 (N_32224,N_31638,N_31621);
or U32225 (N_32225,N_31700,N_31758);
and U32226 (N_32226,N_31703,N_31998);
or U32227 (N_32227,N_31737,N_31782);
nor U32228 (N_32228,N_31810,N_31705);
or U32229 (N_32229,N_31509,N_31820);
nor U32230 (N_32230,N_31860,N_31846);
or U32231 (N_32231,N_31742,N_31841);
nor U32232 (N_32232,N_31795,N_31896);
and U32233 (N_32233,N_31895,N_31809);
xnor U32234 (N_32234,N_31671,N_31527);
nor U32235 (N_32235,N_31600,N_31943);
and U32236 (N_32236,N_31789,N_31736);
or U32237 (N_32237,N_31877,N_31783);
or U32238 (N_32238,N_31990,N_31823);
nor U32239 (N_32239,N_31868,N_31582);
nor U32240 (N_32240,N_31762,N_31996);
nor U32241 (N_32241,N_31778,N_31648);
nor U32242 (N_32242,N_31588,N_31511);
nand U32243 (N_32243,N_31953,N_31776);
xor U32244 (N_32244,N_31870,N_31508);
nor U32245 (N_32245,N_31831,N_31771);
nor U32246 (N_32246,N_31599,N_31983);
nor U32247 (N_32247,N_31981,N_31579);
nand U32248 (N_32248,N_31871,N_31785);
xor U32249 (N_32249,N_31597,N_31922);
nand U32250 (N_32250,N_31949,N_31740);
or U32251 (N_32251,N_31588,N_31635);
nor U32252 (N_32252,N_31780,N_31965);
and U32253 (N_32253,N_31604,N_31541);
xnor U32254 (N_32254,N_31672,N_31944);
xor U32255 (N_32255,N_31948,N_31972);
and U32256 (N_32256,N_31640,N_31585);
nor U32257 (N_32257,N_31717,N_31809);
nand U32258 (N_32258,N_31980,N_31851);
or U32259 (N_32259,N_31675,N_31689);
nor U32260 (N_32260,N_31709,N_31767);
and U32261 (N_32261,N_31752,N_31845);
nand U32262 (N_32262,N_31944,N_31947);
or U32263 (N_32263,N_31705,N_31770);
or U32264 (N_32264,N_31768,N_31889);
or U32265 (N_32265,N_31646,N_31876);
nor U32266 (N_32266,N_31922,N_31933);
nand U32267 (N_32267,N_31604,N_31513);
or U32268 (N_32268,N_31697,N_31559);
and U32269 (N_32269,N_31541,N_31961);
nand U32270 (N_32270,N_31650,N_31686);
nand U32271 (N_32271,N_31503,N_31861);
xnor U32272 (N_32272,N_31954,N_31673);
xor U32273 (N_32273,N_31931,N_31866);
nand U32274 (N_32274,N_31657,N_31645);
nor U32275 (N_32275,N_31609,N_31556);
or U32276 (N_32276,N_31756,N_31789);
and U32277 (N_32277,N_31596,N_31967);
xnor U32278 (N_32278,N_31807,N_31821);
nand U32279 (N_32279,N_31873,N_31775);
xor U32280 (N_32280,N_31834,N_31611);
xor U32281 (N_32281,N_31606,N_31773);
and U32282 (N_32282,N_31584,N_31933);
xnor U32283 (N_32283,N_31648,N_31656);
or U32284 (N_32284,N_31759,N_31659);
or U32285 (N_32285,N_31864,N_31813);
or U32286 (N_32286,N_31632,N_31857);
and U32287 (N_32287,N_31858,N_31594);
nor U32288 (N_32288,N_31902,N_31530);
nor U32289 (N_32289,N_31865,N_31637);
or U32290 (N_32290,N_31846,N_31895);
or U32291 (N_32291,N_31821,N_31970);
and U32292 (N_32292,N_31649,N_31850);
nand U32293 (N_32293,N_31683,N_31584);
nor U32294 (N_32294,N_31775,N_31514);
and U32295 (N_32295,N_31604,N_31849);
or U32296 (N_32296,N_31581,N_31926);
and U32297 (N_32297,N_31723,N_31659);
nor U32298 (N_32298,N_31685,N_31578);
or U32299 (N_32299,N_31619,N_31844);
nor U32300 (N_32300,N_31849,N_31848);
and U32301 (N_32301,N_31862,N_31595);
nor U32302 (N_32302,N_31832,N_31969);
and U32303 (N_32303,N_31574,N_31823);
nand U32304 (N_32304,N_31787,N_31916);
and U32305 (N_32305,N_31808,N_31500);
and U32306 (N_32306,N_31768,N_31927);
nor U32307 (N_32307,N_31508,N_31632);
nand U32308 (N_32308,N_31573,N_31767);
and U32309 (N_32309,N_31606,N_31695);
or U32310 (N_32310,N_31820,N_31885);
nand U32311 (N_32311,N_31570,N_31992);
nand U32312 (N_32312,N_31898,N_31676);
xor U32313 (N_32313,N_31589,N_31662);
nand U32314 (N_32314,N_31994,N_31584);
xor U32315 (N_32315,N_31538,N_31697);
nor U32316 (N_32316,N_31705,N_31550);
or U32317 (N_32317,N_31971,N_31773);
nor U32318 (N_32318,N_31857,N_31915);
nand U32319 (N_32319,N_31920,N_31735);
nor U32320 (N_32320,N_31826,N_31564);
nand U32321 (N_32321,N_31839,N_31986);
nor U32322 (N_32322,N_31718,N_31658);
xor U32323 (N_32323,N_31654,N_31799);
nor U32324 (N_32324,N_31822,N_31942);
nor U32325 (N_32325,N_31706,N_31767);
nor U32326 (N_32326,N_31663,N_31524);
and U32327 (N_32327,N_31854,N_31637);
and U32328 (N_32328,N_31621,N_31825);
and U32329 (N_32329,N_31982,N_31592);
and U32330 (N_32330,N_31612,N_31621);
or U32331 (N_32331,N_31559,N_31534);
nand U32332 (N_32332,N_31777,N_31574);
nand U32333 (N_32333,N_31706,N_31541);
xnor U32334 (N_32334,N_31541,N_31923);
nand U32335 (N_32335,N_31574,N_31975);
and U32336 (N_32336,N_31933,N_31893);
or U32337 (N_32337,N_31811,N_31919);
and U32338 (N_32338,N_31834,N_31907);
or U32339 (N_32339,N_31593,N_31861);
or U32340 (N_32340,N_31972,N_31903);
nor U32341 (N_32341,N_31554,N_31687);
nand U32342 (N_32342,N_31971,N_31927);
nand U32343 (N_32343,N_31807,N_31571);
nand U32344 (N_32344,N_31919,N_31592);
or U32345 (N_32345,N_31589,N_31958);
nand U32346 (N_32346,N_31891,N_31551);
nand U32347 (N_32347,N_31717,N_31574);
xnor U32348 (N_32348,N_31934,N_31530);
nor U32349 (N_32349,N_31563,N_31835);
and U32350 (N_32350,N_31963,N_31936);
or U32351 (N_32351,N_31651,N_31898);
nand U32352 (N_32352,N_31775,N_31749);
and U32353 (N_32353,N_31634,N_31957);
and U32354 (N_32354,N_31848,N_31979);
or U32355 (N_32355,N_31502,N_31985);
nand U32356 (N_32356,N_31922,N_31741);
and U32357 (N_32357,N_31886,N_31733);
nor U32358 (N_32358,N_31500,N_31961);
nand U32359 (N_32359,N_31888,N_31507);
and U32360 (N_32360,N_31542,N_31717);
nand U32361 (N_32361,N_31842,N_31521);
nand U32362 (N_32362,N_31614,N_31911);
or U32363 (N_32363,N_31845,N_31595);
nor U32364 (N_32364,N_31917,N_31828);
nor U32365 (N_32365,N_31937,N_31814);
nor U32366 (N_32366,N_31616,N_31948);
nor U32367 (N_32367,N_31568,N_31836);
nand U32368 (N_32368,N_31833,N_31661);
and U32369 (N_32369,N_31543,N_31571);
and U32370 (N_32370,N_31602,N_31774);
nor U32371 (N_32371,N_31970,N_31549);
nand U32372 (N_32372,N_31985,N_31585);
xor U32373 (N_32373,N_31742,N_31882);
and U32374 (N_32374,N_31543,N_31978);
nor U32375 (N_32375,N_31540,N_31534);
xnor U32376 (N_32376,N_31892,N_31661);
xor U32377 (N_32377,N_31510,N_31931);
nand U32378 (N_32378,N_31871,N_31969);
xnor U32379 (N_32379,N_31814,N_31628);
xor U32380 (N_32380,N_31897,N_31720);
or U32381 (N_32381,N_31733,N_31854);
xnor U32382 (N_32382,N_31672,N_31533);
and U32383 (N_32383,N_31660,N_31594);
nor U32384 (N_32384,N_31525,N_31931);
or U32385 (N_32385,N_31687,N_31998);
nor U32386 (N_32386,N_31619,N_31835);
or U32387 (N_32387,N_31695,N_31941);
or U32388 (N_32388,N_31871,N_31694);
and U32389 (N_32389,N_31705,N_31566);
or U32390 (N_32390,N_31534,N_31774);
and U32391 (N_32391,N_31625,N_31800);
nand U32392 (N_32392,N_31516,N_31924);
nand U32393 (N_32393,N_31916,N_31828);
nand U32394 (N_32394,N_31965,N_31901);
or U32395 (N_32395,N_31884,N_31872);
nand U32396 (N_32396,N_31924,N_31511);
or U32397 (N_32397,N_31986,N_31665);
or U32398 (N_32398,N_31849,N_31828);
and U32399 (N_32399,N_31857,N_31652);
nand U32400 (N_32400,N_31860,N_31523);
xnor U32401 (N_32401,N_31516,N_31972);
or U32402 (N_32402,N_31626,N_31683);
and U32403 (N_32403,N_31643,N_31533);
or U32404 (N_32404,N_31718,N_31678);
or U32405 (N_32405,N_31822,N_31657);
nor U32406 (N_32406,N_31895,N_31743);
and U32407 (N_32407,N_31681,N_31577);
nand U32408 (N_32408,N_31560,N_31911);
nand U32409 (N_32409,N_31909,N_31636);
and U32410 (N_32410,N_31637,N_31648);
nor U32411 (N_32411,N_31596,N_31723);
and U32412 (N_32412,N_31740,N_31698);
nand U32413 (N_32413,N_31824,N_31822);
xor U32414 (N_32414,N_31617,N_31527);
nor U32415 (N_32415,N_31878,N_31524);
nor U32416 (N_32416,N_31701,N_31892);
and U32417 (N_32417,N_31685,N_31551);
nand U32418 (N_32418,N_31508,N_31959);
or U32419 (N_32419,N_31717,N_31679);
and U32420 (N_32420,N_31572,N_31886);
nor U32421 (N_32421,N_31987,N_31583);
or U32422 (N_32422,N_31512,N_31905);
or U32423 (N_32423,N_31840,N_31670);
or U32424 (N_32424,N_31640,N_31508);
nand U32425 (N_32425,N_31864,N_31611);
and U32426 (N_32426,N_31815,N_31963);
nand U32427 (N_32427,N_31861,N_31799);
nand U32428 (N_32428,N_31730,N_31699);
nor U32429 (N_32429,N_31836,N_31739);
or U32430 (N_32430,N_31685,N_31580);
nand U32431 (N_32431,N_31788,N_31647);
nor U32432 (N_32432,N_31645,N_31698);
nand U32433 (N_32433,N_31888,N_31979);
and U32434 (N_32434,N_31786,N_31956);
nor U32435 (N_32435,N_31838,N_31575);
and U32436 (N_32436,N_31953,N_31684);
xnor U32437 (N_32437,N_31650,N_31853);
or U32438 (N_32438,N_31943,N_31553);
nor U32439 (N_32439,N_31919,N_31796);
and U32440 (N_32440,N_31739,N_31975);
or U32441 (N_32441,N_31679,N_31546);
and U32442 (N_32442,N_31520,N_31708);
nor U32443 (N_32443,N_31776,N_31650);
nand U32444 (N_32444,N_31787,N_31645);
nand U32445 (N_32445,N_31957,N_31695);
nor U32446 (N_32446,N_31810,N_31697);
or U32447 (N_32447,N_31511,N_31731);
nor U32448 (N_32448,N_31671,N_31619);
nand U32449 (N_32449,N_31553,N_31767);
nand U32450 (N_32450,N_31637,N_31954);
nor U32451 (N_32451,N_31607,N_31913);
nand U32452 (N_32452,N_31667,N_31803);
nor U32453 (N_32453,N_31519,N_31544);
and U32454 (N_32454,N_31941,N_31596);
nand U32455 (N_32455,N_31989,N_31915);
and U32456 (N_32456,N_31705,N_31639);
xnor U32457 (N_32457,N_31601,N_31881);
nor U32458 (N_32458,N_31794,N_31987);
nor U32459 (N_32459,N_31959,N_31771);
nor U32460 (N_32460,N_31820,N_31999);
or U32461 (N_32461,N_31601,N_31597);
nor U32462 (N_32462,N_31898,N_31912);
and U32463 (N_32463,N_31884,N_31926);
nand U32464 (N_32464,N_31741,N_31657);
and U32465 (N_32465,N_31951,N_31747);
and U32466 (N_32466,N_31759,N_31789);
xor U32467 (N_32467,N_31665,N_31758);
nor U32468 (N_32468,N_31644,N_31979);
nor U32469 (N_32469,N_31505,N_31676);
or U32470 (N_32470,N_31511,N_31894);
and U32471 (N_32471,N_31738,N_31946);
nor U32472 (N_32472,N_31807,N_31914);
xnor U32473 (N_32473,N_31706,N_31726);
or U32474 (N_32474,N_31857,N_31663);
xnor U32475 (N_32475,N_31918,N_31910);
xor U32476 (N_32476,N_31870,N_31540);
or U32477 (N_32477,N_31662,N_31808);
and U32478 (N_32478,N_31804,N_31978);
or U32479 (N_32479,N_31580,N_31766);
nand U32480 (N_32480,N_31953,N_31777);
nand U32481 (N_32481,N_31833,N_31556);
and U32482 (N_32482,N_31616,N_31508);
nor U32483 (N_32483,N_31642,N_31983);
nand U32484 (N_32484,N_31712,N_31998);
nand U32485 (N_32485,N_31799,N_31883);
nor U32486 (N_32486,N_31993,N_31876);
or U32487 (N_32487,N_31976,N_31885);
and U32488 (N_32488,N_31656,N_31592);
and U32489 (N_32489,N_31716,N_31778);
nor U32490 (N_32490,N_31862,N_31574);
nor U32491 (N_32491,N_31788,N_31927);
nand U32492 (N_32492,N_31502,N_31705);
nor U32493 (N_32493,N_31993,N_31852);
or U32494 (N_32494,N_31978,N_31513);
nand U32495 (N_32495,N_31771,N_31961);
and U32496 (N_32496,N_31548,N_31948);
nor U32497 (N_32497,N_31890,N_31840);
or U32498 (N_32498,N_31830,N_31897);
nand U32499 (N_32499,N_31879,N_31832);
or U32500 (N_32500,N_32401,N_32074);
and U32501 (N_32501,N_32333,N_32043);
xnor U32502 (N_32502,N_32453,N_32263);
and U32503 (N_32503,N_32146,N_32148);
nand U32504 (N_32504,N_32203,N_32116);
and U32505 (N_32505,N_32448,N_32212);
and U32506 (N_32506,N_32032,N_32051);
nor U32507 (N_32507,N_32187,N_32122);
or U32508 (N_32508,N_32101,N_32443);
nor U32509 (N_32509,N_32308,N_32123);
nor U32510 (N_32510,N_32049,N_32325);
nor U32511 (N_32511,N_32319,N_32292);
nand U32512 (N_32512,N_32246,N_32073);
nand U32513 (N_32513,N_32423,N_32429);
nor U32514 (N_32514,N_32035,N_32458);
nand U32515 (N_32515,N_32283,N_32001);
nor U32516 (N_32516,N_32222,N_32274);
and U32517 (N_32517,N_32268,N_32430);
or U32518 (N_32518,N_32113,N_32277);
nor U32519 (N_32519,N_32321,N_32295);
nor U32520 (N_32520,N_32008,N_32027);
xor U32521 (N_32521,N_32312,N_32299);
or U32522 (N_32522,N_32219,N_32172);
or U32523 (N_32523,N_32488,N_32346);
or U32524 (N_32524,N_32270,N_32403);
and U32525 (N_32525,N_32190,N_32002);
and U32526 (N_32526,N_32075,N_32197);
and U32527 (N_32527,N_32249,N_32230);
nor U32528 (N_32528,N_32064,N_32413);
nand U32529 (N_32529,N_32210,N_32260);
nor U32530 (N_32530,N_32377,N_32454);
nand U32531 (N_32531,N_32490,N_32486);
or U32532 (N_32532,N_32004,N_32478);
xor U32533 (N_32533,N_32300,N_32067);
nand U32534 (N_32534,N_32056,N_32119);
xnor U32535 (N_32535,N_32361,N_32176);
or U32536 (N_32536,N_32223,N_32129);
or U32537 (N_32537,N_32435,N_32449);
and U32538 (N_32538,N_32163,N_32297);
and U32539 (N_32539,N_32467,N_32406);
nor U32540 (N_32540,N_32144,N_32010);
and U32541 (N_32541,N_32434,N_32477);
and U32542 (N_32542,N_32348,N_32293);
or U32543 (N_32543,N_32284,N_32093);
nand U32544 (N_32544,N_32217,N_32017);
nor U32545 (N_32545,N_32438,N_32427);
nor U32546 (N_32546,N_32152,N_32385);
or U32547 (N_32547,N_32095,N_32294);
or U32548 (N_32548,N_32341,N_32173);
or U32549 (N_32549,N_32311,N_32276);
nor U32550 (N_32550,N_32344,N_32232);
nor U32551 (N_32551,N_32159,N_32376);
xnor U32552 (N_32552,N_32359,N_32240);
nand U32553 (N_32553,N_32349,N_32039);
nor U32554 (N_32554,N_32331,N_32416);
nor U32555 (N_32555,N_32302,N_32171);
xnor U32556 (N_32556,N_32329,N_32492);
nand U32557 (N_32557,N_32424,N_32023);
xor U32558 (N_32558,N_32214,N_32247);
and U32559 (N_32559,N_32257,N_32459);
xnor U32560 (N_32560,N_32288,N_32233);
xor U32561 (N_32561,N_32388,N_32220);
nand U32562 (N_32562,N_32087,N_32314);
and U32563 (N_32563,N_32269,N_32266);
or U32564 (N_32564,N_32041,N_32273);
and U32565 (N_32565,N_32397,N_32353);
nor U32566 (N_32566,N_32379,N_32243);
xnor U32567 (N_32567,N_32252,N_32370);
or U32568 (N_32568,N_32339,N_32211);
nand U32569 (N_32569,N_32307,N_32238);
and U32570 (N_32570,N_32468,N_32383);
nand U32571 (N_32571,N_32200,N_32470);
nand U32572 (N_32572,N_32225,N_32418);
nand U32573 (N_32573,N_32355,N_32209);
and U32574 (N_32574,N_32042,N_32461);
and U32575 (N_32575,N_32352,N_32272);
and U32576 (N_32576,N_32045,N_32196);
or U32577 (N_32577,N_32262,N_32466);
or U32578 (N_32578,N_32054,N_32395);
nor U32579 (N_32579,N_32491,N_32237);
or U32580 (N_32580,N_32180,N_32104);
xnor U32581 (N_32581,N_32132,N_32324);
and U32582 (N_32582,N_32071,N_32065);
nor U32583 (N_32583,N_32231,N_32439);
nand U32584 (N_32584,N_32115,N_32070);
xor U32585 (N_32585,N_32018,N_32033);
xor U32586 (N_32586,N_32289,N_32186);
nand U32587 (N_32587,N_32326,N_32137);
nor U32588 (N_32588,N_32412,N_32494);
nand U32589 (N_32589,N_32474,N_32128);
nand U32590 (N_32590,N_32382,N_32384);
or U32591 (N_32591,N_32082,N_32356);
nor U32592 (N_32592,N_32169,N_32052);
or U32593 (N_32593,N_32059,N_32265);
and U32594 (N_32594,N_32369,N_32437);
nor U32595 (N_32595,N_32487,N_32207);
nand U32596 (N_32596,N_32114,N_32178);
nand U32597 (N_32597,N_32389,N_32436);
and U32598 (N_32598,N_32096,N_32399);
nor U32599 (N_32599,N_32166,N_32112);
or U32600 (N_32600,N_32304,N_32358);
nand U32601 (N_32601,N_32130,N_32183);
xnor U32602 (N_32602,N_32134,N_32414);
and U32603 (N_32603,N_32425,N_32189);
nand U32604 (N_32604,N_32241,N_32310);
and U32605 (N_32605,N_32154,N_32174);
nand U32606 (N_32606,N_32029,N_32165);
nand U32607 (N_32607,N_32221,N_32267);
or U32608 (N_32608,N_32090,N_32179);
nand U32609 (N_32609,N_32242,N_32374);
nor U32610 (N_32610,N_32167,N_32380);
nor U32611 (N_32611,N_32139,N_32484);
nand U32612 (N_32612,N_32164,N_32024);
or U32613 (N_32613,N_32422,N_32386);
nor U32614 (N_32614,N_32083,N_32199);
nand U32615 (N_32615,N_32026,N_32431);
nand U32616 (N_32616,N_32206,N_32100);
and U32617 (N_32617,N_32005,N_32444);
or U32618 (N_32618,N_32396,N_32485);
and U32619 (N_32619,N_32481,N_32031);
nor U32620 (N_32620,N_32244,N_32404);
nor U32621 (N_32621,N_32475,N_32205);
nand U32622 (N_32622,N_32372,N_32428);
or U32623 (N_32623,N_32036,N_32442);
and U32624 (N_32624,N_32080,N_32079);
nand U32625 (N_32625,N_32473,N_32131);
and U32626 (N_32626,N_32105,N_32327);
nor U32627 (N_32627,N_32050,N_32400);
and U32628 (N_32628,N_32493,N_32019);
nand U32629 (N_32629,N_32275,N_32127);
and U32630 (N_32630,N_32016,N_32140);
and U32631 (N_32631,N_32381,N_32126);
nand U32632 (N_32632,N_32149,N_32342);
and U32633 (N_32633,N_32097,N_32234);
nand U32634 (N_32634,N_32495,N_32499);
and U32635 (N_32635,N_32394,N_32102);
nor U32636 (N_32636,N_32250,N_32084);
nor U32637 (N_32637,N_32248,N_32462);
nor U32638 (N_32638,N_32099,N_32253);
xor U32639 (N_32639,N_32347,N_32103);
or U32640 (N_32640,N_32120,N_32088);
nor U32641 (N_32641,N_32440,N_32204);
and U32642 (N_32642,N_32280,N_32390);
or U32643 (N_32643,N_32066,N_32061);
and U32644 (N_32644,N_32463,N_32142);
nand U32645 (N_32645,N_32315,N_32184);
or U32646 (N_32646,N_32335,N_32188);
and U32647 (N_32647,N_32322,N_32046);
xor U32648 (N_32648,N_32021,N_32245);
and U32649 (N_32649,N_32063,N_32393);
nand U32650 (N_32650,N_32398,N_32483);
and U32651 (N_32651,N_32201,N_32391);
nor U32652 (N_32652,N_32278,N_32290);
or U32653 (N_32653,N_32057,N_32141);
nand U32654 (N_32654,N_32020,N_32330);
nand U32655 (N_32655,N_32281,N_32472);
and U32656 (N_32656,N_32215,N_32089);
nand U32657 (N_32657,N_32415,N_32072);
nand U32658 (N_32658,N_32236,N_32455);
nand U32659 (N_32659,N_32058,N_32261);
nor U32660 (N_32660,N_32360,N_32150);
and U32661 (N_32661,N_32037,N_32371);
and U32662 (N_32662,N_32086,N_32471);
and U32663 (N_32663,N_32125,N_32313);
nand U32664 (N_32664,N_32153,N_32226);
and U32665 (N_32665,N_32402,N_32447);
and U32666 (N_32666,N_32162,N_32177);
and U32667 (N_32667,N_32405,N_32194);
nand U32668 (N_32668,N_32218,N_32121);
nand U32669 (N_32669,N_32191,N_32345);
nand U32670 (N_32670,N_32465,N_32069);
or U32671 (N_32671,N_32055,N_32147);
nor U32672 (N_32672,N_32279,N_32091);
nand U32673 (N_32673,N_32239,N_32181);
and U32674 (N_32674,N_32048,N_32441);
nor U32675 (N_32675,N_32014,N_32337);
nor U32676 (N_32676,N_32098,N_32003);
or U32677 (N_32677,N_32497,N_32192);
nor U32678 (N_32678,N_32062,N_32417);
nor U32679 (N_32679,N_32175,N_32138);
and U32680 (N_32680,N_32053,N_32108);
xnor U32681 (N_32681,N_32158,N_32482);
or U32682 (N_32682,N_32317,N_32354);
and U32683 (N_32683,N_32258,N_32316);
nor U32684 (N_32684,N_32452,N_32111);
or U32685 (N_32685,N_32336,N_32198);
nand U32686 (N_32686,N_32480,N_32419);
or U32687 (N_32687,N_32022,N_32170);
and U32688 (N_32688,N_32498,N_32264);
or U32689 (N_32689,N_32025,N_32124);
nand U32690 (N_32690,N_32328,N_32076);
nor U32691 (N_32691,N_32350,N_32034);
or U32692 (N_32692,N_32216,N_32410);
xnor U32693 (N_32693,N_32421,N_32012);
or U32694 (N_32694,N_32068,N_32185);
nor U32695 (N_32695,N_32285,N_32365);
and U32696 (N_32696,N_32457,N_32161);
and U32697 (N_32697,N_32496,N_32451);
and U32698 (N_32698,N_32081,N_32409);
nand U32699 (N_32699,N_32291,N_32015);
or U32700 (N_32700,N_32368,N_32030);
or U32701 (N_32701,N_32117,N_32133);
nand U32702 (N_32702,N_32182,N_32426);
nor U32703 (N_32703,N_32286,N_32092);
and U32704 (N_32704,N_32318,N_32375);
nand U32705 (N_32705,N_32298,N_32110);
nor U32706 (N_32706,N_32251,N_32392);
and U32707 (N_32707,N_32135,N_32078);
nand U32708 (N_32708,N_32202,N_32469);
nor U32709 (N_32709,N_32228,N_32044);
or U32710 (N_32710,N_32456,N_32373);
and U32711 (N_32711,N_32143,N_32408);
nand U32712 (N_32712,N_32040,N_32038);
and U32713 (N_32713,N_32028,N_32107);
and U32714 (N_32714,N_32464,N_32343);
or U32715 (N_32715,N_32476,N_32094);
or U32716 (N_32716,N_32450,N_32287);
and U32717 (N_32717,N_32168,N_32323);
and U32718 (N_32718,N_32145,N_32256);
nand U32719 (N_32719,N_32193,N_32151);
and U32720 (N_32720,N_32378,N_32433);
and U32721 (N_32721,N_32109,N_32364);
nand U32722 (N_32722,N_32009,N_32432);
nand U32723 (N_32723,N_32208,N_32338);
or U32724 (N_32724,N_32411,N_32213);
and U32725 (N_32725,N_32254,N_32332);
or U32726 (N_32726,N_32387,N_32007);
or U32727 (N_32727,N_32155,N_32306);
or U32728 (N_32728,N_32460,N_32334);
nor U32729 (N_32729,N_32047,N_32000);
or U32730 (N_32730,N_32157,N_32271);
or U32731 (N_32731,N_32077,N_32106);
nor U32732 (N_32732,N_32445,N_32305);
or U32733 (N_32733,N_32259,N_32296);
nand U32734 (N_32734,N_32006,N_32301);
or U32735 (N_32735,N_32011,N_32357);
and U32736 (N_32736,N_32013,N_32227);
or U32737 (N_32737,N_32235,N_32340);
xor U32738 (N_32738,N_32160,N_32136);
nor U32739 (N_32739,N_32489,N_32362);
and U32740 (N_32740,N_32320,N_32363);
and U32741 (N_32741,N_32282,N_32351);
nor U32742 (N_32742,N_32367,N_32309);
and U32743 (N_32743,N_32060,N_32229);
nor U32744 (N_32744,N_32085,N_32255);
or U32745 (N_32745,N_32303,N_32446);
nor U32746 (N_32746,N_32224,N_32479);
or U32747 (N_32747,N_32195,N_32407);
nor U32748 (N_32748,N_32156,N_32118);
or U32749 (N_32749,N_32420,N_32366);
nor U32750 (N_32750,N_32085,N_32496);
nand U32751 (N_32751,N_32087,N_32293);
nor U32752 (N_32752,N_32116,N_32083);
xnor U32753 (N_32753,N_32333,N_32229);
nor U32754 (N_32754,N_32095,N_32169);
nand U32755 (N_32755,N_32133,N_32391);
nor U32756 (N_32756,N_32454,N_32192);
xor U32757 (N_32757,N_32454,N_32364);
or U32758 (N_32758,N_32275,N_32036);
or U32759 (N_32759,N_32429,N_32241);
nand U32760 (N_32760,N_32293,N_32152);
nand U32761 (N_32761,N_32203,N_32361);
or U32762 (N_32762,N_32059,N_32257);
or U32763 (N_32763,N_32273,N_32220);
or U32764 (N_32764,N_32272,N_32372);
nand U32765 (N_32765,N_32154,N_32390);
nor U32766 (N_32766,N_32154,N_32441);
nand U32767 (N_32767,N_32384,N_32118);
nand U32768 (N_32768,N_32457,N_32186);
nor U32769 (N_32769,N_32087,N_32062);
or U32770 (N_32770,N_32294,N_32396);
or U32771 (N_32771,N_32007,N_32416);
or U32772 (N_32772,N_32127,N_32339);
nand U32773 (N_32773,N_32218,N_32164);
nor U32774 (N_32774,N_32087,N_32138);
or U32775 (N_32775,N_32379,N_32205);
or U32776 (N_32776,N_32351,N_32363);
or U32777 (N_32777,N_32295,N_32317);
nand U32778 (N_32778,N_32155,N_32192);
nand U32779 (N_32779,N_32146,N_32116);
and U32780 (N_32780,N_32487,N_32316);
nor U32781 (N_32781,N_32184,N_32401);
nor U32782 (N_32782,N_32045,N_32331);
or U32783 (N_32783,N_32133,N_32020);
or U32784 (N_32784,N_32484,N_32488);
nor U32785 (N_32785,N_32273,N_32188);
nor U32786 (N_32786,N_32268,N_32247);
or U32787 (N_32787,N_32305,N_32091);
and U32788 (N_32788,N_32014,N_32104);
and U32789 (N_32789,N_32171,N_32236);
xor U32790 (N_32790,N_32203,N_32267);
or U32791 (N_32791,N_32286,N_32220);
or U32792 (N_32792,N_32423,N_32086);
nand U32793 (N_32793,N_32395,N_32068);
nand U32794 (N_32794,N_32393,N_32243);
and U32795 (N_32795,N_32068,N_32061);
nand U32796 (N_32796,N_32385,N_32311);
nor U32797 (N_32797,N_32205,N_32020);
and U32798 (N_32798,N_32330,N_32438);
and U32799 (N_32799,N_32376,N_32035);
or U32800 (N_32800,N_32498,N_32047);
or U32801 (N_32801,N_32147,N_32451);
nor U32802 (N_32802,N_32119,N_32392);
nor U32803 (N_32803,N_32220,N_32342);
and U32804 (N_32804,N_32357,N_32372);
or U32805 (N_32805,N_32446,N_32205);
or U32806 (N_32806,N_32170,N_32210);
and U32807 (N_32807,N_32172,N_32182);
xor U32808 (N_32808,N_32425,N_32459);
nand U32809 (N_32809,N_32415,N_32235);
or U32810 (N_32810,N_32299,N_32086);
and U32811 (N_32811,N_32306,N_32399);
nand U32812 (N_32812,N_32272,N_32156);
nor U32813 (N_32813,N_32376,N_32283);
or U32814 (N_32814,N_32411,N_32124);
or U32815 (N_32815,N_32429,N_32125);
and U32816 (N_32816,N_32491,N_32137);
or U32817 (N_32817,N_32411,N_32091);
xnor U32818 (N_32818,N_32096,N_32442);
nand U32819 (N_32819,N_32296,N_32278);
and U32820 (N_32820,N_32486,N_32311);
and U32821 (N_32821,N_32411,N_32210);
or U32822 (N_32822,N_32248,N_32268);
xnor U32823 (N_32823,N_32101,N_32163);
xnor U32824 (N_32824,N_32151,N_32249);
nand U32825 (N_32825,N_32298,N_32028);
nand U32826 (N_32826,N_32477,N_32362);
or U32827 (N_32827,N_32142,N_32442);
or U32828 (N_32828,N_32474,N_32045);
nor U32829 (N_32829,N_32367,N_32115);
nand U32830 (N_32830,N_32001,N_32184);
nor U32831 (N_32831,N_32357,N_32166);
nor U32832 (N_32832,N_32130,N_32123);
xnor U32833 (N_32833,N_32427,N_32229);
nand U32834 (N_32834,N_32117,N_32067);
or U32835 (N_32835,N_32039,N_32065);
xnor U32836 (N_32836,N_32202,N_32116);
nor U32837 (N_32837,N_32340,N_32017);
or U32838 (N_32838,N_32185,N_32490);
nand U32839 (N_32839,N_32051,N_32368);
xnor U32840 (N_32840,N_32164,N_32489);
or U32841 (N_32841,N_32299,N_32380);
and U32842 (N_32842,N_32118,N_32442);
nor U32843 (N_32843,N_32026,N_32079);
nor U32844 (N_32844,N_32056,N_32084);
and U32845 (N_32845,N_32376,N_32046);
nand U32846 (N_32846,N_32024,N_32221);
nand U32847 (N_32847,N_32258,N_32261);
nand U32848 (N_32848,N_32021,N_32053);
or U32849 (N_32849,N_32213,N_32062);
or U32850 (N_32850,N_32096,N_32336);
nand U32851 (N_32851,N_32207,N_32291);
nor U32852 (N_32852,N_32486,N_32235);
xnor U32853 (N_32853,N_32381,N_32049);
xnor U32854 (N_32854,N_32173,N_32248);
xnor U32855 (N_32855,N_32333,N_32363);
nand U32856 (N_32856,N_32276,N_32056);
nor U32857 (N_32857,N_32428,N_32414);
or U32858 (N_32858,N_32362,N_32161);
nor U32859 (N_32859,N_32029,N_32125);
nand U32860 (N_32860,N_32459,N_32355);
or U32861 (N_32861,N_32260,N_32350);
and U32862 (N_32862,N_32207,N_32119);
or U32863 (N_32863,N_32304,N_32035);
and U32864 (N_32864,N_32301,N_32198);
and U32865 (N_32865,N_32334,N_32276);
nand U32866 (N_32866,N_32214,N_32396);
nand U32867 (N_32867,N_32112,N_32052);
and U32868 (N_32868,N_32230,N_32100);
and U32869 (N_32869,N_32146,N_32487);
or U32870 (N_32870,N_32356,N_32453);
nand U32871 (N_32871,N_32452,N_32395);
nor U32872 (N_32872,N_32140,N_32290);
or U32873 (N_32873,N_32461,N_32089);
nor U32874 (N_32874,N_32492,N_32437);
or U32875 (N_32875,N_32091,N_32359);
and U32876 (N_32876,N_32343,N_32049);
and U32877 (N_32877,N_32084,N_32307);
or U32878 (N_32878,N_32199,N_32020);
nand U32879 (N_32879,N_32125,N_32188);
or U32880 (N_32880,N_32363,N_32015);
and U32881 (N_32881,N_32064,N_32285);
or U32882 (N_32882,N_32246,N_32431);
nand U32883 (N_32883,N_32132,N_32052);
and U32884 (N_32884,N_32165,N_32420);
or U32885 (N_32885,N_32026,N_32258);
nor U32886 (N_32886,N_32296,N_32379);
xor U32887 (N_32887,N_32372,N_32196);
and U32888 (N_32888,N_32078,N_32210);
nand U32889 (N_32889,N_32103,N_32445);
and U32890 (N_32890,N_32217,N_32250);
nand U32891 (N_32891,N_32319,N_32497);
xnor U32892 (N_32892,N_32347,N_32284);
xnor U32893 (N_32893,N_32089,N_32253);
and U32894 (N_32894,N_32344,N_32082);
xnor U32895 (N_32895,N_32082,N_32485);
nand U32896 (N_32896,N_32441,N_32275);
xnor U32897 (N_32897,N_32424,N_32380);
nand U32898 (N_32898,N_32270,N_32494);
and U32899 (N_32899,N_32179,N_32402);
nor U32900 (N_32900,N_32100,N_32026);
nand U32901 (N_32901,N_32392,N_32101);
nand U32902 (N_32902,N_32257,N_32229);
and U32903 (N_32903,N_32355,N_32468);
and U32904 (N_32904,N_32171,N_32303);
nand U32905 (N_32905,N_32115,N_32253);
nand U32906 (N_32906,N_32170,N_32031);
or U32907 (N_32907,N_32277,N_32496);
nand U32908 (N_32908,N_32455,N_32123);
or U32909 (N_32909,N_32183,N_32438);
nor U32910 (N_32910,N_32324,N_32333);
nor U32911 (N_32911,N_32213,N_32450);
nor U32912 (N_32912,N_32359,N_32141);
and U32913 (N_32913,N_32292,N_32066);
nor U32914 (N_32914,N_32393,N_32446);
or U32915 (N_32915,N_32343,N_32296);
or U32916 (N_32916,N_32458,N_32240);
nand U32917 (N_32917,N_32389,N_32063);
xor U32918 (N_32918,N_32265,N_32006);
or U32919 (N_32919,N_32102,N_32362);
and U32920 (N_32920,N_32431,N_32381);
nor U32921 (N_32921,N_32413,N_32102);
or U32922 (N_32922,N_32440,N_32241);
or U32923 (N_32923,N_32129,N_32032);
and U32924 (N_32924,N_32224,N_32218);
nor U32925 (N_32925,N_32003,N_32211);
and U32926 (N_32926,N_32191,N_32101);
nor U32927 (N_32927,N_32177,N_32071);
or U32928 (N_32928,N_32441,N_32408);
nor U32929 (N_32929,N_32290,N_32133);
or U32930 (N_32930,N_32089,N_32329);
or U32931 (N_32931,N_32085,N_32102);
or U32932 (N_32932,N_32234,N_32238);
nor U32933 (N_32933,N_32086,N_32391);
and U32934 (N_32934,N_32291,N_32496);
or U32935 (N_32935,N_32058,N_32122);
and U32936 (N_32936,N_32107,N_32330);
nand U32937 (N_32937,N_32360,N_32375);
nand U32938 (N_32938,N_32324,N_32437);
or U32939 (N_32939,N_32391,N_32403);
or U32940 (N_32940,N_32304,N_32375);
nand U32941 (N_32941,N_32300,N_32096);
and U32942 (N_32942,N_32346,N_32052);
nor U32943 (N_32943,N_32343,N_32131);
nand U32944 (N_32944,N_32119,N_32102);
nand U32945 (N_32945,N_32347,N_32402);
nand U32946 (N_32946,N_32045,N_32057);
nand U32947 (N_32947,N_32377,N_32116);
nand U32948 (N_32948,N_32176,N_32309);
or U32949 (N_32949,N_32026,N_32044);
nor U32950 (N_32950,N_32314,N_32453);
nor U32951 (N_32951,N_32393,N_32009);
nand U32952 (N_32952,N_32283,N_32298);
xor U32953 (N_32953,N_32019,N_32379);
xnor U32954 (N_32954,N_32083,N_32000);
xor U32955 (N_32955,N_32421,N_32087);
nand U32956 (N_32956,N_32267,N_32040);
and U32957 (N_32957,N_32452,N_32212);
and U32958 (N_32958,N_32353,N_32392);
xor U32959 (N_32959,N_32226,N_32014);
nand U32960 (N_32960,N_32246,N_32103);
nand U32961 (N_32961,N_32131,N_32139);
or U32962 (N_32962,N_32177,N_32169);
or U32963 (N_32963,N_32023,N_32439);
nand U32964 (N_32964,N_32462,N_32464);
nand U32965 (N_32965,N_32194,N_32233);
or U32966 (N_32966,N_32295,N_32456);
nor U32967 (N_32967,N_32465,N_32066);
or U32968 (N_32968,N_32359,N_32400);
and U32969 (N_32969,N_32438,N_32485);
or U32970 (N_32970,N_32433,N_32483);
nand U32971 (N_32971,N_32438,N_32253);
xor U32972 (N_32972,N_32231,N_32042);
nor U32973 (N_32973,N_32134,N_32072);
or U32974 (N_32974,N_32123,N_32100);
xnor U32975 (N_32975,N_32134,N_32451);
or U32976 (N_32976,N_32370,N_32154);
nor U32977 (N_32977,N_32282,N_32129);
or U32978 (N_32978,N_32242,N_32081);
and U32979 (N_32979,N_32210,N_32053);
nand U32980 (N_32980,N_32212,N_32025);
nor U32981 (N_32981,N_32458,N_32176);
nand U32982 (N_32982,N_32180,N_32305);
or U32983 (N_32983,N_32461,N_32341);
or U32984 (N_32984,N_32200,N_32086);
nor U32985 (N_32985,N_32003,N_32461);
and U32986 (N_32986,N_32478,N_32167);
and U32987 (N_32987,N_32340,N_32112);
and U32988 (N_32988,N_32051,N_32405);
nand U32989 (N_32989,N_32065,N_32472);
xor U32990 (N_32990,N_32063,N_32457);
nand U32991 (N_32991,N_32323,N_32398);
nand U32992 (N_32992,N_32145,N_32189);
nand U32993 (N_32993,N_32491,N_32438);
nand U32994 (N_32994,N_32085,N_32196);
xor U32995 (N_32995,N_32018,N_32053);
or U32996 (N_32996,N_32060,N_32486);
and U32997 (N_32997,N_32110,N_32496);
and U32998 (N_32998,N_32093,N_32374);
or U32999 (N_32999,N_32101,N_32365);
xor U33000 (N_33000,N_32696,N_32562);
and U33001 (N_33001,N_32888,N_32845);
nor U33002 (N_33002,N_32789,N_32852);
nand U33003 (N_33003,N_32720,N_32620);
and U33004 (N_33004,N_32790,N_32531);
nor U33005 (N_33005,N_32936,N_32887);
nor U33006 (N_33006,N_32842,N_32932);
nor U33007 (N_33007,N_32925,N_32642);
nand U33008 (N_33008,N_32804,N_32638);
or U33009 (N_33009,N_32816,N_32998);
nor U33010 (N_33010,N_32666,N_32954);
and U33011 (N_33011,N_32651,N_32873);
or U33012 (N_33012,N_32840,N_32534);
and U33013 (N_33013,N_32911,N_32568);
nand U33014 (N_33014,N_32935,N_32918);
nand U33015 (N_33015,N_32754,N_32828);
nor U33016 (N_33016,N_32793,N_32853);
or U33017 (N_33017,N_32509,N_32897);
nor U33018 (N_33018,N_32519,N_32709);
nor U33019 (N_33019,N_32907,N_32612);
xnor U33020 (N_33020,N_32841,N_32871);
and U33021 (N_33021,N_32619,N_32506);
and U33022 (N_33022,N_32933,N_32719);
and U33023 (N_33023,N_32737,N_32717);
or U33024 (N_33024,N_32515,N_32953);
and U33025 (N_33025,N_32715,N_32997);
and U33026 (N_33026,N_32712,N_32780);
nand U33027 (N_33027,N_32652,N_32859);
and U33028 (N_33028,N_32673,N_32931);
nand U33029 (N_33029,N_32617,N_32872);
nand U33030 (N_33030,N_32661,N_32710);
nand U33031 (N_33031,N_32885,N_32960);
nor U33032 (N_33032,N_32849,N_32536);
or U33033 (N_33033,N_32810,N_32660);
nor U33034 (N_33034,N_32833,N_32518);
and U33035 (N_33035,N_32641,N_32805);
nand U33036 (N_33036,N_32613,N_32606);
nand U33037 (N_33037,N_32870,N_32922);
nor U33038 (N_33038,N_32713,N_32502);
nor U33039 (N_33039,N_32543,N_32995);
nand U33040 (N_33040,N_32700,N_32544);
and U33041 (N_33041,N_32899,N_32827);
and U33042 (N_33042,N_32671,N_32588);
nand U33043 (N_33043,N_32733,N_32591);
and U33044 (N_33044,N_32572,N_32803);
or U33045 (N_33045,N_32831,N_32799);
or U33046 (N_33046,N_32996,N_32843);
nand U33047 (N_33047,N_32917,N_32622);
nand U33048 (N_33048,N_32795,N_32743);
or U33049 (N_33049,N_32756,N_32898);
xnor U33050 (N_33050,N_32824,N_32635);
and U33051 (N_33051,N_32614,N_32627);
or U33052 (N_33052,N_32958,N_32658);
nand U33053 (N_33053,N_32758,N_32526);
and U33054 (N_33054,N_32869,N_32787);
nand U33055 (N_33055,N_32556,N_32516);
and U33056 (N_33056,N_32991,N_32848);
nor U33057 (N_33057,N_32929,N_32744);
nor U33058 (N_33058,N_32639,N_32826);
nor U33059 (N_33059,N_32592,N_32708);
and U33060 (N_33060,N_32863,N_32631);
or U33061 (N_33061,N_32574,N_32867);
and U33062 (N_33062,N_32818,N_32610);
nor U33063 (N_33063,N_32988,N_32676);
and U33064 (N_33064,N_32747,N_32906);
and U33065 (N_33065,N_32584,N_32711);
nand U33066 (N_33066,N_32763,N_32669);
nor U33067 (N_33067,N_32728,N_32880);
nand U33068 (N_33068,N_32674,N_32655);
nor U33069 (N_33069,N_32821,N_32685);
nor U33070 (N_33070,N_32510,N_32861);
and U33071 (N_33071,N_32974,N_32616);
nor U33072 (N_33072,N_32981,N_32830);
nand U33073 (N_33073,N_32800,N_32894);
nor U33074 (N_33074,N_32521,N_32792);
xnor U33075 (N_33075,N_32788,N_32844);
and U33076 (N_33076,N_32999,N_32607);
nand U33077 (N_33077,N_32942,N_32694);
nand U33078 (N_33078,N_32774,N_32908);
nor U33079 (N_33079,N_32739,N_32905);
and U33080 (N_33080,N_32609,N_32555);
nand U33081 (N_33081,N_32811,N_32773);
nor U33082 (N_33082,N_32689,N_32862);
xor U33083 (N_33083,N_32921,N_32893);
nand U33084 (N_33084,N_32702,N_32883);
nand U33085 (N_33085,N_32626,N_32819);
and U33086 (N_33086,N_32847,N_32570);
or U33087 (N_33087,N_32505,N_32923);
nor U33088 (N_33088,N_32913,N_32822);
nor U33089 (N_33089,N_32820,N_32663);
nand U33090 (N_33090,N_32692,N_32881);
and U33091 (N_33091,N_32538,N_32909);
and U33092 (N_33092,N_32926,N_32734);
nor U33093 (N_33093,N_32767,N_32884);
nor U33094 (N_33094,N_32973,N_32864);
or U33095 (N_33095,N_32672,N_32813);
or U33096 (N_33096,N_32546,N_32966);
nor U33097 (N_33097,N_32762,N_32511);
nand U33098 (N_33098,N_32624,N_32784);
nor U33099 (N_33099,N_32961,N_32984);
nor U33100 (N_33100,N_32545,N_32508);
nor U33101 (N_33101,N_32723,N_32523);
and U33102 (N_33102,N_32777,N_32633);
nand U33103 (N_33103,N_32527,N_32731);
nor U33104 (N_33104,N_32751,N_32697);
and U33105 (N_33105,N_32722,N_32992);
nor U33106 (N_33106,N_32794,N_32892);
and U33107 (N_33107,N_32769,N_32920);
nor U33108 (N_33108,N_32732,N_32834);
xnor U33109 (N_33109,N_32979,N_32916);
nor U33110 (N_33110,N_32569,N_32559);
and U33111 (N_33111,N_32659,N_32928);
nor U33112 (N_33112,N_32947,N_32977);
or U33113 (N_33113,N_32962,N_32703);
and U33114 (N_33114,N_32890,N_32832);
or U33115 (N_33115,N_32736,N_32782);
or U33116 (N_33116,N_32567,N_32698);
nor U33117 (N_33117,N_32576,N_32677);
and U33118 (N_33118,N_32781,N_32707);
and U33119 (N_33119,N_32989,N_32740);
nand U33120 (N_33120,N_32771,N_32955);
nand U33121 (N_33121,N_32725,N_32786);
xnor U33122 (N_33122,N_32726,N_32939);
nand U33123 (N_33123,N_32640,N_32968);
nand U33124 (N_33124,N_32500,N_32839);
or U33125 (N_33125,N_32687,N_32772);
or U33126 (N_33126,N_32889,N_32730);
or U33127 (N_33127,N_32653,N_32539);
or U33128 (N_33128,N_32682,N_32625);
nor U33129 (N_33129,N_32757,N_32667);
nand U33130 (N_33130,N_32552,N_32943);
or U33131 (N_33131,N_32716,N_32656);
and U33132 (N_33132,N_32724,N_32927);
nand U33133 (N_33133,N_32577,N_32980);
nand U33134 (N_33134,N_32578,N_32650);
nor U33135 (N_33135,N_32860,N_32948);
nand U33136 (N_33136,N_32895,N_32851);
and U33137 (N_33137,N_32823,N_32742);
nor U33138 (N_33138,N_32985,N_32611);
nand U33139 (N_33139,N_32814,N_32681);
nand U33140 (N_33140,N_32746,N_32603);
nor U33141 (N_33141,N_32530,N_32798);
or U33142 (N_33142,N_32680,N_32657);
and U33143 (N_33143,N_32541,N_32678);
and U33144 (N_33144,N_32951,N_32874);
or U33145 (N_33145,N_32587,N_32778);
or U33146 (N_33146,N_32704,N_32670);
nand U33147 (N_33147,N_32718,N_32558);
xnor U33148 (N_33148,N_32665,N_32924);
and U33149 (N_33149,N_32561,N_32982);
and U33150 (N_33150,N_32914,N_32598);
xnor U33151 (N_33151,N_32815,N_32886);
nand U33152 (N_33152,N_32934,N_32634);
nor U33153 (N_33153,N_32632,N_32972);
or U33154 (N_33154,N_32801,N_32808);
nand U33155 (N_33155,N_32532,N_32683);
nand U33156 (N_33156,N_32593,N_32735);
or U33157 (N_33157,N_32866,N_32940);
or U33158 (N_33158,N_32791,N_32891);
nor U33159 (N_33159,N_32507,N_32595);
nor U33160 (N_33160,N_32965,N_32668);
or U33161 (N_33161,N_32761,N_32759);
and U33162 (N_33162,N_32684,N_32802);
or U33163 (N_33163,N_32705,N_32952);
nand U33164 (N_33164,N_32590,N_32949);
or U33165 (N_33165,N_32994,N_32749);
and U33166 (N_33166,N_32957,N_32812);
and U33167 (N_33167,N_32797,N_32528);
or U33168 (N_33168,N_32706,N_32693);
and U33169 (N_33169,N_32760,N_32904);
or U33170 (N_33170,N_32540,N_32875);
and U33171 (N_33171,N_32636,N_32548);
and U33172 (N_33172,N_32647,N_32535);
nor U33173 (N_33173,N_32838,N_32876);
nand U33174 (N_33174,N_32770,N_32741);
and U33175 (N_33175,N_32857,N_32501);
or U33176 (N_33176,N_32643,N_32686);
xnor U33177 (N_33177,N_32779,N_32542);
and U33178 (N_33178,N_32504,N_32768);
or U33179 (N_33179,N_32855,N_32571);
and U33180 (N_33180,N_32529,N_32560);
nor U33181 (N_33181,N_32817,N_32554);
and U33182 (N_33182,N_32628,N_32941);
or U33183 (N_33183,N_32604,N_32945);
and U33184 (N_33184,N_32512,N_32664);
nand U33185 (N_33185,N_32878,N_32902);
and U33186 (N_33186,N_32695,N_32806);
nor U33187 (N_33187,N_32675,N_32919);
xnor U33188 (N_33188,N_32573,N_32755);
xnor U33189 (N_33189,N_32944,N_32809);
nor U33190 (N_33190,N_32580,N_32901);
nor U33191 (N_33191,N_32721,N_32608);
and U33192 (N_33192,N_32752,N_32796);
or U33193 (N_33193,N_32856,N_32564);
nand U33194 (N_33194,N_32950,N_32594);
and U33195 (N_33195,N_32766,N_32986);
xor U33196 (N_33196,N_32550,N_32520);
and U33197 (N_33197,N_32525,N_32637);
and U33198 (N_33198,N_32835,N_32978);
and U33199 (N_33199,N_32727,N_32644);
nand U33200 (N_33200,N_32753,N_32524);
nor U33201 (N_33201,N_32836,N_32618);
and U33202 (N_33202,N_32900,N_32621);
nor U33203 (N_33203,N_32854,N_32937);
xor U33204 (N_33204,N_32589,N_32990);
nand U33205 (N_33205,N_32956,N_32879);
xor U33206 (N_33206,N_32522,N_32701);
nor U33207 (N_33207,N_32581,N_32970);
nand U33208 (N_33208,N_32547,N_32776);
xor U33209 (N_33209,N_32691,N_32969);
nand U33210 (N_33210,N_32513,N_32976);
and U33211 (N_33211,N_32865,N_32582);
or U33212 (N_33212,N_32915,N_32565);
or U33213 (N_33213,N_32764,N_32649);
and U33214 (N_33214,N_32983,N_32785);
and U33215 (N_33215,N_32971,N_32585);
nand U33216 (N_33216,N_32583,N_32517);
nor U33217 (N_33217,N_32605,N_32930);
nor U33218 (N_33218,N_32553,N_32600);
or U33219 (N_33219,N_32783,N_32503);
nor U33220 (N_33220,N_32690,N_32679);
xor U33221 (N_33221,N_32745,N_32748);
and U33222 (N_33222,N_32596,N_32896);
nand U33223 (N_33223,N_32699,N_32566);
and U33224 (N_33224,N_32597,N_32575);
or U33225 (N_33225,N_32825,N_32903);
and U33226 (N_33226,N_32630,N_32714);
nand U33227 (N_33227,N_32563,N_32551);
nor U33228 (N_33228,N_32579,N_32537);
and U33229 (N_33229,N_32750,N_32601);
xor U33230 (N_33230,N_32645,N_32615);
and U33231 (N_33231,N_32557,N_32858);
nor U33232 (N_33232,N_32602,N_32646);
and U33233 (N_33233,N_32837,N_32738);
and U33234 (N_33234,N_32963,N_32882);
and U33235 (N_33235,N_32533,N_32549);
nand U33236 (N_33236,N_32868,N_32623);
or U33237 (N_33237,N_32846,N_32912);
or U33238 (N_33238,N_32877,N_32688);
or U33239 (N_33239,N_32662,N_32514);
nor U33240 (N_33240,N_32946,N_32829);
nand U33241 (N_33241,N_32775,N_32967);
and U33242 (N_33242,N_32910,N_32729);
or U33243 (N_33243,N_32959,N_32648);
or U33244 (N_33244,N_32993,N_32964);
and U33245 (N_33245,N_32850,N_32807);
or U33246 (N_33246,N_32987,N_32599);
nor U33247 (N_33247,N_32629,N_32938);
nand U33248 (N_33248,N_32654,N_32765);
nor U33249 (N_33249,N_32586,N_32975);
nand U33250 (N_33250,N_32848,N_32861);
nor U33251 (N_33251,N_32651,N_32865);
or U33252 (N_33252,N_32611,N_32927);
xnor U33253 (N_33253,N_32906,N_32656);
or U33254 (N_33254,N_32794,N_32788);
and U33255 (N_33255,N_32782,N_32953);
xor U33256 (N_33256,N_32848,N_32871);
and U33257 (N_33257,N_32501,N_32929);
and U33258 (N_33258,N_32816,N_32933);
xnor U33259 (N_33259,N_32542,N_32720);
nand U33260 (N_33260,N_32556,N_32923);
nor U33261 (N_33261,N_32637,N_32871);
or U33262 (N_33262,N_32926,N_32981);
nand U33263 (N_33263,N_32909,N_32569);
and U33264 (N_33264,N_32953,N_32879);
or U33265 (N_33265,N_32620,N_32547);
and U33266 (N_33266,N_32728,N_32833);
xor U33267 (N_33267,N_32788,N_32886);
or U33268 (N_33268,N_32725,N_32700);
nor U33269 (N_33269,N_32864,N_32946);
and U33270 (N_33270,N_32767,N_32987);
and U33271 (N_33271,N_32644,N_32531);
xor U33272 (N_33272,N_32557,N_32763);
or U33273 (N_33273,N_32999,N_32632);
or U33274 (N_33274,N_32890,N_32540);
nor U33275 (N_33275,N_32793,N_32640);
nand U33276 (N_33276,N_32540,N_32541);
or U33277 (N_33277,N_32893,N_32804);
nor U33278 (N_33278,N_32847,N_32578);
nor U33279 (N_33279,N_32972,N_32859);
xor U33280 (N_33280,N_32990,N_32912);
xor U33281 (N_33281,N_32756,N_32716);
nor U33282 (N_33282,N_32747,N_32567);
or U33283 (N_33283,N_32750,N_32822);
and U33284 (N_33284,N_32618,N_32592);
and U33285 (N_33285,N_32612,N_32915);
nor U33286 (N_33286,N_32748,N_32916);
and U33287 (N_33287,N_32645,N_32945);
nand U33288 (N_33288,N_32955,N_32881);
or U33289 (N_33289,N_32811,N_32641);
nor U33290 (N_33290,N_32777,N_32647);
nand U33291 (N_33291,N_32948,N_32547);
nand U33292 (N_33292,N_32611,N_32508);
nand U33293 (N_33293,N_32643,N_32645);
nor U33294 (N_33294,N_32980,N_32563);
nand U33295 (N_33295,N_32641,N_32818);
and U33296 (N_33296,N_32809,N_32606);
or U33297 (N_33297,N_32757,N_32712);
and U33298 (N_33298,N_32952,N_32636);
nand U33299 (N_33299,N_32703,N_32860);
and U33300 (N_33300,N_32845,N_32517);
or U33301 (N_33301,N_32725,N_32939);
nand U33302 (N_33302,N_32978,N_32548);
and U33303 (N_33303,N_32659,N_32600);
xor U33304 (N_33304,N_32589,N_32912);
nor U33305 (N_33305,N_32646,N_32690);
xor U33306 (N_33306,N_32704,N_32861);
nor U33307 (N_33307,N_32799,N_32910);
nor U33308 (N_33308,N_32960,N_32838);
nor U33309 (N_33309,N_32514,N_32660);
nor U33310 (N_33310,N_32678,N_32727);
xnor U33311 (N_33311,N_32894,N_32803);
and U33312 (N_33312,N_32792,N_32658);
nor U33313 (N_33313,N_32962,N_32690);
or U33314 (N_33314,N_32699,N_32937);
nor U33315 (N_33315,N_32563,N_32930);
and U33316 (N_33316,N_32933,N_32910);
nand U33317 (N_33317,N_32624,N_32927);
and U33318 (N_33318,N_32738,N_32739);
nor U33319 (N_33319,N_32849,N_32875);
nand U33320 (N_33320,N_32632,N_32855);
nor U33321 (N_33321,N_32551,N_32702);
nand U33322 (N_33322,N_32664,N_32947);
nand U33323 (N_33323,N_32774,N_32582);
nor U33324 (N_33324,N_32873,N_32948);
and U33325 (N_33325,N_32607,N_32603);
nor U33326 (N_33326,N_32831,N_32687);
nor U33327 (N_33327,N_32888,N_32727);
nor U33328 (N_33328,N_32904,N_32738);
and U33329 (N_33329,N_32955,N_32521);
or U33330 (N_33330,N_32877,N_32642);
and U33331 (N_33331,N_32573,N_32738);
nor U33332 (N_33332,N_32585,N_32808);
and U33333 (N_33333,N_32828,N_32992);
nor U33334 (N_33334,N_32567,N_32963);
and U33335 (N_33335,N_32905,N_32676);
or U33336 (N_33336,N_32752,N_32776);
or U33337 (N_33337,N_32721,N_32578);
and U33338 (N_33338,N_32871,N_32726);
nand U33339 (N_33339,N_32899,N_32615);
xnor U33340 (N_33340,N_32611,N_32612);
nor U33341 (N_33341,N_32737,N_32857);
xor U33342 (N_33342,N_32666,N_32723);
or U33343 (N_33343,N_32706,N_32837);
nand U33344 (N_33344,N_32581,N_32910);
or U33345 (N_33345,N_32975,N_32984);
nor U33346 (N_33346,N_32585,N_32985);
nand U33347 (N_33347,N_32663,N_32556);
nand U33348 (N_33348,N_32968,N_32679);
nor U33349 (N_33349,N_32848,N_32777);
nand U33350 (N_33350,N_32694,N_32675);
xnor U33351 (N_33351,N_32710,N_32737);
xnor U33352 (N_33352,N_32674,N_32504);
or U33353 (N_33353,N_32713,N_32938);
xnor U33354 (N_33354,N_32861,N_32839);
xor U33355 (N_33355,N_32924,N_32844);
nor U33356 (N_33356,N_32976,N_32788);
or U33357 (N_33357,N_32937,N_32728);
or U33358 (N_33358,N_32900,N_32962);
or U33359 (N_33359,N_32887,N_32775);
and U33360 (N_33360,N_32869,N_32909);
nand U33361 (N_33361,N_32896,N_32981);
nor U33362 (N_33362,N_32793,N_32795);
nand U33363 (N_33363,N_32999,N_32567);
nand U33364 (N_33364,N_32859,N_32838);
nor U33365 (N_33365,N_32679,N_32824);
nor U33366 (N_33366,N_32721,N_32685);
and U33367 (N_33367,N_32505,N_32805);
or U33368 (N_33368,N_32940,N_32950);
nor U33369 (N_33369,N_32644,N_32713);
or U33370 (N_33370,N_32539,N_32980);
nand U33371 (N_33371,N_32849,N_32722);
nand U33372 (N_33372,N_32954,N_32527);
nand U33373 (N_33373,N_32513,N_32920);
nand U33374 (N_33374,N_32560,N_32690);
or U33375 (N_33375,N_32507,N_32774);
nor U33376 (N_33376,N_32848,N_32705);
nor U33377 (N_33377,N_32565,N_32585);
and U33378 (N_33378,N_32962,N_32598);
or U33379 (N_33379,N_32625,N_32534);
xor U33380 (N_33380,N_32565,N_32600);
and U33381 (N_33381,N_32566,N_32602);
nand U33382 (N_33382,N_32811,N_32642);
nand U33383 (N_33383,N_32740,N_32504);
nand U33384 (N_33384,N_32508,N_32841);
nor U33385 (N_33385,N_32615,N_32987);
and U33386 (N_33386,N_32679,N_32532);
and U33387 (N_33387,N_32649,N_32573);
or U33388 (N_33388,N_32647,N_32747);
nand U33389 (N_33389,N_32882,N_32709);
and U33390 (N_33390,N_32525,N_32972);
nand U33391 (N_33391,N_32628,N_32687);
xor U33392 (N_33392,N_32885,N_32991);
nand U33393 (N_33393,N_32786,N_32665);
and U33394 (N_33394,N_32771,N_32746);
nor U33395 (N_33395,N_32536,N_32718);
nor U33396 (N_33396,N_32640,N_32825);
or U33397 (N_33397,N_32979,N_32676);
and U33398 (N_33398,N_32606,N_32906);
nor U33399 (N_33399,N_32687,N_32996);
or U33400 (N_33400,N_32809,N_32855);
or U33401 (N_33401,N_32945,N_32640);
and U33402 (N_33402,N_32762,N_32687);
and U33403 (N_33403,N_32858,N_32776);
and U33404 (N_33404,N_32995,N_32911);
or U33405 (N_33405,N_32873,N_32706);
or U33406 (N_33406,N_32522,N_32675);
nand U33407 (N_33407,N_32755,N_32761);
or U33408 (N_33408,N_32645,N_32627);
nand U33409 (N_33409,N_32523,N_32797);
nand U33410 (N_33410,N_32573,N_32864);
nor U33411 (N_33411,N_32789,N_32914);
nor U33412 (N_33412,N_32794,N_32930);
or U33413 (N_33413,N_32548,N_32910);
nand U33414 (N_33414,N_32529,N_32567);
nor U33415 (N_33415,N_32526,N_32947);
xor U33416 (N_33416,N_32953,N_32899);
or U33417 (N_33417,N_32841,N_32687);
nor U33418 (N_33418,N_32953,N_32927);
nor U33419 (N_33419,N_32787,N_32770);
and U33420 (N_33420,N_32856,N_32788);
and U33421 (N_33421,N_32900,N_32523);
nand U33422 (N_33422,N_32649,N_32724);
nor U33423 (N_33423,N_32929,N_32683);
nand U33424 (N_33424,N_32794,N_32822);
and U33425 (N_33425,N_32702,N_32900);
nor U33426 (N_33426,N_32654,N_32706);
nand U33427 (N_33427,N_32726,N_32873);
nor U33428 (N_33428,N_32989,N_32573);
nor U33429 (N_33429,N_32752,N_32912);
and U33430 (N_33430,N_32900,N_32530);
and U33431 (N_33431,N_32601,N_32652);
nand U33432 (N_33432,N_32844,N_32906);
nand U33433 (N_33433,N_32555,N_32653);
and U33434 (N_33434,N_32680,N_32660);
xor U33435 (N_33435,N_32965,N_32595);
nand U33436 (N_33436,N_32813,N_32907);
nor U33437 (N_33437,N_32714,N_32774);
nor U33438 (N_33438,N_32932,N_32946);
or U33439 (N_33439,N_32979,N_32574);
nor U33440 (N_33440,N_32806,N_32675);
xnor U33441 (N_33441,N_32633,N_32766);
and U33442 (N_33442,N_32967,N_32840);
and U33443 (N_33443,N_32993,N_32596);
or U33444 (N_33444,N_32937,N_32711);
and U33445 (N_33445,N_32990,N_32779);
nor U33446 (N_33446,N_32508,N_32959);
nand U33447 (N_33447,N_32502,N_32925);
or U33448 (N_33448,N_32789,N_32785);
xnor U33449 (N_33449,N_32892,N_32504);
or U33450 (N_33450,N_32682,N_32651);
or U33451 (N_33451,N_32645,N_32508);
nor U33452 (N_33452,N_32818,N_32763);
nor U33453 (N_33453,N_32645,N_32613);
or U33454 (N_33454,N_32982,N_32991);
and U33455 (N_33455,N_32710,N_32892);
nand U33456 (N_33456,N_32861,N_32823);
nand U33457 (N_33457,N_32510,N_32899);
nand U33458 (N_33458,N_32797,N_32823);
nor U33459 (N_33459,N_32973,N_32950);
and U33460 (N_33460,N_32773,N_32644);
nand U33461 (N_33461,N_32866,N_32553);
or U33462 (N_33462,N_32633,N_32533);
nand U33463 (N_33463,N_32623,N_32987);
nand U33464 (N_33464,N_32532,N_32537);
nor U33465 (N_33465,N_32854,N_32955);
or U33466 (N_33466,N_32557,N_32829);
and U33467 (N_33467,N_32570,N_32507);
or U33468 (N_33468,N_32789,N_32572);
nand U33469 (N_33469,N_32575,N_32795);
nand U33470 (N_33470,N_32987,N_32867);
nor U33471 (N_33471,N_32599,N_32725);
or U33472 (N_33472,N_32594,N_32863);
nand U33473 (N_33473,N_32648,N_32838);
or U33474 (N_33474,N_32922,N_32931);
nand U33475 (N_33475,N_32548,N_32678);
xor U33476 (N_33476,N_32902,N_32714);
and U33477 (N_33477,N_32507,N_32617);
nor U33478 (N_33478,N_32947,N_32593);
nor U33479 (N_33479,N_32857,N_32840);
nand U33480 (N_33480,N_32919,N_32636);
xnor U33481 (N_33481,N_32976,N_32702);
nor U33482 (N_33482,N_32579,N_32754);
nand U33483 (N_33483,N_32590,N_32607);
nor U33484 (N_33484,N_32907,N_32534);
nor U33485 (N_33485,N_32722,N_32753);
nor U33486 (N_33486,N_32937,N_32659);
nand U33487 (N_33487,N_32863,N_32814);
and U33488 (N_33488,N_32704,N_32767);
or U33489 (N_33489,N_32952,N_32796);
or U33490 (N_33490,N_32523,N_32540);
nor U33491 (N_33491,N_32776,N_32839);
nand U33492 (N_33492,N_32792,N_32867);
nor U33493 (N_33493,N_32858,N_32555);
nor U33494 (N_33494,N_32664,N_32579);
nor U33495 (N_33495,N_32743,N_32756);
or U33496 (N_33496,N_32600,N_32603);
or U33497 (N_33497,N_32695,N_32582);
nand U33498 (N_33498,N_32880,N_32625);
or U33499 (N_33499,N_32698,N_32605);
or U33500 (N_33500,N_33272,N_33481);
or U33501 (N_33501,N_33038,N_33154);
nand U33502 (N_33502,N_33152,N_33412);
or U33503 (N_33503,N_33078,N_33309);
nor U33504 (N_33504,N_33146,N_33379);
nand U33505 (N_33505,N_33418,N_33112);
nand U33506 (N_33506,N_33307,N_33016);
or U33507 (N_33507,N_33298,N_33422);
or U33508 (N_33508,N_33389,N_33092);
and U33509 (N_33509,N_33275,N_33181);
and U33510 (N_33510,N_33281,N_33252);
nand U33511 (N_33511,N_33297,N_33363);
and U33512 (N_33512,N_33405,N_33101);
nand U33513 (N_33513,N_33273,N_33163);
nor U33514 (N_33514,N_33324,N_33359);
or U33515 (N_33515,N_33185,N_33180);
and U33516 (N_33516,N_33401,N_33436);
nand U33517 (N_33517,N_33126,N_33372);
or U33518 (N_33518,N_33010,N_33404);
and U33519 (N_33519,N_33202,N_33391);
nand U33520 (N_33520,N_33117,N_33216);
nor U33521 (N_33521,N_33162,N_33168);
or U33522 (N_33522,N_33308,N_33222);
nor U33523 (N_33523,N_33393,N_33083);
nor U33524 (N_33524,N_33094,N_33084);
and U33525 (N_33525,N_33258,N_33348);
and U33526 (N_33526,N_33043,N_33477);
xor U33527 (N_33527,N_33350,N_33210);
nand U33528 (N_33528,N_33194,N_33417);
nor U33529 (N_33529,N_33499,N_33476);
and U33530 (N_33530,N_33110,N_33342);
nor U33531 (N_33531,N_33454,N_33019);
nor U33532 (N_33532,N_33322,N_33314);
or U33533 (N_33533,N_33229,N_33142);
nor U33534 (N_33534,N_33471,N_33075);
xor U33535 (N_33535,N_33257,N_33030);
nor U33536 (N_33536,N_33265,N_33459);
nor U33537 (N_33537,N_33150,N_33289);
nor U33538 (N_33538,N_33279,N_33005);
nand U33539 (N_33539,N_33259,N_33169);
nor U33540 (N_33540,N_33134,N_33247);
or U33541 (N_33541,N_33042,N_33285);
and U33542 (N_33542,N_33218,N_33356);
and U33543 (N_33543,N_33413,N_33173);
nor U33544 (N_33544,N_33012,N_33123);
xor U33545 (N_33545,N_33014,N_33208);
and U33546 (N_33546,N_33450,N_33211);
and U33547 (N_33547,N_33122,N_33377);
or U33548 (N_33548,N_33028,N_33193);
xnor U33549 (N_33549,N_33018,N_33400);
and U33550 (N_33550,N_33430,N_33473);
nor U33551 (N_33551,N_33296,N_33396);
nand U33552 (N_33552,N_33423,N_33260);
or U33553 (N_33553,N_33214,N_33468);
and U33554 (N_33554,N_33330,N_33474);
nor U33555 (N_33555,N_33431,N_33428);
and U33556 (N_33556,N_33219,N_33097);
and U33557 (N_33557,N_33161,N_33306);
and U33558 (N_33558,N_33262,N_33147);
nor U33559 (N_33559,N_33192,N_33266);
nand U33560 (N_33560,N_33250,N_33299);
nor U33561 (N_33561,N_33230,N_33354);
nor U33562 (N_33562,N_33015,N_33489);
xor U33563 (N_33563,N_33371,N_33165);
nor U33564 (N_33564,N_33105,N_33292);
nand U33565 (N_33565,N_33199,N_33243);
and U33566 (N_33566,N_33261,N_33357);
or U33567 (N_33567,N_33201,N_33321);
and U33568 (N_33568,N_33407,N_33191);
nand U33569 (N_33569,N_33268,N_33382);
and U33570 (N_33570,N_33061,N_33461);
or U33571 (N_33571,N_33066,N_33234);
xor U33572 (N_33572,N_33031,N_33291);
nor U33573 (N_33573,N_33411,N_33233);
and U33574 (N_33574,N_33145,N_33434);
and U33575 (N_33575,N_33249,N_33323);
and U33576 (N_33576,N_33280,N_33100);
nand U33577 (N_33577,N_33335,N_33020);
or U33578 (N_33578,N_33264,N_33485);
nor U33579 (N_33579,N_33334,N_33060);
or U33580 (N_33580,N_33288,N_33133);
nand U33581 (N_33581,N_33093,N_33119);
nand U33582 (N_33582,N_33277,N_33046);
nor U33583 (N_33583,N_33344,N_33302);
nand U33584 (N_33584,N_33072,N_33036);
nor U33585 (N_33585,N_33044,N_33059);
and U33586 (N_33586,N_33300,N_33429);
or U33587 (N_33587,N_33080,N_33108);
or U33588 (N_33588,N_33140,N_33338);
or U33589 (N_33589,N_33183,N_33220);
nor U33590 (N_33590,N_33365,N_33057);
nand U33591 (N_33591,N_33231,N_33496);
nand U33592 (N_33592,N_33443,N_33009);
or U33593 (N_33593,N_33386,N_33148);
nand U33594 (N_33594,N_33164,N_33002);
nor U33595 (N_33595,N_33131,N_33053);
or U33596 (N_33596,N_33432,N_33227);
and U33597 (N_33597,N_33244,N_33099);
xor U33598 (N_33598,N_33033,N_33158);
and U33599 (N_33599,N_33421,N_33346);
nor U33600 (N_33600,N_33236,N_33052);
nor U33601 (N_33601,N_33349,N_33017);
or U33602 (N_33602,N_33384,N_33113);
and U33603 (N_33603,N_33156,N_33465);
or U33604 (N_33604,N_33364,N_33064);
or U33605 (N_33605,N_33424,N_33114);
or U33606 (N_33606,N_33301,N_33392);
xnor U33607 (N_33607,N_33118,N_33182);
nand U33608 (N_33608,N_33077,N_33427);
nor U33609 (N_33609,N_33318,N_33171);
nor U33610 (N_33610,N_33143,N_33151);
and U33611 (N_33611,N_33253,N_33337);
nand U33612 (N_33612,N_33425,N_33209);
and U33613 (N_33613,N_33339,N_33287);
nand U33614 (N_33614,N_33091,N_33245);
nand U33615 (N_33615,N_33495,N_33029);
xnor U33616 (N_33616,N_33284,N_33482);
and U33617 (N_33617,N_33196,N_33035);
or U33618 (N_33618,N_33374,N_33469);
xnor U33619 (N_33619,N_33343,N_33098);
nor U33620 (N_33620,N_33013,N_33204);
nand U33621 (N_33621,N_33466,N_33089);
or U33622 (N_33622,N_33488,N_33303);
or U33623 (N_33623,N_33203,N_33132);
or U33624 (N_33624,N_33149,N_33449);
nor U33625 (N_33625,N_33341,N_33115);
nor U33626 (N_33626,N_33256,N_33437);
or U33627 (N_33627,N_33007,N_33478);
nor U33628 (N_33628,N_33049,N_33483);
nor U33629 (N_33629,N_33305,N_33088);
and U33630 (N_33630,N_33027,N_33087);
and U33631 (N_33631,N_33025,N_33095);
nor U33632 (N_33632,N_33130,N_33074);
or U33633 (N_33633,N_33063,N_33408);
nor U33634 (N_33634,N_33457,N_33189);
nand U33635 (N_33635,N_33458,N_33024);
xor U33636 (N_33636,N_33237,N_33283);
or U33637 (N_33637,N_33420,N_33167);
or U33638 (N_33638,N_33388,N_33276);
nor U33639 (N_33639,N_33492,N_33001);
nor U33640 (N_33640,N_33021,N_33336);
and U33641 (N_33641,N_33232,N_33472);
nor U33642 (N_33642,N_33082,N_33416);
nand U33643 (N_33643,N_33484,N_33419);
or U33644 (N_33644,N_33463,N_33190);
nand U33645 (N_33645,N_33467,N_33240);
and U33646 (N_33646,N_33228,N_33355);
and U33647 (N_33647,N_33317,N_33267);
nand U33648 (N_33648,N_33447,N_33373);
nand U33649 (N_33649,N_33340,N_33414);
and U33650 (N_33650,N_33206,N_33294);
xnor U33651 (N_33651,N_33102,N_33313);
and U33652 (N_33652,N_33332,N_33041);
or U33653 (N_33653,N_33248,N_33109);
or U33654 (N_33654,N_33310,N_33226);
nand U33655 (N_33655,N_33159,N_33380);
or U33656 (N_33656,N_33006,N_33076);
nor U33657 (N_33657,N_33069,N_33406);
and U33658 (N_33658,N_33116,N_33464);
nor U33659 (N_33659,N_33205,N_33022);
nor U33660 (N_33660,N_33435,N_33178);
xnor U33661 (N_33661,N_33103,N_33000);
or U33662 (N_33662,N_33451,N_33155);
and U33663 (N_33663,N_33086,N_33304);
or U33664 (N_33664,N_33225,N_33085);
nand U33665 (N_33665,N_33125,N_33070);
nor U33666 (N_33666,N_33129,N_33139);
xor U33667 (N_33667,N_33370,N_33456);
or U33668 (N_33668,N_33312,N_33058);
or U33669 (N_33669,N_33290,N_33120);
or U33670 (N_33670,N_33316,N_33480);
and U33671 (N_33671,N_33184,N_33254);
and U33672 (N_33672,N_33215,N_33366);
and U33673 (N_33673,N_33319,N_33135);
nor U33674 (N_33674,N_33269,N_33186);
xor U33675 (N_33675,N_33455,N_33221);
and U33676 (N_33676,N_33270,N_33040);
or U33677 (N_33677,N_33172,N_33198);
nand U33678 (N_33678,N_33263,N_33497);
nand U33679 (N_33679,N_33278,N_33107);
or U33680 (N_33680,N_33003,N_33399);
and U33681 (N_33681,N_33136,N_33071);
nand U33682 (N_33682,N_33111,N_33498);
or U33683 (N_33683,N_33376,N_33039);
and U33684 (N_33684,N_33068,N_33462);
nor U33685 (N_33685,N_33241,N_33438);
nand U33686 (N_33686,N_33460,N_33056);
and U33687 (N_33687,N_33157,N_33179);
nand U33688 (N_33688,N_33446,N_33493);
and U33689 (N_33689,N_33491,N_33032);
or U33690 (N_33690,N_33175,N_33368);
nor U33691 (N_33691,N_33274,N_33286);
nor U33692 (N_33692,N_33315,N_33200);
and U33693 (N_33693,N_33442,N_33403);
nor U33694 (N_33694,N_33433,N_33328);
nand U33695 (N_33695,N_33255,N_33195);
or U33696 (N_33696,N_33353,N_33475);
or U33697 (N_33697,N_33367,N_33397);
or U33698 (N_33698,N_33352,N_33235);
and U33699 (N_33699,N_33378,N_33479);
nor U33700 (N_33700,N_33008,N_33239);
or U33701 (N_33701,N_33360,N_33034);
or U33702 (N_33702,N_33141,N_33320);
xor U33703 (N_33703,N_33048,N_33213);
xnor U33704 (N_33704,N_33090,N_33486);
nor U33705 (N_33705,N_33137,N_33188);
nand U33706 (N_33706,N_33079,N_33383);
and U33707 (N_33707,N_33050,N_33047);
or U33708 (N_33708,N_33453,N_33490);
or U33709 (N_33709,N_33345,N_33104);
nand U33710 (N_33710,N_33452,N_33023);
nand U33711 (N_33711,N_33065,N_33067);
or U33712 (N_33712,N_33166,N_33361);
nand U33713 (N_33713,N_33121,N_33326);
nand U33714 (N_33714,N_33293,N_33004);
or U33715 (N_33715,N_33385,N_33045);
nor U33716 (N_33716,N_33224,N_33212);
or U33717 (N_33717,N_33242,N_33295);
nand U33718 (N_33718,N_33081,N_33426);
nor U33719 (N_33719,N_33441,N_33197);
nand U33720 (N_33720,N_33444,N_33124);
nand U33721 (N_33721,N_33223,N_33448);
and U33722 (N_33722,N_33174,N_33398);
and U33723 (N_33723,N_33409,N_33054);
or U33724 (N_33724,N_33351,N_33402);
and U33725 (N_33725,N_33106,N_33375);
and U33726 (N_33726,N_33144,N_33331);
nand U33727 (N_33727,N_33153,N_33217);
or U33728 (N_33728,N_33440,N_33026);
nand U33729 (N_33729,N_33395,N_33176);
or U33730 (N_33730,N_33487,N_33347);
nand U33731 (N_33731,N_33271,N_33381);
xor U33732 (N_33732,N_33415,N_33062);
and U33733 (N_33733,N_33439,N_33073);
nor U33734 (N_33734,N_33128,N_33390);
nor U33735 (N_33735,N_33037,N_33362);
nor U33736 (N_33736,N_33494,N_33358);
and U33737 (N_33737,N_33410,N_33311);
or U33738 (N_33738,N_33177,N_33394);
nand U33739 (N_33739,N_33387,N_33170);
nor U33740 (N_33740,N_33282,N_33238);
and U33741 (N_33741,N_33207,N_33055);
nand U33742 (N_33742,N_33011,N_33138);
or U33743 (N_33743,N_33127,N_33187);
and U33744 (N_33744,N_33470,N_33445);
nand U33745 (N_33745,N_33325,N_33246);
or U33746 (N_33746,N_33329,N_33160);
nand U33747 (N_33747,N_33251,N_33051);
nor U33748 (N_33748,N_33096,N_33327);
and U33749 (N_33749,N_33369,N_33333);
nor U33750 (N_33750,N_33495,N_33020);
or U33751 (N_33751,N_33483,N_33309);
and U33752 (N_33752,N_33468,N_33112);
nand U33753 (N_33753,N_33432,N_33205);
or U33754 (N_33754,N_33246,N_33146);
nor U33755 (N_33755,N_33286,N_33166);
nand U33756 (N_33756,N_33395,N_33213);
nor U33757 (N_33757,N_33016,N_33330);
and U33758 (N_33758,N_33232,N_33344);
xnor U33759 (N_33759,N_33409,N_33488);
xnor U33760 (N_33760,N_33372,N_33313);
and U33761 (N_33761,N_33199,N_33406);
or U33762 (N_33762,N_33375,N_33481);
nor U33763 (N_33763,N_33425,N_33366);
nor U33764 (N_33764,N_33472,N_33399);
nor U33765 (N_33765,N_33411,N_33237);
xnor U33766 (N_33766,N_33128,N_33279);
nor U33767 (N_33767,N_33202,N_33364);
and U33768 (N_33768,N_33161,N_33114);
or U33769 (N_33769,N_33374,N_33360);
and U33770 (N_33770,N_33006,N_33430);
nand U33771 (N_33771,N_33276,N_33005);
and U33772 (N_33772,N_33014,N_33247);
nor U33773 (N_33773,N_33320,N_33113);
nand U33774 (N_33774,N_33319,N_33188);
nor U33775 (N_33775,N_33494,N_33438);
nand U33776 (N_33776,N_33195,N_33431);
and U33777 (N_33777,N_33197,N_33173);
and U33778 (N_33778,N_33440,N_33412);
or U33779 (N_33779,N_33177,N_33276);
xnor U33780 (N_33780,N_33401,N_33183);
or U33781 (N_33781,N_33284,N_33043);
or U33782 (N_33782,N_33116,N_33197);
nor U33783 (N_33783,N_33322,N_33276);
xor U33784 (N_33784,N_33062,N_33090);
xnor U33785 (N_33785,N_33494,N_33184);
nor U33786 (N_33786,N_33450,N_33389);
or U33787 (N_33787,N_33376,N_33395);
or U33788 (N_33788,N_33079,N_33331);
nand U33789 (N_33789,N_33448,N_33301);
xor U33790 (N_33790,N_33130,N_33449);
nand U33791 (N_33791,N_33263,N_33239);
nor U33792 (N_33792,N_33010,N_33445);
or U33793 (N_33793,N_33123,N_33144);
or U33794 (N_33794,N_33321,N_33163);
nand U33795 (N_33795,N_33253,N_33060);
or U33796 (N_33796,N_33020,N_33003);
nor U33797 (N_33797,N_33340,N_33334);
nand U33798 (N_33798,N_33365,N_33079);
xnor U33799 (N_33799,N_33213,N_33469);
and U33800 (N_33800,N_33226,N_33393);
nor U33801 (N_33801,N_33126,N_33002);
and U33802 (N_33802,N_33171,N_33173);
or U33803 (N_33803,N_33382,N_33434);
nor U33804 (N_33804,N_33038,N_33213);
nand U33805 (N_33805,N_33482,N_33238);
or U33806 (N_33806,N_33436,N_33474);
nor U33807 (N_33807,N_33158,N_33194);
nand U33808 (N_33808,N_33159,N_33174);
nor U33809 (N_33809,N_33276,N_33219);
or U33810 (N_33810,N_33195,N_33087);
and U33811 (N_33811,N_33484,N_33454);
nand U33812 (N_33812,N_33262,N_33162);
and U33813 (N_33813,N_33396,N_33375);
nand U33814 (N_33814,N_33121,N_33152);
nand U33815 (N_33815,N_33297,N_33147);
nor U33816 (N_33816,N_33313,N_33015);
nor U33817 (N_33817,N_33102,N_33411);
nor U33818 (N_33818,N_33184,N_33279);
nor U33819 (N_33819,N_33147,N_33098);
nor U33820 (N_33820,N_33023,N_33038);
xnor U33821 (N_33821,N_33373,N_33113);
or U33822 (N_33822,N_33304,N_33213);
or U33823 (N_33823,N_33418,N_33338);
or U33824 (N_33824,N_33022,N_33179);
nor U33825 (N_33825,N_33234,N_33212);
or U33826 (N_33826,N_33277,N_33476);
or U33827 (N_33827,N_33103,N_33313);
nand U33828 (N_33828,N_33367,N_33306);
or U33829 (N_33829,N_33440,N_33022);
or U33830 (N_33830,N_33374,N_33483);
nor U33831 (N_33831,N_33212,N_33096);
or U33832 (N_33832,N_33137,N_33044);
xnor U33833 (N_33833,N_33389,N_33312);
or U33834 (N_33834,N_33240,N_33118);
or U33835 (N_33835,N_33191,N_33386);
or U33836 (N_33836,N_33455,N_33429);
and U33837 (N_33837,N_33180,N_33350);
and U33838 (N_33838,N_33020,N_33311);
nor U33839 (N_33839,N_33158,N_33228);
nor U33840 (N_33840,N_33236,N_33004);
and U33841 (N_33841,N_33294,N_33115);
or U33842 (N_33842,N_33082,N_33280);
nand U33843 (N_33843,N_33290,N_33387);
nor U33844 (N_33844,N_33462,N_33216);
nor U33845 (N_33845,N_33101,N_33275);
nand U33846 (N_33846,N_33457,N_33207);
nor U33847 (N_33847,N_33019,N_33146);
or U33848 (N_33848,N_33244,N_33274);
nor U33849 (N_33849,N_33322,N_33027);
xor U33850 (N_33850,N_33051,N_33136);
or U33851 (N_33851,N_33082,N_33423);
and U33852 (N_33852,N_33213,N_33055);
nor U33853 (N_33853,N_33395,N_33190);
nand U33854 (N_33854,N_33243,N_33396);
and U33855 (N_33855,N_33065,N_33114);
nand U33856 (N_33856,N_33305,N_33443);
or U33857 (N_33857,N_33487,N_33013);
nor U33858 (N_33858,N_33418,N_33350);
or U33859 (N_33859,N_33496,N_33385);
or U33860 (N_33860,N_33369,N_33179);
nand U33861 (N_33861,N_33472,N_33080);
nand U33862 (N_33862,N_33000,N_33493);
nor U33863 (N_33863,N_33031,N_33365);
xor U33864 (N_33864,N_33251,N_33255);
and U33865 (N_33865,N_33198,N_33360);
and U33866 (N_33866,N_33279,N_33150);
and U33867 (N_33867,N_33165,N_33235);
or U33868 (N_33868,N_33427,N_33407);
nand U33869 (N_33869,N_33452,N_33333);
xor U33870 (N_33870,N_33252,N_33074);
nor U33871 (N_33871,N_33210,N_33375);
xnor U33872 (N_33872,N_33486,N_33421);
or U33873 (N_33873,N_33476,N_33059);
and U33874 (N_33874,N_33238,N_33333);
nor U33875 (N_33875,N_33217,N_33167);
nor U33876 (N_33876,N_33071,N_33152);
nor U33877 (N_33877,N_33143,N_33409);
and U33878 (N_33878,N_33082,N_33120);
and U33879 (N_33879,N_33041,N_33438);
and U33880 (N_33880,N_33386,N_33347);
nand U33881 (N_33881,N_33119,N_33190);
xnor U33882 (N_33882,N_33361,N_33406);
and U33883 (N_33883,N_33370,N_33109);
or U33884 (N_33884,N_33496,N_33178);
and U33885 (N_33885,N_33065,N_33051);
or U33886 (N_33886,N_33347,N_33415);
nand U33887 (N_33887,N_33181,N_33320);
and U33888 (N_33888,N_33314,N_33145);
nand U33889 (N_33889,N_33121,N_33479);
or U33890 (N_33890,N_33056,N_33192);
nor U33891 (N_33891,N_33303,N_33101);
nand U33892 (N_33892,N_33060,N_33117);
nor U33893 (N_33893,N_33257,N_33277);
nand U33894 (N_33894,N_33180,N_33356);
or U33895 (N_33895,N_33308,N_33080);
nor U33896 (N_33896,N_33129,N_33055);
and U33897 (N_33897,N_33168,N_33339);
and U33898 (N_33898,N_33467,N_33208);
and U33899 (N_33899,N_33471,N_33310);
or U33900 (N_33900,N_33301,N_33185);
nand U33901 (N_33901,N_33496,N_33179);
or U33902 (N_33902,N_33395,N_33018);
nor U33903 (N_33903,N_33272,N_33253);
xnor U33904 (N_33904,N_33263,N_33129);
nor U33905 (N_33905,N_33314,N_33446);
nand U33906 (N_33906,N_33442,N_33231);
nand U33907 (N_33907,N_33364,N_33014);
and U33908 (N_33908,N_33444,N_33190);
and U33909 (N_33909,N_33294,N_33328);
nand U33910 (N_33910,N_33354,N_33268);
nand U33911 (N_33911,N_33391,N_33228);
nor U33912 (N_33912,N_33293,N_33182);
nor U33913 (N_33913,N_33348,N_33193);
or U33914 (N_33914,N_33016,N_33411);
or U33915 (N_33915,N_33007,N_33217);
xor U33916 (N_33916,N_33459,N_33103);
nor U33917 (N_33917,N_33368,N_33116);
and U33918 (N_33918,N_33054,N_33273);
or U33919 (N_33919,N_33213,N_33082);
or U33920 (N_33920,N_33499,N_33036);
nand U33921 (N_33921,N_33228,N_33265);
or U33922 (N_33922,N_33252,N_33467);
and U33923 (N_33923,N_33340,N_33188);
or U33924 (N_33924,N_33145,N_33382);
or U33925 (N_33925,N_33040,N_33302);
nor U33926 (N_33926,N_33437,N_33069);
and U33927 (N_33927,N_33326,N_33011);
nand U33928 (N_33928,N_33326,N_33276);
or U33929 (N_33929,N_33039,N_33238);
nor U33930 (N_33930,N_33017,N_33181);
or U33931 (N_33931,N_33132,N_33041);
nor U33932 (N_33932,N_33271,N_33043);
nand U33933 (N_33933,N_33015,N_33151);
and U33934 (N_33934,N_33283,N_33071);
nor U33935 (N_33935,N_33349,N_33348);
nor U33936 (N_33936,N_33229,N_33086);
and U33937 (N_33937,N_33170,N_33250);
nor U33938 (N_33938,N_33236,N_33025);
or U33939 (N_33939,N_33067,N_33463);
nor U33940 (N_33940,N_33375,N_33330);
nand U33941 (N_33941,N_33293,N_33062);
nor U33942 (N_33942,N_33368,N_33263);
nand U33943 (N_33943,N_33451,N_33122);
and U33944 (N_33944,N_33136,N_33110);
and U33945 (N_33945,N_33376,N_33111);
or U33946 (N_33946,N_33407,N_33214);
nand U33947 (N_33947,N_33147,N_33203);
nor U33948 (N_33948,N_33098,N_33240);
xor U33949 (N_33949,N_33326,N_33231);
nor U33950 (N_33950,N_33320,N_33032);
nor U33951 (N_33951,N_33099,N_33247);
or U33952 (N_33952,N_33254,N_33432);
nor U33953 (N_33953,N_33365,N_33203);
nor U33954 (N_33954,N_33257,N_33054);
xor U33955 (N_33955,N_33289,N_33016);
or U33956 (N_33956,N_33396,N_33330);
nand U33957 (N_33957,N_33240,N_33208);
or U33958 (N_33958,N_33065,N_33007);
nand U33959 (N_33959,N_33365,N_33485);
nand U33960 (N_33960,N_33105,N_33360);
nor U33961 (N_33961,N_33314,N_33091);
xor U33962 (N_33962,N_33169,N_33081);
and U33963 (N_33963,N_33425,N_33481);
and U33964 (N_33964,N_33052,N_33143);
nand U33965 (N_33965,N_33004,N_33102);
nor U33966 (N_33966,N_33011,N_33195);
nand U33967 (N_33967,N_33131,N_33103);
and U33968 (N_33968,N_33124,N_33225);
or U33969 (N_33969,N_33361,N_33327);
and U33970 (N_33970,N_33340,N_33129);
nand U33971 (N_33971,N_33484,N_33271);
nor U33972 (N_33972,N_33473,N_33384);
xor U33973 (N_33973,N_33218,N_33208);
xor U33974 (N_33974,N_33198,N_33065);
or U33975 (N_33975,N_33146,N_33388);
nand U33976 (N_33976,N_33156,N_33103);
and U33977 (N_33977,N_33083,N_33201);
nor U33978 (N_33978,N_33102,N_33186);
or U33979 (N_33979,N_33324,N_33223);
nor U33980 (N_33980,N_33225,N_33140);
and U33981 (N_33981,N_33271,N_33080);
or U33982 (N_33982,N_33140,N_33205);
nor U33983 (N_33983,N_33032,N_33122);
or U33984 (N_33984,N_33092,N_33424);
nor U33985 (N_33985,N_33286,N_33175);
or U33986 (N_33986,N_33168,N_33366);
nand U33987 (N_33987,N_33102,N_33249);
and U33988 (N_33988,N_33312,N_33477);
nand U33989 (N_33989,N_33436,N_33109);
and U33990 (N_33990,N_33252,N_33291);
and U33991 (N_33991,N_33132,N_33070);
and U33992 (N_33992,N_33347,N_33234);
nor U33993 (N_33993,N_33181,N_33151);
nor U33994 (N_33994,N_33295,N_33355);
and U33995 (N_33995,N_33276,N_33094);
nor U33996 (N_33996,N_33473,N_33337);
nor U33997 (N_33997,N_33197,N_33274);
nor U33998 (N_33998,N_33293,N_33307);
nor U33999 (N_33999,N_33471,N_33217);
and U34000 (N_34000,N_33661,N_33639);
and U34001 (N_34001,N_33568,N_33987);
nor U34002 (N_34002,N_33957,N_33986);
nand U34003 (N_34003,N_33556,N_33577);
or U34004 (N_34004,N_33635,N_33591);
nor U34005 (N_34005,N_33849,N_33921);
and U34006 (N_34006,N_33904,N_33959);
or U34007 (N_34007,N_33745,N_33694);
nor U34008 (N_34008,N_33695,N_33737);
nand U34009 (N_34009,N_33867,N_33801);
xnor U34010 (N_34010,N_33804,N_33792);
nor U34011 (N_34011,N_33637,N_33561);
and U34012 (N_34012,N_33786,N_33946);
nor U34013 (N_34013,N_33732,N_33559);
and U34014 (N_34014,N_33582,N_33671);
nor U34015 (N_34015,N_33859,N_33852);
or U34016 (N_34016,N_33756,N_33779);
and U34017 (N_34017,N_33798,N_33578);
and U34018 (N_34018,N_33612,N_33597);
nand U34019 (N_34019,N_33564,N_33646);
or U34020 (N_34020,N_33660,N_33830);
nor U34021 (N_34021,N_33731,N_33656);
nand U34022 (N_34022,N_33836,N_33738);
nor U34023 (N_34023,N_33647,N_33901);
and U34024 (N_34024,N_33598,N_33596);
nor U34025 (N_34025,N_33817,N_33933);
nand U34026 (N_34026,N_33811,N_33932);
nand U34027 (N_34027,N_33668,N_33523);
or U34028 (N_34028,N_33733,N_33968);
and U34029 (N_34029,N_33951,N_33949);
nand U34030 (N_34030,N_33897,N_33624);
or U34031 (N_34031,N_33814,N_33683);
nand U34032 (N_34032,N_33760,N_33713);
or U34033 (N_34033,N_33799,N_33928);
or U34034 (N_34034,N_33956,N_33751);
nand U34035 (N_34035,N_33815,N_33991);
and U34036 (N_34036,N_33504,N_33877);
or U34037 (N_34037,N_33831,N_33995);
nor U34038 (N_34038,N_33544,N_33664);
and U34039 (N_34039,N_33613,N_33687);
nor U34040 (N_34040,N_33657,N_33906);
or U34041 (N_34041,N_33676,N_33778);
nand U34042 (N_34042,N_33607,N_33746);
nor U34043 (N_34043,N_33808,N_33528);
nor U34044 (N_34044,N_33641,N_33819);
and U34045 (N_34045,N_33510,N_33672);
and U34046 (N_34046,N_33922,N_33684);
or U34047 (N_34047,N_33663,N_33763);
nor U34048 (N_34048,N_33707,N_33574);
or U34049 (N_34049,N_33709,N_33856);
and U34050 (N_34050,N_33530,N_33610);
nand U34051 (N_34051,N_33827,N_33615);
or U34052 (N_34052,N_33702,N_33592);
or U34053 (N_34053,N_33710,N_33711);
or U34054 (N_34054,N_33543,N_33513);
xor U34055 (N_34055,N_33809,N_33572);
and U34056 (N_34056,N_33525,N_33547);
nand U34057 (N_34057,N_33651,N_33990);
xor U34058 (N_34058,N_33963,N_33998);
and U34059 (N_34059,N_33820,N_33908);
nor U34060 (N_34060,N_33649,N_33652);
nor U34061 (N_34061,N_33782,N_33653);
xnor U34062 (N_34062,N_33873,N_33757);
nor U34063 (N_34063,N_33674,N_33871);
nor U34064 (N_34064,N_33557,N_33680);
nor U34065 (N_34065,N_33717,N_33911);
and U34066 (N_34066,N_33627,N_33948);
nand U34067 (N_34067,N_33854,N_33862);
nand U34068 (N_34068,N_33725,N_33805);
nor U34069 (N_34069,N_33935,N_33728);
nand U34070 (N_34070,N_33699,N_33993);
nor U34071 (N_34071,N_33883,N_33984);
or U34072 (N_34072,N_33693,N_33669);
or U34073 (N_34073,N_33758,N_33500);
nor U34074 (N_34074,N_33881,N_33531);
nor U34075 (N_34075,N_33917,N_33878);
and U34076 (N_34076,N_33560,N_33795);
nand U34077 (N_34077,N_33807,N_33580);
and U34078 (N_34078,N_33762,N_33611);
nand U34079 (N_34079,N_33551,N_33952);
and U34080 (N_34080,N_33910,N_33983);
or U34081 (N_34081,N_33902,N_33979);
xnor U34082 (N_34082,N_33539,N_33512);
nand U34083 (N_34083,N_33519,N_33631);
nor U34084 (N_34084,N_33973,N_33994);
nor U34085 (N_34085,N_33934,N_33643);
or U34086 (N_34086,N_33810,N_33761);
and U34087 (N_34087,N_33718,N_33834);
or U34088 (N_34088,N_33744,N_33617);
xnor U34089 (N_34089,N_33835,N_33675);
or U34090 (N_34090,N_33923,N_33784);
nand U34091 (N_34091,N_33593,N_33654);
nor U34092 (N_34092,N_33570,N_33723);
nor U34093 (N_34093,N_33588,N_33925);
nand U34094 (N_34094,N_33868,N_33650);
nand U34095 (N_34095,N_33503,N_33941);
and U34096 (N_34096,N_33636,N_33940);
nand U34097 (N_34097,N_33860,N_33909);
and U34098 (N_34098,N_33748,N_33939);
xor U34099 (N_34099,N_33621,N_33843);
nor U34100 (N_34100,N_33943,N_33685);
and U34101 (N_34101,N_33887,N_33703);
or U34102 (N_34102,N_33541,N_33715);
nand U34103 (N_34103,N_33833,N_33599);
and U34104 (N_34104,N_33945,N_33700);
or U34105 (N_34105,N_33749,N_33955);
nor U34106 (N_34106,N_33623,N_33806);
nor U34107 (N_34107,N_33975,N_33704);
nand U34108 (N_34108,N_33775,N_33882);
and U34109 (N_34109,N_33538,N_33851);
or U34110 (N_34110,N_33886,N_33648);
nor U34111 (N_34111,N_33858,N_33579);
nor U34112 (N_34112,N_33754,N_33619);
nand U34113 (N_34113,N_33888,N_33938);
xor U34114 (N_34114,N_33961,N_33774);
nand U34115 (N_34115,N_33644,N_33770);
nor U34116 (N_34116,N_33900,N_33507);
and U34117 (N_34117,N_33581,N_33616);
or U34118 (N_34118,N_33781,N_33918);
nor U34119 (N_34119,N_33947,N_33665);
xnor U34120 (N_34120,N_33874,N_33594);
or U34121 (N_34121,N_33773,N_33569);
and U34122 (N_34122,N_33790,N_33855);
and U34123 (N_34123,N_33772,N_33903);
nand U34124 (N_34124,N_33502,N_33662);
or U34125 (N_34125,N_33802,N_33822);
and U34126 (N_34126,N_33629,N_33850);
or U34127 (N_34127,N_33527,N_33585);
or U34128 (N_34128,N_33666,N_33840);
nand U34129 (N_34129,N_33590,N_33894);
nor U34130 (N_34130,N_33747,N_33803);
or U34131 (N_34131,N_33832,N_33677);
and U34132 (N_34132,N_33965,N_33857);
nand U34133 (N_34133,N_33566,N_33630);
and U34134 (N_34134,N_33678,N_33706);
nor U34135 (N_34135,N_33537,N_33927);
nor U34136 (N_34136,N_33766,N_33863);
or U34137 (N_34137,N_33912,N_33509);
and U34138 (N_34138,N_33866,N_33769);
and U34139 (N_34139,N_33576,N_33587);
and U34140 (N_34140,N_33930,N_33960);
and U34141 (N_34141,N_33896,N_33899);
nand U34142 (N_34142,N_33589,N_33787);
xnor U34143 (N_34143,N_33976,N_33734);
nor U34144 (N_34144,N_33848,N_33869);
and U34145 (N_34145,N_33658,N_33905);
xnor U34146 (N_34146,N_33954,N_33937);
nand U34147 (N_34147,N_33812,N_33988);
nand U34148 (N_34148,N_33601,N_33696);
nor U34149 (N_34149,N_33562,N_33545);
and U34150 (N_34150,N_33893,N_33727);
nor U34151 (N_34151,N_33555,N_33885);
or U34152 (N_34152,N_33518,N_33926);
and U34153 (N_34153,N_33950,N_33853);
and U34154 (N_34154,N_33506,N_33996);
xnor U34155 (N_34155,N_33516,N_33549);
nor U34156 (N_34156,N_33521,N_33608);
or U34157 (N_34157,N_33529,N_33971);
or U34158 (N_34158,N_33755,N_33701);
and U34159 (N_34159,N_33546,N_33841);
nand U34160 (N_34160,N_33604,N_33767);
or U34161 (N_34161,N_33821,N_33978);
or U34162 (N_34162,N_33916,N_33913);
nor U34163 (N_34163,N_33789,N_33768);
or U34164 (N_34164,N_33823,N_33889);
or U34165 (N_34165,N_33826,N_33697);
and U34166 (N_34166,N_33536,N_33907);
nor U34167 (N_34167,N_33837,N_33844);
nor U34168 (N_34168,N_33719,N_33565);
nand U34169 (N_34169,N_33981,N_33708);
xor U34170 (N_34170,N_33534,N_33839);
and U34171 (N_34171,N_33655,N_33729);
nor U34172 (N_34172,N_33997,N_33548);
nand U34173 (N_34173,N_33875,N_33505);
or U34174 (N_34174,N_33989,N_33524);
nand U34175 (N_34175,N_33796,N_33879);
or U34176 (N_34176,N_33673,N_33895);
nor U34177 (N_34177,N_33642,N_33722);
or U34178 (N_34178,N_33550,N_33919);
or U34179 (N_34179,N_33776,N_33793);
or U34180 (N_34180,N_33872,N_33645);
or U34181 (N_34181,N_33972,N_33682);
or U34182 (N_34182,N_33759,N_33845);
nor U34183 (N_34183,N_33563,N_33953);
nor U34184 (N_34184,N_33777,N_33667);
xnor U34185 (N_34185,N_33522,N_33977);
xor U34186 (N_34186,N_33752,N_33533);
or U34187 (N_34187,N_33753,N_33785);
and U34188 (N_34188,N_33780,N_33681);
or U34189 (N_34189,N_33898,N_33892);
nand U34190 (N_34190,N_33740,N_33842);
or U34191 (N_34191,N_33942,N_33962);
nor U34192 (N_34192,N_33861,N_33553);
and U34193 (N_34193,N_33966,N_33816);
and U34194 (N_34194,N_33735,N_33964);
xor U34195 (N_34195,N_33692,N_33724);
nor U34196 (N_34196,N_33794,N_33828);
or U34197 (N_34197,N_33638,N_33931);
nor U34198 (N_34198,N_33765,N_33618);
and U34199 (N_34199,N_33985,N_33967);
nor U34200 (N_34200,N_33813,N_33511);
xor U34201 (N_34201,N_33573,N_33606);
xor U34202 (N_34202,N_33742,N_33532);
and U34203 (N_34203,N_33688,N_33640);
or U34204 (N_34204,N_33632,N_33720);
or U34205 (N_34205,N_33535,N_33891);
xnor U34206 (N_34206,N_33730,N_33824);
and U34207 (N_34207,N_33501,N_33958);
or U34208 (N_34208,N_33721,N_33864);
nand U34209 (N_34209,N_33771,N_33517);
and U34210 (N_34210,N_33791,N_33540);
nor U34211 (N_34211,N_33880,N_33884);
and U34212 (N_34212,N_33865,N_33614);
nor U34213 (N_34213,N_33603,N_33980);
nor U34214 (N_34214,N_33969,N_33670);
nand U34215 (N_34215,N_33690,N_33739);
nor U34216 (N_34216,N_33609,N_33520);
and U34217 (N_34217,N_33554,N_33583);
nor U34218 (N_34218,N_33625,N_33838);
or U34219 (N_34219,N_33929,N_33508);
or U34220 (N_34220,N_33689,N_33783);
and U34221 (N_34221,N_33691,N_33800);
xnor U34222 (N_34222,N_33595,N_33605);
nand U34223 (N_34223,N_33716,N_33712);
nor U34224 (N_34224,N_33714,N_33999);
nand U34225 (N_34225,N_33992,N_33974);
or U34226 (N_34226,N_33633,N_33825);
or U34227 (N_34227,N_33602,N_33558);
nand U34228 (N_34228,N_33847,N_33970);
xor U34229 (N_34229,N_33741,N_33797);
and U34230 (N_34230,N_33846,N_33736);
nor U34231 (N_34231,N_33526,N_33705);
nor U34232 (N_34232,N_33890,N_33622);
nor U34233 (N_34233,N_33634,N_33571);
nand U34234 (N_34234,N_33743,N_33659);
nor U34235 (N_34235,N_33914,N_33818);
and U34236 (N_34236,N_33514,N_33620);
nand U34237 (N_34237,N_33920,N_33764);
nor U34238 (N_34238,N_33552,N_33575);
and U34239 (N_34239,N_33628,N_33542);
or U34240 (N_34240,N_33788,N_33515);
nand U34241 (N_34241,N_33626,N_33876);
or U34242 (N_34242,N_33698,N_33982);
nor U34243 (N_34243,N_33600,N_33936);
nor U34244 (N_34244,N_33870,N_33726);
nand U34245 (N_34245,N_33584,N_33915);
or U34246 (N_34246,N_33679,N_33750);
or U34247 (N_34247,N_33686,N_33586);
nand U34248 (N_34248,N_33567,N_33924);
nand U34249 (N_34249,N_33829,N_33944);
xnor U34250 (N_34250,N_33770,N_33508);
nand U34251 (N_34251,N_33776,N_33732);
or U34252 (N_34252,N_33801,N_33846);
xor U34253 (N_34253,N_33719,N_33669);
and U34254 (N_34254,N_33736,N_33955);
xor U34255 (N_34255,N_33827,N_33747);
nor U34256 (N_34256,N_33525,N_33708);
nand U34257 (N_34257,N_33731,N_33588);
nand U34258 (N_34258,N_33711,N_33863);
or U34259 (N_34259,N_33990,N_33770);
nand U34260 (N_34260,N_33583,N_33903);
nand U34261 (N_34261,N_33637,N_33636);
xnor U34262 (N_34262,N_33655,N_33734);
nor U34263 (N_34263,N_33957,N_33881);
and U34264 (N_34264,N_33707,N_33871);
nand U34265 (N_34265,N_33601,N_33855);
or U34266 (N_34266,N_33865,N_33547);
nor U34267 (N_34267,N_33902,N_33796);
and U34268 (N_34268,N_33800,N_33781);
nor U34269 (N_34269,N_33520,N_33950);
and U34270 (N_34270,N_33991,N_33524);
and U34271 (N_34271,N_33579,N_33866);
or U34272 (N_34272,N_33514,N_33536);
nand U34273 (N_34273,N_33937,N_33555);
xor U34274 (N_34274,N_33768,N_33986);
and U34275 (N_34275,N_33604,N_33645);
xnor U34276 (N_34276,N_33820,N_33809);
nand U34277 (N_34277,N_33805,N_33830);
or U34278 (N_34278,N_33513,N_33641);
and U34279 (N_34279,N_33747,N_33554);
or U34280 (N_34280,N_33516,N_33669);
nor U34281 (N_34281,N_33718,N_33633);
and U34282 (N_34282,N_33746,N_33999);
or U34283 (N_34283,N_33525,N_33510);
or U34284 (N_34284,N_33994,N_33786);
nor U34285 (N_34285,N_33828,N_33680);
and U34286 (N_34286,N_33561,N_33834);
or U34287 (N_34287,N_33709,N_33775);
and U34288 (N_34288,N_33907,N_33923);
or U34289 (N_34289,N_33898,N_33949);
xnor U34290 (N_34290,N_33947,N_33613);
nor U34291 (N_34291,N_33789,N_33890);
nand U34292 (N_34292,N_33642,N_33781);
nor U34293 (N_34293,N_33839,N_33601);
or U34294 (N_34294,N_33758,N_33747);
or U34295 (N_34295,N_33921,N_33865);
xor U34296 (N_34296,N_33947,N_33973);
and U34297 (N_34297,N_33574,N_33569);
xor U34298 (N_34298,N_33574,N_33688);
nand U34299 (N_34299,N_33867,N_33773);
and U34300 (N_34300,N_33540,N_33633);
xnor U34301 (N_34301,N_33794,N_33553);
nand U34302 (N_34302,N_33911,N_33824);
nor U34303 (N_34303,N_33848,N_33680);
or U34304 (N_34304,N_33684,N_33744);
nand U34305 (N_34305,N_33613,N_33688);
xnor U34306 (N_34306,N_33846,N_33558);
or U34307 (N_34307,N_33781,N_33846);
and U34308 (N_34308,N_33836,N_33670);
nand U34309 (N_34309,N_33817,N_33578);
or U34310 (N_34310,N_33801,N_33957);
nand U34311 (N_34311,N_33901,N_33785);
and U34312 (N_34312,N_33892,N_33698);
nand U34313 (N_34313,N_33657,N_33578);
xor U34314 (N_34314,N_33783,N_33533);
nand U34315 (N_34315,N_33750,N_33680);
nand U34316 (N_34316,N_33635,N_33649);
nor U34317 (N_34317,N_33509,N_33971);
or U34318 (N_34318,N_33860,N_33897);
and U34319 (N_34319,N_33780,N_33857);
nor U34320 (N_34320,N_33721,N_33826);
and U34321 (N_34321,N_33557,N_33900);
nand U34322 (N_34322,N_33812,N_33712);
nor U34323 (N_34323,N_33732,N_33922);
and U34324 (N_34324,N_33804,N_33808);
or U34325 (N_34325,N_33744,N_33512);
and U34326 (N_34326,N_33641,N_33994);
xnor U34327 (N_34327,N_33856,N_33550);
nand U34328 (N_34328,N_33990,N_33710);
nor U34329 (N_34329,N_33561,N_33619);
nor U34330 (N_34330,N_33548,N_33554);
and U34331 (N_34331,N_33962,N_33953);
or U34332 (N_34332,N_33607,N_33808);
or U34333 (N_34333,N_33672,N_33868);
nand U34334 (N_34334,N_33652,N_33977);
nand U34335 (N_34335,N_33662,N_33752);
or U34336 (N_34336,N_33848,N_33625);
or U34337 (N_34337,N_33669,N_33597);
nand U34338 (N_34338,N_33700,N_33669);
nand U34339 (N_34339,N_33828,N_33818);
or U34340 (N_34340,N_33546,N_33562);
nand U34341 (N_34341,N_33586,N_33547);
or U34342 (N_34342,N_33534,N_33569);
xor U34343 (N_34343,N_33953,N_33608);
or U34344 (N_34344,N_33524,N_33613);
xnor U34345 (N_34345,N_33672,N_33808);
or U34346 (N_34346,N_33608,N_33951);
xor U34347 (N_34347,N_33562,N_33954);
or U34348 (N_34348,N_33619,N_33951);
xor U34349 (N_34349,N_33781,N_33562);
nor U34350 (N_34350,N_33701,N_33641);
nor U34351 (N_34351,N_33530,N_33963);
nor U34352 (N_34352,N_33581,N_33534);
or U34353 (N_34353,N_33789,N_33898);
and U34354 (N_34354,N_33740,N_33501);
and U34355 (N_34355,N_33655,N_33526);
nand U34356 (N_34356,N_33792,N_33889);
and U34357 (N_34357,N_33846,N_33674);
xor U34358 (N_34358,N_33731,N_33578);
or U34359 (N_34359,N_33909,N_33769);
and U34360 (N_34360,N_33853,N_33736);
nand U34361 (N_34361,N_33730,N_33739);
nor U34362 (N_34362,N_33959,N_33912);
and U34363 (N_34363,N_33953,N_33914);
nand U34364 (N_34364,N_33516,N_33961);
nor U34365 (N_34365,N_33773,N_33599);
and U34366 (N_34366,N_33520,N_33607);
nor U34367 (N_34367,N_33705,N_33719);
and U34368 (N_34368,N_33587,N_33724);
nor U34369 (N_34369,N_33733,N_33623);
and U34370 (N_34370,N_33550,N_33570);
nor U34371 (N_34371,N_33772,N_33868);
and U34372 (N_34372,N_33507,N_33595);
nand U34373 (N_34373,N_33770,N_33561);
nor U34374 (N_34374,N_33992,N_33954);
and U34375 (N_34375,N_33918,N_33706);
xor U34376 (N_34376,N_33995,N_33929);
xnor U34377 (N_34377,N_33529,N_33506);
and U34378 (N_34378,N_33683,N_33883);
nor U34379 (N_34379,N_33727,N_33931);
nor U34380 (N_34380,N_33633,N_33830);
nand U34381 (N_34381,N_33881,N_33971);
and U34382 (N_34382,N_33742,N_33538);
nand U34383 (N_34383,N_33662,N_33833);
and U34384 (N_34384,N_33536,N_33619);
and U34385 (N_34385,N_33792,N_33983);
or U34386 (N_34386,N_33822,N_33658);
and U34387 (N_34387,N_33697,N_33554);
and U34388 (N_34388,N_33714,N_33629);
and U34389 (N_34389,N_33915,N_33783);
nor U34390 (N_34390,N_33914,N_33683);
nor U34391 (N_34391,N_33651,N_33781);
nor U34392 (N_34392,N_33551,N_33816);
nand U34393 (N_34393,N_33737,N_33533);
nand U34394 (N_34394,N_33647,N_33676);
and U34395 (N_34395,N_33502,N_33630);
or U34396 (N_34396,N_33751,N_33699);
nor U34397 (N_34397,N_33856,N_33936);
and U34398 (N_34398,N_33767,N_33789);
and U34399 (N_34399,N_33681,N_33852);
nor U34400 (N_34400,N_33545,N_33832);
and U34401 (N_34401,N_33583,N_33800);
nand U34402 (N_34402,N_33943,N_33794);
and U34403 (N_34403,N_33623,N_33783);
nor U34404 (N_34404,N_33675,N_33972);
and U34405 (N_34405,N_33898,N_33649);
nor U34406 (N_34406,N_33903,N_33886);
or U34407 (N_34407,N_33633,N_33622);
nor U34408 (N_34408,N_33571,N_33754);
or U34409 (N_34409,N_33924,N_33774);
and U34410 (N_34410,N_33608,N_33518);
or U34411 (N_34411,N_33547,N_33574);
and U34412 (N_34412,N_33543,N_33974);
or U34413 (N_34413,N_33755,N_33752);
nand U34414 (N_34414,N_33506,N_33655);
nand U34415 (N_34415,N_33536,N_33840);
xor U34416 (N_34416,N_33941,N_33506);
nor U34417 (N_34417,N_33928,N_33827);
nor U34418 (N_34418,N_33813,N_33951);
or U34419 (N_34419,N_33901,N_33855);
nor U34420 (N_34420,N_33716,N_33620);
nor U34421 (N_34421,N_33924,N_33820);
nor U34422 (N_34422,N_33748,N_33830);
nor U34423 (N_34423,N_33718,N_33570);
nor U34424 (N_34424,N_33617,N_33783);
nor U34425 (N_34425,N_33534,N_33772);
nor U34426 (N_34426,N_33609,N_33535);
or U34427 (N_34427,N_33807,N_33619);
nand U34428 (N_34428,N_33671,N_33699);
nor U34429 (N_34429,N_33788,N_33814);
nor U34430 (N_34430,N_33869,N_33836);
xor U34431 (N_34431,N_33792,N_33813);
nand U34432 (N_34432,N_33946,N_33878);
xor U34433 (N_34433,N_33796,N_33719);
or U34434 (N_34434,N_33506,N_33785);
or U34435 (N_34435,N_33811,N_33931);
xnor U34436 (N_34436,N_33622,N_33519);
or U34437 (N_34437,N_33561,N_33782);
or U34438 (N_34438,N_33876,N_33955);
and U34439 (N_34439,N_33837,N_33708);
nor U34440 (N_34440,N_33857,N_33986);
xnor U34441 (N_34441,N_33923,N_33837);
nor U34442 (N_34442,N_33941,N_33970);
and U34443 (N_34443,N_33653,N_33615);
nand U34444 (N_34444,N_33877,N_33959);
nand U34445 (N_34445,N_33828,N_33532);
nor U34446 (N_34446,N_33632,N_33615);
and U34447 (N_34447,N_33763,N_33513);
nand U34448 (N_34448,N_33826,N_33564);
nand U34449 (N_34449,N_33907,N_33722);
and U34450 (N_34450,N_33663,N_33747);
nand U34451 (N_34451,N_33630,N_33801);
and U34452 (N_34452,N_33608,N_33781);
and U34453 (N_34453,N_33831,N_33757);
and U34454 (N_34454,N_33630,N_33704);
nor U34455 (N_34455,N_33512,N_33644);
and U34456 (N_34456,N_33592,N_33807);
nand U34457 (N_34457,N_33713,N_33769);
nand U34458 (N_34458,N_33818,N_33607);
or U34459 (N_34459,N_33686,N_33981);
nor U34460 (N_34460,N_33701,N_33885);
nor U34461 (N_34461,N_33832,N_33982);
nand U34462 (N_34462,N_33897,N_33652);
nand U34463 (N_34463,N_33701,N_33906);
and U34464 (N_34464,N_33976,N_33874);
and U34465 (N_34465,N_33761,N_33631);
and U34466 (N_34466,N_33816,N_33601);
or U34467 (N_34467,N_33609,N_33812);
and U34468 (N_34468,N_33879,N_33940);
nor U34469 (N_34469,N_33827,N_33663);
nand U34470 (N_34470,N_33721,N_33825);
or U34471 (N_34471,N_33881,N_33512);
or U34472 (N_34472,N_33755,N_33531);
or U34473 (N_34473,N_33626,N_33993);
nand U34474 (N_34474,N_33886,N_33706);
and U34475 (N_34475,N_33800,N_33747);
nor U34476 (N_34476,N_33806,N_33991);
or U34477 (N_34477,N_33970,N_33927);
and U34478 (N_34478,N_33531,N_33791);
nor U34479 (N_34479,N_33984,N_33535);
nand U34480 (N_34480,N_33916,N_33784);
and U34481 (N_34481,N_33805,N_33557);
nor U34482 (N_34482,N_33978,N_33953);
or U34483 (N_34483,N_33893,N_33673);
nand U34484 (N_34484,N_33631,N_33561);
xor U34485 (N_34485,N_33688,N_33528);
and U34486 (N_34486,N_33872,N_33510);
and U34487 (N_34487,N_33894,N_33652);
xor U34488 (N_34488,N_33853,N_33711);
and U34489 (N_34489,N_33871,N_33704);
and U34490 (N_34490,N_33605,N_33798);
and U34491 (N_34491,N_33674,N_33630);
or U34492 (N_34492,N_33837,N_33690);
nor U34493 (N_34493,N_33640,N_33511);
or U34494 (N_34494,N_33907,N_33573);
nand U34495 (N_34495,N_33967,N_33756);
or U34496 (N_34496,N_33690,N_33768);
and U34497 (N_34497,N_33901,N_33969);
or U34498 (N_34498,N_33514,N_33887);
nand U34499 (N_34499,N_33649,N_33994);
and U34500 (N_34500,N_34286,N_34225);
and U34501 (N_34501,N_34018,N_34039);
or U34502 (N_34502,N_34396,N_34269);
and U34503 (N_34503,N_34005,N_34118);
or U34504 (N_34504,N_34265,N_34348);
nor U34505 (N_34505,N_34121,N_34357);
or U34506 (N_34506,N_34312,N_34015);
nor U34507 (N_34507,N_34239,N_34026);
nand U34508 (N_34508,N_34494,N_34088);
or U34509 (N_34509,N_34046,N_34110);
nor U34510 (N_34510,N_34421,N_34168);
or U34511 (N_34511,N_34449,N_34413);
nand U34512 (N_34512,N_34107,N_34364);
xor U34513 (N_34513,N_34346,N_34493);
nand U34514 (N_34514,N_34272,N_34343);
nor U34515 (N_34515,N_34479,N_34254);
xor U34516 (N_34516,N_34114,N_34440);
and U34517 (N_34517,N_34474,N_34020);
and U34518 (N_34518,N_34124,N_34125);
and U34519 (N_34519,N_34313,N_34288);
nand U34520 (N_34520,N_34260,N_34289);
or U34521 (N_34521,N_34037,N_34367);
and U34522 (N_34522,N_34459,N_34383);
and U34523 (N_34523,N_34024,N_34098);
nor U34524 (N_34524,N_34056,N_34063);
nand U34525 (N_34525,N_34036,N_34399);
nor U34526 (N_34526,N_34149,N_34170);
and U34527 (N_34527,N_34464,N_34298);
nand U34528 (N_34528,N_34089,N_34495);
nor U34529 (N_34529,N_34200,N_34453);
xor U34530 (N_34530,N_34096,N_34309);
or U34531 (N_34531,N_34277,N_34323);
or U34532 (N_34532,N_34368,N_34404);
or U34533 (N_34533,N_34185,N_34101);
or U34534 (N_34534,N_34009,N_34183);
and U34535 (N_34535,N_34195,N_34403);
or U34536 (N_34536,N_34223,N_34167);
and U34537 (N_34537,N_34190,N_34146);
xnor U34538 (N_34538,N_34245,N_34384);
xnor U34539 (N_34539,N_34405,N_34262);
nand U34540 (N_34540,N_34447,N_34355);
xnor U34541 (N_34541,N_34028,N_34490);
nand U34542 (N_34542,N_34010,N_34377);
or U34543 (N_34543,N_34233,N_34071);
and U34544 (N_34544,N_34428,N_34086);
and U34545 (N_34545,N_34394,N_34406);
xnor U34546 (N_34546,N_34158,N_34485);
xor U34547 (N_34547,N_34261,N_34173);
nand U34548 (N_34548,N_34441,N_34252);
nand U34549 (N_34549,N_34450,N_34317);
nor U34550 (N_34550,N_34475,N_34270);
xnor U34551 (N_34551,N_34235,N_34305);
xor U34552 (N_34552,N_34267,N_34287);
and U34553 (N_34553,N_34029,N_34285);
and U34554 (N_34554,N_34220,N_34231);
and U34555 (N_34555,N_34201,N_34238);
and U34556 (N_34556,N_34359,N_34087);
nand U34557 (N_34557,N_34412,N_34470);
nor U34558 (N_34558,N_34085,N_34194);
or U34559 (N_34559,N_34137,N_34294);
nor U34560 (N_34560,N_34092,N_34148);
or U34561 (N_34561,N_34152,N_34079);
or U34562 (N_34562,N_34478,N_34042);
xor U34563 (N_34563,N_34236,N_34308);
nor U34564 (N_34564,N_34492,N_34103);
or U34565 (N_34565,N_34356,N_34160);
nor U34566 (N_34566,N_34295,N_34419);
xnor U34567 (N_34567,N_34388,N_34488);
nor U34568 (N_34568,N_34402,N_34435);
nand U34569 (N_34569,N_34221,N_34145);
and U34570 (N_34570,N_34438,N_34059);
nand U34571 (N_34571,N_34444,N_34140);
nor U34572 (N_34572,N_34242,N_34400);
nand U34573 (N_34573,N_34090,N_34093);
and U34574 (N_34574,N_34001,N_34136);
and U34575 (N_34575,N_34337,N_34176);
nor U34576 (N_34576,N_34186,N_34328);
or U34577 (N_34577,N_34246,N_34048);
nand U34578 (N_34578,N_34410,N_34210);
nand U34579 (N_34579,N_34393,N_34151);
and U34580 (N_34580,N_34213,N_34351);
nand U34581 (N_34581,N_34360,N_34380);
or U34582 (N_34582,N_34062,N_34131);
or U34583 (N_34583,N_34171,N_34060);
nand U34584 (N_34584,N_34455,N_34011);
or U34585 (N_34585,N_34104,N_34442);
nand U34586 (N_34586,N_34255,N_34016);
nor U34587 (N_34587,N_34325,N_34266);
nand U34588 (N_34588,N_34179,N_34466);
and U34589 (N_34589,N_34240,N_34352);
or U34590 (N_34590,N_34499,N_34358);
or U34591 (N_34591,N_34373,N_34003);
or U34592 (N_34592,N_34301,N_34209);
xor U34593 (N_34593,N_34398,N_34297);
nor U34594 (N_34594,N_34392,N_34248);
or U34595 (N_34595,N_34156,N_34243);
nand U34596 (N_34596,N_34117,N_34461);
and U34597 (N_34597,N_34497,N_34423);
nand U34598 (N_34598,N_34030,N_34211);
nor U34599 (N_34599,N_34049,N_34331);
nand U34600 (N_34600,N_34047,N_34381);
nor U34601 (N_34601,N_34227,N_34468);
nor U34602 (N_34602,N_34203,N_34119);
and U34603 (N_34603,N_34418,N_34083);
nand U34604 (N_34604,N_34465,N_34126);
or U34605 (N_34605,N_34228,N_34143);
or U34606 (N_34606,N_34329,N_34105);
nand U34607 (N_34607,N_34379,N_34256);
nor U34608 (N_34608,N_34006,N_34161);
nor U34609 (N_34609,N_34075,N_34296);
or U34610 (N_34610,N_34031,N_34106);
and U34611 (N_34611,N_34330,N_34004);
and U34612 (N_34612,N_34123,N_34275);
xnor U34613 (N_34613,N_34467,N_34417);
or U34614 (N_34614,N_34451,N_34350);
or U34615 (N_34615,N_34054,N_34202);
and U34616 (N_34616,N_34489,N_34369);
or U34617 (N_34617,N_34385,N_34002);
nand U34618 (N_34618,N_34073,N_34147);
nand U34619 (N_34619,N_34250,N_34065);
nand U34620 (N_34620,N_34244,N_34375);
xnor U34621 (N_34621,N_34322,N_34342);
nor U34622 (N_34622,N_34382,N_34184);
nor U34623 (N_34623,N_34333,N_34276);
nand U34624 (N_34624,N_34182,N_34376);
nand U34625 (N_34625,N_34080,N_34074);
nand U34626 (N_34626,N_34469,N_34477);
nor U34627 (N_34627,N_34045,N_34259);
or U34628 (N_34628,N_34249,N_34290);
and U34629 (N_34629,N_34483,N_34043);
and U34630 (N_34630,N_34061,N_34055);
nand U34631 (N_34631,N_34051,N_34226);
and U34632 (N_34632,N_34353,N_34361);
and U34633 (N_34633,N_34278,N_34332);
nor U34634 (N_34634,N_34021,N_34281);
or U34635 (N_34635,N_34484,N_34439);
or U34636 (N_34636,N_34437,N_34033);
nor U34637 (N_34637,N_34111,N_34133);
nor U34638 (N_34638,N_34197,N_34432);
or U34639 (N_34639,N_34409,N_34099);
and U34640 (N_34640,N_34335,N_34268);
nand U34641 (N_34641,N_34371,N_34094);
nor U34642 (N_34642,N_34035,N_34191);
or U34643 (N_34643,N_34081,N_34053);
xor U34644 (N_34644,N_34273,N_34472);
nand U34645 (N_34645,N_34164,N_34155);
nand U34646 (N_34646,N_34034,N_34012);
nor U34647 (N_34647,N_34189,N_34067);
xor U34648 (N_34648,N_34341,N_34362);
nand U34649 (N_34649,N_34222,N_34247);
nor U34650 (N_34650,N_34116,N_34068);
nand U34651 (N_34651,N_34407,N_34443);
nor U34652 (N_34652,N_34387,N_34175);
nor U34653 (N_34653,N_34072,N_34154);
nand U34654 (N_34654,N_34165,N_34122);
and U34655 (N_34655,N_34416,N_34293);
xor U34656 (N_34656,N_34425,N_34013);
nor U34657 (N_34657,N_34304,N_34199);
xnor U34658 (N_34658,N_34306,N_34138);
and U34659 (N_34659,N_34386,N_34084);
nand U34660 (N_34660,N_34253,N_34095);
nor U34661 (N_34661,N_34232,N_34082);
and U34662 (N_34662,N_34206,N_34354);
or U34663 (N_34663,N_34291,N_34128);
or U34664 (N_34664,N_34480,N_34066);
and U34665 (N_34665,N_34284,N_34041);
nand U34666 (N_34666,N_34311,N_34019);
or U34667 (N_34667,N_34365,N_34415);
or U34668 (N_34668,N_34032,N_34193);
nor U34669 (N_34669,N_34132,N_34395);
xor U34670 (N_34670,N_34198,N_34129);
and U34671 (N_34671,N_34241,N_34141);
nand U34672 (N_34672,N_34336,N_34144);
or U34673 (N_34673,N_34397,N_34205);
nand U34674 (N_34674,N_34378,N_34216);
xnor U34675 (N_34675,N_34109,N_34257);
or U34676 (N_34676,N_34345,N_34052);
or U34677 (N_34677,N_34411,N_34163);
nand U34678 (N_34678,N_34091,N_34264);
xor U34679 (N_34679,N_34169,N_34230);
or U34680 (N_34680,N_34139,N_34481);
nor U34681 (N_34681,N_34120,N_34338);
and U34682 (N_34682,N_34431,N_34251);
nand U34683 (N_34683,N_34401,N_34000);
nand U34684 (N_34684,N_34057,N_34436);
and U34685 (N_34685,N_34460,N_34319);
and U34686 (N_34686,N_34040,N_34282);
or U34687 (N_34687,N_34462,N_34188);
or U34688 (N_34688,N_34487,N_34007);
nor U34689 (N_34689,N_34274,N_34192);
nand U34690 (N_34690,N_34280,N_34370);
and U34691 (N_34691,N_34166,N_34058);
and U34692 (N_34692,N_34344,N_34292);
nand U34693 (N_34693,N_34008,N_34321);
nand U34694 (N_34694,N_34314,N_34130);
xnor U34695 (N_34695,N_34318,N_34363);
and U34696 (N_34696,N_34347,N_34457);
nor U34697 (N_34697,N_34215,N_34196);
or U34698 (N_34698,N_34446,N_34022);
nor U34699 (N_34699,N_34180,N_34070);
nor U34700 (N_34700,N_34429,N_34157);
nand U34701 (N_34701,N_34339,N_34300);
xor U34702 (N_34702,N_34486,N_34374);
nor U34703 (N_34703,N_34476,N_34414);
nand U34704 (N_34704,N_34112,N_34498);
or U34705 (N_34705,N_34204,N_34097);
or U34706 (N_34706,N_34064,N_34324);
or U34707 (N_34707,N_34482,N_34208);
xor U34708 (N_34708,N_34150,N_34433);
or U34709 (N_34709,N_34366,N_34229);
xnor U34710 (N_34710,N_34219,N_34263);
nor U34711 (N_34711,N_34320,N_34408);
nand U34712 (N_34712,N_34217,N_34315);
and U34713 (N_34713,N_34237,N_34113);
or U34714 (N_34714,N_34434,N_34496);
nand U34715 (N_34715,N_34426,N_34224);
and U34716 (N_34716,N_34181,N_34178);
nand U34717 (N_34717,N_34038,N_34372);
nand U34718 (N_34718,N_34271,N_34108);
or U34719 (N_34719,N_34310,N_34214);
or U34720 (N_34720,N_34027,N_34102);
nand U34721 (N_34721,N_34340,N_34044);
and U34722 (N_34722,N_34127,N_34078);
nand U34723 (N_34723,N_34299,N_34177);
or U34724 (N_34724,N_34473,N_34279);
nand U34725 (N_34725,N_34427,N_34076);
nor U34726 (N_34726,N_34187,N_34017);
nand U34727 (N_34727,N_34069,N_34135);
and U34728 (N_34728,N_34430,N_34162);
or U34729 (N_34729,N_34218,N_34115);
nand U34730 (N_34730,N_34454,N_34389);
nand U34731 (N_34731,N_34174,N_34303);
and U34732 (N_34732,N_34234,N_34471);
xor U34733 (N_34733,N_34349,N_34452);
xor U34734 (N_34734,N_34458,N_34326);
or U34735 (N_34735,N_34327,N_34014);
nand U34736 (N_34736,N_34077,N_34390);
nand U34737 (N_34737,N_34172,N_34134);
xor U34738 (N_34738,N_34422,N_34153);
and U34739 (N_34739,N_34302,N_34258);
and U34740 (N_34740,N_34025,N_34334);
xor U34741 (N_34741,N_34391,N_34159);
xnor U34742 (N_34742,N_34207,N_34283);
nand U34743 (N_34743,N_34448,N_34316);
or U34744 (N_34744,N_34424,N_34456);
xor U34745 (N_34745,N_34050,N_34445);
and U34746 (N_34746,N_34307,N_34463);
nor U34747 (N_34747,N_34023,N_34491);
nor U34748 (N_34748,N_34100,N_34420);
or U34749 (N_34749,N_34142,N_34212);
nand U34750 (N_34750,N_34205,N_34210);
or U34751 (N_34751,N_34125,N_34400);
or U34752 (N_34752,N_34420,N_34164);
nor U34753 (N_34753,N_34159,N_34100);
nor U34754 (N_34754,N_34125,N_34191);
or U34755 (N_34755,N_34144,N_34415);
or U34756 (N_34756,N_34165,N_34479);
nor U34757 (N_34757,N_34071,N_34292);
or U34758 (N_34758,N_34055,N_34300);
xnor U34759 (N_34759,N_34373,N_34039);
nand U34760 (N_34760,N_34195,N_34410);
and U34761 (N_34761,N_34217,N_34225);
nor U34762 (N_34762,N_34117,N_34370);
nand U34763 (N_34763,N_34322,N_34327);
nand U34764 (N_34764,N_34412,N_34268);
or U34765 (N_34765,N_34210,N_34056);
xnor U34766 (N_34766,N_34039,N_34341);
nand U34767 (N_34767,N_34004,N_34368);
xor U34768 (N_34768,N_34451,N_34096);
xnor U34769 (N_34769,N_34025,N_34307);
or U34770 (N_34770,N_34438,N_34467);
and U34771 (N_34771,N_34427,N_34007);
nand U34772 (N_34772,N_34391,N_34171);
nor U34773 (N_34773,N_34164,N_34015);
or U34774 (N_34774,N_34481,N_34224);
or U34775 (N_34775,N_34260,N_34027);
and U34776 (N_34776,N_34446,N_34405);
nand U34777 (N_34777,N_34484,N_34471);
or U34778 (N_34778,N_34477,N_34323);
nor U34779 (N_34779,N_34387,N_34410);
and U34780 (N_34780,N_34138,N_34486);
or U34781 (N_34781,N_34166,N_34403);
and U34782 (N_34782,N_34345,N_34143);
nand U34783 (N_34783,N_34034,N_34321);
and U34784 (N_34784,N_34323,N_34417);
nand U34785 (N_34785,N_34161,N_34080);
nand U34786 (N_34786,N_34455,N_34150);
nor U34787 (N_34787,N_34473,N_34138);
or U34788 (N_34788,N_34278,N_34005);
or U34789 (N_34789,N_34427,N_34472);
and U34790 (N_34790,N_34096,N_34028);
and U34791 (N_34791,N_34079,N_34310);
nand U34792 (N_34792,N_34252,N_34151);
xnor U34793 (N_34793,N_34045,N_34360);
nand U34794 (N_34794,N_34055,N_34276);
nand U34795 (N_34795,N_34191,N_34255);
nand U34796 (N_34796,N_34150,N_34358);
nor U34797 (N_34797,N_34175,N_34099);
and U34798 (N_34798,N_34146,N_34051);
and U34799 (N_34799,N_34258,N_34265);
and U34800 (N_34800,N_34201,N_34303);
nand U34801 (N_34801,N_34042,N_34309);
or U34802 (N_34802,N_34116,N_34373);
nand U34803 (N_34803,N_34006,N_34079);
nand U34804 (N_34804,N_34023,N_34004);
nand U34805 (N_34805,N_34233,N_34457);
nand U34806 (N_34806,N_34264,N_34000);
and U34807 (N_34807,N_34466,N_34064);
or U34808 (N_34808,N_34345,N_34072);
nor U34809 (N_34809,N_34439,N_34165);
nand U34810 (N_34810,N_34420,N_34314);
nand U34811 (N_34811,N_34223,N_34426);
nand U34812 (N_34812,N_34496,N_34257);
nor U34813 (N_34813,N_34438,N_34271);
nor U34814 (N_34814,N_34127,N_34432);
nor U34815 (N_34815,N_34236,N_34046);
and U34816 (N_34816,N_34462,N_34427);
nor U34817 (N_34817,N_34300,N_34467);
nand U34818 (N_34818,N_34225,N_34381);
nand U34819 (N_34819,N_34469,N_34348);
nand U34820 (N_34820,N_34296,N_34309);
xor U34821 (N_34821,N_34413,N_34148);
or U34822 (N_34822,N_34322,N_34347);
nand U34823 (N_34823,N_34191,N_34002);
and U34824 (N_34824,N_34426,N_34300);
nand U34825 (N_34825,N_34159,N_34086);
xor U34826 (N_34826,N_34472,N_34424);
and U34827 (N_34827,N_34468,N_34423);
nor U34828 (N_34828,N_34270,N_34055);
nor U34829 (N_34829,N_34448,N_34112);
nor U34830 (N_34830,N_34188,N_34063);
and U34831 (N_34831,N_34225,N_34455);
nand U34832 (N_34832,N_34329,N_34142);
nor U34833 (N_34833,N_34486,N_34029);
or U34834 (N_34834,N_34038,N_34018);
nand U34835 (N_34835,N_34262,N_34113);
and U34836 (N_34836,N_34432,N_34148);
nand U34837 (N_34837,N_34257,N_34081);
nand U34838 (N_34838,N_34236,N_34237);
nor U34839 (N_34839,N_34372,N_34370);
nor U34840 (N_34840,N_34247,N_34237);
nor U34841 (N_34841,N_34318,N_34059);
or U34842 (N_34842,N_34463,N_34320);
nor U34843 (N_34843,N_34249,N_34094);
nor U34844 (N_34844,N_34185,N_34168);
xnor U34845 (N_34845,N_34422,N_34413);
nand U34846 (N_34846,N_34293,N_34349);
and U34847 (N_34847,N_34327,N_34389);
and U34848 (N_34848,N_34491,N_34124);
nand U34849 (N_34849,N_34413,N_34284);
nor U34850 (N_34850,N_34319,N_34294);
or U34851 (N_34851,N_34213,N_34459);
or U34852 (N_34852,N_34240,N_34386);
nand U34853 (N_34853,N_34374,N_34077);
and U34854 (N_34854,N_34075,N_34037);
and U34855 (N_34855,N_34272,N_34002);
and U34856 (N_34856,N_34145,N_34057);
or U34857 (N_34857,N_34090,N_34486);
or U34858 (N_34858,N_34231,N_34166);
or U34859 (N_34859,N_34165,N_34049);
nor U34860 (N_34860,N_34211,N_34302);
or U34861 (N_34861,N_34260,N_34309);
or U34862 (N_34862,N_34169,N_34017);
or U34863 (N_34863,N_34411,N_34432);
nand U34864 (N_34864,N_34051,N_34209);
or U34865 (N_34865,N_34209,N_34391);
and U34866 (N_34866,N_34054,N_34320);
or U34867 (N_34867,N_34291,N_34447);
and U34868 (N_34868,N_34025,N_34283);
and U34869 (N_34869,N_34204,N_34210);
nand U34870 (N_34870,N_34319,N_34075);
or U34871 (N_34871,N_34167,N_34439);
and U34872 (N_34872,N_34218,N_34162);
or U34873 (N_34873,N_34164,N_34480);
xor U34874 (N_34874,N_34100,N_34030);
nor U34875 (N_34875,N_34000,N_34471);
nor U34876 (N_34876,N_34203,N_34356);
nand U34877 (N_34877,N_34484,N_34257);
nand U34878 (N_34878,N_34110,N_34057);
and U34879 (N_34879,N_34460,N_34162);
nor U34880 (N_34880,N_34162,N_34264);
nand U34881 (N_34881,N_34190,N_34332);
or U34882 (N_34882,N_34153,N_34310);
or U34883 (N_34883,N_34166,N_34473);
xnor U34884 (N_34884,N_34104,N_34395);
or U34885 (N_34885,N_34202,N_34356);
nand U34886 (N_34886,N_34176,N_34180);
and U34887 (N_34887,N_34499,N_34464);
and U34888 (N_34888,N_34026,N_34005);
or U34889 (N_34889,N_34409,N_34435);
or U34890 (N_34890,N_34151,N_34200);
nor U34891 (N_34891,N_34099,N_34365);
and U34892 (N_34892,N_34245,N_34101);
or U34893 (N_34893,N_34288,N_34457);
or U34894 (N_34894,N_34208,N_34111);
nor U34895 (N_34895,N_34141,N_34325);
nor U34896 (N_34896,N_34061,N_34458);
and U34897 (N_34897,N_34038,N_34412);
and U34898 (N_34898,N_34372,N_34192);
nor U34899 (N_34899,N_34382,N_34379);
nor U34900 (N_34900,N_34041,N_34439);
and U34901 (N_34901,N_34409,N_34076);
and U34902 (N_34902,N_34215,N_34488);
and U34903 (N_34903,N_34274,N_34356);
and U34904 (N_34904,N_34130,N_34188);
xor U34905 (N_34905,N_34083,N_34130);
nand U34906 (N_34906,N_34307,N_34019);
and U34907 (N_34907,N_34190,N_34205);
nor U34908 (N_34908,N_34182,N_34031);
nor U34909 (N_34909,N_34318,N_34405);
and U34910 (N_34910,N_34295,N_34390);
or U34911 (N_34911,N_34470,N_34198);
xnor U34912 (N_34912,N_34178,N_34096);
nor U34913 (N_34913,N_34380,N_34116);
nand U34914 (N_34914,N_34483,N_34106);
nand U34915 (N_34915,N_34079,N_34067);
nor U34916 (N_34916,N_34393,N_34284);
nand U34917 (N_34917,N_34241,N_34266);
and U34918 (N_34918,N_34024,N_34050);
and U34919 (N_34919,N_34141,N_34363);
and U34920 (N_34920,N_34487,N_34185);
nand U34921 (N_34921,N_34028,N_34453);
nand U34922 (N_34922,N_34439,N_34091);
nor U34923 (N_34923,N_34353,N_34460);
nor U34924 (N_34924,N_34456,N_34301);
xor U34925 (N_34925,N_34127,N_34285);
and U34926 (N_34926,N_34258,N_34128);
or U34927 (N_34927,N_34249,N_34337);
nand U34928 (N_34928,N_34098,N_34300);
or U34929 (N_34929,N_34084,N_34068);
or U34930 (N_34930,N_34038,N_34444);
nand U34931 (N_34931,N_34052,N_34134);
nand U34932 (N_34932,N_34217,N_34168);
xor U34933 (N_34933,N_34391,N_34145);
nand U34934 (N_34934,N_34406,N_34488);
and U34935 (N_34935,N_34034,N_34281);
and U34936 (N_34936,N_34473,N_34211);
nand U34937 (N_34937,N_34108,N_34134);
or U34938 (N_34938,N_34421,N_34329);
or U34939 (N_34939,N_34021,N_34415);
xnor U34940 (N_34940,N_34154,N_34354);
and U34941 (N_34941,N_34164,N_34171);
nand U34942 (N_34942,N_34069,N_34074);
and U34943 (N_34943,N_34115,N_34482);
or U34944 (N_34944,N_34165,N_34119);
nor U34945 (N_34945,N_34241,N_34094);
and U34946 (N_34946,N_34107,N_34270);
and U34947 (N_34947,N_34437,N_34144);
xor U34948 (N_34948,N_34381,N_34414);
nand U34949 (N_34949,N_34458,N_34016);
nand U34950 (N_34950,N_34281,N_34415);
or U34951 (N_34951,N_34262,N_34007);
xnor U34952 (N_34952,N_34366,N_34083);
or U34953 (N_34953,N_34329,N_34215);
nor U34954 (N_34954,N_34245,N_34460);
and U34955 (N_34955,N_34357,N_34431);
or U34956 (N_34956,N_34397,N_34372);
or U34957 (N_34957,N_34160,N_34171);
xor U34958 (N_34958,N_34374,N_34454);
and U34959 (N_34959,N_34160,N_34180);
or U34960 (N_34960,N_34354,N_34317);
xnor U34961 (N_34961,N_34180,N_34164);
or U34962 (N_34962,N_34403,N_34016);
and U34963 (N_34963,N_34177,N_34072);
or U34964 (N_34964,N_34235,N_34035);
or U34965 (N_34965,N_34359,N_34298);
and U34966 (N_34966,N_34195,N_34070);
or U34967 (N_34967,N_34428,N_34178);
or U34968 (N_34968,N_34279,N_34041);
and U34969 (N_34969,N_34082,N_34383);
or U34970 (N_34970,N_34083,N_34012);
nand U34971 (N_34971,N_34300,N_34465);
xnor U34972 (N_34972,N_34294,N_34147);
nor U34973 (N_34973,N_34437,N_34404);
or U34974 (N_34974,N_34381,N_34034);
or U34975 (N_34975,N_34418,N_34453);
and U34976 (N_34976,N_34451,N_34059);
nand U34977 (N_34977,N_34431,N_34287);
nor U34978 (N_34978,N_34477,N_34160);
xnor U34979 (N_34979,N_34159,N_34341);
nor U34980 (N_34980,N_34077,N_34313);
and U34981 (N_34981,N_34208,N_34164);
or U34982 (N_34982,N_34397,N_34365);
xnor U34983 (N_34983,N_34121,N_34397);
nor U34984 (N_34984,N_34202,N_34340);
nand U34985 (N_34985,N_34087,N_34153);
and U34986 (N_34986,N_34200,N_34123);
or U34987 (N_34987,N_34096,N_34091);
nand U34988 (N_34988,N_34201,N_34373);
or U34989 (N_34989,N_34078,N_34270);
nor U34990 (N_34990,N_34314,N_34251);
xor U34991 (N_34991,N_34144,N_34203);
or U34992 (N_34992,N_34359,N_34162);
and U34993 (N_34993,N_34139,N_34162);
nand U34994 (N_34994,N_34166,N_34097);
nand U34995 (N_34995,N_34088,N_34210);
xnor U34996 (N_34996,N_34420,N_34369);
nor U34997 (N_34997,N_34422,N_34070);
xnor U34998 (N_34998,N_34464,N_34495);
nand U34999 (N_34999,N_34255,N_34468);
nand U35000 (N_35000,N_34563,N_34903);
or U35001 (N_35001,N_34800,N_34684);
or U35002 (N_35002,N_34588,N_34523);
nand U35003 (N_35003,N_34815,N_34947);
and U35004 (N_35004,N_34782,N_34937);
xor U35005 (N_35005,N_34678,N_34925);
nor U35006 (N_35006,N_34956,N_34935);
or U35007 (N_35007,N_34944,N_34907);
nand U35008 (N_35008,N_34810,N_34963);
xor U35009 (N_35009,N_34960,N_34735);
xor U35010 (N_35010,N_34856,N_34738);
nor U35011 (N_35011,N_34999,N_34527);
or U35012 (N_35012,N_34559,N_34704);
or U35013 (N_35013,N_34662,N_34982);
and U35014 (N_35014,N_34598,N_34534);
or U35015 (N_35015,N_34505,N_34711);
nor U35016 (N_35016,N_34819,N_34813);
or U35017 (N_35017,N_34546,N_34801);
nand U35018 (N_35018,N_34622,N_34790);
xnor U35019 (N_35019,N_34737,N_34826);
and U35020 (N_35020,N_34605,N_34632);
nor U35021 (N_35021,N_34986,N_34607);
nor U35022 (N_35022,N_34503,N_34770);
and U35023 (N_35023,N_34971,N_34649);
nand U35024 (N_35024,N_34761,N_34663);
nor U35025 (N_35025,N_34660,N_34859);
and U35026 (N_35026,N_34549,N_34570);
and U35027 (N_35027,N_34830,N_34988);
nand U35028 (N_35028,N_34510,N_34927);
or U35029 (N_35029,N_34843,N_34928);
nor U35030 (N_35030,N_34697,N_34825);
or U35031 (N_35031,N_34789,N_34943);
or U35032 (N_35032,N_34541,N_34729);
nor U35033 (N_35033,N_34533,N_34781);
or U35034 (N_35034,N_34899,N_34721);
nand U35035 (N_35035,N_34783,N_34579);
and U35036 (N_35036,N_34981,N_34672);
and U35037 (N_35037,N_34516,N_34525);
and U35038 (N_35038,N_34917,N_34728);
and U35039 (N_35039,N_34998,N_34734);
or U35040 (N_35040,N_34718,N_34809);
nand U35041 (N_35041,N_34773,N_34805);
nor U35042 (N_35042,N_34689,N_34876);
xnor U35043 (N_35043,N_34506,N_34707);
nor U35044 (N_35044,N_34582,N_34572);
xnor U35045 (N_35045,N_34724,N_34987);
and U35046 (N_35046,N_34675,N_34544);
and U35047 (N_35047,N_34817,N_34847);
or U35048 (N_35048,N_34871,N_34958);
and U35049 (N_35049,N_34867,N_34824);
nor U35050 (N_35050,N_34716,N_34554);
xnor U35051 (N_35051,N_34528,N_34698);
and U35052 (N_35052,N_34575,N_34553);
or U35053 (N_35053,N_34633,N_34539);
and U35054 (N_35054,N_34621,N_34974);
or U35055 (N_35055,N_34984,N_34746);
nand U35056 (N_35056,N_34569,N_34644);
xor U35057 (N_35057,N_34901,N_34552);
or U35058 (N_35058,N_34788,N_34518);
nand U35059 (N_35059,N_34545,N_34751);
nor U35060 (N_35060,N_34612,N_34994);
nand U35061 (N_35061,N_34926,N_34640);
nand U35062 (N_35062,N_34769,N_34509);
and U35063 (N_35063,N_34702,N_34708);
nor U35064 (N_35064,N_34855,N_34714);
or U35065 (N_35065,N_34722,N_34645);
nand U35066 (N_35066,N_34993,N_34804);
or U35067 (N_35067,N_34604,N_34831);
xnor U35068 (N_35068,N_34587,N_34693);
and U35069 (N_35069,N_34748,N_34918);
nor U35070 (N_35070,N_34667,N_34564);
xor U35071 (N_35071,N_34688,N_34661);
or U35072 (N_35072,N_34565,N_34583);
or U35073 (N_35073,N_34754,N_34940);
xnor U35074 (N_35074,N_34609,N_34853);
or U35075 (N_35075,N_34566,N_34669);
nand U35076 (N_35076,N_34975,N_34623);
nand U35077 (N_35077,N_34705,N_34823);
nand U35078 (N_35078,N_34652,N_34530);
or U35079 (N_35079,N_34627,N_34578);
and U35080 (N_35080,N_34873,N_34683);
nor U35081 (N_35081,N_34886,N_34765);
or U35082 (N_35082,N_34794,N_34908);
nor U35083 (N_35083,N_34655,N_34514);
and U35084 (N_35084,N_34931,N_34685);
and U35085 (N_35085,N_34548,N_34648);
and U35086 (N_35086,N_34979,N_34513);
nand U35087 (N_35087,N_34610,N_34653);
and U35088 (N_35088,N_34763,N_34691);
and U35089 (N_35089,N_34658,N_34750);
nand U35090 (N_35090,N_34639,N_34512);
nand U35091 (N_35091,N_34555,N_34600);
nor U35092 (N_35092,N_34538,N_34665);
nand U35093 (N_35093,N_34797,N_34628);
or U35094 (N_35094,N_34910,N_34690);
and U35095 (N_35095,N_34571,N_34580);
and U35096 (N_35096,N_34715,N_34573);
nor U35097 (N_35097,N_34758,N_34837);
xnor U35098 (N_35098,N_34786,N_34517);
nor U35099 (N_35099,N_34756,N_34972);
or U35100 (N_35100,N_34619,N_34537);
nor U35101 (N_35101,N_34501,N_34818);
nor U35102 (N_35102,N_34515,N_34779);
nor U35103 (N_35103,N_34923,N_34577);
or U35104 (N_35104,N_34753,N_34919);
xnor U35105 (N_35105,N_34832,N_34835);
and U35106 (N_35106,N_34706,N_34952);
and U35107 (N_35107,N_34865,N_34879);
and U35108 (N_35108,N_34868,N_34858);
nand U35109 (N_35109,N_34803,N_34860);
nor U35110 (N_35110,N_34841,N_34976);
and U35111 (N_35111,N_34504,N_34666);
nor U35112 (N_35112,N_34829,N_34641);
and U35113 (N_35113,N_34955,N_34995);
and U35114 (N_35114,N_34852,N_34590);
xnor U35115 (N_35115,N_34732,N_34887);
nand U35116 (N_35116,N_34681,N_34500);
nor U35117 (N_35117,N_34816,N_34664);
and U35118 (N_35118,N_34922,N_34726);
nor U35119 (N_35119,N_34551,N_34961);
or U35120 (N_35120,N_34740,N_34932);
nand U35121 (N_35121,N_34713,N_34620);
nand U35122 (N_35122,N_34890,N_34814);
xnor U35123 (N_35123,N_34793,N_34921);
xnor U35124 (N_35124,N_34954,N_34507);
and U35125 (N_35125,N_34864,N_34776);
nor U35126 (N_35126,N_34970,N_34616);
and U35127 (N_35127,N_34977,N_34766);
or U35128 (N_35128,N_34840,N_34597);
nand U35129 (N_35129,N_34771,N_34808);
nor U35130 (N_35130,N_34897,N_34836);
or U35131 (N_35131,N_34912,N_34877);
nand U35132 (N_35132,N_34557,N_34791);
nor U35133 (N_35133,N_34625,N_34601);
nand U35134 (N_35134,N_34558,N_34703);
nand U35135 (N_35135,N_34668,N_34895);
xor U35136 (N_35136,N_34957,N_34670);
nor U35137 (N_35137,N_34615,N_34888);
nor U35138 (N_35138,N_34866,N_34593);
nand U35139 (N_35139,N_34906,N_34827);
and U35140 (N_35140,N_34820,N_34889);
nor U35141 (N_35141,N_34991,N_34772);
or U35142 (N_35142,N_34629,N_34798);
and U35143 (N_35143,N_34784,N_34787);
and U35144 (N_35144,N_34696,N_34802);
xnor U35145 (N_35145,N_34743,N_34892);
or U35146 (N_35146,N_34594,N_34916);
nand U35147 (N_35147,N_34780,N_34965);
or U35148 (N_35148,N_34673,N_34581);
nand U35149 (N_35149,N_34744,N_34821);
and U35150 (N_35150,N_34973,N_34915);
nand U35151 (N_35151,N_34733,N_34929);
nand U35152 (N_35152,N_34562,N_34768);
and U35153 (N_35153,N_34651,N_34574);
nand U35154 (N_35154,N_34591,N_34812);
nand U35155 (N_35155,N_34978,N_34677);
and U35156 (N_35156,N_34885,N_34996);
or U35157 (N_35157,N_34904,N_34959);
nand U35158 (N_35158,N_34861,N_34624);
or U35159 (N_35159,N_34893,N_34898);
nand U35160 (N_35160,N_34595,N_34914);
xor U35161 (N_35161,N_34694,N_34606);
xnor U35162 (N_35162,N_34757,N_34671);
nor U35163 (N_35163,N_34796,N_34951);
or U35164 (N_35164,N_34950,N_34945);
and U35165 (N_35165,N_34964,N_34626);
nor U35166 (N_35166,N_34568,N_34851);
nand U35167 (N_35167,N_34646,N_34882);
and U35168 (N_35168,N_34967,N_34521);
nor U35169 (N_35169,N_34532,N_34739);
nand U35170 (N_35170,N_34567,N_34842);
or U35171 (N_35171,N_34700,N_34881);
nor U35172 (N_35172,N_34969,N_34550);
or U35173 (N_35173,N_34529,N_34701);
nor U35174 (N_35174,N_34682,N_34520);
and U35175 (N_35175,N_34602,N_34634);
nand U35176 (N_35176,N_34936,N_34613);
nor U35177 (N_35177,N_34799,N_34762);
nand U35178 (N_35178,N_34942,N_34725);
nor U35179 (N_35179,N_34792,N_34778);
nand U35180 (N_35180,N_34949,N_34997);
nand U35181 (N_35181,N_34849,N_34542);
nor U35182 (N_35182,N_34647,N_34611);
xor U35183 (N_35183,N_34966,N_34775);
nand U35184 (N_35184,N_34980,N_34930);
and U35185 (N_35185,N_34913,N_34747);
nor U35186 (N_35186,N_34862,N_34642);
nor U35187 (N_35187,N_34695,N_34723);
nand U35188 (N_35188,N_34745,N_34556);
or U35189 (N_35189,N_34968,N_34508);
nand U35190 (N_35190,N_34526,N_34584);
nor U35191 (N_35191,N_34680,N_34511);
nor U35192 (N_35192,N_34618,N_34777);
or U35193 (N_35193,N_34717,N_34767);
nand U35194 (N_35194,N_34828,N_34643);
or U35195 (N_35195,N_34719,N_34630);
xor U35196 (N_35196,N_34731,N_34502);
and U35197 (N_35197,N_34659,N_34948);
or U35198 (N_35198,N_34522,N_34692);
and U35199 (N_35199,N_34576,N_34811);
xor U35200 (N_35200,N_34806,N_34759);
or U35201 (N_35201,N_34845,N_34720);
nand U35202 (N_35202,N_34872,N_34760);
and U35203 (N_35203,N_34985,N_34938);
nand U35204 (N_35204,N_34547,N_34874);
and U35205 (N_35205,N_34933,N_34686);
and U35206 (N_35206,N_34631,N_34900);
nor U35207 (N_35207,N_34863,N_34953);
or U35208 (N_35208,N_34774,N_34585);
or U35209 (N_35209,N_34730,N_34838);
and U35210 (N_35210,N_34636,N_34749);
nor U35211 (N_35211,N_34848,N_34727);
or U35212 (N_35212,N_34909,N_34608);
and U35213 (N_35213,N_34833,N_34752);
nor U35214 (N_35214,N_34617,N_34846);
or U35215 (N_35215,N_34884,N_34650);
and U35216 (N_35216,N_34599,N_34712);
and U35217 (N_35217,N_34962,N_34637);
nor U35218 (N_35218,N_34687,N_34795);
or U35219 (N_35219,N_34894,N_34990);
and U35220 (N_35220,N_34592,N_34920);
nand U35221 (N_35221,N_34586,N_34764);
nand U35222 (N_35222,N_34875,N_34561);
and U35223 (N_35223,N_34883,N_34896);
nand U35224 (N_35224,N_34785,N_34857);
nand U35225 (N_35225,N_34635,N_34905);
nor U35226 (N_35226,N_34854,N_34589);
nand U35227 (N_35227,N_34531,N_34989);
or U35228 (N_35228,N_34709,N_34850);
or U35229 (N_35229,N_34679,N_34755);
nand U35230 (N_35230,N_34674,N_34924);
xor U35231 (N_35231,N_34710,N_34941);
nand U35232 (N_35232,N_34939,N_34543);
xor U35233 (N_35233,N_34880,N_34911);
or U35234 (N_35234,N_34869,N_34614);
or U35235 (N_35235,N_34844,N_34878);
and U35236 (N_35236,N_34536,N_34741);
nor U35237 (N_35237,N_34676,N_34519);
nand U35238 (N_35238,N_34934,N_34870);
nand U35239 (N_35239,N_34699,N_34524);
or U35240 (N_35240,N_34891,N_34657);
and U35241 (N_35241,N_34638,N_34560);
nor U35242 (N_35242,N_34596,N_34822);
nor U35243 (N_35243,N_34656,N_34983);
nand U35244 (N_35244,N_34807,N_34992);
or U35245 (N_35245,N_34603,N_34535);
nand U35246 (N_35246,N_34946,N_34540);
or U35247 (N_35247,N_34736,N_34834);
nor U35248 (N_35248,N_34742,N_34902);
or U35249 (N_35249,N_34654,N_34839);
nor U35250 (N_35250,N_34575,N_34780);
and U35251 (N_35251,N_34914,N_34771);
and U35252 (N_35252,N_34664,N_34880);
or U35253 (N_35253,N_34761,N_34843);
xnor U35254 (N_35254,N_34715,N_34581);
and U35255 (N_35255,N_34846,N_34587);
nor U35256 (N_35256,N_34605,N_34704);
or U35257 (N_35257,N_34821,N_34845);
nor U35258 (N_35258,N_34654,N_34650);
xnor U35259 (N_35259,N_34851,N_34739);
nand U35260 (N_35260,N_34782,N_34962);
nor U35261 (N_35261,N_34711,N_34586);
or U35262 (N_35262,N_34780,N_34642);
nand U35263 (N_35263,N_34835,N_34694);
nor U35264 (N_35264,N_34850,N_34630);
or U35265 (N_35265,N_34795,N_34875);
nor U35266 (N_35266,N_34932,N_34785);
nand U35267 (N_35267,N_34948,N_34570);
nand U35268 (N_35268,N_34617,N_34620);
xnor U35269 (N_35269,N_34660,N_34822);
and U35270 (N_35270,N_34557,N_34708);
nor U35271 (N_35271,N_34781,N_34719);
nand U35272 (N_35272,N_34797,N_34643);
nand U35273 (N_35273,N_34664,N_34540);
nor U35274 (N_35274,N_34736,N_34885);
and U35275 (N_35275,N_34847,N_34639);
or U35276 (N_35276,N_34794,N_34965);
nand U35277 (N_35277,N_34827,N_34753);
nor U35278 (N_35278,N_34757,N_34695);
or U35279 (N_35279,N_34827,N_34953);
and U35280 (N_35280,N_34511,N_34915);
nand U35281 (N_35281,N_34784,N_34765);
and U35282 (N_35282,N_34866,N_34689);
nand U35283 (N_35283,N_34844,N_34987);
nand U35284 (N_35284,N_34753,N_34953);
xor U35285 (N_35285,N_34904,N_34814);
nor U35286 (N_35286,N_34844,N_34606);
xor U35287 (N_35287,N_34997,N_34580);
nor U35288 (N_35288,N_34513,N_34854);
nand U35289 (N_35289,N_34639,N_34781);
nor U35290 (N_35290,N_34866,N_34730);
nand U35291 (N_35291,N_34946,N_34800);
xor U35292 (N_35292,N_34988,N_34601);
xor U35293 (N_35293,N_34988,N_34651);
and U35294 (N_35294,N_34520,N_34879);
and U35295 (N_35295,N_34680,N_34512);
nor U35296 (N_35296,N_34893,N_34731);
and U35297 (N_35297,N_34996,N_34500);
and U35298 (N_35298,N_34527,N_34739);
nor U35299 (N_35299,N_34846,N_34863);
or U35300 (N_35300,N_34997,N_34729);
and U35301 (N_35301,N_34715,N_34661);
or U35302 (N_35302,N_34635,N_34962);
or U35303 (N_35303,N_34733,N_34576);
nor U35304 (N_35304,N_34848,N_34537);
or U35305 (N_35305,N_34893,N_34844);
xnor U35306 (N_35306,N_34900,N_34535);
and U35307 (N_35307,N_34716,N_34994);
or U35308 (N_35308,N_34840,N_34907);
nand U35309 (N_35309,N_34544,N_34618);
or U35310 (N_35310,N_34742,N_34711);
nor U35311 (N_35311,N_34919,N_34627);
xnor U35312 (N_35312,N_34507,N_34722);
xor U35313 (N_35313,N_34721,N_34841);
or U35314 (N_35314,N_34989,N_34943);
and U35315 (N_35315,N_34693,N_34965);
and U35316 (N_35316,N_34763,N_34651);
nand U35317 (N_35317,N_34583,N_34903);
and U35318 (N_35318,N_34539,N_34925);
or U35319 (N_35319,N_34579,N_34565);
and U35320 (N_35320,N_34921,N_34710);
or U35321 (N_35321,N_34682,N_34963);
and U35322 (N_35322,N_34534,N_34973);
nor U35323 (N_35323,N_34723,N_34692);
nor U35324 (N_35324,N_34919,N_34761);
or U35325 (N_35325,N_34701,N_34873);
nor U35326 (N_35326,N_34774,N_34633);
xor U35327 (N_35327,N_34963,N_34932);
nor U35328 (N_35328,N_34720,N_34568);
and U35329 (N_35329,N_34583,N_34837);
and U35330 (N_35330,N_34687,N_34508);
nor U35331 (N_35331,N_34625,N_34540);
and U35332 (N_35332,N_34659,N_34533);
nand U35333 (N_35333,N_34972,N_34653);
and U35334 (N_35334,N_34651,N_34979);
or U35335 (N_35335,N_34768,N_34520);
nand U35336 (N_35336,N_34979,N_34509);
and U35337 (N_35337,N_34632,N_34520);
nor U35338 (N_35338,N_34507,N_34858);
nor U35339 (N_35339,N_34712,N_34644);
and U35340 (N_35340,N_34942,N_34890);
or U35341 (N_35341,N_34996,N_34713);
nor U35342 (N_35342,N_34848,N_34542);
nor U35343 (N_35343,N_34710,N_34589);
or U35344 (N_35344,N_34914,N_34789);
nor U35345 (N_35345,N_34575,N_34889);
and U35346 (N_35346,N_34693,N_34526);
and U35347 (N_35347,N_34740,N_34966);
nand U35348 (N_35348,N_34590,N_34900);
nor U35349 (N_35349,N_34593,N_34749);
xor U35350 (N_35350,N_34747,N_34939);
nor U35351 (N_35351,N_34566,N_34692);
or U35352 (N_35352,N_34895,N_34663);
nor U35353 (N_35353,N_34519,N_34951);
xor U35354 (N_35354,N_34985,N_34853);
or U35355 (N_35355,N_34691,N_34909);
nand U35356 (N_35356,N_34737,N_34980);
nor U35357 (N_35357,N_34836,N_34843);
and U35358 (N_35358,N_34566,N_34806);
and U35359 (N_35359,N_34958,N_34763);
nand U35360 (N_35360,N_34670,N_34599);
nand U35361 (N_35361,N_34779,N_34544);
nand U35362 (N_35362,N_34802,N_34525);
nand U35363 (N_35363,N_34636,N_34625);
and U35364 (N_35364,N_34986,N_34698);
xor U35365 (N_35365,N_34905,N_34759);
nand U35366 (N_35366,N_34893,N_34546);
nand U35367 (N_35367,N_34920,N_34622);
xor U35368 (N_35368,N_34866,N_34776);
and U35369 (N_35369,N_34564,N_34899);
xnor U35370 (N_35370,N_34658,N_34943);
xnor U35371 (N_35371,N_34752,N_34618);
and U35372 (N_35372,N_34760,N_34547);
nand U35373 (N_35373,N_34671,N_34688);
and U35374 (N_35374,N_34718,N_34896);
or U35375 (N_35375,N_34981,N_34896);
and U35376 (N_35376,N_34954,N_34625);
xor U35377 (N_35377,N_34584,N_34830);
nor U35378 (N_35378,N_34802,N_34772);
and U35379 (N_35379,N_34897,N_34893);
nor U35380 (N_35380,N_34904,N_34998);
nand U35381 (N_35381,N_34997,N_34857);
or U35382 (N_35382,N_34687,N_34925);
xnor U35383 (N_35383,N_34993,N_34588);
nor U35384 (N_35384,N_34524,N_34526);
nor U35385 (N_35385,N_34804,N_34746);
nand U35386 (N_35386,N_34877,N_34956);
nand U35387 (N_35387,N_34904,N_34917);
nand U35388 (N_35388,N_34756,N_34524);
and U35389 (N_35389,N_34772,N_34558);
nor U35390 (N_35390,N_34534,N_34720);
nand U35391 (N_35391,N_34514,N_34899);
and U35392 (N_35392,N_34570,N_34858);
or U35393 (N_35393,N_34557,N_34631);
nor U35394 (N_35394,N_34524,N_34513);
or U35395 (N_35395,N_34678,N_34931);
xnor U35396 (N_35396,N_34585,N_34764);
nand U35397 (N_35397,N_34593,N_34522);
nor U35398 (N_35398,N_34763,N_34969);
xnor U35399 (N_35399,N_34969,N_34707);
and U35400 (N_35400,N_34527,N_34554);
or U35401 (N_35401,N_34919,N_34821);
nand U35402 (N_35402,N_34524,N_34760);
nor U35403 (N_35403,N_34630,N_34683);
nor U35404 (N_35404,N_34739,N_34584);
and U35405 (N_35405,N_34688,N_34905);
or U35406 (N_35406,N_34934,N_34574);
nand U35407 (N_35407,N_34946,N_34508);
nand U35408 (N_35408,N_34647,N_34523);
and U35409 (N_35409,N_34632,N_34818);
nand U35410 (N_35410,N_34541,N_34527);
or U35411 (N_35411,N_34769,N_34935);
and U35412 (N_35412,N_34944,N_34563);
nor U35413 (N_35413,N_34859,N_34725);
or U35414 (N_35414,N_34706,N_34878);
and U35415 (N_35415,N_34582,N_34660);
or U35416 (N_35416,N_34719,N_34760);
nand U35417 (N_35417,N_34820,N_34543);
nand U35418 (N_35418,N_34588,N_34942);
nand U35419 (N_35419,N_34801,N_34703);
nor U35420 (N_35420,N_34777,N_34570);
nor U35421 (N_35421,N_34957,N_34674);
xnor U35422 (N_35422,N_34909,N_34738);
xor U35423 (N_35423,N_34927,N_34990);
or U35424 (N_35424,N_34613,N_34771);
and U35425 (N_35425,N_34544,N_34884);
nand U35426 (N_35426,N_34913,N_34814);
and U35427 (N_35427,N_34976,N_34908);
nand U35428 (N_35428,N_34891,N_34904);
and U35429 (N_35429,N_34696,N_34711);
nand U35430 (N_35430,N_34971,N_34597);
nand U35431 (N_35431,N_34835,N_34763);
or U35432 (N_35432,N_34585,N_34643);
and U35433 (N_35433,N_34937,N_34728);
nor U35434 (N_35434,N_34780,N_34868);
or U35435 (N_35435,N_34939,N_34704);
and U35436 (N_35436,N_34711,N_34882);
and U35437 (N_35437,N_34769,N_34848);
and U35438 (N_35438,N_34758,N_34990);
or U35439 (N_35439,N_34778,N_34737);
and U35440 (N_35440,N_34529,N_34918);
nor U35441 (N_35441,N_34986,N_34782);
or U35442 (N_35442,N_34970,N_34759);
or U35443 (N_35443,N_34728,N_34562);
xor U35444 (N_35444,N_34825,N_34531);
or U35445 (N_35445,N_34784,N_34705);
xor U35446 (N_35446,N_34931,N_34569);
and U35447 (N_35447,N_34613,N_34725);
and U35448 (N_35448,N_34952,N_34863);
or U35449 (N_35449,N_34819,N_34888);
nor U35450 (N_35450,N_34899,N_34907);
or U35451 (N_35451,N_34617,N_34803);
nand U35452 (N_35452,N_34874,N_34755);
nor U35453 (N_35453,N_34720,N_34867);
or U35454 (N_35454,N_34912,N_34829);
nor U35455 (N_35455,N_34642,N_34749);
nor U35456 (N_35456,N_34608,N_34586);
nand U35457 (N_35457,N_34909,N_34692);
or U35458 (N_35458,N_34807,N_34872);
nor U35459 (N_35459,N_34818,N_34565);
and U35460 (N_35460,N_34587,N_34788);
or U35461 (N_35461,N_34551,N_34990);
nor U35462 (N_35462,N_34946,N_34911);
nor U35463 (N_35463,N_34908,N_34885);
nor U35464 (N_35464,N_34540,N_34870);
or U35465 (N_35465,N_34769,N_34775);
nand U35466 (N_35466,N_34825,N_34522);
xnor U35467 (N_35467,N_34899,N_34600);
and U35468 (N_35468,N_34756,N_34904);
and U35469 (N_35469,N_34919,N_34965);
or U35470 (N_35470,N_34642,N_34794);
nand U35471 (N_35471,N_34563,N_34609);
nand U35472 (N_35472,N_34781,N_34993);
and U35473 (N_35473,N_34784,N_34529);
xnor U35474 (N_35474,N_34879,N_34633);
and U35475 (N_35475,N_34909,N_34647);
xor U35476 (N_35476,N_34657,N_34712);
and U35477 (N_35477,N_34913,N_34917);
xnor U35478 (N_35478,N_34603,N_34526);
and U35479 (N_35479,N_34907,N_34524);
nand U35480 (N_35480,N_34609,N_34804);
xnor U35481 (N_35481,N_34565,N_34994);
nor U35482 (N_35482,N_34633,N_34565);
or U35483 (N_35483,N_34904,N_34771);
nor U35484 (N_35484,N_34675,N_34885);
and U35485 (N_35485,N_34824,N_34830);
nor U35486 (N_35486,N_34937,N_34968);
and U35487 (N_35487,N_34710,N_34994);
xor U35488 (N_35488,N_34704,N_34814);
nor U35489 (N_35489,N_34624,N_34737);
nor U35490 (N_35490,N_34832,N_34528);
xnor U35491 (N_35491,N_34992,N_34663);
and U35492 (N_35492,N_34862,N_34652);
or U35493 (N_35493,N_34529,N_34821);
and U35494 (N_35494,N_34691,N_34510);
and U35495 (N_35495,N_34959,N_34540);
or U35496 (N_35496,N_34992,N_34830);
nand U35497 (N_35497,N_34904,N_34979);
and U35498 (N_35498,N_34595,N_34627);
nor U35499 (N_35499,N_34697,N_34643);
nand U35500 (N_35500,N_35008,N_35454);
nor U35501 (N_35501,N_35348,N_35121);
and U35502 (N_35502,N_35272,N_35016);
or U35503 (N_35503,N_35015,N_35284);
xor U35504 (N_35504,N_35104,N_35266);
nor U35505 (N_35505,N_35241,N_35071);
nor U35506 (N_35506,N_35084,N_35079);
or U35507 (N_35507,N_35080,N_35423);
nand U35508 (N_35508,N_35384,N_35294);
or U35509 (N_35509,N_35356,N_35263);
nand U35510 (N_35510,N_35486,N_35339);
and U35511 (N_35511,N_35493,N_35017);
nand U35512 (N_35512,N_35029,N_35236);
and U35513 (N_35513,N_35329,N_35485);
or U35514 (N_35514,N_35393,N_35099);
nand U35515 (N_35515,N_35377,N_35221);
or U35516 (N_35516,N_35004,N_35176);
or U35517 (N_35517,N_35380,N_35499);
nand U35518 (N_35518,N_35042,N_35212);
nor U35519 (N_35519,N_35434,N_35382);
or U35520 (N_35520,N_35129,N_35445);
nor U35521 (N_35521,N_35220,N_35180);
nor U35522 (N_35522,N_35480,N_35412);
and U35523 (N_35523,N_35208,N_35170);
xor U35524 (N_35524,N_35298,N_35025);
nor U35525 (N_35525,N_35333,N_35438);
nor U35526 (N_35526,N_35216,N_35268);
xnor U35527 (N_35527,N_35363,N_35094);
or U35528 (N_35528,N_35245,N_35228);
and U35529 (N_35529,N_35422,N_35488);
and U35530 (N_35530,N_35058,N_35087);
nor U35531 (N_35531,N_35355,N_35137);
nand U35532 (N_35532,N_35000,N_35197);
xor U35533 (N_35533,N_35336,N_35174);
or U35534 (N_35534,N_35239,N_35051);
or U35535 (N_35535,N_35097,N_35037);
nor U35536 (N_35536,N_35184,N_35354);
nand U35537 (N_35537,N_35478,N_35307);
xor U35538 (N_35538,N_35372,N_35319);
and U35539 (N_35539,N_35277,N_35128);
or U35540 (N_35540,N_35096,N_35046);
and U35541 (N_35541,N_35479,N_35052);
and U35542 (N_35542,N_35295,N_35158);
or U35543 (N_35543,N_35160,N_35491);
or U35544 (N_35544,N_35067,N_35142);
and U35545 (N_35545,N_35040,N_35113);
nand U35546 (N_35546,N_35278,N_35374);
nand U35547 (N_35547,N_35111,N_35465);
nor U35548 (N_35548,N_35243,N_35078);
and U35549 (N_35549,N_35464,N_35282);
nand U35550 (N_35550,N_35033,N_35381);
nor U35551 (N_35551,N_35256,N_35063);
nor U35552 (N_35552,N_35392,N_35118);
or U35553 (N_35553,N_35152,N_35075);
nand U35554 (N_35554,N_35300,N_35274);
and U35555 (N_35555,N_35035,N_35145);
or U35556 (N_35556,N_35162,N_35312);
and U35557 (N_35557,N_35141,N_35291);
xor U35558 (N_35558,N_35270,N_35386);
and U35559 (N_35559,N_35007,N_35242);
and U35560 (N_35560,N_35472,N_35189);
nand U35561 (N_35561,N_35019,N_35108);
xnor U35562 (N_35562,N_35202,N_35313);
nor U35563 (N_35563,N_35124,N_35191);
and U35564 (N_35564,N_35089,N_35116);
xnor U35565 (N_35565,N_35461,N_35012);
nor U35566 (N_35566,N_35367,N_35062);
nor U35567 (N_35567,N_35166,N_35290);
nand U35568 (N_35568,N_35095,N_35205);
nand U35569 (N_35569,N_35093,N_35168);
or U35570 (N_35570,N_35332,N_35181);
nand U35571 (N_35571,N_35059,N_35149);
xnor U35572 (N_35572,N_35352,N_35322);
and U35573 (N_35573,N_35287,N_35458);
xnor U35574 (N_35574,N_35143,N_35098);
nor U35575 (N_35575,N_35131,N_35450);
nand U35576 (N_35576,N_35110,N_35135);
nand U35577 (N_35577,N_35378,N_35476);
or U35578 (N_35578,N_35482,N_35020);
and U35579 (N_35579,N_35224,N_35413);
and U35580 (N_35580,N_35171,N_35253);
nand U35581 (N_35581,N_35473,N_35144);
and U35582 (N_35582,N_35292,N_35267);
and U35583 (N_35583,N_35195,N_35314);
xor U35584 (N_35584,N_35351,N_35342);
nor U35585 (N_35585,N_35315,N_35361);
or U35586 (N_35586,N_35109,N_35090);
or U35587 (N_35587,N_35250,N_35402);
and U35588 (N_35588,N_35177,N_35261);
or U35589 (N_35589,N_35376,N_35030);
nor U35590 (N_35590,N_35349,N_35249);
nor U35591 (N_35591,N_35350,N_35320);
nand U35592 (N_35592,N_35390,N_35061);
nand U35593 (N_35593,N_35175,N_35417);
xor U35594 (N_35594,N_35193,N_35082);
nor U35595 (N_35595,N_35383,N_35182);
or U35596 (N_35596,N_35070,N_35091);
and U35597 (N_35597,N_35188,N_35123);
nor U35598 (N_35598,N_35229,N_35130);
or U35599 (N_35599,N_35397,N_35132);
or U35600 (N_35600,N_35173,N_35011);
nor U35601 (N_35601,N_35436,N_35023);
and U35602 (N_35602,N_35009,N_35178);
and U35603 (N_35603,N_35254,N_35214);
nor U35604 (N_35604,N_35013,N_35448);
or U35605 (N_35605,N_35153,N_35271);
or U35606 (N_35606,N_35306,N_35244);
nand U35607 (N_35607,N_35446,N_35398);
nor U35608 (N_35608,N_35433,N_35022);
nand U35609 (N_35609,N_35334,N_35498);
nor U35610 (N_35610,N_35474,N_35321);
or U35611 (N_35611,N_35369,N_35150);
and U35612 (N_35612,N_35497,N_35155);
nor U35613 (N_35613,N_35200,N_35201);
and U35614 (N_35614,N_35204,N_35437);
and U35615 (N_35615,N_35154,N_35257);
nand U35616 (N_35616,N_35086,N_35100);
nor U35617 (N_35617,N_35006,N_35400);
nor U35618 (N_35618,N_35072,N_35440);
nor U35619 (N_35619,N_35330,N_35183);
nand U35620 (N_35620,N_35134,N_35347);
nor U35621 (N_35621,N_35368,N_35186);
nand U35622 (N_35622,N_35489,N_35353);
or U35623 (N_35623,N_35388,N_35280);
xor U35624 (N_35624,N_35206,N_35238);
nor U35625 (N_35625,N_35112,N_35260);
xnor U35626 (N_35626,N_35456,N_35496);
nor U35627 (N_35627,N_35466,N_35223);
or U35628 (N_35628,N_35428,N_35467);
or U35629 (N_35629,N_35408,N_35389);
nor U35630 (N_35630,N_35230,N_35199);
nand U35631 (N_35631,N_35039,N_35288);
nor U35632 (N_35632,N_35275,N_35069);
nor U35633 (N_35633,N_35045,N_35081);
xor U35634 (N_35634,N_35021,N_35165);
nand U35635 (N_35635,N_35407,N_35049);
nand U35636 (N_35636,N_35136,N_35379);
nor U35637 (N_35637,N_35126,N_35034);
or U35638 (N_35638,N_35430,N_35431);
xnor U35639 (N_35639,N_35140,N_35117);
nor U35640 (N_35640,N_35327,N_35451);
nand U35641 (N_35641,N_35146,N_35262);
and U35642 (N_35642,N_35296,N_35490);
nand U35643 (N_35643,N_35005,N_35439);
or U35644 (N_35644,N_35305,N_35010);
and U35645 (N_35645,N_35289,N_35370);
nor U35646 (N_35646,N_35442,N_35432);
nor U35647 (N_35647,N_35304,N_35470);
or U35648 (N_35648,N_35255,N_35391);
nand U35649 (N_35649,N_35102,N_35452);
nand U35650 (N_35650,N_35163,N_35032);
and U35651 (N_35651,N_35138,N_35198);
xnor U35652 (N_35652,N_35468,N_35222);
and U35653 (N_35653,N_35418,N_35416);
and U35654 (N_35654,N_35366,N_35215);
nor U35655 (N_35655,N_35043,N_35469);
nand U35656 (N_35656,N_35429,N_35317);
xor U35657 (N_35657,N_35285,N_35399);
nand U35658 (N_35658,N_35056,N_35237);
and U35659 (N_35659,N_35073,N_35065);
nand U35660 (N_35660,N_35234,N_35101);
and U35661 (N_35661,N_35068,N_35394);
nand U35662 (N_35662,N_35028,N_35139);
or U35663 (N_35663,N_35103,N_35167);
xnor U35664 (N_35664,N_35323,N_35457);
nand U35665 (N_35665,N_35328,N_35106);
and U35666 (N_35666,N_35425,N_35147);
nand U35667 (N_35667,N_35447,N_35460);
nor U35668 (N_35668,N_35325,N_35246);
nand U35669 (N_35669,N_35083,N_35259);
nand U35670 (N_35670,N_35455,N_35481);
nor U35671 (N_35671,N_35395,N_35148);
xor U35672 (N_35672,N_35426,N_35341);
and U35673 (N_35673,N_35211,N_35053);
and U35674 (N_35674,N_35286,N_35415);
xor U35675 (N_35675,N_35044,N_35459);
or U35676 (N_35676,N_35401,N_35258);
nand U35677 (N_35677,N_35346,N_35210);
nand U35678 (N_35678,N_35421,N_35494);
and U35679 (N_35679,N_35419,N_35269);
and U35680 (N_35680,N_35424,N_35218);
or U35681 (N_35681,N_35396,N_35427);
or U35682 (N_35682,N_35151,N_35406);
nand U35683 (N_35683,N_35303,N_35443);
nand U35684 (N_35684,N_35105,N_35156);
or U35685 (N_35685,N_35337,N_35060);
nand U35686 (N_35686,N_35283,N_35157);
and U35687 (N_35687,N_35179,N_35027);
xnor U35688 (N_35688,N_35302,N_35054);
or U35689 (N_35689,N_35127,N_35308);
nand U35690 (N_35690,N_35038,N_35492);
xnor U35691 (N_35691,N_35092,N_35251);
and U35692 (N_35692,N_35227,N_35207);
nor U35693 (N_35693,N_35014,N_35326);
nor U35694 (N_35694,N_35233,N_35344);
xor U35695 (N_35695,N_35047,N_35331);
nand U35696 (N_35696,N_35190,N_35196);
xnor U35697 (N_35697,N_35114,N_35001);
or U35698 (N_35698,N_35194,N_35404);
xor U35699 (N_35699,N_35225,N_35281);
nand U35700 (N_35700,N_35273,N_35219);
nand U35701 (N_35701,N_35449,N_35265);
nor U35702 (N_35702,N_35172,N_35018);
or U35703 (N_35703,N_35226,N_35301);
nand U35704 (N_35704,N_35159,N_35324);
and U35705 (N_35705,N_35115,N_35343);
xnor U35706 (N_35706,N_35362,N_35483);
or U35707 (N_35707,N_35041,N_35463);
and U35708 (N_35708,N_35293,N_35252);
and U35709 (N_35709,N_35475,N_35373);
or U35710 (N_35710,N_35318,N_35192);
nand U35711 (N_35711,N_35066,N_35119);
nor U35712 (N_35712,N_35164,N_35232);
nand U35713 (N_35713,N_35125,N_35364);
or U35714 (N_35714,N_35310,N_35085);
and U35715 (N_35715,N_35345,N_35120);
and U35716 (N_35716,N_35185,N_35161);
nand U35717 (N_35717,N_35031,N_35240);
and U35718 (N_35718,N_35088,N_35409);
nand U35719 (N_35719,N_35444,N_35371);
nor U35720 (N_35720,N_35385,N_35477);
and U35721 (N_35721,N_35203,N_35375);
or U35722 (N_35722,N_35026,N_35435);
and U35723 (N_35723,N_35122,N_35403);
nand U35724 (N_35724,N_35471,N_35169);
nand U35725 (N_35725,N_35024,N_35420);
nand U35726 (N_35726,N_35410,N_35359);
or U35727 (N_35727,N_35076,N_35003);
or U35728 (N_35728,N_35235,N_35411);
nand U35729 (N_35729,N_35050,N_35484);
nand U35730 (N_35730,N_35209,N_35487);
and U35731 (N_35731,N_35358,N_35231);
nand U35732 (N_35732,N_35365,N_35357);
xnor U35733 (N_35733,N_35248,N_35002);
or U35734 (N_35734,N_35405,N_35187);
or U35735 (N_35735,N_35335,N_35338);
xnor U35736 (N_35736,N_35495,N_35048);
and U35737 (N_35737,N_35453,N_35064);
nor U35738 (N_35738,N_35213,N_35360);
or U35739 (N_35739,N_35036,N_35299);
and U35740 (N_35740,N_35441,N_35340);
nor U35741 (N_35741,N_35311,N_35217);
nand U35742 (N_35742,N_35057,N_35414);
nor U35743 (N_35743,N_35264,N_35055);
xnor U35744 (N_35744,N_35279,N_35462);
xor U35745 (N_35745,N_35133,N_35387);
nand U35746 (N_35746,N_35077,N_35074);
and U35747 (N_35747,N_35107,N_35297);
or U35748 (N_35748,N_35276,N_35247);
xor U35749 (N_35749,N_35309,N_35316);
xor U35750 (N_35750,N_35249,N_35264);
and U35751 (N_35751,N_35381,N_35052);
and U35752 (N_35752,N_35269,N_35175);
xor U35753 (N_35753,N_35068,N_35353);
nor U35754 (N_35754,N_35475,N_35009);
nor U35755 (N_35755,N_35155,N_35241);
and U35756 (N_35756,N_35276,N_35174);
or U35757 (N_35757,N_35328,N_35488);
or U35758 (N_35758,N_35223,N_35326);
and U35759 (N_35759,N_35112,N_35412);
nand U35760 (N_35760,N_35022,N_35358);
nor U35761 (N_35761,N_35213,N_35059);
or U35762 (N_35762,N_35261,N_35359);
nand U35763 (N_35763,N_35278,N_35196);
nor U35764 (N_35764,N_35282,N_35237);
nand U35765 (N_35765,N_35272,N_35298);
xor U35766 (N_35766,N_35339,N_35194);
nor U35767 (N_35767,N_35354,N_35428);
xnor U35768 (N_35768,N_35207,N_35433);
and U35769 (N_35769,N_35378,N_35047);
xor U35770 (N_35770,N_35416,N_35005);
nand U35771 (N_35771,N_35247,N_35295);
or U35772 (N_35772,N_35373,N_35376);
and U35773 (N_35773,N_35250,N_35398);
nor U35774 (N_35774,N_35045,N_35199);
and U35775 (N_35775,N_35449,N_35101);
and U35776 (N_35776,N_35048,N_35323);
nand U35777 (N_35777,N_35408,N_35172);
nor U35778 (N_35778,N_35233,N_35493);
or U35779 (N_35779,N_35494,N_35134);
nor U35780 (N_35780,N_35443,N_35322);
nor U35781 (N_35781,N_35230,N_35469);
or U35782 (N_35782,N_35403,N_35493);
nor U35783 (N_35783,N_35299,N_35497);
nor U35784 (N_35784,N_35072,N_35450);
and U35785 (N_35785,N_35116,N_35115);
xor U35786 (N_35786,N_35094,N_35358);
xor U35787 (N_35787,N_35385,N_35258);
nand U35788 (N_35788,N_35019,N_35012);
nand U35789 (N_35789,N_35070,N_35499);
xnor U35790 (N_35790,N_35092,N_35398);
or U35791 (N_35791,N_35433,N_35333);
nand U35792 (N_35792,N_35090,N_35076);
xor U35793 (N_35793,N_35000,N_35454);
or U35794 (N_35794,N_35235,N_35206);
or U35795 (N_35795,N_35256,N_35045);
xnor U35796 (N_35796,N_35328,N_35353);
nor U35797 (N_35797,N_35052,N_35400);
or U35798 (N_35798,N_35385,N_35412);
nor U35799 (N_35799,N_35379,N_35493);
nor U35800 (N_35800,N_35267,N_35457);
nand U35801 (N_35801,N_35094,N_35446);
nor U35802 (N_35802,N_35486,N_35227);
nor U35803 (N_35803,N_35212,N_35275);
and U35804 (N_35804,N_35089,N_35321);
xor U35805 (N_35805,N_35226,N_35259);
or U35806 (N_35806,N_35107,N_35016);
or U35807 (N_35807,N_35325,N_35168);
nand U35808 (N_35808,N_35071,N_35382);
nand U35809 (N_35809,N_35121,N_35265);
and U35810 (N_35810,N_35120,N_35193);
nor U35811 (N_35811,N_35427,N_35288);
nor U35812 (N_35812,N_35487,N_35138);
xnor U35813 (N_35813,N_35153,N_35484);
nand U35814 (N_35814,N_35147,N_35284);
and U35815 (N_35815,N_35417,N_35086);
and U35816 (N_35816,N_35119,N_35498);
or U35817 (N_35817,N_35375,N_35119);
nand U35818 (N_35818,N_35047,N_35274);
and U35819 (N_35819,N_35156,N_35041);
and U35820 (N_35820,N_35421,N_35428);
xor U35821 (N_35821,N_35279,N_35411);
nand U35822 (N_35822,N_35447,N_35168);
or U35823 (N_35823,N_35291,N_35441);
and U35824 (N_35824,N_35464,N_35032);
nor U35825 (N_35825,N_35351,N_35272);
nand U35826 (N_35826,N_35066,N_35168);
nand U35827 (N_35827,N_35032,N_35422);
xor U35828 (N_35828,N_35126,N_35452);
or U35829 (N_35829,N_35413,N_35086);
and U35830 (N_35830,N_35033,N_35478);
and U35831 (N_35831,N_35364,N_35051);
xnor U35832 (N_35832,N_35240,N_35313);
nor U35833 (N_35833,N_35284,N_35282);
and U35834 (N_35834,N_35257,N_35368);
or U35835 (N_35835,N_35242,N_35089);
nand U35836 (N_35836,N_35048,N_35307);
and U35837 (N_35837,N_35235,N_35483);
and U35838 (N_35838,N_35445,N_35314);
and U35839 (N_35839,N_35035,N_35311);
and U35840 (N_35840,N_35287,N_35305);
nor U35841 (N_35841,N_35470,N_35145);
or U35842 (N_35842,N_35383,N_35193);
nand U35843 (N_35843,N_35253,N_35243);
or U35844 (N_35844,N_35449,N_35016);
and U35845 (N_35845,N_35163,N_35105);
nor U35846 (N_35846,N_35154,N_35089);
nor U35847 (N_35847,N_35057,N_35253);
and U35848 (N_35848,N_35439,N_35133);
or U35849 (N_35849,N_35026,N_35339);
and U35850 (N_35850,N_35340,N_35162);
nor U35851 (N_35851,N_35271,N_35129);
xor U35852 (N_35852,N_35366,N_35254);
nand U35853 (N_35853,N_35189,N_35041);
nor U35854 (N_35854,N_35253,N_35261);
or U35855 (N_35855,N_35465,N_35213);
nand U35856 (N_35856,N_35246,N_35130);
and U35857 (N_35857,N_35096,N_35198);
xor U35858 (N_35858,N_35203,N_35159);
and U35859 (N_35859,N_35407,N_35036);
and U35860 (N_35860,N_35247,N_35468);
nand U35861 (N_35861,N_35453,N_35406);
nand U35862 (N_35862,N_35021,N_35472);
and U35863 (N_35863,N_35015,N_35140);
or U35864 (N_35864,N_35032,N_35266);
nor U35865 (N_35865,N_35402,N_35063);
nor U35866 (N_35866,N_35033,N_35094);
or U35867 (N_35867,N_35249,N_35031);
nand U35868 (N_35868,N_35058,N_35021);
or U35869 (N_35869,N_35347,N_35138);
nor U35870 (N_35870,N_35069,N_35000);
nand U35871 (N_35871,N_35462,N_35484);
or U35872 (N_35872,N_35276,N_35216);
nand U35873 (N_35873,N_35407,N_35171);
xnor U35874 (N_35874,N_35206,N_35325);
nor U35875 (N_35875,N_35025,N_35419);
nor U35876 (N_35876,N_35123,N_35267);
nand U35877 (N_35877,N_35070,N_35107);
or U35878 (N_35878,N_35056,N_35029);
and U35879 (N_35879,N_35018,N_35492);
nand U35880 (N_35880,N_35314,N_35046);
and U35881 (N_35881,N_35475,N_35361);
and U35882 (N_35882,N_35120,N_35323);
and U35883 (N_35883,N_35499,N_35275);
and U35884 (N_35884,N_35029,N_35309);
nor U35885 (N_35885,N_35276,N_35115);
and U35886 (N_35886,N_35172,N_35226);
or U35887 (N_35887,N_35342,N_35260);
or U35888 (N_35888,N_35226,N_35169);
xnor U35889 (N_35889,N_35373,N_35427);
or U35890 (N_35890,N_35045,N_35308);
nand U35891 (N_35891,N_35440,N_35335);
xor U35892 (N_35892,N_35266,N_35466);
nor U35893 (N_35893,N_35163,N_35264);
nand U35894 (N_35894,N_35080,N_35171);
nor U35895 (N_35895,N_35391,N_35038);
or U35896 (N_35896,N_35353,N_35089);
and U35897 (N_35897,N_35290,N_35410);
or U35898 (N_35898,N_35000,N_35442);
xnor U35899 (N_35899,N_35393,N_35019);
or U35900 (N_35900,N_35379,N_35010);
or U35901 (N_35901,N_35076,N_35186);
and U35902 (N_35902,N_35292,N_35201);
and U35903 (N_35903,N_35139,N_35188);
and U35904 (N_35904,N_35262,N_35466);
nand U35905 (N_35905,N_35219,N_35445);
or U35906 (N_35906,N_35478,N_35077);
nor U35907 (N_35907,N_35381,N_35069);
nand U35908 (N_35908,N_35329,N_35454);
nand U35909 (N_35909,N_35494,N_35130);
nand U35910 (N_35910,N_35381,N_35439);
xor U35911 (N_35911,N_35357,N_35014);
nand U35912 (N_35912,N_35144,N_35378);
nand U35913 (N_35913,N_35396,N_35381);
and U35914 (N_35914,N_35315,N_35485);
or U35915 (N_35915,N_35442,N_35320);
or U35916 (N_35916,N_35057,N_35015);
xor U35917 (N_35917,N_35298,N_35279);
and U35918 (N_35918,N_35058,N_35129);
xnor U35919 (N_35919,N_35464,N_35098);
and U35920 (N_35920,N_35093,N_35386);
and U35921 (N_35921,N_35223,N_35289);
nor U35922 (N_35922,N_35186,N_35134);
or U35923 (N_35923,N_35450,N_35067);
and U35924 (N_35924,N_35032,N_35087);
or U35925 (N_35925,N_35187,N_35213);
nand U35926 (N_35926,N_35333,N_35014);
nor U35927 (N_35927,N_35447,N_35144);
or U35928 (N_35928,N_35295,N_35117);
and U35929 (N_35929,N_35469,N_35170);
nand U35930 (N_35930,N_35326,N_35200);
nor U35931 (N_35931,N_35174,N_35354);
or U35932 (N_35932,N_35031,N_35371);
and U35933 (N_35933,N_35170,N_35227);
nor U35934 (N_35934,N_35366,N_35127);
nor U35935 (N_35935,N_35300,N_35012);
nand U35936 (N_35936,N_35254,N_35352);
and U35937 (N_35937,N_35366,N_35315);
nor U35938 (N_35938,N_35281,N_35411);
and U35939 (N_35939,N_35427,N_35472);
or U35940 (N_35940,N_35058,N_35015);
nand U35941 (N_35941,N_35498,N_35073);
or U35942 (N_35942,N_35105,N_35394);
nand U35943 (N_35943,N_35421,N_35478);
nor U35944 (N_35944,N_35392,N_35005);
nor U35945 (N_35945,N_35114,N_35486);
or U35946 (N_35946,N_35353,N_35376);
nand U35947 (N_35947,N_35062,N_35070);
xor U35948 (N_35948,N_35489,N_35127);
or U35949 (N_35949,N_35496,N_35418);
nor U35950 (N_35950,N_35183,N_35123);
nor U35951 (N_35951,N_35340,N_35392);
and U35952 (N_35952,N_35454,N_35209);
or U35953 (N_35953,N_35407,N_35206);
and U35954 (N_35954,N_35213,N_35474);
and U35955 (N_35955,N_35037,N_35380);
and U35956 (N_35956,N_35149,N_35232);
nand U35957 (N_35957,N_35371,N_35000);
nor U35958 (N_35958,N_35414,N_35233);
nand U35959 (N_35959,N_35314,N_35448);
nor U35960 (N_35960,N_35383,N_35423);
and U35961 (N_35961,N_35036,N_35019);
nor U35962 (N_35962,N_35011,N_35022);
nand U35963 (N_35963,N_35014,N_35187);
and U35964 (N_35964,N_35176,N_35425);
nor U35965 (N_35965,N_35341,N_35003);
nand U35966 (N_35966,N_35028,N_35150);
nor U35967 (N_35967,N_35358,N_35215);
nor U35968 (N_35968,N_35269,N_35130);
xnor U35969 (N_35969,N_35493,N_35078);
and U35970 (N_35970,N_35141,N_35357);
and U35971 (N_35971,N_35127,N_35377);
nor U35972 (N_35972,N_35455,N_35257);
nand U35973 (N_35973,N_35157,N_35073);
nand U35974 (N_35974,N_35480,N_35128);
and U35975 (N_35975,N_35316,N_35176);
and U35976 (N_35976,N_35214,N_35489);
nand U35977 (N_35977,N_35233,N_35094);
and U35978 (N_35978,N_35381,N_35228);
and U35979 (N_35979,N_35344,N_35206);
xnor U35980 (N_35980,N_35497,N_35465);
xnor U35981 (N_35981,N_35374,N_35038);
or U35982 (N_35982,N_35220,N_35331);
nor U35983 (N_35983,N_35172,N_35372);
and U35984 (N_35984,N_35206,N_35160);
and U35985 (N_35985,N_35171,N_35373);
nand U35986 (N_35986,N_35199,N_35257);
nand U35987 (N_35987,N_35037,N_35455);
or U35988 (N_35988,N_35097,N_35165);
xor U35989 (N_35989,N_35113,N_35241);
or U35990 (N_35990,N_35212,N_35048);
or U35991 (N_35991,N_35187,N_35197);
nor U35992 (N_35992,N_35192,N_35241);
nand U35993 (N_35993,N_35489,N_35067);
nand U35994 (N_35994,N_35313,N_35394);
nand U35995 (N_35995,N_35365,N_35488);
and U35996 (N_35996,N_35277,N_35076);
nor U35997 (N_35997,N_35124,N_35119);
and U35998 (N_35998,N_35373,N_35332);
xor U35999 (N_35999,N_35377,N_35408);
nand U36000 (N_36000,N_35884,N_35753);
or U36001 (N_36001,N_35575,N_35903);
nor U36002 (N_36002,N_35501,N_35837);
or U36003 (N_36003,N_35504,N_35990);
and U36004 (N_36004,N_35984,N_35864);
nor U36005 (N_36005,N_35907,N_35646);
xnor U36006 (N_36006,N_35834,N_35861);
or U36007 (N_36007,N_35761,N_35820);
or U36008 (N_36008,N_35957,N_35977);
nor U36009 (N_36009,N_35866,N_35705);
nand U36010 (N_36010,N_35641,N_35602);
and U36011 (N_36011,N_35595,N_35663);
and U36012 (N_36012,N_35952,N_35686);
or U36013 (N_36013,N_35623,N_35515);
nor U36014 (N_36014,N_35905,N_35792);
xnor U36015 (N_36015,N_35956,N_35614);
or U36016 (N_36016,N_35958,N_35598);
xnor U36017 (N_36017,N_35567,N_35606);
nand U36018 (N_36018,N_35645,N_35604);
nand U36019 (N_36019,N_35513,N_35772);
nor U36020 (N_36020,N_35555,N_35719);
nor U36021 (N_36021,N_35895,N_35640);
nand U36022 (N_36022,N_35767,N_35796);
and U36023 (N_36023,N_35998,N_35927);
or U36024 (N_36024,N_35754,N_35643);
nor U36025 (N_36025,N_35676,N_35695);
nand U36026 (N_36026,N_35847,N_35890);
nor U36027 (N_36027,N_35524,N_35827);
or U36028 (N_36028,N_35625,N_35500);
or U36029 (N_36029,N_35770,N_35732);
nand U36030 (N_36030,N_35605,N_35620);
and U36031 (N_36031,N_35918,N_35526);
or U36032 (N_36032,N_35691,N_35855);
nor U36033 (N_36033,N_35896,N_35985);
nor U36034 (N_36034,N_35624,N_35774);
nand U36035 (N_36035,N_35906,N_35789);
or U36036 (N_36036,N_35523,N_35911);
nand U36037 (N_36037,N_35653,N_35502);
or U36038 (N_36038,N_35781,N_35955);
nand U36039 (N_36039,N_35739,N_35817);
or U36040 (N_36040,N_35887,N_35871);
and U36041 (N_36041,N_35878,N_35997);
xor U36042 (N_36042,N_35972,N_35565);
nand U36043 (N_36043,N_35692,N_35829);
nand U36044 (N_36044,N_35876,N_35613);
nand U36045 (N_36045,N_35718,N_35704);
nor U36046 (N_36046,N_35994,N_35745);
or U36047 (N_36047,N_35549,N_35540);
and U36048 (N_36048,N_35594,N_35910);
nor U36049 (N_36049,N_35617,N_35978);
xor U36050 (N_36050,N_35930,N_35803);
nand U36051 (N_36051,N_35703,N_35870);
and U36052 (N_36052,N_35706,N_35882);
nor U36053 (N_36053,N_35681,N_35647);
nor U36054 (N_36054,N_35800,N_35714);
nand U36055 (N_36055,N_35755,N_35971);
or U36056 (N_36056,N_35631,N_35889);
nor U36057 (N_36057,N_35669,N_35582);
nor U36058 (N_36058,N_35938,N_35945);
nor U36059 (N_36059,N_35746,N_35768);
or U36060 (N_36060,N_35959,N_35917);
nor U36061 (N_36061,N_35799,N_35844);
nor U36062 (N_36062,N_35923,N_35630);
nand U36063 (N_36063,N_35782,N_35697);
or U36064 (N_36064,N_35702,N_35852);
nand U36065 (N_36065,N_35939,N_35811);
nand U36066 (N_36066,N_35675,N_35795);
nand U36067 (N_36067,N_35726,N_35912);
and U36068 (N_36068,N_35699,N_35881);
and U36069 (N_36069,N_35875,N_35762);
nor U36070 (N_36070,N_35758,N_35727);
nor U36071 (N_36071,N_35514,N_35824);
and U36072 (N_36072,N_35892,N_35966);
or U36073 (N_36073,N_35511,N_35813);
or U36074 (N_36074,N_35672,N_35995);
xnor U36075 (N_36075,N_35693,N_35833);
nand U36076 (N_36076,N_35585,N_35748);
and U36077 (N_36077,N_35724,N_35788);
or U36078 (N_36078,N_35583,N_35544);
xor U36079 (N_36079,N_35969,N_35763);
nor U36080 (N_36080,N_35948,N_35859);
nand U36081 (N_36081,N_35668,N_35836);
or U36082 (N_36082,N_35532,N_35991);
and U36083 (N_36083,N_35557,N_35798);
and U36084 (N_36084,N_35596,N_35964);
or U36085 (N_36085,N_35783,N_35553);
nor U36086 (N_36086,N_35715,N_35729);
nor U36087 (N_36087,N_35636,N_35562);
nor U36088 (N_36088,N_35518,N_35684);
and U36089 (N_36089,N_35778,N_35944);
nand U36090 (N_36090,N_35909,N_35512);
and U36091 (N_36091,N_35850,N_35510);
and U36092 (N_36092,N_35541,N_35527);
or U36093 (N_36093,N_35935,N_35588);
nor U36094 (N_36094,N_35552,N_35635);
nor U36095 (N_36095,N_35913,N_35577);
and U36096 (N_36096,N_35794,N_35741);
nor U36097 (N_36097,N_35670,N_35973);
nand U36098 (N_36098,N_35872,N_35776);
or U36099 (N_36099,N_35825,N_35603);
nor U36100 (N_36100,N_35786,N_35908);
or U36101 (N_36101,N_35769,N_35550);
nor U36102 (N_36102,N_35943,N_35810);
nor U36103 (N_36103,N_35738,N_35722);
and U36104 (N_36104,N_35520,N_35733);
and U36105 (N_36105,N_35611,N_35534);
nor U36106 (N_36106,N_35900,N_35656);
nor U36107 (N_36107,N_35951,N_35965);
and U36108 (N_36108,N_35785,N_35961);
and U36109 (N_36109,N_35728,N_35919);
and U36110 (N_36110,N_35560,N_35987);
or U36111 (N_36111,N_35655,N_35673);
or U36112 (N_36112,N_35559,N_35982);
nor U36113 (N_36113,N_35659,N_35954);
nand U36114 (N_36114,N_35507,N_35897);
or U36115 (N_36115,N_35581,N_35642);
nor U36116 (N_36116,N_35516,N_35519);
or U36117 (N_36117,N_35937,N_35626);
nor U36118 (N_36118,N_35573,N_35536);
nand U36119 (N_36119,N_35627,N_35902);
or U36120 (N_36120,N_35723,N_35926);
or U36121 (N_36121,N_35616,N_35815);
nand U36122 (N_36122,N_35946,N_35886);
nor U36123 (N_36123,N_35531,N_35894);
nor U36124 (N_36124,N_35563,N_35752);
nand U36125 (N_36125,N_35537,N_35868);
nor U36126 (N_36126,N_35806,N_35853);
nand U36127 (N_36127,N_35564,N_35717);
or U36128 (N_36128,N_35849,N_35891);
nor U36129 (N_36129,N_35637,N_35931);
or U36130 (N_36130,N_35867,N_35747);
nand U36131 (N_36131,N_35708,N_35694);
nor U36132 (N_36132,N_35962,N_35974);
or U36133 (N_36133,N_35545,N_35830);
nand U36134 (N_36134,N_35756,N_35947);
xor U36135 (N_36135,N_35671,N_35713);
and U36136 (N_36136,N_35734,N_35873);
nor U36137 (N_36137,N_35780,N_35683);
nor U36138 (N_36138,N_35760,N_35509);
nand U36139 (N_36139,N_35993,N_35765);
or U36140 (N_36140,N_35571,N_35757);
nor U36141 (N_36141,N_35576,N_35766);
and U36142 (N_36142,N_35899,N_35814);
xnor U36143 (N_36143,N_35856,N_35823);
or U36144 (N_36144,N_35579,N_35690);
nor U36145 (N_36145,N_35816,N_35660);
or U36146 (N_36146,N_35775,N_35835);
nor U36147 (N_36147,N_35615,N_35589);
nor U36148 (N_36148,N_35628,N_35858);
and U36149 (N_36149,N_35933,N_35644);
or U36150 (N_36150,N_35929,N_35879);
nor U36151 (N_36151,N_35790,N_35779);
or U36152 (N_36152,N_35578,N_35593);
nand U36153 (N_36153,N_35530,N_35730);
xor U36154 (N_36154,N_35970,N_35546);
and U36155 (N_36155,N_35880,N_35522);
nand U36156 (N_36156,N_35677,N_35904);
nor U36157 (N_36157,N_35877,N_35983);
xor U36158 (N_36158,N_35716,N_35701);
and U36159 (N_36159,N_35901,N_35561);
or U36160 (N_36160,N_35648,N_35821);
or U36161 (N_36161,N_35700,N_35934);
nor U36162 (N_36162,N_35942,N_35740);
nand U36163 (N_36163,N_35538,N_35865);
or U36164 (N_36164,N_35771,N_35601);
or U36165 (N_36165,N_35689,N_35525);
nor U36166 (N_36166,N_35976,N_35953);
nor U36167 (N_36167,N_35967,N_35529);
or U36168 (N_36168,N_35711,N_35822);
nand U36169 (N_36169,N_35725,N_35869);
or U36170 (N_36170,N_35599,N_35721);
and U36171 (N_36171,N_35570,N_35787);
xor U36172 (N_36172,N_35652,N_35916);
nor U36173 (N_36173,N_35503,N_35543);
nor U36174 (N_36174,N_35720,N_35517);
nand U36175 (N_36175,N_35883,N_35674);
or U36176 (N_36176,N_35742,N_35936);
nand U36177 (N_36177,N_35622,N_35940);
or U36178 (N_36178,N_35651,N_35558);
nand U36179 (N_36179,N_35857,N_35840);
or U36180 (N_36180,N_35922,N_35506);
or U36181 (N_36181,N_35841,N_35664);
and U36182 (N_36182,N_35678,N_35609);
xor U36183 (N_36183,N_35914,N_35759);
nor U36184 (N_36184,N_35547,N_35851);
nand U36185 (N_36185,N_35839,N_35633);
nor U36186 (N_36186,N_35709,N_35793);
or U36187 (N_36187,N_35863,N_35791);
nor U36188 (N_36188,N_35736,N_35542);
or U36189 (N_36189,N_35607,N_35963);
and U36190 (N_36190,N_35621,N_35843);
nor U36191 (N_36191,N_35666,N_35584);
nor U36192 (N_36192,N_35764,N_35854);
nand U36193 (N_36193,N_35554,N_35826);
xnor U36194 (N_36194,N_35924,N_35528);
nor U36195 (N_36195,N_35950,N_35805);
nor U36196 (N_36196,N_35587,N_35960);
or U36197 (N_36197,N_35680,N_35928);
nand U36198 (N_36198,N_35650,N_35612);
nand U36199 (N_36199,N_35750,N_35797);
nor U36200 (N_36200,N_35744,N_35975);
xor U36201 (N_36201,N_35634,N_35662);
and U36202 (N_36202,N_35777,N_35932);
and U36203 (N_36203,N_35749,N_35521);
and U36204 (N_36204,N_35862,N_35986);
nand U36205 (N_36205,N_35737,N_35539);
xnor U36206 (N_36206,N_35572,N_35888);
or U36207 (N_36207,N_35743,N_35846);
and U36208 (N_36208,N_35941,N_35619);
or U36209 (N_36209,N_35980,N_35949);
nor U36210 (N_36210,N_35979,N_35688);
or U36211 (N_36211,N_35838,N_35569);
xnor U36212 (N_36212,N_35535,N_35679);
nor U36213 (N_36213,N_35848,N_35874);
nor U36214 (N_36214,N_35784,N_35592);
nor U36215 (N_36215,N_35710,N_35731);
or U36216 (N_36216,N_35808,N_35566);
nor U36217 (N_36217,N_35845,N_35807);
nor U36218 (N_36218,N_35996,N_35885);
nor U36219 (N_36219,N_35801,N_35586);
nand U36220 (N_36220,N_35812,N_35551);
nor U36221 (N_36221,N_35773,N_35574);
and U36222 (N_36222,N_35988,N_35639);
nor U36223 (N_36223,N_35696,N_35802);
and U36224 (N_36224,N_35999,N_35981);
nor U36225 (N_36225,N_35632,N_35860);
nor U36226 (N_36226,N_35508,N_35638);
or U36227 (N_36227,N_35608,N_35590);
or U36228 (N_36228,N_35667,N_35735);
nor U36229 (N_36229,N_35533,N_35600);
or U36230 (N_36230,N_35832,N_35685);
nand U36231 (N_36231,N_35893,N_35898);
or U36232 (N_36232,N_35556,N_35818);
or U36233 (N_36233,N_35618,N_35654);
or U36234 (N_36234,N_35687,N_35828);
nor U36235 (N_36235,N_35665,N_35809);
nand U36236 (N_36236,N_35580,N_35649);
or U36237 (N_36237,N_35568,N_35597);
nand U36238 (N_36238,N_35712,N_35751);
nand U36239 (N_36239,N_35548,N_35505);
nor U36240 (N_36240,N_35989,N_35707);
nand U36241 (N_36241,N_35819,N_35915);
xor U36242 (N_36242,N_35661,N_35610);
or U36243 (N_36243,N_35921,N_35920);
nor U36244 (N_36244,N_35698,N_35658);
nand U36245 (N_36245,N_35968,N_35842);
or U36246 (N_36246,N_35992,N_35925);
xor U36247 (N_36247,N_35831,N_35804);
and U36248 (N_36248,N_35682,N_35591);
nand U36249 (N_36249,N_35657,N_35629);
nand U36250 (N_36250,N_35995,N_35979);
or U36251 (N_36251,N_35554,N_35926);
or U36252 (N_36252,N_35766,N_35545);
and U36253 (N_36253,N_35676,N_35840);
or U36254 (N_36254,N_35841,N_35850);
xnor U36255 (N_36255,N_35825,N_35833);
or U36256 (N_36256,N_35894,N_35518);
nand U36257 (N_36257,N_35669,N_35662);
xor U36258 (N_36258,N_35670,N_35981);
and U36259 (N_36259,N_35622,N_35782);
or U36260 (N_36260,N_35601,N_35783);
and U36261 (N_36261,N_35835,N_35870);
nor U36262 (N_36262,N_35514,N_35841);
or U36263 (N_36263,N_35798,N_35544);
xor U36264 (N_36264,N_35934,N_35815);
nor U36265 (N_36265,N_35692,N_35593);
nand U36266 (N_36266,N_35884,N_35974);
nor U36267 (N_36267,N_35599,N_35953);
nand U36268 (N_36268,N_35551,N_35861);
and U36269 (N_36269,N_35978,N_35675);
nor U36270 (N_36270,N_35701,N_35567);
nand U36271 (N_36271,N_35552,N_35781);
nand U36272 (N_36272,N_35618,N_35511);
and U36273 (N_36273,N_35645,N_35671);
xnor U36274 (N_36274,N_35702,N_35657);
nor U36275 (N_36275,N_35747,N_35899);
and U36276 (N_36276,N_35650,N_35786);
nand U36277 (N_36277,N_35549,N_35512);
nor U36278 (N_36278,N_35987,N_35813);
and U36279 (N_36279,N_35631,N_35761);
nand U36280 (N_36280,N_35970,N_35729);
and U36281 (N_36281,N_35546,N_35551);
and U36282 (N_36282,N_35915,N_35834);
or U36283 (N_36283,N_35942,N_35666);
nand U36284 (N_36284,N_35778,N_35925);
and U36285 (N_36285,N_35770,N_35726);
nand U36286 (N_36286,N_35851,N_35672);
nor U36287 (N_36287,N_35863,N_35820);
nor U36288 (N_36288,N_35762,N_35546);
nor U36289 (N_36289,N_35895,N_35557);
nor U36290 (N_36290,N_35592,N_35509);
or U36291 (N_36291,N_35796,N_35835);
and U36292 (N_36292,N_35813,N_35904);
nand U36293 (N_36293,N_35926,N_35933);
and U36294 (N_36294,N_35571,N_35929);
nor U36295 (N_36295,N_35844,N_35630);
or U36296 (N_36296,N_35726,N_35537);
nand U36297 (N_36297,N_35980,N_35863);
and U36298 (N_36298,N_35902,N_35867);
nand U36299 (N_36299,N_35731,N_35541);
and U36300 (N_36300,N_35858,N_35904);
nor U36301 (N_36301,N_35644,N_35757);
nor U36302 (N_36302,N_35814,N_35658);
and U36303 (N_36303,N_35690,N_35572);
or U36304 (N_36304,N_35991,N_35738);
and U36305 (N_36305,N_35685,N_35874);
and U36306 (N_36306,N_35765,N_35716);
or U36307 (N_36307,N_35888,N_35815);
or U36308 (N_36308,N_35547,N_35622);
and U36309 (N_36309,N_35892,N_35896);
or U36310 (N_36310,N_35707,N_35534);
or U36311 (N_36311,N_35925,N_35761);
nand U36312 (N_36312,N_35721,N_35867);
and U36313 (N_36313,N_35835,N_35623);
or U36314 (N_36314,N_35826,N_35896);
or U36315 (N_36315,N_35809,N_35843);
nor U36316 (N_36316,N_35785,N_35957);
xor U36317 (N_36317,N_35642,N_35622);
nand U36318 (N_36318,N_35694,N_35943);
and U36319 (N_36319,N_35605,N_35842);
xnor U36320 (N_36320,N_35544,N_35667);
nand U36321 (N_36321,N_35778,N_35890);
and U36322 (N_36322,N_35922,N_35645);
or U36323 (N_36323,N_35807,N_35618);
nand U36324 (N_36324,N_35916,N_35819);
or U36325 (N_36325,N_35935,N_35696);
nand U36326 (N_36326,N_35877,N_35757);
xor U36327 (N_36327,N_35677,N_35839);
nor U36328 (N_36328,N_35976,N_35982);
or U36329 (N_36329,N_35544,N_35576);
xnor U36330 (N_36330,N_35958,N_35860);
and U36331 (N_36331,N_35669,N_35816);
nand U36332 (N_36332,N_35624,N_35600);
xnor U36333 (N_36333,N_35944,N_35933);
or U36334 (N_36334,N_35789,N_35661);
nand U36335 (N_36335,N_35809,N_35620);
or U36336 (N_36336,N_35997,N_35753);
and U36337 (N_36337,N_35840,N_35628);
nor U36338 (N_36338,N_35718,N_35504);
and U36339 (N_36339,N_35729,N_35687);
nand U36340 (N_36340,N_35692,N_35567);
nand U36341 (N_36341,N_35680,N_35766);
nand U36342 (N_36342,N_35666,N_35790);
nand U36343 (N_36343,N_35544,N_35795);
nor U36344 (N_36344,N_35875,N_35789);
nor U36345 (N_36345,N_35945,N_35809);
xnor U36346 (N_36346,N_35635,N_35627);
and U36347 (N_36347,N_35701,N_35846);
nand U36348 (N_36348,N_35520,N_35994);
or U36349 (N_36349,N_35879,N_35882);
nor U36350 (N_36350,N_35983,N_35949);
and U36351 (N_36351,N_35619,N_35714);
nor U36352 (N_36352,N_35936,N_35609);
or U36353 (N_36353,N_35622,N_35596);
xnor U36354 (N_36354,N_35656,N_35852);
nor U36355 (N_36355,N_35504,N_35698);
and U36356 (N_36356,N_35621,N_35811);
and U36357 (N_36357,N_35847,N_35637);
nor U36358 (N_36358,N_35630,N_35720);
nand U36359 (N_36359,N_35905,N_35902);
xnor U36360 (N_36360,N_35964,N_35682);
and U36361 (N_36361,N_35515,N_35868);
or U36362 (N_36362,N_35757,N_35516);
or U36363 (N_36363,N_35735,N_35528);
nand U36364 (N_36364,N_35608,N_35678);
or U36365 (N_36365,N_35920,N_35669);
and U36366 (N_36366,N_35735,N_35763);
nor U36367 (N_36367,N_35816,N_35915);
and U36368 (N_36368,N_35708,N_35767);
or U36369 (N_36369,N_35624,N_35521);
and U36370 (N_36370,N_35769,N_35992);
or U36371 (N_36371,N_35778,N_35749);
or U36372 (N_36372,N_35538,N_35708);
nor U36373 (N_36373,N_35622,N_35789);
nor U36374 (N_36374,N_35734,N_35956);
xor U36375 (N_36375,N_35639,N_35803);
nand U36376 (N_36376,N_35931,N_35885);
nand U36377 (N_36377,N_35957,N_35953);
nand U36378 (N_36378,N_35763,N_35724);
and U36379 (N_36379,N_35902,N_35643);
and U36380 (N_36380,N_35658,N_35883);
or U36381 (N_36381,N_35956,N_35525);
or U36382 (N_36382,N_35866,N_35876);
nand U36383 (N_36383,N_35719,N_35895);
or U36384 (N_36384,N_35921,N_35568);
and U36385 (N_36385,N_35828,N_35536);
nor U36386 (N_36386,N_35946,N_35653);
and U36387 (N_36387,N_35918,N_35852);
or U36388 (N_36388,N_35920,N_35838);
nand U36389 (N_36389,N_35562,N_35962);
xnor U36390 (N_36390,N_35577,N_35787);
nand U36391 (N_36391,N_35954,N_35641);
and U36392 (N_36392,N_35573,N_35907);
nand U36393 (N_36393,N_35790,N_35966);
or U36394 (N_36394,N_35514,N_35653);
or U36395 (N_36395,N_35560,N_35613);
and U36396 (N_36396,N_35868,N_35701);
and U36397 (N_36397,N_35952,N_35663);
or U36398 (N_36398,N_35800,N_35778);
or U36399 (N_36399,N_35578,N_35846);
or U36400 (N_36400,N_35909,N_35629);
nand U36401 (N_36401,N_35817,N_35750);
nand U36402 (N_36402,N_35992,N_35606);
or U36403 (N_36403,N_35761,N_35863);
xor U36404 (N_36404,N_35987,N_35899);
nor U36405 (N_36405,N_35673,N_35727);
xnor U36406 (N_36406,N_35665,N_35874);
nor U36407 (N_36407,N_35547,N_35986);
nand U36408 (N_36408,N_35905,N_35827);
xor U36409 (N_36409,N_35935,N_35812);
or U36410 (N_36410,N_35891,N_35609);
nand U36411 (N_36411,N_35793,N_35732);
nand U36412 (N_36412,N_35619,N_35883);
or U36413 (N_36413,N_35967,N_35770);
and U36414 (N_36414,N_35781,N_35895);
or U36415 (N_36415,N_35884,N_35726);
xnor U36416 (N_36416,N_35554,N_35954);
and U36417 (N_36417,N_35563,N_35970);
and U36418 (N_36418,N_35801,N_35507);
nand U36419 (N_36419,N_35641,N_35934);
nand U36420 (N_36420,N_35527,N_35644);
and U36421 (N_36421,N_35958,N_35789);
and U36422 (N_36422,N_35905,N_35864);
nor U36423 (N_36423,N_35864,N_35942);
and U36424 (N_36424,N_35929,N_35871);
nor U36425 (N_36425,N_35619,N_35983);
and U36426 (N_36426,N_35563,N_35652);
nand U36427 (N_36427,N_35647,N_35954);
nand U36428 (N_36428,N_35785,N_35650);
nand U36429 (N_36429,N_35574,N_35593);
or U36430 (N_36430,N_35593,N_35583);
and U36431 (N_36431,N_35557,N_35879);
nor U36432 (N_36432,N_35615,N_35926);
nand U36433 (N_36433,N_35852,N_35760);
nor U36434 (N_36434,N_35960,N_35925);
nor U36435 (N_36435,N_35803,N_35815);
and U36436 (N_36436,N_35885,N_35737);
nor U36437 (N_36437,N_35849,N_35837);
xnor U36438 (N_36438,N_35522,N_35609);
and U36439 (N_36439,N_35871,N_35942);
and U36440 (N_36440,N_35513,N_35501);
xor U36441 (N_36441,N_35687,N_35787);
nor U36442 (N_36442,N_35941,N_35688);
nor U36443 (N_36443,N_35533,N_35983);
and U36444 (N_36444,N_35735,N_35982);
nor U36445 (N_36445,N_35990,N_35567);
nor U36446 (N_36446,N_35646,N_35533);
nor U36447 (N_36447,N_35505,N_35659);
or U36448 (N_36448,N_35617,N_35523);
nand U36449 (N_36449,N_35823,N_35840);
and U36450 (N_36450,N_35791,N_35891);
and U36451 (N_36451,N_35686,N_35846);
or U36452 (N_36452,N_35615,N_35733);
nor U36453 (N_36453,N_35989,N_35664);
nor U36454 (N_36454,N_35902,N_35607);
nor U36455 (N_36455,N_35523,N_35884);
or U36456 (N_36456,N_35863,N_35849);
xor U36457 (N_36457,N_35531,N_35658);
or U36458 (N_36458,N_35918,N_35529);
xor U36459 (N_36459,N_35961,N_35849);
nor U36460 (N_36460,N_35985,N_35881);
nor U36461 (N_36461,N_35894,N_35843);
or U36462 (N_36462,N_35626,N_35989);
nor U36463 (N_36463,N_35777,N_35694);
nand U36464 (N_36464,N_35788,N_35834);
xnor U36465 (N_36465,N_35685,N_35527);
or U36466 (N_36466,N_35554,N_35702);
and U36467 (N_36467,N_35731,N_35600);
nor U36468 (N_36468,N_35937,N_35906);
and U36469 (N_36469,N_35506,N_35654);
nand U36470 (N_36470,N_35500,N_35668);
nand U36471 (N_36471,N_35680,N_35825);
nor U36472 (N_36472,N_35568,N_35904);
and U36473 (N_36473,N_35652,N_35938);
and U36474 (N_36474,N_35566,N_35978);
xor U36475 (N_36475,N_35854,N_35832);
or U36476 (N_36476,N_35917,N_35735);
and U36477 (N_36477,N_35814,N_35529);
and U36478 (N_36478,N_35638,N_35897);
nand U36479 (N_36479,N_35578,N_35658);
nor U36480 (N_36480,N_35518,N_35743);
nor U36481 (N_36481,N_35880,N_35701);
xnor U36482 (N_36482,N_35932,N_35870);
xor U36483 (N_36483,N_35719,N_35981);
nor U36484 (N_36484,N_35524,N_35780);
xor U36485 (N_36485,N_35791,N_35522);
nand U36486 (N_36486,N_35680,N_35962);
nand U36487 (N_36487,N_35709,N_35567);
or U36488 (N_36488,N_35766,N_35716);
xor U36489 (N_36489,N_35594,N_35712);
xor U36490 (N_36490,N_35581,N_35712);
or U36491 (N_36491,N_35987,N_35903);
or U36492 (N_36492,N_35999,N_35855);
and U36493 (N_36493,N_35970,N_35635);
and U36494 (N_36494,N_35902,N_35616);
nor U36495 (N_36495,N_35811,N_35792);
xnor U36496 (N_36496,N_35592,N_35581);
or U36497 (N_36497,N_35501,N_35945);
xnor U36498 (N_36498,N_35568,N_35641);
nand U36499 (N_36499,N_35539,N_35533);
nor U36500 (N_36500,N_36492,N_36131);
or U36501 (N_36501,N_36379,N_36347);
xor U36502 (N_36502,N_36285,N_36461);
nand U36503 (N_36503,N_36414,N_36313);
nand U36504 (N_36504,N_36489,N_36399);
or U36505 (N_36505,N_36188,N_36151);
or U36506 (N_36506,N_36137,N_36231);
and U36507 (N_36507,N_36145,N_36040);
nor U36508 (N_36508,N_36247,N_36423);
or U36509 (N_36509,N_36445,N_36368);
or U36510 (N_36510,N_36475,N_36408);
or U36511 (N_36511,N_36012,N_36404);
nor U36512 (N_36512,N_36187,N_36350);
or U36513 (N_36513,N_36225,N_36339);
xnor U36514 (N_36514,N_36364,N_36221);
or U36515 (N_36515,N_36323,N_36232);
and U36516 (N_36516,N_36165,N_36054);
xor U36517 (N_36517,N_36147,N_36381);
nand U36518 (N_36518,N_36268,N_36245);
nand U36519 (N_36519,N_36412,N_36395);
xnor U36520 (N_36520,N_36069,N_36214);
nor U36521 (N_36521,N_36167,N_36374);
xor U36522 (N_36522,N_36371,N_36393);
nor U36523 (N_36523,N_36209,N_36417);
nor U36524 (N_36524,N_36171,N_36019);
nand U36525 (N_36525,N_36181,N_36168);
xor U36526 (N_36526,N_36169,N_36306);
nand U36527 (N_36527,N_36474,N_36483);
or U36528 (N_36528,N_36104,N_36139);
nor U36529 (N_36529,N_36159,N_36194);
or U36530 (N_36530,N_36071,N_36200);
nand U36531 (N_36531,N_36222,N_36266);
and U36532 (N_36532,N_36466,N_36327);
or U36533 (N_36533,N_36416,N_36411);
nor U36534 (N_36534,N_36198,N_36084);
and U36535 (N_36535,N_36119,N_36065);
nor U36536 (N_36536,N_36383,N_36469);
or U36537 (N_36537,N_36025,N_36080);
and U36538 (N_36538,N_36047,N_36264);
or U36539 (N_36539,N_36287,N_36237);
nand U36540 (N_36540,N_36488,N_36108);
or U36541 (N_36541,N_36004,N_36079);
nor U36542 (N_36542,N_36008,N_36128);
nand U36543 (N_36543,N_36360,N_36230);
nor U36544 (N_36544,N_36367,N_36491);
or U36545 (N_36545,N_36369,N_36366);
nand U36546 (N_36546,N_36096,N_36238);
nor U36547 (N_36547,N_36068,N_36303);
nand U36548 (N_36548,N_36044,N_36278);
nand U36549 (N_36549,N_36038,N_36111);
and U36550 (N_36550,N_36223,N_36090);
xnor U36551 (N_36551,N_36336,N_36456);
and U36552 (N_36552,N_36149,N_36267);
nor U36553 (N_36553,N_36280,N_36075);
and U36554 (N_36554,N_36311,N_36122);
nor U36555 (N_36555,N_36333,N_36319);
and U36556 (N_36556,N_36471,N_36452);
nor U36557 (N_36557,N_36190,N_36256);
nor U36558 (N_36558,N_36255,N_36195);
xor U36559 (N_36559,N_36284,N_36130);
nand U36560 (N_36560,N_36449,N_36430);
or U36561 (N_36561,N_36252,N_36121);
or U36562 (N_36562,N_36039,N_36402);
and U36563 (N_36563,N_36477,N_36113);
and U36564 (N_36564,N_36372,N_36192);
or U36565 (N_36565,N_36403,N_36175);
and U36566 (N_36566,N_36353,N_36028);
or U36567 (N_36567,N_36196,N_36386);
and U36568 (N_36568,N_36010,N_36308);
nand U36569 (N_36569,N_36193,N_36092);
and U36570 (N_36570,N_36472,N_36027);
and U36571 (N_36571,N_36265,N_36493);
nor U36572 (N_36572,N_36435,N_36453);
nor U36573 (N_36573,N_36217,N_36447);
nand U36574 (N_36574,N_36455,N_36468);
or U36575 (N_36575,N_36085,N_36126);
or U36576 (N_36576,N_36338,N_36304);
xnor U36577 (N_36577,N_36021,N_36272);
nor U36578 (N_36578,N_36114,N_36076);
nand U36579 (N_36579,N_36312,N_36301);
nand U36580 (N_36580,N_36166,N_36117);
nand U36581 (N_36581,N_36003,N_36398);
xor U36582 (N_36582,N_36129,N_36275);
and U36583 (N_36583,N_36426,N_36061);
and U36584 (N_36584,N_36227,N_36125);
and U36585 (N_36585,N_36315,N_36201);
nand U36586 (N_36586,N_36332,N_36026);
nor U36587 (N_36587,N_36391,N_36116);
or U36588 (N_36588,N_36378,N_36156);
nor U36589 (N_36589,N_36006,N_36329);
and U36590 (N_36590,N_36377,N_36174);
nand U36591 (N_36591,N_36286,N_36011);
nor U36592 (N_36592,N_36279,N_36320);
nor U36593 (N_36593,N_36425,N_36127);
xor U36594 (N_36594,N_36486,N_36224);
and U36595 (N_36595,N_36354,N_36326);
nand U36596 (N_36596,N_36334,N_36219);
xor U36597 (N_36597,N_36148,N_36042);
nor U36598 (N_36598,N_36433,N_36001);
or U36599 (N_36599,N_36294,N_36482);
xnor U36600 (N_36600,N_36300,N_36182);
nand U36601 (N_36601,N_36093,N_36299);
nor U36602 (N_36602,N_36462,N_36056);
nor U36603 (N_36603,N_36115,N_36322);
nand U36604 (N_36604,N_36205,N_36218);
xor U36605 (N_36605,N_36380,N_36282);
nor U36606 (N_36606,N_36152,N_36109);
nor U36607 (N_36607,N_36390,N_36053);
or U36608 (N_36608,N_36259,N_36409);
and U36609 (N_36609,N_36202,N_36173);
or U36610 (N_36610,N_36153,N_36438);
nand U36611 (N_36611,N_36178,N_36496);
xor U36612 (N_36612,N_36233,N_36197);
xnor U36613 (N_36613,N_36176,N_36242);
and U36614 (N_36614,N_36274,N_36249);
nor U36615 (N_36615,N_36094,N_36144);
nand U36616 (N_36616,N_36234,N_36022);
nand U36617 (N_36617,N_36066,N_36018);
nor U36618 (N_36618,N_36376,N_36045);
nor U36619 (N_36619,N_36133,N_36289);
nor U36620 (N_36620,N_36446,N_36213);
nor U36621 (N_36621,N_36363,N_36046);
and U36622 (N_36622,N_36273,N_36292);
nand U36623 (N_36623,N_36296,N_36002);
or U36624 (N_36624,N_36321,N_36077);
and U36625 (N_36625,N_36101,N_36310);
or U36626 (N_36626,N_36024,N_36208);
nand U36627 (N_36627,N_36087,N_36494);
and U36628 (N_36628,N_36465,N_36450);
nand U36629 (N_36629,N_36457,N_36244);
or U36630 (N_36630,N_36100,N_36162);
or U36631 (N_36631,N_36210,N_36072);
and U36632 (N_36632,N_36269,N_36330);
nor U36633 (N_36633,N_36184,N_36436);
nor U36634 (N_36634,N_36032,N_36307);
nor U36635 (N_36635,N_36388,N_36142);
nor U36636 (N_36636,N_36443,N_36120);
and U36637 (N_36637,N_36070,N_36016);
nand U36638 (N_36638,N_36052,N_36155);
nor U36639 (N_36639,N_36358,N_36207);
and U36640 (N_36640,N_36460,N_36023);
nor U36641 (N_36641,N_36355,N_36083);
nor U36642 (N_36642,N_36324,N_36241);
and U36643 (N_36643,N_36017,N_36211);
or U36644 (N_36644,N_36497,N_36110);
or U36645 (N_36645,N_36318,N_36464);
nand U36646 (N_36646,N_36373,N_36473);
and U36647 (N_36647,N_36146,N_36103);
and U36648 (N_36648,N_36365,N_36243);
nor U36649 (N_36649,N_36035,N_36419);
or U36650 (N_36650,N_36470,N_36031);
nand U36651 (N_36651,N_36328,N_36410);
nor U36652 (N_36652,N_36226,N_36432);
nor U36653 (N_36653,N_36490,N_36009);
or U36654 (N_36654,N_36257,N_36246);
or U36655 (N_36655,N_36451,N_36078);
nand U36656 (N_36656,N_36458,N_36135);
and U36657 (N_36657,N_36160,N_36191);
nand U36658 (N_36658,N_36479,N_36123);
or U36659 (N_36659,N_36206,N_36033);
nor U36660 (N_36660,N_36005,N_36351);
and U36661 (N_36661,N_36041,N_36424);
and U36662 (N_36662,N_36389,N_36034);
or U36663 (N_36663,N_36480,N_36349);
nand U36664 (N_36664,N_36189,N_36098);
or U36665 (N_36665,N_36014,N_36401);
or U36666 (N_36666,N_36060,N_36013);
nand U36667 (N_36667,N_36420,N_36050);
or U36668 (N_36668,N_36406,N_36442);
nor U36669 (N_36669,N_36281,N_36260);
and U36670 (N_36670,N_36112,N_36143);
and U36671 (N_36671,N_36236,N_36164);
or U36672 (N_36672,N_36343,N_36258);
and U36673 (N_36673,N_36212,N_36362);
or U36674 (N_36674,N_36440,N_36463);
or U36675 (N_36675,N_36089,N_36150);
nand U36676 (N_36676,N_36158,N_36172);
and U36677 (N_36677,N_36356,N_36185);
nor U36678 (N_36678,N_36276,N_36251);
and U36679 (N_36679,N_36297,N_36495);
or U36680 (N_36680,N_36270,N_36074);
nor U36681 (N_36681,N_36239,N_36263);
or U36682 (N_36682,N_36478,N_36295);
nor U36683 (N_36683,N_36049,N_36124);
xnor U36684 (N_36684,N_36394,N_36291);
xor U36685 (N_36685,N_36439,N_36203);
or U36686 (N_36686,N_36067,N_36062);
and U36687 (N_36687,N_36082,N_36361);
nor U36688 (N_36688,N_36317,N_36298);
and U36689 (N_36689,N_36170,N_36359);
nor U36690 (N_36690,N_36341,N_36385);
xor U36691 (N_36691,N_36498,N_36413);
nor U36692 (N_36692,N_36015,N_36370);
xnor U36693 (N_36693,N_36254,N_36397);
nor U36694 (N_36694,N_36396,N_36064);
and U36695 (N_36695,N_36407,N_36086);
nand U36696 (N_36696,N_36487,N_36037);
nand U36697 (N_36697,N_36309,N_36102);
xnor U36698 (N_36698,N_36020,N_36000);
nor U36699 (N_36699,N_36387,N_36138);
and U36700 (N_36700,N_36421,N_36346);
nor U36701 (N_36701,N_36283,N_36325);
nand U36702 (N_36702,N_36476,N_36136);
and U36703 (N_36703,N_36204,N_36342);
nand U36704 (N_36704,N_36099,N_36029);
nand U36705 (N_36705,N_36337,N_36097);
nor U36706 (N_36706,N_36186,N_36180);
nor U36707 (N_36707,N_36448,N_36248);
nand U36708 (N_36708,N_36467,N_36441);
and U36709 (N_36709,N_36405,N_36088);
nand U36710 (N_36710,N_36216,N_36392);
nand U36711 (N_36711,N_36352,N_36059);
xor U36712 (N_36712,N_36434,N_36277);
or U36713 (N_36713,N_36177,N_36454);
and U36714 (N_36714,N_36481,N_36427);
nor U36715 (N_36715,N_36007,N_36345);
and U36716 (N_36716,N_36063,N_36107);
nor U36717 (N_36717,N_36459,N_36140);
xor U36718 (N_36718,N_36081,N_36288);
xor U36719 (N_36719,N_36428,N_36235);
and U36720 (N_36720,N_36199,N_36485);
nand U36721 (N_36721,N_36400,N_36240);
nor U36722 (N_36722,N_36384,N_36179);
and U36723 (N_36723,N_36073,N_36431);
and U36724 (N_36724,N_36271,N_36183);
nand U36725 (N_36725,N_36444,N_36091);
nor U36726 (N_36726,N_36141,N_36132);
xnor U36727 (N_36727,N_36302,N_36422);
xnor U36728 (N_36728,N_36105,N_36030);
nand U36729 (N_36729,N_36118,N_36344);
nand U36730 (N_36730,N_36228,N_36043);
or U36731 (N_36731,N_36484,N_36290);
nand U36732 (N_36732,N_36375,N_36415);
nand U36733 (N_36733,N_36154,N_36229);
and U36734 (N_36734,N_36262,N_36357);
and U36735 (N_36735,N_36253,N_36499);
or U36736 (N_36736,N_36293,N_36305);
or U36737 (N_36737,N_36250,N_36220);
and U36738 (N_36738,N_36418,N_36036);
nand U36739 (N_36739,N_36055,N_36348);
or U36740 (N_36740,N_36157,N_36134);
or U36741 (N_36741,N_36163,N_36051);
nor U36742 (N_36742,N_36340,N_36048);
nand U36743 (N_36743,N_36429,N_36261);
or U36744 (N_36744,N_36382,N_36331);
or U36745 (N_36745,N_36335,N_36058);
nor U36746 (N_36746,N_36161,N_36057);
or U36747 (N_36747,N_36316,N_36095);
nand U36748 (N_36748,N_36437,N_36314);
xor U36749 (N_36749,N_36106,N_36215);
nand U36750 (N_36750,N_36365,N_36393);
nand U36751 (N_36751,N_36137,N_36306);
nand U36752 (N_36752,N_36049,N_36453);
or U36753 (N_36753,N_36021,N_36105);
nand U36754 (N_36754,N_36127,N_36456);
and U36755 (N_36755,N_36332,N_36086);
or U36756 (N_36756,N_36228,N_36422);
and U36757 (N_36757,N_36333,N_36377);
or U36758 (N_36758,N_36081,N_36233);
or U36759 (N_36759,N_36066,N_36014);
or U36760 (N_36760,N_36216,N_36331);
or U36761 (N_36761,N_36427,N_36322);
nand U36762 (N_36762,N_36310,N_36151);
and U36763 (N_36763,N_36169,N_36393);
nor U36764 (N_36764,N_36402,N_36116);
xor U36765 (N_36765,N_36066,N_36015);
nor U36766 (N_36766,N_36273,N_36379);
nand U36767 (N_36767,N_36302,N_36186);
and U36768 (N_36768,N_36135,N_36425);
and U36769 (N_36769,N_36499,N_36409);
and U36770 (N_36770,N_36106,N_36279);
and U36771 (N_36771,N_36303,N_36113);
nand U36772 (N_36772,N_36478,N_36270);
nor U36773 (N_36773,N_36389,N_36172);
or U36774 (N_36774,N_36407,N_36045);
or U36775 (N_36775,N_36434,N_36482);
and U36776 (N_36776,N_36403,N_36440);
nand U36777 (N_36777,N_36391,N_36244);
nor U36778 (N_36778,N_36462,N_36322);
nand U36779 (N_36779,N_36378,N_36314);
xor U36780 (N_36780,N_36201,N_36464);
nand U36781 (N_36781,N_36494,N_36364);
or U36782 (N_36782,N_36417,N_36021);
nor U36783 (N_36783,N_36142,N_36109);
nand U36784 (N_36784,N_36262,N_36056);
nor U36785 (N_36785,N_36350,N_36063);
xor U36786 (N_36786,N_36425,N_36393);
or U36787 (N_36787,N_36248,N_36019);
nor U36788 (N_36788,N_36026,N_36274);
or U36789 (N_36789,N_36171,N_36459);
and U36790 (N_36790,N_36424,N_36258);
xor U36791 (N_36791,N_36457,N_36173);
nor U36792 (N_36792,N_36357,N_36188);
nand U36793 (N_36793,N_36055,N_36276);
nor U36794 (N_36794,N_36343,N_36005);
nor U36795 (N_36795,N_36354,N_36301);
nand U36796 (N_36796,N_36109,N_36069);
nor U36797 (N_36797,N_36232,N_36118);
or U36798 (N_36798,N_36394,N_36344);
nor U36799 (N_36799,N_36115,N_36159);
nor U36800 (N_36800,N_36481,N_36470);
nor U36801 (N_36801,N_36412,N_36289);
xor U36802 (N_36802,N_36138,N_36061);
nor U36803 (N_36803,N_36209,N_36344);
nand U36804 (N_36804,N_36019,N_36339);
nand U36805 (N_36805,N_36437,N_36405);
nand U36806 (N_36806,N_36224,N_36366);
xnor U36807 (N_36807,N_36059,N_36457);
nand U36808 (N_36808,N_36010,N_36136);
and U36809 (N_36809,N_36460,N_36369);
and U36810 (N_36810,N_36242,N_36395);
xnor U36811 (N_36811,N_36193,N_36198);
or U36812 (N_36812,N_36447,N_36287);
nor U36813 (N_36813,N_36269,N_36184);
nor U36814 (N_36814,N_36330,N_36456);
nor U36815 (N_36815,N_36027,N_36445);
xor U36816 (N_36816,N_36395,N_36231);
nor U36817 (N_36817,N_36102,N_36301);
nand U36818 (N_36818,N_36387,N_36020);
or U36819 (N_36819,N_36300,N_36011);
nand U36820 (N_36820,N_36317,N_36432);
nor U36821 (N_36821,N_36180,N_36071);
and U36822 (N_36822,N_36111,N_36240);
and U36823 (N_36823,N_36349,N_36390);
and U36824 (N_36824,N_36329,N_36102);
nand U36825 (N_36825,N_36499,N_36300);
nor U36826 (N_36826,N_36006,N_36170);
nor U36827 (N_36827,N_36301,N_36472);
or U36828 (N_36828,N_36147,N_36214);
nand U36829 (N_36829,N_36286,N_36178);
or U36830 (N_36830,N_36024,N_36186);
and U36831 (N_36831,N_36414,N_36450);
xnor U36832 (N_36832,N_36015,N_36295);
nand U36833 (N_36833,N_36254,N_36460);
xnor U36834 (N_36834,N_36474,N_36040);
nand U36835 (N_36835,N_36454,N_36329);
nor U36836 (N_36836,N_36113,N_36127);
and U36837 (N_36837,N_36482,N_36249);
nand U36838 (N_36838,N_36378,N_36146);
xor U36839 (N_36839,N_36356,N_36389);
nor U36840 (N_36840,N_36086,N_36459);
nor U36841 (N_36841,N_36261,N_36229);
nor U36842 (N_36842,N_36241,N_36327);
xnor U36843 (N_36843,N_36261,N_36111);
or U36844 (N_36844,N_36361,N_36451);
nand U36845 (N_36845,N_36375,N_36205);
xnor U36846 (N_36846,N_36137,N_36187);
nor U36847 (N_36847,N_36092,N_36156);
nand U36848 (N_36848,N_36311,N_36433);
nor U36849 (N_36849,N_36234,N_36157);
and U36850 (N_36850,N_36382,N_36131);
and U36851 (N_36851,N_36233,N_36405);
or U36852 (N_36852,N_36021,N_36070);
nand U36853 (N_36853,N_36049,N_36130);
xnor U36854 (N_36854,N_36131,N_36299);
nand U36855 (N_36855,N_36044,N_36071);
nand U36856 (N_36856,N_36485,N_36099);
xnor U36857 (N_36857,N_36161,N_36251);
nand U36858 (N_36858,N_36026,N_36472);
nor U36859 (N_36859,N_36467,N_36440);
nor U36860 (N_36860,N_36373,N_36108);
and U36861 (N_36861,N_36496,N_36424);
or U36862 (N_36862,N_36065,N_36188);
nor U36863 (N_36863,N_36106,N_36298);
or U36864 (N_36864,N_36488,N_36341);
or U36865 (N_36865,N_36382,N_36168);
or U36866 (N_36866,N_36291,N_36369);
nor U36867 (N_36867,N_36418,N_36174);
or U36868 (N_36868,N_36068,N_36417);
and U36869 (N_36869,N_36155,N_36469);
nand U36870 (N_36870,N_36301,N_36443);
and U36871 (N_36871,N_36082,N_36376);
xor U36872 (N_36872,N_36361,N_36248);
and U36873 (N_36873,N_36298,N_36487);
or U36874 (N_36874,N_36015,N_36094);
nand U36875 (N_36875,N_36313,N_36015);
and U36876 (N_36876,N_36232,N_36405);
nor U36877 (N_36877,N_36117,N_36317);
and U36878 (N_36878,N_36421,N_36290);
nand U36879 (N_36879,N_36027,N_36350);
nand U36880 (N_36880,N_36213,N_36168);
or U36881 (N_36881,N_36144,N_36049);
nor U36882 (N_36882,N_36446,N_36410);
nor U36883 (N_36883,N_36258,N_36038);
and U36884 (N_36884,N_36028,N_36181);
nand U36885 (N_36885,N_36392,N_36044);
xnor U36886 (N_36886,N_36355,N_36062);
nor U36887 (N_36887,N_36156,N_36196);
xor U36888 (N_36888,N_36101,N_36298);
nand U36889 (N_36889,N_36372,N_36321);
xnor U36890 (N_36890,N_36243,N_36018);
or U36891 (N_36891,N_36271,N_36021);
and U36892 (N_36892,N_36257,N_36199);
and U36893 (N_36893,N_36129,N_36083);
and U36894 (N_36894,N_36140,N_36292);
and U36895 (N_36895,N_36262,N_36321);
nor U36896 (N_36896,N_36464,N_36128);
nor U36897 (N_36897,N_36270,N_36427);
or U36898 (N_36898,N_36403,N_36415);
nor U36899 (N_36899,N_36046,N_36113);
or U36900 (N_36900,N_36440,N_36364);
or U36901 (N_36901,N_36173,N_36498);
xor U36902 (N_36902,N_36411,N_36331);
or U36903 (N_36903,N_36190,N_36485);
or U36904 (N_36904,N_36318,N_36487);
nor U36905 (N_36905,N_36233,N_36316);
xnor U36906 (N_36906,N_36227,N_36191);
nor U36907 (N_36907,N_36078,N_36051);
nand U36908 (N_36908,N_36190,N_36427);
and U36909 (N_36909,N_36394,N_36098);
and U36910 (N_36910,N_36100,N_36183);
xnor U36911 (N_36911,N_36134,N_36405);
nand U36912 (N_36912,N_36390,N_36032);
nand U36913 (N_36913,N_36170,N_36255);
nand U36914 (N_36914,N_36497,N_36313);
nor U36915 (N_36915,N_36485,N_36309);
nor U36916 (N_36916,N_36007,N_36340);
xor U36917 (N_36917,N_36039,N_36419);
and U36918 (N_36918,N_36065,N_36076);
and U36919 (N_36919,N_36403,N_36490);
or U36920 (N_36920,N_36351,N_36245);
nor U36921 (N_36921,N_36238,N_36362);
nand U36922 (N_36922,N_36033,N_36013);
or U36923 (N_36923,N_36097,N_36240);
nand U36924 (N_36924,N_36106,N_36332);
nor U36925 (N_36925,N_36404,N_36124);
and U36926 (N_36926,N_36116,N_36047);
nor U36927 (N_36927,N_36068,N_36285);
nand U36928 (N_36928,N_36180,N_36356);
xor U36929 (N_36929,N_36132,N_36450);
and U36930 (N_36930,N_36019,N_36495);
and U36931 (N_36931,N_36204,N_36288);
and U36932 (N_36932,N_36002,N_36097);
nor U36933 (N_36933,N_36271,N_36266);
xnor U36934 (N_36934,N_36350,N_36298);
nand U36935 (N_36935,N_36386,N_36349);
nor U36936 (N_36936,N_36473,N_36003);
xnor U36937 (N_36937,N_36439,N_36056);
and U36938 (N_36938,N_36386,N_36234);
and U36939 (N_36939,N_36202,N_36220);
and U36940 (N_36940,N_36487,N_36334);
or U36941 (N_36941,N_36112,N_36029);
or U36942 (N_36942,N_36147,N_36158);
or U36943 (N_36943,N_36377,N_36203);
nand U36944 (N_36944,N_36090,N_36061);
nand U36945 (N_36945,N_36272,N_36277);
nand U36946 (N_36946,N_36311,N_36440);
and U36947 (N_36947,N_36197,N_36073);
nand U36948 (N_36948,N_36459,N_36412);
nor U36949 (N_36949,N_36258,N_36253);
and U36950 (N_36950,N_36096,N_36415);
nand U36951 (N_36951,N_36041,N_36353);
and U36952 (N_36952,N_36014,N_36237);
and U36953 (N_36953,N_36493,N_36065);
xor U36954 (N_36954,N_36147,N_36086);
nor U36955 (N_36955,N_36498,N_36376);
and U36956 (N_36956,N_36000,N_36101);
or U36957 (N_36957,N_36274,N_36105);
nand U36958 (N_36958,N_36448,N_36305);
or U36959 (N_36959,N_36270,N_36228);
or U36960 (N_36960,N_36167,N_36165);
nor U36961 (N_36961,N_36290,N_36203);
nor U36962 (N_36962,N_36404,N_36057);
nand U36963 (N_36963,N_36143,N_36275);
and U36964 (N_36964,N_36330,N_36398);
and U36965 (N_36965,N_36216,N_36290);
nor U36966 (N_36966,N_36260,N_36251);
and U36967 (N_36967,N_36187,N_36017);
nand U36968 (N_36968,N_36095,N_36103);
and U36969 (N_36969,N_36134,N_36315);
nand U36970 (N_36970,N_36039,N_36031);
nand U36971 (N_36971,N_36224,N_36045);
nand U36972 (N_36972,N_36304,N_36480);
and U36973 (N_36973,N_36324,N_36255);
or U36974 (N_36974,N_36027,N_36010);
nor U36975 (N_36975,N_36466,N_36075);
and U36976 (N_36976,N_36141,N_36112);
or U36977 (N_36977,N_36227,N_36360);
nand U36978 (N_36978,N_36362,N_36287);
or U36979 (N_36979,N_36178,N_36243);
xnor U36980 (N_36980,N_36354,N_36302);
nand U36981 (N_36981,N_36342,N_36192);
nor U36982 (N_36982,N_36443,N_36312);
nor U36983 (N_36983,N_36177,N_36260);
nand U36984 (N_36984,N_36246,N_36127);
or U36985 (N_36985,N_36381,N_36127);
or U36986 (N_36986,N_36158,N_36406);
or U36987 (N_36987,N_36114,N_36415);
and U36988 (N_36988,N_36155,N_36383);
or U36989 (N_36989,N_36495,N_36391);
or U36990 (N_36990,N_36308,N_36320);
or U36991 (N_36991,N_36122,N_36399);
and U36992 (N_36992,N_36372,N_36086);
nand U36993 (N_36993,N_36090,N_36446);
xnor U36994 (N_36994,N_36389,N_36094);
nor U36995 (N_36995,N_36346,N_36223);
and U36996 (N_36996,N_36438,N_36154);
nor U36997 (N_36997,N_36001,N_36075);
or U36998 (N_36998,N_36145,N_36308);
and U36999 (N_36999,N_36379,N_36017);
or U37000 (N_37000,N_36741,N_36564);
nor U37001 (N_37001,N_36713,N_36732);
and U37002 (N_37002,N_36971,N_36687);
xor U37003 (N_37003,N_36511,N_36724);
nand U37004 (N_37004,N_36685,N_36800);
nand U37005 (N_37005,N_36743,N_36575);
xor U37006 (N_37006,N_36683,N_36990);
and U37007 (N_37007,N_36705,N_36832);
nand U37008 (N_37008,N_36817,N_36695);
xor U37009 (N_37009,N_36974,N_36653);
nand U37010 (N_37010,N_36907,N_36877);
nand U37011 (N_37011,N_36969,N_36898);
and U37012 (N_37012,N_36917,N_36759);
and U37013 (N_37013,N_36966,N_36748);
xor U37014 (N_37014,N_36649,N_36532);
and U37015 (N_37015,N_36622,N_36987);
and U37016 (N_37016,N_36651,N_36775);
nor U37017 (N_37017,N_36854,N_36998);
or U37018 (N_37018,N_36804,N_36659);
or U37019 (N_37019,N_36814,N_36562);
and U37020 (N_37020,N_36860,N_36984);
nand U37021 (N_37021,N_36618,N_36568);
or U37022 (N_37022,N_36662,N_36897);
xnor U37023 (N_37023,N_36903,N_36566);
and U37024 (N_37024,N_36892,N_36760);
and U37025 (N_37025,N_36671,N_36818);
nand U37026 (N_37026,N_36738,N_36955);
or U37027 (N_37027,N_36584,N_36587);
nand U37028 (N_37028,N_36936,N_36747);
nand U37029 (N_37029,N_36650,N_36600);
nor U37030 (N_37030,N_36961,N_36951);
nor U37031 (N_37031,N_36585,N_36824);
nor U37032 (N_37032,N_36553,N_36534);
nor U37033 (N_37033,N_36710,N_36613);
and U37034 (N_37034,N_36932,N_36661);
or U37035 (N_37035,N_36709,N_36792);
nand U37036 (N_37036,N_36597,N_36993);
nor U37037 (N_37037,N_36595,N_36776);
nand U37038 (N_37038,N_36522,N_36931);
or U37039 (N_37039,N_36642,N_36889);
nand U37040 (N_37040,N_36561,N_36972);
and U37041 (N_37041,N_36894,N_36546);
and U37042 (N_37042,N_36576,N_36670);
nand U37043 (N_37043,N_36949,N_36608);
and U37044 (N_37044,N_36664,N_36714);
nand U37045 (N_37045,N_36537,N_36803);
xnor U37046 (N_37046,N_36719,N_36797);
nor U37047 (N_37047,N_36866,N_36787);
nand U37048 (N_37048,N_36698,N_36864);
and U37049 (N_37049,N_36855,N_36862);
xnor U37050 (N_37050,N_36846,N_36810);
or U37051 (N_37051,N_36588,N_36943);
nand U37052 (N_37052,N_36711,N_36723);
nand U37053 (N_37053,N_36682,N_36833);
or U37054 (N_37054,N_36909,N_36733);
nor U37055 (N_37055,N_36875,N_36934);
and U37056 (N_37056,N_36629,N_36594);
or U37057 (N_37057,N_36782,N_36563);
or U37058 (N_37058,N_36997,N_36857);
nand U37059 (N_37059,N_36908,N_36541);
nor U37060 (N_37060,N_36874,N_36539);
nor U37061 (N_37061,N_36633,N_36829);
xnor U37062 (N_37062,N_36995,N_36948);
nor U37063 (N_37063,N_36550,N_36796);
and U37064 (N_37064,N_36774,N_36603);
xor U37065 (N_37065,N_36837,N_36675);
nand U37066 (N_37066,N_36820,N_36580);
nor U37067 (N_37067,N_36996,N_36935);
and U37068 (N_37068,N_36836,N_36918);
and U37069 (N_37069,N_36913,N_36569);
or U37070 (N_37070,N_36611,N_36668);
nor U37071 (N_37071,N_36788,N_36933);
or U37072 (N_37072,N_36765,N_36612);
nor U37073 (N_37073,N_36910,N_36731);
or U37074 (N_37074,N_36989,N_36921);
nor U37075 (N_37075,N_36519,N_36601);
and U37076 (N_37076,N_36880,N_36663);
nand U37077 (N_37077,N_36544,N_36925);
nor U37078 (N_37078,N_36763,N_36531);
and U37079 (N_37079,N_36841,N_36556);
xor U37080 (N_37080,N_36527,N_36644);
nor U37081 (N_37081,N_36795,N_36500);
nand U37082 (N_37082,N_36703,N_36545);
xnor U37083 (N_37083,N_36916,N_36609);
xnor U37084 (N_37084,N_36736,N_36808);
nand U37085 (N_37085,N_36838,N_36999);
xnor U37086 (N_37086,N_36507,N_36845);
or U37087 (N_37087,N_36548,N_36956);
nand U37088 (N_37088,N_36677,N_36596);
and U37089 (N_37089,N_36952,N_36586);
xnor U37090 (N_37090,N_36706,N_36915);
or U37091 (N_37091,N_36988,N_36669);
nand U37092 (N_37092,N_36912,N_36926);
xor U37093 (N_37093,N_36885,N_36791);
nand U37094 (N_37094,N_36528,N_36821);
nand U37095 (N_37095,N_36872,N_36930);
nand U37096 (N_37096,N_36764,N_36652);
nor U37097 (N_37097,N_36666,N_36807);
or U37098 (N_37098,N_36890,N_36637);
nor U37099 (N_37099,N_36606,N_36794);
or U37100 (N_37100,N_36784,N_36513);
or U37101 (N_37101,N_36887,N_36624);
or U37102 (N_37102,N_36630,N_36578);
or U37103 (N_37103,N_36766,N_36826);
nand U37104 (N_37104,N_36542,N_36945);
nor U37105 (N_37105,N_36802,N_36986);
nand U37106 (N_37106,N_36660,N_36806);
and U37107 (N_37107,N_36757,N_36602);
or U37108 (N_37108,N_36726,N_36905);
and U37109 (N_37109,N_36684,N_36750);
xor U37110 (N_37110,N_36508,N_36924);
and U37111 (N_37111,N_36657,N_36967);
or U37112 (N_37112,N_36737,N_36769);
nor U37113 (N_37113,N_36786,N_36780);
nor U37114 (N_37114,N_36538,N_36883);
and U37115 (N_37115,N_36623,N_36673);
nand U37116 (N_37116,N_36589,N_36886);
nand U37117 (N_37117,N_36746,N_36979);
nand U37118 (N_37118,N_36565,N_36842);
and U37119 (N_37119,N_36767,N_36783);
nand U37120 (N_37120,N_36557,N_36621);
nor U37121 (N_37121,N_36728,N_36648);
xor U37122 (N_37122,N_36672,N_36515);
and U37123 (N_37123,N_36983,N_36771);
and U37124 (N_37124,N_36516,N_36535);
nand U37125 (N_37125,N_36923,N_36893);
or U37126 (N_37126,N_36811,N_36559);
and U37127 (N_37127,N_36902,N_36975);
nand U37128 (N_37128,N_36610,N_36526);
and U37129 (N_37129,N_36571,N_36579);
or U37130 (N_37130,N_36701,N_36744);
nor U37131 (N_37131,N_36994,N_36730);
and U37132 (N_37132,N_36740,N_36963);
and U37133 (N_37133,N_36859,N_36968);
or U37134 (N_37134,N_36843,N_36679);
nor U37135 (N_37135,N_36506,N_36828);
or U37136 (N_37136,N_36977,N_36614);
or U37137 (N_37137,N_36944,N_36911);
xnor U37138 (N_37138,N_36693,N_36754);
nand U37139 (N_37139,N_36965,N_36779);
and U37140 (N_37140,N_36697,N_36840);
or U37141 (N_37141,N_36947,N_36639);
and U37142 (N_37142,N_36888,N_36715);
nor U37143 (N_37143,N_36985,N_36593);
nand U37144 (N_37144,N_36941,N_36950);
nor U37145 (N_37145,N_36552,N_36980);
nor U37146 (N_37146,N_36708,N_36895);
nand U37147 (N_37147,N_36667,N_36848);
and U37148 (N_37148,N_36899,N_36962);
nor U37149 (N_37149,N_36574,N_36785);
xor U37150 (N_37150,N_36772,N_36896);
nand U37151 (N_37151,N_36768,N_36938);
nor U37152 (N_37152,N_36521,N_36745);
or U37153 (N_37153,N_36958,N_36599);
or U37154 (N_37154,N_36819,N_36647);
nand U37155 (N_37155,N_36646,N_36725);
or U37156 (N_37156,N_36640,N_36635);
nor U37157 (N_37157,N_36879,N_36619);
xnor U37158 (N_37158,N_36835,N_36702);
or U37159 (N_37159,N_36581,N_36834);
and U37160 (N_37160,N_36954,N_36805);
nor U37161 (N_37161,N_36505,N_36827);
and U37162 (N_37162,N_36973,N_36781);
or U37163 (N_37163,N_36816,N_36825);
and U37164 (N_37164,N_36856,N_36823);
nand U37165 (N_37165,N_36699,N_36970);
nor U37166 (N_37166,N_36616,N_36929);
and U37167 (N_37167,N_36605,N_36525);
xor U37168 (N_37168,N_36940,N_36676);
nand U37169 (N_37169,N_36632,N_36844);
and U37170 (N_37170,N_36543,N_36577);
nand U37171 (N_37171,N_36517,N_36761);
and U37172 (N_37172,N_36549,N_36716);
nor U37173 (N_37173,N_36991,N_36873);
nand U37174 (N_37174,N_36801,N_36690);
or U37175 (N_37175,N_36555,N_36688);
and U37176 (N_37176,N_36536,N_36900);
and U37177 (N_37177,N_36793,N_36582);
nand U37178 (N_37178,N_36604,N_36798);
nor U37179 (N_37179,N_36689,N_36529);
and U37180 (N_37180,N_36729,N_36778);
nor U37181 (N_37181,N_36554,N_36937);
xor U37182 (N_37182,N_36533,N_36830);
or U37183 (N_37183,N_36878,N_36674);
and U37184 (N_37184,N_36501,N_36572);
or U37185 (N_37185,N_36510,N_36583);
and U37186 (N_37186,N_36520,N_36678);
and U37187 (N_37187,N_36720,N_36755);
nor U37188 (N_37188,N_36964,N_36919);
or U37189 (N_37189,N_36904,N_36869);
nand U37190 (N_37190,N_36598,N_36863);
and U37191 (N_37191,N_36634,N_36686);
xor U37192 (N_37192,N_36502,N_36680);
or U37193 (N_37193,N_36927,N_36751);
nand U37194 (N_37194,N_36812,N_36858);
nor U37195 (N_37195,N_36920,N_36981);
or U37196 (N_37196,N_36882,N_36628);
or U37197 (N_37197,N_36512,N_36960);
or U37198 (N_37198,N_36839,N_36617);
and U37199 (N_37199,N_36762,N_36742);
nor U37200 (N_37200,N_36691,N_36645);
or U37201 (N_37201,N_36749,N_36727);
and U37202 (N_37202,N_36692,N_36939);
nor U37203 (N_37203,N_36734,N_36551);
nor U37204 (N_37204,N_36503,N_36957);
nand U37205 (N_37205,N_36570,N_36643);
nand U37206 (N_37206,N_36607,N_36567);
or U37207 (N_37207,N_36540,N_36770);
nor U37208 (N_37208,N_36753,N_36959);
or U37209 (N_37209,N_36922,N_36704);
and U37210 (N_37210,N_36906,N_36871);
or U37211 (N_37211,N_36658,N_36853);
nor U37212 (N_37212,N_36636,N_36815);
and U37213 (N_37213,N_36809,N_36694);
or U37214 (N_37214,N_36847,N_36928);
and U37215 (N_37215,N_36756,N_36504);
and U37216 (N_37216,N_36573,N_36831);
nand U37217 (N_37217,N_36790,N_36758);
nor U37218 (N_37218,N_36631,N_36591);
or U37219 (N_37219,N_36615,N_36558);
nand U37220 (N_37220,N_36681,N_36982);
nor U37221 (N_37221,N_36696,N_36739);
nor U37222 (N_37222,N_36722,N_36777);
or U37223 (N_37223,N_36861,N_36865);
xor U37224 (N_37224,N_36656,N_36665);
xnor U37225 (N_37225,N_36946,N_36813);
nor U37226 (N_37226,N_36707,N_36735);
or U37227 (N_37227,N_36914,N_36752);
nand U37228 (N_37228,N_36530,N_36626);
or U37229 (N_37229,N_36891,N_36868);
and U37230 (N_37230,N_36822,N_36547);
and U37231 (N_37231,N_36942,N_36884);
and U37232 (N_37232,N_36592,N_36976);
nand U37233 (N_37233,N_36712,N_36718);
nor U37234 (N_37234,N_36620,N_36849);
nand U37235 (N_37235,N_36992,N_36509);
nand U37236 (N_37236,N_36627,N_36717);
or U37237 (N_37237,N_36876,N_36978);
or U37238 (N_37238,N_36773,N_36789);
nor U37239 (N_37239,N_36590,N_36625);
nor U37240 (N_37240,N_36654,N_36523);
nand U37241 (N_37241,N_36655,N_36852);
nor U37242 (N_37242,N_36721,N_36870);
nand U37243 (N_37243,N_36518,N_36851);
nand U37244 (N_37244,N_36524,N_36514);
nand U37245 (N_37245,N_36638,N_36799);
or U37246 (N_37246,N_36881,N_36560);
and U37247 (N_37247,N_36641,N_36700);
or U37248 (N_37248,N_36850,N_36901);
or U37249 (N_37249,N_36953,N_36867);
or U37250 (N_37250,N_36590,N_36618);
nand U37251 (N_37251,N_36669,N_36512);
xor U37252 (N_37252,N_36692,N_36834);
or U37253 (N_37253,N_36640,N_36774);
xnor U37254 (N_37254,N_36953,N_36776);
and U37255 (N_37255,N_36838,N_36873);
or U37256 (N_37256,N_36821,N_36786);
nor U37257 (N_37257,N_36538,N_36953);
or U37258 (N_37258,N_36932,N_36575);
nand U37259 (N_37259,N_36704,N_36880);
and U37260 (N_37260,N_36936,N_36824);
and U37261 (N_37261,N_36513,N_36665);
or U37262 (N_37262,N_36907,N_36992);
and U37263 (N_37263,N_36845,N_36879);
nand U37264 (N_37264,N_36553,N_36533);
nor U37265 (N_37265,N_36762,N_36638);
nor U37266 (N_37266,N_36600,N_36839);
nand U37267 (N_37267,N_36517,N_36853);
nand U37268 (N_37268,N_36635,N_36942);
nor U37269 (N_37269,N_36690,N_36607);
and U37270 (N_37270,N_36731,N_36839);
xnor U37271 (N_37271,N_36749,N_36942);
nand U37272 (N_37272,N_36569,N_36955);
nand U37273 (N_37273,N_36857,N_36780);
xnor U37274 (N_37274,N_36700,N_36537);
nor U37275 (N_37275,N_36605,N_36812);
or U37276 (N_37276,N_36539,N_36562);
nor U37277 (N_37277,N_36905,N_36559);
or U37278 (N_37278,N_36630,N_36924);
nand U37279 (N_37279,N_36928,N_36543);
or U37280 (N_37280,N_36512,N_36862);
or U37281 (N_37281,N_36796,N_36710);
nor U37282 (N_37282,N_36634,N_36663);
or U37283 (N_37283,N_36657,N_36554);
or U37284 (N_37284,N_36694,N_36551);
nor U37285 (N_37285,N_36932,N_36765);
or U37286 (N_37286,N_36595,N_36974);
or U37287 (N_37287,N_36504,N_36589);
nand U37288 (N_37288,N_36773,N_36921);
and U37289 (N_37289,N_36518,N_36794);
nand U37290 (N_37290,N_36941,N_36574);
and U37291 (N_37291,N_36739,N_36611);
nor U37292 (N_37292,N_36520,N_36971);
or U37293 (N_37293,N_36891,N_36602);
nor U37294 (N_37294,N_36792,N_36968);
and U37295 (N_37295,N_36634,N_36564);
xor U37296 (N_37296,N_36775,N_36840);
nand U37297 (N_37297,N_36828,N_36936);
or U37298 (N_37298,N_36912,N_36637);
nand U37299 (N_37299,N_36717,N_36571);
or U37300 (N_37300,N_36672,N_36957);
and U37301 (N_37301,N_36743,N_36559);
nand U37302 (N_37302,N_36696,N_36989);
or U37303 (N_37303,N_36739,N_36947);
nor U37304 (N_37304,N_36951,N_36610);
nand U37305 (N_37305,N_36573,N_36528);
or U37306 (N_37306,N_36848,N_36766);
nand U37307 (N_37307,N_36754,N_36898);
nand U37308 (N_37308,N_36508,N_36916);
nor U37309 (N_37309,N_36566,N_36603);
nor U37310 (N_37310,N_36800,N_36736);
or U37311 (N_37311,N_36621,N_36726);
and U37312 (N_37312,N_36707,N_36573);
nand U37313 (N_37313,N_36897,N_36559);
and U37314 (N_37314,N_36797,N_36679);
nor U37315 (N_37315,N_36708,N_36781);
nor U37316 (N_37316,N_36796,N_36834);
nand U37317 (N_37317,N_36560,N_36755);
nor U37318 (N_37318,N_36955,N_36728);
nor U37319 (N_37319,N_36885,N_36952);
nor U37320 (N_37320,N_36922,N_36548);
and U37321 (N_37321,N_36744,N_36646);
nor U37322 (N_37322,N_36566,N_36910);
nor U37323 (N_37323,N_36566,N_36757);
or U37324 (N_37324,N_36830,N_36777);
or U37325 (N_37325,N_36945,N_36776);
nor U37326 (N_37326,N_36947,N_36541);
xor U37327 (N_37327,N_36939,N_36863);
nor U37328 (N_37328,N_36514,N_36660);
or U37329 (N_37329,N_36996,N_36617);
nor U37330 (N_37330,N_36554,N_36764);
or U37331 (N_37331,N_36740,N_36749);
nand U37332 (N_37332,N_36953,N_36626);
nand U37333 (N_37333,N_36545,N_36939);
and U37334 (N_37334,N_36872,N_36746);
or U37335 (N_37335,N_36676,N_36672);
and U37336 (N_37336,N_36671,N_36911);
or U37337 (N_37337,N_36502,N_36859);
nor U37338 (N_37338,N_36700,N_36855);
nand U37339 (N_37339,N_36863,N_36693);
xor U37340 (N_37340,N_36735,N_36503);
nand U37341 (N_37341,N_36803,N_36681);
or U37342 (N_37342,N_36847,N_36783);
xor U37343 (N_37343,N_36917,N_36774);
and U37344 (N_37344,N_36848,N_36864);
nor U37345 (N_37345,N_36801,N_36652);
or U37346 (N_37346,N_36889,N_36918);
nor U37347 (N_37347,N_36987,N_36606);
nand U37348 (N_37348,N_36700,N_36750);
or U37349 (N_37349,N_36876,N_36582);
nor U37350 (N_37350,N_36867,N_36891);
or U37351 (N_37351,N_36990,N_36563);
or U37352 (N_37352,N_36877,N_36978);
nand U37353 (N_37353,N_36678,N_36620);
or U37354 (N_37354,N_36954,N_36705);
xnor U37355 (N_37355,N_36878,N_36555);
or U37356 (N_37356,N_36944,N_36839);
nor U37357 (N_37357,N_36673,N_36564);
or U37358 (N_37358,N_36960,N_36778);
nand U37359 (N_37359,N_36863,N_36787);
nor U37360 (N_37360,N_36511,N_36850);
and U37361 (N_37361,N_36754,N_36839);
and U37362 (N_37362,N_36698,N_36546);
or U37363 (N_37363,N_36770,N_36788);
and U37364 (N_37364,N_36829,N_36994);
and U37365 (N_37365,N_36949,N_36819);
nand U37366 (N_37366,N_36779,N_36702);
nor U37367 (N_37367,N_36815,N_36659);
and U37368 (N_37368,N_36975,N_36712);
nor U37369 (N_37369,N_36850,N_36763);
and U37370 (N_37370,N_36864,N_36557);
nor U37371 (N_37371,N_36794,N_36779);
and U37372 (N_37372,N_36584,N_36885);
xor U37373 (N_37373,N_36575,N_36521);
or U37374 (N_37374,N_36513,N_36957);
nand U37375 (N_37375,N_36831,N_36782);
or U37376 (N_37376,N_36945,N_36835);
or U37377 (N_37377,N_36602,N_36796);
nor U37378 (N_37378,N_36910,N_36684);
and U37379 (N_37379,N_36831,N_36899);
and U37380 (N_37380,N_36594,N_36633);
and U37381 (N_37381,N_36776,N_36635);
nor U37382 (N_37382,N_36988,N_36689);
nor U37383 (N_37383,N_36931,N_36915);
nor U37384 (N_37384,N_36518,N_36829);
nor U37385 (N_37385,N_36784,N_36708);
or U37386 (N_37386,N_36765,N_36954);
nor U37387 (N_37387,N_36825,N_36833);
or U37388 (N_37388,N_36977,N_36759);
nor U37389 (N_37389,N_36789,N_36976);
nand U37390 (N_37390,N_36503,N_36669);
and U37391 (N_37391,N_36917,N_36964);
or U37392 (N_37392,N_36864,N_36699);
nor U37393 (N_37393,N_36854,N_36907);
or U37394 (N_37394,N_36532,N_36766);
or U37395 (N_37395,N_36862,N_36732);
nand U37396 (N_37396,N_36526,N_36621);
and U37397 (N_37397,N_36910,N_36517);
or U37398 (N_37398,N_36638,N_36656);
and U37399 (N_37399,N_36928,N_36923);
and U37400 (N_37400,N_36517,N_36746);
and U37401 (N_37401,N_36602,N_36779);
and U37402 (N_37402,N_36523,N_36888);
and U37403 (N_37403,N_36646,N_36522);
or U37404 (N_37404,N_36988,N_36975);
or U37405 (N_37405,N_36574,N_36871);
nand U37406 (N_37406,N_36810,N_36874);
and U37407 (N_37407,N_36539,N_36689);
and U37408 (N_37408,N_36542,N_36730);
xnor U37409 (N_37409,N_36617,N_36896);
nand U37410 (N_37410,N_36964,N_36775);
nand U37411 (N_37411,N_36535,N_36765);
nor U37412 (N_37412,N_36555,N_36788);
and U37413 (N_37413,N_36927,N_36506);
nor U37414 (N_37414,N_36723,N_36945);
nand U37415 (N_37415,N_36512,N_36526);
and U37416 (N_37416,N_36527,N_36997);
and U37417 (N_37417,N_36975,N_36721);
nor U37418 (N_37418,N_36601,N_36983);
xnor U37419 (N_37419,N_36676,N_36818);
or U37420 (N_37420,N_36879,N_36687);
and U37421 (N_37421,N_36648,N_36993);
or U37422 (N_37422,N_36858,N_36534);
nor U37423 (N_37423,N_36935,N_36870);
and U37424 (N_37424,N_36822,N_36952);
nand U37425 (N_37425,N_36907,N_36772);
and U37426 (N_37426,N_36554,N_36880);
and U37427 (N_37427,N_36639,N_36885);
nand U37428 (N_37428,N_36748,N_36803);
nor U37429 (N_37429,N_36825,N_36821);
nand U37430 (N_37430,N_36699,N_36870);
and U37431 (N_37431,N_36832,N_36720);
nand U37432 (N_37432,N_36806,N_36693);
and U37433 (N_37433,N_36602,N_36848);
or U37434 (N_37434,N_36751,N_36613);
nand U37435 (N_37435,N_36674,N_36876);
and U37436 (N_37436,N_36961,N_36892);
nor U37437 (N_37437,N_36705,N_36658);
nand U37438 (N_37438,N_36629,N_36656);
nor U37439 (N_37439,N_36671,N_36904);
and U37440 (N_37440,N_36840,N_36784);
or U37441 (N_37441,N_36982,N_36698);
nand U37442 (N_37442,N_36542,N_36535);
and U37443 (N_37443,N_36677,N_36517);
xor U37444 (N_37444,N_36638,N_36579);
xor U37445 (N_37445,N_36847,N_36648);
nand U37446 (N_37446,N_36639,N_36907);
nor U37447 (N_37447,N_36813,N_36509);
and U37448 (N_37448,N_36911,N_36718);
nand U37449 (N_37449,N_36574,N_36680);
and U37450 (N_37450,N_36656,N_36735);
xor U37451 (N_37451,N_36507,N_36613);
and U37452 (N_37452,N_36559,N_36695);
nor U37453 (N_37453,N_36769,N_36859);
nand U37454 (N_37454,N_36634,N_36506);
xor U37455 (N_37455,N_36752,N_36712);
nor U37456 (N_37456,N_36978,N_36962);
or U37457 (N_37457,N_36588,N_36602);
xor U37458 (N_37458,N_36630,N_36881);
and U37459 (N_37459,N_36885,N_36611);
or U37460 (N_37460,N_36545,N_36601);
and U37461 (N_37461,N_36833,N_36989);
xnor U37462 (N_37462,N_36725,N_36829);
nand U37463 (N_37463,N_36880,N_36652);
and U37464 (N_37464,N_36578,N_36795);
xnor U37465 (N_37465,N_36957,N_36819);
xnor U37466 (N_37466,N_36880,N_36545);
nor U37467 (N_37467,N_36821,N_36871);
nor U37468 (N_37468,N_36859,N_36854);
and U37469 (N_37469,N_36707,N_36774);
nand U37470 (N_37470,N_36919,N_36906);
and U37471 (N_37471,N_36909,N_36843);
nand U37472 (N_37472,N_36722,N_36925);
nand U37473 (N_37473,N_36854,N_36601);
nor U37474 (N_37474,N_36622,N_36628);
and U37475 (N_37475,N_36939,N_36841);
and U37476 (N_37476,N_36915,N_36636);
nor U37477 (N_37477,N_36639,N_36831);
and U37478 (N_37478,N_36908,N_36603);
nor U37479 (N_37479,N_36650,N_36967);
and U37480 (N_37480,N_36651,N_36819);
nand U37481 (N_37481,N_36589,N_36675);
or U37482 (N_37482,N_36828,N_36658);
nor U37483 (N_37483,N_36598,N_36643);
and U37484 (N_37484,N_36840,N_36685);
or U37485 (N_37485,N_36562,N_36747);
and U37486 (N_37486,N_36754,N_36807);
nor U37487 (N_37487,N_36922,N_36709);
and U37488 (N_37488,N_36785,N_36595);
xnor U37489 (N_37489,N_36740,N_36572);
and U37490 (N_37490,N_36527,N_36906);
or U37491 (N_37491,N_36840,N_36734);
nand U37492 (N_37492,N_36607,N_36500);
or U37493 (N_37493,N_36996,N_36872);
or U37494 (N_37494,N_36794,N_36817);
nand U37495 (N_37495,N_36942,N_36680);
and U37496 (N_37496,N_36572,N_36515);
and U37497 (N_37497,N_36761,N_36608);
nand U37498 (N_37498,N_36989,N_36949);
nand U37499 (N_37499,N_36847,N_36673);
nor U37500 (N_37500,N_37075,N_37379);
or U37501 (N_37501,N_37090,N_37372);
or U37502 (N_37502,N_37324,N_37469);
nor U37503 (N_37503,N_37449,N_37097);
and U37504 (N_37504,N_37129,N_37254);
or U37505 (N_37505,N_37438,N_37119);
and U37506 (N_37506,N_37441,N_37237);
or U37507 (N_37507,N_37258,N_37122);
xnor U37508 (N_37508,N_37384,N_37305);
nand U37509 (N_37509,N_37420,N_37195);
nand U37510 (N_37510,N_37034,N_37040);
and U37511 (N_37511,N_37033,N_37247);
and U37512 (N_37512,N_37087,N_37472);
and U37513 (N_37513,N_37493,N_37068);
nor U37514 (N_37514,N_37021,N_37459);
nand U37515 (N_37515,N_37363,N_37158);
and U37516 (N_37516,N_37104,N_37130);
nor U37517 (N_37517,N_37489,N_37440);
nor U37518 (N_37518,N_37264,N_37125);
nor U37519 (N_37519,N_37446,N_37020);
nand U37520 (N_37520,N_37396,N_37289);
or U37521 (N_37521,N_37200,N_37037);
and U37522 (N_37522,N_37394,N_37418);
nand U37523 (N_37523,N_37393,N_37266);
and U37524 (N_37524,N_37273,N_37380);
and U37525 (N_37525,N_37412,N_37454);
nor U37526 (N_37526,N_37225,N_37271);
nor U37527 (N_37527,N_37285,N_37259);
or U37528 (N_37528,N_37265,N_37452);
nand U37529 (N_37529,N_37278,N_37096);
or U37530 (N_37530,N_37220,N_37343);
nand U37531 (N_37531,N_37052,N_37132);
nor U37532 (N_37532,N_37407,N_37221);
or U37533 (N_37533,N_37240,N_37084);
nor U37534 (N_37534,N_37042,N_37198);
xor U37535 (N_37535,N_37082,N_37382);
xor U37536 (N_37536,N_37408,N_37288);
nor U37537 (N_37537,N_37373,N_37491);
or U37538 (N_37538,N_37235,N_37092);
or U37539 (N_37539,N_37284,N_37071);
and U37540 (N_37540,N_37135,N_37444);
or U37541 (N_37541,N_37045,N_37048);
xnor U37542 (N_37542,N_37074,N_37333);
nor U37543 (N_37543,N_37361,N_37012);
xnor U37544 (N_37544,N_37003,N_37005);
or U37545 (N_37545,N_37138,N_37080);
nor U37546 (N_37546,N_37476,N_37173);
nor U37547 (N_37547,N_37405,N_37117);
nand U37548 (N_37548,N_37088,N_37283);
nand U37549 (N_37549,N_37267,N_37229);
nand U37550 (N_37550,N_37498,N_37432);
and U37551 (N_37551,N_37103,N_37035);
or U37552 (N_37552,N_37159,N_37185);
nand U37553 (N_37553,N_37487,N_37114);
and U37554 (N_37554,N_37126,N_37248);
or U37555 (N_37555,N_37176,N_37057);
or U37556 (N_37556,N_37344,N_37197);
nand U37557 (N_37557,N_37133,N_37011);
and U37558 (N_37558,N_37029,N_37314);
or U37559 (N_37559,N_37317,N_37112);
and U37560 (N_37560,N_37059,N_37019);
xnor U37561 (N_37561,N_37147,N_37014);
nor U37562 (N_37562,N_37190,N_37111);
and U37563 (N_37563,N_37322,N_37142);
and U37564 (N_37564,N_37089,N_37083);
xnor U37565 (N_37565,N_37300,N_37479);
nand U37566 (N_37566,N_37272,N_37047);
nand U37567 (N_37567,N_37329,N_37004);
or U37568 (N_37568,N_37417,N_37468);
and U37569 (N_37569,N_37152,N_37341);
and U37570 (N_37570,N_37465,N_37389);
nand U37571 (N_37571,N_37091,N_37348);
nand U37572 (N_37572,N_37471,N_37213);
nand U37573 (N_37573,N_37072,N_37025);
and U37574 (N_37574,N_37447,N_37257);
or U37575 (N_37575,N_37340,N_37419);
or U37576 (N_37576,N_37427,N_37275);
xnor U37577 (N_37577,N_37162,N_37167);
xor U37578 (N_37578,N_37354,N_37141);
nand U37579 (N_37579,N_37450,N_37243);
nor U37580 (N_37580,N_37378,N_37064);
or U37581 (N_37581,N_37430,N_37001);
and U37582 (N_37582,N_37186,N_37388);
or U37583 (N_37583,N_37073,N_37172);
nand U37584 (N_37584,N_37295,N_37118);
xor U37585 (N_37585,N_37274,N_37208);
or U37586 (N_37586,N_37255,N_37262);
or U37587 (N_37587,N_37281,N_37397);
nand U37588 (N_37588,N_37050,N_37453);
and U37589 (N_37589,N_37303,N_37320);
nand U37590 (N_37590,N_37007,N_37425);
and U37591 (N_37591,N_37106,N_37279);
and U37592 (N_37592,N_37239,N_37386);
or U37593 (N_37593,N_37157,N_37124);
nand U37594 (N_37594,N_37325,N_37110);
and U37595 (N_37595,N_37194,N_37480);
or U37596 (N_37596,N_37401,N_37352);
nand U37597 (N_37597,N_37013,N_37413);
nand U37598 (N_37598,N_37306,N_37346);
nor U37599 (N_37599,N_37426,N_37457);
or U37600 (N_37600,N_37137,N_37353);
nor U37601 (N_37601,N_37339,N_37252);
and U37602 (N_37602,N_37335,N_37085);
or U37603 (N_37603,N_37381,N_37038);
xnor U37604 (N_37604,N_37277,N_37250);
and U37605 (N_37605,N_37219,N_37403);
and U37606 (N_37606,N_37392,N_37364);
nor U37607 (N_37607,N_37230,N_37188);
and U37608 (N_37608,N_37307,N_37140);
and U37609 (N_37609,N_37251,N_37431);
or U37610 (N_37610,N_37349,N_37345);
nand U37611 (N_37611,N_37054,N_37107);
and U37612 (N_37612,N_37144,N_37365);
nand U37613 (N_37613,N_37460,N_37475);
nand U37614 (N_37614,N_37357,N_37256);
xnor U37615 (N_37615,N_37253,N_37336);
nand U37616 (N_37616,N_37398,N_37016);
xnor U37617 (N_37617,N_37227,N_37318);
xor U37618 (N_37618,N_37411,N_37293);
or U37619 (N_37619,N_37051,N_37448);
nor U37620 (N_37620,N_37436,N_37136);
nand U37621 (N_37621,N_37299,N_37234);
nand U37622 (N_37622,N_37070,N_37242);
xor U37623 (N_37623,N_37120,N_37205);
xnor U37624 (N_37624,N_37095,N_37212);
or U37625 (N_37625,N_37467,N_37215);
nor U37626 (N_37626,N_37296,N_37406);
and U37627 (N_37627,N_37287,N_37433);
or U37628 (N_37628,N_37105,N_37323);
and U37629 (N_37629,N_37169,N_37017);
nand U37630 (N_37630,N_37202,N_37312);
and U37631 (N_37631,N_37218,N_37171);
nor U37632 (N_37632,N_37199,N_37423);
nand U37633 (N_37633,N_37470,N_37164);
nor U37634 (N_37634,N_37370,N_37055);
nor U37635 (N_37635,N_37216,N_37161);
nor U37636 (N_37636,N_37187,N_37477);
nor U37637 (N_37637,N_37223,N_37244);
and U37638 (N_37638,N_37414,N_37139);
nor U37639 (N_37639,N_37214,N_37154);
nand U37640 (N_37640,N_37209,N_37018);
and U37641 (N_37641,N_37065,N_37163);
or U37642 (N_37642,N_37099,N_37443);
xnor U37643 (N_37643,N_37400,N_37466);
nor U37644 (N_37644,N_37000,N_37367);
nand U37645 (N_37645,N_37490,N_37094);
and U37646 (N_37646,N_37063,N_37207);
nand U37647 (N_37647,N_37192,N_37113);
nand U37648 (N_37648,N_37321,N_37023);
nand U37649 (N_37649,N_37175,N_37410);
and U37650 (N_37650,N_37148,N_37399);
nor U37651 (N_37651,N_37098,N_37276);
and U37652 (N_37652,N_37290,N_37043);
and U37653 (N_37653,N_37168,N_37351);
nor U37654 (N_37654,N_37217,N_37002);
or U37655 (N_37655,N_37494,N_37066);
and U37656 (N_37656,N_37422,N_37053);
and U37657 (N_37657,N_37309,N_37455);
xnor U37658 (N_37658,N_37328,N_37304);
nor U37659 (N_37659,N_37030,N_37182);
nor U37660 (N_37660,N_37404,N_37385);
nand U37661 (N_37661,N_37102,N_37006);
nand U37662 (N_37662,N_37009,N_37041);
nand U37663 (N_37663,N_37058,N_37246);
nand U37664 (N_37664,N_37143,N_37330);
nand U37665 (N_37665,N_37474,N_37180);
or U37666 (N_37666,N_37039,N_37236);
nor U37667 (N_37667,N_37391,N_37429);
or U37668 (N_37668,N_37486,N_37131);
and U37669 (N_37669,N_37191,N_37086);
xnor U37670 (N_37670,N_37189,N_37245);
xnor U37671 (N_37671,N_37473,N_37297);
nor U37672 (N_37672,N_37456,N_37056);
and U37673 (N_37673,N_37260,N_37093);
xnor U37674 (N_37674,N_37116,N_37231);
nor U37675 (N_37675,N_37478,N_37496);
or U37676 (N_37676,N_37206,N_37462);
nand U37677 (N_37677,N_37108,N_37435);
or U37678 (N_37678,N_37311,N_37282);
and U37679 (N_37679,N_37360,N_37109);
nor U37680 (N_37680,N_37374,N_37319);
or U37681 (N_37681,N_37268,N_37326);
or U37682 (N_37682,N_37165,N_37269);
nand U37683 (N_37683,N_37008,N_37376);
xnor U37684 (N_37684,N_37177,N_37184);
nand U37685 (N_37685,N_37298,N_37224);
nand U37686 (N_37686,N_37123,N_37334);
or U37687 (N_37687,N_37036,N_37201);
nand U37688 (N_37688,N_37358,N_37128);
nand U37689 (N_37689,N_37415,N_37222);
or U37690 (N_37690,N_37156,N_37439);
nor U37691 (N_37691,N_37359,N_37368);
and U37692 (N_37692,N_37150,N_37369);
nand U37693 (N_37693,N_37145,N_37155);
or U37694 (N_37694,N_37424,N_37482);
nand U37695 (N_37695,N_37232,N_37077);
and U37696 (N_37696,N_37210,N_37280);
nor U37697 (N_37697,N_37355,N_37302);
or U37698 (N_37698,N_37313,N_37026);
nor U37699 (N_37699,N_37463,N_37451);
or U37700 (N_37700,N_37183,N_37204);
or U37701 (N_37701,N_37179,N_37121);
and U37702 (N_37702,N_37375,N_37263);
or U37703 (N_37703,N_37024,N_37338);
nor U37704 (N_37704,N_37178,N_37485);
and U37705 (N_37705,N_37228,N_37170);
and U37706 (N_37706,N_37492,N_37115);
and U37707 (N_37707,N_37100,N_37153);
and U37708 (N_37708,N_37387,N_37481);
nand U37709 (N_37709,N_37174,N_37069);
nand U37710 (N_37710,N_37062,N_37067);
and U37711 (N_37711,N_37046,N_37044);
or U37712 (N_37712,N_37127,N_37181);
nor U37713 (N_37713,N_37437,N_37060);
xnor U37714 (N_37714,N_37031,N_37196);
nor U37715 (N_37715,N_37294,N_37028);
or U37716 (N_37716,N_37331,N_37315);
nor U37717 (N_37717,N_37327,N_37061);
and U37718 (N_37718,N_37010,N_37497);
or U37719 (N_37719,N_37249,N_37022);
and U37720 (N_37720,N_37015,N_37149);
or U37721 (N_37721,N_37337,N_37409);
nor U37722 (N_37722,N_37241,N_37027);
or U37723 (N_37723,N_37134,N_37261);
xor U37724 (N_37724,N_37166,N_37371);
nor U37725 (N_37725,N_37488,N_37342);
and U37726 (N_37726,N_37332,N_37316);
nand U37727 (N_37727,N_37233,N_37499);
or U37728 (N_37728,N_37416,N_37076);
nor U37729 (N_37729,N_37079,N_37458);
and U37730 (N_37730,N_37146,N_37286);
and U37731 (N_37731,N_37350,N_37151);
and U37732 (N_37732,N_37032,N_37270);
nor U37733 (N_37733,N_37211,N_37428);
nor U37734 (N_37734,N_37226,N_37366);
and U37735 (N_37735,N_37495,N_37461);
xor U37736 (N_37736,N_37356,N_37383);
nand U37737 (N_37737,N_37395,N_37308);
xor U37738 (N_37738,N_37203,N_37292);
or U37739 (N_37739,N_37301,N_37445);
nor U37740 (N_37740,N_37377,N_37362);
or U37741 (N_37741,N_37078,N_37402);
or U37742 (N_37742,N_37238,N_37049);
nand U37743 (N_37743,N_37442,N_37464);
nor U37744 (N_37744,N_37081,N_37390);
nand U37745 (N_37745,N_37310,N_37421);
nand U37746 (N_37746,N_37101,N_37347);
and U37747 (N_37747,N_37484,N_37193);
or U37748 (N_37748,N_37434,N_37483);
and U37749 (N_37749,N_37160,N_37291);
nand U37750 (N_37750,N_37354,N_37468);
nor U37751 (N_37751,N_37248,N_37220);
nor U37752 (N_37752,N_37268,N_37016);
and U37753 (N_37753,N_37175,N_37304);
and U37754 (N_37754,N_37395,N_37447);
nor U37755 (N_37755,N_37221,N_37340);
or U37756 (N_37756,N_37231,N_37345);
nor U37757 (N_37757,N_37478,N_37446);
or U37758 (N_37758,N_37178,N_37194);
or U37759 (N_37759,N_37460,N_37408);
nand U37760 (N_37760,N_37492,N_37389);
nor U37761 (N_37761,N_37136,N_37343);
or U37762 (N_37762,N_37308,N_37281);
or U37763 (N_37763,N_37129,N_37123);
and U37764 (N_37764,N_37276,N_37203);
and U37765 (N_37765,N_37041,N_37062);
and U37766 (N_37766,N_37158,N_37097);
nand U37767 (N_37767,N_37190,N_37007);
and U37768 (N_37768,N_37354,N_37075);
and U37769 (N_37769,N_37010,N_37112);
nand U37770 (N_37770,N_37475,N_37411);
or U37771 (N_37771,N_37217,N_37455);
nand U37772 (N_37772,N_37396,N_37023);
nor U37773 (N_37773,N_37058,N_37386);
or U37774 (N_37774,N_37093,N_37312);
nor U37775 (N_37775,N_37071,N_37131);
nor U37776 (N_37776,N_37230,N_37369);
and U37777 (N_37777,N_37097,N_37215);
nand U37778 (N_37778,N_37224,N_37246);
nand U37779 (N_37779,N_37067,N_37025);
and U37780 (N_37780,N_37235,N_37254);
or U37781 (N_37781,N_37292,N_37415);
nand U37782 (N_37782,N_37185,N_37332);
xnor U37783 (N_37783,N_37499,N_37073);
xnor U37784 (N_37784,N_37262,N_37468);
xnor U37785 (N_37785,N_37336,N_37342);
or U37786 (N_37786,N_37311,N_37397);
and U37787 (N_37787,N_37260,N_37282);
nand U37788 (N_37788,N_37281,N_37147);
nor U37789 (N_37789,N_37233,N_37454);
or U37790 (N_37790,N_37422,N_37441);
and U37791 (N_37791,N_37026,N_37398);
nand U37792 (N_37792,N_37280,N_37231);
or U37793 (N_37793,N_37297,N_37191);
xnor U37794 (N_37794,N_37348,N_37198);
nand U37795 (N_37795,N_37150,N_37482);
nand U37796 (N_37796,N_37493,N_37065);
nor U37797 (N_37797,N_37209,N_37449);
or U37798 (N_37798,N_37397,N_37403);
xnor U37799 (N_37799,N_37390,N_37344);
and U37800 (N_37800,N_37093,N_37463);
xnor U37801 (N_37801,N_37306,N_37456);
nor U37802 (N_37802,N_37266,N_37004);
and U37803 (N_37803,N_37088,N_37200);
and U37804 (N_37804,N_37267,N_37060);
and U37805 (N_37805,N_37037,N_37066);
xor U37806 (N_37806,N_37329,N_37064);
or U37807 (N_37807,N_37256,N_37144);
xnor U37808 (N_37808,N_37441,N_37221);
nand U37809 (N_37809,N_37163,N_37261);
xnor U37810 (N_37810,N_37001,N_37462);
or U37811 (N_37811,N_37461,N_37343);
or U37812 (N_37812,N_37218,N_37045);
nand U37813 (N_37813,N_37449,N_37038);
nand U37814 (N_37814,N_37334,N_37300);
xor U37815 (N_37815,N_37167,N_37317);
and U37816 (N_37816,N_37260,N_37239);
and U37817 (N_37817,N_37343,N_37018);
or U37818 (N_37818,N_37431,N_37264);
nor U37819 (N_37819,N_37491,N_37380);
xnor U37820 (N_37820,N_37440,N_37483);
nand U37821 (N_37821,N_37365,N_37322);
nand U37822 (N_37822,N_37207,N_37008);
nor U37823 (N_37823,N_37362,N_37073);
nand U37824 (N_37824,N_37015,N_37171);
nand U37825 (N_37825,N_37008,N_37331);
and U37826 (N_37826,N_37190,N_37477);
or U37827 (N_37827,N_37199,N_37416);
or U37828 (N_37828,N_37394,N_37382);
or U37829 (N_37829,N_37188,N_37165);
or U37830 (N_37830,N_37217,N_37465);
nand U37831 (N_37831,N_37457,N_37209);
or U37832 (N_37832,N_37450,N_37468);
nand U37833 (N_37833,N_37076,N_37382);
and U37834 (N_37834,N_37317,N_37078);
or U37835 (N_37835,N_37028,N_37011);
xor U37836 (N_37836,N_37090,N_37225);
and U37837 (N_37837,N_37449,N_37178);
nand U37838 (N_37838,N_37077,N_37279);
nor U37839 (N_37839,N_37339,N_37220);
nor U37840 (N_37840,N_37255,N_37005);
nand U37841 (N_37841,N_37479,N_37259);
or U37842 (N_37842,N_37343,N_37188);
or U37843 (N_37843,N_37028,N_37418);
and U37844 (N_37844,N_37195,N_37372);
or U37845 (N_37845,N_37043,N_37258);
nand U37846 (N_37846,N_37244,N_37199);
and U37847 (N_37847,N_37250,N_37292);
nand U37848 (N_37848,N_37409,N_37165);
and U37849 (N_37849,N_37435,N_37247);
nor U37850 (N_37850,N_37499,N_37169);
xnor U37851 (N_37851,N_37301,N_37079);
nand U37852 (N_37852,N_37231,N_37027);
or U37853 (N_37853,N_37247,N_37431);
and U37854 (N_37854,N_37396,N_37475);
or U37855 (N_37855,N_37491,N_37240);
or U37856 (N_37856,N_37098,N_37391);
xor U37857 (N_37857,N_37493,N_37269);
or U37858 (N_37858,N_37419,N_37008);
nor U37859 (N_37859,N_37123,N_37095);
or U37860 (N_37860,N_37064,N_37236);
or U37861 (N_37861,N_37236,N_37471);
nand U37862 (N_37862,N_37400,N_37103);
nand U37863 (N_37863,N_37333,N_37491);
or U37864 (N_37864,N_37144,N_37312);
xor U37865 (N_37865,N_37083,N_37441);
nor U37866 (N_37866,N_37494,N_37332);
nor U37867 (N_37867,N_37347,N_37450);
nand U37868 (N_37868,N_37000,N_37136);
and U37869 (N_37869,N_37020,N_37108);
and U37870 (N_37870,N_37440,N_37306);
and U37871 (N_37871,N_37318,N_37111);
nand U37872 (N_37872,N_37186,N_37430);
nor U37873 (N_37873,N_37290,N_37432);
and U37874 (N_37874,N_37158,N_37172);
nor U37875 (N_37875,N_37379,N_37081);
nor U37876 (N_37876,N_37353,N_37018);
nor U37877 (N_37877,N_37010,N_37446);
and U37878 (N_37878,N_37478,N_37424);
nand U37879 (N_37879,N_37081,N_37244);
xnor U37880 (N_37880,N_37154,N_37002);
or U37881 (N_37881,N_37331,N_37403);
or U37882 (N_37882,N_37159,N_37108);
nor U37883 (N_37883,N_37232,N_37020);
or U37884 (N_37884,N_37112,N_37470);
nand U37885 (N_37885,N_37062,N_37381);
or U37886 (N_37886,N_37158,N_37031);
nand U37887 (N_37887,N_37395,N_37423);
nand U37888 (N_37888,N_37495,N_37335);
and U37889 (N_37889,N_37128,N_37426);
nand U37890 (N_37890,N_37213,N_37253);
or U37891 (N_37891,N_37098,N_37153);
and U37892 (N_37892,N_37335,N_37156);
or U37893 (N_37893,N_37195,N_37348);
nand U37894 (N_37894,N_37032,N_37194);
nand U37895 (N_37895,N_37217,N_37039);
or U37896 (N_37896,N_37382,N_37167);
or U37897 (N_37897,N_37352,N_37366);
or U37898 (N_37898,N_37231,N_37239);
nand U37899 (N_37899,N_37415,N_37124);
nor U37900 (N_37900,N_37162,N_37461);
and U37901 (N_37901,N_37481,N_37459);
and U37902 (N_37902,N_37443,N_37496);
or U37903 (N_37903,N_37202,N_37185);
xnor U37904 (N_37904,N_37343,N_37453);
xor U37905 (N_37905,N_37379,N_37198);
and U37906 (N_37906,N_37395,N_37307);
nand U37907 (N_37907,N_37292,N_37251);
or U37908 (N_37908,N_37299,N_37075);
and U37909 (N_37909,N_37486,N_37238);
and U37910 (N_37910,N_37055,N_37124);
and U37911 (N_37911,N_37185,N_37174);
and U37912 (N_37912,N_37286,N_37336);
and U37913 (N_37913,N_37213,N_37286);
and U37914 (N_37914,N_37479,N_37226);
nand U37915 (N_37915,N_37330,N_37215);
and U37916 (N_37916,N_37030,N_37436);
nor U37917 (N_37917,N_37284,N_37120);
nand U37918 (N_37918,N_37436,N_37403);
nor U37919 (N_37919,N_37155,N_37382);
or U37920 (N_37920,N_37411,N_37429);
or U37921 (N_37921,N_37218,N_37120);
nor U37922 (N_37922,N_37213,N_37086);
nand U37923 (N_37923,N_37102,N_37150);
and U37924 (N_37924,N_37173,N_37053);
nor U37925 (N_37925,N_37417,N_37236);
and U37926 (N_37926,N_37014,N_37124);
or U37927 (N_37927,N_37288,N_37115);
nand U37928 (N_37928,N_37168,N_37223);
or U37929 (N_37929,N_37207,N_37062);
nand U37930 (N_37930,N_37185,N_37078);
nor U37931 (N_37931,N_37279,N_37422);
or U37932 (N_37932,N_37087,N_37311);
xor U37933 (N_37933,N_37117,N_37145);
and U37934 (N_37934,N_37177,N_37210);
and U37935 (N_37935,N_37351,N_37299);
nor U37936 (N_37936,N_37181,N_37488);
and U37937 (N_37937,N_37485,N_37037);
nor U37938 (N_37938,N_37020,N_37270);
nor U37939 (N_37939,N_37240,N_37410);
nand U37940 (N_37940,N_37153,N_37143);
and U37941 (N_37941,N_37107,N_37003);
and U37942 (N_37942,N_37277,N_37360);
and U37943 (N_37943,N_37227,N_37484);
and U37944 (N_37944,N_37287,N_37164);
or U37945 (N_37945,N_37289,N_37390);
or U37946 (N_37946,N_37034,N_37326);
nand U37947 (N_37947,N_37278,N_37006);
nand U37948 (N_37948,N_37465,N_37376);
and U37949 (N_37949,N_37446,N_37229);
nand U37950 (N_37950,N_37124,N_37409);
or U37951 (N_37951,N_37427,N_37014);
nand U37952 (N_37952,N_37401,N_37008);
or U37953 (N_37953,N_37004,N_37470);
xor U37954 (N_37954,N_37283,N_37004);
and U37955 (N_37955,N_37091,N_37142);
and U37956 (N_37956,N_37143,N_37284);
or U37957 (N_37957,N_37179,N_37023);
nor U37958 (N_37958,N_37070,N_37167);
or U37959 (N_37959,N_37357,N_37457);
or U37960 (N_37960,N_37260,N_37139);
nor U37961 (N_37961,N_37383,N_37306);
nor U37962 (N_37962,N_37229,N_37434);
nor U37963 (N_37963,N_37148,N_37277);
or U37964 (N_37964,N_37135,N_37301);
nor U37965 (N_37965,N_37174,N_37383);
and U37966 (N_37966,N_37028,N_37344);
xnor U37967 (N_37967,N_37173,N_37163);
nor U37968 (N_37968,N_37183,N_37417);
and U37969 (N_37969,N_37122,N_37182);
or U37970 (N_37970,N_37205,N_37268);
nand U37971 (N_37971,N_37425,N_37423);
and U37972 (N_37972,N_37257,N_37285);
nand U37973 (N_37973,N_37340,N_37194);
nor U37974 (N_37974,N_37456,N_37104);
or U37975 (N_37975,N_37157,N_37197);
nor U37976 (N_37976,N_37131,N_37408);
or U37977 (N_37977,N_37405,N_37491);
and U37978 (N_37978,N_37346,N_37022);
nand U37979 (N_37979,N_37440,N_37148);
nor U37980 (N_37980,N_37153,N_37151);
xnor U37981 (N_37981,N_37466,N_37430);
or U37982 (N_37982,N_37239,N_37192);
and U37983 (N_37983,N_37107,N_37386);
nand U37984 (N_37984,N_37161,N_37423);
or U37985 (N_37985,N_37302,N_37284);
xor U37986 (N_37986,N_37137,N_37489);
and U37987 (N_37987,N_37033,N_37128);
nor U37988 (N_37988,N_37391,N_37462);
nand U37989 (N_37989,N_37424,N_37416);
nand U37990 (N_37990,N_37012,N_37464);
nand U37991 (N_37991,N_37400,N_37462);
nand U37992 (N_37992,N_37212,N_37324);
or U37993 (N_37993,N_37148,N_37052);
nand U37994 (N_37994,N_37421,N_37380);
nor U37995 (N_37995,N_37136,N_37163);
nor U37996 (N_37996,N_37125,N_37303);
nor U37997 (N_37997,N_37083,N_37054);
xor U37998 (N_37998,N_37245,N_37366);
and U37999 (N_37999,N_37087,N_37330);
and U38000 (N_38000,N_37639,N_37763);
nor U38001 (N_38001,N_37783,N_37928);
or U38002 (N_38002,N_37730,N_37883);
nand U38003 (N_38003,N_37696,N_37732);
and U38004 (N_38004,N_37669,N_37784);
nor U38005 (N_38005,N_37720,N_37515);
nor U38006 (N_38006,N_37907,N_37828);
and U38007 (N_38007,N_37504,N_37864);
nor U38008 (N_38008,N_37599,N_37704);
or U38009 (N_38009,N_37586,N_37935);
nor U38010 (N_38010,N_37653,N_37826);
or U38011 (N_38011,N_37874,N_37633);
and U38012 (N_38012,N_37713,N_37844);
nand U38013 (N_38013,N_37718,N_37894);
nor U38014 (N_38014,N_37862,N_37878);
xnor U38015 (N_38015,N_37535,N_37646);
or U38016 (N_38016,N_37758,N_37970);
nand U38017 (N_38017,N_37792,N_37789);
and U38018 (N_38018,N_37772,N_37742);
nand U38019 (N_38019,N_37971,N_37904);
xor U38020 (N_38020,N_37965,N_37906);
nor U38021 (N_38021,N_37961,N_37505);
nor U38022 (N_38022,N_37807,N_37652);
nand U38023 (N_38023,N_37649,N_37876);
and U38024 (N_38024,N_37525,N_37825);
nand U38025 (N_38025,N_37921,N_37985);
nand U38026 (N_38026,N_37725,N_37848);
and U38027 (N_38027,N_37684,N_37685);
or U38028 (N_38028,N_37542,N_37768);
and U38029 (N_38029,N_37637,N_37788);
nor U38030 (N_38030,N_37818,N_37700);
nand U38031 (N_38031,N_37994,N_37714);
nor U38032 (N_38032,N_37527,N_37560);
and U38033 (N_38033,N_37645,N_37659);
xor U38034 (N_38034,N_37651,N_37990);
nor U38035 (N_38035,N_37621,N_37954);
and U38036 (N_38036,N_37899,N_37889);
nand U38037 (N_38037,N_37623,N_37592);
nand U38038 (N_38038,N_37922,N_37891);
xnor U38039 (N_38039,N_37740,N_37625);
xnor U38040 (N_38040,N_37723,N_37948);
nor U38041 (N_38041,N_37810,N_37748);
nand U38042 (N_38042,N_37642,N_37927);
and U38043 (N_38043,N_37752,N_37692);
nor U38044 (N_38044,N_37983,N_37664);
nor U38045 (N_38045,N_37829,N_37675);
and U38046 (N_38046,N_37967,N_37538);
nor U38047 (N_38047,N_37662,N_37676);
nor U38048 (N_38048,N_37885,N_37850);
and U38049 (N_38049,N_37902,N_37608);
nor U38050 (N_38050,N_37619,N_37524);
nand U38051 (N_38051,N_37981,N_37607);
nand U38052 (N_38052,N_37979,N_37797);
or U38053 (N_38053,N_37877,N_37531);
nand U38054 (N_38054,N_37544,N_37936);
or U38055 (N_38055,N_37736,N_37701);
or U38056 (N_38056,N_37728,N_37762);
and U38057 (N_38057,N_37968,N_37931);
nor U38058 (N_38058,N_37916,N_37858);
nand U38059 (N_38059,N_37791,N_37893);
nor U38060 (N_38060,N_37629,N_37579);
or U38061 (N_38061,N_37521,N_37978);
or U38062 (N_38062,N_37919,N_37787);
nand U38063 (N_38063,N_37947,N_37860);
or U38064 (N_38064,N_37924,N_37707);
and U38065 (N_38065,N_37849,N_37754);
or U38066 (N_38066,N_37604,N_37972);
nor U38067 (N_38067,N_37612,N_37926);
or U38068 (N_38068,N_37843,N_37838);
or U38069 (N_38069,N_37562,N_37749);
and U38070 (N_38070,N_37753,N_37566);
xor U38071 (N_38071,N_37512,N_37903);
and U38072 (N_38072,N_37563,N_37991);
nor U38073 (N_38073,N_37875,N_37997);
nand U38074 (N_38074,N_37678,N_37568);
and U38075 (N_38075,N_37811,N_37949);
and U38076 (N_38076,N_37553,N_37613);
nand U38077 (N_38077,N_37995,N_37945);
and U38078 (N_38078,N_37594,N_37816);
and U38079 (N_38079,N_37672,N_37556);
nand U38080 (N_38080,N_37577,N_37661);
or U38081 (N_38081,N_37522,N_37694);
and U38082 (N_38082,N_37636,N_37695);
and U38083 (N_38083,N_37564,N_37782);
and U38084 (N_38084,N_37777,N_37630);
nand U38085 (N_38085,N_37781,N_37969);
and U38086 (N_38086,N_37729,N_37999);
nand U38087 (N_38087,N_37790,N_37955);
xnor U38088 (N_38088,N_37510,N_37745);
and U38089 (N_38089,N_37809,N_37832);
xnor U38090 (N_38090,N_37541,N_37833);
nand U38091 (N_38091,N_37799,N_37548);
nand U38092 (N_38092,N_37744,N_37958);
or U38093 (N_38093,N_37666,N_37567);
or U38094 (N_38094,N_37549,N_37731);
or U38095 (N_38095,N_37658,N_37598);
nand U38096 (N_38096,N_37712,N_37839);
nor U38097 (N_38097,N_37561,N_37980);
nor U38098 (N_38098,N_37973,N_37546);
nand U38099 (N_38099,N_37721,N_37528);
and U38100 (N_38100,N_37974,N_37640);
nand U38101 (N_38101,N_37545,N_37866);
and U38102 (N_38102,N_37892,N_37603);
nand U38103 (N_38103,N_37670,N_37609);
or U38104 (N_38104,N_37942,N_37778);
or U38105 (N_38105,N_37509,N_37761);
and U38106 (N_38106,N_37727,N_37517);
and U38107 (N_38107,N_37911,N_37737);
or U38108 (N_38108,N_37890,N_37597);
nand U38109 (N_38109,N_37845,N_37726);
nor U38110 (N_38110,N_37870,N_37932);
and U38111 (N_38111,N_37526,N_37764);
or U38112 (N_38112,N_37815,N_37993);
or U38113 (N_38113,N_37508,N_37578);
xnor U38114 (N_38114,N_37937,N_37705);
and U38115 (N_38115,N_37532,N_37741);
nor U38116 (N_38116,N_37677,N_37998);
nand U38117 (N_38117,N_37767,N_37626);
nor U38118 (N_38118,N_37668,N_37536);
or U38119 (N_38119,N_37984,N_37638);
nand U38120 (N_38120,N_37812,N_37596);
and U38121 (N_38121,N_37751,N_37831);
xnor U38122 (N_38122,N_37715,N_37618);
nand U38123 (N_38123,N_37909,N_37801);
xnor U38124 (N_38124,N_37861,N_37632);
or U38125 (N_38125,N_37939,N_37855);
nor U38126 (N_38126,N_37750,N_37952);
nor U38127 (N_38127,N_37755,N_37820);
nand U38128 (N_38128,N_37837,N_37550);
nor U38129 (N_38129,N_37863,N_37688);
nand U38130 (N_38130,N_37614,N_37895);
nor U38131 (N_38131,N_37882,N_37734);
nand U38132 (N_38132,N_37709,N_37940);
or U38133 (N_38133,N_37600,N_37769);
or U38134 (N_38134,N_37773,N_37643);
and U38135 (N_38135,N_37582,N_37519);
nand U38136 (N_38136,N_37917,N_37591);
and U38137 (N_38137,N_37827,N_37756);
and U38138 (N_38138,N_37933,N_37690);
or U38139 (N_38139,N_37836,N_37975);
or U38140 (N_38140,N_37765,N_37691);
or U38141 (N_38141,N_37501,N_37610);
and U38142 (N_38142,N_37842,N_37918);
or U38143 (N_38143,N_37667,N_37552);
and U38144 (N_38144,N_37996,N_37823);
or U38145 (N_38145,N_37914,N_37905);
nand U38146 (N_38146,N_37533,N_37840);
or U38147 (N_38147,N_37779,N_37795);
or U38148 (N_38148,N_37500,N_37898);
xor U38149 (N_38149,N_37571,N_37558);
or U38150 (N_38150,N_37957,N_37681);
or U38151 (N_38151,N_37956,N_37655);
nand U38152 (N_38152,N_37516,N_37786);
or U38153 (N_38153,N_37941,N_37554);
xor U38154 (N_38154,N_37605,N_37648);
or U38155 (N_38155,N_37798,N_37513);
and U38156 (N_38156,N_37673,N_37853);
nand U38157 (N_38157,N_37938,N_37951);
xnor U38158 (N_38158,N_37910,N_37775);
nand U38159 (N_38159,N_37506,N_37627);
and U38160 (N_38160,N_37766,N_37593);
and U38161 (N_38161,N_37869,N_37835);
or U38162 (N_38162,N_37871,N_37539);
nand U38163 (N_38163,N_37915,N_37682);
and U38164 (N_38164,N_37817,N_37735);
and U38165 (N_38165,N_37929,N_37896);
nor U38166 (N_38166,N_37803,N_37529);
and U38167 (N_38167,N_37872,N_37628);
and U38168 (N_38168,N_37588,N_37986);
nand U38169 (N_38169,N_37551,N_37644);
or U38170 (N_38170,N_37540,N_37846);
nor U38171 (N_38171,N_37616,N_37654);
or U38172 (N_38172,N_37583,N_37759);
nand U38173 (N_38173,N_37617,N_37834);
xor U38174 (N_38174,N_37988,N_37534);
xnor U38175 (N_38175,N_37572,N_37717);
nand U38176 (N_38176,N_37887,N_37523);
and U38177 (N_38177,N_37857,N_37689);
and U38178 (N_38178,N_37770,N_37511);
xnor U38179 (N_38179,N_37964,N_37854);
or U38180 (N_38180,N_37913,N_37602);
or U38181 (N_38181,N_37960,N_37514);
nor U38182 (N_38182,N_37879,N_37587);
nor U38183 (N_38183,N_37865,N_37635);
nor U38184 (N_38184,N_37611,N_37868);
or U38185 (N_38185,N_37747,N_37719);
and U38186 (N_38186,N_37706,N_37698);
and U38187 (N_38187,N_37992,N_37543);
or U38188 (N_38188,N_37581,N_37656);
or U38189 (N_38189,N_37589,N_37841);
xnor U38190 (N_38190,N_37738,N_37859);
nand U38191 (N_38191,N_37650,N_37743);
xnor U38192 (N_38192,N_37520,N_37912);
and U38193 (N_38193,N_37760,N_37813);
and U38194 (N_38194,N_37590,N_37557);
nor U38195 (N_38195,N_37805,N_37989);
and U38196 (N_38196,N_37873,N_37663);
and U38197 (N_38197,N_37923,N_37697);
and U38198 (N_38198,N_37780,N_37606);
nand U38199 (N_38199,N_37674,N_37710);
nand U38200 (N_38200,N_37722,N_37953);
nand U38201 (N_38201,N_37819,N_37950);
and U38202 (N_38202,N_37641,N_37555);
or U38203 (N_38203,N_37699,N_37631);
nand U38204 (N_38204,N_37822,N_37507);
nand U38205 (N_38205,N_37518,N_37615);
and U38206 (N_38206,N_37852,N_37679);
nor U38207 (N_38207,N_37576,N_37595);
nor U38208 (N_38208,N_37647,N_37897);
or U38209 (N_38209,N_37806,N_37962);
and U38210 (N_38210,N_37908,N_37944);
and U38211 (N_38211,N_37794,N_37702);
or U38212 (N_38212,N_37585,N_37982);
nor U38213 (N_38213,N_37601,N_37537);
nand U38214 (N_38214,N_37693,N_37793);
or U38215 (N_38215,N_37884,N_37776);
or U38216 (N_38216,N_37821,N_37796);
and U38217 (N_38217,N_37569,N_37671);
nand U38218 (N_38218,N_37660,N_37665);
nor U38219 (N_38219,N_37943,N_37624);
and U38220 (N_38220,N_37934,N_37502);
and U38221 (N_38221,N_37930,N_37867);
xnor U38222 (N_38222,N_37503,N_37771);
and U38223 (N_38223,N_37620,N_37856);
nand U38224 (N_38224,N_37757,N_37976);
or U38225 (N_38225,N_37724,N_37959);
or U38226 (N_38226,N_37963,N_37739);
nor U38227 (N_38227,N_37687,N_37683);
and U38228 (N_38228,N_37565,N_37886);
nor U38229 (N_38229,N_37733,N_37580);
nand U38230 (N_38230,N_37851,N_37622);
or U38231 (N_38231,N_37746,N_37824);
and U38232 (N_38232,N_37711,N_37530);
or U38233 (N_38233,N_37977,N_37901);
nand U38234 (N_38234,N_37703,N_37847);
xnor U38235 (N_38235,N_37946,N_37634);
and U38236 (N_38236,N_37657,N_37966);
nor U38237 (N_38237,N_37880,N_37774);
or U38238 (N_38238,N_37925,N_37716);
or U38239 (N_38239,N_37547,N_37559);
xnor U38240 (N_38240,N_37573,N_37804);
xnor U38241 (N_38241,N_37800,N_37584);
xor U38242 (N_38242,N_37575,N_37686);
nor U38243 (N_38243,N_37814,N_37802);
nand U38244 (N_38244,N_37808,N_37574);
or U38245 (N_38245,N_37987,N_37785);
or U38246 (N_38246,N_37830,N_37570);
and U38247 (N_38247,N_37680,N_37920);
and U38248 (N_38248,N_37900,N_37881);
nor U38249 (N_38249,N_37888,N_37708);
xor U38250 (N_38250,N_37936,N_37800);
nor U38251 (N_38251,N_37893,N_37977);
nor U38252 (N_38252,N_37887,N_37989);
nor U38253 (N_38253,N_37806,N_37588);
or U38254 (N_38254,N_37884,N_37619);
nand U38255 (N_38255,N_37944,N_37967);
and U38256 (N_38256,N_37947,N_37803);
or U38257 (N_38257,N_37772,N_37620);
nand U38258 (N_38258,N_37550,N_37919);
nor U38259 (N_38259,N_37736,N_37710);
or U38260 (N_38260,N_37674,N_37697);
and U38261 (N_38261,N_37880,N_37860);
nor U38262 (N_38262,N_37863,N_37589);
or U38263 (N_38263,N_37962,N_37567);
nand U38264 (N_38264,N_37856,N_37845);
and U38265 (N_38265,N_37788,N_37830);
and U38266 (N_38266,N_37520,N_37603);
or U38267 (N_38267,N_37757,N_37844);
nor U38268 (N_38268,N_37595,N_37730);
nand U38269 (N_38269,N_37600,N_37504);
nor U38270 (N_38270,N_37759,N_37641);
nand U38271 (N_38271,N_37508,N_37561);
and U38272 (N_38272,N_37635,N_37875);
and U38273 (N_38273,N_37998,N_37949);
nor U38274 (N_38274,N_37827,N_37731);
nand U38275 (N_38275,N_37707,N_37755);
or U38276 (N_38276,N_37633,N_37530);
nand U38277 (N_38277,N_37587,N_37785);
or U38278 (N_38278,N_37717,N_37834);
or U38279 (N_38279,N_37646,N_37769);
nand U38280 (N_38280,N_37570,N_37810);
nor U38281 (N_38281,N_37939,N_37741);
and U38282 (N_38282,N_37547,N_37676);
and U38283 (N_38283,N_37649,N_37808);
nand U38284 (N_38284,N_37978,N_37998);
nor U38285 (N_38285,N_37934,N_37890);
and U38286 (N_38286,N_37548,N_37666);
or U38287 (N_38287,N_37626,N_37954);
or U38288 (N_38288,N_37951,N_37907);
xnor U38289 (N_38289,N_37589,N_37885);
or U38290 (N_38290,N_37652,N_37610);
or U38291 (N_38291,N_37791,N_37655);
nand U38292 (N_38292,N_37953,N_37519);
nor U38293 (N_38293,N_37596,N_37813);
or U38294 (N_38294,N_37829,N_37640);
xnor U38295 (N_38295,N_37571,N_37772);
and U38296 (N_38296,N_37954,N_37956);
nand U38297 (N_38297,N_37992,N_37931);
and U38298 (N_38298,N_37559,N_37833);
xor U38299 (N_38299,N_37648,N_37703);
or U38300 (N_38300,N_37873,N_37884);
and U38301 (N_38301,N_37838,N_37712);
nor U38302 (N_38302,N_37876,N_37828);
nand U38303 (N_38303,N_37552,N_37531);
nand U38304 (N_38304,N_37925,N_37502);
and U38305 (N_38305,N_37792,N_37946);
nor U38306 (N_38306,N_37739,N_37851);
nand U38307 (N_38307,N_37922,N_37690);
xnor U38308 (N_38308,N_37514,N_37705);
nand U38309 (N_38309,N_37581,N_37807);
nor U38310 (N_38310,N_37505,N_37841);
and U38311 (N_38311,N_37756,N_37607);
xor U38312 (N_38312,N_37791,N_37577);
or U38313 (N_38313,N_37795,N_37891);
and U38314 (N_38314,N_37922,N_37862);
nand U38315 (N_38315,N_37588,N_37782);
nand U38316 (N_38316,N_37837,N_37790);
or U38317 (N_38317,N_37694,N_37585);
or U38318 (N_38318,N_37996,N_37594);
nor U38319 (N_38319,N_37542,N_37620);
or U38320 (N_38320,N_37539,N_37750);
or U38321 (N_38321,N_37704,N_37819);
nand U38322 (N_38322,N_37821,N_37856);
nand U38323 (N_38323,N_37792,N_37985);
or U38324 (N_38324,N_37836,N_37942);
nand U38325 (N_38325,N_37604,N_37575);
and U38326 (N_38326,N_37784,N_37632);
xor U38327 (N_38327,N_37953,N_37885);
or U38328 (N_38328,N_37670,N_37574);
and U38329 (N_38329,N_37772,N_37815);
and U38330 (N_38330,N_37545,N_37805);
nor U38331 (N_38331,N_37953,N_37603);
nand U38332 (N_38332,N_37700,N_37744);
nor U38333 (N_38333,N_37793,N_37812);
nand U38334 (N_38334,N_37572,N_37634);
or U38335 (N_38335,N_37726,N_37772);
nand U38336 (N_38336,N_37981,N_37562);
nor U38337 (N_38337,N_37867,N_37917);
xor U38338 (N_38338,N_37898,N_37874);
nand U38339 (N_38339,N_37909,N_37611);
or U38340 (N_38340,N_37987,N_37687);
nor U38341 (N_38341,N_37736,N_37589);
nor U38342 (N_38342,N_37777,N_37919);
or U38343 (N_38343,N_37974,N_37788);
nor U38344 (N_38344,N_37818,N_37691);
or U38345 (N_38345,N_37511,N_37936);
or U38346 (N_38346,N_37957,N_37871);
and U38347 (N_38347,N_37801,N_37735);
nand U38348 (N_38348,N_37849,N_37936);
or U38349 (N_38349,N_37860,N_37591);
and U38350 (N_38350,N_37522,N_37555);
nor U38351 (N_38351,N_37849,N_37948);
and U38352 (N_38352,N_37836,N_37563);
or U38353 (N_38353,N_37973,N_37840);
or U38354 (N_38354,N_37757,N_37503);
xor U38355 (N_38355,N_37559,N_37947);
nor U38356 (N_38356,N_37757,N_37702);
nand U38357 (N_38357,N_37608,N_37668);
nand U38358 (N_38358,N_37746,N_37725);
or U38359 (N_38359,N_37913,N_37981);
and U38360 (N_38360,N_37799,N_37671);
xor U38361 (N_38361,N_37523,N_37643);
and U38362 (N_38362,N_37652,N_37677);
or U38363 (N_38363,N_37975,N_37654);
nor U38364 (N_38364,N_37665,N_37563);
and U38365 (N_38365,N_37749,N_37929);
or U38366 (N_38366,N_37832,N_37764);
xnor U38367 (N_38367,N_37786,N_37753);
nand U38368 (N_38368,N_37745,N_37685);
nand U38369 (N_38369,N_37507,N_37542);
or U38370 (N_38370,N_37958,N_37933);
or U38371 (N_38371,N_37569,N_37660);
and U38372 (N_38372,N_37741,N_37962);
or U38373 (N_38373,N_37586,N_37745);
nand U38374 (N_38374,N_37752,N_37884);
xnor U38375 (N_38375,N_37732,N_37979);
or U38376 (N_38376,N_37869,N_37673);
or U38377 (N_38377,N_37737,N_37656);
nor U38378 (N_38378,N_37813,N_37914);
nor U38379 (N_38379,N_37686,N_37664);
nand U38380 (N_38380,N_37645,N_37649);
nor U38381 (N_38381,N_37922,N_37542);
and U38382 (N_38382,N_37514,N_37726);
xor U38383 (N_38383,N_37895,N_37716);
and U38384 (N_38384,N_37809,N_37695);
and U38385 (N_38385,N_37713,N_37674);
and U38386 (N_38386,N_37711,N_37606);
or U38387 (N_38387,N_37959,N_37773);
nand U38388 (N_38388,N_37975,N_37911);
nand U38389 (N_38389,N_37714,N_37621);
and U38390 (N_38390,N_37526,N_37786);
nor U38391 (N_38391,N_37653,N_37571);
and U38392 (N_38392,N_37684,N_37800);
nor U38393 (N_38393,N_37505,N_37587);
or U38394 (N_38394,N_37519,N_37913);
nor U38395 (N_38395,N_37911,N_37645);
nand U38396 (N_38396,N_37575,N_37694);
or U38397 (N_38397,N_37920,N_37552);
nand U38398 (N_38398,N_37904,N_37786);
xor U38399 (N_38399,N_37869,N_37528);
or U38400 (N_38400,N_37926,N_37983);
or U38401 (N_38401,N_37581,N_37684);
nand U38402 (N_38402,N_37971,N_37696);
or U38403 (N_38403,N_37993,N_37707);
nand U38404 (N_38404,N_37692,N_37572);
nor U38405 (N_38405,N_37908,N_37572);
xor U38406 (N_38406,N_37933,N_37560);
and U38407 (N_38407,N_37906,N_37901);
nor U38408 (N_38408,N_37627,N_37871);
or U38409 (N_38409,N_37881,N_37960);
and U38410 (N_38410,N_37809,N_37710);
or U38411 (N_38411,N_37904,N_37587);
nand U38412 (N_38412,N_37640,N_37914);
nand U38413 (N_38413,N_37982,N_37805);
nand U38414 (N_38414,N_37551,N_37736);
or U38415 (N_38415,N_37657,N_37704);
xor U38416 (N_38416,N_37523,N_37824);
and U38417 (N_38417,N_37548,N_37755);
nor U38418 (N_38418,N_37553,N_37590);
or U38419 (N_38419,N_37701,N_37663);
nand U38420 (N_38420,N_37854,N_37984);
or U38421 (N_38421,N_37837,N_37602);
nand U38422 (N_38422,N_37517,N_37796);
or U38423 (N_38423,N_37608,N_37548);
and U38424 (N_38424,N_37591,N_37936);
or U38425 (N_38425,N_37559,N_37750);
and U38426 (N_38426,N_37827,N_37715);
and U38427 (N_38427,N_37993,N_37973);
nor U38428 (N_38428,N_37811,N_37674);
or U38429 (N_38429,N_37999,N_37899);
nand U38430 (N_38430,N_37974,N_37835);
and U38431 (N_38431,N_37874,N_37881);
and U38432 (N_38432,N_37898,N_37523);
or U38433 (N_38433,N_37808,N_37775);
nor U38434 (N_38434,N_37684,N_37539);
and U38435 (N_38435,N_37822,N_37794);
or U38436 (N_38436,N_37595,N_37956);
and U38437 (N_38437,N_37762,N_37834);
and U38438 (N_38438,N_37825,N_37554);
nand U38439 (N_38439,N_37531,N_37920);
or U38440 (N_38440,N_37526,N_37979);
nor U38441 (N_38441,N_37583,N_37991);
nand U38442 (N_38442,N_37881,N_37895);
nand U38443 (N_38443,N_37770,N_37925);
or U38444 (N_38444,N_37668,N_37564);
xor U38445 (N_38445,N_37927,N_37920);
nand U38446 (N_38446,N_37518,N_37768);
nand U38447 (N_38447,N_37937,N_37598);
nand U38448 (N_38448,N_37635,N_37798);
and U38449 (N_38449,N_37721,N_37966);
nor U38450 (N_38450,N_37992,N_37742);
nand U38451 (N_38451,N_37897,N_37913);
nor U38452 (N_38452,N_37814,N_37819);
and U38453 (N_38453,N_37881,N_37977);
or U38454 (N_38454,N_37858,N_37569);
nand U38455 (N_38455,N_37658,N_37851);
xor U38456 (N_38456,N_37910,N_37840);
xor U38457 (N_38457,N_37695,N_37909);
or U38458 (N_38458,N_37855,N_37969);
or U38459 (N_38459,N_37842,N_37732);
and U38460 (N_38460,N_37903,N_37836);
nor U38461 (N_38461,N_37594,N_37591);
and U38462 (N_38462,N_37667,N_37823);
nand U38463 (N_38463,N_37904,N_37547);
and U38464 (N_38464,N_37601,N_37793);
and U38465 (N_38465,N_37994,N_37573);
and U38466 (N_38466,N_37900,N_37864);
and U38467 (N_38467,N_37722,N_37653);
or U38468 (N_38468,N_37958,N_37560);
nor U38469 (N_38469,N_37607,N_37564);
and U38470 (N_38470,N_37969,N_37733);
or U38471 (N_38471,N_37655,N_37521);
and U38472 (N_38472,N_37900,N_37558);
and U38473 (N_38473,N_37819,N_37625);
nor U38474 (N_38474,N_37528,N_37581);
and U38475 (N_38475,N_37685,N_37833);
nand U38476 (N_38476,N_37652,N_37502);
or U38477 (N_38477,N_37925,N_37777);
nand U38478 (N_38478,N_37864,N_37576);
nor U38479 (N_38479,N_37597,N_37514);
nor U38480 (N_38480,N_37582,N_37783);
nor U38481 (N_38481,N_37609,N_37887);
nor U38482 (N_38482,N_37676,N_37534);
and U38483 (N_38483,N_37951,N_37646);
and U38484 (N_38484,N_37717,N_37817);
and U38485 (N_38485,N_37733,N_37649);
or U38486 (N_38486,N_37974,N_37643);
nor U38487 (N_38487,N_37741,N_37775);
nand U38488 (N_38488,N_37946,N_37570);
nor U38489 (N_38489,N_37505,N_37819);
nor U38490 (N_38490,N_37715,N_37881);
and U38491 (N_38491,N_37907,N_37723);
nor U38492 (N_38492,N_37952,N_37690);
and U38493 (N_38493,N_37818,N_37719);
or U38494 (N_38494,N_37830,N_37692);
nand U38495 (N_38495,N_37558,N_37689);
and U38496 (N_38496,N_37902,N_37988);
nor U38497 (N_38497,N_37921,N_37639);
and U38498 (N_38498,N_37577,N_37783);
xnor U38499 (N_38499,N_37759,N_37635);
and U38500 (N_38500,N_38269,N_38299);
or U38501 (N_38501,N_38079,N_38489);
and U38502 (N_38502,N_38128,N_38172);
and U38503 (N_38503,N_38228,N_38349);
or U38504 (N_38504,N_38167,N_38458);
or U38505 (N_38505,N_38445,N_38483);
nand U38506 (N_38506,N_38036,N_38065);
nand U38507 (N_38507,N_38005,N_38461);
and U38508 (N_38508,N_38348,N_38108);
or U38509 (N_38509,N_38045,N_38278);
nor U38510 (N_38510,N_38055,N_38466);
and U38511 (N_38511,N_38161,N_38311);
nand U38512 (N_38512,N_38424,N_38366);
and U38513 (N_38513,N_38451,N_38460);
nor U38514 (N_38514,N_38174,N_38314);
nor U38515 (N_38515,N_38485,N_38302);
or U38516 (N_38516,N_38277,N_38417);
nor U38517 (N_38517,N_38064,N_38247);
nor U38518 (N_38518,N_38390,N_38257);
nor U38519 (N_38519,N_38249,N_38238);
nor U38520 (N_38520,N_38153,N_38215);
nand U38521 (N_38521,N_38450,N_38355);
and U38522 (N_38522,N_38404,N_38300);
or U38523 (N_38523,N_38356,N_38431);
nand U38524 (N_38524,N_38075,N_38376);
nand U38525 (N_38525,N_38180,N_38041);
nor U38526 (N_38526,N_38371,N_38114);
nor U38527 (N_38527,N_38382,N_38230);
and U38528 (N_38528,N_38132,N_38321);
nand U38529 (N_38529,N_38234,N_38429);
nand U38530 (N_38530,N_38198,N_38194);
and U38531 (N_38531,N_38202,N_38177);
nor U38532 (N_38532,N_38140,N_38059);
and U38533 (N_38533,N_38078,N_38393);
or U38534 (N_38534,N_38354,N_38440);
nand U38535 (N_38535,N_38439,N_38057);
or U38536 (N_38536,N_38329,N_38490);
nor U38537 (N_38537,N_38368,N_38038);
nand U38538 (N_38538,N_38492,N_38449);
and U38539 (N_38539,N_38255,N_38345);
nor U38540 (N_38540,N_38120,N_38350);
and U38541 (N_38541,N_38318,N_38124);
and U38542 (N_38542,N_38015,N_38465);
and U38543 (N_38543,N_38373,N_38009);
nand U38544 (N_38544,N_38474,N_38284);
and U38545 (N_38545,N_38040,N_38452);
and U38546 (N_38546,N_38491,N_38205);
nand U38547 (N_38547,N_38006,N_38496);
nor U38548 (N_38548,N_38196,N_38096);
nand U38549 (N_38549,N_38233,N_38054);
nand U38550 (N_38550,N_38212,N_38332);
and U38551 (N_38551,N_38358,N_38438);
and U38552 (N_38552,N_38080,N_38051);
or U38553 (N_38553,N_38187,N_38229);
nand U38554 (N_38554,N_38303,N_38252);
and U38555 (N_38555,N_38024,N_38346);
nand U38556 (N_38556,N_38216,N_38169);
or U38557 (N_38557,N_38105,N_38495);
nor U38558 (N_38558,N_38192,N_38432);
or U38559 (N_38559,N_38185,N_38218);
or U38560 (N_38560,N_38135,N_38068);
or U38561 (N_38561,N_38004,N_38082);
nor U38562 (N_38562,N_38282,N_38372);
or U38563 (N_38563,N_38377,N_38408);
nand U38564 (N_38564,N_38352,N_38443);
nor U38565 (N_38565,N_38281,N_38103);
and U38566 (N_38566,N_38179,N_38220);
xnor U38567 (N_38567,N_38034,N_38428);
nor U38568 (N_38568,N_38025,N_38046);
or U38569 (N_38569,N_38239,N_38380);
xor U38570 (N_38570,N_38379,N_38037);
nor U38571 (N_38571,N_38028,N_38478);
and U38572 (N_38572,N_38016,N_38280);
nand U38573 (N_38573,N_38092,N_38325);
or U38574 (N_38574,N_38117,N_38471);
or U38575 (N_38575,N_38305,N_38433);
and U38576 (N_38576,N_38316,N_38422);
and U38577 (N_38577,N_38126,N_38406);
or U38578 (N_38578,N_38367,N_38195);
and U38579 (N_38579,N_38219,N_38044);
or U38580 (N_38580,N_38060,N_38023);
nor U38581 (N_38581,N_38137,N_38214);
nor U38582 (N_38582,N_38070,N_38254);
nor U38583 (N_38583,N_38479,N_38351);
or U38584 (N_38584,N_38335,N_38416);
or U38585 (N_38585,N_38245,N_38014);
and U38586 (N_38586,N_38116,N_38336);
nand U38587 (N_38587,N_38222,N_38298);
and U38588 (N_38588,N_38119,N_38125);
xor U38589 (N_38589,N_38149,N_38306);
nor U38590 (N_38590,N_38112,N_38344);
or U38591 (N_38591,N_38110,N_38083);
xor U38592 (N_38592,N_38468,N_38235);
and U38593 (N_38593,N_38413,N_38000);
nor U38594 (N_38594,N_38211,N_38181);
and U38595 (N_38595,N_38176,N_38436);
or U38596 (N_38596,N_38320,N_38020);
xor U38597 (N_38597,N_38189,N_38190);
or U38598 (N_38598,N_38292,N_38442);
nand U38599 (N_38599,N_38401,N_38476);
and U38600 (N_38600,N_38093,N_38236);
xor U38601 (N_38601,N_38488,N_38455);
nand U38602 (N_38602,N_38084,N_38317);
or U38603 (N_38603,N_38164,N_38111);
nand U38604 (N_38604,N_38012,N_38165);
nand U38605 (N_38605,N_38262,N_38266);
nand U38606 (N_38606,N_38201,N_38410);
and U38607 (N_38607,N_38069,N_38204);
or U38608 (N_38608,N_38099,N_38173);
and U38609 (N_38609,N_38243,N_38077);
or U38610 (N_38610,N_38293,N_38066);
nand U38611 (N_38611,N_38338,N_38131);
and U38612 (N_38612,N_38425,N_38319);
nor U38613 (N_38613,N_38133,N_38363);
or U38614 (N_38614,N_38400,N_38050);
nand U38615 (N_38615,N_38019,N_38203);
nand U38616 (N_38616,N_38237,N_38018);
xnor U38617 (N_38617,N_38147,N_38271);
nand U38618 (N_38618,N_38397,N_38261);
and U38619 (N_38619,N_38049,N_38396);
or U38620 (N_38620,N_38275,N_38043);
nor U38621 (N_38621,N_38441,N_38274);
xnor U38622 (N_38622,N_38289,N_38146);
or U38623 (N_38623,N_38134,N_38369);
and U38624 (N_38624,N_38056,N_38091);
and U38625 (N_38625,N_38227,N_38033);
or U38626 (N_38626,N_38208,N_38370);
nand U38627 (N_38627,N_38224,N_38324);
nand U38628 (N_38628,N_38463,N_38343);
and U38629 (N_38629,N_38326,N_38145);
or U38630 (N_38630,N_38076,N_38086);
and U38631 (N_38631,N_38472,N_38297);
nand U38632 (N_38632,N_38072,N_38158);
xnor U38633 (N_38633,N_38427,N_38094);
or U38634 (N_38634,N_38081,N_38402);
or U38635 (N_38635,N_38029,N_38008);
xnor U38636 (N_38636,N_38193,N_38225);
xor U38637 (N_38637,N_38328,N_38118);
and U38638 (N_38638,N_38394,N_38484);
nand U38639 (N_38639,N_38499,N_38285);
nor U38640 (N_38640,N_38323,N_38063);
nor U38641 (N_38641,N_38213,N_38264);
or U38642 (N_38642,N_38183,N_38223);
nand U38643 (N_38643,N_38333,N_38154);
nor U38644 (N_38644,N_38210,N_38088);
xor U38645 (N_38645,N_38418,N_38122);
or U38646 (N_38646,N_38374,N_38378);
nor U38647 (N_38647,N_38327,N_38085);
nor U38648 (N_38648,N_38209,N_38337);
nor U38649 (N_38649,N_38434,N_38206);
nand U38650 (N_38650,N_38453,N_38426);
nand U38651 (N_38651,N_38121,N_38184);
and U38652 (N_38652,N_38389,N_38113);
nand U38653 (N_38653,N_38494,N_38221);
nand U38654 (N_38654,N_38392,N_38260);
nor U38655 (N_38655,N_38309,N_38334);
and U38656 (N_38656,N_38365,N_38256);
and U38657 (N_38657,N_38097,N_38010);
nor U38658 (N_38658,N_38270,N_38062);
nor U38659 (N_38659,N_38267,N_38032);
or U38660 (N_38660,N_38159,N_38375);
and U38661 (N_38661,N_38002,N_38163);
nor U38662 (N_38662,N_38359,N_38246);
nand U38663 (N_38663,N_38331,N_38160);
nand U38664 (N_38664,N_38420,N_38007);
nor U38665 (N_38665,N_38482,N_38272);
nand U38666 (N_38666,N_38437,N_38409);
and U38667 (N_38667,N_38415,N_38360);
nand U38668 (N_38668,N_38361,N_38498);
nand U38669 (N_38669,N_38313,N_38178);
nand U38670 (N_38670,N_38250,N_38170);
and U38671 (N_38671,N_38251,N_38444);
nor U38672 (N_38672,N_38253,N_38232);
nand U38673 (N_38673,N_38357,N_38188);
nor U38674 (N_38674,N_38138,N_38136);
nand U38675 (N_38675,N_38090,N_38291);
and U38676 (N_38676,N_38315,N_38383);
nand U38677 (N_38677,N_38242,N_38286);
nand U38678 (N_38678,N_38405,N_38398);
and U38679 (N_38679,N_38330,N_38109);
and U38680 (N_38680,N_38186,N_38486);
or U38681 (N_38681,N_38342,N_38011);
and U38682 (N_38682,N_38407,N_38039);
and U38683 (N_38683,N_38130,N_38030);
and U38684 (N_38684,N_38481,N_38384);
nand U38685 (N_38685,N_38175,N_38106);
nand U38686 (N_38686,N_38456,N_38279);
and U38687 (N_38687,N_38027,N_38244);
or U38688 (N_38688,N_38248,N_38058);
xnor U38689 (N_38689,N_38258,N_38052);
nand U38690 (N_38690,N_38104,N_38207);
and U38691 (N_38691,N_38150,N_38493);
nor U38692 (N_38692,N_38089,N_38414);
and U38693 (N_38693,N_38151,N_38074);
nand U38694 (N_38694,N_38362,N_38464);
nor U38695 (N_38695,N_38031,N_38421);
and U38696 (N_38696,N_38100,N_38123);
and U38697 (N_38697,N_38430,N_38017);
nor U38698 (N_38698,N_38459,N_38295);
nand U38699 (N_38699,N_38182,N_38107);
or U38700 (N_38700,N_38241,N_38448);
nor U38701 (N_38701,N_38047,N_38347);
xnor U38702 (N_38702,N_38473,N_38021);
or U38703 (N_38703,N_38001,N_38386);
or U38704 (N_38704,N_38162,N_38226);
or U38705 (N_38705,N_38143,N_38301);
or U38706 (N_38706,N_38399,N_38477);
nand U38707 (N_38707,N_38388,N_38067);
nand U38708 (N_38708,N_38391,N_38102);
xnor U38709 (N_38709,N_38013,N_38087);
xnor U38710 (N_38710,N_38322,N_38156);
nor U38711 (N_38711,N_38155,N_38061);
and U38712 (N_38712,N_38035,N_38364);
nor U38713 (N_38713,N_38423,N_38101);
nand U38714 (N_38714,N_38307,N_38497);
or U38715 (N_38715,N_38296,N_38259);
nor U38716 (N_38716,N_38148,N_38129);
nor U38717 (N_38717,N_38288,N_38310);
or U38718 (N_38718,N_38480,N_38265);
or U38719 (N_38719,N_38166,N_38191);
and U38720 (N_38720,N_38273,N_38053);
nand U38721 (N_38721,N_38294,N_38412);
nand U38722 (N_38722,N_38411,N_38071);
nor U38723 (N_38723,N_38144,N_38312);
or U38724 (N_38724,N_38467,N_38469);
and U38725 (N_38725,N_38240,N_38385);
and U38726 (N_38726,N_38287,N_38340);
nand U38727 (N_38727,N_38200,N_38095);
and U38728 (N_38728,N_38454,N_38462);
and U38729 (N_38729,N_38142,N_38197);
nand U38730 (N_38730,N_38457,N_38276);
nand U38731 (N_38731,N_38470,N_38042);
or U38732 (N_38732,N_38022,N_38003);
or U38733 (N_38733,N_38268,N_38290);
nor U38734 (N_38734,N_38403,N_38446);
and U38735 (N_38735,N_38304,N_38217);
and U38736 (N_38736,N_38141,N_38115);
or U38737 (N_38737,N_38263,N_38419);
nor U38738 (N_38738,N_38339,N_38139);
nand U38739 (N_38739,N_38152,N_38341);
or U38740 (N_38740,N_38447,N_38026);
and U38741 (N_38741,N_38308,N_38475);
and U38742 (N_38742,N_38199,N_38387);
and U38743 (N_38743,N_38435,N_38098);
or U38744 (N_38744,N_38171,N_38231);
nor U38745 (N_38745,N_38073,N_38283);
nor U38746 (N_38746,N_38048,N_38353);
nand U38747 (N_38747,N_38127,N_38381);
or U38748 (N_38748,N_38157,N_38168);
nand U38749 (N_38749,N_38487,N_38395);
or U38750 (N_38750,N_38439,N_38094);
or U38751 (N_38751,N_38466,N_38183);
and U38752 (N_38752,N_38233,N_38022);
and U38753 (N_38753,N_38258,N_38114);
and U38754 (N_38754,N_38092,N_38403);
nor U38755 (N_38755,N_38204,N_38182);
and U38756 (N_38756,N_38462,N_38181);
or U38757 (N_38757,N_38156,N_38416);
and U38758 (N_38758,N_38441,N_38061);
and U38759 (N_38759,N_38215,N_38132);
nor U38760 (N_38760,N_38018,N_38354);
nor U38761 (N_38761,N_38155,N_38076);
and U38762 (N_38762,N_38242,N_38413);
nand U38763 (N_38763,N_38056,N_38131);
nand U38764 (N_38764,N_38420,N_38463);
nand U38765 (N_38765,N_38393,N_38251);
or U38766 (N_38766,N_38117,N_38028);
nand U38767 (N_38767,N_38004,N_38407);
or U38768 (N_38768,N_38204,N_38011);
xor U38769 (N_38769,N_38074,N_38103);
or U38770 (N_38770,N_38334,N_38322);
nand U38771 (N_38771,N_38098,N_38450);
nand U38772 (N_38772,N_38375,N_38289);
nand U38773 (N_38773,N_38343,N_38271);
or U38774 (N_38774,N_38088,N_38461);
nor U38775 (N_38775,N_38329,N_38178);
nor U38776 (N_38776,N_38165,N_38400);
nand U38777 (N_38777,N_38165,N_38249);
or U38778 (N_38778,N_38204,N_38032);
xor U38779 (N_38779,N_38238,N_38008);
and U38780 (N_38780,N_38394,N_38028);
or U38781 (N_38781,N_38316,N_38342);
xor U38782 (N_38782,N_38089,N_38083);
and U38783 (N_38783,N_38439,N_38150);
and U38784 (N_38784,N_38307,N_38033);
nor U38785 (N_38785,N_38349,N_38472);
or U38786 (N_38786,N_38290,N_38018);
nor U38787 (N_38787,N_38208,N_38122);
nand U38788 (N_38788,N_38488,N_38154);
or U38789 (N_38789,N_38137,N_38106);
nor U38790 (N_38790,N_38180,N_38404);
and U38791 (N_38791,N_38308,N_38111);
or U38792 (N_38792,N_38106,N_38231);
nor U38793 (N_38793,N_38238,N_38240);
nand U38794 (N_38794,N_38425,N_38302);
nor U38795 (N_38795,N_38484,N_38055);
nor U38796 (N_38796,N_38261,N_38463);
and U38797 (N_38797,N_38354,N_38171);
nor U38798 (N_38798,N_38292,N_38144);
nand U38799 (N_38799,N_38434,N_38409);
nor U38800 (N_38800,N_38484,N_38422);
xor U38801 (N_38801,N_38330,N_38292);
xnor U38802 (N_38802,N_38436,N_38388);
nand U38803 (N_38803,N_38405,N_38157);
nor U38804 (N_38804,N_38292,N_38074);
or U38805 (N_38805,N_38161,N_38007);
nor U38806 (N_38806,N_38187,N_38048);
nand U38807 (N_38807,N_38411,N_38177);
nor U38808 (N_38808,N_38330,N_38088);
nor U38809 (N_38809,N_38278,N_38490);
nor U38810 (N_38810,N_38245,N_38395);
or U38811 (N_38811,N_38117,N_38201);
xnor U38812 (N_38812,N_38130,N_38315);
and U38813 (N_38813,N_38448,N_38088);
and U38814 (N_38814,N_38194,N_38413);
nor U38815 (N_38815,N_38499,N_38491);
nand U38816 (N_38816,N_38099,N_38391);
nand U38817 (N_38817,N_38268,N_38111);
nand U38818 (N_38818,N_38463,N_38168);
nand U38819 (N_38819,N_38461,N_38154);
and U38820 (N_38820,N_38275,N_38337);
or U38821 (N_38821,N_38336,N_38408);
or U38822 (N_38822,N_38314,N_38013);
nand U38823 (N_38823,N_38046,N_38262);
nor U38824 (N_38824,N_38179,N_38489);
xnor U38825 (N_38825,N_38362,N_38434);
nand U38826 (N_38826,N_38350,N_38065);
or U38827 (N_38827,N_38473,N_38066);
nor U38828 (N_38828,N_38439,N_38160);
nand U38829 (N_38829,N_38232,N_38441);
nor U38830 (N_38830,N_38227,N_38236);
or U38831 (N_38831,N_38163,N_38116);
nand U38832 (N_38832,N_38069,N_38347);
and U38833 (N_38833,N_38060,N_38257);
xnor U38834 (N_38834,N_38338,N_38466);
and U38835 (N_38835,N_38026,N_38262);
and U38836 (N_38836,N_38452,N_38461);
or U38837 (N_38837,N_38131,N_38416);
and U38838 (N_38838,N_38198,N_38062);
nand U38839 (N_38839,N_38024,N_38414);
and U38840 (N_38840,N_38441,N_38081);
nor U38841 (N_38841,N_38499,N_38462);
xnor U38842 (N_38842,N_38271,N_38228);
or U38843 (N_38843,N_38233,N_38413);
and U38844 (N_38844,N_38336,N_38158);
xor U38845 (N_38845,N_38445,N_38008);
and U38846 (N_38846,N_38193,N_38263);
nand U38847 (N_38847,N_38073,N_38490);
or U38848 (N_38848,N_38311,N_38260);
nand U38849 (N_38849,N_38137,N_38162);
nor U38850 (N_38850,N_38281,N_38405);
and U38851 (N_38851,N_38131,N_38058);
nor U38852 (N_38852,N_38044,N_38102);
nor U38853 (N_38853,N_38447,N_38332);
nor U38854 (N_38854,N_38197,N_38387);
or U38855 (N_38855,N_38204,N_38302);
or U38856 (N_38856,N_38219,N_38259);
nor U38857 (N_38857,N_38356,N_38304);
xnor U38858 (N_38858,N_38072,N_38375);
nor U38859 (N_38859,N_38142,N_38336);
nand U38860 (N_38860,N_38366,N_38290);
nor U38861 (N_38861,N_38420,N_38391);
or U38862 (N_38862,N_38078,N_38425);
nor U38863 (N_38863,N_38023,N_38218);
or U38864 (N_38864,N_38080,N_38438);
nor U38865 (N_38865,N_38255,N_38443);
xnor U38866 (N_38866,N_38195,N_38359);
or U38867 (N_38867,N_38467,N_38241);
nand U38868 (N_38868,N_38092,N_38123);
nor U38869 (N_38869,N_38361,N_38006);
nand U38870 (N_38870,N_38146,N_38138);
and U38871 (N_38871,N_38245,N_38027);
and U38872 (N_38872,N_38351,N_38348);
or U38873 (N_38873,N_38242,N_38388);
and U38874 (N_38874,N_38281,N_38179);
or U38875 (N_38875,N_38067,N_38273);
xor U38876 (N_38876,N_38063,N_38262);
or U38877 (N_38877,N_38427,N_38471);
and U38878 (N_38878,N_38196,N_38407);
nor U38879 (N_38879,N_38247,N_38258);
or U38880 (N_38880,N_38248,N_38052);
nand U38881 (N_38881,N_38450,N_38178);
nor U38882 (N_38882,N_38329,N_38354);
and U38883 (N_38883,N_38404,N_38249);
or U38884 (N_38884,N_38158,N_38439);
and U38885 (N_38885,N_38075,N_38150);
nand U38886 (N_38886,N_38174,N_38230);
and U38887 (N_38887,N_38142,N_38411);
nand U38888 (N_38888,N_38413,N_38145);
and U38889 (N_38889,N_38025,N_38031);
nor U38890 (N_38890,N_38330,N_38137);
and U38891 (N_38891,N_38303,N_38074);
nor U38892 (N_38892,N_38408,N_38209);
nor U38893 (N_38893,N_38110,N_38337);
nor U38894 (N_38894,N_38292,N_38343);
nand U38895 (N_38895,N_38463,N_38331);
or U38896 (N_38896,N_38328,N_38161);
nand U38897 (N_38897,N_38356,N_38278);
nor U38898 (N_38898,N_38387,N_38431);
xor U38899 (N_38899,N_38087,N_38393);
and U38900 (N_38900,N_38332,N_38001);
or U38901 (N_38901,N_38488,N_38019);
and U38902 (N_38902,N_38272,N_38144);
nand U38903 (N_38903,N_38108,N_38063);
nand U38904 (N_38904,N_38205,N_38252);
and U38905 (N_38905,N_38465,N_38407);
xnor U38906 (N_38906,N_38283,N_38261);
and U38907 (N_38907,N_38336,N_38169);
and U38908 (N_38908,N_38019,N_38080);
nand U38909 (N_38909,N_38210,N_38118);
and U38910 (N_38910,N_38084,N_38278);
or U38911 (N_38911,N_38498,N_38364);
nor U38912 (N_38912,N_38117,N_38156);
or U38913 (N_38913,N_38320,N_38155);
xnor U38914 (N_38914,N_38482,N_38210);
xnor U38915 (N_38915,N_38253,N_38408);
or U38916 (N_38916,N_38365,N_38009);
xnor U38917 (N_38917,N_38340,N_38166);
nand U38918 (N_38918,N_38243,N_38410);
nand U38919 (N_38919,N_38163,N_38028);
or U38920 (N_38920,N_38437,N_38126);
nor U38921 (N_38921,N_38447,N_38194);
or U38922 (N_38922,N_38125,N_38472);
nand U38923 (N_38923,N_38017,N_38377);
or U38924 (N_38924,N_38310,N_38080);
and U38925 (N_38925,N_38190,N_38324);
nor U38926 (N_38926,N_38142,N_38398);
or U38927 (N_38927,N_38354,N_38312);
nor U38928 (N_38928,N_38205,N_38055);
and U38929 (N_38929,N_38057,N_38187);
nand U38930 (N_38930,N_38188,N_38232);
or U38931 (N_38931,N_38245,N_38347);
or U38932 (N_38932,N_38384,N_38447);
nor U38933 (N_38933,N_38460,N_38115);
and U38934 (N_38934,N_38038,N_38098);
and U38935 (N_38935,N_38077,N_38353);
nor U38936 (N_38936,N_38220,N_38369);
nand U38937 (N_38937,N_38149,N_38157);
nor U38938 (N_38938,N_38375,N_38139);
xnor U38939 (N_38939,N_38140,N_38082);
nand U38940 (N_38940,N_38205,N_38105);
or U38941 (N_38941,N_38217,N_38319);
or U38942 (N_38942,N_38378,N_38000);
nand U38943 (N_38943,N_38209,N_38109);
or U38944 (N_38944,N_38089,N_38292);
and U38945 (N_38945,N_38034,N_38182);
xor U38946 (N_38946,N_38234,N_38286);
nand U38947 (N_38947,N_38401,N_38038);
or U38948 (N_38948,N_38016,N_38452);
and U38949 (N_38949,N_38350,N_38073);
nand U38950 (N_38950,N_38069,N_38363);
nor U38951 (N_38951,N_38246,N_38238);
nor U38952 (N_38952,N_38156,N_38292);
and U38953 (N_38953,N_38018,N_38478);
and U38954 (N_38954,N_38069,N_38271);
and U38955 (N_38955,N_38069,N_38093);
nand U38956 (N_38956,N_38363,N_38352);
nand U38957 (N_38957,N_38006,N_38160);
nand U38958 (N_38958,N_38267,N_38049);
xor U38959 (N_38959,N_38216,N_38210);
xor U38960 (N_38960,N_38067,N_38226);
or U38961 (N_38961,N_38374,N_38270);
and U38962 (N_38962,N_38255,N_38220);
and U38963 (N_38963,N_38304,N_38023);
and U38964 (N_38964,N_38293,N_38313);
or U38965 (N_38965,N_38334,N_38068);
or U38966 (N_38966,N_38475,N_38117);
nand U38967 (N_38967,N_38058,N_38092);
nor U38968 (N_38968,N_38496,N_38380);
nor U38969 (N_38969,N_38182,N_38014);
nor U38970 (N_38970,N_38246,N_38194);
and U38971 (N_38971,N_38168,N_38061);
nor U38972 (N_38972,N_38153,N_38365);
and U38973 (N_38973,N_38070,N_38257);
nand U38974 (N_38974,N_38134,N_38060);
and U38975 (N_38975,N_38095,N_38174);
nor U38976 (N_38976,N_38095,N_38230);
xnor U38977 (N_38977,N_38215,N_38352);
and U38978 (N_38978,N_38415,N_38469);
nor U38979 (N_38979,N_38421,N_38111);
nor U38980 (N_38980,N_38053,N_38361);
nor U38981 (N_38981,N_38269,N_38439);
and U38982 (N_38982,N_38166,N_38000);
nand U38983 (N_38983,N_38094,N_38362);
xnor U38984 (N_38984,N_38417,N_38447);
and U38985 (N_38985,N_38366,N_38338);
and U38986 (N_38986,N_38474,N_38335);
nor U38987 (N_38987,N_38259,N_38025);
nand U38988 (N_38988,N_38015,N_38056);
or U38989 (N_38989,N_38461,N_38176);
or U38990 (N_38990,N_38074,N_38483);
or U38991 (N_38991,N_38132,N_38050);
nor U38992 (N_38992,N_38178,N_38078);
nand U38993 (N_38993,N_38198,N_38291);
or U38994 (N_38994,N_38054,N_38037);
xnor U38995 (N_38995,N_38221,N_38312);
or U38996 (N_38996,N_38433,N_38233);
nand U38997 (N_38997,N_38352,N_38470);
nand U38998 (N_38998,N_38398,N_38325);
xor U38999 (N_38999,N_38438,N_38492);
nand U39000 (N_39000,N_38698,N_38800);
nor U39001 (N_39001,N_38908,N_38557);
nor U39002 (N_39002,N_38885,N_38627);
nand U39003 (N_39003,N_38608,N_38537);
and U39004 (N_39004,N_38682,N_38662);
xor U39005 (N_39005,N_38701,N_38536);
nor U39006 (N_39006,N_38630,N_38962);
and U39007 (N_39007,N_38747,N_38754);
nor U39008 (N_39008,N_38953,N_38526);
xnor U39009 (N_39009,N_38591,N_38650);
nor U39010 (N_39010,N_38805,N_38809);
and U39011 (N_39011,N_38581,N_38862);
and U39012 (N_39012,N_38788,N_38714);
nor U39013 (N_39013,N_38795,N_38705);
or U39014 (N_39014,N_38769,N_38540);
or U39015 (N_39015,N_38741,N_38589);
and U39016 (N_39016,N_38811,N_38645);
or U39017 (N_39017,N_38657,N_38851);
and U39018 (N_39018,N_38571,N_38525);
nor U39019 (N_39019,N_38959,N_38804);
and U39020 (N_39020,N_38562,N_38738);
nand U39021 (N_39021,N_38577,N_38995);
xnor U39022 (N_39022,N_38950,N_38726);
nand U39023 (N_39023,N_38825,N_38952);
and U39024 (N_39024,N_38944,N_38846);
xnor U39025 (N_39025,N_38934,N_38822);
nand U39026 (N_39026,N_38896,N_38632);
and U39027 (N_39027,N_38585,N_38672);
and U39028 (N_39028,N_38764,N_38559);
or U39029 (N_39029,N_38860,N_38920);
and U39030 (N_39030,N_38816,N_38633);
nor U39031 (N_39031,N_38879,N_38979);
nand U39032 (N_39032,N_38622,N_38919);
and U39033 (N_39033,N_38721,N_38617);
nor U39034 (N_39034,N_38936,N_38693);
or U39035 (N_39035,N_38579,N_38775);
and U39036 (N_39036,N_38539,N_38659);
nor U39037 (N_39037,N_38960,N_38977);
nor U39038 (N_39038,N_38907,N_38667);
nand U39039 (N_39039,N_38821,N_38828);
nand U39040 (N_39040,N_38678,N_38763);
and U39041 (N_39041,N_38778,N_38558);
nor U39042 (N_39042,N_38786,N_38875);
nor U39043 (N_39043,N_38947,N_38859);
nand U39044 (N_39044,N_38887,N_38724);
and U39045 (N_39045,N_38757,N_38722);
and U39046 (N_39046,N_38535,N_38787);
nand U39047 (N_39047,N_38899,N_38845);
xor U39048 (N_39048,N_38553,N_38538);
nand U39049 (N_39049,N_38695,N_38694);
or U39050 (N_39050,N_38915,N_38855);
xor U39051 (N_39051,N_38761,N_38576);
and U39052 (N_39052,N_38731,N_38543);
nor U39053 (N_39053,N_38864,N_38756);
or U39054 (N_39054,N_38813,N_38911);
and U39055 (N_39055,N_38565,N_38753);
nor U39056 (N_39056,N_38856,N_38969);
nor U39057 (N_39057,N_38938,N_38502);
or U39058 (N_39058,N_38767,N_38729);
or U39059 (N_39059,N_38623,N_38643);
xor U39060 (N_39060,N_38651,N_38642);
and U39061 (N_39061,N_38710,N_38897);
nor U39062 (N_39062,N_38863,N_38857);
nor U39063 (N_39063,N_38532,N_38886);
and U39064 (N_39064,N_38586,N_38774);
or U39065 (N_39065,N_38981,N_38734);
nand U39066 (N_39066,N_38574,N_38575);
or U39067 (N_39067,N_38626,N_38777);
nor U39068 (N_39068,N_38758,N_38797);
or U39069 (N_39069,N_38573,N_38604);
or U39070 (N_39070,N_38928,N_38620);
xnor U39071 (N_39071,N_38964,N_38906);
or U39072 (N_39072,N_38718,N_38904);
or U39073 (N_39073,N_38689,N_38831);
nor U39074 (N_39074,N_38900,N_38834);
or U39075 (N_39075,N_38635,N_38599);
and U39076 (N_39076,N_38658,N_38618);
nand U39077 (N_39077,N_38654,N_38823);
or U39078 (N_39078,N_38880,N_38973);
nand U39079 (N_39079,N_38739,N_38641);
or U39080 (N_39080,N_38621,N_38740);
nand U39081 (N_39081,N_38556,N_38554);
nand U39082 (N_39082,N_38592,N_38649);
nand U39083 (N_39083,N_38607,N_38692);
nand U39084 (N_39084,N_38771,N_38597);
nor U39085 (N_39085,N_38884,N_38807);
nand U39086 (N_39086,N_38600,N_38636);
or U39087 (N_39087,N_38660,N_38712);
xnor U39088 (N_39088,N_38541,N_38515);
or U39089 (N_39089,N_38700,N_38681);
nor U39090 (N_39090,N_38531,N_38970);
xnor U39091 (N_39091,N_38798,N_38792);
nand U39092 (N_39092,N_38588,N_38951);
nand U39093 (N_39093,N_38910,N_38527);
nor U39094 (N_39094,N_38683,N_38655);
nor U39095 (N_39095,N_38796,N_38877);
nand U39096 (N_39096,N_38881,N_38967);
xnor U39097 (N_39097,N_38567,N_38566);
nor U39098 (N_39098,N_38595,N_38814);
or U39099 (N_39099,N_38521,N_38609);
or U39100 (N_39100,N_38716,N_38986);
nor U39101 (N_39101,N_38582,N_38522);
or U39102 (N_39102,N_38760,N_38918);
nand U39103 (N_39103,N_38820,N_38590);
or U39104 (N_39104,N_38612,N_38839);
or U39105 (N_39105,N_38686,N_38883);
nor U39106 (N_39106,N_38916,N_38765);
nand U39107 (N_39107,N_38614,N_38790);
and U39108 (N_39108,N_38932,N_38512);
nand U39109 (N_39109,N_38530,N_38974);
nand U39110 (N_39110,N_38817,N_38941);
and U39111 (N_39111,N_38991,N_38561);
or U39112 (N_39112,N_38687,N_38545);
and U39113 (N_39113,N_38968,N_38815);
xor U39114 (N_39114,N_38544,N_38909);
and U39115 (N_39115,N_38746,N_38664);
and U39116 (N_39116,N_38519,N_38983);
nand U39117 (N_39117,N_38997,N_38848);
and U39118 (N_39118,N_38528,N_38925);
nor U39119 (N_39119,N_38546,N_38755);
nand U39120 (N_39120,N_38893,N_38615);
nand U39121 (N_39121,N_38870,N_38598);
nor U39122 (N_39122,N_38963,N_38781);
or U39123 (N_39123,N_38929,N_38580);
and U39124 (N_39124,N_38549,N_38830);
nand U39125 (N_39125,N_38652,N_38542);
and U39126 (N_39126,N_38513,N_38719);
nand U39127 (N_39127,N_38674,N_38924);
nand U39128 (N_39128,N_38836,N_38616);
nor U39129 (N_39129,N_38569,N_38534);
nor U39130 (N_39130,N_38751,N_38661);
xnor U39131 (N_39131,N_38782,N_38587);
or U39132 (N_39132,N_38677,N_38989);
nand U39133 (N_39133,N_38946,N_38610);
or U39134 (N_39134,N_38961,N_38762);
xor U39135 (N_39135,N_38637,N_38551);
nand U39136 (N_39136,N_38844,N_38752);
and U39137 (N_39137,N_38560,N_38759);
nand U39138 (N_39138,N_38978,N_38696);
or U39139 (N_39139,N_38669,N_38665);
or U39140 (N_39140,N_38921,N_38980);
nand U39141 (N_39141,N_38913,N_38745);
xor U39142 (N_39142,N_38548,N_38985);
or U39143 (N_39143,N_38776,N_38976);
or U39144 (N_39144,N_38824,N_38748);
and U39145 (N_39145,N_38998,N_38902);
nand U39146 (N_39146,N_38602,N_38835);
and U39147 (N_39147,N_38939,N_38987);
and U39148 (N_39148,N_38930,N_38994);
xnor U39149 (N_39149,N_38866,N_38671);
and U39150 (N_39150,N_38605,N_38517);
xnor U39151 (N_39151,N_38680,N_38601);
xnor U39152 (N_39152,N_38647,N_38653);
nor U39153 (N_39153,N_38518,N_38720);
nor U39154 (N_39154,N_38699,N_38849);
xnor U39155 (N_39155,N_38572,N_38793);
nand U39156 (N_39156,N_38940,N_38794);
and U39157 (N_39157,N_38727,N_38503);
and U39158 (N_39158,N_38768,N_38744);
nand U39159 (N_39159,N_38933,N_38841);
and U39160 (N_39160,N_38993,N_38914);
or U39161 (N_39161,N_38890,N_38583);
nor U39162 (N_39162,N_38871,N_38770);
and U39163 (N_39163,N_38837,N_38827);
or U39164 (N_39164,N_38780,N_38552);
and U39165 (N_39165,N_38766,N_38949);
and U39166 (N_39166,N_38818,N_38711);
or U39167 (N_39167,N_38802,N_38533);
xnor U39168 (N_39168,N_38903,N_38840);
or U39169 (N_39169,N_38688,N_38555);
nand U39170 (N_39170,N_38510,N_38882);
and U39171 (N_39171,N_38666,N_38500);
and U39172 (N_39172,N_38889,N_38843);
xnor U39173 (N_39173,N_38584,N_38594);
and U39174 (N_39174,N_38975,N_38892);
nor U39175 (N_39175,N_38613,N_38656);
nand U39176 (N_39176,N_38803,N_38808);
nor U39177 (N_39177,N_38966,N_38878);
xor U39178 (N_39178,N_38873,N_38861);
and U39179 (N_39179,N_38958,N_38676);
nand U39180 (N_39180,N_38965,N_38888);
or U39181 (N_39181,N_38988,N_38876);
or U39182 (N_39182,N_38663,N_38631);
nand U39183 (N_39183,N_38628,N_38838);
xor U39184 (N_39184,N_38749,N_38514);
and U39185 (N_39185,N_38593,N_38772);
nor U39186 (N_39186,N_38506,N_38673);
or U39187 (N_39187,N_38955,N_38791);
and U39188 (N_39188,N_38894,N_38806);
and U39189 (N_39189,N_38625,N_38773);
xor U39190 (N_39190,N_38564,N_38634);
and U39191 (N_39191,N_38723,N_38927);
nor U39192 (N_39192,N_38853,N_38709);
or U39193 (N_39193,N_38685,N_38922);
and U39194 (N_39194,N_38736,N_38708);
nor U39195 (N_39195,N_38697,N_38784);
and U39196 (N_39196,N_38703,N_38619);
nor U39197 (N_39197,N_38799,N_38702);
xnor U39198 (N_39198,N_38743,N_38812);
nor U39199 (N_39199,N_38905,N_38629);
or U39200 (N_39200,N_38606,N_38735);
or U39201 (N_39201,N_38639,N_38730);
xor U39202 (N_39202,N_38520,N_38529);
xnor U39203 (N_39203,N_38996,N_38874);
or U39204 (N_39204,N_38507,N_38644);
and U39205 (N_39205,N_38640,N_38842);
and U39206 (N_39206,N_38789,N_38670);
or U39207 (N_39207,N_38847,N_38937);
and U39208 (N_39208,N_38713,N_38819);
or U39209 (N_39209,N_38972,N_38717);
xnor U39210 (N_39210,N_38728,N_38706);
nor U39211 (N_39211,N_38898,N_38523);
or U39212 (N_39212,N_38971,N_38783);
xnor U39213 (N_39213,N_38511,N_38984);
and U39214 (N_39214,N_38854,N_38917);
nor U39215 (N_39215,N_38829,N_38948);
or U39216 (N_39216,N_38691,N_38690);
or U39217 (N_39217,N_38750,N_38779);
nand U39218 (N_39218,N_38675,N_38869);
or U39219 (N_39219,N_38923,N_38872);
xor U39220 (N_39220,N_38684,N_38679);
xnor U39221 (N_39221,N_38570,N_38935);
or U39222 (N_39222,N_38508,N_38603);
nand U39223 (N_39223,N_38668,N_38926);
or U39224 (N_39224,N_38638,N_38785);
nor U39225 (N_39225,N_38868,N_38715);
nor U39226 (N_39226,N_38982,N_38833);
or U39227 (N_39227,N_38563,N_38596);
or U39228 (N_39228,N_38826,N_38624);
nand U39229 (N_39229,N_38867,N_38707);
or U39230 (N_39230,N_38578,N_38505);
nand U39231 (N_39231,N_38852,N_38992);
nor U39232 (N_39232,N_38954,N_38901);
nor U39233 (N_39233,N_38832,N_38858);
and U39234 (N_39234,N_38568,N_38865);
xnor U39235 (N_39235,N_38547,N_38524);
or U39236 (N_39236,N_38931,N_38732);
nor U39237 (N_39237,N_38891,N_38516);
or U39238 (N_39238,N_38550,N_38810);
nand U39239 (N_39239,N_38611,N_38725);
nor U39240 (N_39240,N_38742,N_38895);
nand U39241 (N_39241,N_38504,N_38850);
and U39242 (N_39242,N_38646,N_38945);
xor U39243 (N_39243,N_38943,N_38801);
nand U39244 (N_39244,N_38956,N_38999);
or U39245 (N_39245,N_38648,N_38942);
xor U39246 (N_39246,N_38509,N_38733);
nand U39247 (N_39247,N_38957,N_38704);
nand U39248 (N_39248,N_38501,N_38912);
nor U39249 (N_39249,N_38990,N_38737);
nand U39250 (N_39250,N_38685,N_38961);
and U39251 (N_39251,N_38935,N_38910);
xor U39252 (N_39252,N_38613,N_38622);
nand U39253 (N_39253,N_38717,N_38964);
and U39254 (N_39254,N_38634,N_38963);
nor U39255 (N_39255,N_38515,N_38596);
or U39256 (N_39256,N_38808,N_38880);
nor U39257 (N_39257,N_38732,N_38733);
nand U39258 (N_39258,N_38891,N_38873);
and U39259 (N_39259,N_38737,N_38742);
nand U39260 (N_39260,N_38971,N_38758);
and U39261 (N_39261,N_38736,N_38641);
nor U39262 (N_39262,N_38771,N_38940);
nor U39263 (N_39263,N_38540,N_38923);
nor U39264 (N_39264,N_38521,N_38660);
nand U39265 (N_39265,N_38500,N_38592);
or U39266 (N_39266,N_38581,N_38768);
xor U39267 (N_39267,N_38848,N_38587);
or U39268 (N_39268,N_38895,N_38775);
and U39269 (N_39269,N_38559,N_38670);
nand U39270 (N_39270,N_38553,N_38697);
nor U39271 (N_39271,N_38831,N_38995);
nor U39272 (N_39272,N_38808,N_38568);
or U39273 (N_39273,N_38741,N_38922);
nor U39274 (N_39274,N_38714,N_38673);
nor U39275 (N_39275,N_38978,N_38798);
nor U39276 (N_39276,N_38519,N_38824);
nand U39277 (N_39277,N_38698,N_38504);
and U39278 (N_39278,N_38612,N_38698);
or U39279 (N_39279,N_38593,N_38975);
or U39280 (N_39280,N_38897,N_38707);
nor U39281 (N_39281,N_38874,N_38670);
or U39282 (N_39282,N_38854,N_38726);
or U39283 (N_39283,N_38594,N_38780);
and U39284 (N_39284,N_38814,N_38824);
nand U39285 (N_39285,N_38656,N_38605);
nor U39286 (N_39286,N_38693,N_38975);
xnor U39287 (N_39287,N_38828,N_38721);
nor U39288 (N_39288,N_38840,N_38727);
and U39289 (N_39289,N_38824,N_38605);
or U39290 (N_39290,N_38909,N_38722);
nor U39291 (N_39291,N_38815,N_38571);
and U39292 (N_39292,N_38751,N_38530);
and U39293 (N_39293,N_38611,N_38939);
or U39294 (N_39294,N_38844,N_38931);
nand U39295 (N_39295,N_38995,N_38723);
xnor U39296 (N_39296,N_38518,N_38622);
nor U39297 (N_39297,N_38942,N_38888);
or U39298 (N_39298,N_38752,N_38771);
nand U39299 (N_39299,N_38845,N_38551);
or U39300 (N_39300,N_38908,N_38539);
nor U39301 (N_39301,N_38954,N_38894);
or U39302 (N_39302,N_38660,N_38675);
nand U39303 (N_39303,N_38840,N_38531);
nor U39304 (N_39304,N_38774,N_38537);
and U39305 (N_39305,N_38770,N_38536);
nand U39306 (N_39306,N_38895,N_38735);
nand U39307 (N_39307,N_38870,N_38830);
and U39308 (N_39308,N_38928,N_38992);
nor U39309 (N_39309,N_38746,N_38514);
nand U39310 (N_39310,N_38864,N_38614);
nand U39311 (N_39311,N_38637,N_38504);
nor U39312 (N_39312,N_38658,N_38837);
nor U39313 (N_39313,N_38891,N_38657);
or U39314 (N_39314,N_38936,N_38504);
xnor U39315 (N_39315,N_38794,N_38587);
or U39316 (N_39316,N_38854,N_38737);
nor U39317 (N_39317,N_38613,N_38815);
and U39318 (N_39318,N_38584,N_38784);
nand U39319 (N_39319,N_38597,N_38681);
and U39320 (N_39320,N_38732,N_38935);
or U39321 (N_39321,N_38525,N_38555);
nor U39322 (N_39322,N_38886,N_38981);
and U39323 (N_39323,N_38552,N_38923);
and U39324 (N_39324,N_38530,N_38706);
xor U39325 (N_39325,N_38887,N_38734);
xnor U39326 (N_39326,N_38537,N_38540);
nand U39327 (N_39327,N_38992,N_38603);
nor U39328 (N_39328,N_38984,N_38914);
nand U39329 (N_39329,N_38933,N_38840);
or U39330 (N_39330,N_38757,N_38977);
and U39331 (N_39331,N_38545,N_38841);
or U39332 (N_39332,N_38697,N_38852);
and U39333 (N_39333,N_38943,N_38950);
and U39334 (N_39334,N_38700,N_38712);
xor U39335 (N_39335,N_38701,N_38887);
nand U39336 (N_39336,N_38663,N_38521);
and U39337 (N_39337,N_38771,N_38798);
nor U39338 (N_39338,N_38666,N_38515);
or U39339 (N_39339,N_38933,N_38665);
and U39340 (N_39340,N_38941,N_38888);
xnor U39341 (N_39341,N_38701,N_38915);
or U39342 (N_39342,N_38802,N_38978);
or U39343 (N_39343,N_38902,N_38865);
nand U39344 (N_39344,N_38670,N_38654);
nand U39345 (N_39345,N_38823,N_38825);
and U39346 (N_39346,N_38629,N_38809);
or U39347 (N_39347,N_38550,N_38700);
nor U39348 (N_39348,N_38873,N_38741);
and U39349 (N_39349,N_38887,N_38995);
nand U39350 (N_39350,N_38859,N_38791);
nor U39351 (N_39351,N_38671,N_38532);
nor U39352 (N_39352,N_38931,N_38707);
nand U39353 (N_39353,N_38805,N_38714);
and U39354 (N_39354,N_38763,N_38751);
or U39355 (N_39355,N_38979,N_38618);
nand U39356 (N_39356,N_38501,N_38544);
and U39357 (N_39357,N_38842,N_38622);
xnor U39358 (N_39358,N_38662,N_38775);
and U39359 (N_39359,N_38990,N_38811);
nor U39360 (N_39360,N_38535,N_38608);
nand U39361 (N_39361,N_38650,N_38592);
and U39362 (N_39362,N_38758,N_38563);
nor U39363 (N_39363,N_38878,N_38668);
nor U39364 (N_39364,N_38586,N_38678);
or U39365 (N_39365,N_38894,N_38843);
nand U39366 (N_39366,N_38967,N_38682);
or U39367 (N_39367,N_38682,N_38807);
or U39368 (N_39368,N_38941,N_38872);
nor U39369 (N_39369,N_38924,N_38549);
nor U39370 (N_39370,N_38862,N_38767);
or U39371 (N_39371,N_38693,N_38667);
xnor U39372 (N_39372,N_38851,N_38923);
nand U39373 (N_39373,N_38858,N_38804);
nand U39374 (N_39374,N_38961,N_38797);
or U39375 (N_39375,N_38615,N_38830);
nor U39376 (N_39376,N_38792,N_38636);
nand U39377 (N_39377,N_38543,N_38734);
and U39378 (N_39378,N_38691,N_38581);
or U39379 (N_39379,N_38730,N_38836);
nor U39380 (N_39380,N_38694,N_38657);
nor U39381 (N_39381,N_38572,N_38531);
nor U39382 (N_39382,N_38838,N_38627);
nand U39383 (N_39383,N_38677,N_38923);
nand U39384 (N_39384,N_38750,N_38959);
and U39385 (N_39385,N_38676,N_38749);
and U39386 (N_39386,N_38952,N_38841);
nand U39387 (N_39387,N_38961,N_38560);
or U39388 (N_39388,N_38792,N_38752);
or U39389 (N_39389,N_38736,N_38697);
or U39390 (N_39390,N_38903,N_38654);
nand U39391 (N_39391,N_38864,N_38764);
or U39392 (N_39392,N_38600,N_38869);
nor U39393 (N_39393,N_38820,N_38700);
nand U39394 (N_39394,N_38862,N_38784);
nand U39395 (N_39395,N_38945,N_38803);
or U39396 (N_39396,N_38528,N_38957);
nor U39397 (N_39397,N_38613,N_38800);
or U39398 (N_39398,N_38941,N_38658);
nand U39399 (N_39399,N_38744,N_38946);
or U39400 (N_39400,N_38785,N_38654);
nand U39401 (N_39401,N_38581,N_38783);
or U39402 (N_39402,N_38749,N_38882);
or U39403 (N_39403,N_38964,N_38913);
and U39404 (N_39404,N_38922,N_38611);
and U39405 (N_39405,N_38899,N_38849);
xor U39406 (N_39406,N_38726,N_38707);
nor U39407 (N_39407,N_38582,N_38887);
nor U39408 (N_39408,N_38554,N_38796);
and U39409 (N_39409,N_38608,N_38733);
nor U39410 (N_39410,N_38685,N_38969);
or U39411 (N_39411,N_38668,N_38501);
nor U39412 (N_39412,N_38913,N_38831);
nor U39413 (N_39413,N_38639,N_38605);
and U39414 (N_39414,N_38981,N_38931);
or U39415 (N_39415,N_38921,N_38863);
and U39416 (N_39416,N_38588,N_38885);
nor U39417 (N_39417,N_38607,N_38716);
nand U39418 (N_39418,N_38594,N_38912);
nor U39419 (N_39419,N_38543,N_38826);
or U39420 (N_39420,N_38672,N_38734);
and U39421 (N_39421,N_38828,N_38664);
nor U39422 (N_39422,N_38740,N_38512);
or U39423 (N_39423,N_38980,N_38677);
nand U39424 (N_39424,N_38753,N_38995);
xnor U39425 (N_39425,N_38728,N_38896);
or U39426 (N_39426,N_38955,N_38986);
or U39427 (N_39427,N_38828,N_38991);
and U39428 (N_39428,N_38519,N_38808);
nand U39429 (N_39429,N_38555,N_38644);
nand U39430 (N_39430,N_38897,N_38686);
xnor U39431 (N_39431,N_38766,N_38902);
xnor U39432 (N_39432,N_38862,N_38821);
and U39433 (N_39433,N_38863,N_38917);
nor U39434 (N_39434,N_38551,N_38542);
and U39435 (N_39435,N_38946,N_38957);
nor U39436 (N_39436,N_38954,N_38524);
xor U39437 (N_39437,N_38714,N_38819);
nor U39438 (N_39438,N_38617,N_38717);
or U39439 (N_39439,N_38620,N_38821);
nor U39440 (N_39440,N_38897,N_38656);
or U39441 (N_39441,N_38726,N_38719);
and U39442 (N_39442,N_38793,N_38679);
nand U39443 (N_39443,N_38726,N_38692);
nor U39444 (N_39444,N_38601,N_38527);
nor U39445 (N_39445,N_38878,N_38725);
or U39446 (N_39446,N_38563,N_38722);
xor U39447 (N_39447,N_38523,N_38760);
nor U39448 (N_39448,N_38710,N_38847);
or U39449 (N_39449,N_38842,N_38757);
or U39450 (N_39450,N_38869,N_38832);
nor U39451 (N_39451,N_38525,N_38591);
nor U39452 (N_39452,N_38874,N_38667);
or U39453 (N_39453,N_38509,N_38505);
xnor U39454 (N_39454,N_38963,N_38661);
nand U39455 (N_39455,N_38527,N_38609);
nand U39456 (N_39456,N_38570,N_38837);
or U39457 (N_39457,N_38653,N_38923);
nor U39458 (N_39458,N_38725,N_38869);
nor U39459 (N_39459,N_38992,N_38904);
nand U39460 (N_39460,N_38873,N_38930);
or U39461 (N_39461,N_38700,N_38892);
nand U39462 (N_39462,N_38895,N_38502);
nor U39463 (N_39463,N_38666,N_38806);
and U39464 (N_39464,N_38818,N_38513);
or U39465 (N_39465,N_38665,N_38796);
nor U39466 (N_39466,N_38944,N_38929);
and U39467 (N_39467,N_38983,N_38998);
or U39468 (N_39468,N_38509,N_38608);
nor U39469 (N_39469,N_38681,N_38814);
and U39470 (N_39470,N_38547,N_38726);
and U39471 (N_39471,N_38912,N_38504);
nand U39472 (N_39472,N_38584,N_38949);
or U39473 (N_39473,N_38747,N_38828);
or U39474 (N_39474,N_38765,N_38589);
nand U39475 (N_39475,N_38674,N_38910);
xor U39476 (N_39476,N_38740,N_38535);
or U39477 (N_39477,N_38812,N_38911);
nand U39478 (N_39478,N_38654,N_38933);
nand U39479 (N_39479,N_38744,N_38755);
nor U39480 (N_39480,N_38538,N_38608);
nand U39481 (N_39481,N_38504,N_38651);
nor U39482 (N_39482,N_38977,N_38905);
or U39483 (N_39483,N_38841,N_38963);
nand U39484 (N_39484,N_38688,N_38590);
or U39485 (N_39485,N_38968,N_38644);
and U39486 (N_39486,N_38622,N_38531);
nor U39487 (N_39487,N_38972,N_38639);
and U39488 (N_39488,N_38748,N_38563);
or U39489 (N_39489,N_38611,N_38668);
nand U39490 (N_39490,N_38920,N_38800);
or U39491 (N_39491,N_38606,N_38776);
nor U39492 (N_39492,N_38789,N_38741);
nor U39493 (N_39493,N_38542,N_38568);
nand U39494 (N_39494,N_38557,N_38901);
or U39495 (N_39495,N_38938,N_38910);
xor U39496 (N_39496,N_38666,N_38645);
or U39497 (N_39497,N_38813,N_38887);
xnor U39498 (N_39498,N_38605,N_38953);
or U39499 (N_39499,N_38791,N_38589);
nand U39500 (N_39500,N_39023,N_39290);
nand U39501 (N_39501,N_39407,N_39411);
nand U39502 (N_39502,N_39034,N_39471);
xnor U39503 (N_39503,N_39463,N_39244);
nor U39504 (N_39504,N_39044,N_39350);
and U39505 (N_39505,N_39067,N_39490);
or U39506 (N_39506,N_39381,N_39439);
nor U39507 (N_39507,N_39013,N_39349);
or U39508 (N_39508,N_39408,N_39230);
nor U39509 (N_39509,N_39243,N_39309);
and U39510 (N_39510,N_39142,N_39080);
and U39511 (N_39511,N_39178,N_39160);
and U39512 (N_39512,N_39491,N_39311);
or U39513 (N_39513,N_39330,N_39380);
nor U39514 (N_39514,N_39064,N_39006);
nor U39515 (N_39515,N_39271,N_39338);
nor U39516 (N_39516,N_39263,N_39074);
or U39517 (N_39517,N_39340,N_39397);
xor U39518 (N_39518,N_39337,N_39334);
nor U39519 (N_39519,N_39120,N_39116);
nand U39520 (N_39520,N_39379,N_39363);
or U39521 (N_39521,N_39409,N_39358);
or U39522 (N_39522,N_39398,N_39422);
or U39523 (N_39523,N_39322,N_39180);
nor U39524 (N_39524,N_39113,N_39227);
and U39525 (N_39525,N_39216,N_39470);
or U39526 (N_39526,N_39351,N_39445);
or U39527 (N_39527,N_39114,N_39012);
or U39528 (N_39528,N_39028,N_39466);
and U39529 (N_39529,N_39049,N_39265);
nand U39530 (N_39530,N_39159,N_39220);
and U39531 (N_39531,N_39250,N_39026);
and U39532 (N_39532,N_39177,N_39193);
or U39533 (N_39533,N_39373,N_39016);
or U39534 (N_39534,N_39268,N_39229);
nand U39535 (N_39535,N_39137,N_39007);
nand U39536 (N_39536,N_39254,N_39295);
and U39537 (N_39537,N_39121,N_39175);
and U39538 (N_39538,N_39155,N_39205);
or U39539 (N_39539,N_39460,N_39454);
and U39540 (N_39540,N_39434,N_39017);
nand U39541 (N_39541,N_39371,N_39222);
nor U39542 (N_39542,N_39069,N_39102);
or U39543 (N_39543,N_39435,N_39468);
nor U39544 (N_39544,N_39019,N_39405);
xor U39545 (N_39545,N_39276,N_39267);
or U39546 (N_39546,N_39071,N_39415);
nand U39547 (N_39547,N_39496,N_39047);
nand U39548 (N_39548,N_39237,N_39057);
nor U39549 (N_39549,N_39200,N_39369);
nor U39550 (N_39550,N_39106,N_39467);
nor U39551 (N_39551,N_39241,N_39027);
nor U39552 (N_39552,N_39386,N_39084);
nor U39553 (N_39553,N_39425,N_39077);
xor U39554 (N_39554,N_39412,N_39389);
and U39555 (N_39555,N_39487,N_39148);
and U39556 (N_39556,N_39211,N_39005);
or U39557 (N_39557,N_39426,N_39157);
xor U39558 (N_39558,N_39210,N_39105);
xor U39559 (N_39559,N_39011,N_39300);
nand U39560 (N_39560,N_39251,N_39192);
xor U39561 (N_39561,N_39461,N_39119);
nand U39562 (N_39562,N_39286,N_39372);
nor U39563 (N_39563,N_39219,N_39225);
xor U39564 (N_39564,N_39394,N_39194);
nand U39565 (N_39565,N_39070,N_39449);
or U39566 (N_39566,N_39094,N_39335);
nor U39567 (N_39567,N_39145,N_39190);
nor U39568 (N_39568,N_39202,N_39072);
nand U39569 (N_39569,N_39401,N_39383);
xor U39570 (N_39570,N_39078,N_39499);
nor U39571 (N_39571,N_39170,N_39498);
or U39572 (N_39572,N_39296,N_39400);
nor U39573 (N_39573,N_39103,N_39260);
or U39574 (N_39574,N_39326,N_39274);
and U39575 (N_39575,N_39485,N_39087);
or U39576 (N_39576,N_39109,N_39442);
nand U39577 (N_39577,N_39493,N_39127);
nand U39578 (N_39578,N_39291,N_39390);
nor U39579 (N_39579,N_39388,N_39325);
or U39580 (N_39580,N_39375,N_39030);
nand U39581 (N_39581,N_39317,N_39336);
and U39582 (N_39582,N_39098,N_39089);
xor U39583 (N_39583,N_39421,N_39320);
and U39584 (N_39584,N_39059,N_39416);
nor U39585 (N_39585,N_39393,N_39134);
nor U39586 (N_39586,N_39060,N_39152);
or U39587 (N_39587,N_39143,N_39451);
nor U39588 (N_39588,N_39199,N_39303);
nor U39589 (N_39589,N_39450,N_39359);
or U39590 (N_39590,N_39289,N_39298);
and U39591 (N_39591,N_39437,N_39304);
or U39592 (N_39592,N_39189,N_39203);
nor U39593 (N_39593,N_39124,N_39443);
xnor U39594 (N_39594,N_39208,N_39294);
nor U39595 (N_39595,N_39021,N_39112);
or U39596 (N_39596,N_39306,N_39333);
nor U39597 (N_39597,N_39231,N_39139);
and U39598 (N_39598,N_39420,N_39249);
nand U39599 (N_39599,N_39036,N_39083);
nor U39600 (N_39600,N_39436,N_39462);
or U39601 (N_39601,N_39419,N_39051);
nand U39602 (N_39602,N_39004,N_39223);
nand U39603 (N_39603,N_39275,N_39088);
and U39604 (N_39604,N_39272,N_39031);
and U39605 (N_39605,N_39014,N_39423);
or U39606 (N_39606,N_39050,N_39187);
nor U39607 (N_39607,N_39154,N_39475);
and U39608 (N_39608,N_39151,N_39236);
and U39609 (N_39609,N_39032,N_39431);
nor U39610 (N_39610,N_39488,N_39346);
and U39611 (N_39611,N_39201,N_39195);
nor U39612 (N_39612,N_39446,N_39438);
nor U39613 (N_39613,N_39108,N_39062);
nor U39614 (N_39614,N_39280,N_39022);
and U39615 (N_39615,N_39406,N_39384);
nand U39616 (N_39616,N_39395,N_39055);
nand U39617 (N_39617,N_39382,N_39115);
nand U39618 (N_39618,N_39003,N_39374);
or U39619 (N_39619,N_39361,N_39182);
nand U39620 (N_39620,N_39345,N_39138);
or U39621 (N_39621,N_39213,N_39186);
nand U39622 (N_39622,N_39489,N_39125);
and U39623 (N_39623,N_39433,N_39258);
and U39624 (N_39624,N_39215,N_39314);
nor U39625 (N_39625,N_39302,N_39339);
and U39626 (N_39626,N_39344,N_39206);
and U39627 (N_39627,N_39262,N_39226);
xor U39628 (N_39628,N_39224,N_39081);
or U39629 (N_39629,N_39355,N_39166);
nand U39630 (N_39630,N_39357,N_39188);
or U39631 (N_39631,N_39378,N_39473);
nor U39632 (N_39632,N_39207,N_39129);
nand U39633 (N_39633,N_39284,N_39347);
nor U39634 (N_39634,N_39441,N_39135);
or U39635 (N_39635,N_39354,N_39247);
or U39636 (N_39636,N_39292,N_39196);
or U39637 (N_39637,N_39429,N_39097);
or U39638 (N_39638,N_39174,N_39456);
or U39639 (N_39639,N_39048,N_39353);
nor U39640 (N_39640,N_39283,N_39368);
nand U39641 (N_39641,N_39252,N_39301);
nand U39642 (N_39642,N_39130,N_39043);
or U39643 (N_39643,N_39321,N_39136);
nand U39644 (N_39644,N_39474,N_39418);
nand U39645 (N_39645,N_39492,N_39144);
xnor U39646 (N_39646,N_39000,N_39107);
xnor U39647 (N_39647,N_39399,N_39233);
or U39648 (N_39648,N_39288,N_39458);
nand U39649 (N_39649,N_39269,N_39327);
or U39650 (N_39650,N_39008,N_39168);
and U39651 (N_39651,N_39228,N_39480);
xor U39652 (N_39652,N_39118,N_39217);
nand U39653 (N_39653,N_39285,N_39141);
or U39654 (N_39654,N_39185,N_39090);
xor U39655 (N_39655,N_39482,N_39156);
and U39656 (N_39656,N_39058,N_39246);
nor U39657 (N_39657,N_39056,N_39366);
nand U39658 (N_39658,N_39101,N_39305);
xor U39659 (N_39659,N_39128,N_39024);
nand U39660 (N_39660,N_39033,N_39015);
nor U39661 (N_39661,N_39427,N_39315);
nand U39662 (N_39662,N_39029,N_39256);
nor U39663 (N_39663,N_39172,N_39075);
nand U39664 (N_39664,N_39093,N_39095);
or U39665 (N_39665,N_39150,N_39001);
nand U39666 (N_39666,N_39387,N_39037);
nand U39667 (N_39667,N_39328,N_39440);
nand U39668 (N_39668,N_39171,N_39356);
and U39669 (N_39669,N_39376,N_39495);
nand U39670 (N_39670,N_39221,N_39279);
or U39671 (N_39671,N_39117,N_39483);
and U39672 (N_39672,N_39323,N_39486);
or U39673 (N_39673,N_39402,N_39164);
or U39674 (N_39674,N_39153,N_39253);
xor U39675 (N_39675,N_39140,N_39478);
nor U39676 (N_39676,N_39497,N_39410);
or U39677 (N_39677,N_39391,N_39133);
and U39678 (N_39678,N_39061,N_39257);
or U39679 (N_39679,N_39179,N_39082);
and U39680 (N_39680,N_39424,N_39099);
or U39681 (N_39681,N_39111,N_39010);
nor U39682 (N_39682,N_39018,N_39100);
xnor U39683 (N_39683,N_39123,N_39341);
or U39684 (N_39684,N_39161,N_39162);
and U39685 (N_39685,N_39293,N_39053);
or U39686 (N_39686,N_39131,N_39169);
xor U39687 (N_39687,N_39167,N_39039);
xor U39688 (N_39688,N_39181,N_39240);
and U39689 (N_39689,N_39417,N_39204);
nand U39690 (N_39690,N_39476,N_39319);
xor U39691 (N_39691,N_39209,N_39085);
or U39692 (N_39692,N_39430,N_39183);
or U39693 (N_39693,N_39038,N_39273);
nor U39694 (N_39694,N_39277,N_39362);
nor U39695 (N_39695,N_39367,N_39132);
nand U39696 (N_39696,N_39479,N_39104);
or U39697 (N_39697,N_39197,N_39270);
nand U39698 (N_39698,N_39232,N_39238);
nand U39699 (N_39699,N_39310,N_39235);
or U39700 (N_39700,N_39264,N_39191);
nor U39701 (N_39701,N_39299,N_39176);
nor U39702 (N_39702,N_39494,N_39052);
nor U39703 (N_39703,N_39234,N_39348);
and U39704 (N_39704,N_39365,N_39068);
and U39705 (N_39705,N_39477,N_39079);
xor U39706 (N_39706,N_39364,N_39464);
nor U39707 (N_39707,N_39149,N_39009);
and U39708 (N_39708,N_39331,N_39184);
nand U39709 (N_39709,N_39459,N_39042);
nand U39710 (N_39710,N_39020,N_39396);
nor U39711 (N_39711,N_39282,N_39096);
or U39712 (N_39712,N_39329,N_39242);
and U39713 (N_39713,N_39481,N_39414);
nand U39714 (N_39714,N_39122,N_39352);
nand U39715 (N_39715,N_39092,N_39469);
nand U39716 (N_39716,N_39370,N_39447);
or U39717 (N_39717,N_39248,N_39046);
nor U39718 (N_39718,N_39403,N_39035);
xnor U39719 (N_39719,N_39360,N_39472);
or U39720 (N_39720,N_39266,N_39218);
nand U39721 (N_39721,N_39065,N_39040);
nand U39722 (N_39722,N_39214,N_39324);
and U39723 (N_39723,N_39444,N_39054);
and U39724 (N_39724,N_39255,N_39281);
or U39725 (N_39725,N_39392,N_39428);
nand U39726 (N_39726,N_39312,N_39484);
and U39727 (N_39727,N_39147,N_39198);
or U39728 (N_39728,N_39158,N_39432);
nand U39729 (N_39729,N_39318,N_39342);
or U39730 (N_39730,N_39146,N_39041);
xnor U39731 (N_39731,N_39278,N_39073);
nor U39732 (N_39732,N_39091,N_39465);
nand U39733 (N_39733,N_39453,N_39126);
nor U39734 (N_39734,N_39110,N_39212);
xnor U39735 (N_39735,N_39457,N_39287);
nand U39736 (N_39736,N_39076,N_39413);
or U39737 (N_39737,N_39332,N_39343);
and U39738 (N_39738,N_39448,N_39002);
nand U39739 (N_39739,N_39045,N_39259);
nor U39740 (N_39740,N_39239,N_39163);
nor U39741 (N_39741,N_39452,N_39377);
nor U39742 (N_39742,N_39025,N_39404);
and U39743 (N_39743,N_39308,N_39316);
nor U39744 (N_39744,N_39063,N_39455);
nand U39745 (N_39745,N_39313,N_39385);
nand U39746 (N_39746,N_39297,N_39307);
and U39747 (N_39747,N_39066,N_39245);
and U39748 (N_39748,N_39173,N_39261);
nand U39749 (N_39749,N_39086,N_39165);
nor U39750 (N_39750,N_39187,N_39165);
or U39751 (N_39751,N_39499,N_39216);
nand U39752 (N_39752,N_39342,N_39141);
or U39753 (N_39753,N_39147,N_39274);
nor U39754 (N_39754,N_39346,N_39221);
nor U39755 (N_39755,N_39182,N_39452);
nand U39756 (N_39756,N_39204,N_39432);
nor U39757 (N_39757,N_39412,N_39050);
and U39758 (N_39758,N_39111,N_39206);
or U39759 (N_39759,N_39303,N_39134);
and U39760 (N_39760,N_39425,N_39442);
and U39761 (N_39761,N_39175,N_39084);
nor U39762 (N_39762,N_39313,N_39310);
nor U39763 (N_39763,N_39270,N_39485);
xnor U39764 (N_39764,N_39152,N_39326);
nor U39765 (N_39765,N_39134,N_39180);
or U39766 (N_39766,N_39370,N_39140);
or U39767 (N_39767,N_39240,N_39381);
and U39768 (N_39768,N_39173,N_39373);
or U39769 (N_39769,N_39406,N_39495);
nand U39770 (N_39770,N_39066,N_39145);
or U39771 (N_39771,N_39109,N_39040);
and U39772 (N_39772,N_39453,N_39050);
nand U39773 (N_39773,N_39469,N_39379);
and U39774 (N_39774,N_39276,N_39363);
or U39775 (N_39775,N_39284,N_39298);
and U39776 (N_39776,N_39470,N_39032);
or U39777 (N_39777,N_39161,N_39337);
or U39778 (N_39778,N_39296,N_39052);
nor U39779 (N_39779,N_39374,N_39054);
nand U39780 (N_39780,N_39262,N_39368);
and U39781 (N_39781,N_39049,N_39272);
or U39782 (N_39782,N_39267,N_39422);
nand U39783 (N_39783,N_39447,N_39153);
or U39784 (N_39784,N_39139,N_39128);
or U39785 (N_39785,N_39240,N_39026);
nand U39786 (N_39786,N_39439,N_39369);
and U39787 (N_39787,N_39265,N_39108);
nand U39788 (N_39788,N_39166,N_39226);
nor U39789 (N_39789,N_39441,N_39208);
or U39790 (N_39790,N_39053,N_39369);
and U39791 (N_39791,N_39078,N_39021);
or U39792 (N_39792,N_39377,N_39406);
or U39793 (N_39793,N_39152,N_39433);
nand U39794 (N_39794,N_39061,N_39187);
nor U39795 (N_39795,N_39431,N_39418);
and U39796 (N_39796,N_39105,N_39439);
nand U39797 (N_39797,N_39091,N_39325);
xor U39798 (N_39798,N_39077,N_39258);
nand U39799 (N_39799,N_39359,N_39495);
xnor U39800 (N_39800,N_39475,N_39133);
nand U39801 (N_39801,N_39384,N_39415);
nand U39802 (N_39802,N_39409,N_39477);
and U39803 (N_39803,N_39161,N_39467);
and U39804 (N_39804,N_39255,N_39153);
and U39805 (N_39805,N_39152,N_39171);
or U39806 (N_39806,N_39226,N_39101);
xor U39807 (N_39807,N_39309,N_39286);
nor U39808 (N_39808,N_39339,N_39095);
xor U39809 (N_39809,N_39112,N_39448);
xor U39810 (N_39810,N_39415,N_39077);
or U39811 (N_39811,N_39436,N_39397);
nor U39812 (N_39812,N_39217,N_39009);
or U39813 (N_39813,N_39335,N_39482);
xor U39814 (N_39814,N_39444,N_39172);
or U39815 (N_39815,N_39067,N_39121);
nand U39816 (N_39816,N_39406,N_39378);
or U39817 (N_39817,N_39237,N_39248);
or U39818 (N_39818,N_39159,N_39326);
nand U39819 (N_39819,N_39466,N_39473);
nor U39820 (N_39820,N_39364,N_39435);
nand U39821 (N_39821,N_39397,N_39169);
or U39822 (N_39822,N_39176,N_39207);
and U39823 (N_39823,N_39105,N_39076);
and U39824 (N_39824,N_39485,N_39138);
or U39825 (N_39825,N_39294,N_39103);
nor U39826 (N_39826,N_39456,N_39074);
nor U39827 (N_39827,N_39114,N_39080);
nand U39828 (N_39828,N_39228,N_39369);
and U39829 (N_39829,N_39030,N_39118);
or U39830 (N_39830,N_39263,N_39327);
nand U39831 (N_39831,N_39052,N_39144);
or U39832 (N_39832,N_39124,N_39298);
nor U39833 (N_39833,N_39368,N_39033);
nor U39834 (N_39834,N_39186,N_39040);
nor U39835 (N_39835,N_39177,N_39067);
nor U39836 (N_39836,N_39422,N_39216);
xnor U39837 (N_39837,N_39252,N_39150);
nand U39838 (N_39838,N_39289,N_39477);
xnor U39839 (N_39839,N_39139,N_39482);
or U39840 (N_39840,N_39264,N_39110);
nand U39841 (N_39841,N_39063,N_39350);
nor U39842 (N_39842,N_39431,N_39274);
or U39843 (N_39843,N_39309,N_39406);
xnor U39844 (N_39844,N_39079,N_39478);
and U39845 (N_39845,N_39229,N_39259);
nand U39846 (N_39846,N_39145,N_39027);
nand U39847 (N_39847,N_39318,N_39199);
nor U39848 (N_39848,N_39175,N_39076);
or U39849 (N_39849,N_39388,N_39444);
and U39850 (N_39850,N_39040,N_39488);
or U39851 (N_39851,N_39176,N_39032);
nand U39852 (N_39852,N_39074,N_39353);
xnor U39853 (N_39853,N_39052,N_39241);
or U39854 (N_39854,N_39234,N_39437);
nor U39855 (N_39855,N_39456,N_39284);
nand U39856 (N_39856,N_39013,N_39177);
nand U39857 (N_39857,N_39415,N_39390);
and U39858 (N_39858,N_39375,N_39259);
or U39859 (N_39859,N_39439,N_39033);
nor U39860 (N_39860,N_39453,N_39404);
nand U39861 (N_39861,N_39232,N_39226);
or U39862 (N_39862,N_39088,N_39373);
nand U39863 (N_39863,N_39102,N_39153);
nor U39864 (N_39864,N_39062,N_39348);
nand U39865 (N_39865,N_39091,N_39385);
nor U39866 (N_39866,N_39304,N_39045);
or U39867 (N_39867,N_39194,N_39047);
nand U39868 (N_39868,N_39384,N_39131);
nor U39869 (N_39869,N_39285,N_39267);
and U39870 (N_39870,N_39210,N_39487);
or U39871 (N_39871,N_39483,N_39297);
and U39872 (N_39872,N_39410,N_39106);
nor U39873 (N_39873,N_39312,N_39265);
nand U39874 (N_39874,N_39309,N_39378);
nor U39875 (N_39875,N_39069,N_39046);
or U39876 (N_39876,N_39059,N_39228);
and U39877 (N_39877,N_39000,N_39054);
nand U39878 (N_39878,N_39027,N_39015);
nor U39879 (N_39879,N_39043,N_39107);
nand U39880 (N_39880,N_39177,N_39348);
nor U39881 (N_39881,N_39143,N_39199);
xor U39882 (N_39882,N_39419,N_39000);
xor U39883 (N_39883,N_39224,N_39082);
and U39884 (N_39884,N_39123,N_39221);
and U39885 (N_39885,N_39232,N_39228);
nand U39886 (N_39886,N_39287,N_39431);
nor U39887 (N_39887,N_39352,N_39135);
and U39888 (N_39888,N_39077,N_39231);
or U39889 (N_39889,N_39247,N_39216);
or U39890 (N_39890,N_39058,N_39253);
or U39891 (N_39891,N_39007,N_39051);
nand U39892 (N_39892,N_39289,N_39170);
and U39893 (N_39893,N_39354,N_39269);
or U39894 (N_39894,N_39100,N_39231);
nand U39895 (N_39895,N_39118,N_39322);
and U39896 (N_39896,N_39019,N_39479);
nand U39897 (N_39897,N_39386,N_39024);
and U39898 (N_39898,N_39084,N_39225);
xor U39899 (N_39899,N_39412,N_39303);
xnor U39900 (N_39900,N_39389,N_39322);
nand U39901 (N_39901,N_39165,N_39048);
or U39902 (N_39902,N_39073,N_39045);
or U39903 (N_39903,N_39313,N_39395);
nand U39904 (N_39904,N_39241,N_39153);
or U39905 (N_39905,N_39208,N_39494);
and U39906 (N_39906,N_39378,N_39349);
and U39907 (N_39907,N_39296,N_39096);
xnor U39908 (N_39908,N_39093,N_39311);
nor U39909 (N_39909,N_39100,N_39282);
and U39910 (N_39910,N_39332,N_39180);
and U39911 (N_39911,N_39050,N_39247);
xnor U39912 (N_39912,N_39169,N_39250);
nor U39913 (N_39913,N_39070,N_39220);
or U39914 (N_39914,N_39395,N_39176);
or U39915 (N_39915,N_39179,N_39072);
nor U39916 (N_39916,N_39055,N_39086);
or U39917 (N_39917,N_39170,N_39393);
or U39918 (N_39918,N_39009,N_39175);
and U39919 (N_39919,N_39056,N_39000);
xor U39920 (N_39920,N_39063,N_39368);
or U39921 (N_39921,N_39262,N_39162);
nor U39922 (N_39922,N_39466,N_39096);
nand U39923 (N_39923,N_39447,N_39166);
nor U39924 (N_39924,N_39118,N_39491);
nand U39925 (N_39925,N_39370,N_39253);
nand U39926 (N_39926,N_39434,N_39038);
xnor U39927 (N_39927,N_39023,N_39038);
nor U39928 (N_39928,N_39428,N_39284);
nand U39929 (N_39929,N_39070,N_39054);
nand U39930 (N_39930,N_39461,N_39131);
and U39931 (N_39931,N_39192,N_39475);
xor U39932 (N_39932,N_39243,N_39151);
nand U39933 (N_39933,N_39256,N_39333);
nor U39934 (N_39934,N_39367,N_39306);
nand U39935 (N_39935,N_39279,N_39007);
and U39936 (N_39936,N_39473,N_39125);
and U39937 (N_39937,N_39335,N_39193);
nor U39938 (N_39938,N_39262,N_39388);
or U39939 (N_39939,N_39207,N_39292);
or U39940 (N_39940,N_39259,N_39063);
nor U39941 (N_39941,N_39208,N_39194);
or U39942 (N_39942,N_39454,N_39085);
nand U39943 (N_39943,N_39003,N_39454);
and U39944 (N_39944,N_39271,N_39021);
and U39945 (N_39945,N_39476,N_39257);
xnor U39946 (N_39946,N_39244,N_39314);
nand U39947 (N_39947,N_39167,N_39112);
and U39948 (N_39948,N_39332,N_39123);
nand U39949 (N_39949,N_39450,N_39290);
or U39950 (N_39950,N_39250,N_39491);
or U39951 (N_39951,N_39475,N_39072);
nand U39952 (N_39952,N_39198,N_39431);
nor U39953 (N_39953,N_39462,N_39370);
nand U39954 (N_39954,N_39308,N_39045);
and U39955 (N_39955,N_39183,N_39027);
or U39956 (N_39956,N_39118,N_39086);
or U39957 (N_39957,N_39375,N_39456);
nor U39958 (N_39958,N_39463,N_39250);
nand U39959 (N_39959,N_39070,N_39436);
xnor U39960 (N_39960,N_39468,N_39003);
or U39961 (N_39961,N_39341,N_39027);
xnor U39962 (N_39962,N_39311,N_39280);
or U39963 (N_39963,N_39004,N_39130);
or U39964 (N_39964,N_39467,N_39316);
nor U39965 (N_39965,N_39004,N_39164);
xor U39966 (N_39966,N_39045,N_39058);
nand U39967 (N_39967,N_39130,N_39073);
nand U39968 (N_39968,N_39167,N_39492);
xnor U39969 (N_39969,N_39414,N_39031);
nor U39970 (N_39970,N_39418,N_39337);
nand U39971 (N_39971,N_39360,N_39375);
xnor U39972 (N_39972,N_39159,N_39020);
nand U39973 (N_39973,N_39188,N_39102);
nor U39974 (N_39974,N_39428,N_39114);
nand U39975 (N_39975,N_39056,N_39032);
and U39976 (N_39976,N_39431,N_39486);
nand U39977 (N_39977,N_39478,N_39331);
and U39978 (N_39978,N_39480,N_39402);
nor U39979 (N_39979,N_39298,N_39204);
or U39980 (N_39980,N_39200,N_39419);
xor U39981 (N_39981,N_39130,N_39187);
xor U39982 (N_39982,N_39369,N_39120);
nand U39983 (N_39983,N_39382,N_39206);
or U39984 (N_39984,N_39239,N_39475);
or U39985 (N_39985,N_39289,N_39305);
nor U39986 (N_39986,N_39405,N_39477);
nor U39987 (N_39987,N_39216,N_39129);
and U39988 (N_39988,N_39310,N_39058);
and U39989 (N_39989,N_39276,N_39033);
nand U39990 (N_39990,N_39449,N_39095);
or U39991 (N_39991,N_39265,N_39248);
nor U39992 (N_39992,N_39218,N_39322);
nor U39993 (N_39993,N_39390,N_39161);
nor U39994 (N_39994,N_39114,N_39065);
or U39995 (N_39995,N_39429,N_39093);
nand U39996 (N_39996,N_39043,N_39069);
or U39997 (N_39997,N_39340,N_39336);
and U39998 (N_39998,N_39001,N_39334);
and U39999 (N_39999,N_39380,N_39170);
nor U40000 (N_40000,N_39789,N_39715);
nand U40001 (N_40001,N_39756,N_39565);
nor U40002 (N_40002,N_39670,N_39511);
and U40003 (N_40003,N_39945,N_39628);
or U40004 (N_40004,N_39871,N_39588);
nor U40005 (N_40005,N_39958,N_39865);
or U40006 (N_40006,N_39859,N_39621);
nand U40007 (N_40007,N_39584,N_39652);
and U40008 (N_40008,N_39528,N_39925);
nand U40009 (N_40009,N_39981,N_39940);
or U40010 (N_40010,N_39881,N_39897);
or U40011 (N_40011,N_39807,N_39610);
or U40012 (N_40012,N_39513,N_39933);
xor U40013 (N_40013,N_39998,N_39919);
nor U40014 (N_40014,N_39834,N_39839);
and U40015 (N_40015,N_39913,N_39855);
or U40016 (N_40016,N_39591,N_39814);
nand U40017 (N_40017,N_39861,N_39990);
or U40018 (N_40018,N_39595,N_39809);
and U40019 (N_40019,N_39792,N_39550);
nand U40020 (N_40020,N_39930,N_39651);
and U40021 (N_40021,N_39934,N_39680);
nor U40022 (N_40022,N_39711,N_39972);
and U40023 (N_40023,N_39667,N_39587);
xor U40024 (N_40024,N_39509,N_39841);
or U40025 (N_40025,N_39574,N_39596);
xnor U40026 (N_40026,N_39902,N_39782);
or U40027 (N_40027,N_39936,N_39806);
nor U40028 (N_40028,N_39776,N_39532);
nor U40029 (N_40029,N_39863,N_39672);
nor U40030 (N_40030,N_39744,N_39818);
xnor U40031 (N_40031,N_39552,N_39837);
or U40032 (N_40032,N_39766,N_39907);
nor U40033 (N_40033,N_39567,N_39770);
nor U40034 (N_40034,N_39916,N_39838);
xor U40035 (N_40035,N_39617,N_39531);
or U40036 (N_40036,N_39835,N_39649);
nor U40037 (N_40037,N_39583,N_39971);
nor U40038 (N_40038,N_39741,N_39592);
nor U40039 (N_40039,N_39943,N_39718);
xnor U40040 (N_40040,N_39955,N_39903);
or U40041 (N_40041,N_39501,N_39740);
or U40042 (N_40042,N_39638,N_39753);
and U40043 (N_40043,N_39864,N_39954);
or U40044 (N_40044,N_39962,N_39856);
nand U40045 (N_40045,N_39696,N_39573);
nor U40046 (N_40046,N_39685,N_39602);
or U40047 (N_40047,N_39643,N_39904);
or U40048 (N_40048,N_39576,N_39558);
and U40049 (N_40049,N_39822,N_39815);
xor U40050 (N_40050,N_39735,N_39580);
nor U40051 (N_40051,N_39849,N_39798);
nand U40052 (N_40052,N_39830,N_39537);
nand U40053 (N_40053,N_39957,N_39797);
and U40054 (N_40054,N_39547,N_39745);
nand U40055 (N_40055,N_39877,N_39706);
nand U40056 (N_40056,N_39542,N_39688);
nor U40057 (N_40057,N_39662,N_39655);
xnor U40058 (N_40058,N_39534,N_39812);
and U40059 (N_40059,N_39844,N_39700);
nor U40060 (N_40060,N_39641,N_39951);
and U40061 (N_40061,N_39761,N_39612);
or U40062 (N_40062,N_39909,N_39613);
nor U40063 (N_40063,N_39698,N_39999);
nor U40064 (N_40064,N_39654,N_39701);
or U40065 (N_40065,N_39887,N_39663);
nor U40066 (N_40066,N_39626,N_39977);
nor U40067 (N_40067,N_39799,N_39647);
nand U40068 (N_40068,N_39950,N_39772);
or U40069 (N_40069,N_39522,N_39979);
and U40070 (N_40070,N_39608,N_39607);
nand U40071 (N_40071,N_39948,N_39747);
or U40072 (N_40072,N_39586,N_39773);
nand U40073 (N_40073,N_39525,N_39828);
and U40074 (N_40074,N_39676,N_39743);
nand U40075 (N_40075,N_39635,N_39899);
nand U40076 (N_40076,N_39751,N_39765);
or U40077 (N_40077,N_39679,N_39755);
nor U40078 (N_40078,N_39976,N_39619);
nor U40079 (N_40079,N_39504,N_39546);
nor U40080 (N_40080,N_39920,N_39896);
nor U40081 (N_40081,N_39737,N_39533);
nor U40082 (N_40082,N_39923,N_39924);
nor U40083 (N_40083,N_39529,N_39989);
nand U40084 (N_40084,N_39736,N_39823);
and U40085 (N_40085,N_39796,N_39598);
nor U40086 (N_40086,N_39867,N_39569);
xnor U40087 (N_40087,N_39810,N_39568);
xor U40088 (N_40088,N_39660,N_39536);
nor U40089 (N_40089,N_39911,N_39926);
or U40090 (N_40090,N_39702,N_39526);
and U40091 (N_40091,N_39746,N_39575);
and U40092 (N_40092,N_39886,N_39754);
nor U40093 (N_40093,N_39769,N_39614);
or U40094 (N_40094,N_39778,N_39921);
or U40095 (N_40095,N_39973,N_39703);
nor U40096 (N_40096,N_39601,N_39952);
nor U40097 (N_40097,N_39553,N_39514);
nand U40098 (N_40098,N_39953,N_39554);
or U40099 (N_40099,N_39787,N_39616);
and U40100 (N_40100,N_39908,N_39800);
and U40101 (N_40101,N_39767,N_39704);
nand U40102 (N_40102,N_39738,N_39975);
nand U40103 (N_40103,N_39960,N_39517);
nand U40104 (N_40104,N_39648,N_39712);
nand U40105 (N_40105,N_39503,N_39816);
xnor U40106 (N_40106,N_39846,N_39560);
or U40107 (N_40107,N_39803,N_39716);
nand U40108 (N_40108,N_39632,N_39611);
or U40109 (N_40109,N_39862,N_39910);
or U40110 (N_40110,N_39543,N_39980);
nor U40111 (N_40111,N_39956,N_39941);
nor U40112 (N_40112,N_39727,N_39931);
and U40113 (N_40113,N_39829,N_39914);
and U40114 (N_40114,N_39985,N_39674);
or U40115 (N_40115,N_39893,N_39771);
and U40116 (N_40116,N_39917,N_39997);
nand U40117 (N_40117,N_39637,N_39524);
nor U40118 (N_40118,N_39944,N_39555);
nor U40119 (N_40119,N_39545,N_39512);
xnor U40120 (N_40120,N_39656,N_39764);
nor U40121 (N_40121,N_39984,N_39840);
nand U40122 (N_40122,N_39996,N_39959);
nand U40123 (N_40123,N_39734,N_39889);
and U40124 (N_40124,N_39683,N_39847);
nor U40125 (N_40125,N_39857,N_39992);
and U40126 (N_40126,N_39538,N_39817);
and U40127 (N_40127,N_39609,N_39915);
nor U40128 (N_40128,N_39549,N_39686);
and U40129 (N_40129,N_39724,N_39901);
or U40130 (N_40130,N_39732,N_39681);
nand U40131 (N_40131,N_39579,N_39832);
nor U40132 (N_40132,N_39774,N_39742);
and U40133 (N_40133,N_39629,N_39988);
and U40134 (N_40134,N_39721,N_39819);
or U40135 (N_40135,N_39781,N_39780);
nand U40136 (N_40136,N_39882,N_39644);
and U40137 (N_40137,N_39697,N_39993);
xor U40138 (N_40138,N_39939,N_39577);
and U40139 (N_40139,N_39786,N_39821);
or U40140 (N_40140,N_39581,N_39946);
xor U40141 (N_40141,N_39891,N_39860);
nor U40142 (N_40142,N_39918,N_39539);
xor U40143 (N_40143,N_39603,N_39620);
nand U40144 (N_40144,N_39748,N_39827);
nand U40145 (N_40145,N_39604,N_39678);
nor U40146 (N_40146,N_39880,N_39937);
xor U40147 (N_40147,N_39804,N_39708);
xnor U40148 (N_40148,N_39883,N_39802);
nor U40149 (N_40149,N_39669,N_39605);
nor U40150 (N_40150,N_39873,N_39725);
xor U40151 (N_40151,N_39540,N_39673);
and U40152 (N_40152,N_39890,N_39661);
and U40153 (N_40153,N_39653,N_39878);
xnor U40154 (N_40154,N_39559,N_39983);
or U40155 (N_40155,N_39942,N_39659);
nor U40156 (N_40156,N_39900,N_39717);
nand U40157 (N_40157,N_39582,N_39790);
xnor U40158 (N_40158,N_39530,N_39518);
nor U40159 (N_40159,N_39723,N_39500);
xnor U40160 (N_40160,N_39801,N_39519);
or U40161 (N_40161,N_39675,N_39845);
or U40162 (N_40162,N_39947,N_39820);
xor U40163 (N_40163,N_39759,N_39594);
and U40164 (N_40164,N_39833,N_39692);
xor U40165 (N_40165,N_39720,N_39710);
nand U40166 (N_40166,N_39589,N_39929);
and U40167 (N_40167,N_39965,N_39788);
or U40168 (N_40168,N_39968,N_39969);
or U40169 (N_40169,N_39624,N_39987);
nor U40170 (N_40170,N_39775,N_39922);
or U40171 (N_40171,N_39682,N_39876);
or U40172 (N_40172,N_39777,N_39668);
and U40173 (N_40173,N_39763,N_39728);
or U40174 (N_40174,N_39813,N_39510);
nor U40175 (N_40175,N_39515,N_39694);
nor U40176 (N_40176,N_39695,N_39749);
nor U40177 (N_40177,N_39986,N_39758);
and U40178 (N_40178,N_39562,N_39677);
or U40179 (N_40179,N_39645,N_39808);
and U40180 (N_40180,N_39585,N_39627);
xnor U40181 (N_40181,N_39831,N_39722);
nand U40182 (N_40182,N_39507,N_39684);
nor U40183 (N_40183,N_39625,N_39851);
and U40184 (N_40184,N_39731,N_39634);
nor U40185 (N_40185,N_39600,N_39666);
nor U40186 (N_40186,N_39689,N_39599);
and U40187 (N_40187,N_39884,N_39785);
or U40188 (N_40188,N_39633,N_39646);
nor U40189 (N_40189,N_39615,N_39779);
and U40190 (N_40190,N_39978,N_39564);
and U40191 (N_40191,N_39557,N_39793);
nor U40192 (N_40192,N_39502,N_39892);
nor U40193 (N_40193,N_39687,N_39719);
nor U40194 (N_40194,N_39966,N_39826);
nand U40195 (N_40195,N_39571,N_39665);
xor U40196 (N_40196,N_39853,N_39794);
nand U40197 (N_40197,N_39898,N_39894);
and U40198 (N_40198,N_39824,N_39709);
nor U40199 (N_40199,N_39578,N_39825);
xor U40200 (N_40200,N_39768,N_39527);
and U40201 (N_40201,N_39650,N_39693);
and U40202 (N_40202,N_39874,N_39872);
nand U40203 (N_40203,N_39606,N_39563);
or U40204 (N_40204,N_39783,N_39795);
nand U40205 (N_40205,N_39690,N_39691);
or U40206 (N_40206,N_39508,N_39566);
nand U40207 (N_40207,N_39854,N_39964);
nor U40208 (N_40208,N_39590,N_39805);
nand U40209 (N_40209,N_39593,N_39726);
and U40210 (N_40210,N_39705,N_39597);
nand U40211 (N_40211,N_39895,N_39982);
or U40212 (N_40212,N_39870,N_39762);
nor U40213 (N_40213,N_39963,N_39843);
xor U40214 (N_40214,N_39935,N_39888);
nor U40215 (N_40215,N_39505,N_39791);
or U40216 (N_40216,N_39561,N_39879);
xnor U40217 (N_40217,N_39636,N_39760);
or U40218 (N_40218,N_39961,N_39630);
or U40219 (N_40219,N_39535,N_39730);
and U40220 (N_40220,N_39967,N_39657);
nand U40221 (N_40221,N_39622,N_39750);
xnor U40222 (N_40222,N_39548,N_39906);
nor U40223 (N_40223,N_39739,N_39875);
nand U40224 (N_40224,N_39752,N_39928);
or U40225 (N_40225,N_39811,N_39784);
nor U40226 (N_40226,N_39905,N_39506);
or U40227 (N_40227,N_39885,N_39541);
and U40228 (N_40228,N_39848,N_39938);
or U40229 (N_40229,N_39713,N_39572);
xor U40230 (N_40230,N_39842,N_39836);
and U40231 (N_40231,N_39699,N_39757);
nor U40232 (N_40232,N_39714,N_39642);
xnor U40233 (N_40233,N_39664,N_39994);
nor U40234 (N_40234,N_39623,N_39974);
nor U40235 (N_40235,N_39516,N_39869);
and U40236 (N_40236,N_39631,N_39852);
or U40237 (N_40237,N_39521,N_39927);
and U40238 (N_40238,N_39556,N_39912);
xnor U40239 (N_40239,N_39850,N_39544);
nand U40240 (N_40240,N_39729,N_39671);
and U40241 (N_40241,N_39551,N_39970);
nand U40242 (N_40242,N_39570,N_39733);
nand U40243 (N_40243,N_39991,N_39858);
nand U40244 (N_40244,N_39868,N_39949);
nand U40245 (N_40245,N_39640,N_39523);
nor U40246 (N_40246,N_39707,N_39866);
or U40247 (N_40247,N_39658,N_39639);
or U40248 (N_40248,N_39618,N_39995);
and U40249 (N_40249,N_39932,N_39520);
nor U40250 (N_40250,N_39658,N_39599);
or U40251 (N_40251,N_39809,N_39728);
and U40252 (N_40252,N_39799,N_39954);
nand U40253 (N_40253,N_39569,N_39720);
or U40254 (N_40254,N_39714,N_39552);
nor U40255 (N_40255,N_39713,N_39947);
nor U40256 (N_40256,N_39886,N_39682);
nand U40257 (N_40257,N_39732,N_39946);
and U40258 (N_40258,N_39789,N_39887);
nor U40259 (N_40259,N_39992,N_39840);
xor U40260 (N_40260,N_39791,N_39609);
and U40261 (N_40261,N_39739,N_39519);
or U40262 (N_40262,N_39678,N_39652);
or U40263 (N_40263,N_39957,N_39833);
and U40264 (N_40264,N_39864,N_39710);
xor U40265 (N_40265,N_39770,N_39968);
or U40266 (N_40266,N_39586,N_39933);
and U40267 (N_40267,N_39953,N_39643);
xnor U40268 (N_40268,N_39877,N_39725);
or U40269 (N_40269,N_39743,N_39639);
nor U40270 (N_40270,N_39895,N_39988);
and U40271 (N_40271,N_39671,N_39878);
nor U40272 (N_40272,N_39561,N_39547);
nor U40273 (N_40273,N_39851,N_39888);
nand U40274 (N_40274,N_39701,N_39986);
xor U40275 (N_40275,N_39736,N_39579);
and U40276 (N_40276,N_39725,N_39992);
and U40277 (N_40277,N_39758,N_39558);
nand U40278 (N_40278,N_39851,N_39798);
and U40279 (N_40279,N_39535,N_39980);
or U40280 (N_40280,N_39955,N_39663);
nand U40281 (N_40281,N_39530,N_39813);
or U40282 (N_40282,N_39846,N_39951);
or U40283 (N_40283,N_39896,N_39966);
nor U40284 (N_40284,N_39674,N_39500);
nor U40285 (N_40285,N_39735,N_39622);
nor U40286 (N_40286,N_39530,N_39648);
and U40287 (N_40287,N_39522,N_39727);
nand U40288 (N_40288,N_39673,N_39815);
nand U40289 (N_40289,N_39923,N_39894);
or U40290 (N_40290,N_39709,N_39835);
or U40291 (N_40291,N_39687,N_39660);
or U40292 (N_40292,N_39792,N_39725);
nor U40293 (N_40293,N_39528,N_39708);
or U40294 (N_40294,N_39848,N_39752);
and U40295 (N_40295,N_39677,N_39710);
or U40296 (N_40296,N_39519,N_39753);
or U40297 (N_40297,N_39836,N_39701);
nand U40298 (N_40298,N_39561,N_39712);
and U40299 (N_40299,N_39631,N_39963);
and U40300 (N_40300,N_39616,N_39519);
nand U40301 (N_40301,N_39783,N_39623);
and U40302 (N_40302,N_39631,N_39954);
nand U40303 (N_40303,N_39958,N_39699);
nor U40304 (N_40304,N_39981,N_39625);
and U40305 (N_40305,N_39633,N_39518);
nor U40306 (N_40306,N_39687,N_39989);
and U40307 (N_40307,N_39653,N_39917);
nand U40308 (N_40308,N_39625,N_39861);
nand U40309 (N_40309,N_39976,N_39700);
and U40310 (N_40310,N_39600,N_39537);
nand U40311 (N_40311,N_39857,N_39906);
nor U40312 (N_40312,N_39852,N_39691);
or U40313 (N_40313,N_39899,N_39753);
nor U40314 (N_40314,N_39569,N_39577);
or U40315 (N_40315,N_39805,N_39648);
or U40316 (N_40316,N_39526,N_39904);
xnor U40317 (N_40317,N_39561,N_39748);
nand U40318 (N_40318,N_39660,N_39560);
and U40319 (N_40319,N_39513,N_39762);
nand U40320 (N_40320,N_39831,N_39546);
or U40321 (N_40321,N_39989,N_39779);
or U40322 (N_40322,N_39653,N_39569);
nand U40323 (N_40323,N_39659,N_39884);
nand U40324 (N_40324,N_39749,N_39859);
nand U40325 (N_40325,N_39843,N_39956);
or U40326 (N_40326,N_39762,N_39926);
nor U40327 (N_40327,N_39765,N_39792);
or U40328 (N_40328,N_39845,N_39735);
nor U40329 (N_40329,N_39858,N_39865);
nand U40330 (N_40330,N_39717,N_39911);
nor U40331 (N_40331,N_39635,N_39853);
and U40332 (N_40332,N_39783,N_39745);
nor U40333 (N_40333,N_39833,N_39583);
and U40334 (N_40334,N_39710,N_39899);
nor U40335 (N_40335,N_39622,N_39542);
and U40336 (N_40336,N_39624,N_39704);
xor U40337 (N_40337,N_39650,N_39642);
or U40338 (N_40338,N_39551,N_39920);
nand U40339 (N_40339,N_39780,N_39963);
nor U40340 (N_40340,N_39670,N_39636);
nand U40341 (N_40341,N_39855,N_39518);
nor U40342 (N_40342,N_39841,N_39982);
or U40343 (N_40343,N_39747,N_39748);
nand U40344 (N_40344,N_39568,N_39738);
nand U40345 (N_40345,N_39692,N_39895);
nand U40346 (N_40346,N_39884,N_39989);
or U40347 (N_40347,N_39661,N_39779);
xor U40348 (N_40348,N_39584,N_39839);
or U40349 (N_40349,N_39761,N_39791);
or U40350 (N_40350,N_39710,N_39698);
nand U40351 (N_40351,N_39779,N_39967);
or U40352 (N_40352,N_39689,N_39656);
or U40353 (N_40353,N_39890,N_39639);
and U40354 (N_40354,N_39600,N_39760);
nand U40355 (N_40355,N_39521,N_39920);
nor U40356 (N_40356,N_39926,N_39905);
or U40357 (N_40357,N_39986,N_39604);
nand U40358 (N_40358,N_39955,N_39645);
nand U40359 (N_40359,N_39795,N_39587);
nor U40360 (N_40360,N_39618,N_39915);
nand U40361 (N_40361,N_39520,N_39638);
or U40362 (N_40362,N_39608,N_39881);
or U40363 (N_40363,N_39642,N_39647);
and U40364 (N_40364,N_39994,N_39951);
or U40365 (N_40365,N_39686,N_39541);
or U40366 (N_40366,N_39895,N_39738);
or U40367 (N_40367,N_39951,N_39531);
or U40368 (N_40368,N_39835,N_39508);
nand U40369 (N_40369,N_39946,N_39608);
nor U40370 (N_40370,N_39813,N_39564);
or U40371 (N_40371,N_39873,N_39711);
or U40372 (N_40372,N_39810,N_39549);
nor U40373 (N_40373,N_39714,N_39812);
nor U40374 (N_40374,N_39870,N_39564);
nand U40375 (N_40375,N_39909,N_39571);
nor U40376 (N_40376,N_39733,N_39911);
and U40377 (N_40377,N_39658,N_39510);
xor U40378 (N_40378,N_39861,N_39940);
xor U40379 (N_40379,N_39994,N_39648);
nor U40380 (N_40380,N_39789,N_39763);
and U40381 (N_40381,N_39909,N_39911);
or U40382 (N_40382,N_39587,N_39564);
nor U40383 (N_40383,N_39815,N_39828);
and U40384 (N_40384,N_39920,N_39796);
xnor U40385 (N_40385,N_39783,N_39590);
or U40386 (N_40386,N_39609,N_39674);
nor U40387 (N_40387,N_39859,N_39593);
nor U40388 (N_40388,N_39813,N_39663);
or U40389 (N_40389,N_39865,N_39762);
or U40390 (N_40390,N_39593,N_39641);
nor U40391 (N_40391,N_39573,N_39811);
xor U40392 (N_40392,N_39891,N_39927);
xnor U40393 (N_40393,N_39534,N_39690);
and U40394 (N_40394,N_39944,N_39553);
nor U40395 (N_40395,N_39713,N_39887);
nand U40396 (N_40396,N_39567,N_39573);
nor U40397 (N_40397,N_39544,N_39971);
xor U40398 (N_40398,N_39916,N_39735);
xnor U40399 (N_40399,N_39760,N_39888);
nand U40400 (N_40400,N_39623,N_39918);
or U40401 (N_40401,N_39726,N_39883);
and U40402 (N_40402,N_39798,N_39980);
or U40403 (N_40403,N_39829,N_39951);
xor U40404 (N_40404,N_39716,N_39844);
nand U40405 (N_40405,N_39868,N_39558);
or U40406 (N_40406,N_39608,N_39969);
xor U40407 (N_40407,N_39903,N_39554);
and U40408 (N_40408,N_39891,N_39612);
and U40409 (N_40409,N_39838,N_39729);
nand U40410 (N_40410,N_39882,N_39688);
or U40411 (N_40411,N_39656,N_39810);
or U40412 (N_40412,N_39642,N_39560);
xor U40413 (N_40413,N_39902,N_39856);
or U40414 (N_40414,N_39730,N_39635);
nor U40415 (N_40415,N_39640,N_39594);
nand U40416 (N_40416,N_39705,N_39793);
and U40417 (N_40417,N_39706,N_39827);
and U40418 (N_40418,N_39693,N_39800);
and U40419 (N_40419,N_39598,N_39724);
and U40420 (N_40420,N_39646,N_39612);
or U40421 (N_40421,N_39663,N_39994);
and U40422 (N_40422,N_39666,N_39765);
and U40423 (N_40423,N_39582,N_39535);
nor U40424 (N_40424,N_39659,N_39686);
nand U40425 (N_40425,N_39594,N_39883);
xnor U40426 (N_40426,N_39950,N_39764);
xnor U40427 (N_40427,N_39931,N_39717);
and U40428 (N_40428,N_39793,N_39685);
and U40429 (N_40429,N_39841,N_39740);
or U40430 (N_40430,N_39805,N_39906);
nand U40431 (N_40431,N_39823,N_39963);
or U40432 (N_40432,N_39917,N_39553);
xor U40433 (N_40433,N_39906,N_39581);
and U40434 (N_40434,N_39562,N_39836);
nand U40435 (N_40435,N_39759,N_39680);
nand U40436 (N_40436,N_39612,N_39949);
or U40437 (N_40437,N_39889,N_39745);
or U40438 (N_40438,N_39601,N_39716);
or U40439 (N_40439,N_39744,N_39804);
xor U40440 (N_40440,N_39982,N_39761);
or U40441 (N_40441,N_39983,N_39632);
and U40442 (N_40442,N_39757,N_39538);
or U40443 (N_40443,N_39828,N_39734);
nor U40444 (N_40444,N_39975,N_39686);
and U40445 (N_40445,N_39776,N_39910);
nand U40446 (N_40446,N_39550,N_39874);
nor U40447 (N_40447,N_39730,N_39697);
or U40448 (N_40448,N_39692,N_39675);
or U40449 (N_40449,N_39534,N_39728);
and U40450 (N_40450,N_39546,N_39733);
xor U40451 (N_40451,N_39773,N_39745);
or U40452 (N_40452,N_39682,N_39671);
and U40453 (N_40453,N_39828,N_39609);
nand U40454 (N_40454,N_39740,N_39991);
nor U40455 (N_40455,N_39572,N_39879);
and U40456 (N_40456,N_39573,N_39533);
and U40457 (N_40457,N_39906,N_39684);
or U40458 (N_40458,N_39941,N_39636);
nor U40459 (N_40459,N_39725,N_39501);
xor U40460 (N_40460,N_39911,N_39685);
and U40461 (N_40461,N_39736,N_39617);
nand U40462 (N_40462,N_39978,N_39595);
or U40463 (N_40463,N_39613,N_39720);
nand U40464 (N_40464,N_39995,N_39773);
nor U40465 (N_40465,N_39518,N_39526);
nor U40466 (N_40466,N_39769,N_39795);
nor U40467 (N_40467,N_39694,N_39689);
or U40468 (N_40468,N_39819,N_39816);
nand U40469 (N_40469,N_39752,N_39724);
or U40470 (N_40470,N_39871,N_39800);
nor U40471 (N_40471,N_39979,N_39701);
xor U40472 (N_40472,N_39744,N_39928);
or U40473 (N_40473,N_39614,N_39561);
or U40474 (N_40474,N_39821,N_39502);
nor U40475 (N_40475,N_39909,N_39963);
xnor U40476 (N_40476,N_39561,N_39686);
nor U40477 (N_40477,N_39787,N_39501);
and U40478 (N_40478,N_39795,N_39570);
or U40479 (N_40479,N_39517,N_39741);
and U40480 (N_40480,N_39807,N_39993);
or U40481 (N_40481,N_39672,N_39746);
and U40482 (N_40482,N_39825,N_39963);
nand U40483 (N_40483,N_39550,N_39996);
or U40484 (N_40484,N_39618,N_39956);
nand U40485 (N_40485,N_39506,N_39960);
nand U40486 (N_40486,N_39869,N_39530);
nand U40487 (N_40487,N_39532,N_39762);
and U40488 (N_40488,N_39800,N_39596);
or U40489 (N_40489,N_39753,N_39583);
nor U40490 (N_40490,N_39794,N_39823);
and U40491 (N_40491,N_39630,N_39760);
and U40492 (N_40492,N_39954,N_39846);
nand U40493 (N_40493,N_39865,N_39649);
xnor U40494 (N_40494,N_39939,N_39919);
xnor U40495 (N_40495,N_39547,N_39870);
and U40496 (N_40496,N_39672,N_39655);
or U40497 (N_40497,N_39608,N_39506);
xnor U40498 (N_40498,N_39711,N_39941);
nor U40499 (N_40499,N_39729,N_39775);
nand U40500 (N_40500,N_40220,N_40302);
and U40501 (N_40501,N_40197,N_40296);
and U40502 (N_40502,N_40451,N_40295);
and U40503 (N_40503,N_40486,N_40400);
or U40504 (N_40504,N_40181,N_40315);
and U40505 (N_40505,N_40301,N_40361);
or U40506 (N_40506,N_40059,N_40484);
xnor U40507 (N_40507,N_40180,N_40353);
nand U40508 (N_40508,N_40282,N_40122);
xor U40509 (N_40509,N_40178,N_40412);
xnor U40510 (N_40510,N_40456,N_40097);
or U40511 (N_40511,N_40209,N_40455);
and U40512 (N_40512,N_40072,N_40288);
or U40513 (N_40513,N_40357,N_40092);
or U40514 (N_40514,N_40174,N_40336);
or U40515 (N_40515,N_40261,N_40099);
nor U40516 (N_40516,N_40397,N_40290);
or U40517 (N_40517,N_40441,N_40137);
xor U40518 (N_40518,N_40044,N_40101);
and U40519 (N_40519,N_40165,N_40482);
and U40520 (N_40520,N_40319,N_40067);
and U40521 (N_40521,N_40047,N_40138);
nor U40522 (N_40522,N_40338,N_40024);
nor U40523 (N_40523,N_40233,N_40422);
nor U40524 (N_40524,N_40387,N_40184);
nor U40525 (N_40525,N_40027,N_40415);
nand U40526 (N_40526,N_40308,N_40100);
or U40527 (N_40527,N_40170,N_40445);
and U40528 (N_40528,N_40251,N_40121);
nor U40529 (N_40529,N_40452,N_40468);
nor U40530 (N_40530,N_40034,N_40068);
nand U40531 (N_40531,N_40476,N_40407);
xnor U40532 (N_40532,N_40304,N_40351);
or U40533 (N_40533,N_40252,N_40320);
and U40534 (N_40534,N_40048,N_40466);
and U40535 (N_40535,N_40129,N_40194);
nor U40536 (N_40536,N_40454,N_40139);
nand U40537 (N_40537,N_40028,N_40250);
and U40538 (N_40538,N_40461,N_40405);
and U40539 (N_40539,N_40439,N_40009);
or U40540 (N_40540,N_40313,N_40164);
xnor U40541 (N_40541,N_40431,N_40402);
or U40542 (N_40542,N_40172,N_40231);
nor U40543 (N_40543,N_40001,N_40131);
nor U40544 (N_40544,N_40305,N_40041);
nor U40545 (N_40545,N_40065,N_40488);
or U40546 (N_40546,N_40142,N_40136);
xor U40547 (N_40547,N_40260,N_40003);
xor U40548 (N_40548,N_40469,N_40359);
nand U40549 (N_40549,N_40462,N_40085);
or U40550 (N_40550,N_40325,N_40205);
nand U40551 (N_40551,N_40109,N_40303);
and U40552 (N_40552,N_40354,N_40388);
and U40553 (N_40553,N_40273,N_40262);
nor U40554 (N_40554,N_40457,N_40020);
xnor U40555 (N_40555,N_40449,N_40378);
and U40556 (N_40556,N_40426,N_40348);
nor U40557 (N_40557,N_40289,N_40370);
or U40558 (N_40558,N_40298,N_40022);
and U40559 (N_40559,N_40311,N_40398);
nand U40560 (N_40560,N_40343,N_40210);
and U40561 (N_40561,N_40384,N_40106);
nand U40562 (N_40562,N_40277,N_40185);
or U40563 (N_40563,N_40019,N_40372);
nand U40564 (N_40564,N_40366,N_40183);
nand U40565 (N_40565,N_40271,N_40341);
xor U40566 (N_40566,N_40025,N_40151);
and U40567 (N_40567,N_40406,N_40005);
nor U40568 (N_40568,N_40135,N_40429);
and U40569 (N_40569,N_40331,N_40498);
or U40570 (N_40570,N_40073,N_40011);
xnor U40571 (N_40571,N_40224,N_40225);
and U40572 (N_40572,N_40458,N_40226);
xnor U40573 (N_40573,N_40230,N_40435);
or U40574 (N_40574,N_40327,N_40023);
and U40575 (N_40575,N_40291,N_40050);
nor U40576 (N_40576,N_40091,N_40175);
nor U40577 (N_40577,N_40167,N_40247);
or U40578 (N_40578,N_40032,N_40096);
and U40579 (N_40579,N_40453,N_40399);
and U40580 (N_40580,N_40013,N_40212);
or U40581 (N_40581,N_40246,N_40186);
nand U40582 (N_40582,N_40150,N_40293);
or U40583 (N_40583,N_40071,N_40440);
and U40584 (N_40584,N_40401,N_40093);
and U40585 (N_40585,N_40264,N_40054);
nor U40586 (N_40586,N_40064,N_40483);
and U40587 (N_40587,N_40248,N_40083);
or U40588 (N_40588,N_40095,N_40104);
and U40589 (N_40589,N_40021,N_40118);
xor U40590 (N_40590,N_40113,N_40045);
or U40591 (N_40591,N_40000,N_40029);
nand U40592 (N_40592,N_40190,N_40166);
nand U40593 (N_40593,N_40385,N_40408);
xor U40594 (N_40594,N_40227,N_40499);
or U40595 (N_40595,N_40177,N_40254);
nor U40596 (N_40596,N_40160,N_40103);
or U40597 (N_40597,N_40423,N_40344);
or U40598 (N_40598,N_40058,N_40424);
and U40599 (N_40599,N_40031,N_40240);
or U40600 (N_40600,N_40245,N_40496);
nand U40601 (N_40601,N_40014,N_40347);
and U40602 (N_40602,N_40195,N_40187);
nand U40603 (N_40603,N_40446,N_40314);
and U40604 (N_40604,N_40442,N_40259);
or U40605 (N_40605,N_40263,N_40253);
or U40606 (N_40606,N_40006,N_40409);
or U40607 (N_40607,N_40218,N_40464);
nor U40608 (N_40608,N_40215,N_40123);
xnor U40609 (N_40609,N_40272,N_40368);
nor U40610 (N_40610,N_40074,N_40493);
nand U40611 (N_40611,N_40152,N_40102);
and U40612 (N_40612,N_40242,N_40004);
nand U40613 (N_40613,N_40202,N_40244);
nand U40614 (N_40614,N_40081,N_40480);
and U40615 (N_40615,N_40249,N_40299);
nand U40616 (N_40616,N_40278,N_40376);
nor U40617 (N_40617,N_40403,N_40076);
nand U40618 (N_40618,N_40080,N_40030);
nand U40619 (N_40619,N_40168,N_40460);
xnor U40620 (N_40620,N_40459,N_40036);
nor U40621 (N_40621,N_40437,N_40307);
or U40622 (N_40622,N_40116,N_40062);
or U40623 (N_40623,N_40443,N_40265);
or U40624 (N_40624,N_40140,N_40479);
and U40625 (N_40625,N_40395,N_40267);
nor U40626 (N_40626,N_40056,N_40330);
or U40627 (N_40627,N_40478,N_40356);
nand U40628 (N_40628,N_40084,N_40367);
nor U40629 (N_40629,N_40274,N_40176);
nand U40630 (N_40630,N_40127,N_40219);
and U40631 (N_40631,N_40485,N_40410);
nand U40632 (N_40632,N_40199,N_40217);
and U40633 (N_40633,N_40337,N_40352);
nor U40634 (N_40634,N_40444,N_40369);
and U40635 (N_40635,N_40326,N_40494);
and U40636 (N_40636,N_40200,N_40432);
and U40637 (N_40637,N_40179,N_40257);
and U40638 (N_40638,N_40203,N_40196);
nand U40639 (N_40639,N_40171,N_40132);
xor U40640 (N_40640,N_40292,N_40236);
and U40641 (N_40641,N_40365,N_40404);
or U40642 (N_40642,N_40390,N_40420);
and U40643 (N_40643,N_40279,N_40204);
and U40644 (N_40644,N_40329,N_40317);
and U40645 (N_40645,N_40155,N_40018);
nand U40646 (N_40646,N_40037,N_40110);
xnor U40647 (N_40647,N_40427,N_40055);
nand U40648 (N_40648,N_40039,N_40283);
nor U40649 (N_40649,N_40223,N_40382);
and U40650 (N_40650,N_40383,N_40321);
nor U40651 (N_40651,N_40360,N_40222);
nor U40652 (N_40652,N_40294,N_40173);
nand U40653 (N_40653,N_40335,N_40284);
nand U40654 (N_40654,N_40130,N_40216);
xnor U40655 (N_40655,N_40038,N_40470);
and U40656 (N_40656,N_40143,N_40276);
and U40657 (N_40657,N_40375,N_40475);
and U40658 (N_40658,N_40077,N_40323);
xor U40659 (N_40659,N_40381,N_40312);
nand U40660 (N_40660,N_40318,N_40355);
xnor U40661 (N_40661,N_40207,N_40235);
and U40662 (N_40662,N_40211,N_40350);
nand U40663 (N_40663,N_40125,N_40421);
nand U40664 (N_40664,N_40070,N_40489);
and U40665 (N_40665,N_40269,N_40141);
xor U40666 (N_40666,N_40472,N_40002);
and U40667 (N_40667,N_40477,N_40281);
nand U40668 (N_40668,N_40087,N_40391);
nand U40669 (N_40669,N_40474,N_40239);
or U40670 (N_40670,N_40088,N_40287);
nand U40671 (N_40671,N_40094,N_40492);
nor U40672 (N_40672,N_40465,N_40026);
nor U40673 (N_40673,N_40017,N_40069);
nor U40674 (N_40674,N_40238,N_40115);
and U40675 (N_40675,N_40286,N_40414);
xnor U40676 (N_40676,N_40371,N_40149);
and U40677 (N_40677,N_40322,N_40234);
nand U40678 (N_40678,N_40188,N_40053);
nor U40679 (N_40679,N_40316,N_40035);
or U40680 (N_40680,N_40364,N_40214);
or U40681 (N_40681,N_40189,N_40413);
nor U40682 (N_40682,N_40089,N_40066);
or U40683 (N_40683,N_40487,N_40256);
or U40684 (N_40684,N_40363,N_40016);
xnor U40685 (N_40685,N_40430,N_40471);
and U40686 (N_40686,N_40436,N_40208);
nor U40687 (N_40687,N_40148,N_40008);
and U40688 (N_40688,N_40374,N_40417);
nor U40689 (N_40689,N_40154,N_40119);
or U40690 (N_40690,N_40126,N_40057);
and U40691 (N_40691,N_40112,N_40120);
nor U40692 (N_40692,N_40258,N_40147);
nand U40693 (N_40693,N_40270,N_40108);
nand U40694 (N_40694,N_40389,N_40419);
nor U40695 (N_40695,N_40111,N_40243);
nor U40696 (N_40696,N_40051,N_40333);
or U40697 (N_40697,N_40463,N_40161);
xor U40698 (N_40698,N_40297,N_40310);
nand U40699 (N_40699,N_40192,N_40362);
or U40700 (N_40700,N_40124,N_40346);
or U40701 (N_40701,N_40163,N_40345);
nand U40702 (N_40702,N_40467,N_40339);
and U40703 (N_40703,N_40090,N_40153);
or U40704 (N_40704,N_40491,N_40380);
nor U40705 (N_40705,N_40328,N_40114);
and U40706 (N_40706,N_40393,N_40280);
xor U40707 (N_40707,N_40255,N_40232);
xor U40708 (N_40708,N_40144,N_40373);
nand U40709 (N_40709,N_40193,N_40411);
nand U40710 (N_40710,N_40241,N_40349);
nor U40711 (N_40711,N_40146,N_40300);
or U40712 (N_40712,N_40052,N_40334);
or U40713 (N_40713,N_40182,N_40438);
nor U40714 (N_40714,N_40046,N_40158);
nand U40715 (N_40715,N_40162,N_40117);
nor U40716 (N_40716,N_40105,N_40379);
nor U40717 (N_40717,N_40206,N_40340);
or U40718 (N_40718,N_40237,N_40309);
nand U40719 (N_40719,N_40043,N_40007);
nor U40720 (N_40720,N_40306,N_40213);
and U40721 (N_40721,N_40473,N_40266);
or U40722 (N_40722,N_40447,N_40201);
xnor U40723 (N_40723,N_40229,N_40082);
nor U40724 (N_40724,N_40060,N_40015);
and U40725 (N_40725,N_40394,N_40033);
and U40726 (N_40726,N_40157,N_40040);
nand U40727 (N_40727,N_40497,N_40332);
or U40728 (N_40728,N_40145,N_40063);
and U40729 (N_40729,N_40490,N_40450);
and U40730 (N_40730,N_40107,N_40396);
nand U40731 (N_40731,N_40078,N_40434);
nor U40732 (N_40732,N_40128,N_40061);
nand U40733 (N_40733,N_40342,N_40134);
xor U40734 (N_40734,N_40133,N_40268);
or U40735 (N_40735,N_40079,N_40042);
nor U40736 (N_40736,N_40418,N_40169);
or U40737 (N_40737,N_40012,N_40428);
nand U40738 (N_40738,N_40159,N_40416);
and U40739 (N_40739,N_40392,N_40228);
or U40740 (N_40740,N_40285,N_40049);
or U40741 (N_40741,N_40198,N_40377);
or U40742 (N_40742,N_40425,N_40075);
or U40743 (N_40743,N_40086,N_40324);
nor U40744 (N_40744,N_40010,N_40358);
nor U40745 (N_40745,N_40275,N_40495);
nor U40746 (N_40746,N_40433,N_40448);
and U40747 (N_40747,N_40386,N_40191);
nor U40748 (N_40748,N_40221,N_40098);
or U40749 (N_40749,N_40156,N_40481);
nand U40750 (N_40750,N_40069,N_40009);
or U40751 (N_40751,N_40114,N_40406);
or U40752 (N_40752,N_40146,N_40373);
or U40753 (N_40753,N_40081,N_40199);
nand U40754 (N_40754,N_40487,N_40456);
nor U40755 (N_40755,N_40477,N_40210);
xnor U40756 (N_40756,N_40117,N_40218);
and U40757 (N_40757,N_40314,N_40378);
nor U40758 (N_40758,N_40468,N_40211);
nor U40759 (N_40759,N_40297,N_40009);
nand U40760 (N_40760,N_40026,N_40108);
nand U40761 (N_40761,N_40397,N_40036);
and U40762 (N_40762,N_40195,N_40451);
or U40763 (N_40763,N_40282,N_40214);
nor U40764 (N_40764,N_40140,N_40027);
and U40765 (N_40765,N_40052,N_40155);
nor U40766 (N_40766,N_40445,N_40257);
nand U40767 (N_40767,N_40346,N_40059);
nand U40768 (N_40768,N_40389,N_40014);
nand U40769 (N_40769,N_40290,N_40407);
xor U40770 (N_40770,N_40055,N_40141);
and U40771 (N_40771,N_40375,N_40472);
or U40772 (N_40772,N_40369,N_40179);
nor U40773 (N_40773,N_40483,N_40476);
and U40774 (N_40774,N_40269,N_40125);
nand U40775 (N_40775,N_40287,N_40270);
or U40776 (N_40776,N_40478,N_40299);
or U40777 (N_40777,N_40272,N_40024);
or U40778 (N_40778,N_40006,N_40173);
and U40779 (N_40779,N_40282,N_40053);
or U40780 (N_40780,N_40361,N_40499);
xnor U40781 (N_40781,N_40357,N_40361);
and U40782 (N_40782,N_40170,N_40406);
nor U40783 (N_40783,N_40061,N_40073);
nor U40784 (N_40784,N_40433,N_40125);
xor U40785 (N_40785,N_40401,N_40286);
nor U40786 (N_40786,N_40301,N_40250);
xnor U40787 (N_40787,N_40407,N_40198);
or U40788 (N_40788,N_40302,N_40380);
nor U40789 (N_40789,N_40277,N_40311);
or U40790 (N_40790,N_40234,N_40355);
nand U40791 (N_40791,N_40250,N_40437);
or U40792 (N_40792,N_40291,N_40343);
nand U40793 (N_40793,N_40311,N_40207);
xor U40794 (N_40794,N_40440,N_40457);
or U40795 (N_40795,N_40071,N_40428);
nor U40796 (N_40796,N_40208,N_40339);
nor U40797 (N_40797,N_40067,N_40475);
nand U40798 (N_40798,N_40468,N_40256);
nor U40799 (N_40799,N_40409,N_40343);
nor U40800 (N_40800,N_40309,N_40181);
nor U40801 (N_40801,N_40245,N_40412);
or U40802 (N_40802,N_40369,N_40155);
or U40803 (N_40803,N_40487,N_40448);
and U40804 (N_40804,N_40243,N_40063);
nor U40805 (N_40805,N_40257,N_40460);
xnor U40806 (N_40806,N_40191,N_40199);
nand U40807 (N_40807,N_40152,N_40187);
and U40808 (N_40808,N_40458,N_40387);
and U40809 (N_40809,N_40258,N_40150);
nor U40810 (N_40810,N_40343,N_40450);
nand U40811 (N_40811,N_40253,N_40468);
xor U40812 (N_40812,N_40011,N_40084);
nor U40813 (N_40813,N_40315,N_40155);
or U40814 (N_40814,N_40317,N_40367);
nand U40815 (N_40815,N_40442,N_40123);
and U40816 (N_40816,N_40122,N_40246);
or U40817 (N_40817,N_40384,N_40262);
nor U40818 (N_40818,N_40037,N_40264);
or U40819 (N_40819,N_40193,N_40087);
nand U40820 (N_40820,N_40441,N_40476);
or U40821 (N_40821,N_40111,N_40359);
nor U40822 (N_40822,N_40476,N_40215);
and U40823 (N_40823,N_40387,N_40195);
nor U40824 (N_40824,N_40151,N_40241);
nor U40825 (N_40825,N_40317,N_40269);
nor U40826 (N_40826,N_40000,N_40290);
nand U40827 (N_40827,N_40025,N_40432);
or U40828 (N_40828,N_40083,N_40409);
nand U40829 (N_40829,N_40212,N_40423);
nor U40830 (N_40830,N_40069,N_40347);
nand U40831 (N_40831,N_40131,N_40149);
nand U40832 (N_40832,N_40222,N_40247);
xor U40833 (N_40833,N_40357,N_40007);
and U40834 (N_40834,N_40412,N_40413);
xor U40835 (N_40835,N_40200,N_40283);
nand U40836 (N_40836,N_40231,N_40200);
nor U40837 (N_40837,N_40400,N_40086);
and U40838 (N_40838,N_40398,N_40424);
nand U40839 (N_40839,N_40134,N_40438);
nor U40840 (N_40840,N_40084,N_40021);
or U40841 (N_40841,N_40331,N_40438);
nor U40842 (N_40842,N_40363,N_40215);
nor U40843 (N_40843,N_40278,N_40032);
xor U40844 (N_40844,N_40048,N_40045);
nor U40845 (N_40845,N_40216,N_40383);
or U40846 (N_40846,N_40017,N_40425);
nand U40847 (N_40847,N_40352,N_40210);
or U40848 (N_40848,N_40035,N_40322);
nor U40849 (N_40849,N_40299,N_40489);
and U40850 (N_40850,N_40416,N_40214);
nor U40851 (N_40851,N_40467,N_40464);
and U40852 (N_40852,N_40000,N_40215);
nand U40853 (N_40853,N_40136,N_40141);
or U40854 (N_40854,N_40036,N_40222);
nand U40855 (N_40855,N_40276,N_40060);
and U40856 (N_40856,N_40328,N_40370);
and U40857 (N_40857,N_40456,N_40047);
or U40858 (N_40858,N_40203,N_40268);
or U40859 (N_40859,N_40005,N_40022);
or U40860 (N_40860,N_40012,N_40465);
nor U40861 (N_40861,N_40145,N_40263);
xor U40862 (N_40862,N_40426,N_40347);
nand U40863 (N_40863,N_40441,N_40259);
and U40864 (N_40864,N_40233,N_40265);
or U40865 (N_40865,N_40182,N_40319);
xor U40866 (N_40866,N_40329,N_40351);
xor U40867 (N_40867,N_40060,N_40236);
and U40868 (N_40868,N_40138,N_40059);
nand U40869 (N_40869,N_40492,N_40386);
nand U40870 (N_40870,N_40073,N_40453);
nor U40871 (N_40871,N_40388,N_40120);
and U40872 (N_40872,N_40162,N_40197);
and U40873 (N_40873,N_40063,N_40291);
and U40874 (N_40874,N_40269,N_40408);
xnor U40875 (N_40875,N_40366,N_40450);
or U40876 (N_40876,N_40081,N_40031);
xnor U40877 (N_40877,N_40035,N_40053);
xnor U40878 (N_40878,N_40245,N_40499);
and U40879 (N_40879,N_40326,N_40176);
nor U40880 (N_40880,N_40157,N_40144);
nand U40881 (N_40881,N_40086,N_40406);
nor U40882 (N_40882,N_40255,N_40388);
and U40883 (N_40883,N_40304,N_40039);
nor U40884 (N_40884,N_40339,N_40364);
and U40885 (N_40885,N_40391,N_40473);
or U40886 (N_40886,N_40451,N_40081);
nor U40887 (N_40887,N_40039,N_40145);
and U40888 (N_40888,N_40325,N_40374);
nor U40889 (N_40889,N_40181,N_40147);
xnor U40890 (N_40890,N_40016,N_40300);
xnor U40891 (N_40891,N_40078,N_40234);
nor U40892 (N_40892,N_40368,N_40134);
or U40893 (N_40893,N_40172,N_40179);
nor U40894 (N_40894,N_40109,N_40036);
nor U40895 (N_40895,N_40281,N_40427);
or U40896 (N_40896,N_40165,N_40282);
or U40897 (N_40897,N_40384,N_40136);
and U40898 (N_40898,N_40498,N_40155);
xor U40899 (N_40899,N_40235,N_40159);
and U40900 (N_40900,N_40340,N_40014);
nand U40901 (N_40901,N_40499,N_40237);
nand U40902 (N_40902,N_40439,N_40226);
nand U40903 (N_40903,N_40234,N_40140);
xor U40904 (N_40904,N_40265,N_40121);
nand U40905 (N_40905,N_40479,N_40069);
nor U40906 (N_40906,N_40144,N_40422);
nor U40907 (N_40907,N_40178,N_40000);
or U40908 (N_40908,N_40300,N_40381);
and U40909 (N_40909,N_40197,N_40055);
or U40910 (N_40910,N_40371,N_40023);
nand U40911 (N_40911,N_40458,N_40217);
and U40912 (N_40912,N_40417,N_40096);
nand U40913 (N_40913,N_40427,N_40402);
nand U40914 (N_40914,N_40143,N_40345);
nand U40915 (N_40915,N_40075,N_40428);
or U40916 (N_40916,N_40291,N_40130);
nor U40917 (N_40917,N_40393,N_40479);
nand U40918 (N_40918,N_40439,N_40026);
and U40919 (N_40919,N_40376,N_40196);
or U40920 (N_40920,N_40442,N_40132);
and U40921 (N_40921,N_40089,N_40379);
and U40922 (N_40922,N_40105,N_40280);
nor U40923 (N_40923,N_40464,N_40056);
nand U40924 (N_40924,N_40017,N_40181);
or U40925 (N_40925,N_40143,N_40013);
nand U40926 (N_40926,N_40143,N_40108);
xor U40927 (N_40927,N_40297,N_40124);
and U40928 (N_40928,N_40441,N_40036);
and U40929 (N_40929,N_40379,N_40431);
nand U40930 (N_40930,N_40082,N_40409);
or U40931 (N_40931,N_40372,N_40444);
xnor U40932 (N_40932,N_40130,N_40051);
nand U40933 (N_40933,N_40050,N_40434);
and U40934 (N_40934,N_40215,N_40033);
nor U40935 (N_40935,N_40245,N_40421);
or U40936 (N_40936,N_40257,N_40496);
or U40937 (N_40937,N_40295,N_40405);
and U40938 (N_40938,N_40360,N_40405);
and U40939 (N_40939,N_40437,N_40465);
and U40940 (N_40940,N_40022,N_40094);
or U40941 (N_40941,N_40313,N_40197);
or U40942 (N_40942,N_40418,N_40457);
and U40943 (N_40943,N_40161,N_40131);
xor U40944 (N_40944,N_40018,N_40086);
nand U40945 (N_40945,N_40014,N_40062);
or U40946 (N_40946,N_40375,N_40354);
xor U40947 (N_40947,N_40230,N_40077);
nand U40948 (N_40948,N_40156,N_40202);
xor U40949 (N_40949,N_40010,N_40215);
and U40950 (N_40950,N_40301,N_40092);
nand U40951 (N_40951,N_40339,N_40151);
xnor U40952 (N_40952,N_40314,N_40445);
nand U40953 (N_40953,N_40477,N_40238);
or U40954 (N_40954,N_40059,N_40212);
nor U40955 (N_40955,N_40069,N_40160);
and U40956 (N_40956,N_40058,N_40437);
or U40957 (N_40957,N_40356,N_40313);
nor U40958 (N_40958,N_40379,N_40004);
and U40959 (N_40959,N_40496,N_40453);
nor U40960 (N_40960,N_40209,N_40269);
or U40961 (N_40961,N_40485,N_40052);
nor U40962 (N_40962,N_40029,N_40045);
nor U40963 (N_40963,N_40048,N_40443);
nand U40964 (N_40964,N_40230,N_40209);
or U40965 (N_40965,N_40178,N_40261);
nand U40966 (N_40966,N_40402,N_40403);
xor U40967 (N_40967,N_40064,N_40268);
nand U40968 (N_40968,N_40046,N_40283);
or U40969 (N_40969,N_40486,N_40089);
nand U40970 (N_40970,N_40248,N_40459);
or U40971 (N_40971,N_40134,N_40218);
nand U40972 (N_40972,N_40181,N_40303);
and U40973 (N_40973,N_40424,N_40074);
and U40974 (N_40974,N_40083,N_40316);
or U40975 (N_40975,N_40157,N_40153);
and U40976 (N_40976,N_40179,N_40298);
and U40977 (N_40977,N_40416,N_40464);
and U40978 (N_40978,N_40138,N_40362);
or U40979 (N_40979,N_40424,N_40375);
or U40980 (N_40980,N_40238,N_40480);
and U40981 (N_40981,N_40270,N_40173);
or U40982 (N_40982,N_40095,N_40402);
nand U40983 (N_40983,N_40044,N_40434);
nand U40984 (N_40984,N_40327,N_40084);
and U40985 (N_40985,N_40124,N_40018);
or U40986 (N_40986,N_40279,N_40430);
and U40987 (N_40987,N_40139,N_40222);
or U40988 (N_40988,N_40457,N_40208);
and U40989 (N_40989,N_40111,N_40286);
nand U40990 (N_40990,N_40370,N_40030);
nor U40991 (N_40991,N_40431,N_40403);
and U40992 (N_40992,N_40244,N_40389);
or U40993 (N_40993,N_40315,N_40072);
and U40994 (N_40994,N_40335,N_40394);
nand U40995 (N_40995,N_40262,N_40161);
nand U40996 (N_40996,N_40426,N_40280);
nor U40997 (N_40997,N_40425,N_40263);
or U40998 (N_40998,N_40323,N_40128);
or U40999 (N_40999,N_40392,N_40277);
and U41000 (N_41000,N_40629,N_40501);
xor U41001 (N_41001,N_40849,N_40766);
nand U41002 (N_41002,N_40974,N_40738);
xnor U41003 (N_41003,N_40533,N_40746);
or U41004 (N_41004,N_40751,N_40511);
and U41005 (N_41005,N_40556,N_40702);
nand U41006 (N_41006,N_40528,N_40730);
or U41007 (N_41007,N_40805,N_40674);
nand U41008 (N_41008,N_40548,N_40837);
nand U41009 (N_41009,N_40831,N_40981);
and U41010 (N_41010,N_40723,N_40506);
nor U41011 (N_41011,N_40543,N_40546);
nor U41012 (N_41012,N_40503,N_40798);
nor U41013 (N_41013,N_40948,N_40750);
nor U41014 (N_41014,N_40597,N_40735);
nor U41015 (N_41015,N_40645,N_40971);
or U41016 (N_41016,N_40579,N_40964);
and U41017 (N_41017,N_40539,N_40870);
nor U41018 (N_41018,N_40859,N_40860);
nor U41019 (N_41019,N_40532,N_40536);
and U41020 (N_41020,N_40646,N_40973);
nand U41021 (N_41021,N_40940,N_40567);
and U41022 (N_41022,N_40524,N_40998);
nor U41023 (N_41023,N_40624,N_40685);
or U41024 (N_41024,N_40634,N_40967);
and U41025 (N_41025,N_40801,N_40510);
xor U41026 (N_41026,N_40720,N_40578);
nand U41027 (N_41027,N_40784,N_40789);
nor U41028 (N_41028,N_40507,N_40635);
or U41029 (N_41029,N_40797,N_40905);
xor U41030 (N_41030,N_40976,N_40700);
and U41031 (N_41031,N_40790,N_40653);
nand U41032 (N_41032,N_40871,N_40892);
xnor U41033 (N_41033,N_40935,N_40690);
nor U41034 (N_41034,N_40911,N_40979);
xor U41035 (N_41035,N_40654,N_40897);
nor U41036 (N_41036,N_40584,N_40534);
or U41037 (N_41037,N_40846,N_40963);
nor U41038 (N_41038,N_40585,N_40583);
and U41039 (N_41039,N_40876,N_40555);
or U41040 (N_41040,N_40682,N_40816);
nand U41041 (N_41041,N_40669,N_40921);
nand U41042 (N_41042,N_40713,N_40862);
xor U41043 (N_41043,N_40693,N_40777);
or U41044 (N_41044,N_40626,N_40522);
nand U41045 (N_41045,N_40800,N_40754);
nand U41046 (N_41046,N_40850,N_40719);
nor U41047 (N_41047,N_40678,N_40686);
xor U41048 (N_41048,N_40665,N_40531);
or U41049 (N_41049,N_40550,N_40740);
and U41050 (N_41050,N_40745,N_40553);
xnor U41051 (N_41051,N_40615,N_40959);
and U41052 (N_41052,N_40642,N_40625);
xor U41053 (N_41053,N_40866,N_40826);
nand U41054 (N_41054,N_40612,N_40771);
nor U41055 (N_41055,N_40773,N_40722);
and U41056 (N_41056,N_40966,N_40756);
nand U41057 (N_41057,N_40513,N_40960);
xor U41058 (N_41058,N_40611,N_40622);
nand U41059 (N_41059,N_40558,N_40933);
xnor U41060 (N_41060,N_40747,N_40934);
nand U41061 (N_41061,N_40881,N_40944);
nand U41062 (N_41062,N_40605,N_40736);
and U41063 (N_41063,N_40868,N_40996);
xor U41064 (N_41064,N_40576,N_40643);
nor U41065 (N_41065,N_40886,N_40614);
xor U41066 (N_41066,N_40708,N_40610);
and U41067 (N_41067,N_40600,N_40676);
and U41068 (N_41068,N_40559,N_40759);
nor U41069 (N_41069,N_40637,N_40803);
or U41070 (N_41070,N_40987,N_40995);
or U41071 (N_41071,N_40835,N_40982);
and U41072 (N_41072,N_40906,N_40950);
or U41073 (N_41073,N_40521,N_40814);
and U41074 (N_41074,N_40999,N_40989);
and U41075 (N_41075,N_40591,N_40565);
or U41076 (N_41076,N_40604,N_40581);
nand U41077 (N_41077,N_40658,N_40596);
nor U41078 (N_41078,N_40648,N_40887);
nor U41079 (N_41079,N_40727,N_40725);
xor U41080 (N_41080,N_40962,N_40775);
or U41081 (N_41081,N_40679,N_40840);
nor U41082 (N_41082,N_40502,N_40609);
or U41083 (N_41083,N_40752,N_40717);
or U41084 (N_41084,N_40903,N_40785);
nand U41085 (N_41085,N_40662,N_40660);
nor U41086 (N_41086,N_40841,N_40592);
nor U41087 (N_41087,N_40793,N_40761);
and U41088 (N_41088,N_40970,N_40913);
xor U41089 (N_41089,N_40656,N_40704);
or U41090 (N_41090,N_40683,N_40744);
and U41091 (N_41091,N_40972,N_40701);
and U41092 (N_41092,N_40885,N_40640);
nand U41093 (N_41093,N_40621,N_40542);
or U41094 (N_41094,N_40997,N_40993);
nor U41095 (N_41095,N_40807,N_40724);
and U41096 (N_41096,N_40821,N_40957);
and U41097 (N_41097,N_40762,N_40763);
nor U41098 (N_41098,N_40829,N_40875);
nor U41099 (N_41099,N_40541,N_40666);
nand U41100 (N_41100,N_40882,N_40599);
nand U41101 (N_41101,N_40895,N_40547);
or U41102 (N_41102,N_40718,N_40845);
nand U41103 (N_41103,N_40606,N_40619);
nor U41104 (N_41104,N_40770,N_40842);
or U41105 (N_41105,N_40516,N_40922);
nand U41106 (N_41106,N_40928,N_40650);
nor U41107 (N_41107,N_40817,N_40667);
nor U41108 (N_41108,N_40852,N_40857);
nor U41109 (N_41109,N_40677,N_40582);
nand U41110 (N_41110,N_40739,N_40568);
nand U41111 (N_41111,N_40824,N_40694);
and U41112 (N_41112,N_40737,N_40819);
nand U41113 (N_41113,N_40917,N_40564);
and U41114 (N_41114,N_40574,N_40969);
nor U41115 (N_41115,N_40986,N_40809);
nor U41116 (N_41116,N_40937,N_40909);
nand U41117 (N_41117,N_40955,N_40748);
nor U41118 (N_41118,N_40823,N_40782);
nand U41119 (N_41119,N_40799,N_40743);
nor U41120 (N_41120,N_40525,N_40673);
xor U41121 (N_41121,N_40519,N_40710);
nand U41122 (N_41122,N_40529,N_40815);
nand U41123 (N_41123,N_40791,N_40898);
and U41124 (N_41124,N_40900,N_40569);
nand U41125 (N_41125,N_40983,N_40830);
nand U41126 (N_41126,N_40779,N_40661);
nand U41127 (N_41127,N_40869,N_40958);
or U41128 (N_41128,N_40781,N_40883);
xnor U41129 (N_41129,N_40838,N_40680);
nor U41130 (N_41130,N_40668,N_40908);
nand U41131 (N_41131,N_40716,N_40517);
nor U41132 (N_41132,N_40924,N_40537);
and U41133 (N_41133,N_40570,N_40732);
or U41134 (N_41134,N_40623,N_40627);
nand U41135 (N_41135,N_40602,N_40872);
nand U41136 (N_41136,N_40729,N_40899);
and U41137 (N_41137,N_40956,N_40832);
and U41138 (N_41138,N_40926,N_40863);
nand U41139 (N_41139,N_40749,N_40504);
nor U41140 (N_41140,N_40500,N_40764);
and U41141 (N_41141,N_40776,N_40985);
or U41142 (N_41142,N_40527,N_40616);
or U41143 (N_41143,N_40706,N_40918);
or U41144 (N_41144,N_40879,N_40684);
nand U41145 (N_41145,N_40633,N_40925);
nand U41146 (N_41146,N_40698,N_40889);
nand U41147 (N_41147,N_40540,N_40632);
or U41148 (N_41148,N_40772,N_40721);
nor U41149 (N_41149,N_40932,N_40557);
nor U41150 (N_41150,N_40827,N_40949);
and U41151 (N_41151,N_40641,N_40607);
or U41152 (N_41152,N_40587,N_40795);
xnor U41153 (N_41153,N_40994,N_40663);
xor U41154 (N_41154,N_40590,N_40589);
and U41155 (N_41155,N_40984,N_40545);
nor U41156 (N_41156,N_40755,N_40544);
or U41157 (N_41157,N_40699,N_40774);
nor U41158 (N_41158,N_40808,N_40711);
and U41159 (N_41159,N_40880,N_40915);
and U41160 (N_41160,N_40707,N_40595);
nand U41161 (N_41161,N_40705,N_40952);
nor U41162 (N_41162,N_40520,N_40657);
nor U41163 (N_41163,N_40855,N_40695);
nor U41164 (N_41164,N_40728,N_40851);
nand U41165 (N_41165,N_40977,N_40767);
nand U41166 (N_41166,N_40509,N_40647);
nor U41167 (N_41167,N_40515,N_40874);
nor U41168 (N_41168,N_40907,N_40936);
and U41169 (N_41169,N_40802,N_40820);
or U41170 (N_41170,N_40742,N_40783);
xor U41171 (N_41171,N_40988,N_40942);
nand U41172 (N_41172,N_40618,N_40709);
and U41173 (N_41173,N_40843,N_40978);
nor U41174 (N_41174,N_40526,N_40804);
and U41175 (N_41175,N_40914,N_40975);
nor U41176 (N_41176,N_40636,N_40577);
nand U41177 (N_41177,N_40562,N_40786);
and U41178 (N_41178,N_40916,N_40961);
nand U41179 (N_41179,N_40549,N_40954);
nand U41180 (N_41180,N_40794,N_40649);
or U41181 (N_41181,N_40638,N_40947);
and U41182 (N_41182,N_40965,N_40692);
or U41183 (N_41183,N_40884,N_40630);
nor U41184 (N_41184,N_40873,N_40733);
nor U41185 (N_41185,N_40670,N_40980);
nand U41186 (N_41186,N_40644,N_40938);
and U41187 (N_41187,N_40655,N_40848);
and U41188 (N_41188,N_40941,N_40603);
nor U41189 (N_41189,N_40806,N_40768);
nand U41190 (N_41190,N_40566,N_40672);
xor U41191 (N_41191,N_40575,N_40505);
and U41192 (N_41192,N_40813,N_40811);
xnor U41193 (N_41193,N_40931,N_40757);
nand U41194 (N_41194,N_40580,N_40847);
nor U41195 (N_41195,N_40572,N_40968);
nand U41196 (N_41196,N_40758,N_40586);
or U41197 (N_41197,N_40731,N_40514);
or U41198 (N_41198,N_40760,N_40551);
and U41199 (N_41199,N_40778,N_40671);
or U41200 (N_41200,N_40910,N_40681);
xnor U41201 (N_41201,N_40571,N_40943);
nand U41202 (N_41202,N_40792,N_40687);
and U41203 (N_41203,N_40780,N_40594);
or U41204 (N_41204,N_40864,N_40839);
nor U41205 (N_41205,N_40825,N_40920);
and U41206 (N_41206,N_40788,N_40834);
nor U41207 (N_41207,N_40856,N_40535);
nand U41208 (N_41208,N_40769,N_40664);
nor U41209 (N_41209,N_40812,N_40753);
and U41210 (N_41210,N_40854,N_40512);
nor U41211 (N_41211,N_40990,N_40896);
or U41212 (N_41212,N_40691,N_40919);
or U41213 (N_41213,N_40563,N_40741);
nand U41214 (N_41214,N_40844,N_40891);
xnor U41215 (N_41215,N_40893,N_40828);
xnor U41216 (N_41216,N_40715,N_40538);
nand U41217 (N_41217,N_40675,N_40939);
nor U41218 (N_41218,N_40890,N_40508);
nor U41219 (N_41219,N_40523,N_40552);
xnor U41220 (N_41220,N_40639,N_40946);
and U41221 (N_41221,N_40588,N_40651);
nor U41222 (N_41222,N_40601,N_40518);
nand U41223 (N_41223,N_40912,N_40894);
nor U41224 (N_41224,N_40593,N_40712);
nor U41225 (N_41225,N_40923,N_40878);
and U41226 (N_41226,N_40554,N_40530);
and U41227 (N_41227,N_40929,N_40810);
or U41228 (N_41228,N_40697,N_40689);
nor U41229 (N_41229,N_40608,N_40688);
nand U41230 (N_41230,N_40902,N_40945);
nand U41231 (N_41231,N_40927,N_40865);
nand U41232 (N_41232,N_40858,N_40901);
and U41233 (N_41233,N_40696,N_40888);
nor U41234 (N_41234,N_40867,N_40714);
nor U41235 (N_41235,N_40861,N_40822);
nor U41236 (N_41236,N_40726,N_40951);
or U41237 (N_41237,N_40628,N_40734);
nor U41238 (N_41238,N_40631,N_40836);
and U41239 (N_41239,N_40613,N_40617);
and U41240 (N_41240,N_40992,N_40765);
or U41241 (N_41241,N_40659,N_40598);
nand U41242 (N_41242,N_40796,N_40787);
and U41243 (N_41243,N_40877,N_40573);
xnor U41244 (N_41244,N_40652,N_40991);
and U41245 (N_41245,N_40703,N_40904);
and U41246 (N_41246,N_40953,N_40853);
and U41247 (N_41247,N_40561,N_40560);
nand U41248 (N_41248,N_40930,N_40818);
nor U41249 (N_41249,N_40620,N_40833);
nand U41250 (N_41250,N_40754,N_40583);
or U41251 (N_41251,N_40680,N_40936);
or U41252 (N_41252,N_40843,N_40826);
or U41253 (N_41253,N_40831,N_40681);
or U41254 (N_41254,N_40674,N_40538);
or U41255 (N_41255,N_40515,N_40565);
or U41256 (N_41256,N_40507,N_40645);
and U41257 (N_41257,N_40850,N_40737);
xnor U41258 (N_41258,N_40610,N_40730);
nor U41259 (N_41259,N_40809,N_40764);
xnor U41260 (N_41260,N_40591,N_40632);
nor U41261 (N_41261,N_40543,N_40769);
or U41262 (N_41262,N_40900,N_40947);
nor U41263 (N_41263,N_40808,N_40930);
nor U41264 (N_41264,N_40747,N_40632);
or U41265 (N_41265,N_40831,N_40593);
and U41266 (N_41266,N_40825,N_40733);
nand U41267 (N_41267,N_40822,N_40754);
or U41268 (N_41268,N_40674,N_40693);
nand U41269 (N_41269,N_40851,N_40538);
xor U41270 (N_41270,N_40621,N_40879);
nand U41271 (N_41271,N_40905,N_40846);
xor U41272 (N_41272,N_40799,N_40638);
nand U41273 (N_41273,N_40510,N_40550);
and U41274 (N_41274,N_40818,N_40965);
or U41275 (N_41275,N_40692,N_40718);
nand U41276 (N_41276,N_40836,N_40816);
xnor U41277 (N_41277,N_40711,N_40688);
nor U41278 (N_41278,N_40617,N_40905);
and U41279 (N_41279,N_40939,N_40950);
nor U41280 (N_41280,N_40671,N_40942);
nand U41281 (N_41281,N_40629,N_40606);
and U41282 (N_41282,N_40614,N_40800);
nand U41283 (N_41283,N_40920,N_40925);
or U41284 (N_41284,N_40924,N_40900);
and U41285 (N_41285,N_40958,N_40814);
or U41286 (N_41286,N_40535,N_40571);
nor U41287 (N_41287,N_40943,N_40911);
nand U41288 (N_41288,N_40696,N_40601);
nand U41289 (N_41289,N_40572,N_40673);
xnor U41290 (N_41290,N_40522,N_40866);
nand U41291 (N_41291,N_40513,N_40899);
nand U41292 (N_41292,N_40854,N_40799);
nand U41293 (N_41293,N_40739,N_40553);
nor U41294 (N_41294,N_40955,N_40652);
nand U41295 (N_41295,N_40849,N_40654);
xor U41296 (N_41296,N_40539,N_40956);
nand U41297 (N_41297,N_40808,N_40541);
or U41298 (N_41298,N_40970,N_40980);
and U41299 (N_41299,N_40510,N_40788);
nor U41300 (N_41300,N_40501,N_40757);
nand U41301 (N_41301,N_40999,N_40506);
nor U41302 (N_41302,N_40619,N_40921);
nor U41303 (N_41303,N_40649,N_40663);
nor U41304 (N_41304,N_40985,N_40591);
and U41305 (N_41305,N_40615,N_40794);
or U41306 (N_41306,N_40964,N_40952);
or U41307 (N_41307,N_40707,N_40531);
nand U41308 (N_41308,N_40714,N_40643);
nand U41309 (N_41309,N_40525,N_40918);
nand U41310 (N_41310,N_40566,N_40877);
and U41311 (N_41311,N_40815,N_40862);
nor U41312 (N_41312,N_40816,N_40837);
xor U41313 (N_41313,N_40630,N_40710);
or U41314 (N_41314,N_40807,N_40595);
xor U41315 (N_41315,N_40782,N_40721);
nand U41316 (N_41316,N_40774,N_40794);
nor U41317 (N_41317,N_40555,N_40953);
nor U41318 (N_41318,N_40644,N_40575);
and U41319 (N_41319,N_40717,N_40880);
nor U41320 (N_41320,N_40544,N_40969);
or U41321 (N_41321,N_40812,N_40959);
and U41322 (N_41322,N_40802,N_40939);
nand U41323 (N_41323,N_40859,N_40513);
and U41324 (N_41324,N_40818,N_40831);
nand U41325 (N_41325,N_40931,N_40803);
and U41326 (N_41326,N_40606,N_40871);
xor U41327 (N_41327,N_40841,N_40501);
nor U41328 (N_41328,N_40735,N_40583);
and U41329 (N_41329,N_40553,N_40927);
nor U41330 (N_41330,N_40831,N_40767);
xnor U41331 (N_41331,N_40691,N_40834);
nor U41332 (N_41332,N_40871,N_40998);
nor U41333 (N_41333,N_40690,N_40602);
or U41334 (N_41334,N_40763,N_40941);
and U41335 (N_41335,N_40658,N_40627);
xor U41336 (N_41336,N_40974,N_40650);
nand U41337 (N_41337,N_40619,N_40952);
nor U41338 (N_41338,N_40650,N_40689);
or U41339 (N_41339,N_40984,N_40840);
or U41340 (N_41340,N_40843,N_40934);
or U41341 (N_41341,N_40742,N_40612);
nor U41342 (N_41342,N_40900,N_40656);
nand U41343 (N_41343,N_40771,N_40966);
nand U41344 (N_41344,N_40935,N_40819);
nor U41345 (N_41345,N_40767,N_40722);
nor U41346 (N_41346,N_40572,N_40781);
nor U41347 (N_41347,N_40580,N_40747);
xnor U41348 (N_41348,N_40831,N_40752);
nand U41349 (N_41349,N_40644,N_40511);
or U41350 (N_41350,N_40542,N_40924);
or U41351 (N_41351,N_40804,N_40596);
nand U41352 (N_41352,N_40766,N_40871);
nand U41353 (N_41353,N_40535,N_40564);
or U41354 (N_41354,N_40890,N_40616);
or U41355 (N_41355,N_40710,N_40890);
nand U41356 (N_41356,N_40722,N_40985);
nand U41357 (N_41357,N_40883,N_40719);
nand U41358 (N_41358,N_40990,N_40976);
nand U41359 (N_41359,N_40937,N_40811);
nand U41360 (N_41360,N_40688,N_40812);
nand U41361 (N_41361,N_40729,N_40672);
or U41362 (N_41362,N_40633,N_40832);
nor U41363 (N_41363,N_40963,N_40625);
nor U41364 (N_41364,N_40756,N_40702);
and U41365 (N_41365,N_40657,N_40993);
nand U41366 (N_41366,N_40602,N_40641);
nor U41367 (N_41367,N_40982,N_40781);
nor U41368 (N_41368,N_40651,N_40697);
xnor U41369 (N_41369,N_40647,N_40545);
and U41370 (N_41370,N_40969,N_40529);
or U41371 (N_41371,N_40901,N_40650);
nand U41372 (N_41372,N_40644,N_40723);
xor U41373 (N_41373,N_40536,N_40547);
nor U41374 (N_41374,N_40524,N_40520);
nor U41375 (N_41375,N_40894,N_40997);
and U41376 (N_41376,N_40551,N_40591);
or U41377 (N_41377,N_40853,N_40623);
and U41378 (N_41378,N_40893,N_40694);
nand U41379 (N_41379,N_40723,N_40892);
and U41380 (N_41380,N_40734,N_40924);
nor U41381 (N_41381,N_40633,N_40621);
nand U41382 (N_41382,N_40647,N_40751);
xor U41383 (N_41383,N_40907,N_40652);
nor U41384 (N_41384,N_40620,N_40786);
or U41385 (N_41385,N_40712,N_40855);
nor U41386 (N_41386,N_40747,N_40723);
and U41387 (N_41387,N_40813,N_40584);
xnor U41388 (N_41388,N_40931,N_40989);
xor U41389 (N_41389,N_40518,N_40701);
nand U41390 (N_41390,N_40613,N_40606);
nor U41391 (N_41391,N_40679,N_40663);
and U41392 (N_41392,N_40990,N_40507);
and U41393 (N_41393,N_40591,N_40719);
and U41394 (N_41394,N_40992,N_40824);
xor U41395 (N_41395,N_40509,N_40700);
and U41396 (N_41396,N_40806,N_40726);
or U41397 (N_41397,N_40571,N_40965);
or U41398 (N_41398,N_40588,N_40615);
or U41399 (N_41399,N_40883,N_40785);
or U41400 (N_41400,N_40720,N_40505);
nand U41401 (N_41401,N_40837,N_40972);
or U41402 (N_41402,N_40760,N_40593);
and U41403 (N_41403,N_40966,N_40588);
nand U41404 (N_41404,N_40861,N_40770);
and U41405 (N_41405,N_40659,N_40718);
and U41406 (N_41406,N_40665,N_40887);
or U41407 (N_41407,N_40777,N_40605);
and U41408 (N_41408,N_40663,N_40523);
or U41409 (N_41409,N_40685,N_40817);
or U41410 (N_41410,N_40504,N_40924);
nor U41411 (N_41411,N_40953,N_40833);
or U41412 (N_41412,N_40771,N_40881);
or U41413 (N_41413,N_40709,N_40866);
nand U41414 (N_41414,N_40579,N_40551);
or U41415 (N_41415,N_40812,N_40903);
and U41416 (N_41416,N_40765,N_40788);
nor U41417 (N_41417,N_40670,N_40768);
nor U41418 (N_41418,N_40865,N_40941);
or U41419 (N_41419,N_40924,N_40708);
and U41420 (N_41420,N_40612,N_40630);
nand U41421 (N_41421,N_40555,N_40829);
and U41422 (N_41422,N_40689,N_40546);
nand U41423 (N_41423,N_40930,N_40906);
or U41424 (N_41424,N_40821,N_40694);
and U41425 (N_41425,N_40985,N_40830);
and U41426 (N_41426,N_40722,N_40945);
nand U41427 (N_41427,N_40915,N_40585);
xnor U41428 (N_41428,N_40863,N_40743);
and U41429 (N_41429,N_40737,N_40985);
and U41430 (N_41430,N_40733,N_40623);
nor U41431 (N_41431,N_40913,N_40603);
nor U41432 (N_41432,N_40912,N_40838);
or U41433 (N_41433,N_40996,N_40821);
or U41434 (N_41434,N_40975,N_40614);
and U41435 (N_41435,N_40766,N_40708);
nor U41436 (N_41436,N_40957,N_40642);
nor U41437 (N_41437,N_40890,N_40681);
nand U41438 (N_41438,N_40556,N_40596);
nand U41439 (N_41439,N_40882,N_40532);
nand U41440 (N_41440,N_40969,N_40981);
xnor U41441 (N_41441,N_40652,N_40936);
or U41442 (N_41442,N_40961,N_40816);
xnor U41443 (N_41443,N_40849,N_40770);
or U41444 (N_41444,N_40541,N_40645);
or U41445 (N_41445,N_40778,N_40849);
and U41446 (N_41446,N_40671,N_40997);
nand U41447 (N_41447,N_40986,N_40824);
and U41448 (N_41448,N_40782,N_40917);
and U41449 (N_41449,N_40842,N_40974);
or U41450 (N_41450,N_40757,N_40669);
xor U41451 (N_41451,N_40810,N_40504);
nor U41452 (N_41452,N_40790,N_40904);
nand U41453 (N_41453,N_40645,N_40912);
and U41454 (N_41454,N_40812,N_40511);
and U41455 (N_41455,N_40689,N_40969);
and U41456 (N_41456,N_40863,N_40924);
xnor U41457 (N_41457,N_40503,N_40595);
nor U41458 (N_41458,N_40541,N_40529);
nor U41459 (N_41459,N_40585,N_40667);
or U41460 (N_41460,N_40529,N_40854);
nand U41461 (N_41461,N_40650,N_40970);
nor U41462 (N_41462,N_40877,N_40988);
nor U41463 (N_41463,N_40743,N_40724);
and U41464 (N_41464,N_40759,N_40858);
nor U41465 (N_41465,N_40796,N_40644);
nand U41466 (N_41466,N_40740,N_40544);
and U41467 (N_41467,N_40835,N_40744);
or U41468 (N_41468,N_40723,N_40626);
nor U41469 (N_41469,N_40968,N_40600);
or U41470 (N_41470,N_40781,N_40504);
xor U41471 (N_41471,N_40793,N_40833);
nand U41472 (N_41472,N_40996,N_40732);
nor U41473 (N_41473,N_40930,N_40585);
xor U41474 (N_41474,N_40561,N_40564);
nor U41475 (N_41475,N_40614,N_40551);
or U41476 (N_41476,N_40907,N_40638);
xnor U41477 (N_41477,N_40671,N_40524);
nand U41478 (N_41478,N_40513,N_40612);
nor U41479 (N_41479,N_40930,N_40699);
nor U41480 (N_41480,N_40826,N_40716);
nor U41481 (N_41481,N_40527,N_40659);
and U41482 (N_41482,N_40648,N_40602);
or U41483 (N_41483,N_40666,N_40822);
nand U41484 (N_41484,N_40748,N_40614);
or U41485 (N_41485,N_40680,N_40731);
xnor U41486 (N_41486,N_40563,N_40967);
xnor U41487 (N_41487,N_40786,N_40899);
nor U41488 (N_41488,N_40543,N_40656);
nor U41489 (N_41489,N_40618,N_40629);
and U41490 (N_41490,N_40638,N_40860);
nand U41491 (N_41491,N_40974,N_40625);
or U41492 (N_41492,N_40813,N_40581);
nor U41493 (N_41493,N_40533,N_40790);
or U41494 (N_41494,N_40619,N_40820);
nand U41495 (N_41495,N_40635,N_40989);
xnor U41496 (N_41496,N_40978,N_40936);
or U41497 (N_41497,N_40549,N_40836);
nor U41498 (N_41498,N_40911,N_40956);
or U41499 (N_41499,N_40504,N_40797);
and U41500 (N_41500,N_41408,N_41335);
nand U41501 (N_41501,N_41181,N_41109);
and U41502 (N_41502,N_41203,N_41034);
and U41503 (N_41503,N_41345,N_41371);
xnor U41504 (N_41504,N_41451,N_41325);
nor U41505 (N_41505,N_41274,N_41063);
nor U41506 (N_41506,N_41067,N_41084);
nor U41507 (N_41507,N_41483,N_41187);
nand U41508 (N_41508,N_41218,N_41173);
and U41509 (N_41509,N_41272,N_41008);
nor U41510 (N_41510,N_41031,N_41390);
and U41511 (N_41511,N_41275,N_41389);
xor U41512 (N_41512,N_41421,N_41267);
xnor U41513 (N_41513,N_41152,N_41347);
xor U41514 (N_41514,N_41130,N_41230);
or U41515 (N_41515,N_41290,N_41001);
and U41516 (N_41516,N_41201,N_41299);
and U41517 (N_41517,N_41324,N_41418);
nand U41518 (N_41518,N_41160,N_41050);
and U41519 (N_41519,N_41029,N_41461);
nor U41520 (N_41520,N_41204,N_41348);
nor U41521 (N_41521,N_41178,N_41023);
or U41522 (N_41522,N_41256,N_41159);
nand U41523 (N_41523,N_41142,N_41400);
xor U41524 (N_41524,N_41234,N_41077);
nor U41525 (N_41525,N_41409,N_41055);
nor U41526 (N_41526,N_41238,N_41165);
and U41527 (N_41527,N_41496,N_41355);
nand U41528 (N_41528,N_41132,N_41472);
nand U41529 (N_41529,N_41303,N_41412);
nor U41530 (N_41530,N_41378,N_41396);
nand U41531 (N_41531,N_41103,N_41089);
or U41532 (N_41532,N_41148,N_41397);
nor U41533 (N_41533,N_41364,N_41269);
or U41534 (N_41534,N_41490,N_41424);
and U41535 (N_41535,N_41054,N_41282);
or U41536 (N_41536,N_41015,N_41011);
and U41537 (N_41537,N_41014,N_41079);
nor U41538 (N_41538,N_41338,N_41010);
or U41539 (N_41539,N_41381,N_41155);
and U41540 (N_41540,N_41266,N_41487);
and U41541 (N_41541,N_41158,N_41447);
nand U41542 (N_41542,N_41352,N_41175);
xor U41543 (N_41543,N_41006,N_41288);
and U41544 (N_41544,N_41351,N_41313);
nand U41545 (N_41545,N_41212,N_41420);
nand U41546 (N_41546,N_41164,N_41395);
nor U41547 (N_41547,N_41383,N_41277);
or U41548 (N_41548,N_41214,N_41088);
and U41549 (N_41549,N_41041,N_41112);
and U41550 (N_41550,N_41016,N_41291);
nor U41551 (N_41551,N_41194,N_41123);
nor U41552 (N_41552,N_41370,N_41343);
or U41553 (N_41553,N_41000,N_41470);
nor U41554 (N_41554,N_41078,N_41040);
and U41555 (N_41555,N_41136,N_41247);
and U41556 (N_41556,N_41126,N_41166);
xor U41557 (N_41557,N_41252,N_41227);
nand U41558 (N_41558,N_41265,N_41384);
and U41559 (N_41559,N_41388,N_41231);
and U41560 (N_41560,N_41071,N_41353);
nor U41561 (N_41561,N_41319,N_41349);
nand U41562 (N_41562,N_41382,N_41069);
nand U41563 (N_41563,N_41458,N_41206);
or U41564 (N_41564,N_41406,N_41115);
nor U41565 (N_41565,N_41459,N_41191);
nand U41566 (N_41566,N_41200,N_41243);
nor U41567 (N_41567,N_41259,N_41017);
xor U41568 (N_41568,N_41436,N_41321);
nand U41569 (N_41569,N_41425,N_41087);
nor U41570 (N_41570,N_41308,N_41322);
nand U41571 (N_41571,N_41419,N_41043);
xor U41572 (N_41572,N_41138,N_41479);
or U41573 (N_41573,N_41346,N_41305);
and U41574 (N_41574,N_41049,N_41236);
nor U41575 (N_41575,N_41331,N_41150);
or U41576 (N_41576,N_41086,N_41283);
nand U41577 (N_41577,N_41056,N_41416);
or U41578 (N_41578,N_41209,N_41445);
and U41579 (N_41579,N_41053,N_41497);
and U41580 (N_41580,N_41475,N_41156);
or U41581 (N_41581,N_41030,N_41064);
and U41582 (N_41582,N_41198,N_41426);
and U41583 (N_41583,N_41244,N_41310);
nor U41584 (N_41584,N_41466,N_41262);
or U41585 (N_41585,N_41018,N_41494);
xnor U41586 (N_41586,N_41477,N_41362);
or U41587 (N_41587,N_41059,N_41374);
and U41588 (N_41588,N_41060,N_41473);
and U41589 (N_41589,N_41312,N_41220);
nand U41590 (N_41590,N_41270,N_41369);
and U41591 (N_41591,N_41235,N_41340);
nor U41592 (N_41592,N_41344,N_41326);
or U41593 (N_41593,N_41172,N_41075);
or U41594 (N_41594,N_41258,N_41005);
and U41595 (N_41595,N_41309,N_41281);
nand U41596 (N_41596,N_41315,N_41196);
nor U41597 (N_41597,N_41176,N_41491);
or U41598 (N_41598,N_41337,N_41225);
nand U41599 (N_41599,N_41028,N_41435);
nand U41600 (N_41600,N_41415,N_41192);
nand U41601 (N_41601,N_41033,N_41493);
or U41602 (N_41602,N_41062,N_41106);
and U41603 (N_41603,N_41065,N_41202);
nand U41604 (N_41604,N_41167,N_41417);
nand U41605 (N_41605,N_41118,N_41208);
nor U41606 (N_41606,N_41213,N_41217);
or U41607 (N_41607,N_41051,N_41450);
and U41608 (N_41608,N_41284,N_41229);
and U41609 (N_41609,N_41440,N_41365);
or U41610 (N_41610,N_41405,N_41433);
and U41611 (N_41611,N_41226,N_41318);
or U41612 (N_41612,N_41197,N_41422);
and U41613 (N_41613,N_41495,N_41489);
nand U41614 (N_41614,N_41285,N_41264);
and U41615 (N_41615,N_41300,N_41157);
nor U41616 (N_41616,N_41468,N_41414);
nand U41617 (N_41617,N_41042,N_41114);
or U41618 (N_41618,N_41429,N_41081);
or U41619 (N_41619,N_41048,N_41095);
nor U41620 (N_41620,N_41147,N_41398);
nand U41621 (N_41621,N_41108,N_41375);
and U41622 (N_41622,N_41190,N_41237);
or U41623 (N_41623,N_41224,N_41025);
nand U41624 (N_41624,N_41072,N_41452);
and U41625 (N_41625,N_41385,N_41327);
or U41626 (N_41626,N_41428,N_41446);
and U41627 (N_41627,N_41153,N_41100);
and U41628 (N_41628,N_41467,N_41316);
nand U41629 (N_41629,N_41476,N_41210);
and U41630 (N_41630,N_41357,N_41096);
nor U41631 (N_41631,N_41068,N_41180);
or U41632 (N_41632,N_41009,N_41387);
nor U41633 (N_41633,N_41129,N_41135);
and U41634 (N_41634,N_41144,N_41139);
and U41635 (N_41635,N_41151,N_41404);
xor U41636 (N_41636,N_41022,N_41070);
nor U41637 (N_41637,N_41268,N_41019);
xnor U41638 (N_41638,N_41061,N_41304);
nand U41639 (N_41639,N_41254,N_41161);
nor U41640 (N_41640,N_41462,N_41286);
or U41641 (N_41641,N_41205,N_41498);
nor U41642 (N_41642,N_41074,N_41107);
and U41643 (N_41643,N_41314,N_41021);
and U41644 (N_41644,N_41257,N_41038);
and U41645 (N_41645,N_41110,N_41255);
and U41646 (N_41646,N_41113,N_41484);
and U41647 (N_41647,N_41211,N_41124);
or U41648 (N_41648,N_41376,N_41367);
or U41649 (N_41649,N_41298,N_41127);
or U41650 (N_41650,N_41330,N_41117);
or U41651 (N_41651,N_41431,N_41241);
nor U41652 (N_41652,N_41128,N_41092);
nand U41653 (N_41653,N_41463,N_41432);
nand U41654 (N_41654,N_41372,N_41492);
or U41655 (N_41655,N_41469,N_41222);
and U41656 (N_41656,N_41482,N_41004);
xnor U41657 (N_41657,N_41083,N_41278);
nand U41658 (N_41658,N_41441,N_41120);
nand U41659 (N_41659,N_41323,N_41294);
and U41660 (N_41660,N_41295,N_41093);
nor U41661 (N_41661,N_41442,N_41456);
or U41662 (N_41662,N_41311,N_41223);
xor U41663 (N_41663,N_41393,N_41207);
nor U41664 (N_41664,N_41336,N_41350);
xnor U41665 (N_41665,N_41444,N_41007);
nor U41666 (N_41666,N_41177,N_41328);
and U41667 (N_41667,N_41239,N_41003);
nand U41668 (N_41668,N_41358,N_41091);
or U41669 (N_41669,N_41366,N_41329);
nand U41670 (N_41670,N_41199,N_41219);
and U41671 (N_41671,N_41185,N_41013);
nor U41672 (N_41672,N_41342,N_41052);
or U41673 (N_41673,N_41154,N_41057);
or U41674 (N_41674,N_41363,N_41486);
and U41675 (N_41675,N_41453,N_41368);
nand U41676 (N_41676,N_41455,N_41116);
nor U41677 (N_41677,N_41292,N_41423);
xnor U41678 (N_41678,N_41080,N_41131);
nand U41679 (N_41679,N_41039,N_41402);
or U41680 (N_41680,N_41188,N_41403);
and U41681 (N_41681,N_41263,N_41221);
or U41682 (N_41682,N_41232,N_41094);
or U41683 (N_41683,N_41215,N_41301);
xor U41684 (N_41684,N_41119,N_41341);
nor U41685 (N_41685,N_41317,N_41253);
or U41686 (N_41686,N_41171,N_41260);
or U41687 (N_41687,N_41320,N_41133);
or U41688 (N_41688,N_41146,N_41276);
and U41689 (N_41689,N_41134,N_41280);
nand U41690 (N_41690,N_41361,N_41020);
or U41691 (N_41691,N_41386,N_41024);
or U41692 (N_41692,N_41145,N_41140);
and U41693 (N_41693,N_41251,N_41098);
nor U41694 (N_41694,N_41289,N_41111);
or U41695 (N_41695,N_41332,N_41026);
xnor U41696 (N_41696,N_41182,N_41149);
nand U41697 (N_41697,N_41102,N_41193);
nor U41698 (N_41698,N_41141,N_41090);
nor U41699 (N_41699,N_41471,N_41216);
and U41700 (N_41700,N_41162,N_41279);
or U41701 (N_41701,N_41411,N_41073);
or U41702 (N_41702,N_41245,N_41246);
nor U41703 (N_41703,N_41296,N_41401);
nor U41704 (N_41704,N_41125,N_41373);
or U41705 (N_41705,N_41307,N_41066);
xnor U41706 (N_41706,N_41036,N_41271);
nand U41707 (N_41707,N_41168,N_41104);
nand U41708 (N_41708,N_41044,N_41170);
and U41709 (N_41709,N_41240,N_41097);
or U41710 (N_41710,N_41306,N_41058);
and U41711 (N_41711,N_41027,N_41076);
nand U41712 (N_41712,N_41437,N_41228);
or U41713 (N_41713,N_41002,N_41045);
and U41714 (N_41714,N_41359,N_41410);
nor U41715 (N_41715,N_41485,N_41184);
xnor U41716 (N_41716,N_41242,N_41297);
nand U41717 (N_41717,N_41377,N_41121);
nand U41718 (N_41718,N_41105,N_41293);
or U41719 (N_41719,N_41101,N_41248);
nand U41720 (N_41720,N_41448,N_41137);
nor U41721 (N_41721,N_41339,N_41430);
or U41722 (N_41722,N_41488,N_41189);
or U41723 (N_41723,N_41478,N_41334);
xnor U41724 (N_41724,N_41012,N_41032);
nor U41725 (N_41725,N_41250,N_41195);
or U41726 (N_41726,N_41037,N_41457);
xnor U41727 (N_41727,N_41443,N_41046);
and U41728 (N_41728,N_41261,N_41099);
xnor U41729 (N_41729,N_41449,N_41413);
and U41730 (N_41730,N_41354,N_41464);
nand U41731 (N_41731,N_41035,N_41179);
or U41732 (N_41732,N_41174,N_41454);
nand U41733 (N_41733,N_41407,N_41047);
nand U41734 (N_41734,N_41143,N_41480);
nand U41735 (N_41735,N_41460,N_41439);
xor U41736 (N_41736,N_41394,N_41273);
nor U41737 (N_41737,N_41356,N_41186);
or U41738 (N_41738,N_41399,N_41233);
and U41739 (N_41739,N_41438,N_41287);
nor U41740 (N_41740,N_41085,N_41379);
nor U41741 (N_41741,N_41249,N_41481);
nor U41742 (N_41742,N_41163,N_41465);
nand U41743 (N_41743,N_41391,N_41499);
or U41744 (N_41744,N_41427,N_41082);
or U41745 (N_41745,N_41380,N_41392);
and U41746 (N_41746,N_41474,N_41302);
or U41747 (N_41747,N_41122,N_41183);
nand U41748 (N_41748,N_41333,N_41360);
and U41749 (N_41749,N_41434,N_41169);
xnor U41750 (N_41750,N_41393,N_41072);
and U41751 (N_41751,N_41451,N_41304);
xor U41752 (N_41752,N_41243,N_41011);
nand U41753 (N_41753,N_41491,N_41472);
nor U41754 (N_41754,N_41079,N_41159);
nor U41755 (N_41755,N_41138,N_41056);
and U41756 (N_41756,N_41367,N_41212);
and U41757 (N_41757,N_41181,N_41176);
and U41758 (N_41758,N_41047,N_41034);
and U41759 (N_41759,N_41434,N_41462);
and U41760 (N_41760,N_41139,N_41326);
nand U41761 (N_41761,N_41312,N_41182);
and U41762 (N_41762,N_41261,N_41101);
xnor U41763 (N_41763,N_41400,N_41167);
and U41764 (N_41764,N_41122,N_41015);
nor U41765 (N_41765,N_41217,N_41110);
nand U41766 (N_41766,N_41208,N_41127);
nand U41767 (N_41767,N_41370,N_41012);
nand U41768 (N_41768,N_41029,N_41206);
or U41769 (N_41769,N_41219,N_41200);
nor U41770 (N_41770,N_41208,N_41463);
nor U41771 (N_41771,N_41216,N_41240);
or U41772 (N_41772,N_41038,N_41065);
nor U41773 (N_41773,N_41264,N_41358);
nor U41774 (N_41774,N_41384,N_41147);
nor U41775 (N_41775,N_41375,N_41040);
or U41776 (N_41776,N_41288,N_41187);
nor U41777 (N_41777,N_41479,N_41396);
nor U41778 (N_41778,N_41169,N_41007);
or U41779 (N_41779,N_41497,N_41449);
or U41780 (N_41780,N_41104,N_41156);
nor U41781 (N_41781,N_41342,N_41212);
or U41782 (N_41782,N_41380,N_41470);
or U41783 (N_41783,N_41464,N_41341);
nor U41784 (N_41784,N_41296,N_41210);
and U41785 (N_41785,N_41416,N_41219);
nor U41786 (N_41786,N_41333,N_41225);
nor U41787 (N_41787,N_41241,N_41178);
nand U41788 (N_41788,N_41493,N_41203);
xnor U41789 (N_41789,N_41010,N_41438);
or U41790 (N_41790,N_41092,N_41389);
or U41791 (N_41791,N_41170,N_41248);
xnor U41792 (N_41792,N_41204,N_41432);
or U41793 (N_41793,N_41083,N_41359);
xnor U41794 (N_41794,N_41081,N_41278);
nand U41795 (N_41795,N_41242,N_41374);
nor U41796 (N_41796,N_41230,N_41347);
nand U41797 (N_41797,N_41385,N_41365);
nand U41798 (N_41798,N_41163,N_41308);
and U41799 (N_41799,N_41245,N_41015);
nor U41800 (N_41800,N_41147,N_41163);
nand U41801 (N_41801,N_41084,N_41236);
and U41802 (N_41802,N_41199,N_41280);
nor U41803 (N_41803,N_41053,N_41325);
nor U41804 (N_41804,N_41281,N_41371);
and U41805 (N_41805,N_41399,N_41254);
or U41806 (N_41806,N_41028,N_41220);
nand U41807 (N_41807,N_41235,N_41025);
nor U41808 (N_41808,N_41277,N_41350);
nor U41809 (N_41809,N_41485,N_41088);
nand U41810 (N_41810,N_41321,N_41497);
or U41811 (N_41811,N_41358,N_41061);
nand U41812 (N_41812,N_41062,N_41019);
xor U41813 (N_41813,N_41331,N_41193);
and U41814 (N_41814,N_41318,N_41228);
nand U41815 (N_41815,N_41250,N_41123);
nor U41816 (N_41816,N_41487,N_41193);
nor U41817 (N_41817,N_41285,N_41008);
nor U41818 (N_41818,N_41038,N_41052);
nor U41819 (N_41819,N_41490,N_41308);
and U41820 (N_41820,N_41037,N_41204);
and U41821 (N_41821,N_41251,N_41092);
xnor U41822 (N_41822,N_41288,N_41394);
nor U41823 (N_41823,N_41279,N_41240);
or U41824 (N_41824,N_41093,N_41187);
xnor U41825 (N_41825,N_41013,N_41368);
nor U41826 (N_41826,N_41241,N_41497);
or U41827 (N_41827,N_41324,N_41082);
and U41828 (N_41828,N_41498,N_41351);
nor U41829 (N_41829,N_41411,N_41205);
nand U41830 (N_41830,N_41210,N_41273);
and U41831 (N_41831,N_41018,N_41472);
and U41832 (N_41832,N_41248,N_41226);
or U41833 (N_41833,N_41015,N_41151);
nand U41834 (N_41834,N_41452,N_41191);
xor U41835 (N_41835,N_41392,N_41151);
and U41836 (N_41836,N_41183,N_41124);
or U41837 (N_41837,N_41205,N_41382);
nor U41838 (N_41838,N_41114,N_41488);
or U41839 (N_41839,N_41414,N_41044);
xnor U41840 (N_41840,N_41284,N_41455);
or U41841 (N_41841,N_41119,N_41299);
nor U41842 (N_41842,N_41056,N_41131);
nand U41843 (N_41843,N_41281,N_41111);
xnor U41844 (N_41844,N_41375,N_41174);
nor U41845 (N_41845,N_41447,N_41300);
nor U41846 (N_41846,N_41258,N_41300);
xnor U41847 (N_41847,N_41068,N_41202);
or U41848 (N_41848,N_41009,N_41146);
or U41849 (N_41849,N_41418,N_41489);
nor U41850 (N_41850,N_41224,N_41249);
nand U41851 (N_41851,N_41221,N_41444);
nor U41852 (N_41852,N_41052,N_41015);
nor U41853 (N_41853,N_41484,N_41399);
or U41854 (N_41854,N_41042,N_41043);
or U41855 (N_41855,N_41363,N_41038);
and U41856 (N_41856,N_41073,N_41377);
and U41857 (N_41857,N_41017,N_41263);
and U41858 (N_41858,N_41179,N_41487);
or U41859 (N_41859,N_41033,N_41199);
or U41860 (N_41860,N_41481,N_41193);
or U41861 (N_41861,N_41345,N_41027);
or U41862 (N_41862,N_41444,N_41360);
nand U41863 (N_41863,N_41492,N_41383);
or U41864 (N_41864,N_41382,N_41261);
nand U41865 (N_41865,N_41053,N_41447);
nor U41866 (N_41866,N_41283,N_41051);
xor U41867 (N_41867,N_41274,N_41091);
or U41868 (N_41868,N_41377,N_41076);
nand U41869 (N_41869,N_41424,N_41067);
nand U41870 (N_41870,N_41415,N_41467);
nand U41871 (N_41871,N_41139,N_41129);
and U41872 (N_41872,N_41016,N_41188);
or U41873 (N_41873,N_41066,N_41092);
and U41874 (N_41874,N_41133,N_41432);
nor U41875 (N_41875,N_41090,N_41129);
and U41876 (N_41876,N_41226,N_41021);
xor U41877 (N_41877,N_41045,N_41372);
or U41878 (N_41878,N_41376,N_41043);
nand U41879 (N_41879,N_41495,N_41037);
and U41880 (N_41880,N_41425,N_41431);
nand U41881 (N_41881,N_41457,N_41317);
or U41882 (N_41882,N_41167,N_41085);
nor U41883 (N_41883,N_41263,N_41154);
or U41884 (N_41884,N_41191,N_41168);
xnor U41885 (N_41885,N_41037,N_41051);
nor U41886 (N_41886,N_41364,N_41320);
xor U41887 (N_41887,N_41397,N_41045);
nand U41888 (N_41888,N_41484,N_41324);
nand U41889 (N_41889,N_41071,N_41047);
or U41890 (N_41890,N_41429,N_41103);
nand U41891 (N_41891,N_41176,N_41111);
nand U41892 (N_41892,N_41345,N_41087);
nor U41893 (N_41893,N_41012,N_41066);
and U41894 (N_41894,N_41295,N_41212);
or U41895 (N_41895,N_41271,N_41225);
or U41896 (N_41896,N_41333,N_41251);
nor U41897 (N_41897,N_41293,N_41498);
and U41898 (N_41898,N_41474,N_41496);
nor U41899 (N_41899,N_41040,N_41152);
or U41900 (N_41900,N_41386,N_41147);
nor U41901 (N_41901,N_41366,N_41300);
nor U41902 (N_41902,N_41220,N_41022);
xor U41903 (N_41903,N_41386,N_41329);
nor U41904 (N_41904,N_41091,N_41382);
nor U41905 (N_41905,N_41245,N_41440);
and U41906 (N_41906,N_41363,N_41346);
nor U41907 (N_41907,N_41483,N_41452);
and U41908 (N_41908,N_41358,N_41193);
and U41909 (N_41909,N_41261,N_41070);
xor U41910 (N_41910,N_41285,N_41357);
nand U41911 (N_41911,N_41024,N_41416);
and U41912 (N_41912,N_41081,N_41092);
or U41913 (N_41913,N_41148,N_41488);
nor U41914 (N_41914,N_41330,N_41487);
and U41915 (N_41915,N_41456,N_41349);
nor U41916 (N_41916,N_41479,N_41146);
or U41917 (N_41917,N_41299,N_41034);
nor U41918 (N_41918,N_41410,N_41017);
nor U41919 (N_41919,N_41083,N_41325);
or U41920 (N_41920,N_41223,N_41032);
or U41921 (N_41921,N_41078,N_41010);
and U41922 (N_41922,N_41469,N_41248);
xnor U41923 (N_41923,N_41184,N_41220);
or U41924 (N_41924,N_41419,N_41218);
nand U41925 (N_41925,N_41204,N_41478);
nand U41926 (N_41926,N_41393,N_41199);
and U41927 (N_41927,N_41464,N_41329);
nand U41928 (N_41928,N_41363,N_41273);
xor U41929 (N_41929,N_41385,N_41326);
nor U41930 (N_41930,N_41189,N_41122);
or U41931 (N_41931,N_41496,N_41424);
or U41932 (N_41932,N_41456,N_41075);
xor U41933 (N_41933,N_41277,N_41352);
or U41934 (N_41934,N_41314,N_41070);
and U41935 (N_41935,N_41082,N_41316);
or U41936 (N_41936,N_41401,N_41342);
and U41937 (N_41937,N_41120,N_41111);
and U41938 (N_41938,N_41173,N_41166);
and U41939 (N_41939,N_41356,N_41367);
xnor U41940 (N_41940,N_41123,N_41435);
and U41941 (N_41941,N_41135,N_41166);
xnor U41942 (N_41942,N_41038,N_41233);
or U41943 (N_41943,N_41236,N_41198);
or U41944 (N_41944,N_41206,N_41471);
and U41945 (N_41945,N_41024,N_41347);
or U41946 (N_41946,N_41175,N_41481);
nand U41947 (N_41947,N_41419,N_41013);
or U41948 (N_41948,N_41369,N_41333);
nor U41949 (N_41949,N_41483,N_41115);
or U41950 (N_41950,N_41068,N_41428);
and U41951 (N_41951,N_41006,N_41201);
and U41952 (N_41952,N_41454,N_41290);
and U41953 (N_41953,N_41172,N_41197);
nor U41954 (N_41954,N_41350,N_41070);
and U41955 (N_41955,N_41332,N_41393);
and U41956 (N_41956,N_41182,N_41260);
nand U41957 (N_41957,N_41314,N_41121);
nor U41958 (N_41958,N_41190,N_41392);
nor U41959 (N_41959,N_41075,N_41196);
nor U41960 (N_41960,N_41054,N_41024);
and U41961 (N_41961,N_41308,N_41179);
and U41962 (N_41962,N_41229,N_41433);
nand U41963 (N_41963,N_41132,N_41153);
nand U41964 (N_41964,N_41044,N_41491);
nand U41965 (N_41965,N_41297,N_41027);
nor U41966 (N_41966,N_41079,N_41192);
nand U41967 (N_41967,N_41486,N_41219);
xor U41968 (N_41968,N_41445,N_41370);
nor U41969 (N_41969,N_41318,N_41183);
or U41970 (N_41970,N_41074,N_41386);
nor U41971 (N_41971,N_41112,N_41413);
nand U41972 (N_41972,N_41342,N_41346);
nand U41973 (N_41973,N_41499,N_41087);
nor U41974 (N_41974,N_41312,N_41441);
nor U41975 (N_41975,N_41398,N_41373);
nand U41976 (N_41976,N_41370,N_41310);
or U41977 (N_41977,N_41410,N_41181);
nor U41978 (N_41978,N_41023,N_41073);
nand U41979 (N_41979,N_41252,N_41260);
or U41980 (N_41980,N_41399,N_41079);
or U41981 (N_41981,N_41384,N_41158);
nand U41982 (N_41982,N_41231,N_41023);
nand U41983 (N_41983,N_41484,N_41104);
nand U41984 (N_41984,N_41311,N_41221);
and U41985 (N_41985,N_41137,N_41103);
or U41986 (N_41986,N_41321,N_41042);
or U41987 (N_41987,N_41241,N_41205);
nand U41988 (N_41988,N_41166,N_41481);
or U41989 (N_41989,N_41235,N_41407);
nand U41990 (N_41990,N_41443,N_41466);
or U41991 (N_41991,N_41354,N_41429);
and U41992 (N_41992,N_41152,N_41173);
nand U41993 (N_41993,N_41386,N_41269);
nand U41994 (N_41994,N_41129,N_41441);
nand U41995 (N_41995,N_41479,N_41139);
nor U41996 (N_41996,N_41470,N_41388);
nand U41997 (N_41997,N_41416,N_41349);
nand U41998 (N_41998,N_41137,N_41148);
nor U41999 (N_41999,N_41224,N_41169);
nor U42000 (N_42000,N_41845,N_41881);
or U42001 (N_42001,N_41981,N_41975);
and U42002 (N_42002,N_41634,N_41528);
and U42003 (N_42003,N_41710,N_41512);
and U42004 (N_42004,N_41912,N_41660);
nor U42005 (N_42005,N_41958,N_41850);
nor U42006 (N_42006,N_41685,N_41805);
and U42007 (N_42007,N_41521,N_41530);
or U42008 (N_42008,N_41987,N_41852);
nand U42009 (N_42009,N_41918,N_41813);
nand U42010 (N_42010,N_41826,N_41747);
nor U42011 (N_42011,N_41846,N_41992);
nand U42012 (N_42012,N_41500,N_41983);
nand U42013 (N_42013,N_41984,N_41926);
and U42014 (N_42014,N_41879,N_41535);
or U42015 (N_42015,N_41891,N_41777);
and U42016 (N_42016,N_41915,N_41695);
or U42017 (N_42017,N_41865,N_41651);
nand U42018 (N_42018,N_41570,N_41827);
nor U42019 (N_42019,N_41972,N_41741);
nor U42020 (N_42020,N_41682,N_41726);
nand U42021 (N_42021,N_41809,N_41697);
and U42022 (N_42022,N_41783,N_41893);
xor U42023 (N_42023,N_41889,N_41633);
nor U42024 (N_42024,N_41593,N_41626);
or U42025 (N_42025,N_41948,N_41877);
or U42026 (N_42026,N_41995,N_41672);
or U42027 (N_42027,N_41962,N_41637);
or U42028 (N_42028,N_41872,N_41727);
or U42029 (N_42029,N_41774,N_41916);
nor U42030 (N_42030,N_41970,N_41661);
or U42031 (N_42031,N_41990,N_41675);
and U42032 (N_42032,N_41755,N_41834);
or U42033 (N_42033,N_41980,N_41867);
and U42034 (N_42034,N_41770,N_41931);
or U42035 (N_42035,N_41604,N_41577);
nand U42036 (N_42036,N_41533,N_41771);
nor U42037 (N_42037,N_41767,N_41555);
nand U42038 (N_42038,N_41698,N_41804);
or U42039 (N_42039,N_41789,N_41642);
xnor U42040 (N_42040,N_41717,N_41875);
nor U42041 (N_42041,N_41502,N_41572);
and U42042 (N_42042,N_41764,N_41922);
or U42043 (N_42043,N_41700,N_41607);
or U42044 (N_42044,N_41635,N_41947);
or U42045 (N_42045,N_41973,N_41788);
nor U42046 (N_42046,N_41897,N_41745);
nand U42047 (N_42047,N_41649,N_41799);
or U42048 (N_42048,N_41684,N_41861);
and U42049 (N_42049,N_41884,N_41561);
xnor U42050 (N_42050,N_41520,N_41778);
or U42051 (N_42051,N_41559,N_41974);
and U42052 (N_42052,N_41668,N_41539);
nand U42053 (N_42053,N_41587,N_41930);
and U42054 (N_42054,N_41655,N_41993);
nor U42055 (N_42055,N_41686,N_41580);
nand U42056 (N_42056,N_41558,N_41784);
or U42057 (N_42057,N_41526,N_41624);
or U42058 (N_42058,N_41880,N_41927);
nor U42059 (N_42059,N_41696,N_41692);
nor U42060 (N_42060,N_41776,N_41574);
or U42061 (N_42061,N_41951,N_41567);
xor U42062 (N_42062,N_41838,N_41869);
or U42063 (N_42063,N_41605,N_41775);
nand U42064 (N_42064,N_41841,N_41708);
xor U42065 (N_42065,N_41718,N_41803);
nor U42066 (N_42066,N_41669,N_41553);
nor U42067 (N_42067,N_41825,N_41818);
or U42068 (N_42068,N_41627,N_41853);
or U42069 (N_42069,N_41878,N_41608);
nor U42070 (N_42070,N_41966,N_41595);
or U42071 (N_42071,N_41954,N_41596);
nand U42072 (N_42072,N_41597,N_41740);
nor U42073 (N_42073,N_41511,N_41699);
xnor U42074 (N_42074,N_41529,N_41516);
nor U42075 (N_42075,N_41814,N_41819);
nor U42076 (N_42076,N_41901,N_41610);
or U42077 (N_42077,N_41806,N_41899);
and U42078 (N_42078,N_41664,N_41937);
nand U42079 (N_42079,N_41705,N_41736);
and U42080 (N_42080,N_41791,N_41870);
nor U42081 (N_42081,N_41863,N_41681);
nand U42082 (N_42082,N_41653,N_41578);
nor U42083 (N_42083,N_41956,N_41934);
or U42084 (N_42084,N_41792,N_41584);
xor U42085 (N_42085,N_41911,N_41991);
nand U42086 (N_42086,N_41560,N_41601);
or U42087 (N_42087,N_41501,N_41541);
or U42088 (N_42088,N_41965,N_41753);
and U42089 (N_42089,N_41734,N_41543);
nand U42090 (N_42090,N_41657,N_41550);
nor U42091 (N_42091,N_41913,N_41647);
nor U42092 (N_42092,N_41821,N_41998);
nand U42093 (N_42093,N_41706,N_41786);
or U42094 (N_42094,N_41527,N_41517);
and U42095 (N_42095,N_41858,N_41554);
or U42096 (N_42096,N_41942,N_41557);
or U42097 (N_42097,N_41617,N_41831);
nor U42098 (N_42098,N_41976,N_41691);
nor U42099 (N_42099,N_41822,N_41896);
nor U42100 (N_42100,N_41750,N_41670);
or U42101 (N_42101,N_41963,N_41632);
and U42102 (N_42102,N_41645,N_41694);
nor U42103 (N_42103,N_41807,N_41997);
nor U42104 (N_42104,N_41523,N_41795);
or U42105 (N_42105,N_41940,N_41630);
or U42106 (N_42106,N_41882,N_41739);
nor U42107 (N_42107,N_41961,N_41854);
and U42108 (N_42108,N_41599,N_41615);
and U42109 (N_42109,N_41828,N_41644);
nor U42110 (N_42110,N_41728,N_41999);
nand U42111 (N_42111,N_41782,N_41800);
and U42112 (N_42112,N_41503,N_41628);
nor U42113 (N_42113,N_41921,N_41715);
xor U42114 (N_42114,N_41712,N_41967);
and U42115 (N_42115,N_41920,N_41643);
nand U42116 (N_42116,N_41674,N_41876);
or U42117 (N_42117,N_41689,N_41742);
nand U42118 (N_42118,N_41549,N_41659);
or U42119 (N_42119,N_41702,N_41538);
nor U42120 (N_42120,N_41888,N_41725);
xnor U42121 (N_42121,N_41687,N_41908);
nand U42122 (N_42122,N_41514,N_41982);
nand U42123 (N_42123,N_41812,N_41864);
and U42124 (N_42124,N_41576,N_41785);
nand U42125 (N_42125,N_41796,N_41860);
nand U42126 (N_42126,N_41761,N_41534);
or U42127 (N_42127,N_41746,N_41636);
nor U42128 (N_42128,N_41510,N_41840);
nand U42129 (N_42129,N_41646,N_41724);
and U42130 (N_42130,N_41959,N_41760);
or U42131 (N_42131,N_41892,N_41594);
xnor U42132 (N_42132,N_41751,N_41735);
or U42133 (N_42133,N_41671,N_41979);
xnor U42134 (N_42134,N_41569,N_41666);
nor U42135 (N_42135,N_41953,N_41552);
nand U42136 (N_42136,N_41773,N_41787);
nand U42137 (N_42137,N_41903,N_41756);
xor U42138 (N_42138,N_41939,N_41509);
and U42139 (N_42139,N_41568,N_41677);
nor U42140 (N_42140,N_41589,N_41619);
or U42141 (N_42141,N_41588,N_41690);
or U42142 (N_42142,N_41964,N_41754);
nor U42143 (N_42143,N_41829,N_41808);
or U42144 (N_42144,N_41729,N_41547);
nor U42145 (N_42145,N_41525,N_41600);
nor U42146 (N_42146,N_41744,N_41612);
nand U42147 (N_42147,N_41790,N_41551);
nand U42148 (N_42148,N_41874,N_41562);
or U42149 (N_42149,N_41923,N_41978);
nand U42150 (N_42150,N_41842,N_41592);
nand U42151 (N_42151,N_41932,N_41650);
and U42152 (N_42152,N_41943,N_41810);
and U42153 (N_42153,N_41749,N_41855);
or U42154 (N_42154,N_41946,N_41638);
and U42155 (N_42155,N_41917,N_41765);
nor U42156 (N_42156,N_41815,N_41618);
or U42157 (N_42157,N_41909,N_41847);
nand U42158 (N_42158,N_41900,N_41833);
or U42159 (N_42159,N_41679,N_41733);
and U42160 (N_42160,N_41950,N_41641);
or U42161 (N_42161,N_41622,N_41794);
or U42162 (N_42162,N_41748,N_41986);
nand U42163 (N_42163,N_41602,N_41581);
or U42164 (N_42164,N_41971,N_41832);
nor U42165 (N_42165,N_41565,N_41907);
and U42166 (N_42166,N_41656,N_41598);
nor U42167 (N_42167,N_41737,N_41573);
or U42168 (N_42168,N_41563,N_41758);
or U42169 (N_42169,N_41839,N_41835);
and U42170 (N_42170,N_41933,N_41508);
or U42171 (N_42171,N_41658,N_41654);
nor U42172 (N_42172,N_41868,N_41518);
and U42173 (N_42173,N_41722,N_41949);
nor U42174 (N_42174,N_41713,N_41723);
nor U42175 (N_42175,N_41762,N_41779);
or U42176 (N_42176,N_41769,N_41887);
nor U42177 (N_42177,N_41988,N_41614);
nor U42178 (N_42178,N_41556,N_41609);
nand U42179 (N_42179,N_41781,N_41802);
nand U42180 (N_42180,N_41640,N_41851);
nor U42181 (N_42181,N_41575,N_41531);
and U42182 (N_42182,N_41844,N_41603);
nor U42183 (N_42183,N_41537,N_41830);
and U42184 (N_42184,N_41507,N_41583);
nand U42185 (N_42185,N_41902,N_41929);
nor U42186 (N_42186,N_41886,N_41611);
nor U42187 (N_42187,N_41590,N_41925);
or U42188 (N_42188,N_41662,N_41732);
or U42189 (N_42189,N_41629,N_41859);
and U42190 (N_42190,N_41857,N_41673);
or U42191 (N_42191,N_41977,N_41957);
nor U42192 (N_42192,N_41564,N_41969);
or U42193 (N_42193,N_41613,N_41936);
and U42194 (N_42194,N_41836,N_41924);
nor U42195 (N_42195,N_41542,N_41941);
and U42196 (N_42196,N_41620,N_41811);
or U42197 (N_42197,N_41505,N_41890);
nand U42198 (N_42198,N_41904,N_41848);
nor U42199 (N_42199,N_41985,N_41680);
nor U42200 (N_42200,N_41506,N_41793);
nor U42201 (N_42201,N_41519,N_41652);
and U42202 (N_42202,N_41766,N_41823);
xor U42203 (N_42203,N_41738,N_41873);
or U42204 (N_42204,N_41952,N_41616);
or U42205 (N_42205,N_41566,N_41743);
nor U42206 (N_42206,N_41704,N_41955);
or U42207 (N_42207,N_41989,N_41721);
nand U42208 (N_42208,N_41768,N_41678);
nand U42209 (N_42209,N_41910,N_41513);
and U42210 (N_42210,N_41548,N_41663);
xor U42211 (N_42211,N_41591,N_41862);
or U42212 (N_42212,N_41683,N_41763);
or U42213 (N_42213,N_41639,N_41579);
nand U42214 (N_42214,N_41960,N_41504);
or U42215 (N_42215,N_41843,N_41703);
nand U42216 (N_42216,N_41797,N_41667);
nand U42217 (N_42217,N_41898,N_41945);
nor U42218 (N_42218,N_41772,N_41720);
nand U42219 (N_42219,N_41856,N_41895);
nor U42220 (N_42220,N_41544,N_41688);
nand U42221 (N_42221,N_41817,N_41709);
nand U42222 (N_42222,N_41540,N_41707);
nand U42223 (N_42223,N_41801,N_41665);
or U42224 (N_42224,N_41730,N_41515);
xor U42225 (N_42225,N_41935,N_41586);
nand U42226 (N_42226,N_41919,N_41798);
or U42227 (N_42227,N_41522,N_41631);
nor U42228 (N_42228,N_41714,N_41837);
nand U42229 (N_42229,N_41711,N_41994);
nor U42230 (N_42230,N_41582,N_41571);
nand U42231 (N_42231,N_41585,N_41780);
nand U42232 (N_42232,N_41757,N_41536);
xnor U42233 (N_42233,N_41625,N_41623);
or U42234 (N_42234,N_41676,N_41532);
xnor U42235 (N_42235,N_41906,N_41524);
or U42236 (N_42236,N_41871,N_41701);
xnor U42237 (N_42237,N_41546,N_41905);
nand U42238 (N_42238,N_41719,N_41824);
xnor U42239 (N_42239,N_41968,N_41938);
and U42240 (N_42240,N_41885,N_41545);
or U42241 (N_42241,N_41693,N_41928);
or U42242 (N_42242,N_41996,N_41883);
or U42243 (N_42243,N_41866,N_41621);
nor U42244 (N_42244,N_41820,N_41816);
and U42245 (N_42245,N_41606,N_41894);
or U42246 (N_42246,N_41849,N_41752);
xnor U42247 (N_42247,N_41944,N_41716);
nand U42248 (N_42248,N_41648,N_41731);
or U42249 (N_42249,N_41914,N_41759);
or U42250 (N_42250,N_41878,N_41764);
or U42251 (N_42251,N_41772,N_41715);
nand U42252 (N_42252,N_41721,N_41590);
nand U42253 (N_42253,N_41668,N_41767);
and U42254 (N_42254,N_41845,N_41945);
nand U42255 (N_42255,N_41944,N_41769);
nand U42256 (N_42256,N_41828,N_41605);
nand U42257 (N_42257,N_41565,N_41804);
or U42258 (N_42258,N_41697,N_41588);
nor U42259 (N_42259,N_41902,N_41800);
nand U42260 (N_42260,N_41912,N_41668);
or U42261 (N_42261,N_41742,N_41640);
and U42262 (N_42262,N_41753,N_41885);
nor U42263 (N_42263,N_41605,N_41781);
and U42264 (N_42264,N_41541,N_41679);
or U42265 (N_42265,N_41991,N_41970);
and U42266 (N_42266,N_41583,N_41512);
and U42267 (N_42267,N_41603,N_41839);
nor U42268 (N_42268,N_41889,N_41567);
or U42269 (N_42269,N_41823,N_41503);
and U42270 (N_42270,N_41543,N_41583);
nand U42271 (N_42271,N_41648,N_41600);
or U42272 (N_42272,N_41921,N_41714);
nand U42273 (N_42273,N_41558,N_41902);
or U42274 (N_42274,N_41943,N_41966);
or U42275 (N_42275,N_41802,N_41535);
nand U42276 (N_42276,N_41877,N_41717);
and U42277 (N_42277,N_41959,N_41851);
nand U42278 (N_42278,N_41771,N_41736);
nor U42279 (N_42279,N_41525,N_41974);
and U42280 (N_42280,N_41581,N_41579);
and U42281 (N_42281,N_41733,N_41925);
and U42282 (N_42282,N_41940,N_41696);
or U42283 (N_42283,N_41541,N_41763);
and U42284 (N_42284,N_41510,N_41939);
and U42285 (N_42285,N_41852,N_41860);
or U42286 (N_42286,N_41833,N_41770);
nor U42287 (N_42287,N_41780,N_41868);
nor U42288 (N_42288,N_41525,N_41841);
or U42289 (N_42289,N_41944,N_41898);
and U42290 (N_42290,N_41893,N_41659);
and U42291 (N_42291,N_41666,N_41732);
and U42292 (N_42292,N_41828,N_41648);
nor U42293 (N_42293,N_41707,N_41562);
and U42294 (N_42294,N_41929,N_41524);
and U42295 (N_42295,N_41918,N_41540);
and U42296 (N_42296,N_41880,N_41515);
nand U42297 (N_42297,N_41941,N_41931);
nand U42298 (N_42298,N_41688,N_41966);
nand U42299 (N_42299,N_41661,N_41895);
nand U42300 (N_42300,N_41694,N_41684);
nor U42301 (N_42301,N_41588,N_41703);
and U42302 (N_42302,N_41914,N_41714);
and U42303 (N_42303,N_41655,N_41606);
nor U42304 (N_42304,N_41708,N_41574);
nand U42305 (N_42305,N_41807,N_41727);
or U42306 (N_42306,N_41737,N_41789);
or U42307 (N_42307,N_41975,N_41949);
nor U42308 (N_42308,N_41846,N_41644);
nor U42309 (N_42309,N_41603,N_41688);
nand U42310 (N_42310,N_41632,N_41666);
nor U42311 (N_42311,N_41785,N_41672);
nor U42312 (N_42312,N_41932,N_41999);
nand U42313 (N_42313,N_41718,N_41881);
nand U42314 (N_42314,N_41893,N_41719);
or U42315 (N_42315,N_41544,N_41637);
xnor U42316 (N_42316,N_41666,N_41765);
nand U42317 (N_42317,N_41740,N_41552);
nand U42318 (N_42318,N_41695,N_41508);
and U42319 (N_42319,N_41583,N_41523);
xor U42320 (N_42320,N_41654,N_41858);
and U42321 (N_42321,N_41979,N_41871);
and U42322 (N_42322,N_41900,N_41927);
or U42323 (N_42323,N_41611,N_41794);
or U42324 (N_42324,N_41680,N_41833);
or U42325 (N_42325,N_41790,N_41624);
or U42326 (N_42326,N_41987,N_41736);
xnor U42327 (N_42327,N_41555,N_41524);
nand U42328 (N_42328,N_41608,N_41556);
or U42329 (N_42329,N_41790,N_41750);
xnor U42330 (N_42330,N_41870,N_41964);
and U42331 (N_42331,N_41893,N_41689);
or U42332 (N_42332,N_41804,N_41881);
nor U42333 (N_42333,N_41793,N_41966);
and U42334 (N_42334,N_41896,N_41715);
and U42335 (N_42335,N_41771,N_41807);
xnor U42336 (N_42336,N_41616,N_41676);
and U42337 (N_42337,N_41555,N_41567);
or U42338 (N_42338,N_41770,N_41642);
and U42339 (N_42339,N_41960,N_41632);
nand U42340 (N_42340,N_41982,N_41841);
or U42341 (N_42341,N_41960,N_41590);
and U42342 (N_42342,N_41841,N_41970);
and U42343 (N_42343,N_41585,N_41583);
or U42344 (N_42344,N_41753,N_41922);
or U42345 (N_42345,N_41586,N_41937);
nand U42346 (N_42346,N_41629,N_41872);
nor U42347 (N_42347,N_41906,N_41611);
or U42348 (N_42348,N_41865,N_41717);
and U42349 (N_42349,N_41587,N_41708);
xor U42350 (N_42350,N_41522,N_41902);
nand U42351 (N_42351,N_41831,N_41602);
nand U42352 (N_42352,N_41893,N_41761);
nand U42353 (N_42353,N_41997,N_41842);
and U42354 (N_42354,N_41686,N_41888);
or U42355 (N_42355,N_41743,N_41952);
and U42356 (N_42356,N_41896,N_41775);
and U42357 (N_42357,N_41653,N_41851);
xnor U42358 (N_42358,N_41959,N_41879);
nand U42359 (N_42359,N_41672,N_41978);
nor U42360 (N_42360,N_41524,N_41980);
and U42361 (N_42361,N_41663,N_41822);
nand U42362 (N_42362,N_41639,N_41526);
nor U42363 (N_42363,N_41997,N_41932);
xnor U42364 (N_42364,N_41659,N_41554);
and U42365 (N_42365,N_41870,N_41673);
or U42366 (N_42366,N_41547,N_41549);
and U42367 (N_42367,N_41597,N_41962);
and U42368 (N_42368,N_41833,N_41832);
nor U42369 (N_42369,N_41746,N_41955);
and U42370 (N_42370,N_41705,N_41826);
and U42371 (N_42371,N_41580,N_41572);
xnor U42372 (N_42372,N_41992,N_41739);
nor U42373 (N_42373,N_41546,N_41690);
nor U42374 (N_42374,N_41571,N_41950);
nand U42375 (N_42375,N_41512,N_41819);
nor U42376 (N_42376,N_41625,N_41697);
or U42377 (N_42377,N_41620,N_41968);
nand U42378 (N_42378,N_41955,N_41503);
xnor U42379 (N_42379,N_41607,N_41873);
or U42380 (N_42380,N_41570,N_41562);
or U42381 (N_42381,N_41558,N_41670);
nand U42382 (N_42382,N_41531,N_41626);
and U42383 (N_42383,N_41576,N_41861);
nor U42384 (N_42384,N_41604,N_41868);
nand U42385 (N_42385,N_41510,N_41904);
nor U42386 (N_42386,N_41910,N_41598);
nand U42387 (N_42387,N_41965,N_41880);
nor U42388 (N_42388,N_41998,N_41762);
or U42389 (N_42389,N_41804,N_41870);
or U42390 (N_42390,N_41983,N_41726);
or U42391 (N_42391,N_41504,N_41930);
and U42392 (N_42392,N_41800,N_41692);
or U42393 (N_42393,N_41870,N_41994);
nand U42394 (N_42394,N_41709,N_41505);
nand U42395 (N_42395,N_41816,N_41823);
and U42396 (N_42396,N_41672,N_41731);
or U42397 (N_42397,N_41827,N_41523);
nor U42398 (N_42398,N_41768,N_41851);
or U42399 (N_42399,N_41607,N_41898);
and U42400 (N_42400,N_41638,N_41664);
or U42401 (N_42401,N_41561,N_41688);
nand U42402 (N_42402,N_41656,N_41583);
nor U42403 (N_42403,N_41743,N_41712);
and U42404 (N_42404,N_41826,N_41591);
nor U42405 (N_42405,N_41758,N_41617);
nand U42406 (N_42406,N_41876,N_41905);
and U42407 (N_42407,N_41785,N_41541);
and U42408 (N_42408,N_41862,N_41883);
and U42409 (N_42409,N_41879,N_41908);
or U42410 (N_42410,N_41936,N_41634);
and U42411 (N_42411,N_41865,N_41725);
nand U42412 (N_42412,N_41523,N_41683);
nand U42413 (N_42413,N_41732,N_41629);
nand U42414 (N_42414,N_41544,N_41755);
or U42415 (N_42415,N_41666,N_41774);
nor U42416 (N_42416,N_41841,N_41629);
xnor U42417 (N_42417,N_41940,N_41990);
xnor U42418 (N_42418,N_41698,N_41678);
nor U42419 (N_42419,N_41552,N_41532);
and U42420 (N_42420,N_41865,N_41974);
nand U42421 (N_42421,N_41928,N_41677);
or U42422 (N_42422,N_41529,N_41540);
nor U42423 (N_42423,N_41882,N_41546);
nor U42424 (N_42424,N_41784,N_41687);
and U42425 (N_42425,N_41675,N_41994);
nor U42426 (N_42426,N_41704,N_41633);
or U42427 (N_42427,N_41523,N_41685);
or U42428 (N_42428,N_41775,N_41824);
nand U42429 (N_42429,N_41614,N_41544);
and U42430 (N_42430,N_41651,N_41967);
or U42431 (N_42431,N_41588,N_41694);
nand U42432 (N_42432,N_41703,N_41616);
and U42433 (N_42433,N_41684,N_41780);
and U42434 (N_42434,N_41758,N_41985);
xnor U42435 (N_42435,N_41756,N_41830);
nor U42436 (N_42436,N_41847,N_41802);
and U42437 (N_42437,N_41686,N_41756);
nor U42438 (N_42438,N_41677,N_41540);
xor U42439 (N_42439,N_41508,N_41775);
nor U42440 (N_42440,N_41963,N_41903);
xor U42441 (N_42441,N_41734,N_41679);
and U42442 (N_42442,N_41972,N_41600);
nand U42443 (N_42443,N_41625,N_41578);
nor U42444 (N_42444,N_41961,N_41869);
nor U42445 (N_42445,N_41622,N_41609);
nor U42446 (N_42446,N_41959,N_41692);
nand U42447 (N_42447,N_41929,N_41698);
or U42448 (N_42448,N_41948,N_41967);
nand U42449 (N_42449,N_41865,N_41796);
nor U42450 (N_42450,N_41784,N_41707);
or U42451 (N_42451,N_41817,N_41713);
and U42452 (N_42452,N_41554,N_41800);
nor U42453 (N_42453,N_41556,N_41646);
and U42454 (N_42454,N_41689,N_41907);
nand U42455 (N_42455,N_41615,N_41639);
or U42456 (N_42456,N_41773,N_41692);
and U42457 (N_42457,N_41913,N_41793);
or U42458 (N_42458,N_41893,N_41921);
or U42459 (N_42459,N_41819,N_41630);
nor U42460 (N_42460,N_41733,N_41919);
nor U42461 (N_42461,N_41669,N_41885);
and U42462 (N_42462,N_41650,N_41539);
and U42463 (N_42463,N_41732,N_41852);
nor U42464 (N_42464,N_41857,N_41690);
nor U42465 (N_42465,N_41729,N_41826);
xnor U42466 (N_42466,N_41965,N_41606);
nor U42467 (N_42467,N_41860,N_41556);
and U42468 (N_42468,N_41865,N_41794);
nor U42469 (N_42469,N_41730,N_41505);
and U42470 (N_42470,N_41619,N_41862);
nand U42471 (N_42471,N_41817,N_41800);
or U42472 (N_42472,N_41875,N_41586);
and U42473 (N_42473,N_41833,N_41704);
and U42474 (N_42474,N_41692,N_41583);
xor U42475 (N_42475,N_41756,N_41827);
or U42476 (N_42476,N_41546,N_41924);
and U42477 (N_42477,N_41926,N_41758);
nand U42478 (N_42478,N_41737,N_41836);
nor U42479 (N_42479,N_41925,N_41954);
nand U42480 (N_42480,N_41605,N_41509);
and U42481 (N_42481,N_41502,N_41806);
nand U42482 (N_42482,N_41945,N_41729);
or U42483 (N_42483,N_41908,N_41506);
xnor U42484 (N_42484,N_41771,N_41520);
or U42485 (N_42485,N_41531,N_41507);
or U42486 (N_42486,N_41660,N_41974);
and U42487 (N_42487,N_41966,N_41784);
xor U42488 (N_42488,N_41979,N_41991);
or U42489 (N_42489,N_41526,N_41915);
nor U42490 (N_42490,N_41508,N_41620);
nor U42491 (N_42491,N_41561,N_41511);
and U42492 (N_42492,N_41989,N_41622);
nor U42493 (N_42493,N_41965,N_41800);
nand U42494 (N_42494,N_41825,N_41839);
nand U42495 (N_42495,N_41751,N_41823);
xnor U42496 (N_42496,N_41974,N_41904);
or U42497 (N_42497,N_41982,N_41890);
nor U42498 (N_42498,N_41786,N_41634);
or U42499 (N_42499,N_41741,N_41882);
nor U42500 (N_42500,N_42189,N_42204);
nor U42501 (N_42501,N_42058,N_42114);
nand U42502 (N_42502,N_42295,N_42442);
nand U42503 (N_42503,N_42237,N_42335);
nand U42504 (N_42504,N_42112,N_42458);
and U42505 (N_42505,N_42102,N_42141);
and U42506 (N_42506,N_42079,N_42245);
or U42507 (N_42507,N_42020,N_42086);
nand U42508 (N_42508,N_42137,N_42433);
nor U42509 (N_42509,N_42131,N_42121);
xnor U42510 (N_42510,N_42048,N_42468);
and U42511 (N_42511,N_42423,N_42134);
and U42512 (N_42512,N_42057,N_42015);
or U42513 (N_42513,N_42184,N_42139);
and U42514 (N_42514,N_42337,N_42041);
nor U42515 (N_42515,N_42461,N_42357);
and U42516 (N_42516,N_42013,N_42070);
nor U42517 (N_42517,N_42223,N_42331);
or U42518 (N_42518,N_42449,N_42353);
nand U42519 (N_42519,N_42267,N_42087);
and U42520 (N_42520,N_42474,N_42064);
nand U42521 (N_42521,N_42312,N_42333);
or U42522 (N_42522,N_42242,N_42281);
nand U42523 (N_42523,N_42192,N_42481);
nor U42524 (N_42524,N_42196,N_42219);
nand U42525 (N_42525,N_42185,N_42180);
nor U42526 (N_42526,N_42332,N_42172);
nor U42527 (N_42527,N_42347,N_42258);
nand U42528 (N_42528,N_42417,N_42151);
nand U42529 (N_42529,N_42301,N_42021);
xor U42530 (N_42530,N_42165,N_42148);
nor U42531 (N_42531,N_42026,N_42201);
and U42532 (N_42532,N_42138,N_42149);
nand U42533 (N_42533,N_42288,N_42170);
and U42534 (N_42534,N_42345,N_42169);
and U42535 (N_42535,N_42231,N_42044);
or U42536 (N_42536,N_42429,N_42297);
xnor U42537 (N_42537,N_42107,N_42421);
nor U42538 (N_42538,N_42212,N_42430);
nor U42539 (N_42539,N_42375,N_42336);
nand U42540 (N_42540,N_42025,N_42038);
nor U42541 (N_42541,N_42241,N_42240);
nor U42542 (N_42542,N_42164,N_42125);
and U42543 (N_42543,N_42406,N_42418);
nand U42544 (N_42544,N_42454,N_42456);
nand U42545 (N_42545,N_42318,N_42147);
or U42546 (N_42546,N_42052,N_42450);
nor U42547 (N_42547,N_42338,N_42105);
nor U42548 (N_42548,N_42214,N_42284);
and U42549 (N_42549,N_42156,N_42043);
or U42550 (N_42550,N_42253,N_42455);
and U42551 (N_42551,N_42055,N_42329);
nor U42552 (N_42552,N_42202,N_42111);
nor U42553 (N_42553,N_42003,N_42362);
or U42554 (N_42554,N_42399,N_42308);
nand U42555 (N_42555,N_42120,N_42166);
or U42556 (N_42556,N_42190,N_42388);
and U42557 (N_42557,N_42067,N_42299);
and U42558 (N_42558,N_42422,N_42259);
nor U42559 (N_42559,N_42191,N_42311);
and U42560 (N_42560,N_42247,N_42459);
nor U42561 (N_42561,N_42255,N_42088);
or U42562 (N_42562,N_42391,N_42019);
and U42563 (N_42563,N_42271,N_42280);
and U42564 (N_42564,N_42179,N_42061);
or U42565 (N_42565,N_42118,N_42486);
and U42566 (N_42566,N_42465,N_42478);
xor U42567 (N_42567,N_42173,N_42466);
xnor U42568 (N_42568,N_42194,N_42414);
nand U42569 (N_42569,N_42319,N_42424);
or U42570 (N_42570,N_42252,N_42434);
and U42571 (N_42571,N_42250,N_42436);
nor U42572 (N_42572,N_42005,N_42126);
and U42573 (N_42573,N_42389,N_42370);
or U42574 (N_42574,N_42416,N_42049);
nand U42575 (N_42575,N_42000,N_42496);
or U42576 (N_42576,N_42053,N_42144);
or U42577 (N_42577,N_42036,N_42227);
or U42578 (N_42578,N_42060,N_42428);
and U42579 (N_42579,N_42217,N_42328);
or U42580 (N_42580,N_42097,N_42359);
nand U42581 (N_42581,N_42243,N_42136);
nor U42582 (N_42582,N_42146,N_42195);
and U42583 (N_42583,N_42292,N_42076);
xor U42584 (N_42584,N_42492,N_42122);
nand U42585 (N_42585,N_42398,N_42443);
nand U42586 (N_42586,N_42282,N_42068);
or U42587 (N_42587,N_42104,N_42249);
nand U42588 (N_42588,N_42283,N_42404);
nor U42589 (N_42589,N_42346,N_42472);
nor U42590 (N_42590,N_42343,N_42094);
and U42591 (N_42591,N_42409,N_42489);
nand U42592 (N_42592,N_42106,N_42274);
and U42593 (N_42593,N_42029,N_42339);
and U42594 (N_42594,N_42316,N_42369);
nor U42595 (N_42595,N_42206,N_42056);
nand U42596 (N_42596,N_42011,N_42350);
nand U42597 (N_42597,N_42495,N_42322);
nand U42598 (N_42598,N_42415,N_42368);
and U42599 (N_42599,N_42213,N_42177);
nand U42600 (N_42600,N_42168,N_42033);
and U42601 (N_42601,N_42354,N_42300);
xnor U42602 (N_42602,N_42309,N_42188);
nand U42603 (N_42603,N_42447,N_42018);
and U42604 (N_42604,N_42108,N_42098);
or U42605 (N_42605,N_42065,N_42074);
and U42606 (N_42606,N_42187,N_42427);
nand U42607 (N_42607,N_42341,N_42420);
or U42608 (N_42608,N_42066,N_42358);
and U42609 (N_42609,N_42432,N_42497);
nand U42610 (N_42610,N_42470,N_42419);
and U42611 (N_42611,N_42393,N_42487);
nor U42612 (N_42612,N_42035,N_42440);
and U42613 (N_42613,N_42275,N_42103);
xnor U42614 (N_42614,N_42411,N_42027);
nand U42615 (N_42615,N_42342,N_42451);
xnor U42616 (N_42616,N_42225,N_42031);
and U42617 (N_42617,N_42040,N_42367);
or U42618 (N_42618,N_42475,N_42073);
or U42619 (N_42619,N_42349,N_42467);
nand U42620 (N_42620,N_42412,N_42374);
nand U42621 (N_42621,N_42330,N_42163);
or U42622 (N_42622,N_42364,N_42115);
or U42623 (N_42623,N_42310,N_42386);
and U42624 (N_42624,N_42162,N_42384);
or U42625 (N_42625,N_42260,N_42317);
or U42626 (N_42626,N_42326,N_42083);
nand U42627 (N_42627,N_42128,N_42324);
or U42628 (N_42628,N_42046,N_42473);
or U42629 (N_42629,N_42235,N_42376);
or U42630 (N_42630,N_42493,N_42238);
nor U42631 (N_42631,N_42340,N_42334);
nor U42632 (N_42632,N_42426,N_42269);
nand U42633 (N_42633,N_42007,N_42085);
and U42634 (N_42634,N_42159,N_42488);
or U42635 (N_42635,N_42452,N_42477);
or U42636 (N_42636,N_42186,N_42387);
nor U42637 (N_42637,N_42377,N_42279);
or U42638 (N_42638,N_42378,N_42008);
and U42639 (N_42639,N_42032,N_42209);
nor U42640 (N_42640,N_42207,N_42059);
nor U42641 (N_42641,N_42246,N_42482);
nor U42642 (N_42642,N_42265,N_42262);
nand U42643 (N_42643,N_42167,N_42327);
and U42644 (N_42644,N_42444,N_42273);
and U42645 (N_42645,N_42261,N_42101);
nand U42646 (N_42646,N_42010,N_42251);
nand U42647 (N_42647,N_42448,N_42323);
xnor U42648 (N_42648,N_42145,N_42197);
or U42649 (N_42649,N_42069,N_42153);
nor U42650 (N_42650,N_42286,N_42045);
nand U42651 (N_42651,N_42017,N_42290);
nand U42652 (N_42652,N_42022,N_42095);
or U42653 (N_42653,N_42285,N_42483);
and U42654 (N_42654,N_42355,N_42124);
xor U42655 (N_42655,N_42491,N_42132);
nor U42656 (N_42656,N_42200,N_42425);
and U42657 (N_42657,N_42437,N_42037);
or U42658 (N_42658,N_42266,N_42365);
and U42659 (N_42659,N_42325,N_42140);
xnor U42660 (N_42660,N_42127,N_42408);
nand U42661 (N_42661,N_42198,N_42445);
and U42662 (N_42662,N_42152,N_42257);
xor U42663 (N_42663,N_42012,N_42171);
or U42664 (N_42664,N_42226,N_42110);
and U42665 (N_42665,N_42075,N_42160);
xor U42666 (N_42666,N_42371,N_42222);
nor U42667 (N_42667,N_42158,N_42494);
or U42668 (N_42668,N_42228,N_42405);
and U42669 (N_42669,N_42157,N_42314);
xnor U42670 (N_42670,N_42092,N_42203);
or U42671 (N_42671,N_42183,N_42089);
or U42672 (N_42672,N_42034,N_42485);
and U42673 (N_42673,N_42116,N_42302);
or U42674 (N_42674,N_42397,N_42480);
xnor U42675 (N_42675,N_42264,N_42016);
and U42676 (N_42676,N_42352,N_42239);
nand U42677 (N_42677,N_42154,N_42174);
xor U42678 (N_42678,N_42220,N_42460);
nand U42679 (N_42679,N_42082,N_42024);
nor U42680 (N_42680,N_42360,N_42028);
nand U42681 (N_42681,N_42051,N_42023);
xor U42682 (N_42682,N_42351,N_42210);
nand U42683 (N_42683,N_42078,N_42155);
nor U42684 (N_42684,N_42438,N_42109);
xnor U42685 (N_42685,N_42077,N_42268);
nor U42686 (N_42686,N_42390,N_42096);
or U42687 (N_42687,N_42100,N_42009);
or U42688 (N_42688,N_42402,N_42462);
and U42689 (N_42689,N_42244,N_42001);
nor U42690 (N_42690,N_42143,N_42072);
nor U42691 (N_42691,N_42150,N_42410);
nor U42692 (N_42692,N_42401,N_42395);
and U42693 (N_42693,N_42315,N_42313);
and U42694 (N_42694,N_42320,N_42366);
nand U42695 (N_42695,N_42361,N_42230);
nand U42696 (N_42696,N_42081,N_42348);
and U42697 (N_42697,N_42381,N_42063);
or U42698 (N_42698,N_42403,N_42091);
xor U42699 (N_42699,N_42129,N_42270);
or U42700 (N_42700,N_42205,N_42394);
nor U42701 (N_42701,N_42123,N_42004);
and U42702 (N_42702,N_42431,N_42062);
and U42703 (N_42703,N_42090,N_42484);
nor U42704 (N_42704,N_42218,N_42221);
xnor U42705 (N_42705,N_42093,N_42385);
and U42706 (N_42706,N_42463,N_42498);
or U42707 (N_42707,N_42291,N_42236);
or U42708 (N_42708,N_42050,N_42379);
xnor U42709 (N_42709,N_42373,N_42303);
xnor U42710 (N_42710,N_42175,N_42383);
xor U42711 (N_42711,N_42396,N_42142);
xnor U42712 (N_42712,N_42471,N_42296);
and U42713 (N_42713,N_42133,N_42479);
nand U42714 (N_42714,N_42356,N_42435);
nand U42715 (N_42715,N_42298,N_42234);
xor U42716 (N_42716,N_42211,N_42071);
and U42717 (N_42717,N_42272,N_42135);
and U42718 (N_42718,N_42446,N_42130);
nor U42719 (N_42719,N_42117,N_42400);
nand U42720 (N_42720,N_42439,N_42321);
or U42721 (N_42721,N_42304,N_42042);
or U42722 (N_42722,N_42453,N_42006);
nand U42723 (N_42723,N_42248,N_42469);
or U42724 (N_42724,N_42215,N_42182);
nand U42725 (N_42725,N_42382,N_42476);
xnor U42726 (N_42726,N_42002,N_42084);
nor U42727 (N_42727,N_42229,N_42306);
and U42728 (N_42728,N_42161,N_42256);
nor U42729 (N_42729,N_42047,N_42464);
nand U42730 (N_42730,N_42499,N_42294);
or U42731 (N_42731,N_42233,N_42441);
and U42732 (N_42732,N_42232,N_42363);
nand U42733 (N_42733,N_42181,N_42014);
or U42734 (N_42734,N_42413,N_42176);
or U42735 (N_42735,N_42080,N_42287);
or U42736 (N_42736,N_42113,N_42490);
or U42737 (N_42737,N_42039,N_42276);
nor U42738 (N_42738,N_42099,N_42392);
nor U42739 (N_42739,N_42263,N_42224);
and U42740 (N_42740,N_42054,N_42305);
nand U42741 (N_42741,N_42119,N_42277);
xor U42742 (N_42742,N_42307,N_42216);
nor U42743 (N_42743,N_42372,N_42293);
or U42744 (N_42744,N_42278,N_42457);
nand U42745 (N_42745,N_42254,N_42380);
nand U42746 (N_42746,N_42193,N_42407);
and U42747 (N_42747,N_42178,N_42030);
or U42748 (N_42748,N_42199,N_42344);
or U42749 (N_42749,N_42289,N_42208);
and U42750 (N_42750,N_42207,N_42031);
and U42751 (N_42751,N_42023,N_42360);
and U42752 (N_42752,N_42126,N_42364);
xnor U42753 (N_42753,N_42122,N_42036);
nand U42754 (N_42754,N_42015,N_42433);
or U42755 (N_42755,N_42190,N_42077);
and U42756 (N_42756,N_42174,N_42255);
nor U42757 (N_42757,N_42088,N_42263);
and U42758 (N_42758,N_42276,N_42349);
nand U42759 (N_42759,N_42002,N_42387);
nand U42760 (N_42760,N_42369,N_42014);
or U42761 (N_42761,N_42167,N_42130);
nor U42762 (N_42762,N_42484,N_42219);
and U42763 (N_42763,N_42132,N_42308);
and U42764 (N_42764,N_42139,N_42439);
nand U42765 (N_42765,N_42127,N_42052);
nor U42766 (N_42766,N_42070,N_42393);
and U42767 (N_42767,N_42103,N_42137);
nor U42768 (N_42768,N_42421,N_42023);
nand U42769 (N_42769,N_42380,N_42423);
nor U42770 (N_42770,N_42059,N_42426);
and U42771 (N_42771,N_42372,N_42297);
nor U42772 (N_42772,N_42164,N_42329);
and U42773 (N_42773,N_42177,N_42471);
nand U42774 (N_42774,N_42146,N_42314);
nor U42775 (N_42775,N_42220,N_42357);
and U42776 (N_42776,N_42112,N_42412);
or U42777 (N_42777,N_42423,N_42137);
or U42778 (N_42778,N_42175,N_42205);
and U42779 (N_42779,N_42116,N_42212);
nand U42780 (N_42780,N_42158,N_42294);
and U42781 (N_42781,N_42412,N_42024);
and U42782 (N_42782,N_42305,N_42072);
or U42783 (N_42783,N_42288,N_42110);
and U42784 (N_42784,N_42266,N_42414);
nor U42785 (N_42785,N_42034,N_42285);
nor U42786 (N_42786,N_42014,N_42194);
nor U42787 (N_42787,N_42087,N_42061);
and U42788 (N_42788,N_42170,N_42360);
and U42789 (N_42789,N_42036,N_42273);
and U42790 (N_42790,N_42062,N_42139);
and U42791 (N_42791,N_42154,N_42075);
nor U42792 (N_42792,N_42240,N_42273);
nor U42793 (N_42793,N_42396,N_42091);
nand U42794 (N_42794,N_42431,N_42348);
nor U42795 (N_42795,N_42407,N_42470);
or U42796 (N_42796,N_42141,N_42292);
and U42797 (N_42797,N_42140,N_42421);
nor U42798 (N_42798,N_42054,N_42260);
and U42799 (N_42799,N_42161,N_42203);
nand U42800 (N_42800,N_42299,N_42103);
or U42801 (N_42801,N_42019,N_42228);
nand U42802 (N_42802,N_42147,N_42084);
and U42803 (N_42803,N_42108,N_42102);
and U42804 (N_42804,N_42433,N_42272);
nor U42805 (N_42805,N_42343,N_42171);
and U42806 (N_42806,N_42130,N_42113);
nor U42807 (N_42807,N_42063,N_42244);
xnor U42808 (N_42808,N_42030,N_42283);
and U42809 (N_42809,N_42020,N_42120);
nor U42810 (N_42810,N_42236,N_42229);
nor U42811 (N_42811,N_42033,N_42374);
nor U42812 (N_42812,N_42117,N_42115);
xor U42813 (N_42813,N_42274,N_42356);
nor U42814 (N_42814,N_42195,N_42436);
nand U42815 (N_42815,N_42189,N_42407);
or U42816 (N_42816,N_42156,N_42245);
or U42817 (N_42817,N_42192,N_42161);
nor U42818 (N_42818,N_42178,N_42210);
nor U42819 (N_42819,N_42414,N_42052);
nor U42820 (N_42820,N_42243,N_42025);
or U42821 (N_42821,N_42336,N_42052);
and U42822 (N_42822,N_42153,N_42173);
nor U42823 (N_42823,N_42193,N_42489);
nand U42824 (N_42824,N_42061,N_42465);
or U42825 (N_42825,N_42031,N_42096);
or U42826 (N_42826,N_42184,N_42382);
xor U42827 (N_42827,N_42213,N_42463);
or U42828 (N_42828,N_42057,N_42497);
nand U42829 (N_42829,N_42261,N_42190);
or U42830 (N_42830,N_42004,N_42317);
xor U42831 (N_42831,N_42490,N_42166);
xor U42832 (N_42832,N_42431,N_42439);
xnor U42833 (N_42833,N_42121,N_42220);
nor U42834 (N_42834,N_42409,N_42019);
xnor U42835 (N_42835,N_42031,N_42300);
nor U42836 (N_42836,N_42279,N_42042);
nor U42837 (N_42837,N_42494,N_42254);
nor U42838 (N_42838,N_42281,N_42448);
nor U42839 (N_42839,N_42066,N_42328);
nand U42840 (N_42840,N_42304,N_42355);
and U42841 (N_42841,N_42077,N_42335);
xnor U42842 (N_42842,N_42135,N_42228);
and U42843 (N_42843,N_42206,N_42373);
xnor U42844 (N_42844,N_42404,N_42013);
or U42845 (N_42845,N_42206,N_42195);
nor U42846 (N_42846,N_42255,N_42041);
and U42847 (N_42847,N_42281,N_42129);
nor U42848 (N_42848,N_42314,N_42282);
xor U42849 (N_42849,N_42233,N_42278);
nand U42850 (N_42850,N_42351,N_42450);
nor U42851 (N_42851,N_42272,N_42484);
or U42852 (N_42852,N_42481,N_42154);
xnor U42853 (N_42853,N_42272,N_42362);
and U42854 (N_42854,N_42302,N_42157);
nand U42855 (N_42855,N_42078,N_42172);
and U42856 (N_42856,N_42366,N_42398);
nor U42857 (N_42857,N_42231,N_42065);
and U42858 (N_42858,N_42251,N_42121);
nor U42859 (N_42859,N_42171,N_42458);
nand U42860 (N_42860,N_42287,N_42139);
xor U42861 (N_42861,N_42420,N_42372);
nand U42862 (N_42862,N_42072,N_42362);
and U42863 (N_42863,N_42165,N_42145);
or U42864 (N_42864,N_42087,N_42443);
and U42865 (N_42865,N_42049,N_42261);
nand U42866 (N_42866,N_42349,N_42370);
nand U42867 (N_42867,N_42208,N_42013);
and U42868 (N_42868,N_42497,N_42142);
xor U42869 (N_42869,N_42486,N_42229);
nor U42870 (N_42870,N_42279,N_42062);
nand U42871 (N_42871,N_42346,N_42381);
nand U42872 (N_42872,N_42185,N_42365);
or U42873 (N_42873,N_42475,N_42455);
or U42874 (N_42874,N_42322,N_42026);
nor U42875 (N_42875,N_42020,N_42018);
nand U42876 (N_42876,N_42301,N_42251);
nand U42877 (N_42877,N_42086,N_42092);
nor U42878 (N_42878,N_42415,N_42135);
xor U42879 (N_42879,N_42104,N_42330);
nor U42880 (N_42880,N_42194,N_42368);
nand U42881 (N_42881,N_42383,N_42353);
nor U42882 (N_42882,N_42421,N_42244);
nor U42883 (N_42883,N_42092,N_42087);
or U42884 (N_42884,N_42199,N_42188);
nor U42885 (N_42885,N_42378,N_42284);
or U42886 (N_42886,N_42311,N_42137);
nor U42887 (N_42887,N_42183,N_42016);
nor U42888 (N_42888,N_42161,N_42354);
or U42889 (N_42889,N_42277,N_42065);
nor U42890 (N_42890,N_42141,N_42200);
xor U42891 (N_42891,N_42257,N_42107);
nor U42892 (N_42892,N_42161,N_42134);
nor U42893 (N_42893,N_42177,N_42200);
nor U42894 (N_42894,N_42155,N_42405);
nand U42895 (N_42895,N_42334,N_42335);
nand U42896 (N_42896,N_42141,N_42470);
and U42897 (N_42897,N_42089,N_42429);
xor U42898 (N_42898,N_42116,N_42182);
nor U42899 (N_42899,N_42224,N_42442);
and U42900 (N_42900,N_42485,N_42442);
nor U42901 (N_42901,N_42480,N_42287);
or U42902 (N_42902,N_42218,N_42183);
and U42903 (N_42903,N_42185,N_42478);
and U42904 (N_42904,N_42241,N_42242);
or U42905 (N_42905,N_42382,N_42319);
or U42906 (N_42906,N_42378,N_42063);
xnor U42907 (N_42907,N_42022,N_42226);
or U42908 (N_42908,N_42489,N_42320);
nand U42909 (N_42909,N_42337,N_42480);
nand U42910 (N_42910,N_42327,N_42403);
nor U42911 (N_42911,N_42193,N_42154);
nor U42912 (N_42912,N_42244,N_42161);
nand U42913 (N_42913,N_42006,N_42409);
nand U42914 (N_42914,N_42306,N_42043);
and U42915 (N_42915,N_42096,N_42049);
and U42916 (N_42916,N_42337,N_42466);
nor U42917 (N_42917,N_42323,N_42210);
and U42918 (N_42918,N_42383,N_42168);
or U42919 (N_42919,N_42074,N_42299);
xnor U42920 (N_42920,N_42155,N_42249);
nand U42921 (N_42921,N_42432,N_42029);
and U42922 (N_42922,N_42282,N_42334);
xor U42923 (N_42923,N_42102,N_42183);
nand U42924 (N_42924,N_42410,N_42016);
xor U42925 (N_42925,N_42432,N_42253);
nand U42926 (N_42926,N_42490,N_42243);
nand U42927 (N_42927,N_42167,N_42038);
and U42928 (N_42928,N_42361,N_42259);
or U42929 (N_42929,N_42153,N_42498);
or U42930 (N_42930,N_42018,N_42078);
nor U42931 (N_42931,N_42116,N_42260);
nand U42932 (N_42932,N_42036,N_42405);
and U42933 (N_42933,N_42228,N_42209);
or U42934 (N_42934,N_42266,N_42378);
and U42935 (N_42935,N_42347,N_42317);
nand U42936 (N_42936,N_42265,N_42089);
and U42937 (N_42937,N_42483,N_42046);
and U42938 (N_42938,N_42348,N_42215);
nor U42939 (N_42939,N_42226,N_42005);
or U42940 (N_42940,N_42096,N_42452);
nor U42941 (N_42941,N_42488,N_42069);
or U42942 (N_42942,N_42472,N_42214);
or U42943 (N_42943,N_42487,N_42332);
or U42944 (N_42944,N_42471,N_42181);
nand U42945 (N_42945,N_42408,N_42103);
nand U42946 (N_42946,N_42307,N_42023);
xor U42947 (N_42947,N_42214,N_42286);
or U42948 (N_42948,N_42185,N_42292);
nor U42949 (N_42949,N_42458,N_42131);
and U42950 (N_42950,N_42262,N_42349);
nand U42951 (N_42951,N_42368,N_42459);
nand U42952 (N_42952,N_42498,N_42080);
and U42953 (N_42953,N_42303,N_42108);
and U42954 (N_42954,N_42452,N_42074);
and U42955 (N_42955,N_42047,N_42350);
nand U42956 (N_42956,N_42038,N_42227);
nor U42957 (N_42957,N_42273,N_42152);
or U42958 (N_42958,N_42385,N_42106);
or U42959 (N_42959,N_42109,N_42128);
and U42960 (N_42960,N_42442,N_42128);
and U42961 (N_42961,N_42145,N_42240);
or U42962 (N_42962,N_42489,N_42455);
nor U42963 (N_42963,N_42106,N_42152);
or U42964 (N_42964,N_42315,N_42215);
nor U42965 (N_42965,N_42410,N_42070);
nor U42966 (N_42966,N_42205,N_42471);
or U42967 (N_42967,N_42187,N_42278);
xnor U42968 (N_42968,N_42187,N_42174);
or U42969 (N_42969,N_42432,N_42422);
and U42970 (N_42970,N_42071,N_42274);
xnor U42971 (N_42971,N_42035,N_42183);
and U42972 (N_42972,N_42046,N_42184);
or U42973 (N_42973,N_42221,N_42092);
or U42974 (N_42974,N_42261,N_42152);
nand U42975 (N_42975,N_42059,N_42429);
nor U42976 (N_42976,N_42265,N_42088);
or U42977 (N_42977,N_42345,N_42272);
nand U42978 (N_42978,N_42090,N_42210);
nand U42979 (N_42979,N_42358,N_42412);
nand U42980 (N_42980,N_42463,N_42403);
or U42981 (N_42981,N_42210,N_42293);
xor U42982 (N_42982,N_42278,N_42104);
nand U42983 (N_42983,N_42086,N_42152);
nor U42984 (N_42984,N_42229,N_42012);
nand U42985 (N_42985,N_42343,N_42349);
nor U42986 (N_42986,N_42265,N_42438);
nand U42987 (N_42987,N_42206,N_42072);
nand U42988 (N_42988,N_42489,N_42262);
xor U42989 (N_42989,N_42251,N_42283);
and U42990 (N_42990,N_42014,N_42053);
nand U42991 (N_42991,N_42363,N_42266);
nand U42992 (N_42992,N_42206,N_42066);
and U42993 (N_42993,N_42012,N_42019);
and U42994 (N_42994,N_42037,N_42091);
or U42995 (N_42995,N_42367,N_42264);
and U42996 (N_42996,N_42319,N_42096);
nand U42997 (N_42997,N_42330,N_42458);
or U42998 (N_42998,N_42090,N_42456);
and U42999 (N_42999,N_42396,N_42436);
nor U43000 (N_43000,N_42797,N_42579);
and U43001 (N_43001,N_42836,N_42621);
xor U43002 (N_43002,N_42824,N_42918);
and U43003 (N_43003,N_42605,N_42973);
nor U43004 (N_43004,N_42891,N_42720);
or U43005 (N_43005,N_42966,N_42670);
nand U43006 (N_43006,N_42808,N_42627);
xnor U43007 (N_43007,N_42877,N_42513);
nand U43008 (N_43008,N_42777,N_42613);
or U43009 (N_43009,N_42828,N_42640);
or U43010 (N_43010,N_42965,N_42994);
nand U43011 (N_43011,N_42886,N_42521);
nor U43012 (N_43012,N_42747,N_42721);
nand U43013 (N_43013,N_42666,N_42634);
nor U43014 (N_43014,N_42664,N_42970);
nand U43015 (N_43015,N_42568,N_42599);
nor U43016 (N_43016,N_42617,N_42844);
or U43017 (N_43017,N_42745,N_42984);
nand U43018 (N_43018,N_42971,N_42875);
nand U43019 (N_43019,N_42782,N_42942);
or U43020 (N_43020,N_42868,N_42962);
or U43021 (N_43021,N_42622,N_42712);
nor U43022 (N_43022,N_42692,N_42762);
nand U43023 (N_43023,N_42818,N_42563);
nand U43024 (N_43024,N_42688,N_42826);
nand U43025 (N_43025,N_42660,N_42803);
nand U43026 (N_43026,N_42776,N_42752);
nand U43027 (N_43027,N_42872,N_42561);
or U43028 (N_43028,N_42644,N_42933);
or U43029 (N_43029,N_42509,N_42765);
nor U43030 (N_43030,N_42880,N_42545);
or U43031 (N_43031,N_42645,N_42680);
nor U43032 (N_43032,N_42620,N_42811);
nand U43033 (N_43033,N_42806,N_42921);
nand U43034 (N_43034,N_42998,N_42780);
nand U43035 (N_43035,N_42618,N_42691);
or U43036 (N_43036,N_42746,N_42841);
nand U43037 (N_43037,N_42584,N_42676);
nand U43038 (N_43038,N_42739,N_42560);
xnor U43039 (N_43039,N_42591,N_42772);
xor U43040 (N_43040,N_42592,N_42631);
or U43041 (N_43041,N_42802,N_42922);
or U43042 (N_43042,N_42825,N_42601);
and U43043 (N_43043,N_42732,N_42514);
nand U43044 (N_43044,N_42536,N_42804);
nor U43045 (N_43045,N_42959,N_42517);
nand U43046 (N_43046,N_42682,N_42717);
and U43047 (N_43047,N_42566,N_42755);
nand U43048 (N_43048,N_42650,N_42558);
nor U43049 (N_43049,N_42871,N_42763);
or U43050 (N_43050,N_42928,N_42914);
and U43051 (N_43051,N_42540,N_42958);
nor U43052 (N_43052,N_42529,N_42503);
or U43053 (N_43053,N_42524,N_42799);
and U43054 (N_43054,N_42667,N_42787);
or U43055 (N_43055,N_42541,N_42904);
or U43056 (N_43056,N_42699,N_42674);
nand U43057 (N_43057,N_42654,N_42955);
xnor U43058 (N_43058,N_42805,N_42862);
or U43059 (N_43059,N_42728,N_42507);
and U43060 (N_43060,N_42542,N_42646);
nor U43061 (N_43061,N_42576,N_42757);
nor U43062 (N_43062,N_42936,N_42741);
and U43063 (N_43063,N_42539,N_42953);
nor U43064 (N_43064,N_42833,N_42581);
and U43065 (N_43065,N_42882,N_42684);
and U43066 (N_43066,N_42945,N_42768);
and U43067 (N_43067,N_42870,N_42593);
and U43068 (N_43068,N_42547,N_42504);
nand U43069 (N_43069,N_42832,N_42719);
xor U43070 (N_43070,N_42960,N_42625);
or U43071 (N_43071,N_42711,N_42678);
nand U43072 (N_43072,N_42864,N_42830);
and U43073 (N_43073,N_42683,N_42764);
nor U43074 (N_43074,N_42855,N_42642);
nor U43075 (N_43075,N_42885,N_42919);
nand U43076 (N_43076,N_42759,N_42733);
xor U43077 (N_43077,N_42927,N_42743);
xnor U43078 (N_43078,N_42651,N_42929);
nand U43079 (N_43079,N_42907,N_42569);
and U43080 (N_43080,N_42594,N_42750);
or U43081 (N_43081,N_42520,N_42814);
or U43082 (N_43082,N_42989,N_42532);
or U43083 (N_43083,N_42573,N_42730);
and U43084 (N_43084,N_42500,N_42952);
nor U43085 (N_43085,N_42744,N_42923);
and U43086 (N_43086,N_42990,N_42845);
nand U43087 (N_43087,N_42546,N_42794);
nor U43088 (N_43088,N_42789,N_42713);
or U43089 (N_43089,N_42636,N_42821);
and U43090 (N_43090,N_42829,N_42858);
nand U43091 (N_43091,N_42901,N_42810);
xnor U43092 (N_43092,N_42624,N_42781);
or U43093 (N_43093,N_42761,N_42550);
or U43094 (N_43094,N_42552,N_42876);
and U43095 (N_43095,N_42838,N_42586);
nand U43096 (N_43096,N_42548,N_42944);
xor U43097 (N_43097,N_42724,N_42641);
xor U43098 (N_43098,N_42567,N_42917);
nand U43099 (N_43099,N_42846,N_42512);
or U43100 (N_43100,N_42587,N_42769);
nand U43101 (N_43101,N_42849,N_42900);
nand U43102 (N_43102,N_42979,N_42537);
nand U43103 (N_43103,N_42506,N_42510);
or U43104 (N_43104,N_42898,N_42515);
nand U43105 (N_43105,N_42822,N_42600);
xor U43106 (N_43106,N_42656,N_42502);
or U43107 (N_43107,N_42616,N_42854);
xor U43108 (N_43108,N_42954,N_42975);
nor U43109 (N_43109,N_42638,N_42931);
or U43110 (N_43110,N_42580,N_42530);
nand U43111 (N_43111,N_42926,N_42675);
nand U43112 (N_43112,N_42707,N_42796);
nor U43113 (N_43113,N_42767,N_42939);
nand U43114 (N_43114,N_42588,N_42735);
nand U43115 (N_43115,N_42977,N_42816);
or U43116 (N_43116,N_42597,N_42582);
nor U43117 (N_43117,N_42800,N_42890);
xor U43118 (N_43118,N_42749,N_42525);
and U43119 (N_43119,N_42710,N_42701);
nand U43120 (N_43120,N_42974,N_42982);
and U43121 (N_43121,N_42635,N_42551);
nor U43122 (N_43122,N_42623,N_42834);
nor U43123 (N_43123,N_42788,N_42689);
nand U43124 (N_43124,N_42867,N_42538);
xnor U43125 (N_43125,N_42756,N_42912);
nand U43126 (N_43126,N_42827,N_42686);
nand U43127 (N_43127,N_42941,N_42861);
xor U43128 (N_43128,N_42511,N_42714);
nor U43129 (N_43129,N_42610,N_42925);
nor U43130 (N_43130,N_42673,N_42878);
and U43131 (N_43131,N_42869,N_42629);
or U43132 (N_43132,N_42798,N_42595);
nand U43133 (N_43133,N_42578,N_42531);
and U43134 (N_43134,N_42813,N_42725);
nand U43135 (N_43135,N_42742,N_42700);
nand U43136 (N_43136,N_42708,N_42961);
or U43137 (N_43137,N_42779,N_42856);
and U43138 (N_43138,N_42771,N_42791);
nor U43139 (N_43139,N_42612,N_42737);
and U43140 (N_43140,N_42718,N_42848);
nor U43141 (N_43141,N_42895,N_42934);
nand U43142 (N_43142,N_42685,N_42792);
and U43143 (N_43143,N_42793,N_42723);
nand U43144 (N_43144,N_42948,N_42554);
nor U43145 (N_43145,N_42709,N_42949);
nor U43146 (N_43146,N_42785,N_42703);
and U43147 (N_43147,N_42694,N_42860);
nor U43148 (N_43148,N_42817,N_42562);
nand U43149 (N_43149,N_42611,N_42992);
and U43150 (N_43150,N_42614,N_42736);
and U43151 (N_43151,N_42956,N_42851);
nor U43152 (N_43152,N_42853,N_42863);
and U43153 (N_43153,N_42873,N_42639);
and U43154 (N_43154,N_42555,N_42697);
nand U43155 (N_43155,N_42659,N_42696);
or U43156 (N_43156,N_42596,N_42702);
nor U43157 (N_43157,N_42671,N_42894);
or U43158 (N_43158,N_42831,N_42715);
xor U43159 (N_43159,N_42658,N_42643);
xnor U43160 (N_43160,N_42859,N_42968);
or U43161 (N_43161,N_42501,N_42559);
or U43162 (N_43162,N_42910,N_42758);
or U43163 (N_43163,N_42839,N_42893);
and U43164 (N_43164,N_42690,N_42903);
or U43165 (N_43165,N_42556,N_42874);
nor U43166 (N_43166,N_42790,N_42572);
nor U43167 (N_43167,N_42522,N_42906);
and U43168 (N_43168,N_42980,N_42661);
or U43169 (N_43169,N_42987,N_42774);
nor U43170 (N_43170,N_42662,N_42693);
or U43171 (N_43171,N_42937,N_42812);
nand U43172 (N_43172,N_42571,N_42669);
nor U43173 (N_43173,N_42657,N_42991);
nor U43174 (N_43174,N_42534,N_42518);
and U43175 (N_43175,N_42698,N_42677);
or U43176 (N_43176,N_42823,N_42795);
nor U43177 (N_43177,N_42528,N_42920);
and U43178 (N_43178,N_42583,N_42896);
nor U43179 (N_43179,N_42883,N_42866);
nand U43180 (N_43180,N_42681,N_42967);
xnor U43181 (N_43181,N_42951,N_42783);
nor U43182 (N_43182,N_42647,N_42705);
or U43183 (N_43183,N_42716,N_42607);
nand U43184 (N_43184,N_42628,N_42653);
nor U43185 (N_43185,N_42663,N_42835);
nand U43186 (N_43186,N_42606,N_42760);
and U43187 (N_43187,N_42748,N_42574);
or U43188 (N_43188,N_42604,N_42753);
or U43189 (N_43189,N_42888,N_42523);
nor U43190 (N_43190,N_42649,N_42915);
and U43191 (N_43191,N_42519,N_42946);
nor U43192 (N_43192,N_42905,N_42972);
and U43193 (N_43193,N_42809,N_42902);
nor U43194 (N_43194,N_42751,N_42527);
and U43195 (N_43195,N_42985,N_42897);
nor U43196 (N_43196,N_42943,N_42516);
nand U43197 (N_43197,N_42801,N_42608);
or U43198 (N_43198,N_42996,N_42603);
and U43199 (N_43199,N_42932,N_42963);
nor U43200 (N_43200,N_42879,N_42577);
nand U43201 (N_43201,N_42981,N_42598);
nor U43202 (N_43202,N_42935,N_42526);
nand U43203 (N_43203,N_42731,N_42911);
and U43204 (N_43204,N_42766,N_42999);
or U43205 (N_43205,N_42820,N_42544);
nand U43206 (N_43206,N_42722,N_42609);
nand U43207 (N_43207,N_42983,N_42807);
or U43208 (N_43208,N_42754,N_42899);
and U43209 (N_43209,N_42957,N_42652);
and U43210 (N_43210,N_42770,N_42857);
and U43211 (N_43211,N_42575,N_42986);
nor U43212 (N_43212,N_42940,N_42726);
and U43213 (N_43213,N_42729,N_42619);
xnor U43214 (N_43214,N_42837,N_42589);
and U43215 (N_43215,N_42602,N_42993);
and U43216 (N_43216,N_42533,N_42727);
and U43217 (N_43217,N_42679,N_42687);
nor U43218 (N_43218,N_42924,N_42648);
nor U43219 (N_43219,N_42630,N_42976);
xor U43220 (N_43220,N_42889,N_42665);
or U43221 (N_43221,N_42543,N_42887);
nand U43222 (N_43222,N_42850,N_42978);
and U43223 (N_43223,N_42740,N_42775);
nor U43224 (N_43224,N_42508,N_42852);
nor U43225 (N_43225,N_42637,N_42842);
xnor U43226 (N_43226,N_42633,N_42913);
and U43227 (N_43227,N_42565,N_42570);
nand U43228 (N_43228,N_42930,N_42734);
nor U43229 (N_43229,N_42632,N_42892);
nand U43230 (N_43230,N_42615,N_42819);
nor U43231 (N_43231,N_42590,N_42997);
xor U43232 (N_43232,N_42964,N_42884);
or U43233 (N_43233,N_42995,N_42843);
or U43234 (N_43234,N_42695,N_42784);
xor U43235 (N_43235,N_42549,N_42668);
nand U43236 (N_43236,N_42778,N_42564);
and U43237 (N_43237,N_42557,N_42847);
nor U43238 (N_43238,N_42773,N_42881);
xnor U43239 (N_43239,N_42655,N_42950);
or U43240 (N_43240,N_42916,N_42865);
nand U43241 (N_43241,N_42738,N_42815);
and U43242 (N_43242,N_42947,N_42672);
and U43243 (N_43243,N_42505,N_42938);
and U43244 (N_43244,N_42840,N_42988);
nand U43245 (N_43245,N_42969,N_42706);
xnor U43246 (N_43246,N_42626,N_42786);
and U43247 (N_43247,N_42553,N_42908);
nor U43248 (N_43248,N_42535,N_42909);
nor U43249 (N_43249,N_42704,N_42585);
xor U43250 (N_43250,N_42706,N_42694);
xnor U43251 (N_43251,N_42558,N_42676);
nand U43252 (N_43252,N_42851,N_42776);
nor U43253 (N_43253,N_42600,N_42987);
xnor U43254 (N_43254,N_42548,N_42617);
nor U43255 (N_43255,N_42503,N_42537);
or U43256 (N_43256,N_42880,N_42802);
or U43257 (N_43257,N_42738,N_42549);
or U43258 (N_43258,N_42580,N_42551);
nand U43259 (N_43259,N_42767,N_42969);
and U43260 (N_43260,N_42645,N_42737);
or U43261 (N_43261,N_42503,N_42811);
and U43262 (N_43262,N_42568,N_42882);
or U43263 (N_43263,N_42676,N_42593);
nor U43264 (N_43264,N_42667,N_42577);
and U43265 (N_43265,N_42845,N_42719);
or U43266 (N_43266,N_42937,N_42711);
nor U43267 (N_43267,N_42715,N_42512);
xnor U43268 (N_43268,N_42574,N_42981);
nand U43269 (N_43269,N_42870,N_42571);
and U43270 (N_43270,N_42785,N_42884);
nor U43271 (N_43271,N_42870,N_42910);
nand U43272 (N_43272,N_42530,N_42587);
or U43273 (N_43273,N_42862,N_42753);
or U43274 (N_43274,N_42521,N_42621);
or U43275 (N_43275,N_42799,N_42804);
nor U43276 (N_43276,N_42809,N_42668);
nor U43277 (N_43277,N_42936,N_42542);
or U43278 (N_43278,N_42537,N_42788);
xor U43279 (N_43279,N_42922,N_42899);
nand U43280 (N_43280,N_42660,N_42729);
nor U43281 (N_43281,N_42839,N_42715);
and U43282 (N_43282,N_42834,N_42712);
xor U43283 (N_43283,N_42650,N_42789);
nand U43284 (N_43284,N_42535,N_42924);
xor U43285 (N_43285,N_42963,N_42572);
or U43286 (N_43286,N_42525,N_42868);
or U43287 (N_43287,N_42802,N_42580);
or U43288 (N_43288,N_42790,N_42893);
nand U43289 (N_43289,N_42726,N_42930);
xnor U43290 (N_43290,N_42676,N_42675);
nor U43291 (N_43291,N_42984,N_42916);
nor U43292 (N_43292,N_42999,N_42646);
or U43293 (N_43293,N_42929,N_42539);
nand U43294 (N_43294,N_42507,N_42950);
nor U43295 (N_43295,N_42804,N_42578);
xor U43296 (N_43296,N_42524,N_42601);
nor U43297 (N_43297,N_42819,N_42740);
xnor U43298 (N_43298,N_42539,N_42756);
nand U43299 (N_43299,N_42915,N_42644);
nand U43300 (N_43300,N_42917,N_42541);
nand U43301 (N_43301,N_42978,N_42765);
nor U43302 (N_43302,N_42789,N_42564);
nand U43303 (N_43303,N_42653,N_42635);
or U43304 (N_43304,N_42744,N_42582);
nor U43305 (N_43305,N_42691,N_42653);
and U43306 (N_43306,N_42782,N_42527);
nand U43307 (N_43307,N_42882,N_42849);
or U43308 (N_43308,N_42957,N_42556);
nor U43309 (N_43309,N_42845,N_42799);
and U43310 (N_43310,N_42972,N_42817);
nor U43311 (N_43311,N_42943,N_42728);
nand U43312 (N_43312,N_42519,N_42994);
and U43313 (N_43313,N_42622,N_42995);
and U43314 (N_43314,N_42858,N_42936);
xnor U43315 (N_43315,N_42829,N_42807);
or U43316 (N_43316,N_42854,N_42958);
and U43317 (N_43317,N_42567,N_42852);
nand U43318 (N_43318,N_42954,N_42642);
nand U43319 (N_43319,N_42983,N_42568);
and U43320 (N_43320,N_42707,N_42940);
or U43321 (N_43321,N_42721,N_42944);
nand U43322 (N_43322,N_42776,N_42741);
and U43323 (N_43323,N_42516,N_42687);
and U43324 (N_43324,N_42548,N_42872);
nor U43325 (N_43325,N_42578,N_42762);
or U43326 (N_43326,N_42730,N_42752);
and U43327 (N_43327,N_42939,N_42958);
nand U43328 (N_43328,N_42979,N_42554);
and U43329 (N_43329,N_42987,N_42527);
nor U43330 (N_43330,N_42711,N_42922);
nor U43331 (N_43331,N_42869,N_42503);
xnor U43332 (N_43332,N_42510,N_42738);
xnor U43333 (N_43333,N_42527,N_42920);
or U43334 (N_43334,N_42710,N_42684);
nor U43335 (N_43335,N_42615,N_42803);
and U43336 (N_43336,N_42717,N_42802);
or U43337 (N_43337,N_42902,N_42628);
nand U43338 (N_43338,N_42594,N_42511);
and U43339 (N_43339,N_42915,N_42586);
nand U43340 (N_43340,N_42770,N_42689);
nor U43341 (N_43341,N_42786,N_42756);
nor U43342 (N_43342,N_42580,N_42887);
or U43343 (N_43343,N_42544,N_42886);
nand U43344 (N_43344,N_42729,N_42852);
and U43345 (N_43345,N_42918,N_42706);
or U43346 (N_43346,N_42947,N_42686);
or U43347 (N_43347,N_42716,N_42635);
and U43348 (N_43348,N_42671,N_42648);
nor U43349 (N_43349,N_42664,N_42519);
or U43350 (N_43350,N_42985,N_42534);
xnor U43351 (N_43351,N_42987,N_42627);
xor U43352 (N_43352,N_42601,N_42567);
nor U43353 (N_43353,N_42852,N_42921);
nor U43354 (N_43354,N_42634,N_42805);
nand U43355 (N_43355,N_42779,N_42910);
nand U43356 (N_43356,N_42903,N_42615);
xor U43357 (N_43357,N_42941,N_42655);
and U43358 (N_43358,N_42848,N_42562);
and U43359 (N_43359,N_42865,N_42588);
and U43360 (N_43360,N_42572,N_42624);
nand U43361 (N_43361,N_42664,N_42851);
nand U43362 (N_43362,N_42798,N_42711);
xor U43363 (N_43363,N_42788,N_42573);
nand U43364 (N_43364,N_42746,N_42873);
nand U43365 (N_43365,N_42828,N_42829);
and U43366 (N_43366,N_42858,N_42764);
nor U43367 (N_43367,N_42934,N_42993);
nor U43368 (N_43368,N_42691,N_42646);
nor U43369 (N_43369,N_42786,N_42544);
nor U43370 (N_43370,N_42975,N_42515);
and U43371 (N_43371,N_42705,N_42868);
nor U43372 (N_43372,N_42565,N_42726);
or U43373 (N_43373,N_42727,N_42651);
xnor U43374 (N_43374,N_42830,N_42526);
nand U43375 (N_43375,N_42693,N_42638);
or U43376 (N_43376,N_42692,N_42727);
xnor U43377 (N_43377,N_42793,N_42975);
or U43378 (N_43378,N_42776,N_42945);
nand U43379 (N_43379,N_42738,N_42584);
or U43380 (N_43380,N_42946,N_42972);
nor U43381 (N_43381,N_42624,N_42712);
and U43382 (N_43382,N_42642,N_42699);
nand U43383 (N_43383,N_42662,N_42512);
or U43384 (N_43384,N_42518,N_42709);
nand U43385 (N_43385,N_42570,N_42734);
or U43386 (N_43386,N_42664,N_42814);
nor U43387 (N_43387,N_42961,N_42621);
and U43388 (N_43388,N_42560,N_42856);
nor U43389 (N_43389,N_42867,N_42721);
and U43390 (N_43390,N_42896,N_42704);
and U43391 (N_43391,N_42654,N_42777);
xor U43392 (N_43392,N_42799,N_42884);
and U43393 (N_43393,N_42942,N_42632);
nand U43394 (N_43394,N_42922,N_42510);
xor U43395 (N_43395,N_42872,N_42877);
and U43396 (N_43396,N_42882,N_42558);
nand U43397 (N_43397,N_42581,N_42518);
xor U43398 (N_43398,N_42517,N_42502);
and U43399 (N_43399,N_42716,N_42896);
xor U43400 (N_43400,N_42998,N_42816);
nor U43401 (N_43401,N_42849,N_42945);
nor U43402 (N_43402,N_42792,N_42684);
nor U43403 (N_43403,N_42973,N_42980);
nor U43404 (N_43404,N_42831,N_42540);
nor U43405 (N_43405,N_42765,N_42739);
nor U43406 (N_43406,N_42991,N_42809);
or U43407 (N_43407,N_42634,N_42564);
nand U43408 (N_43408,N_42929,N_42923);
nand U43409 (N_43409,N_42751,N_42836);
nor U43410 (N_43410,N_42521,N_42756);
xnor U43411 (N_43411,N_42754,N_42551);
and U43412 (N_43412,N_42682,N_42535);
nand U43413 (N_43413,N_42800,N_42946);
or U43414 (N_43414,N_42740,N_42774);
or U43415 (N_43415,N_42561,N_42591);
nor U43416 (N_43416,N_42716,N_42795);
nand U43417 (N_43417,N_42870,N_42902);
xor U43418 (N_43418,N_42774,N_42828);
nor U43419 (N_43419,N_42585,N_42672);
nor U43420 (N_43420,N_42801,N_42728);
xor U43421 (N_43421,N_42607,N_42728);
nand U43422 (N_43422,N_42861,N_42506);
nor U43423 (N_43423,N_42885,N_42524);
or U43424 (N_43424,N_42679,N_42572);
and U43425 (N_43425,N_42783,N_42944);
or U43426 (N_43426,N_42525,N_42625);
nor U43427 (N_43427,N_42701,N_42573);
or U43428 (N_43428,N_42969,N_42548);
or U43429 (N_43429,N_42903,N_42635);
or U43430 (N_43430,N_42824,N_42902);
and U43431 (N_43431,N_42913,N_42870);
or U43432 (N_43432,N_42595,N_42759);
nor U43433 (N_43433,N_42678,N_42563);
nand U43434 (N_43434,N_42838,N_42818);
and U43435 (N_43435,N_42872,N_42753);
or U43436 (N_43436,N_42747,N_42907);
and U43437 (N_43437,N_42534,N_42588);
or U43438 (N_43438,N_42999,N_42561);
nand U43439 (N_43439,N_42508,N_42912);
and U43440 (N_43440,N_42789,N_42550);
and U43441 (N_43441,N_42960,N_42684);
nand U43442 (N_43442,N_42519,N_42996);
or U43443 (N_43443,N_42897,N_42920);
or U43444 (N_43444,N_42962,N_42857);
or U43445 (N_43445,N_42508,N_42524);
and U43446 (N_43446,N_42719,N_42897);
or U43447 (N_43447,N_42698,N_42563);
and U43448 (N_43448,N_42819,N_42854);
xnor U43449 (N_43449,N_42673,N_42839);
nand U43450 (N_43450,N_42797,N_42974);
nand U43451 (N_43451,N_42620,N_42781);
nand U43452 (N_43452,N_42534,N_42851);
nand U43453 (N_43453,N_42515,N_42672);
nor U43454 (N_43454,N_42790,N_42842);
and U43455 (N_43455,N_42910,N_42588);
nand U43456 (N_43456,N_42523,N_42924);
nor U43457 (N_43457,N_42767,N_42661);
and U43458 (N_43458,N_42751,N_42564);
nand U43459 (N_43459,N_42941,N_42699);
and U43460 (N_43460,N_42611,N_42942);
nand U43461 (N_43461,N_42692,N_42594);
nor U43462 (N_43462,N_42711,N_42815);
nor U43463 (N_43463,N_42552,N_42609);
nor U43464 (N_43464,N_42735,N_42712);
and U43465 (N_43465,N_42558,N_42579);
nand U43466 (N_43466,N_42709,N_42838);
nor U43467 (N_43467,N_42671,N_42532);
or U43468 (N_43468,N_42916,N_42535);
nand U43469 (N_43469,N_42871,N_42583);
nor U43470 (N_43470,N_42849,N_42663);
nand U43471 (N_43471,N_42583,N_42861);
and U43472 (N_43472,N_42627,N_42535);
nand U43473 (N_43473,N_42609,N_42897);
and U43474 (N_43474,N_42594,N_42955);
and U43475 (N_43475,N_42973,N_42688);
nand U43476 (N_43476,N_42702,N_42683);
nor U43477 (N_43477,N_42560,N_42766);
or U43478 (N_43478,N_42521,N_42614);
and U43479 (N_43479,N_42627,N_42533);
nand U43480 (N_43480,N_42811,N_42949);
or U43481 (N_43481,N_42825,N_42554);
nor U43482 (N_43482,N_42607,N_42905);
xnor U43483 (N_43483,N_42744,N_42990);
xnor U43484 (N_43484,N_42513,N_42913);
xor U43485 (N_43485,N_42899,N_42895);
and U43486 (N_43486,N_42997,N_42976);
and U43487 (N_43487,N_42648,N_42668);
and U43488 (N_43488,N_42955,N_42871);
xnor U43489 (N_43489,N_42814,N_42504);
or U43490 (N_43490,N_42914,N_42868);
or U43491 (N_43491,N_42704,N_42904);
and U43492 (N_43492,N_42858,N_42684);
and U43493 (N_43493,N_42602,N_42606);
nor U43494 (N_43494,N_42835,N_42894);
and U43495 (N_43495,N_42834,N_42700);
nand U43496 (N_43496,N_42644,N_42611);
xnor U43497 (N_43497,N_42648,N_42950);
or U43498 (N_43498,N_42920,N_42523);
and U43499 (N_43499,N_42748,N_42553);
and U43500 (N_43500,N_43445,N_43259);
nand U43501 (N_43501,N_43085,N_43488);
nand U43502 (N_43502,N_43431,N_43385);
or U43503 (N_43503,N_43012,N_43243);
nor U43504 (N_43504,N_43163,N_43175);
or U43505 (N_43505,N_43348,N_43466);
and U43506 (N_43506,N_43467,N_43063);
nor U43507 (N_43507,N_43202,N_43160);
xor U43508 (N_43508,N_43275,N_43357);
xor U43509 (N_43509,N_43210,N_43475);
xnor U43510 (N_43510,N_43456,N_43271);
and U43511 (N_43511,N_43113,N_43123);
nor U43512 (N_43512,N_43036,N_43443);
nand U43513 (N_43513,N_43343,N_43109);
or U43514 (N_43514,N_43489,N_43070);
and U43515 (N_43515,N_43487,N_43222);
xor U43516 (N_43516,N_43016,N_43238);
and U43517 (N_43517,N_43153,N_43345);
and U43518 (N_43518,N_43252,N_43095);
nor U43519 (N_43519,N_43342,N_43365);
nand U43520 (N_43520,N_43239,N_43077);
and U43521 (N_43521,N_43082,N_43097);
nand U43522 (N_43522,N_43090,N_43376);
and U43523 (N_43523,N_43112,N_43284);
and U43524 (N_43524,N_43008,N_43439);
nor U43525 (N_43525,N_43178,N_43071);
nand U43526 (N_43526,N_43381,N_43476);
and U43527 (N_43527,N_43287,N_43330);
nand U43528 (N_43528,N_43293,N_43303);
and U43529 (N_43529,N_43069,N_43135);
and U43530 (N_43530,N_43392,N_43360);
nor U43531 (N_43531,N_43370,N_43413);
nand U43532 (N_43532,N_43223,N_43276);
nand U43533 (N_43533,N_43044,N_43025);
and U43534 (N_43534,N_43468,N_43408);
nand U43535 (N_43535,N_43384,N_43405);
nand U43536 (N_43536,N_43282,N_43083);
nand U43537 (N_43537,N_43427,N_43249);
nand U43538 (N_43538,N_43074,N_43010);
or U43539 (N_43539,N_43161,N_43213);
nor U43540 (N_43540,N_43358,N_43434);
nand U43541 (N_43541,N_43004,N_43087);
nor U43542 (N_43542,N_43079,N_43354);
and U43543 (N_43543,N_43349,N_43352);
nor U43544 (N_43544,N_43228,N_43084);
and U43545 (N_43545,N_43355,N_43438);
or U43546 (N_43546,N_43067,N_43286);
or U43547 (N_43547,N_43054,N_43493);
and U43548 (N_43548,N_43245,N_43347);
xnor U43549 (N_43549,N_43028,N_43191);
or U43550 (N_43550,N_43449,N_43435);
nand U43551 (N_43551,N_43143,N_43418);
or U43552 (N_43552,N_43061,N_43402);
and U43553 (N_43553,N_43041,N_43096);
nor U43554 (N_43554,N_43151,N_43369);
nor U43555 (N_43555,N_43133,N_43307);
nor U43556 (N_43556,N_43164,N_43207);
nor U43557 (N_43557,N_43062,N_43137);
nor U43558 (N_43558,N_43289,N_43270);
or U43559 (N_43559,N_43410,N_43005);
or U43560 (N_43560,N_43395,N_43377);
or U43561 (N_43561,N_43183,N_43339);
nor U43562 (N_43562,N_43327,N_43350);
xor U43563 (N_43563,N_43317,N_43333);
or U43564 (N_43564,N_43409,N_43242);
and U43565 (N_43565,N_43219,N_43233);
or U43566 (N_43566,N_43174,N_43383);
and U43567 (N_43567,N_43320,N_43454);
nand U43568 (N_43568,N_43332,N_43417);
nand U43569 (N_43569,N_43460,N_43046);
and U43570 (N_43570,N_43230,N_43144);
nor U43571 (N_43571,N_43396,N_43181);
and U43572 (N_43572,N_43400,N_43263);
and U43573 (N_43573,N_43121,N_43053);
xor U43574 (N_43574,N_43186,N_43102);
or U43575 (N_43575,N_43462,N_43173);
and U43576 (N_43576,N_43057,N_43406);
xnor U43577 (N_43577,N_43127,N_43148);
nor U43578 (N_43578,N_43124,N_43318);
or U43579 (N_43579,N_43000,N_43037);
or U43580 (N_43580,N_43017,N_43457);
nand U43581 (N_43581,N_43356,N_43106);
and U43582 (N_43582,N_43442,N_43166);
or U43583 (N_43583,N_43193,N_43407);
nor U43584 (N_43584,N_43221,N_43027);
and U43585 (N_43585,N_43363,N_43308);
nor U43586 (N_43586,N_43478,N_43300);
or U43587 (N_43587,N_43170,N_43091);
nand U43588 (N_43588,N_43055,N_43440);
nor U43589 (N_43589,N_43051,N_43255);
and U43590 (N_43590,N_43394,N_43180);
xnor U43591 (N_43591,N_43229,N_43296);
and U43592 (N_43592,N_43262,N_43452);
or U43593 (N_43593,N_43007,N_43038);
nand U43594 (N_43594,N_43331,N_43251);
nand U43595 (N_43595,N_43236,N_43294);
xnor U43596 (N_43596,N_43313,N_43011);
or U43597 (N_43597,N_43120,N_43423);
nand U43598 (N_43598,N_43098,N_43056);
or U43599 (N_43599,N_43129,N_43072);
and U43600 (N_43600,N_43156,N_43366);
nor U43601 (N_43601,N_43244,N_43188);
or U43602 (N_43602,N_43225,N_43465);
xnor U43603 (N_43603,N_43494,N_43379);
xor U43604 (N_43604,N_43103,N_43277);
nand U43605 (N_43605,N_43099,N_43246);
xor U43606 (N_43606,N_43105,N_43136);
or U43607 (N_43607,N_43147,N_43450);
or U43608 (N_43608,N_43260,N_43240);
nand U43609 (N_43609,N_43059,N_43073);
nand U43610 (N_43610,N_43177,N_43375);
or U43611 (N_43611,N_43162,N_43032);
and U43612 (N_43612,N_43304,N_43159);
and U43613 (N_43613,N_43328,N_43272);
nand U43614 (N_43614,N_43309,N_43248);
nor U43615 (N_43615,N_43204,N_43437);
and U43616 (N_43616,N_43171,N_43104);
nand U43617 (N_43617,N_43321,N_43026);
nor U43618 (N_43618,N_43316,N_43145);
nor U43619 (N_43619,N_43430,N_43482);
or U43620 (N_43620,N_43196,N_43201);
or U43621 (N_43621,N_43344,N_43002);
nand U43622 (N_43622,N_43471,N_43458);
nand U43623 (N_43623,N_43372,N_43288);
xor U43624 (N_43624,N_43283,N_43310);
xor U43625 (N_43625,N_43444,N_43432);
and U43626 (N_43626,N_43269,N_43088);
and U43627 (N_43627,N_43401,N_43022);
and U43628 (N_43628,N_43206,N_43371);
xor U43629 (N_43629,N_43388,N_43362);
or U43630 (N_43630,N_43257,N_43092);
and U43631 (N_43631,N_43337,N_43322);
nand U43632 (N_43632,N_43134,N_43498);
and U43633 (N_43633,N_43179,N_43305);
xnor U43634 (N_43634,N_43009,N_43336);
nor U43635 (N_43635,N_43235,N_43013);
nor U43636 (N_43636,N_43312,N_43224);
and U43637 (N_43637,N_43464,N_43266);
or U43638 (N_43638,N_43326,N_43264);
and U43639 (N_43639,N_43131,N_43481);
or U43640 (N_43640,N_43126,N_43157);
nand U43641 (N_43641,N_43324,N_43014);
xnor U43642 (N_43642,N_43267,N_43338);
or U43643 (N_43643,N_43185,N_43469);
and U43644 (N_43644,N_43479,N_43003);
nand U43645 (N_43645,N_43066,N_43043);
nand U43646 (N_43646,N_43380,N_43411);
or U43647 (N_43647,N_43404,N_43382);
and U43648 (N_43648,N_43295,N_43033);
nand U43649 (N_43649,N_43024,N_43335);
and U43650 (N_43650,N_43428,N_43499);
nor U43651 (N_43651,N_43253,N_43397);
or U43652 (N_43652,N_43039,N_43361);
and U43653 (N_43653,N_43029,N_43064);
nand U43654 (N_43654,N_43459,N_43215);
xor U43655 (N_43655,N_43353,N_43128);
or U43656 (N_43656,N_43232,N_43107);
nor U43657 (N_43657,N_43281,N_43047);
or U43658 (N_43658,N_43403,N_43473);
nor U43659 (N_43659,N_43198,N_43485);
and U43660 (N_43660,N_43019,N_43101);
nand U43661 (N_43661,N_43089,N_43285);
or U43662 (N_43662,N_43472,N_43075);
or U43663 (N_43663,N_43455,N_43297);
nand U43664 (N_43664,N_43190,N_43194);
and U43665 (N_43665,N_43378,N_43416);
nand U43666 (N_43666,N_43076,N_43218);
and U43667 (N_43667,N_43167,N_43448);
nor U43668 (N_43668,N_43042,N_43226);
nand U43669 (N_43669,N_43424,N_43274);
or U43670 (N_43670,N_43292,N_43031);
and U43671 (N_43671,N_43386,N_43374);
nand U43672 (N_43672,N_43149,N_43182);
nand U43673 (N_43673,N_43214,N_43419);
nor U43674 (N_43674,N_43393,N_43414);
nand U43675 (N_43675,N_43023,N_43425);
and U43676 (N_43676,N_43209,N_43203);
nor U43677 (N_43677,N_43483,N_43018);
and U43678 (N_43678,N_43329,N_43118);
or U43679 (N_43679,N_43168,N_43030);
or U43680 (N_43680,N_43006,N_43122);
and U43681 (N_43681,N_43197,N_43187);
nand U43682 (N_43682,N_43453,N_43052);
nand U43683 (N_43683,N_43130,N_43373);
or U43684 (N_43684,N_43421,N_43492);
and U43685 (N_43685,N_43477,N_43346);
and U43686 (N_43686,N_43315,N_43094);
and U43687 (N_43687,N_43306,N_43115);
nand U43688 (N_43688,N_43290,N_43265);
nor U43689 (N_43689,N_43110,N_43058);
and U43690 (N_43690,N_43132,N_43298);
nand U43691 (N_43691,N_43340,N_43020);
nor U43692 (N_43692,N_43351,N_43184);
or U43693 (N_43693,N_43474,N_43189);
or U43694 (N_43694,N_43045,N_43389);
nor U43695 (N_43695,N_43176,N_43050);
nor U43696 (N_43696,N_43195,N_43436);
nand U43697 (N_43697,N_43391,N_43341);
nor U43698 (N_43698,N_43268,N_43470);
nor U43699 (N_43699,N_43359,N_43490);
nand U43700 (N_43700,N_43446,N_43139);
and U43701 (N_43701,N_43461,N_43495);
or U43702 (N_43702,N_43001,N_43319);
xnor U43703 (N_43703,N_43314,N_43108);
or U43704 (N_43704,N_43415,N_43412);
nor U43705 (N_43705,N_43142,N_43368);
nor U43706 (N_43706,N_43119,N_43390);
or U43707 (N_43707,N_43241,N_43200);
xnor U43708 (N_43708,N_43068,N_43152);
or U43709 (N_43709,N_43093,N_43258);
xor U43710 (N_43710,N_43302,N_43100);
nor U43711 (N_43711,N_43078,N_43015);
nand U43712 (N_43712,N_43220,N_43497);
nor U43713 (N_43713,N_43199,N_43155);
nor U43714 (N_43714,N_43060,N_43429);
or U43715 (N_43715,N_43280,N_43146);
xnor U43716 (N_43716,N_43114,N_43212);
xor U43717 (N_43717,N_43048,N_43141);
and U43718 (N_43718,N_43165,N_43116);
nor U43719 (N_43719,N_43138,N_43211);
and U43720 (N_43720,N_43311,N_43441);
nor U43721 (N_43721,N_43169,N_43398);
and U43722 (N_43722,N_43422,N_43291);
nand U43723 (N_43723,N_43420,N_43065);
or U43724 (N_43724,N_43081,N_43172);
or U43725 (N_43725,N_43334,N_43080);
nand U43726 (N_43726,N_43256,N_43299);
nand U43727 (N_43727,N_43426,N_43034);
and U43728 (N_43728,N_43447,N_43021);
nor U43729 (N_43729,N_43254,N_43208);
and U43730 (N_43730,N_43250,N_43279);
and U43731 (N_43731,N_43231,N_43247);
nor U43732 (N_43732,N_43301,N_43192);
nand U43733 (N_43733,N_43158,N_43261);
nand U43734 (N_43734,N_43387,N_43480);
nand U43735 (N_43735,N_43463,N_43323);
nand U43736 (N_43736,N_43140,N_43117);
and U43737 (N_43737,N_43496,N_43278);
nand U43738 (N_43738,N_43049,N_43150);
and U43739 (N_43739,N_43237,N_43205);
or U43740 (N_43740,N_43491,N_43125);
nor U43741 (N_43741,N_43035,N_43040);
xnor U43742 (N_43742,N_43227,N_43484);
or U43743 (N_43743,N_43399,N_43111);
or U43744 (N_43744,N_43325,N_43217);
nand U43745 (N_43745,N_43451,N_43367);
nor U43746 (N_43746,N_43154,N_43364);
or U43747 (N_43747,N_43086,N_43273);
xnor U43748 (N_43748,N_43234,N_43486);
or U43749 (N_43749,N_43433,N_43216);
or U43750 (N_43750,N_43484,N_43219);
and U43751 (N_43751,N_43411,N_43463);
xor U43752 (N_43752,N_43148,N_43024);
nor U43753 (N_43753,N_43278,N_43222);
or U43754 (N_43754,N_43327,N_43244);
xnor U43755 (N_43755,N_43304,N_43058);
nor U43756 (N_43756,N_43125,N_43340);
nand U43757 (N_43757,N_43346,N_43003);
and U43758 (N_43758,N_43133,N_43365);
nor U43759 (N_43759,N_43107,N_43065);
nor U43760 (N_43760,N_43027,N_43377);
and U43761 (N_43761,N_43429,N_43008);
nor U43762 (N_43762,N_43108,N_43028);
or U43763 (N_43763,N_43433,N_43395);
and U43764 (N_43764,N_43392,N_43104);
xnor U43765 (N_43765,N_43246,N_43412);
nand U43766 (N_43766,N_43435,N_43350);
nor U43767 (N_43767,N_43495,N_43032);
and U43768 (N_43768,N_43256,N_43468);
nor U43769 (N_43769,N_43190,N_43181);
nand U43770 (N_43770,N_43097,N_43359);
nand U43771 (N_43771,N_43400,N_43151);
nand U43772 (N_43772,N_43372,N_43066);
or U43773 (N_43773,N_43130,N_43274);
nor U43774 (N_43774,N_43199,N_43105);
nor U43775 (N_43775,N_43025,N_43286);
and U43776 (N_43776,N_43098,N_43166);
nand U43777 (N_43777,N_43408,N_43416);
or U43778 (N_43778,N_43003,N_43222);
nand U43779 (N_43779,N_43435,N_43310);
or U43780 (N_43780,N_43170,N_43447);
nand U43781 (N_43781,N_43277,N_43135);
or U43782 (N_43782,N_43043,N_43285);
and U43783 (N_43783,N_43111,N_43482);
and U43784 (N_43784,N_43352,N_43479);
nor U43785 (N_43785,N_43346,N_43259);
nor U43786 (N_43786,N_43379,N_43010);
or U43787 (N_43787,N_43035,N_43317);
or U43788 (N_43788,N_43059,N_43348);
nor U43789 (N_43789,N_43456,N_43238);
nand U43790 (N_43790,N_43068,N_43349);
xor U43791 (N_43791,N_43202,N_43032);
or U43792 (N_43792,N_43063,N_43421);
nand U43793 (N_43793,N_43015,N_43150);
and U43794 (N_43794,N_43003,N_43011);
nor U43795 (N_43795,N_43074,N_43289);
nand U43796 (N_43796,N_43139,N_43175);
or U43797 (N_43797,N_43091,N_43143);
xor U43798 (N_43798,N_43266,N_43475);
or U43799 (N_43799,N_43454,N_43169);
nor U43800 (N_43800,N_43073,N_43423);
and U43801 (N_43801,N_43055,N_43256);
xor U43802 (N_43802,N_43057,N_43169);
and U43803 (N_43803,N_43251,N_43278);
and U43804 (N_43804,N_43028,N_43060);
xor U43805 (N_43805,N_43264,N_43015);
nand U43806 (N_43806,N_43017,N_43233);
nor U43807 (N_43807,N_43342,N_43094);
nor U43808 (N_43808,N_43332,N_43140);
nor U43809 (N_43809,N_43375,N_43248);
nand U43810 (N_43810,N_43175,N_43193);
nand U43811 (N_43811,N_43129,N_43184);
nor U43812 (N_43812,N_43223,N_43173);
nor U43813 (N_43813,N_43016,N_43089);
nand U43814 (N_43814,N_43073,N_43153);
and U43815 (N_43815,N_43169,N_43380);
xnor U43816 (N_43816,N_43132,N_43300);
or U43817 (N_43817,N_43007,N_43152);
xnor U43818 (N_43818,N_43347,N_43150);
and U43819 (N_43819,N_43165,N_43050);
nand U43820 (N_43820,N_43439,N_43096);
and U43821 (N_43821,N_43212,N_43205);
and U43822 (N_43822,N_43325,N_43299);
nor U43823 (N_43823,N_43301,N_43310);
or U43824 (N_43824,N_43183,N_43368);
nor U43825 (N_43825,N_43003,N_43378);
xnor U43826 (N_43826,N_43470,N_43161);
and U43827 (N_43827,N_43221,N_43236);
and U43828 (N_43828,N_43062,N_43471);
nor U43829 (N_43829,N_43062,N_43338);
nand U43830 (N_43830,N_43066,N_43268);
nor U43831 (N_43831,N_43239,N_43128);
and U43832 (N_43832,N_43435,N_43420);
xor U43833 (N_43833,N_43161,N_43101);
or U43834 (N_43834,N_43026,N_43069);
and U43835 (N_43835,N_43403,N_43362);
or U43836 (N_43836,N_43065,N_43475);
or U43837 (N_43837,N_43285,N_43257);
nand U43838 (N_43838,N_43002,N_43024);
and U43839 (N_43839,N_43199,N_43248);
and U43840 (N_43840,N_43426,N_43480);
xnor U43841 (N_43841,N_43167,N_43252);
and U43842 (N_43842,N_43121,N_43339);
nand U43843 (N_43843,N_43118,N_43108);
or U43844 (N_43844,N_43419,N_43436);
nand U43845 (N_43845,N_43140,N_43407);
nor U43846 (N_43846,N_43469,N_43022);
nand U43847 (N_43847,N_43182,N_43000);
nor U43848 (N_43848,N_43338,N_43109);
or U43849 (N_43849,N_43356,N_43043);
or U43850 (N_43850,N_43468,N_43488);
xnor U43851 (N_43851,N_43264,N_43390);
nor U43852 (N_43852,N_43269,N_43160);
nor U43853 (N_43853,N_43032,N_43109);
xor U43854 (N_43854,N_43087,N_43198);
or U43855 (N_43855,N_43062,N_43281);
and U43856 (N_43856,N_43489,N_43377);
xor U43857 (N_43857,N_43084,N_43499);
nand U43858 (N_43858,N_43373,N_43367);
nor U43859 (N_43859,N_43355,N_43022);
nand U43860 (N_43860,N_43362,N_43077);
nor U43861 (N_43861,N_43490,N_43421);
and U43862 (N_43862,N_43281,N_43107);
nand U43863 (N_43863,N_43202,N_43107);
nand U43864 (N_43864,N_43441,N_43010);
or U43865 (N_43865,N_43125,N_43317);
and U43866 (N_43866,N_43437,N_43024);
or U43867 (N_43867,N_43114,N_43008);
nand U43868 (N_43868,N_43281,N_43364);
nor U43869 (N_43869,N_43216,N_43266);
or U43870 (N_43870,N_43278,N_43495);
and U43871 (N_43871,N_43015,N_43401);
nand U43872 (N_43872,N_43402,N_43391);
and U43873 (N_43873,N_43488,N_43370);
nor U43874 (N_43874,N_43036,N_43009);
nand U43875 (N_43875,N_43300,N_43397);
or U43876 (N_43876,N_43302,N_43285);
and U43877 (N_43877,N_43354,N_43054);
nor U43878 (N_43878,N_43030,N_43312);
and U43879 (N_43879,N_43279,N_43383);
and U43880 (N_43880,N_43351,N_43389);
or U43881 (N_43881,N_43459,N_43237);
nor U43882 (N_43882,N_43303,N_43061);
nor U43883 (N_43883,N_43433,N_43183);
or U43884 (N_43884,N_43112,N_43015);
nand U43885 (N_43885,N_43234,N_43223);
xnor U43886 (N_43886,N_43039,N_43394);
and U43887 (N_43887,N_43021,N_43257);
nand U43888 (N_43888,N_43275,N_43133);
xor U43889 (N_43889,N_43244,N_43030);
and U43890 (N_43890,N_43333,N_43015);
xnor U43891 (N_43891,N_43306,N_43411);
or U43892 (N_43892,N_43200,N_43022);
nand U43893 (N_43893,N_43321,N_43312);
and U43894 (N_43894,N_43238,N_43004);
or U43895 (N_43895,N_43435,N_43044);
or U43896 (N_43896,N_43088,N_43128);
nor U43897 (N_43897,N_43398,N_43489);
and U43898 (N_43898,N_43133,N_43447);
or U43899 (N_43899,N_43073,N_43284);
nor U43900 (N_43900,N_43324,N_43355);
nand U43901 (N_43901,N_43148,N_43044);
xor U43902 (N_43902,N_43061,N_43426);
nand U43903 (N_43903,N_43313,N_43124);
and U43904 (N_43904,N_43308,N_43097);
or U43905 (N_43905,N_43253,N_43204);
nor U43906 (N_43906,N_43354,N_43467);
xor U43907 (N_43907,N_43383,N_43257);
nand U43908 (N_43908,N_43136,N_43374);
or U43909 (N_43909,N_43083,N_43377);
nor U43910 (N_43910,N_43096,N_43292);
or U43911 (N_43911,N_43384,N_43161);
xor U43912 (N_43912,N_43013,N_43181);
and U43913 (N_43913,N_43468,N_43303);
nand U43914 (N_43914,N_43391,N_43300);
nor U43915 (N_43915,N_43017,N_43382);
or U43916 (N_43916,N_43016,N_43129);
or U43917 (N_43917,N_43047,N_43417);
nor U43918 (N_43918,N_43101,N_43433);
and U43919 (N_43919,N_43186,N_43205);
nand U43920 (N_43920,N_43169,N_43394);
and U43921 (N_43921,N_43028,N_43310);
nand U43922 (N_43922,N_43076,N_43065);
xor U43923 (N_43923,N_43018,N_43232);
nand U43924 (N_43924,N_43455,N_43462);
nand U43925 (N_43925,N_43293,N_43286);
and U43926 (N_43926,N_43485,N_43478);
or U43927 (N_43927,N_43431,N_43286);
nor U43928 (N_43928,N_43427,N_43101);
or U43929 (N_43929,N_43311,N_43195);
or U43930 (N_43930,N_43476,N_43262);
and U43931 (N_43931,N_43224,N_43333);
nand U43932 (N_43932,N_43323,N_43380);
nor U43933 (N_43933,N_43267,N_43262);
nand U43934 (N_43934,N_43333,N_43098);
nand U43935 (N_43935,N_43402,N_43290);
or U43936 (N_43936,N_43464,N_43257);
xnor U43937 (N_43937,N_43183,N_43301);
nand U43938 (N_43938,N_43033,N_43113);
and U43939 (N_43939,N_43026,N_43320);
nand U43940 (N_43940,N_43232,N_43313);
xor U43941 (N_43941,N_43080,N_43460);
xnor U43942 (N_43942,N_43261,N_43020);
nand U43943 (N_43943,N_43013,N_43077);
xor U43944 (N_43944,N_43436,N_43189);
nand U43945 (N_43945,N_43418,N_43172);
and U43946 (N_43946,N_43178,N_43079);
nand U43947 (N_43947,N_43375,N_43489);
and U43948 (N_43948,N_43292,N_43490);
or U43949 (N_43949,N_43222,N_43247);
or U43950 (N_43950,N_43331,N_43246);
or U43951 (N_43951,N_43054,N_43042);
xnor U43952 (N_43952,N_43472,N_43155);
xnor U43953 (N_43953,N_43258,N_43081);
nand U43954 (N_43954,N_43458,N_43193);
or U43955 (N_43955,N_43359,N_43406);
xor U43956 (N_43956,N_43261,N_43427);
nor U43957 (N_43957,N_43183,N_43054);
xnor U43958 (N_43958,N_43442,N_43497);
xor U43959 (N_43959,N_43375,N_43030);
nand U43960 (N_43960,N_43104,N_43484);
and U43961 (N_43961,N_43194,N_43424);
nand U43962 (N_43962,N_43358,N_43268);
or U43963 (N_43963,N_43207,N_43440);
xnor U43964 (N_43964,N_43200,N_43393);
or U43965 (N_43965,N_43303,N_43138);
and U43966 (N_43966,N_43348,N_43306);
nand U43967 (N_43967,N_43322,N_43499);
or U43968 (N_43968,N_43358,N_43463);
and U43969 (N_43969,N_43205,N_43213);
or U43970 (N_43970,N_43136,N_43333);
and U43971 (N_43971,N_43474,N_43270);
nand U43972 (N_43972,N_43412,N_43251);
nand U43973 (N_43973,N_43216,N_43420);
and U43974 (N_43974,N_43404,N_43223);
and U43975 (N_43975,N_43056,N_43106);
nand U43976 (N_43976,N_43471,N_43181);
or U43977 (N_43977,N_43323,N_43468);
or U43978 (N_43978,N_43224,N_43456);
and U43979 (N_43979,N_43030,N_43445);
nor U43980 (N_43980,N_43300,N_43207);
nor U43981 (N_43981,N_43316,N_43295);
nand U43982 (N_43982,N_43146,N_43019);
or U43983 (N_43983,N_43440,N_43410);
and U43984 (N_43984,N_43471,N_43442);
xor U43985 (N_43985,N_43032,N_43262);
nor U43986 (N_43986,N_43481,N_43051);
and U43987 (N_43987,N_43426,N_43046);
xor U43988 (N_43988,N_43262,N_43330);
or U43989 (N_43989,N_43400,N_43449);
nand U43990 (N_43990,N_43012,N_43120);
or U43991 (N_43991,N_43149,N_43053);
or U43992 (N_43992,N_43386,N_43491);
xnor U43993 (N_43993,N_43069,N_43090);
and U43994 (N_43994,N_43261,N_43304);
or U43995 (N_43995,N_43319,N_43219);
nand U43996 (N_43996,N_43318,N_43265);
nor U43997 (N_43997,N_43434,N_43490);
and U43998 (N_43998,N_43240,N_43329);
or U43999 (N_43999,N_43067,N_43052);
and U44000 (N_44000,N_43779,N_43763);
nor U44001 (N_44001,N_43969,N_43932);
nand U44002 (N_44002,N_43709,N_43597);
nand U44003 (N_44003,N_43582,N_43974);
nand U44004 (N_44004,N_43961,N_43819);
or U44005 (N_44005,N_43717,N_43915);
nand U44006 (N_44006,N_43617,N_43786);
or U44007 (N_44007,N_43569,N_43897);
or U44008 (N_44008,N_43892,N_43669);
nand U44009 (N_44009,N_43814,N_43829);
or U44010 (N_44010,N_43784,N_43524);
nand U44011 (N_44011,N_43735,N_43861);
nand U44012 (N_44012,N_43837,N_43713);
nand U44013 (N_44013,N_43677,N_43531);
nand U44014 (N_44014,N_43654,N_43951);
or U44015 (N_44015,N_43976,N_43873);
nand U44016 (N_44016,N_43935,N_43817);
and U44017 (N_44017,N_43884,N_43648);
xor U44018 (N_44018,N_43908,N_43880);
nor U44019 (N_44019,N_43722,N_43872);
or U44020 (N_44020,N_43902,N_43664);
and U44021 (N_44021,N_43962,N_43813);
nand U44022 (N_44022,N_43668,N_43665);
or U44023 (N_44023,N_43930,N_43611);
or U44024 (N_44024,N_43538,N_43893);
or U44025 (N_44025,N_43938,N_43724);
nor U44026 (N_44026,N_43841,N_43711);
and U44027 (N_44027,N_43656,N_43737);
or U44028 (N_44028,N_43614,N_43972);
and U44029 (N_44029,N_43719,N_43681);
and U44030 (N_44030,N_43781,N_43583);
nand U44031 (N_44031,N_43996,N_43761);
nor U44032 (N_44032,N_43522,N_43682);
or U44033 (N_44033,N_43562,N_43639);
nand U44034 (N_44034,N_43580,N_43793);
nor U44035 (N_44035,N_43822,N_43621);
xnor U44036 (N_44036,N_43785,N_43868);
xor U44037 (N_44037,N_43846,N_43758);
or U44038 (N_44038,N_43762,N_43710);
nand U44039 (N_44039,N_43997,N_43848);
nor U44040 (N_44040,N_43864,N_43802);
nand U44041 (N_44041,N_43800,N_43771);
or U44042 (N_44042,N_43678,N_43593);
nor U44043 (N_44043,N_43657,N_43693);
nor U44044 (N_44044,N_43586,N_43827);
or U44045 (N_44045,N_43756,N_43749);
or U44046 (N_44046,N_43699,N_43752);
xnor U44047 (N_44047,N_43843,N_43518);
or U44048 (N_44048,N_43670,N_43831);
nand U44049 (N_44049,N_43615,N_43564);
nand U44050 (N_44050,N_43501,N_43940);
or U44051 (N_44051,N_43759,N_43547);
nand U44052 (N_44052,N_43772,N_43943);
and U44053 (N_44053,N_43592,N_43673);
nand U44054 (N_44054,N_43859,N_43515);
nor U44055 (N_44055,N_43568,N_43557);
or U44056 (N_44056,N_43643,N_43730);
and U44057 (N_44057,N_43548,N_43584);
and U44058 (N_44058,N_43971,N_43700);
nand U44059 (N_44059,N_43856,N_43550);
xor U44060 (N_44060,N_43746,N_43581);
and U44061 (N_44061,N_43714,N_43929);
nor U44062 (N_44062,N_43979,N_43513);
nand U44063 (N_44063,N_43606,N_43750);
nor U44064 (N_44064,N_43543,N_43958);
and U44065 (N_44065,N_43502,N_43875);
xnor U44066 (N_44066,N_43900,N_43903);
or U44067 (N_44067,N_43888,N_43671);
and U44068 (N_44068,N_43980,N_43815);
nand U44069 (N_44069,N_43808,N_43939);
xnor U44070 (N_44070,N_43733,N_43532);
nor U44071 (N_44071,N_43994,N_43944);
nand U44072 (N_44072,N_43936,N_43744);
or U44073 (N_44073,N_43645,N_43517);
or U44074 (N_44074,N_43541,N_43504);
and U44075 (N_44075,N_43916,N_43701);
nor U44076 (N_44076,N_43540,N_43549);
or U44077 (N_44077,N_43818,N_43858);
or U44078 (N_44078,N_43596,N_43866);
nand U44079 (N_44079,N_43616,N_43847);
nor U44080 (N_44080,N_43716,N_43707);
nand U44081 (N_44081,N_43839,N_43807);
and U44082 (N_44082,N_43732,N_43528);
or U44083 (N_44083,N_43613,N_43925);
nor U44084 (N_44084,N_43955,N_43926);
nor U44085 (N_44085,N_43765,N_43742);
or U44086 (N_44086,N_43680,N_43816);
or U44087 (N_44087,N_43510,N_43555);
xor U44088 (N_44088,N_43505,N_43977);
and U44089 (N_44089,N_43529,N_43834);
nand U44090 (N_44090,N_43798,N_43795);
and U44091 (N_44091,N_43948,N_43525);
nor U44092 (N_44092,N_43629,N_43849);
or U44093 (N_44093,N_43684,N_43715);
and U44094 (N_44094,N_43566,N_43556);
or U44095 (N_44095,N_43734,N_43533);
or U44096 (N_44096,N_43877,N_43745);
and U44097 (N_44097,N_43953,N_43706);
nand U44098 (N_44098,N_43791,N_43917);
nor U44099 (N_44099,N_43904,N_43991);
and U44100 (N_44100,N_43981,N_43812);
nand U44101 (N_44101,N_43530,N_43627);
and U44102 (N_44102,N_43828,N_43600);
xor U44103 (N_44103,N_43565,N_43898);
nand U44104 (N_44104,N_43728,N_43782);
and U44105 (N_44105,N_43747,N_43512);
or U44106 (N_44106,N_43748,N_43883);
nor U44107 (N_44107,N_43650,N_43686);
nand U44108 (N_44108,N_43865,N_43623);
xor U44109 (N_44109,N_43907,N_43960);
or U44110 (N_44110,N_43850,N_43878);
or U44111 (N_44111,N_43952,N_43690);
and U44112 (N_44112,N_43889,N_43712);
and U44113 (N_44113,N_43990,N_43726);
nand U44114 (N_44114,N_43914,N_43601);
and U44115 (N_44115,N_43937,N_43637);
nand U44116 (N_44116,N_43918,N_43704);
and U44117 (N_44117,N_43574,N_43723);
nand U44118 (N_44118,N_43797,N_43545);
and U44119 (N_44119,N_43635,N_43634);
or U44120 (N_44120,N_43824,N_43519);
nand U44121 (N_44121,N_43661,N_43941);
nor U44122 (N_44122,N_43741,N_43571);
or U44123 (N_44123,N_43942,N_43927);
nor U44124 (N_44124,N_43626,N_43516);
and U44125 (N_44125,N_43973,N_43867);
nand U44126 (N_44126,N_43810,N_43691);
nand U44127 (N_44127,N_43823,N_43546);
and U44128 (N_44128,N_43780,N_43755);
or U44129 (N_44129,N_43983,N_43886);
or U44130 (N_44130,N_43905,N_43685);
or U44131 (N_44131,N_43820,N_43636);
and U44132 (N_44132,N_43933,N_43663);
nand U44133 (N_44133,N_43885,N_43804);
and U44134 (N_44134,N_43508,N_43870);
and U44135 (N_44135,N_43854,N_43551);
or U44136 (N_44136,N_43595,N_43975);
xor U44137 (N_44137,N_43922,N_43598);
or U44138 (N_44138,N_43862,N_43766);
nand U44139 (N_44139,N_43590,N_43777);
nand U44140 (N_44140,N_43662,N_43570);
xor U44141 (N_44141,N_43934,N_43567);
xor U44142 (N_44142,N_43931,N_43835);
or U44143 (N_44143,N_43845,N_43842);
nand U44144 (N_44144,N_43840,N_43695);
or U44145 (N_44145,N_43891,N_43985);
nor U44146 (N_44146,N_43901,N_43751);
nor U44147 (N_44147,N_43638,N_43949);
xnor U44148 (N_44148,N_43694,N_43632);
nand U44149 (N_44149,N_43855,N_43954);
xor U44150 (N_44150,N_43527,N_43988);
nand U44151 (N_44151,N_43956,N_43725);
nand U44152 (N_44152,N_43757,N_43882);
nand U44153 (N_44153,N_43760,N_43575);
nor U44154 (N_44154,N_43640,N_43633);
or U44155 (N_44155,N_43853,N_43628);
or U44156 (N_44156,N_43890,N_43544);
nor U44157 (N_44157,N_43676,N_43964);
nor U44158 (N_44158,N_43836,N_43776);
or U44159 (N_44159,N_43579,N_43563);
or U44160 (N_44160,N_43651,N_43683);
nand U44161 (N_44161,N_43622,N_43561);
and U44162 (N_44162,N_43687,N_43619);
and U44163 (N_44163,N_43799,N_43718);
xor U44164 (N_44164,N_43618,N_43796);
nor U44165 (N_44165,N_43803,N_43863);
and U44166 (N_44166,N_43604,N_43659);
xnor U44167 (N_44167,N_43801,N_43610);
or U44168 (N_44168,N_43652,N_43558);
or U44169 (N_44169,N_43790,N_43999);
nor U44170 (N_44170,N_43692,N_43526);
nor U44171 (N_44171,N_43774,N_43511);
and U44172 (N_44172,N_43647,N_43646);
nand U44173 (N_44173,N_43989,N_43675);
and U44174 (N_44174,N_43993,N_43894);
and U44175 (N_44175,N_43642,N_43767);
and U44176 (N_44176,N_43624,N_43631);
or U44177 (N_44177,N_43572,N_43920);
or U44178 (N_44178,N_43871,N_43775);
nor U44179 (N_44179,N_43738,N_43832);
nor U44180 (N_44180,N_43950,N_43912);
xnor U44181 (N_44181,N_43923,N_43919);
or U44182 (N_44182,N_43874,N_43553);
nand U44183 (N_44183,N_43599,N_43587);
xor U44184 (N_44184,N_43753,N_43844);
nand U44185 (N_44185,N_43708,N_43591);
and U44186 (N_44186,N_43968,N_43559);
or U44187 (N_44187,N_43739,N_43852);
nor U44188 (N_44188,N_43794,N_43913);
nand U44189 (N_44189,N_43788,N_43509);
nand U44190 (N_44190,N_43560,N_43523);
xor U44191 (N_44191,N_43731,N_43928);
or U44192 (N_44192,N_43982,N_43674);
or U44193 (N_44193,N_43653,N_43605);
and U44194 (N_44194,N_43768,N_43965);
and U44195 (N_44195,N_43698,N_43946);
nand U44196 (N_44196,N_43536,N_43537);
and U44197 (N_44197,N_43881,N_43506);
or U44198 (N_44198,N_43589,N_43860);
or U44199 (N_44199,N_43658,N_43585);
and U44200 (N_44200,N_43770,N_43998);
nand U44201 (N_44201,N_43821,N_43500);
and U44202 (N_44202,N_43727,N_43966);
nand U44203 (N_44203,N_43655,N_43970);
nand U44204 (N_44204,N_43641,N_43825);
nor U44205 (N_44205,N_43666,N_43667);
and U44206 (N_44206,N_43729,N_43895);
nand U44207 (N_44207,N_43534,N_43987);
and U44208 (N_44208,N_43539,N_43764);
or U44209 (N_44209,N_43924,N_43521);
and U44210 (N_44210,N_43743,N_43705);
and U44211 (N_44211,N_43688,N_43789);
and U44212 (N_44212,N_43672,N_43826);
nor U44213 (N_44213,N_43702,N_43769);
and U44214 (N_44214,N_43887,N_43910);
and U44215 (N_44215,N_43554,N_43503);
xnor U44216 (N_44216,N_43911,N_43876);
nor U44217 (N_44217,N_43754,N_43602);
nor U44218 (N_44218,N_43806,N_43805);
nand U44219 (N_44219,N_43899,N_43620);
or U44220 (N_44220,N_43857,N_43736);
xnor U44221 (N_44221,N_43535,N_43609);
and U44222 (N_44222,N_43607,N_43573);
nor U44223 (N_44223,N_43740,N_43959);
and U44224 (N_44224,N_43689,N_43957);
nor U44225 (N_44225,N_43612,N_43514);
or U44226 (N_44226,N_43588,N_43869);
or U44227 (N_44227,N_43603,N_43967);
and U44228 (N_44228,N_43906,N_43995);
nand U44229 (N_44229,N_43721,N_43696);
nand U44230 (N_44230,N_43703,N_43552);
and U44231 (N_44231,N_43625,N_43644);
or U44232 (N_44232,N_43921,N_43578);
and U44233 (N_44233,N_43792,N_43720);
and U44234 (N_44234,N_43778,N_43909);
nand U44235 (N_44235,N_43660,N_43992);
and U44236 (N_44236,N_43833,N_43838);
or U44237 (N_44237,N_43945,N_43947);
or U44238 (N_44238,N_43576,N_43879);
xor U44239 (N_44239,N_43608,N_43630);
or U44240 (N_44240,N_43679,N_43809);
nor U44241 (N_44241,N_43787,N_43811);
nor U44242 (N_44242,N_43963,N_43594);
nand U44243 (N_44243,N_43697,N_43649);
or U44244 (N_44244,N_43978,N_43542);
and U44245 (N_44245,N_43577,N_43896);
nand U44246 (N_44246,N_43520,N_43830);
or U44247 (N_44247,N_43851,N_43773);
nor U44248 (N_44248,N_43986,N_43507);
nor U44249 (N_44249,N_43984,N_43783);
or U44250 (N_44250,N_43604,N_43741);
nand U44251 (N_44251,N_43530,N_43712);
xor U44252 (N_44252,N_43522,N_43516);
and U44253 (N_44253,N_43911,N_43572);
nand U44254 (N_44254,N_43828,N_43919);
xnor U44255 (N_44255,N_43991,N_43925);
nor U44256 (N_44256,N_43984,N_43988);
and U44257 (N_44257,N_43959,N_43504);
or U44258 (N_44258,N_43602,N_43847);
nor U44259 (N_44259,N_43716,N_43809);
nor U44260 (N_44260,N_43652,N_43790);
xnor U44261 (N_44261,N_43831,N_43882);
nand U44262 (N_44262,N_43866,N_43658);
nor U44263 (N_44263,N_43876,N_43835);
nand U44264 (N_44264,N_43999,N_43750);
nand U44265 (N_44265,N_43819,N_43603);
or U44266 (N_44266,N_43742,N_43697);
nor U44267 (N_44267,N_43850,N_43531);
or U44268 (N_44268,N_43688,N_43677);
nand U44269 (N_44269,N_43839,N_43627);
or U44270 (N_44270,N_43642,N_43866);
and U44271 (N_44271,N_43827,N_43674);
nand U44272 (N_44272,N_43849,N_43848);
xnor U44273 (N_44273,N_43561,N_43775);
nand U44274 (N_44274,N_43585,N_43604);
or U44275 (N_44275,N_43858,N_43944);
and U44276 (N_44276,N_43579,N_43526);
nand U44277 (N_44277,N_43750,N_43715);
xor U44278 (N_44278,N_43817,N_43877);
or U44279 (N_44279,N_43564,N_43757);
xor U44280 (N_44280,N_43569,N_43666);
or U44281 (N_44281,N_43703,N_43715);
or U44282 (N_44282,N_43811,N_43927);
nand U44283 (N_44283,N_43714,N_43516);
and U44284 (N_44284,N_43676,N_43783);
or U44285 (N_44285,N_43689,N_43708);
nand U44286 (N_44286,N_43736,N_43830);
nor U44287 (N_44287,N_43641,N_43716);
nor U44288 (N_44288,N_43961,N_43987);
nor U44289 (N_44289,N_43524,N_43732);
or U44290 (N_44290,N_43504,N_43774);
nor U44291 (N_44291,N_43939,N_43833);
and U44292 (N_44292,N_43955,N_43947);
and U44293 (N_44293,N_43545,N_43984);
nor U44294 (N_44294,N_43637,N_43758);
or U44295 (N_44295,N_43793,N_43845);
or U44296 (N_44296,N_43704,N_43643);
nor U44297 (N_44297,N_43659,N_43579);
or U44298 (N_44298,N_43690,N_43936);
xnor U44299 (N_44299,N_43501,N_43583);
nor U44300 (N_44300,N_43874,N_43981);
nand U44301 (N_44301,N_43888,N_43732);
xnor U44302 (N_44302,N_43541,N_43903);
or U44303 (N_44303,N_43806,N_43634);
nor U44304 (N_44304,N_43541,N_43615);
nor U44305 (N_44305,N_43988,N_43827);
and U44306 (N_44306,N_43615,N_43585);
or U44307 (N_44307,N_43687,N_43801);
or U44308 (N_44308,N_43556,N_43637);
or U44309 (N_44309,N_43736,N_43718);
xnor U44310 (N_44310,N_43954,N_43666);
and U44311 (N_44311,N_43579,N_43999);
nor U44312 (N_44312,N_43978,N_43850);
xnor U44313 (N_44313,N_43871,N_43725);
and U44314 (N_44314,N_43839,N_43706);
and U44315 (N_44315,N_43876,N_43542);
xnor U44316 (N_44316,N_43595,N_43925);
and U44317 (N_44317,N_43708,N_43756);
nor U44318 (N_44318,N_43587,N_43755);
nand U44319 (N_44319,N_43743,N_43735);
and U44320 (N_44320,N_43763,N_43703);
nor U44321 (N_44321,N_43657,N_43625);
nand U44322 (N_44322,N_43522,N_43872);
or U44323 (N_44323,N_43876,N_43526);
nand U44324 (N_44324,N_43549,N_43638);
xor U44325 (N_44325,N_43551,N_43527);
nor U44326 (N_44326,N_43990,N_43782);
or U44327 (N_44327,N_43551,N_43619);
and U44328 (N_44328,N_43982,N_43912);
nand U44329 (N_44329,N_43896,N_43943);
nand U44330 (N_44330,N_43939,N_43651);
and U44331 (N_44331,N_43834,N_43601);
nand U44332 (N_44332,N_43762,N_43769);
or U44333 (N_44333,N_43526,N_43686);
nor U44334 (N_44334,N_43678,N_43557);
nand U44335 (N_44335,N_43778,N_43818);
or U44336 (N_44336,N_43675,N_43554);
or U44337 (N_44337,N_43706,N_43680);
nor U44338 (N_44338,N_43607,N_43722);
nand U44339 (N_44339,N_43991,N_43659);
or U44340 (N_44340,N_43766,N_43979);
nand U44341 (N_44341,N_43865,N_43921);
xnor U44342 (N_44342,N_43610,N_43716);
nand U44343 (N_44343,N_43678,N_43568);
nand U44344 (N_44344,N_43560,N_43647);
or U44345 (N_44345,N_43785,N_43900);
or U44346 (N_44346,N_43600,N_43733);
and U44347 (N_44347,N_43577,N_43728);
or U44348 (N_44348,N_43544,N_43763);
and U44349 (N_44349,N_43539,N_43585);
and U44350 (N_44350,N_43800,N_43630);
and U44351 (N_44351,N_43762,N_43897);
nor U44352 (N_44352,N_43582,N_43701);
nor U44353 (N_44353,N_43997,N_43882);
or U44354 (N_44354,N_43789,N_43572);
nand U44355 (N_44355,N_43846,N_43502);
nor U44356 (N_44356,N_43719,N_43710);
nand U44357 (N_44357,N_43983,N_43621);
nand U44358 (N_44358,N_43748,N_43539);
or U44359 (N_44359,N_43838,N_43733);
nand U44360 (N_44360,N_43916,N_43666);
and U44361 (N_44361,N_43821,N_43967);
nor U44362 (N_44362,N_43588,N_43823);
nand U44363 (N_44363,N_43515,N_43843);
nor U44364 (N_44364,N_43628,N_43778);
and U44365 (N_44365,N_43963,N_43758);
nor U44366 (N_44366,N_43806,N_43742);
or U44367 (N_44367,N_43827,N_43629);
and U44368 (N_44368,N_43933,N_43718);
xor U44369 (N_44369,N_43582,N_43699);
nor U44370 (N_44370,N_43729,N_43633);
nor U44371 (N_44371,N_43785,N_43621);
nand U44372 (N_44372,N_43657,N_43530);
nor U44373 (N_44373,N_43813,N_43817);
and U44374 (N_44374,N_43940,N_43916);
nor U44375 (N_44375,N_43909,N_43930);
nor U44376 (N_44376,N_43885,N_43584);
nor U44377 (N_44377,N_43805,N_43515);
nand U44378 (N_44378,N_43697,N_43637);
nor U44379 (N_44379,N_43883,N_43911);
or U44380 (N_44380,N_43535,N_43661);
xor U44381 (N_44381,N_43889,N_43552);
nand U44382 (N_44382,N_43674,N_43797);
nor U44383 (N_44383,N_43772,N_43576);
xnor U44384 (N_44384,N_43599,N_43826);
nor U44385 (N_44385,N_43724,N_43895);
nand U44386 (N_44386,N_43537,N_43830);
or U44387 (N_44387,N_43675,N_43652);
or U44388 (N_44388,N_43667,N_43590);
and U44389 (N_44389,N_43923,N_43834);
nand U44390 (N_44390,N_43703,N_43923);
nand U44391 (N_44391,N_43696,N_43671);
nor U44392 (N_44392,N_43665,N_43893);
and U44393 (N_44393,N_43841,N_43800);
nor U44394 (N_44394,N_43951,N_43969);
nor U44395 (N_44395,N_43610,N_43762);
nand U44396 (N_44396,N_43556,N_43616);
nor U44397 (N_44397,N_43792,N_43863);
and U44398 (N_44398,N_43857,N_43902);
nor U44399 (N_44399,N_43610,N_43731);
nand U44400 (N_44400,N_43789,N_43584);
and U44401 (N_44401,N_43833,N_43613);
nand U44402 (N_44402,N_43500,N_43815);
and U44403 (N_44403,N_43712,N_43645);
nor U44404 (N_44404,N_43825,N_43672);
and U44405 (N_44405,N_43637,N_43806);
nor U44406 (N_44406,N_43932,N_43885);
nor U44407 (N_44407,N_43844,N_43911);
and U44408 (N_44408,N_43562,N_43668);
nor U44409 (N_44409,N_43939,N_43759);
xnor U44410 (N_44410,N_43729,N_43717);
or U44411 (N_44411,N_43896,N_43569);
xor U44412 (N_44412,N_43659,N_43795);
and U44413 (N_44413,N_43609,N_43695);
and U44414 (N_44414,N_43881,N_43610);
nor U44415 (N_44415,N_43977,N_43563);
nand U44416 (N_44416,N_43520,N_43816);
nand U44417 (N_44417,N_43652,N_43576);
or U44418 (N_44418,N_43937,N_43993);
nand U44419 (N_44419,N_43708,N_43776);
nor U44420 (N_44420,N_43714,N_43579);
nor U44421 (N_44421,N_43505,N_43764);
nor U44422 (N_44422,N_43962,N_43632);
or U44423 (N_44423,N_43976,N_43574);
nand U44424 (N_44424,N_43974,N_43954);
or U44425 (N_44425,N_43658,N_43841);
or U44426 (N_44426,N_43858,N_43779);
nand U44427 (N_44427,N_43561,N_43828);
and U44428 (N_44428,N_43928,N_43531);
and U44429 (N_44429,N_43691,N_43503);
nand U44430 (N_44430,N_43848,N_43940);
and U44431 (N_44431,N_43785,N_43897);
nor U44432 (N_44432,N_43780,N_43846);
and U44433 (N_44433,N_43518,N_43539);
and U44434 (N_44434,N_43841,N_43805);
nor U44435 (N_44435,N_43744,N_43963);
and U44436 (N_44436,N_43921,N_43738);
nor U44437 (N_44437,N_43767,N_43910);
and U44438 (N_44438,N_43669,N_43567);
and U44439 (N_44439,N_43626,N_43944);
and U44440 (N_44440,N_43774,N_43627);
and U44441 (N_44441,N_43534,N_43749);
and U44442 (N_44442,N_43528,N_43526);
and U44443 (N_44443,N_43785,N_43977);
nand U44444 (N_44444,N_43876,N_43600);
nor U44445 (N_44445,N_43753,N_43597);
nand U44446 (N_44446,N_43987,N_43624);
nor U44447 (N_44447,N_43857,N_43567);
and U44448 (N_44448,N_43600,N_43902);
nor U44449 (N_44449,N_43785,N_43641);
and U44450 (N_44450,N_43978,N_43710);
and U44451 (N_44451,N_43851,N_43799);
xor U44452 (N_44452,N_43582,N_43857);
nor U44453 (N_44453,N_43504,N_43882);
nor U44454 (N_44454,N_43974,N_43695);
or U44455 (N_44455,N_43979,N_43907);
or U44456 (N_44456,N_43553,N_43664);
or U44457 (N_44457,N_43802,N_43868);
and U44458 (N_44458,N_43711,N_43906);
xnor U44459 (N_44459,N_43749,N_43791);
or U44460 (N_44460,N_43888,N_43664);
and U44461 (N_44461,N_43756,N_43640);
nor U44462 (N_44462,N_43901,N_43911);
nand U44463 (N_44463,N_43987,N_43890);
or U44464 (N_44464,N_43578,N_43635);
xor U44465 (N_44465,N_43563,N_43957);
nor U44466 (N_44466,N_43941,N_43513);
nand U44467 (N_44467,N_43667,N_43616);
nor U44468 (N_44468,N_43872,N_43699);
nand U44469 (N_44469,N_43624,N_43534);
nor U44470 (N_44470,N_43673,N_43501);
or U44471 (N_44471,N_43747,N_43640);
nor U44472 (N_44472,N_43586,N_43669);
nand U44473 (N_44473,N_43721,N_43722);
and U44474 (N_44474,N_43995,N_43991);
nor U44475 (N_44475,N_43875,N_43710);
and U44476 (N_44476,N_43912,N_43673);
nand U44477 (N_44477,N_43694,N_43838);
and U44478 (N_44478,N_43971,N_43503);
nor U44479 (N_44479,N_43955,N_43950);
or U44480 (N_44480,N_43637,N_43734);
nor U44481 (N_44481,N_43547,N_43748);
and U44482 (N_44482,N_43986,N_43829);
xnor U44483 (N_44483,N_43777,N_43942);
or U44484 (N_44484,N_43519,N_43916);
nand U44485 (N_44485,N_43539,N_43707);
or U44486 (N_44486,N_43692,N_43771);
and U44487 (N_44487,N_43622,N_43858);
and U44488 (N_44488,N_43551,N_43931);
nor U44489 (N_44489,N_43837,N_43864);
or U44490 (N_44490,N_43737,N_43741);
or U44491 (N_44491,N_43591,N_43842);
and U44492 (N_44492,N_43570,N_43914);
nor U44493 (N_44493,N_43837,N_43598);
nor U44494 (N_44494,N_43971,N_43984);
and U44495 (N_44495,N_43784,N_43791);
and U44496 (N_44496,N_43862,N_43784);
and U44497 (N_44497,N_43773,N_43809);
or U44498 (N_44498,N_43890,N_43741);
and U44499 (N_44499,N_43608,N_43500);
nor U44500 (N_44500,N_44091,N_44087);
or U44501 (N_44501,N_44419,N_44041);
nor U44502 (N_44502,N_44317,N_44133);
or U44503 (N_44503,N_44430,N_44411);
nand U44504 (N_44504,N_44273,N_44453);
nor U44505 (N_44505,N_44201,N_44367);
nand U44506 (N_44506,N_44197,N_44018);
nand U44507 (N_44507,N_44167,N_44145);
and U44508 (N_44508,N_44435,N_44375);
or U44509 (N_44509,N_44443,N_44467);
nand U44510 (N_44510,N_44229,N_44011);
or U44511 (N_44511,N_44462,N_44265);
and U44512 (N_44512,N_44387,N_44454);
and U44513 (N_44513,N_44100,N_44422);
or U44514 (N_44514,N_44272,N_44108);
and U44515 (N_44515,N_44464,N_44267);
or U44516 (N_44516,N_44020,N_44045);
or U44517 (N_44517,N_44287,N_44303);
and U44518 (N_44518,N_44295,N_44327);
and U44519 (N_44519,N_44063,N_44074);
xor U44520 (N_44520,N_44230,N_44030);
and U44521 (N_44521,N_44460,N_44234);
and U44522 (N_44522,N_44456,N_44362);
or U44523 (N_44523,N_44266,N_44024);
nor U44524 (N_44524,N_44298,N_44181);
and U44525 (N_44525,N_44421,N_44363);
and U44526 (N_44526,N_44347,N_44242);
nor U44527 (N_44527,N_44006,N_44243);
nor U44528 (N_44528,N_44216,N_44334);
nor U44529 (N_44529,N_44007,N_44301);
nand U44530 (N_44530,N_44379,N_44206);
or U44531 (N_44531,N_44010,N_44195);
nor U44532 (N_44532,N_44068,N_44495);
nor U44533 (N_44533,N_44226,N_44213);
xnor U44534 (N_44534,N_44142,N_44324);
xnor U44535 (N_44535,N_44268,N_44326);
nand U44536 (N_44536,N_44117,N_44075);
nand U44537 (N_44537,N_44439,N_44027);
or U44538 (N_44538,N_44366,N_44188);
xnor U44539 (N_44539,N_44028,N_44121);
or U44540 (N_44540,N_44158,N_44440);
nor U44541 (N_44541,N_44249,N_44048);
and U44542 (N_44542,N_44246,N_44178);
and U44543 (N_44543,N_44135,N_44157);
and U44544 (N_44544,N_44052,N_44138);
nor U44545 (N_44545,N_44002,N_44388);
nand U44546 (N_44546,N_44207,N_44349);
nand U44547 (N_44547,N_44497,N_44047);
nand U44548 (N_44548,N_44170,N_44403);
xor U44549 (N_44549,N_44104,N_44253);
or U44550 (N_44550,N_44164,N_44290);
nor U44551 (N_44551,N_44037,N_44374);
or U44552 (N_44552,N_44154,N_44448);
nand U44553 (N_44553,N_44054,N_44012);
and U44554 (N_44554,N_44199,N_44129);
nor U44555 (N_44555,N_44274,N_44044);
xor U44556 (N_44556,N_44381,N_44466);
and U44557 (N_44557,N_44481,N_44355);
and U44558 (N_44558,N_44364,N_44162);
or U44559 (N_44559,N_44437,N_44203);
nor U44560 (N_44560,N_44306,N_44310);
nor U44561 (N_44561,N_44369,N_44077);
nor U44562 (N_44562,N_44472,N_44341);
or U44563 (N_44563,N_44286,N_44130);
nand U44564 (N_44564,N_44370,N_44008);
xor U44565 (N_44565,N_44088,N_44136);
nand U44566 (N_44566,N_44254,N_44407);
or U44567 (N_44567,N_44311,N_44026);
and U44568 (N_44568,N_44275,N_44185);
and U44569 (N_44569,N_44262,N_44353);
and U44570 (N_44570,N_44478,N_44227);
or U44571 (N_44571,N_44291,N_44480);
xnor U44572 (N_44572,N_44457,N_44050);
nor U44573 (N_44573,N_44248,N_44487);
xnor U44574 (N_44574,N_44269,N_44016);
and U44575 (N_44575,N_44445,N_44289);
nor U44576 (N_44576,N_44413,N_44415);
nand U44577 (N_44577,N_44376,N_44163);
xor U44578 (N_44578,N_44186,N_44198);
nand U44579 (N_44579,N_44228,N_44049);
nor U44580 (N_44580,N_44486,N_44384);
nor U44581 (N_44581,N_44490,N_44083);
nand U44582 (N_44582,N_44488,N_44156);
nand U44583 (N_44583,N_44149,N_44132);
xnor U44584 (N_44584,N_44114,N_44019);
nor U44585 (N_44585,N_44172,N_44250);
nor U44586 (N_44586,N_44238,N_44039);
and U44587 (N_44587,N_44465,N_44321);
nor U44588 (N_44588,N_44471,N_44082);
or U44589 (N_44589,N_44496,N_44498);
and U44590 (N_44590,N_44451,N_44420);
or U44591 (N_44591,N_44015,N_44125);
or U44592 (N_44592,N_44424,N_44463);
nor U44593 (N_44593,N_44279,N_44067);
and U44594 (N_44594,N_44360,N_44492);
xnor U44595 (N_44595,N_44414,N_44078);
and U44596 (N_44596,N_44174,N_44278);
xnor U44597 (N_44597,N_44493,N_44211);
xor U44598 (N_44598,N_44080,N_44389);
nand U44599 (N_44599,N_44373,N_44051);
and U44600 (N_44600,N_44475,N_44412);
or U44601 (N_44601,N_44208,N_44281);
or U44602 (N_44602,N_44426,N_44469);
or U44603 (N_44603,N_44260,N_44022);
or U44604 (N_44604,N_44473,N_44089);
or U44605 (N_44605,N_44292,N_44425);
and U44606 (N_44606,N_44474,N_44252);
nor U44607 (N_44607,N_44461,N_44072);
or U44608 (N_44608,N_44377,N_44476);
and U44609 (N_44609,N_44432,N_44401);
or U44610 (N_44610,N_44479,N_44318);
or U44611 (N_44611,N_44155,N_44299);
and U44612 (N_44612,N_44499,N_44331);
nand U44613 (N_44613,N_44235,N_44031);
nand U44614 (N_44614,N_44337,N_44442);
nand U44615 (N_44615,N_44222,N_44485);
nand U44616 (N_44616,N_44323,N_44137);
nor U44617 (N_44617,N_44231,N_44131);
nand U44618 (N_44618,N_44320,N_44069);
nand U44619 (N_44619,N_44300,N_44212);
or U44620 (N_44620,N_44126,N_44236);
nor U44621 (N_44621,N_44062,N_44304);
nor U44622 (N_44622,N_44245,N_44093);
xnor U44623 (N_44623,N_44055,N_44101);
nor U44624 (N_44624,N_44122,N_44297);
or U44625 (N_44625,N_44204,N_44393);
nor U44626 (N_44626,N_44345,N_44284);
or U44627 (N_44627,N_44309,N_44491);
or U44628 (N_44628,N_44086,N_44308);
and U44629 (N_44629,N_44033,N_44150);
nor U44630 (N_44630,N_44214,N_44111);
nand U44631 (N_44631,N_44009,N_44194);
xor U44632 (N_44632,N_44280,N_44329);
and U44633 (N_44633,N_44179,N_44336);
nand U44634 (N_44634,N_44431,N_44094);
nand U44635 (N_44635,N_44351,N_44056);
xnor U44636 (N_44636,N_44438,N_44118);
or U44637 (N_44637,N_44277,N_44271);
nand U44638 (N_44638,N_44139,N_44200);
nand U44639 (N_44639,N_44017,N_44128);
or U44640 (N_44640,N_44064,N_44410);
nor U44641 (N_44641,N_44209,N_44219);
nand U44642 (N_44642,N_44202,N_44107);
or U44643 (N_44643,N_44258,N_44313);
nor U44644 (N_44644,N_44294,N_44482);
or U44645 (N_44645,N_44160,N_44116);
xnor U44646 (N_44646,N_44084,N_44428);
xnor U44647 (N_44647,N_44434,N_44057);
xnor U44648 (N_44648,N_44354,N_44058);
nor U44649 (N_44649,N_44314,N_44021);
nand U44650 (N_44650,N_44400,N_44240);
xnor U44651 (N_44651,N_44073,N_44099);
or U44652 (N_44652,N_44232,N_44061);
nor U44653 (N_44653,N_44494,N_44447);
nand U44654 (N_44654,N_44293,N_44436);
and U44655 (N_44655,N_44257,N_44040);
or U44656 (N_44656,N_44095,N_44004);
and U44657 (N_44657,N_44459,N_44283);
or U44658 (N_44658,N_44408,N_44023);
nor U44659 (N_44659,N_44070,N_44035);
and U44660 (N_44660,N_44391,N_44405);
xnor U44661 (N_44661,N_44120,N_44263);
nor U44662 (N_44662,N_44344,N_44429);
and U44663 (N_44663,N_44416,N_44098);
and U44664 (N_44664,N_44350,N_44398);
and U44665 (N_44665,N_44319,N_44127);
nor U44666 (N_44666,N_44109,N_44143);
and U44667 (N_44667,N_44288,N_44441);
nand U44668 (N_44668,N_44348,N_44097);
nor U44669 (N_44669,N_44182,N_44307);
nand U44670 (N_44670,N_44103,N_44105);
nand U44671 (N_44671,N_44092,N_44392);
nor U44672 (N_44672,N_44477,N_44333);
and U44673 (N_44673,N_44106,N_44161);
and U44674 (N_44674,N_44404,N_44446);
nor U44675 (N_44675,N_44036,N_44444);
nand U44676 (N_44676,N_44175,N_44261);
nand U44677 (N_44677,N_44169,N_44141);
nor U44678 (N_44678,N_44191,N_44000);
and U44679 (N_44679,N_44399,N_44315);
and U44680 (N_44680,N_44224,N_44335);
nor U44681 (N_44681,N_44147,N_44276);
nor U44682 (N_44682,N_44296,N_44359);
and U44683 (N_44683,N_44096,N_44066);
or U44684 (N_44684,N_44171,N_44071);
nor U44685 (N_44685,N_44455,N_44255);
nor U44686 (N_44686,N_44241,N_44489);
and U44687 (N_44687,N_44146,N_44029);
or U44688 (N_44688,N_44053,N_44330);
or U44689 (N_44689,N_44134,N_44378);
nor U44690 (N_44690,N_44342,N_44217);
nor U44691 (N_44691,N_44372,N_44239);
and U44692 (N_44692,N_44368,N_44144);
nor U44693 (N_44693,N_44102,N_44233);
nand U44694 (N_44694,N_44124,N_44417);
xor U44695 (N_44695,N_44484,N_44450);
nand U44696 (N_44696,N_44340,N_44034);
nand U44697 (N_44697,N_44187,N_44014);
or U44698 (N_44698,N_44302,N_44060);
nor U44699 (N_44699,N_44418,N_44065);
xor U44700 (N_44700,N_44270,N_44190);
nand U44701 (N_44701,N_44123,N_44140);
nand U44702 (N_44702,N_44113,N_44423);
and U44703 (N_44703,N_44119,N_44346);
nand U44704 (N_44704,N_44153,N_44458);
nor U44705 (N_44705,N_44409,N_44218);
and U44706 (N_44706,N_44165,N_44013);
or U44707 (N_44707,N_44328,N_44385);
xor U44708 (N_44708,N_44358,N_44180);
or U44709 (N_44709,N_44402,N_44394);
nor U44710 (N_44710,N_44220,N_44090);
nor U44711 (N_44711,N_44043,N_44357);
nand U44712 (N_44712,N_44380,N_44038);
nor U44713 (N_44713,N_44433,N_44332);
and U44714 (N_44714,N_44152,N_44215);
xnor U44715 (N_44715,N_44110,N_44361);
nor U44716 (N_44716,N_44322,N_44365);
or U44717 (N_44717,N_44059,N_44264);
and U44718 (N_44718,N_44371,N_44151);
or U44719 (N_44719,N_44046,N_44282);
or U44720 (N_44720,N_44173,N_44225);
xnor U44721 (N_44721,N_44193,N_44032);
xor U44722 (N_44722,N_44177,N_44244);
xor U44723 (N_44723,N_44184,N_44325);
and U44724 (N_44724,N_44427,N_44312);
and U44725 (N_44725,N_44183,N_44003);
and U44726 (N_44726,N_44305,N_44076);
xor U44727 (N_44727,N_44339,N_44247);
and U44728 (N_44728,N_44396,N_44205);
xnor U44729 (N_44729,N_44470,N_44256);
nand U44730 (N_44730,N_44115,N_44221);
and U44731 (N_44731,N_44237,N_44343);
and U44732 (N_44732,N_44352,N_44382);
nand U44733 (N_44733,N_44338,N_44166);
or U44734 (N_44734,N_44210,N_44316);
nor U44735 (N_44735,N_44148,N_44259);
nand U44736 (N_44736,N_44085,N_44005);
nand U44737 (N_44737,N_44001,N_44189);
or U44738 (N_44738,N_44483,N_44449);
nand U44739 (N_44739,N_44390,N_44112);
and U44740 (N_44740,N_44251,N_44168);
or U44741 (N_44741,N_44468,N_44176);
and U44742 (N_44742,N_44397,N_44081);
or U44743 (N_44743,N_44386,N_44159);
xnor U44744 (N_44744,N_44025,N_44356);
nor U44745 (N_44745,N_44383,N_44285);
and U44746 (N_44746,N_44079,N_44406);
nand U44747 (N_44747,N_44192,N_44196);
nand U44748 (N_44748,N_44223,N_44395);
or U44749 (N_44749,N_44042,N_44452);
and U44750 (N_44750,N_44176,N_44077);
nor U44751 (N_44751,N_44248,N_44223);
nand U44752 (N_44752,N_44301,N_44024);
and U44753 (N_44753,N_44050,N_44093);
and U44754 (N_44754,N_44219,N_44182);
nand U44755 (N_44755,N_44301,N_44294);
nor U44756 (N_44756,N_44152,N_44030);
nor U44757 (N_44757,N_44197,N_44496);
xor U44758 (N_44758,N_44200,N_44470);
or U44759 (N_44759,N_44093,N_44280);
nand U44760 (N_44760,N_44239,N_44471);
nand U44761 (N_44761,N_44215,N_44284);
or U44762 (N_44762,N_44134,N_44130);
nor U44763 (N_44763,N_44412,N_44061);
xnor U44764 (N_44764,N_44046,N_44315);
nand U44765 (N_44765,N_44288,N_44480);
nand U44766 (N_44766,N_44446,N_44032);
or U44767 (N_44767,N_44007,N_44466);
or U44768 (N_44768,N_44218,N_44068);
nor U44769 (N_44769,N_44120,N_44184);
or U44770 (N_44770,N_44040,N_44442);
nand U44771 (N_44771,N_44491,N_44338);
or U44772 (N_44772,N_44011,N_44078);
nor U44773 (N_44773,N_44116,N_44202);
nand U44774 (N_44774,N_44183,N_44316);
nand U44775 (N_44775,N_44123,N_44078);
and U44776 (N_44776,N_44293,N_44329);
nand U44777 (N_44777,N_44273,N_44479);
nand U44778 (N_44778,N_44112,N_44484);
nand U44779 (N_44779,N_44220,N_44207);
nor U44780 (N_44780,N_44097,N_44259);
nor U44781 (N_44781,N_44156,N_44342);
and U44782 (N_44782,N_44297,N_44068);
nand U44783 (N_44783,N_44030,N_44251);
nand U44784 (N_44784,N_44090,N_44140);
and U44785 (N_44785,N_44111,N_44203);
or U44786 (N_44786,N_44271,N_44432);
nand U44787 (N_44787,N_44472,N_44022);
and U44788 (N_44788,N_44212,N_44085);
xor U44789 (N_44789,N_44058,N_44378);
or U44790 (N_44790,N_44363,N_44171);
nor U44791 (N_44791,N_44107,N_44145);
or U44792 (N_44792,N_44338,N_44378);
xor U44793 (N_44793,N_44095,N_44272);
and U44794 (N_44794,N_44149,N_44290);
or U44795 (N_44795,N_44189,N_44386);
and U44796 (N_44796,N_44097,N_44190);
or U44797 (N_44797,N_44249,N_44239);
or U44798 (N_44798,N_44385,N_44046);
or U44799 (N_44799,N_44345,N_44298);
xnor U44800 (N_44800,N_44029,N_44115);
and U44801 (N_44801,N_44327,N_44410);
and U44802 (N_44802,N_44304,N_44073);
nand U44803 (N_44803,N_44476,N_44157);
xor U44804 (N_44804,N_44439,N_44307);
nand U44805 (N_44805,N_44155,N_44048);
or U44806 (N_44806,N_44004,N_44283);
xnor U44807 (N_44807,N_44189,N_44193);
or U44808 (N_44808,N_44234,N_44358);
or U44809 (N_44809,N_44045,N_44150);
nor U44810 (N_44810,N_44051,N_44181);
and U44811 (N_44811,N_44151,N_44313);
or U44812 (N_44812,N_44438,N_44190);
and U44813 (N_44813,N_44394,N_44104);
xnor U44814 (N_44814,N_44206,N_44402);
nor U44815 (N_44815,N_44119,N_44149);
or U44816 (N_44816,N_44215,N_44266);
and U44817 (N_44817,N_44020,N_44010);
and U44818 (N_44818,N_44402,N_44230);
xnor U44819 (N_44819,N_44498,N_44363);
xnor U44820 (N_44820,N_44416,N_44045);
nor U44821 (N_44821,N_44199,N_44484);
nor U44822 (N_44822,N_44059,N_44458);
xnor U44823 (N_44823,N_44204,N_44479);
or U44824 (N_44824,N_44160,N_44373);
nor U44825 (N_44825,N_44302,N_44097);
or U44826 (N_44826,N_44189,N_44404);
xnor U44827 (N_44827,N_44076,N_44463);
and U44828 (N_44828,N_44260,N_44199);
or U44829 (N_44829,N_44342,N_44040);
nor U44830 (N_44830,N_44054,N_44236);
or U44831 (N_44831,N_44392,N_44483);
and U44832 (N_44832,N_44452,N_44034);
xor U44833 (N_44833,N_44407,N_44185);
or U44834 (N_44834,N_44264,N_44281);
or U44835 (N_44835,N_44010,N_44058);
nand U44836 (N_44836,N_44461,N_44000);
nand U44837 (N_44837,N_44470,N_44344);
and U44838 (N_44838,N_44451,N_44433);
or U44839 (N_44839,N_44173,N_44420);
nand U44840 (N_44840,N_44285,N_44405);
nor U44841 (N_44841,N_44047,N_44281);
and U44842 (N_44842,N_44123,N_44272);
nand U44843 (N_44843,N_44405,N_44481);
and U44844 (N_44844,N_44495,N_44081);
nand U44845 (N_44845,N_44132,N_44341);
nand U44846 (N_44846,N_44028,N_44339);
and U44847 (N_44847,N_44454,N_44248);
or U44848 (N_44848,N_44174,N_44007);
or U44849 (N_44849,N_44149,N_44027);
nand U44850 (N_44850,N_44299,N_44188);
and U44851 (N_44851,N_44091,N_44303);
or U44852 (N_44852,N_44459,N_44206);
xor U44853 (N_44853,N_44464,N_44348);
nor U44854 (N_44854,N_44253,N_44209);
nand U44855 (N_44855,N_44308,N_44040);
and U44856 (N_44856,N_44471,N_44325);
or U44857 (N_44857,N_44130,N_44218);
and U44858 (N_44858,N_44486,N_44209);
nand U44859 (N_44859,N_44157,N_44278);
nor U44860 (N_44860,N_44265,N_44471);
nor U44861 (N_44861,N_44007,N_44258);
nand U44862 (N_44862,N_44400,N_44177);
nor U44863 (N_44863,N_44356,N_44369);
nand U44864 (N_44864,N_44210,N_44141);
nor U44865 (N_44865,N_44307,N_44216);
or U44866 (N_44866,N_44483,N_44342);
nand U44867 (N_44867,N_44275,N_44132);
xnor U44868 (N_44868,N_44011,N_44393);
nor U44869 (N_44869,N_44268,N_44061);
xnor U44870 (N_44870,N_44028,N_44476);
or U44871 (N_44871,N_44424,N_44028);
and U44872 (N_44872,N_44143,N_44137);
xnor U44873 (N_44873,N_44100,N_44275);
nor U44874 (N_44874,N_44345,N_44497);
nor U44875 (N_44875,N_44469,N_44111);
nor U44876 (N_44876,N_44398,N_44468);
nand U44877 (N_44877,N_44297,N_44436);
nor U44878 (N_44878,N_44044,N_44466);
and U44879 (N_44879,N_44370,N_44123);
xor U44880 (N_44880,N_44466,N_44201);
and U44881 (N_44881,N_44211,N_44370);
and U44882 (N_44882,N_44080,N_44230);
and U44883 (N_44883,N_44421,N_44096);
nand U44884 (N_44884,N_44080,N_44089);
nor U44885 (N_44885,N_44340,N_44207);
or U44886 (N_44886,N_44457,N_44129);
nand U44887 (N_44887,N_44155,N_44266);
and U44888 (N_44888,N_44334,N_44092);
and U44889 (N_44889,N_44423,N_44033);
and U44890 (N_44890,N_44252,N_44499);
and U44891 (N_44891,N_44397,N_44116);
or U44892 (N_44892,N_44230,N_44309);
nor U44893 (N_44893,N_44498,N_44257);
and U44894 (N_44894,N_44167,N_44218);
or U44895 (N_44895,N_44052,N_44077);
nand U44896 (N_44896,N_44084,N_44366);
and U44897 (N_44897,N_44317,N_44439);
xor U44898 (N_44898,N_44285,N_44362);
nand U44899 (N_44899,N_44326,N_44479);
nor U44900 (N_44900,N_44006,N_44047);
nor U44901 (N_44901,N_44164,N_44032);
nor U44902 (N_44902,N_44351,N_44475);
xor U44903 (N_44903,N_44035,N_44151);
and U44904 (N_44904,N_44318,N_44425);
or U44905 (N_44905,N_44197,N_44488);
and U44906 (N_44906,N_44052,N_44385);
nand U44907 (N_44907,N_44024,N_44175);
nand U44908 (N_44908,N_44130,N_44413);
nor U44909 (N_44909,N_44460,N_44301);
or U44910 (N_44910,N_44208,N_44444);
xor U44911 (N_44911,N_44177,N_44187);
nor U44912 (N_44912,N_44115,N_44134);
or U44913 (N_44913,N_44418,N_44309);
xnor U44914 (N_44914,N_44254,N_44285);
nand U44915 (N_44915,N_44091,N_44227);
or U44916 (N_44916,N_44187,N_44050);
nand U44917 (N_44917,N_44087,N_44370);
nor U44918 (N_44918,N_44049,N_44369);
nor U44919 (N_44919,N_44063,N_44026);
xnor U44920 (N_44920,N_44482,N_44374);
or U44921 (N_44921,N_44119,N_44067);
or U44922 (N_44922,N_44327,N_44097);
nor U44923 (N_44923,N_44498,N_44378);
and U44924 (N_44924,N_44259,N_44387);
nor U44925 (N_44925,N_44102,N_44083);
or U44926 (N_44926,N_44101,N_44330);
or U44927 (N_44927,N_44072,N_44181);
xor U44928 (N_44928,N_44312,N_44218);
xor U44929 (N_44929,N_44422,N_44447);
and U44930 (N_44930,N_44164,N_44343);
nor U44931 (N_44931,N_44351,N_44078);
and U44932 (N_44932,N_44121,N_44242);
and U44933 (N_44933,N_44408,N_44281);
and U44934 (N_44934,N_44393,N_44344);
and U44935 (N_44935,N_44493,N_44213);
nor U44936 (N_44936,N_44425,N_44139);
xnor U44937 (N_44937,N_44064,N_44384);
and U44938 (N_44938,N_44134,N_44261);
or U44939 (N_44939,N_44227,N_44093);
or U44940 (N_44940,N_44460,N_44414);
and U44941 (N_44941,N_44032,N_44264);
or U44942 (N_44942,N_44032,N_44141);
and U44943 (N_44943,N_44493,N_44200);
nand U44944 (N_44944,N_44248,N_44192);
nand U44945 (N_44945,N_44361,N_44339);
nor U44946 (N_44946,N_44259,N_44402);
nor U44947 (N_44947,N_44427,N_44065);
and U44948 (N_44948,N_44223,N_44098);
nor U44949 (N_44949,N_44158,N_44370);
nand U44950 (N_44950,N_44130,N_44476);
xor U44951 (N_44951,N_44121,N_44460);
xnor U44952 (N_44952,N_44312,N_44207);
and U44953 (N_44953,N_44423,N_44439);
and U44954 (N_44954,N_44100,N_44274);
or U44955 (N_44955,N_44207,N_44441);
and U44956 (N_44956,N_44085,N_44493);
or U44957 (N_44957,N_44248,N_44093);
nor U44958 (N_44958,N_44098,N_44203);
nor U44959 (N_44959,N_44387,N_44094);
or U44960 (N_44960,N_44141,N_44248);
nor U44961 (N_44961,N_44065,N_44461);
and U44962 (N_44962,N_44186,N_44253);
nand U44963 (N_44963,N_44405,N_44042);
nand U44964 (N_44964,N_44394,N_44332);
nand U44965 (N_44965,N_44037,N_44488);
and U44966 (N_44966,N_44173,N_44122);
or U44967 (N_44967,N_44199,N_44385);
and U44968 (N_44968,N_44409,N_44486);
nand U44969 (N_44969,N_44446,N_44289);
nor U44970 (N_44970,N_44254,N_44024);
or U44971 (N_44971,N_44420,N_44416);
xnor U44972 (N_44972,N_44217,N_44373);
nor U44973 (N_44973,N_44208,N_44363);
nor U44974 (N_44974,N_44356,N_44000);
nand U44975 (N_44975,N_44345,N_44122);
or U44976 (N_44976,N_44406,N_44233);
nor U44977 (N_44977,N_44040,N_44198);
nor U44978 (N_44978,N_44134,N_44329);
xor U44979 (N_44979,N_44208,N_44235);
and U44980 (N_44980,N_44433,N_44244);
and U44981 (N_44981,N_44234,N_44108);
nand U44982 (N_44982,N_44147,N_44198);
xnor U44983 (N_44983,N_44239,N_44384);
or U44984 (N_44984,N_44149,N_44442);
nand U44985 (N_44985,N_44026,N_44335);
nor U44986 (N_44986,N_44017,N_44222);
and U44987 (N_44987,N_44105,N_44169);
nor U44988 (N_44988,N_44122,N_44293);
nor U44989 (N_44989,N_44074,N_44271);
nor U44990 (N_44990,N_44274,N_44005);
or U44991 (N_44991,N_44210,N_44166);
and U44992 (N_44992,N_44422,N_44124);
nor U44993 (N_44993,N_44093,N_44032);
nor U44994 (N_44994,N_44043,N_44269);
and U44995 (N_44995,N_44353,N_44158);
nor U44996 (N_44996,N_44027,N_44315);
nor U44997 (N_44997,N_44115,N_44183);
and U44998 (N_44998,N_44478,N_44167);
nand U44999 (N_44999,N_44428,N_44122);
nor U45000 (N_45000,N_44637,N_44734);
or U45001 (N_45001,N_44612,N_44801);
nor U45002 (N_45002,N_44501,N_44769);
or U45003 (N_45003,N_44517,N_44756);
and U45004 (N_45004,N_44996,N_44736);
and U45005 (N_45005,N_44857,N_44726);
nor U45006 (N_45006,N_44840,N_44843);
or U45007 (N_45007,N_44969,N_44902);
nor U45008 (N_45008,N_44853,N_44896);
and U45009 (N_45009,N_44809,N_44936);
nand U45010 (N_45010,N_44695,N_44624);
nor U45011 (N_45011,N_44914,N_44674);
and U45012 (N_45012,N_44942,N_44689);
nand U45013 (N_45013,N_44865,N_44948);
and U45014 (N_45014,N_44753,N_44705);
xor U45015 (N_45015,N_44582,N_44974);
and U45016 (N_45016,N_44667,N_44503);
xnor U45017 (N_45017,N_44947,N_44589);
nand U45018 (N_45018,N_44623,N_44816);
nor U45019 (N_45019,N_44554,N_44610);
nand U45020 (N_45020,N_44613,N_44911);
or U45021 (N_45021,N_44876,N_44837);
and U45022 (N_45022,N_44549,N_44570);
and U45023 (N_45023,N_44930,N_44972);
nor U45024 (N_45024,N_44538,N_44609);
nor U45025 (N_45025,N_44791,N_44861);
or U45026 (N_45026,N_44891,N_44778);
and U45027 (N_45027,N_44761,N_44575);
xnor U45028 (N_45028,N_44619,N_44872);
nand U45029 (N_45029,N_44514,N_44714);
nand U45030 (N_45030,N_44710,N_44810);
or U45031 (N_45031,N_44656,N_44644);
nand U45032 (N_45032,N_44751,N_44935);
nand U45033 (N_45033,N_44924,N_44727);
xor U45034 (N_45034,N_44691,N_44713);
and U45035 (N_45035,N_44573,N_44544);
nand U45036 (N_45036,N_44627,N_44663);
and U45037 (N_45037,N_44817,N_44789);
nand U45038 (N_45038,N_44511,N_44963);
or U45039 (N_45039,N_44567,N_44708);
and U45040 (N_45040,N_44552,N_44550);
nor U45041 (N_45041,N_44966,N_44685);
xor U45042 (N_45042,N_44850,N_44533);
and U45043 (N_45043,N_44918,N_44529);
and U45044 (N_45044,N_44844,N_44693);
or U45045 (N_45045,N_44950,N_44956);
and U45046 (N_45046,N_44738,N_44621);
nand U45047 (N_45047,N_44615,N_44975);
or U45048 (N_45048,N_44586,N_44912);
and U45049 (N_45049,N_44939,N_44764);
nor U45050 (N_45050,N_44908,N_44907);
nor U45051 (N_45051,N_44639,N_44721);
nor U45052 (N_45052,N_44808,N_44945);
or U45053 (N_45053,N_44688,N_44718);
and U45054 (N_45054,N_44702,N_44715);
and U45055 (N_45055,N_44779,N_44851);
or U45056 (N_45056,N_44880,N_44811);
nand U45057 (N_45057,N_44804,N_44643);
or U45058 (N_45058,N_44704,N_44707);
nand U45059 (N_45059,N_44763,N_44893);
and U45060 (N_45060,N_44686,N_44913);
nand U45061 (N_45061,N_44988,N_44858);
and U45062 (N_45062,N_44992,N_44832);
nand U45063 (N_45063,N_44548,N_44971);
xor U45064 (N_45064,N_44754,N_44593);
or U45065 (N_45065,N_44668,N_44919);
xnor U45066 (N_45066,N_44722,N_44985);
and U45067 (N_45067,N_44827,N_44916);
or U45068 (N_45068,N_44968,N_44910);
and U45069 (N_45069,N_44759,N_44821);
xor U45070 (N_45070,N_44665,N_44525);
nor U45071 (N_45071,N_44894,N_44709);
or U45072 (N_45072,N_44859,N_44524);
xnor U45073 (N_45073,N_44530,N_44915);
or U45074 (N_45074,N_44711,N_44792);
nor U45075 (N_45075,N_44601,N_44635);
nor U45076 (N_45076,N_44505,N_44904);
and U45077 (N_45077,N_44502,N_44961);
nand U45078 (N_45078,N_44775,N_44599);
and U45079 (N_45079,N_44798,N_44871);
and U45080 (N_45080,N_44572,N_44760);
nor U45081 (N_45081,N_44606,N_44557);
or U45082 (N_45082,N_44826,N_44943);
nor U45083 (N_45083,N_44651,N_44855);
and U45084 (N_45084,N_44547,N_44854);
nor U45085 (N_45085,N_44700,N_44694);
or U45086 (N_45086,N_44692,N_44928);
nor U45087 (N_45087,N_44820,N_44576);
nand U45088 (N_45088,N_44542,N_44531);
xnor U45089 (N_45089,N_44541,N_44574);
and U45090 (N_45090,N_44981,N_44927);
nor U45091 (N_45091,N_44881,N_44720);
and U45092 (N_45092,N_44535,N_44946);
or U45093 (N_45093,N_44781,N_44829);
or U45094 (N_45094,N_44890,N_44560);
or U45095 (N_45095,N_44770,N_44706);
and U45096 (N_45096,N_44757,N_44540);
nor U45097 (N_45097,N_44940,N_44578);
or U45098 (N_45098,N_44579,N_44640);
nor U45099 (N_45099,N_44614,N_44551);
or U45100 (N_45100,N_44648,N_44543);
nand U45101 (N_45101,N_44521,N_44841);
xor U45102 (N_45102,N_44799,N_44933);
and U45103 (N_45103,N_44508,N_44958);
nor U45104 (N_45104,N_44500,N_44645);
nor U45105 (N_45105,N_44863,N_44980);
nor U45106 (N_45106,N_44660,N_44553);
or U45107 (N_45107,N_44681,N_44874);
nand U45108 (N_45108,N_44546,N_44744);
nor U45109 (N_45109,N_44955,N_44617);
nand U45110 (N_45110,N_44938,N_44828);
nand U45111 (N_45111,N_44979,N_44815);
nand U45112 (N_45112,N_44717,N_44602);
nor U45113 (N_45113,N_44766,N_44862);
nand U45114 (N_45114,N_44830,N_44735);
and U45115 (N_45115,N_44959,N_44802);
nand U45116 (N_45116,N_44646,N_44989);
and U45117 (N_45117,N_44847,N_44604);
or U45118 (N_45118,N_44733,N_44783);
nor U45119 (N_45119,N_44953,N_44591);
nor U45120 (N_45120,N_44728,N_44537);
and U45121 (N_45121,N_44678,N_44774);
nor U45122 (N_45122,N_44558,N_44747);
nor U45123 (N_45123,N_44776,N_44510);
and U45124 (N_45124,N_44905,N_44730);
nand U45125 (N_45125,N_44937,N_44993);
or U45126 (N_45126,N_44750,N_44539);
nor U45127 (N_45127,N_44994,N_44903);
and U45128 (N_45128,N_44749,N_44683);
nor U45129 (N_45129,N_44528,N_44941);
and U45130 (N_45130,N_44823,N_44818);
nor U45131 (N_45131,N_44836,N_44527);
or U45132 (N_45132,N_44856,N_44745);
nor U45133 (N_45133,N_44906,N_44677);
nand U45134 (N_45134,N_44931,N_44620);
nand U45135 (N_45135,N_44652,N_44765);
nor U45136 (N_45136,N_44703,N_44864);
and U45137 (N_45137,N_44509,N_44957);
or U45138 (N_45138,N_44831,N_44842);
nor U45139 (N_45139,N_44987,N_44687);
xnor U45140 (N_45140,N_44867,N_44625);
nand U45141 (N_45141,N_44632,N_44951);
xor U45142 (N_45142,N_44676,N_44852);
nor U45143 (N_45143,N_44900,N_44504);
nand U45144 (N_45144,N_44565,N_44921);
nand U45145 (N_45145,N_44679,N_44748);
or U45146 (N_45146,N_44690,N_44696);
or U45147 (N_45147,N_44870,N_44636);
and U45148 (N_45148,N_44898,N_44559);
nand U45149 (N_45149,N_44758,N_44659);
nor U45150 (N_45150,N_44655,N_44526);
and U45151 (N_45151,N_44569,N_44534);
and U45152 (N_45152,N_44712,N_44922);
xor U45153 (N_45153,N_44807,N_44628);
and U45154 (N_45154,N_44650,N_44884);
nand U45155 (N_45155,N_44675,N_44658);
or U45156 (N_45156,N_44622,N_44653);
or U45157 (N_45157,N_44944,N_44556);
xnor U45158 (N_45158,N_44768,N_44773);
nand U45159 (N_45159,N_44897,N_44767);
nor U45160 (N_45160,N_44697,N_44752);
nand U45161 (N_45161,N_44608,N_44630);
and U45162 (N_45162,N_44782,N_44724);
nor U45163 (N_45163,N_44568,N_44866);
or U45164 (N_45164,N_44626,N_44607);
nand U45165 (N_45165,N_44869,N_44596);
and U45166 (N_45166,N_44684,N_44555);
and U45167 (N_45167,N_44885,N_44592);
nand U45168 (N_45168,N_44984,N_44846);
or U45169 (N_45169,N_44729,N_44584);
xnor U45170 (N_45170,N_44633,N_44520);
nor U45171 (N_45171,N_44616,N_44699);
or U45172 (N_45172,N_44732,N_44701);
xnor U45173 (N_45173,N_44800,N_44895);
and U45174 (N_45174,N_44682,N_44824);
or U45175 (N_45175,N_44967,N_44641);
or U45176 (N_45176,N_44670,N_44848);
nand U45177 (N_45177,N_44962,N_44631);
xor U45178 (N_45178,N_44562,N_44666);
nor U45179 (N_45179,N_44597,N_44788);
and U45180 (N_45180,N_44999,N_44673);
and U45181 (N_45181,N_44965,N_44875);
xnor U45182 (N_45182,N_44545,N_44977);
or U45183 (N_45183,N_44739,N_44581);
nand U45184 (N_45184,N_44796,N_44901);
nor U45185 (N_45185,N_44507,N_44585);
nor U45186 (N_45186,N_44882,N_44838);
nand U45187 (N_45187,N_44762,N_44519);
or U45188 (N_45188,N_44588,N_44982);
or U45189 (N_45189,N_44970,N_44834);
nand U45190 (N_45190,N_44794,N_44662);
or U45191 (N_45191,N_44883,N_44932);
or U45192 (N_45192,N_44803,N_44649);
nand U45193 (N_45193,N_44522,N_44923);
or U45194 (N_45194,N_44719,N_44731);
or U45195 (N_45195,N_44642,N_44580);
nand U45196 (N_45196,N_44600,N_44998);
nand U45197 (N_45197,N_44671,N_44638);
nor U45198 (N_45198,N_44629,N_44755);
or U45199 (N_45199,N_44813,N_44990);
nor U45200 (N_45200,N_44669,N_44909);
xor U45201 (N_45201,N_44786,N_44949);
or U45202 (N_45202,N_44849,N_44716);
nor U45203 (N_45203,N_44805,N_44860);
and U45204 (N_45204,N_44892,N_44563);
nor U45205 (N_45205,N_44790,N_44571);
nand U45206 (N_45206,N_44879,N_44618);
and U45207 (N_45207,N_44973,N_44743);
nand U45208 (N_45208,N_44536,N_44925);
nand U45209 (N_45209,N_44594,N_44784);
and U45210 (N_45210,N_44513,N_44845);
and U45211 (N_45211,N_44587,N_44780);
xor U45212 (N_45212,N_44839,N_44583);
or U45213 (N_45213,N_44833,N_44888);
nor U45214 (N_45214,N_44917,N_44952);
or U45215 (N_45215,N_44590,N_44523);
nor U45216 (N_45216,N_44934,N_44723);
nor U45217 (N_45217,N_44672,N_44986);
and U45218 (N_45218,N_44577,N_44611);
nor U45219 (N_45219,N_44777,N_44899);
and U45220 (N_45220,N_44868,N_44983);
and U45221 (N_45221,N_44825,N_44877);
or U45222 (N_45222,N_44664,N_44741);
nor U45223 (N_45223,N_44680,N_44746);
nor U45224 (N_45224,N_44835,N_44566);
and U45225 (N_45225,N_44926,N_44995);
or U45226 (N_45226,N_44997,N_44742);
and U45227 (N_45227,N_44819,N_44561);
or U45228 (N_45228,N_44797,N_44772);
or U45229 (N_45229,N_44814,N_44920);
nand U45230 (N_45230,N_44506,N_44806);
xnor U45231 (N_45231,N_44740,N_44991);
xor U45232 (N_45232,N_44964,N_44605);
xor U45233 (N_45233,N_44878,N_44598);
or U45234 (N_45234,N_44725,N_44603);
and U45235 (N_45235,N_44793,N_44516);
or U45236 (N_45236,N_44889,N_44795);
and U45237 (N_45237,N_44978,N_44518);
nor U45238 (N_45238,N_44886,N_44512);
nor U45239 (N_45239,N_44785,N_44698);
and U45240 (N_45240,N_44929,N_44661);
nand U45241 (N_45241,N_44873,N_44532);
or U45242 (N_45242,N_44654,N_44887);
nor U45243 (N_45243,N_44657,N_44737);
or U45244 (N_45244,N_44822,N_44564);
nand U45245 (N_45245,N_44515,N_44787);
nand U45246 (N_45246,N_44954,N_44960);
nor U45247 (N_45247,N_44976,N_44595);
or U45248 (N_45248,N_44771,N_44634);
or U45249 (N_45249,N_44647,N_44812);
nor U45250 (N_45250,N_44964,N_44843);
nor U45251 (N_45251,N_44857,N_44932);
nand U45252 (N_45252,N_44832,N_44984);
nor U45253 (N_45253,N_44641,N_44727);
and U45254 (N_45254,N_44643,N_44953);
nor U45255 (N_45255,N_44844,N_44853);
nor U45256 (N_45256,N_44941,N_44737);
and U45257 (N_45257,N_44567,N_44774);
and U45258 (N_45258,N_44723,N_44990);
nand U45259 (N_45259,N_44746,N_44566);
xor U45260 (N_45260,N_44649,N_44572);
and U45261 (N_45261,N_44954,N_44862);
nor U45262 (N_45262,N_44859,N_44769);
nand U45263 (N_45263,N_44793,N_44584);
or U45264 (N_45264,N_44814,N_44940);
nand U45265 (N_45265,N_44711,N_44745);
nor U45266 (N_45266,N_44705,N_44590);
nor U45267 (N_45267,N_44934,N_44786);
xor U45268 (N_45268,N_44701,N_44550);
nand U45269 (N_45269,N_44832,N_44556);
and U45270 (N_45270,N_44903,N_44889);
and U45271 (N_45271,N_44586,N_44719);
nor U45272 (N_45272,N_44600,N_44922);
nand U45273 (N_45273,N_44858,N_44665);
or U45274 (N_45274,N_44769,N_44605);
xor U45275 (N_45275,N_44697,N_44820);
or U45276 (N_45276,N_44962,N_44959);
xor U45277 (N_45277,N_44588,N_44573);
nor U45278 (N_45278,N_44916,N_44559);
or U45279 (N_45279,N_44867,N_44778);
and U45280 (N_45280,N_44912,N_44527);
or U45281 (N_45281,N_44894,N_44770);
nor U45282 (N_45282,N_44677,N_44926);
nand U45283 (N_45283,N_44942,N_44658);
nand U45284 (N_45284,N_44526,N_44947);
nor U45285 (N_45285,N_44931,N_44519);
nor U45286 (N_45286,N_44924,N_44669);
xor U45287 (N_45287,N_44796,N_44768);
nand U45288 (N_45288,N_44520,N_44879);
and U45289 (N_45289,N_44678,N_44846);
and U45290 (N_45290,N_44828,N_44819);
nand U45291 (N_45291,N_44944,N_44609);
nor U45292 (N_45292,N_44702,N_44939);
and U45293 (N_45293,N_44928,N_44648);
and U45294 (N_45294,N_44719,N_44822);
nor U45295 (N_45295,N_44568,N_44786);
nor U45296 (N_45296,N_44855,N_44866);
nor U45297 (N_45297,N_44627,N_44508);
nor U45298 (N_45298,N_44725,N_44556);
and U45299 (N_45299,N_44648,N_44828);
or U45300 (N_45300,N_44980,N_44997);
nand U45301 (N_45301,N_44776,N_44997);
or U45302 (N_45302,N_44517,N_44699);
nor U45303 (N_45303,N_44624,N_44585);
xor U45304 (N_45304,N_44774,N_44892);
or U45305 (N_45305,N_44737,N_44730);
or U45306 (N_45306,N_44902,N_44709);
nand U45307 (N_45307,N_44846,N_44651);
nand U45308 (N_45308,N_44527,N_44573);
or U45309 (N_45309,N_44600,N_44729);
or U45310 (N_45310,N_44549,N_44920);
or U45311 (N_45311,N_44994,N_44546);
xor U45312 (N_45312,N_44836,N_44792);
and U45313 (N_45313,N_44611,N_44813);
or U45314 (N_45314,N_44928,N_44640);
or U45315 (N_45315,N_44559,N_44965);
nand U45316 (N_45316,N_44974,N_44526);
or U45317 (N_45317,N_44965,N_44734);
or U45318 (N_45318,N_44905,N_44725);
nand U45319 (N_45319,N_44810,N_44592);
nor U45320 (N_45320,N_44964,N_44807);
or U45321 (N_45321,N_44664,N_44938);
and U45322 (N_45322,N_44803,N_44855);
and U45323 (N_45323,N_44678,N_44837);
nand U45324 (N_45324,N_44962,N_44930);
nand U45325 (N_45325,N_44610,N_44519);
nor U45326 (N_45326,N_44898,N_44582);
nand U45327 (N_45327,N_44748,N_44883);
nor U45328 (N_45328,N_44690,N_44847);
nand U45329 (N_45329,N_44811,N_44935);
nor U45330 (N_45330,N_44856,N_44679);
nor U45331 (N_45331,N_44886,N_44586);
xnor U45332 (N_45332,N_44936,N_44943);
nor U45333 (N_45333,N_44772,N_44699);
and U45334 (N_45334,N_44806,N_44764);
or U45335 (N_45335,N_44641,N_44916);
or U45336 (N_45336,N_44678,N_44906);
nor U45337 (N_45337,N_44854,N_44544);
and U45338 (N_45338,N_44598,N_44866);
or U45339 (N_45339,N_44667,N_44652);
or U45340 (N_45340,N_44889,N_44785);
or U45341 (N_45341,N_44609,N_44913);
xnor U45342 (N_45342,N_44563,N_44777);
or U45343 (N_45343,N_44836,N_44811);
nand U45344 (N_45344,N_44781,N_44559);
and U45345 (N_45345,N_44764,N_44908);
nand U45346 (N_45346,N_44819,N_44734);
and U45347 (N_45347,N_44764,N_44547);
xor U45348 (N_45348,N_44508,N_44813);
nand U45349 (N_45349,N_44696,N_44742);
and U45350 (N_45350,N_44553,N_44706);
nor U45351 (N_45351,N_44709,N_44726);
nor U45352 (N_45352,N_44806,N_44800);
xnor U45353 (N_45353,N_44863,N_44629);
xnor U45354 (N_45354,N_44998,N_44539);
nand U45355 (N_45355,N_44660,N_44578);
nand U45356 (N_45356,N_44732,N_44896);
and U45357 (N_45357,N_44753,N_44514);
and U45358 (N_45358,N_44876,N_44647);
xor U45359 (N_45359,N_44708,N_44713);
nand U45360 (N_45360,N_44976,N_44599);
nor U45361 (N_45361,N_44761,N_44883);
nand U45362 (N_45362,N_44572,N_44605);
and U45363 (N_45363,N_44553,N_44564);
and U45364 (N_45364,N_44837,N_44743);
or U45365 (N_45365,N_44685,N_44965);
or U45366 (N_45366,N_44942,N_44991);
nor U45367 (N_45367,N_44811,N_44563);
nand U45368 (N_45368,N_44733,N_44655);
nand U45369 (N_45369,N_44827,N_44922);
and U45370 (N_45370,N_44683,N_44626);
and U45371 (N_45371,N_44676,N_44844);
or U45372 (N_45372,N_44518,N_44809);
nand U45373 (N_45373,N_44678,N_44798);
nor U45374 (N_45374,N_44674,N_44763);
nor U45375 (N_45375,N_44618,N_44596);
nor U45376 (N_45376,N_44534,N_44597);
nand U45377 (N_45377,N_44722,N_44906);
and U45378 (N_45378,N_44686,N_44962);
xor U45379 (N_45379,N_44983,N_44747);
and U45380 (N_45380,N_44809,N_44565);
nor U45381 (N_45381,N_44747,N_44599);
and U45382 (N_45382,N_44847,N_44963);
nand U45383 (N_45383,N_44598,N_44839);
nor U45384 (N_45384,N_44738,N_44778);
or U45385 (N_45385,N_44849,N_44773);
nor U45386 (N_45386,N_44726,N_44887);
or U45387 (N_45387,N_44725,N_44740);
nand U45388 (N_45388,N_44676,N_44711);
and U45389 (N_45389,N_44587,N_44974);
and U45390 (N_45390,N_44739,N_44725);
xnor U45391 (N_45391,N_44622,N_44518);
and U45392 (N_45392,N_44823,N_44967);
nand U45393 (N_45393,N_44932,N_44563);
or U45394 (N_45394,N_44867,N_44826);
nor U45395 (N_45395,N_44627,N_44879);
xor U45396 (N_45396,N_44751,N_44708);
nor U45397 (N_45397,N_44867,N_44974);
or U45398 (N_45398,N_44513,N_44871);
and U45399 (N_45399,N_44582,N_44910);
nor U45400 (N_45400,N_44675,N_44960);
nor U45401 (N_45401,N_44864,N_44755);
or U45402 (N_45402,N_44944,N_44872);
nor U45403 (N_45403,N_44578,N_44711);
or U45404 (N_45404,N_44639,N_44837);
or U45405 (N_45405,N_44648,N_44813);
nor U45406 (N_45406,N_44937,N_44697);
or U45407 (N_45407,N_44622,N_44860);
or U45408 (N_45408,N_44821,N_44619);
nand U45409 (N_45409,N_44679,N_44927);
or U45410 (N_45410,N_44584,N_44861);
nand U45411 (N_45411,N_44554,N_44596);
and U45412 (N_45412,N_44993,N_44938);
and U45413 (N_45413,N_44855,N_44777);
and U45414 (N_45414,N_44729,N_44722);
or U45415 (N_45415,N_44502,N_44963);
nand U45416 (N_45416,N_44821,N_44769);
nand U45417 (N_45417,N_44861,N_44852);
nand U45418 (N_45418,N_44767,N_44748);
nor U45419 (N_45419,N_44701,N_44747);
or U45420 (N_45420,N_44866,N_44741);
nor U45421 (N_45421,N_44696,N_44998);
or U45422 (N_45422,N_44575,N_44711);
nor U45423 (N_45423,N_44639,N_44558);
nor U45424 (N_45424,N_44582,N_44516);
nand U45425 (N_45425,N_44622,N_44691);
xor U45426 (N_45426,N_44887,N_44511);
nand U45427 (N_45427,N_44730,N_44918);
or U45428 (N_45428,N_44793,N_44541);
nand U45429 (N_45429,N_44975,N_44651);
nand U45430 (N_45430,N_44922,N_44853);
nand U45431 (N_45431,N_44953,N_44504);
and U45432 (N_45432,N_44995,N_44647);
nor U45433 (N_45433,N_44619,N_44838);
nand U45434 (N_45434,N_44683,N_44902);
and U45435 (N_45435,N_44533,N_44683);
and U45436 (N_45436,N_44797,N_44835);
or U45437 (N_45437,N_44564,N_44838);
or U45438 (N_45438,N_44687,N_44523);
nor U45439 (N_45439,N_44542,N_44732);
or U45440 (N_45440,N_44916,N_44736);
or U45441 (N_45441,N_44631,N_44587);
nor U45442 (N_45442,N_44587,N_44795);
xnor U45443 (N_45443,N_44940,N_44710);
nand U45444 (N_45444,N_44954,N_44901);
or U45445 (N_45445,N_44787,N_44512);
or U45446 (N_45446,N_44561,N_44726);
and U45447 (N_45447,N_44972,N_44739);
or U45448 (N_45448,N_44917,N_44928);
and U45449 (N_45449,N_44730,N_44575);
nand U45450 (N_45450,N_44949,N_44953);
nand U45451 (N_45451,N_44798,N_44758);
xnor U45452 (N_45452,N_44559,N_44800);
xor U45453 (N_45453,N_44868,N_44791);
and U45454 (N_45454,N_44601,N_44849);
and U45455 (N_45455,N_44512,N_44740);
or U45456 (N_45456,N_44539,N_44643);
nand U45457 (N_45457,N_44766,N_44709);
and U45458 (N_45458,N_44603,N_44865);
nand U45459 (N_45459,N_44733,N_44880);
and U45460 (N_45460,N_44591,N_44680);
nand U45461 (N_45461,N_44708,N_44626);
nor U45462 (N_45462,N_44738,N_44830);
nand U45463 (N_45463,N_44595,N_44898);
or U45464 (N_45464,N_44929,N_44623);
nand U45465 (N_45465,N_44536,N_44746);
or U45466 (N_45466,N_44636,N_44763);
and U45467 (N_45467,N_44615,N_44580);
xnor U45468 (N_45468,N_44934,N_44623);
nand U45469 (N_45469,N_44834,N_44839);
nor U45470 (N_45470,N_44819,N_44664);
nor U45471 (N_45471,N_44801,N_44898);
nor U45472 (N_45472,N_44679,N_44913);
and U45473 (N_45473,N_44920,N_44835);
and U45474 (N_45474,N_44967,N_44998);
or U45475 (N_45475,N_44643,N_44652);
nand U45476 (N_45476,N_44948,N_44789);
nand U45477 (N_45477,N_44585,N_44570);
xnor U45478 (N_45478,N_44747,N_44790);
and U45479 (N_45479,N_44652,N_44751);
nand U45480 (N_45480,N_44629,N_44675);
nor U45481 (N_45481,N_44977,N_44896);
nand U45482 (N_45482,N_44696,N_44997);
nor U45483 (N_45483,N_44716,N_44617);
nand U45484 (N_45484,N_44706,N_44724);
nand U45485 (N_45485,N_44524,N_44935);
nor U45486 (N_45486,N_44868,N_44771);
or U45487 (N_45487,N_44819,N_44641);
nand U45488 (N_45488,N_44709,N_44864);
nor U45489 (N_45489,N_44953,N_44542);
or U45490 (N_45490,N_44933,N_44964);
and U45491 (N_45491,N_44947,N_44766);
nor U45492 (N_45492,N_44880,N_44676);
or U45493 (N_45493,N_44661,N_44663);
and U45494 (N_45494,N_44700,N_44807);
or U45495 (N_45495,N_44807,N_44714);
or U45496 (N_45496,N_44578,N_44543);
xor U45497 (N_45497,N_44519,N_44999);
xor U45498 (N_45498,N_44556,N_44667);
or U45499 (N_45499,N_44592,N_44930);
xnor U45500 (N_45500,N_45475,N_45400);
nor U45501 (N_45501,N_45288,N_45256);
xnor U45502 (N_45502,N_45272,N_45432);
nand U45503 (N_45503,N_45042,N_45154);
nand U45504 (N_45504,N_45248,N_45457);
nand U45505 (N_45505,N_45287,N_45341);
or U45506 (N_45506,N_45397,N_45009);
xnor U45507 (N_45507,N_45347,N_45442);
and U45508 (N_45508,N_45132,N_45307);
nand U45509 (N_45509,N_45447,N_45234);
or U45510 (N_45510,N_45486,N_45119);
or U45511 (N_45511,N_45122,N_45253);
nand U45512 (N_45512,N_45106,N_45446);
xor U45513 (N_45513,N_45394,N_45322);
or U45514 (N_45514,N_45359,N_45043);
or U45515 (N_45515,N_45167,N_45343);
nor U45516 (N_45516,N_45279,N_45164);
and U45517 (N_45517,N_45003,N_45078);
and U45518 (N_45518,N_45216,N_45222);
and U45519 (N_45519,N_45246,N_45024);
nand U45520 (N_45520,N_45040,N_45054);
and U45521 (N_45521,N_45370,N_45384);
and U45522 (N_45522,N_45239,N_45252);
nand U45523 (N_45523,N_45381,N_45278);
xor U45524 (N_45524,N_45152,N_45057);
and U45525 (N_45525,N_45125,N_45342);
or U45526 (N_45526,N_45490,N_45206);
nand U45527 (N_45527,N_45310,N_45076);
nor U45528 (N_45528,N_45443,N_45380);
nor U45529 (N_45529,N_45315,N_45105);
xnor U45530 (N_45530,N_45297,N_45464);
and U45531 (N_45531,N_45022,N_45335);
or U45532 (N_45532,N_45188,N_45023);
nand U45533 (N_45533,N_45033,N_45103);
nor U45534 (N_45534,N_45079,N_45269);
nand U45535 (N_45535,N_45485,N_45146);
nor U45536 (N_45536,N_45088,N_45428);
nand U45537 (N_45537,N_45226,N_45121);
or U45538 (N_45538,N_45469,N_45371);
nand U45539 (N_45539,N_45179,N_45283);
nand U45540 (N_45540,N_45368,N_45113);
nand U45541 (N_45541,N_45026,N_45271);
xor U45542 (N_45542,N_45494,N_45225);
nand U45543 (N_45543,N_45006,N_45449);
nand U45544 (N_45544,N_45237,N_45431);
or U45545 (N_45545,N_45410,N_45210);
and U45546 (N_45546,N_45203,N_45304);
xor U45547 (N_45547,N_45060,N_45492);
nor U45548 (N_45548,N_45015,N_45092);
or U45549 (N_45549,N_45392,N_45221);
nand U45550 (N_45550,N_45481,N_45251);
or U45551 (N_45551,N_45303,N_45047);
xor U45552 (N_45552,N_45171,N_45120);
nand U45553 (N_45553,N_45429,N_45032);
nor U45554 (N_45554,N_45435,N_45476);
and U45555 (N_45555,N_45405,N_45067);
and U45556 (N_45556,N_45451,N_45366);
nor U45557 (N_45557,N_45369,N_45401);
and U45558 (N_45558,N_45455,N_45138);
and U45559 (N_45559,N_45045,N_45019);
xnor U45560 (N_45560,N_45229,N_45326);
and U45561 (N_45561,N_45161,N_45263);
and U45562 (N_45562,N_45391,N_45069);
and U45563 (N_45563,N_45160,N_45056);
nand U45564 (N_45564,N_45478,N_45150);
nand U45565 (N_45565,N_45220,N_45257);
and U45566 (N_45566,N_45261,N_45089);
and U45567 (N_45567,N_45389,N_45487);
nand U45568 (N_45568,N_45127,N_45036);
nor U45569 (N_45569,N_45174,N_45473);
and U45570 (N_45570,N_45240,N_45149);
nor U45571 (N_45571,N_45004,N_45095);
and U45572 (N_45572,N_45465,N_45354);
or U45573 (N_45573,N_45139,N_45173);
and U45574 (N_45574,N_45129,N_45262);
nand U45575 (N_45575,N_45403,N_45218);
or U45576 (N_45576,N_45099,N_45062);
and U45577 (N_45577,N_45055,N_45250);
xnor U45578 (N_45578,N_45409,N_45367);
nor U45579 (N_45579,N_45274,N_45422);
nor U45580 (N_45580,N_45375,N_45363);
nor U45581 (N_45581,N_45123,N_45355);
and U45582 (N_45582,N_45273,N_45499);
nor U45583 (N_45583,N_45365,N_45339);
xor U45584 (N_45584,N_45166,N_45493);
and U45585 (N_45585,N_45267,N_45109);
and U45586 (N_45586,N_45311,N_45461);
or U45587 (N_45587,N_45323,N_45212);
nor U45588 (N_45588,N_45051,N_45030);
nand U45589 (N_45589,N_45200,N_45104);
and U45590 (N_45590,N_45018,N_45414);
and U45591 (N_45591,N_45411,N_45087);
and U45592 (N_45592,N_45080,N_45471);
or U45593 (N_45593,N_45313,N_45198);
and U45594 (N_45594,N_45412,N_45182);
xnor U45595 (N_45595,N_45285,N_45223);
xor U45596 (N_45596,N_45268,N_45007);
and U45597 (N_45597,N_45197,N_45484);
and U45598 (N_45598,N_45034,N_45420);
nand U45599 (N_45599,N_45141,N_45002);
nor U45600 (N_45600,N_45314,N_45333);
and U45601 (N_45601,N_45144,N_45390);
xor U45602 (N_45602,N_45441,N_45011);
or U45603 (N_45603,N_45387,N_45438);
nor U45604 (N_45604,N_45459,N_45230);
nor U45605 (N_45605,N_45112,N_45479);
or U45606 (N_45606,N_45180,N_45421);
or U45607 (N_45607,N_45100,N_45065);
xnor U45608 (N_45608,N_45488,N_45136);
nand U45609 (N_45609,N_45094,N_45340);
or U45610 (N_45610,N_45172,N_45073);
and U45611 (N_45611,N_45417,N_45037);
nand U45612 (N_45612,N_45114,N_45133);
nor U45613 (N_45613,N_45027,N_45110);
nor U45614 (N_45614,N_45298,N_45168);
xor U45615 (N_45615,N_45000,N_45423);
and U45616 (N_45616,N_45338,N_45301);
and U45617 (N_45617,N_45293,N_45299);
and U45618 (N_45618,N_45372,N_45064);
nor U45619 (N_45619,N_45021,N_45107);
or U45620 (N_45620,N_45068,N_45005);
nor U45621 (N_45621,N_45195,N_45497);
nor U45622 (N_45622,N_45190,N_45059);
and U45623 (N_45623,N_45482,N_45352);
nand U45624 (N_45624,N_45091,N_45491);
or U45625 (N_45625,N_45325,N_45332);
and U45626 (N_45626,N_45102,N_45219);
or U45627 (N_45627,N_45440,N_45427);
and U45628 (N_45628,N_45364,N_45344);
or U45629 (N_45629,N_45258,N_45236);
nand U45630 (N_45630,N_45238,N_45450);
nor U45631 (N_45631,N_45290,N_45467);
and U45632 (N_45632,N_45373,N_45181);
nand U45633 (N_45633,N_45483,N_45463);
and U45634 (N_45634,N_45124,N_45437);
nor U45635 (N_45635,N_45187,N_45264);
or U45636 (N_45636,N_45406,N_45202);
or U45637 (N_45637,N_45118,N_45041);
nand U45638 (N_45638,N_45211,N_45477);
nand U45639 (N_45639,N_45385,N_45439);
nor U45640 (N_45640,N_45312,N_45294);
nand U45641 (N_45641,N_45194,N_45134);
nor U45642 (N_45642,N_45362,N_45353);
nor U45643 (N_45643,N_45075,N_45308);
nand U45644 (N_45644,N_45396,N_45193);
or U45645 (N_45645,N_45292,N_45346);
or U45646 (N_45646,N_45241,N_45012);
nand U45647 (N_45647,N_45334,N_45260);
nor U45648 (N_45648,N_45245,N_45151);
xor U45649 (N_45649,N_45291,N_45213);
and U45650 (N_45650,N_45046,N_45386);
and U45651 (N_45651,N_45016,N_45472);
xnor U45652 (N_45652,N_45281,N_45084);
nor U45653 (N_45653,N_45070,N_45498);
nand U45654 (N_45654,N_45399,N_45214);
and U45655 (N_45655,N_45284,N_45135);
or U45656 (N_45656,N_45327,N_45224);
nand U45657 (N_45657,N_45116,N_45044);
or U45658 (N_45658,N_45300,N_45331);
or U45659 (N_45659,N_45205,N_45408);
xnor U45660 (N_45660,N_45014,N_45207);
or U45661 (N_45661,N_45480,N_45117);
nor U45662 (N_45662,N_45081,N_45317);
or U45663 (N_45663,N_45376,N_45407);
or U45664 (N_45664,N_45382,N_45178);
nand U45665 (N_45665,N_45128,N_45445);
nand U45666 (N_45666,N_45413,N_45242);
or U45667 (N_45667,N_45316,N_45066);
nor U45668 (N_45668,N_45048,N_45458);
nor U45669 (N_45669,N_45177,N_45115);
nand U45670 (N_45670,N_45402,N_45192);
or U45671 (N_45671,N_45130,N_45049);
nand U45672 (N_45672,N_45145,N_45039);
or U45673 (N_45673,N_45277,N_45415);
xor U45674 (N_45674,N_45108,N_45061);
and U45675 (N_45675,N_45148,N_45289);
or U45676 (N_45676,N_45013,N_45474);
nand U45677 (N_45677,N_45282,N_45140);
or U45678 (N_45678,N_45286,N_45319);
nand U45679 (N_45679,N_45495,N_45184);
nor U45680 (N_45680,N_45489,N_45183);
nor U45681 (N_45681,N_45157,N_45378);
nor U45682 (N_45682,N_45466,N_45433);
nand U45683 (N_45683,N_45001,N_45419);
nor U45684 (N_45684,N_45320,N_45086);
nand U45685 (N_45685,N_45204,N_45008);
xor U45686 (N_45686,N_45452,N_45017);
nor U45687 (N_45687,N_45383,N_45053);
nor U45688 (N_45688,N_45085,N_45050);
nor U45689 (N_45689,N_45275,N_45328);
or U45690 (N_45690,N_45444,N_45404);
or U45691 (N_45691,N_45361,N_45093);
nand U45692 (N_45692,N_45345,N_45097);
nor U45693 (N_45693,N_45233,N_45058);
nand U45694 (N_45694,N_45096,N_45176);
xor U45695 (N_45695,N_45156,N_45249);
nor U45696 (N_45696,N_45031,N_45425);
nand U45697 (N_45697,N_45351,N_45227);
nand U45698 (N_45698,N_45159,N_45185);
nand U45699 (N_45699,N_45337,N_45169);
nor U45700 (N_45700,N_45254,N_45426);
nand U45701 (N_45701,N_45416,N_45191);
nand U45702 (N_45702,N_45357,N_45374);
nand U45703 (N_45703,N_45052,N_45215);
or U45704 (N_45704,N_45083,N_45235);
nand U45705 (N_45705,N_45077,N_45462);
and U45706 (N_45706,N_45358,N_45302);
nand U45707 (N_45707,N_45143,N_45434);
or U45708 (N_45708,N_45020,N_45270);
nor U45709 (N_45709,N_45424,N_45377);
nor U45710 (N_45710,N_45430,N_45329);
nor U45711 (N_45711,N_45255,N_45265);
or U45712 (N_45712,N_45309,N_45072);
nor U45713 (N_45713,N_45330,N_45418);
nor U45714 (N_45714,N_45217,N_45379);
nand U45715 (N_45715,N_45350,N_45231);
and U45716 (N_45716,N_45232,N_45398);
or U45717 (N_45717,N_45090,N_45393);
nand U45718 (N_45718,N_45199,N_45496);
or U45719 (N_45719,N_45388,N_45038);
nand U45720 (N_45720,N_45348,N_45321);
and U45721 (N_45721,N_45454,N_45147);
nor U45722 (N_45722,N_45201,N_45071);
nand U45723 (N_45723,N_45468,N_45453);
nor U45724 (N_45724,N_45186,N_45244);
xor U45725 (N_45725,N_45162,N_45029);
and U45726 (N_45726,N_45010,N_45063);
nor U45727 (N_45727,N_45035,N_45360);
or U45728 (N_45728,N_45111,N_45266);
or U45729 (N_45729,N_45165,N_45470);
nor U45730 (N_45730,N_45456,N_45153);
nand U45731 (N_45731,N_45295,N_45243);
or U45732 (N_45732,N_45276,N_45028);
or U45733 (N_45733,N_45356,N_45098);
or U45734 (N_45734,N_45336,N_45209);
or U45735 (N_45735,N_45349,N_45436);
or U45736 (N_45736,N_45025,N_45247);
and U45737 (N_45737,N_45158,N_45170);
nor U45738 (N_45738,N_45228,N_45208);
or U45739 (N_45739,N_45155,N_45296);
or U45740 (N_45740,N_45324,N_45318);
or U45741 (N_45741,N_45280,N_45306);
xnor U45742 (N_45742,N_45126,N_45082);
xnor U45743 (N_45743,N_45460,N_45137);
and U45744 (N_45744,N_45196,N_45142);
nor U45745 (N_45745,N_45101,N_45395);
nand U45746 (N_45746,N_45163,N_45189);
nor U45747 (N_45747,N_45175,N_45074);
xor U45748 (N_45748,N_45259,N_45448);
nand U45749 (N_45749,N_45305,N_45131);
nand U45750 (N_45750,N_45163,N_45372);
nand U45751 (N_45751,N_45207,N_45454);
nand U45752 (N_45752,N_45400,N_45237);
and U45753 (N_45753,N_45307,N_45011);
nand U45754 (N_45754,N_45055,N_45357);
and U45755 (N_45755,N_45333,N_45459);
xnor U45756 (N_45756,N_45303,N_45406);
and U45757 (N_45757,N_45325,N_45040);
or U45758 (N_45758,N_45331,N_45219);
nor U45759 (N_45759,N_45105,N_45250);
nand U45760 (N_45760,N_45084,N_45414);
nor U45761 (N_45761,N_45348,N_45336);
or U45762 (N_45762,N_45321,N_45410);
nand U45763 (N_45763,N_45362,N_45120);
or U45764 (N_45764,N_45187,N_45330);
and U45765 (N_45765,N_45267,N_45312);
nand U45766 (N_45766,N_45296,N_45149);
or U45767 (N_45767,N_45333,N_45277);
nor U45768 (N_45768,N_45310,N_45290);
nand U45769 (N_45769,N_45222,N_45104);
and U45770 (N_45770,N_45146,N_45324);
or U45771 (N_45771,N_45330,N_45037);
and U45772 (N_45772,N_45341,N_45220);
or U45773 (N_45773,N_45460,N_45424);
and U45774 (N_45774,N_45395,N_45116);
nand U45775 (N_45775,N_45196,N_45272);
xnor U45776 (N_45776,N_45374,N_45491);
and U45777 (N_45777,N_45082,N_45241);
nand U45778 (N_45778,N_45206,N_45426);
nor U45779 (N_45779,N_45373,N_45146);
nor U45780 (N_45780,N_45390,N_45382);
nor U45781 (N_45781,N_45488,N_45026);
nor U45782 (N_45782,N_45135,N_45131);
and U45783 (N_45783,N_45457,N_45139);
and U45784 (N_45784,N_45071,N_45483);
or U45785 (N_45785,N_45325,N_45229);
nor U45786 (N_45786,N_45261,N_45178);
or U45787 (N_45787,N_45268,N_45321);
and U45788 (N_45788,N_45146,N_45194);
and U45789 (N_45789,N_45467,N_45231);
and U45790 (N_45790,N_45274,N_45362);
or U45791 (N_45791,N_45155,N_45444);
or U45792 (N_45792,N_45120,N_45330);
nor U45793 (N_45793,N_45001,N_45491);
or U45794 (N_45794,N_45282,N_45016);
or U45795 (N_45795,N_45402,N_45407);
nand U45796 (N_45796,N_45471,N_45060);
and U45797 (N_45797,N_45023,N_45333);
xnor U45798 (N_45798,N_45467,N_45092);
or U45799 (N_45799,N_45098,N_45185);
and U45800 (N_45800,N_45151,N_45036);
nor U45801 (N_45801,N_45066,N_45122);
nand U45802 (N_45802,N_45257,N_45407);
nand U45803 (N_45803,N_45405,N_45282);
nor U45804 (N_45804,N_45165,N_45068);
nor U45805 (N_45805,N_45034,N_45262);
or U45806 (N_45806,N_45150,N_45187);
nor U45807 (N_45807,N_45286,N_45305);
nor U45808 (N_45808,N_45155,N_45215);
and U45809 (N_45809,N_45338,N_45010);
or U45810 (N_45810,N_45262,N_45178);
xor U45811 (N_45811,N_45365,N_45396);
nor U45812 (N_45812,N_45430,N_45437);
and U45813 (N_45813,N_45044,N_45296);
and U45814 (N_45814,N_45076,N_45326);
and U45815 (N_45815,N_45228,N_45466);
nand U45816 (N_45816,N_45401,N_45459);
xor U45817 (N_45817,N_45235,N_45126);
nor U45818 (N_45818,N_45371,N_45203);
or U45819 (N_45819,N_45445,N_45340);
xnor U45820 (N_45820,N_45102,N_45328);
or U45821 (N_45821,N_45378,N_45487);
or U45822 (N_45822,N_45171,N_45003);
and U45823 (N_45823,N_45249,N_45288);
or U45824 (N_45824,N_45335,N_45165);
or U45825 (N_45825,N_45125,N_45137);
and U45826 (N_45826,N_45168,N_45078);
nor U45827 (N_45827,N_45088,N_45446);
nor U45828 (N_45828,N_45457,N_45198);
or U45829 (N_45829,N_45029,N_45179);
nand U45830 (N_45830,N_45136,N_45185);
and U45831 (N_45831,N_45085,N_45206);
nand U45832 (N_45832,N_45060,N_45486);
nand U45833 (N_45833,N_45346,N_45461);
nor U45834 (N_45834,N_45235,N_45066);
nand U45835 (N_45835,N_45229,N_45395);
or U45836 (N_45836,N_45244,N_45142);
or U45837 (N_45837,N_45085,N_45125);
nor U45838 (N_45838,N_45368,N_45176);
or U45839 (N_45839,N_45042,N_45312);
nor U45840 (N_45840,N_45212,N_45274);
xnor U45841 (N_45841,N_45240,N_45337);
nor U45842 (N_45842,N_45138,N_45452);
nor U45843 (N_45843,N_45086,N_45120);
or U45844 (N_45844,N_45321,N_45312);
and U45845 (N_45845,N_45323,N_45146);
nor U45846 (N_45846,N_45143,N_45124);
xnor U45847 (N_45847,N_45162,N_45327);
nor U45848 (N_45848,N_45342,N_45163);
xor U45849 (N_45849,N_45336,N_45111);
nand U45850 (N_45850,N_45263,N_45430);
and U45851 (N_45851,N_45227,N_45493);
and U45852 (N_45852,N_45235,N_45308);
nor U45853 (N_45853,N_45393,N_45243);
or U45854 (N_45854,N_45350,N_45018);
nand U45855 (N_45855,N_45066,N_45216);
nand U45856 (N_45856,N_45293,N_45497);
and U45857 (N_45857,N_45326,N_45333);
and U45858 (N_45858,N_45083,N_45084);
nand U45859 (N_45859,N_45396,N_45213);
and U45860 (N_45860,N_45119,N_45495);
or U45861 (N_45861,N_45015,N_45429);
or U45862 (N_45862,N_45322,N_45017);
and U45863 (N_45863,N_45214,N_45468);
nand U45864 (N_45864,N_45465,N_45109);
nor U45865 (N_45865,N_45245,N_45294);
or U45866 (N_45866,N_45147,N_45026);
xnor U45867 (N_45867,N_45147,N_45422);
and U45868 (N_45868,N_45311,N_45453);
or U45869 (N_45869,N_45255,N_45396);
xor U45870 (N_45870,N_45191,N_45453);
and U45871 (N_45871,N_45460,N_45016);
or U45872 (N_45872,N_45200,N_45122);
and U45873 (N_45873,N_45225,N_45253);
nand U45874 (N_45874,N_45345,N_45210);
nor U45875 (N_45875,N_45258,N_45390);
nand U45876 (N_45876,N_45358,N_45258);
nor U45877 (N_45877,N_45281,N_45060);
nand U45878 (N_45878,N_45027,N_45078);
nand U45879 (N_45879,N_45283,N_45291);
or U45880 (N_45880,N_45108,N_45014);
and U45881 (N_45881,N_45043,N_45063);
nand U45882 (N_45882,N_45140,N_45206);
nor U45883 (N_45883,N_45330,N_45102);
and U45884 (N_45884,N_45277,N_45287);
and U45885 (N_45885,N_45363,N_45197);
or U45886 (N_45886,N_45466,N_45108);
and U45887 (N_45887,N_45130,N_45397);
and U45888 (N_45888,N_45246,N_45336);
or U45889 (N_45889,N_45098,N_45059);
or U45890 (N_45890,N_45275,N_45488);
and U45891 (N_45891,N_45323,N_45386);
and U45892 (N_45892,N_45304,N_45255);
nand U45893 (N_45893,N_45318,N_45052);
xor U45894 (N_45894,N_45359,N_45284);
or U45895 (N_45895,N_45240,N_45248);
or U45896 (N_45896,N_45306,N_45160);
nand U45897 (N_45897,N_45174,N_45248);
and U45898 (N_45898,N_45199,N_45461);
nor U45899 (N_45899,N_45254,N_45203);
nor U45900 (N_45900,N_45361,N_45231);
nand U45901 (N_45901,N_45472,N_45087);
or U45902 (N_45902,N_45258,N_45479);
nor U45903 (N_45903,N_45354,N_45015);
nor U45904 (N_45904,N_45320,N_45227);
or U45905 (N_45905,N_45301,N_45375);
and U45906 (N_45906,N_45437,N_45429);
xor U45907 (N_45907,N_45232,N_45219);
and U45908 (N_45908,N_45049,N_45409);
and U45909 (N_45909,N_45467,N_45321);
nor U45910 (N_45910,N_45383,N_45218);
or U45911 (N_45911,N_45291,N_45049);
or U45912 (N_45912,N_45200,N_45226);
and U45913 (N_45913,N_45299,N_45181);
nor U45914 (N_45914,N_45193,N_45039);
and U45915 (N_45915,N_45483,N_45111);
and U45916 (N_45916,N_45099,N_45276);
nor U45917 (N_45917,N_45262,N_45387);
or U45918 (N_45918,N_45117,N_45385);
xnor U45919 (N_45919,N_45011,N_45401);
nand U45920 (N_45920,N_45214,N_45254);
nand U45921 (N_45921,N_45338,N_45370);
and U45922 (N_45922,N_45419,N_45446);
and U45923 (N_45923,N_45236,N_45425);
or U45924 (N_45924,N_45410,N_45203);
nand U45925 (N_45925,N_45351,N_45286);
nand U45926 (N_45926,N_45115,N_45183);
nand U45927 (N_45927,N_45191,N_45161);
or U45928 (N_45928,N_45167,N_45379);
nand U45929 (N_45929,N_45209,N_45474);
or U45930 (N_45930,N_45033,N_45227);
and U45931 (N_45931,N_45111,N_45205);
and U45932 (N_45932,N_45077,N_45113);
or U45933 (N_45933,N_45461,N_45359);
and U45934 (N_45934,N_45074,N_45430);
xnor U45935 (N_45935,N_45262,N_45282);
nand U45936 (N_45936,N_45043,N_45251);
xnor U45937 (N_45937,N_45128,N_45034);
and U45938 (N_45938,N_45277,N_45145);
nand U45939 (N_45939,N_45186,N_45203);
and U45940 (N_45940,N_45306,N_45105);
nand U45941 (N_45941,N_45464,N_45305);
or U45942 (N_45942,N_45335,N_45451);
and U45943 (N_45943,N_45451,N_45234);
xor U45944 (N_45944,N_45423,N_45286);
nor U45945 (N_45945,N_45162,N_45473);
nand U45946 (N_45946,N_45171,N_45205);
nand U45947 (N_45947,N_45341,N_45231);
nor U45948 (N_45948,N_45041,N_45268);
nor U45949 (N_45949,N_45353,N_45276);
xnor U45950 (N_45950,N_45098,N_45417);
nor U45951 (N_45951,N_45353,N_45206);
and U45952 (N_45952,N_45370,N_45297);
nor U45953 (N_45953,N_45360,N_45380);
nor U45954 (N_45954,N_45157,N_45049);
xor U45955 (N_45955,N_45331,N_45431);
nor U45956 (N_45956,N_45227,N_45114);
nand U45957 (N_45957,N_45009,N_45330);
nor U45958 (N_45958,N_45181,N_45308);
or U45959 (N_45959,N_45134,N_45234);
nor U45960 (N_45960,N_45261,N_45478);
and U45961 (N_45961,N_45492,N_45353);
or U45962 (N_45962,N_45488,N_45471);
xor U45963 (N_45963,N_45103,N_45260);
and U45964 (N_45964,N_45171,N_45261);
or U45965 (N_45965,N_45115,N_45391);
nand U45966 (N_45966,N_45209,N_45376);
nor U45967 (N_45967,N_45422,N_45308);
or U45968 (N_45968,N_45133,N_45366);
or U45969 (N_45969,N_45084,N_45297);
or U45970 (N_45970,N_45143,N_45349);
or U45971 (N_45971,N_45340,N_45079);
and U45972 (N_45972,N_45436,N_45137);
nand U45973 (N_45973,N_45005,N_45070);
and U45974 (N_45974,N_45061,N_45308);
nor U45975 (N_45975,N_45475,N_45304);
or U45976 (N_45976,N_45281,N_45460);
nor U45977 (N_45977,N_45130,N_45396);
nand U45978 (N_45978,N_45196,N_45269);
and U45979 (N_45979,N_45228,N_45094);
and U45980 (N_45980,N_45169,N_45175);
xor U45981 (N_45981,N_45134,N_45133);
and U45982 (N_45982,N_45047,N_45245);
and U45983 (N_45983,N_45271,N_45084);
nor U45984 (N_45984,N_45151,N_45169);
or U45985 (N_45985,N_45107,N_45231);
nand U45986 (N_45986,N_45233,N_45465);
nand U45987 (N_45987,N_45056,N_45437);
xor U45988 (N_45988,N_45139,N_45037);
nand U45989 (N_45989,N_45316,N_45422);
and U45990 (N_45990,N_45390,N_45462);
and U45991 (N_45991,N_45462,N_45020);
or U45992 (N_45992,N_45205,N_45086);
nand U45993 (N_45993,N_45009,N_45241);
and U45994 (N_45994,N_45051,N_45182);
or U45995 (N_45995,N_45136,N_45355);
or U45996 (N_45996,N_45320,N_45299);
and U45997 (N_45997,N_45161,N_45159);
or U45998 (N_45998,N_45000,N_45487);
or U45999 (N_45999,N_45041,N_45433);
or U46000 (N_46000,N_45932,N_45926);
nor U46001 (N_46001,N_45706,N_45740);
or U46002 (N_46002,N_45798,N_45900);
or U46003 (N_46003,N_45690,N_45726);
nand U46004 (N_46004,N_45974,N_45684);
or U46005 (N_46005,N_45611,N_45579);
and U46006 (N_46006,N_45561,N_45841);
nand U46007 (N_46007,N_45592,N_45959);
nand U46008 (N_46008,N_45615,N_45644);
nor U46009 (N_46009,N_45714,N_45998);
nand U46010 (N_46010,N_45997,N_45890);
or U46011 (N_46011,N_45526,N_45624);
nand U46012 (N_46012,N_45949,N_45565);
or U46013 (N_46013,N_45739,N_45816);
and U46014 (N_46014,N_45529,N_45756);
and U46015 (N_46015,N_45605,N_45977);
and U46016 (N_46016,N_45769,N_45961);
or U46017 (N_46017,N_45658,N_45770);
nand U46018 (N_46018,N_45801,N_45757);
xor U46019 (N_46019,N_45896,N_45534);
and U46020 (N_46020,N_45908,N_45783);
nor U46021 (N_46021,N_45876,N_45987);
or U46022 (N_46022,N_45598,N_45917);
nor U46023 (N_46023,N_45507,N_45652);
and U46024 (N_46024,N_45732,N_45636);
nand U46025 (N_46025,N_45805,N_45952);
or U46026 (N_46026,N_45635,N_45898);
nor U46027 (N_46027,N_45523,N_45905);
or U46028 (N_46028,N_45901,N_45887);
and U46029 (N_46029,N_45707,N_45849);
nor U46030 (N_46030,N_45613,N_45790);
and U46031 (N_46031,N_45914,N_45559);
or U46032 (N_46032,N_45692,N_45623);
or U46033 (N_46033,N_45878,N_45948);
and U46034 (N_46034,N_45577,N_45510);
or U46035 (N_46035,N_45587,N_45681);
and U46036 (N_46036,N_45865,N_45985);
and U46037 (N_46037,N_45567,N_45689);
and U46038 (N_46038,N_45612,N_45674);
or U46039 (N_46039,N_45923,N_45662);
and U46040 (N_46040,N_45767,N_45633);
or U46041 (N_46041,N_45618,N_45826);
nand U46042 (N_46042,N_45676,N_45936);
nor U46043 (N_46043,N_45825,N_45820);
nand U46044 (N_46044,N_45793,N_45713);
and U46045 (N_46045,N_45924,N_45667);
nand U46046 (N_46046,N_45875,N_45728);
nand U46047 (N_46047,N_45734,N_45906);
nand U46048 (N_46048,N_45916,N_45504);
nand U46049 (N_46049,N_45607,N_45913);
nand U46050 (N_46050,N_45555,N_45775);
or U46051 (N_46051,N_45902,N_45649);
or U46052 (N_46052,N_45996,N_45861);
nor U46053 (N_46053,N_45910,N_45854);
or U46054 (N_46054,N_45538,N_45947);
nand U46055 (N_46055,N_45547,N_45549);
nor U46056 (N_46056,N_45711,N_45646);
or U46057 (N_46057,N_45956,N_45893);
xnor U46058 (N_46058,N_45809,N_45620);
nor U46059 (N_46059,N_45621,N_45761);
nand U46060 (N_46060,N_45682,N_45863);
xor U46061 (N_46061,N_45606,N_45812);
nor U46062 (N_46062,N_45528,N_45999);
nand U46063 (N_46063,N_45963,N_45846);
or U46064 (N_46064,N_45982,N_45683);
and U46065 (N_46065,N_45840,N_45870);
nand U46066 (N_46066,N_45837,N_45797);
and U46067 (N_46067,N_45639,N_45753);
nand U46068 (N_46068,N_45604,N_45637);
or U46069 (N_46069,N_45558,N_45920);
or U46070 (N_46070,N_45842,N_45929);
xnor U46071 (N_46071,N_45693,N_45970);
and U46072 (N_46072,N_45839,N_45562);
xor U46073 (N_46073,N_45694,N_45532);
nor U46074 (N_46074,N_45838,N_45943);
or U46075 (N_46075,N_45672,N_45641);
nand U46076 (N_46076,N_45748,N_45852);
nor U46077 (N_46077,N_45551,N_45645);
and U46078 (N_46078,N_45880,N_45502);
nand U46079 (N_46079,N_45819,N_45758);
or U46080 (N_46080,N_45525,N_45979);
xnor U46081 (N_46081,N_45834,N_45955);
xor U46082 (N_46082,N_45744,N_45871);
nor U46083 (N_46083,N_45516,N_45832);
nand U46084 (N_46084,N_45669,N_45655);
nand U46085 (N_46085,N_45716,N_45953);
nand U46086 (N_46086,N_45990,N_45666);
and U46087 (N_46087,N_45600,N_45543);
nor U46088 (N_46088,N_45518,N_45981);
and U46089 (N_46089,N_45991,N_45980);
or U46090 (N_46090,N_45904,N_45671);
and U46091 (N_46091,N_45759,N_45527);
nor U46092 (N_46092,N_45568,N_45622);
nor U46093 (N_46093,N_45608,N_45712);
nand U46094 (N_46094,N_45780,N_45754);
and U46095 (N_46095,N_45934,N_45601);
and U46096 (N_46096,N_45563,N_45836);
and U46097 (N_46097,N_45540,N_45822);
and U46098 (N_46098,N_45668,N_45976);
nand U46099 (N_46099,N_45988,N_45627);
or U46100 (N_46100,N_45511,N_45574);
nand U46101 (N_46101,N_45519,N_45699);
or U46102 (N_46102,N_45771,N_45735);
and U46103 (N_46103,N_45994,N_45588);
xor U46104 (N_46104,N_45553,N_45750);
or U46105 (N_46105,N_45781,N_45686);
nor U46106 (N_46106,N_45866,N_45995);
or U46107 (N_46107,N_45844,N_45892);
nand U46108 (N_46108,N_45556,N_45873);
and U46109 (N_46109,N_45807,N_45872);
nor U46110 (N_46110,N_45856,N_45782);
nor U46111 (N_46111,N_45815,N_45992);
or U46112 (N_46112,N_45894,N_45792);
nor U46113 (N_46113,N_45772,N_45760);
and U46114 (N_46114,N_45550,N_45591);
or U46115 (N_46115,N_45745,N_45680);
or U46116 (N_46116,N_45791,N_45777);
or U46117 (N_46117,N_45886,N_45742);
nor U46118 (N_46118,N_45884,N_45720);
or U46119 (N_46119,N_45544,N_45847);
xor U46120 (N_46120,N_45656,N_45575);
nand U46121 (N_46121,N_45922,N_45500);
xnor U46122 (N_46122,N_45899,N_45560);
or U46123 (N_46123,N_45803,N_45944);
and U46124 (N_46124,N_45535,N_45983);
and U46125 (N_46125,N_45594,N_45640);
and U46126 (N_46126,N_45817,N_45533);
nor U46127 (N_46127,N_45883,N_45648);
nand U46128 (N_46128,N_45675,N_45814);
and U46129 (N_46129,N_45546,N_45521);
or U46130 (N_46130,N_45705,N_45531);
or U46131 (N_46131,N_45524,N_45536);
and U46132 (N_46132,N_45704,N_45984);
nand U46133 (N_46133,N_45653,N_45715);
or U46134 (N_46134,N_45619,N_45566);
xor U46135 (N_46135,N_45741,N_45573);
or U46136 (N_46136,N_45804,N_45788);
and U46137 (N_46137,N_45897,N_45581);
and U46138 (N_46138,N_45643,N_45664);
xor U46139 (N_46139,N_45599,N_45864);
xnor U46140 (N_46140,N_45879,N_45634);
and U46141 (N_46141,N_45794,N_45743);
or U46142 (N_46142,N_45628,N_45749);
or U46143 (N_46143,N_45554,N_45891);
nor U46144 (N_46144,N_45821,N_45729);
nand U46145 (N_46145,N_45935,N_45731);
and U46146 (N_46146,N_45746,N_45933);
nand U46147 (N_46147,N_45765,N_45971);
nor U46148 (N_46148,N_45964,N_45862);
and U46149 (N_46149,N_45708,N_45501);
and U46150 (N_46150,N_45751,N_45576);
and U46151 (N_46151,N_45522,N_45818);
and U46152 (N_46152,N_45539,N_45673);
or U46153 (N_46153,N_45965,N_45806);
or U46154 (N_46154,N_45590,N_45571);
and U46155 (N_46155,N_45657,N_45702);
nor U46156 (N_46156,N_45966,N_45659);
xnor U46157 (N_46157,N_45882,N_45718);
and U46158 (N_46158,N_45677,N_45786);
nor U46159 (N_46159,N_45958,N_45853);
or U46160 (N_46160,N_45651,N_45631);
xnor U46161 (N_46161,N_45730,N_45614);
nand U46162 (N_46162,N_45650,N_45831);
and U46163 (N_46163,N_45810,N_45685);
and U46164 (N_46164,N_45927,N_45530);
nand U46165 (N_46165,N_45795,N_45572);
and U46166 (N_46166,N_45695,N_45957);
or U46167 (N_46167,N_45629,N_45603);
or U46168 (N_46168,N_45787,N_45975);
nand U46169 (N_46169,N_45828,N_45903);
or U46170 (N_46170,N_45915,N_45687);
nor U46171 (N_46171,N_45569,N_45665);
or U46172 (N_46172,N_45578,N_45808);
and U46173 (N_46173,N_45638,N_45691);
or U46174 (N_46174,N_45833,N_45800);
and U46175 (N_46175,N_45940,N_45867);
xnor U46176 (N_46176,N_45513,N_45595);
and U46177 (N_46177,N_45951,N_45796);
xnor U46178 (N_46178,N_45874,N_45950);
nand U46179 (N_46179,N_45938,N_45789);
nor U46180 (N_46180,N_45725,N_45850);
or U46181 (N_46181,N_45552,N_45610);
nand U46182 (N_46182,N_45919,N_45946);
xnor U46183 (N_46183,N_45857,N_45960);
and U46184 (N_46184,N_45654,N_45722);
nand U46185 (N_46185,N_45670,N_45973);
nor U46186 (N_46186,N_45733,N_45738);
and U46187 (N_46187,N_45907,N_45506);
xnor U46188 (N_46188,N_45703,N_45597);
or U46189 (N_46189,N_45773,N_45942);
and U46190 (N_46190,N_45724,N_45514);
nor U46191 (N_46191,N_45700,N_45663);
nand U46192 (N_46192,N_45537,N_45586);
nor U46193 (N_46193,N_45678,N_45564);
nand U46194 (N_46194,N_45911,N_45642);
and U46195 (N_46195,N_45823,N_45617);
and U46196 (N_46196,N_45784,N_45928);
or U46197 (N_46197,N_45517,N_45503);
nand U46198 (N_46198,N_45858,N_45709);
nand U46199 (N_46199,N_45895,N_45557);
nor U46200 (N_46200,N_45602,N_45593);
nor U46201 (N_46201,N_45545,N_45869);
nand U46202 (N_46202,N_45939,N_45515);
nor U46203 (N_46203,N_45993,N_45931);
xnor U46204 (N_46204,N_45888,N_45679);
nand U46205 (N_46205,N_45855,N_45989);
nand U46206 (N_46206,N_45830,N_45727);
or U46207 (N_46207,N_45868,N_45968);
nor U46208 (N_46208,N_45778,N_45717);
nand U46209 (N_46209,N_45583,N_45986);
and U46210 (N_46210,N_45508,N_45736);
and U46211 (N_46211,N_45710,N_45766);
nand U46212 (N_46212,N_45859,N_45877);
nor U46213 (N_46213,N_45918,N_45582);
and U46214 (N_46214,N_45723,N_45829);
or U46215 (N_46215,N_45921,N_45937);
nand U46216 (N_46216,N_45632,N_45776);
and U46217 (N_46217,N_45851,N_45799);
nor U46218 (N_46218,N_45625,N_45762);
nor U46219 (N_46219,N_45811,N_45813);
xor U46220 (N_46220,N_45747,N_45737);
nor U46221 (N_46221,N_45764,N_45945);
and U46222 (N_46222,N_45752,N_45616);
nand U46223 (N_46223,N_45824,N_45580);
nor U46224 (N_46224,N_45962,N_45630);
nand U46225 (N_46225,N_45848,N_45978);
and U46226 (N_46226,N_45688,N_45696);
xnor U46227 (N_46227,N_45570,N_45802);
nand U46228 (N_46228,N_45925,N_45542);
xnor U46229 (N_46229,N_45779,N_45585);
xnor U46230 (N_46230,N_45596,N_45941);
or U46231 (N_46231,N_45860,N_45827);
nor U46232 (N_46232,N_45889,N_45721);
nand U46233 (N_46233,N_45698,N_45505);
xnor U46234 (N_46234,N_45835,N_45520);
xnor U46235 (N_46235,N_45701,N_45763);
and U46236 (N_46236,N_45885,N_45719);
nand U46237 (N_46237,N_45881,N_45509);
nor U46238 (N_46238,N_45755,N_45512);
nand U46239 (N_46239,N_45647,N_45541);
xnor U46240 (N_46240,N_45909,N_45660);
xnor U46241 (N_46241,N_45609,N_45584);
and U46242 (N_46242,N_45845,N_45626);
nand U46243 (N_46243,N_45843,N_45954);
nand U46244 (N_46244,N_45785,N_45774);
xnor U46245 (N_46245,N_45661,N_45967);
nor U46246 (N_46246,N_45930,N_45912);
nor U46247 (N_46247,N_45548,N_45969);
or U46248 (N_46248,N_45768,N_45589);
or U46249 (N_46249,N_45697,N_45972);
nand U46250 (N_46250,N_45714,N_45502);
xor U46251 (N_46251,N_45519,N_45807);
and U46252 (N_46252,N_45544,N_45903);
xor U46253 (N_46253,N_45806,N_45551);
nand U46254 (N_46254,N_45917,N_45977);
nor U46255 (N_46255,N_45879,N_45627);
nor U46256 (N_46256,N_45581,N_45902);
or U46257 (N_46257,N_45943,N_45967);
xnor U46258 (N_46258,N_45527,N_45920);
nor U46259 (N_46259,N_45895,N_45532);
nand U46260 (N_46260,N_45610,N_45882);
and U46261 (N_46261,N_45880,N_45655);
xor U46262 (N_46262,N_45602,N_45905);
nand U46263 (N_46263,N_45559,N_45998);
nor U46264 (N_46264,N_45557,N_45582);
nor U46265 (N_46265,N_45639,N_45812);
or U46266 (N_46266,N_45825,N_45640);
or U46267 (N_46267,N_45625,N_45523);
nand U46268 (N_46268,N_45511,N_45993);
or U46269 (N_46269,N_45723,N_45942);
nor U46270 (N_46270,N_45553,N_45986);
and U46271 (N_46271,N_45978,N_45640);
and U46272 (N_46272,N_45766,N_45508);
nand U46273 (N_46273,N_45732,N_45657);
nand U46274 (N_46274,N_45986,N_45607);
nor U46275 (N_46275,N_45605,N_45694);
xor U46276 (N_46276,N_45751,N_45520);
nor U46277 (N_46277,N_45643,N_45687);
nand U46278 (N_46278,N_45615,N_45960);
nand U46279 (N_46279,N_45915,N_45816);
nand U46280 (N_46280,N_45699,N_45744);
or U46281 (N_46281,N_45612,N_45705);
and U46282 (N_46282,N_45700,N_45674);
nand U46283 (N_46283,N_45915,N_45543);
xnor U46284 (N_46284,N_45777,N_45701);
or U46285 (N_46285,N_45510,N_45603);
and U46286 (N_46286,N_45883,N_45850);
or U46287 (N_46287,N_45574,N_45502);
or U46288 (N_46288,N_45753,N_45709);
and U46289 (N_46289,N_45809,N_45664);
or U46290 (N_46290,N_45575,N_45856);
nand U46291 (N_46291,N_45576,N_45801);
nor U46292 (N_46292,N_45998,N_45607);
nand U46293 (N_46293,N_45864,N_45878);
xor U46294 (N_46294,N_45721,N_45874);
or U46295 (N_46295,N_45634,N_45887);
and U46296 (N_46296,N_45746,N_45822);
nor U46297 (N_46297,N_45832,N_45827);
and U46298 (N_46298,N_45697,N_45632);
and U46299 (N_46299,N_45527,N_45664);
nor U46300 (N_46300,N_45828,N_45906);
and U46301 (N_46301,N_45894,N_45515);
nand U46302 (N_46302,N_45754,N_45638);
nand U46303 (N_46303,N_45919,N_45938);
nand U46304 (N_46304,N_45659,N_45691);
nand U46305 (N_46305,N_45762,N_45891);
nand U46306 (N_46306,N_45989,N_45996);
and U46307 (N_46307,N_45637,N_45841);
and U46308 (N_46308,N_45681,N_45913);
nand U46309 (N_46309,N_45957,N_45740);
nand U46310 (N_46310,N_45618,N_45598);
nor U46311 (N_46311,N_45548,N_45875);
xnor U46312 (N_46312,N_45692,N_45745);
nand U46313 (N_46313,N_45713,N_45768);
xor U46314 (N_46314,N_45525,N_45916);
or U46315 (N_46315,N_45711,N_45523);
or U46316 (N_46316,N_45635,N_45510);
or U46317 (N_46317,N_45523,N_45648);
nor U46318 (N_46318,N_45766,N_45500);
and U46319 (N_46319,N_45554,N_45897);
and U46320 (N_46320,N_45747,N_45790);
and U46321 (N_46321,N_45586,N_45954);
and U46322 (N_46322,N_45717,N_45621);
nor U46323 (N_46323,N_45745,N_45644);
nor U46324 (N_46324,N_45985,N_45824);
or U46325 (N_46325,N_45720,N_45928);
or U46326 (N_46326,N_45804,N_45769);
nand U46327 (N_46327,N_45542,N_45689);
nand U46328 (N_46328,N_45856,N_45744);
or U46329 (N_46329,N_45879,N_45687);
and U46330 (N_46330,N_45590,N_45880);
or U46331 (N_46331,N_45881,N_45662);
or U46332 (N_46332,N_45834,N_45781);
nor U46333 (N_46333,N_45866,N_45519);
and U46334 (N_46334,N_45504,N_45833);
nand U46335 (N_46335,N_45653,N_45865);
nor U46336 (N_46336,N_45796,N_45974);
or U46337 (N_46337,N_45969,N_45500);
or U46338 (N_46338,N_45858,N_45698);
and U46339 (N_46339,N_45601,N_45853);
and U46340 (N_46340,N_45647,N_45784);
or U46341 (N_46341,N_45581,N_45950);
and U46342 (N_46342,N_45730,N_45928);
nand U46343 (N_46343,N_45567,N_45557);
and U46344 (N_46344,N_45995,N_45786);
or U46345 (N_46345,N_45571,N_45531);
and U46346 (N_46346,N_45608,N_45864);
xor U46347 (N_46347,N_45654,N_45810);
or U46348 (N_46348,N_45994,N_45534);
nor U46349 (N_46349,N_45937,N_45933);
and U46350 (N_46350,N_45823,N_45579);
or U46351 (N_46351,N_45796,N_45590);
nor U46352 (N_46352,N_45561,N_45896);
and U46353 (N_46353,N_45814,N_45964);
nand U46354 (N_46354,N_45764,N_45994);
or U46355 (N_46355,N_45629,N_45669);
and U46356 (N_46356,N_45984,N_45698);
nor U46357 (N_46357,N_45841,N_45972);
nand U46358 (N_46358,N_45860,N_45948);
or U46359 (N_46359,N_45920,N_45706);
and U46360 (N_46360,N_45546,N_45924);
nor U46361 (N_46361,N_45617,N_45698);
nor U46362 (N_46362,N_45880,N_45820);
nand U46363 (N_46363,N_45727,N_45594);
or U46364 (N_46364,N_45515,N_45686);
nor U46365 (N_46365,N_45860,N_45779);
and U46366 (N_46366,N_45639,N_45670);
or U46367 (N_46367,N_45736,N_45815);
or U46368 (N_46368,N_45705,N_45920);
nor U46369 (N_46369,N_45898,N_45581);
nand U46370 (N_46370,N_45826,N_45781);
and U46371 (N_46371,N_45668,N_45544);
and U46372 (N_46372,N_45862,N_45998);
or U46373 (N_46373,N_45529,N_45578);
nor U46374 (N_46374,N_45637,N_45677);
nand U46375 (N_46375,N_45986,N_45887);
nand U46376 (N_46376,N_45984,N_45703);
nor U46377 (N_46377,N_45734,N_45634);
nor U46378 (N_46378,N_45763,N_45971);
xnor U46379 (N_46379,N_45849,N_45549);
nor U46380 (N_46380,N_45585,N_45888);
nor U46381 (N_46381,N_45639,N_45928);
nand U46382 (N_46382,N_45700,N_45841);
nor U46383 (N_46383,N_45768,N_45605);
and U46384 (N_46384,N_45791,N_45828);
nor U46385 (N_46385,N_45646,N_45602);
nor U46386 (N_46386,N_45920,N_45543);
or U46387 (N_46387,N_45656,N_45811);
or U46388 (N_46388,N_45693,N_45926);
nor U46389 (N_46389,N_45777,N_45717);
nor U46390 (N_46390,N_45982,N_45872);
nor U46391 (N_46391,N_45517,N_45904);
and U46392 (N_46392,N_45964,N_45823);
nand U46393 (N_46393,N_45899,N_45934);
nor U46394 (N_46394,N_45619,N_45650);
nand U46395 (N_46395,N_45882,N_45756);
and U46396 (N_46396,N_45876,N_45862);
and U46397 (N_46397,N_45609,N_45612);
or U46398 (N_46398,N_45993,N_45534);
and U46399 (N_46399,N_45658,N_45797);
nand U46400 (N_46400,N_45949,N_45684);
and U46401 (N_46401,N_45762,N_45868);
nor U46402 (N_46402,N_45566,N_45578);
or U46403 (N_46403,N_45583,N_45786);
and U46404 (N_46404,N_45862,N_45694);
or U46405 (N_46405,N_45938,N_45677);
or U46406 (N_46406,N_45964,N_45729);
nor U46407 (N_46407,N_45571,N_45880);
nor U46408 (N_46408,N_45766,N_45571);
or U46409 (N_46409,N_45899,N_45619);
nor U46410 (N_46410,N_45907,N_45548);
nand U46411 (N_46411,N_45748,N_45701);
nor U46412 (N_46412,N_45735,N_45561);
or U46413 (N_46413,N_45706,N_45945);
and U46414 (N_46414,N_45778,N_45607);
nand U46415 (N_46415,N_45802,N_45607);
and U46416 (N_46416,N_45566,N_45929);
or U46417 (N_46417,N_45529,N_45775);
xor U46418 (N_46418,N_45565,N_45881);
and U46419 (N_46419,N_45871,N_45831);
or U46420 (N_46420,N_45922,N_45771);
nand U46421 (N_46421,N_45519,N_45785);
nand U46422 (N_46422,N_45575,N_45845);
and U46423 (N_46423,N_45681,N_45837);
nor U46424 (N_46424,N_45692,N_45836);
or U46425 (N_46425,N_45857,N_45854);
nor U46426 (N_46426,N_45566,N_45953);
nand U46427 (N_46427,N_45952,N_45540);
and U46428 (N_46428,N_45786,N_45681);
or U46429 (N_46429,N_45983,N_45940);
or U46430 (N_46430,N_45950,N_45785);
or U46431 (N_46431,N_45526,N_45556);
and U46432 (N_46432,N_45726,N_45530);
or U46433 (N_46433,N_45558,N_45785);
or U46434 (N_46434,N_45947,N_45558);
and U46435 (N_46435,N_45924,N_45506);
or U46436 (N_46436,N_45808,N_45802);
or U46437 (N_46437,N_45543,N_45722);
and U46438 (N_46438,N_45649,N_45845);
and U46439 (N_46439,N_45879,N_45674);
nand U46440 (N_46440,N_45993,N_45942);
or U46441 (N_46441,N_45833,N_45587);
and U46442 (N_46442,N_45807,N_45729);
and U46443 (N_46443,N_45810,N_45604);
or U46444 (N_46444,N_45678,N_45874);
or U46445 (N_46445,N_45743,N_45834);
nand U46446 (N_46446,N_45521,N_45530);
xor U46447 (N_46447,N_45855,N_45634);
nand U46448 (N_46448,N_45590,N_45797);
xor U46449 (N_46449,N_45990,N_45641);
or U46450 (N_46450,N_45960,N_45803);
nor U46451 (N_46451,N_45718,N_45886);
or U46452 (N_46452,N_45788,N_45572);
xor U46453 (N_46453,N_45824,N_45516);
nand U46454 (N_46454,N_45661,N_45503);
nor U46455 (N_46455,N_45514,N_45510);
nand U46456 (N_46456,N_45891,N_45546);
or U46457 (N_46457,N_45781,N_45822);
nor U46458 (N_46458,N_45558,N_45571);
nand U46459 (N_46459,N_45669,N_45829);
nand U46460 (N_46460,N_45505,N_45941);
xor U46461 (N_46461,N_45753,N_45926);
or U46462 (N_46462,N_45750,N_45650);
or U46463 (N_46463,N_45945,N_45791);
nor U46464 (N_46464,N_45702,N_45531);
nand U46465 (N_46465,N_45900,N_45754);
nor U46466 (N_46466,N_45882,N_45568);
or U46467 (N_46467,N_45620,N_45610);
and U46468 (N_46468,N_45871,N_45570);
and U46469 (N_46469,N_45636,N_45553);
and U46470 (N_46470,N_45852,N_45937);
or U46471 (N_46471,N_45562,N_45820);
and U46472 (N_46472,N_45936,N_45848);
nor U46473 (N_46473,N_45889,N_45528);
nor U46474 (N_46474,N_45949,N_45599);
and U46475 (N_46475,N_45915,N_45899);
nor U46476 (N_46476,N_45831,N_45607);
nor U46477 (N_46477,N_45779,N_45757);
xor U46478 (N_46478,N_45644,N_45680);
and U46479 (N_46479,N_45613,N_45838);
nor U46480 (N_46480,N_45999,N_45501);
and U46481 (N_46481,N_45806,N_45577);
nor U46482 (N_46482,N_45919,N_45696);
or U46483 (N_46483,N_45807,N_45797);
or U46484 (N_46484,N_45585,N_45852);
nor U46485 (N_46485,N_45835,N_45822);
or U46486 (N_46486,N_45893,N_45922);
xor U46487 (N_46487,N_45501,N_45723);
and U46488 (N_46488,N_45503,N_45559);
xnor U46489 (N_46489,N_45547,N_45618);
or U46490 (N_46490,N_45875,N_45767);
nor U46491 (N_46491,N_45817,N_45828);
or U46492 (N_46492,N_45681,N_45583);
and U46493 (N_46493,N_45788,N_45784);
nand U46494 (N_46494,N_45667,N_45764);
nor U46495 (N_46495,N_45739,N_45677);
nor U46496 (N_46496,N_45799,N_45757);
nor U46497 (N_46497,N_45616,N_45739);
or U46498 (N_46498,N_45875,N_45785);
and U46499 (N_46499,N_45639,N_45960);
and U46500 (N_46500,N_46035,N_46173);
nand U46501 (N_46501,N_46434,N_46214);
nor U46502 (N_46502,N_46161,N_46144);
and U46503 (N_46503,N_46051,N_46108);
and U46504 (N_46504,N_46203,N_46458);
and U46505 (N_46505,N_46427,N_46360);
nand U46506 (N_46506,N_46482,N_46474);
nor U46507 (N_46507,N_46054,N_46251);
or U46508 (N_46508,N_46055,N_46181);
xor U46509 (N_46509,N_46175,N_46351);
nor U46510 (N_46510,N_46358,N_46262);
nand U46511 (N_46511,N_46118,N_46001);
and U46512 (N_46512,N_46237,N_46371);
and U46513 (N_46513,N_46249,N_46209);
xnor U46514 (N_46514,N_46211,N_46460);
and U46515 (N_46515,N_46115,N_46164);
nand U46516 (N_46516,N_46309,N_46299);
and U46517 (N_46517,N_46403,N_46199);
nor U46518 (N_46518,N_46480,N_46014);
nor U46519 (N_46519,N_46461,N_46133);
or U46520 (N_46520,N_46433,N_46192);
nor U46521 (N_46521,N_46085,N_46442);
nand U46522 (N_46522,N_46229,N_46392);
xnor U46523 (N_46523,N_46241,N_46132);
nor U46524 (N_46524,N_46182,N_46149);
xnor U46525 (N_46525,N_46188,N_46408);
nand U46526 (N_46526,N_46471,N_46201);
or U46527 (N_46527,N_46011,N_46096);
xor U46528 (N_46528,N_46267,N_46289);
or U46529 (N_46529,N_46288,N_46074);
xor U46530 (N_46530,N_46194,N_46105);
or U46531 (N_46531,N_46219,N_46165);
xor U46532 (N_46532,N_46272,N_46270);
nor U46533 (N_46533,N_46489,N_46031);
nor U46534 (N_46534,N_46316,N_46143);
nand U46535 (N_46535,N_46002,N_46378);
nor U46536 (N_46536,N_46359,N_46236);
and U46537 (N_46537,N_46370,N_46135);
or U46538 (N_46538,N_46198,N_46223);
nor U46539 (N_46539,N_46022,N_46399);
nor U46540 (N_46540,N_46231,N_46379);
or U46541 (N_46541,N_46389,N_46017);
or U46542 (N_46542,N_46346,N_46266);
and U46543 (N_46543,N_46490,N_46284);
nand U46544 (N_46544,N_46091,N_46130);
nand U46545 (N_46545,N_46395,N_46107);
nor U46546 (N_46546,N_46010,N_46041);
nor U46547 (N_46547,N_46364,N_46065);
and U46548 (N_46548,N_46340,N_46243);
or U46549 (N_46549,N_46426,N_46225);
xor U46550 (N_46550,N_46400,N_46250);
xnor U46551 (N_46551,N_46467,N_46079);
xor U46552 (N_46552,N_46078,N_46449);
and U46553 (N_46553,N_46230,N_46034);
and U46554 (N_46554,N_46056,N_46007);
xor U46555 (N_46555,N_46363,N_46274);
nand U46556 (N_46556,N_46396,N_46401);
and U46557 (N_46557,N_46071,N_46180);
nor U46558 (N_46558,N_46247,N_46276);
or U46559 (N_46559,N_46431,N_46436);
or U46560 (N_46560,N_46162,N_46006);
and U46561 (N_46561,N_46365,N_46015);
xnor U46562 (N_46562,N_46184,N_46300);
nand U46563 (N_46563,N_46492,N_46140);
or U46564 (N_46564,N_46355,N_46151);
or U46565 (N_46565,N_46382,N_46260);
nand U46566 (N_46566,N_46039,N_46083);
nand U46567 (N_46567,N_46117,N_46259);
nor U46568 (N_46568,N_46104,N_46028);
and U46569 (N_46569,N_46292,N_46344);
or U46570 (N_46570,N_46185,N_46414);
and U46571 (N_46571,N_46275,N_46106);
or U46572 (N_46572,N_46374,N_46304);
or U46573 (N_46573,N_46255,N_46486);
or U46574 (N_46574,N_46322,N_46047);
and U46575 (N_46575,N_46462,N_46146);
and U46576 (N_46576,N_46373,N_46222);
xor U46577 (N_46577,N_46415,N_46261);
nor U46578 (N_46578,N_46348,N_46293);
nand U46579 (N_46579,N_46197,N_46376);
or U46580 (N_46580,N_46451,N_46342);
xnor U46581 (N_46581,N_46439,N_46393);
xor U46582 (N_46582,N_46152,N_46145);
or U46583 (N_46583,N_46290,N_46070);
nor U46584 (N_46584,N_46128,N_46123);
or U46585 (N_46585,N_46210,N_46457);
nor U46586 (N_46586,N_46496,N_46177);
and U46587 (N_46587,N_46148,N_46196);
nor U46588 (N_46588,N_46088,N_46466);
nand U46589 (N_46589,N_46445,N_46361);
or U46590 (N_46590,N_46423,N_46043);
or U46591 (N_46591,N_46429,N_46216);
and U46592 (N_46592,N_46252,N_46150);
nand U46593 (N_46593,N_46470,N_46269);
and U46594 (N_46594,N_46138,N_46330);
nor U46595 (N_46595,N_46495,N_46481);
xor U46596 (N_46596,N_46446,N_46176);
nand U46597 (N_46597,N_46030,N_46411);
nand U46598 (N_46598,N_46334,N_46406);
nand U46599 (N_46599,N_46402,N_46064);
nand U46600 (N_46600,N_46328,N_46310);
and U46601 (N_46601,N_46326,N_46450);
nor U46602 (N_46602,N_46422,N_46092);
or U46603 (N_46603,N_46318,N_46263);
nor U46604 (N_46604,N_46120,N_46084);
or U46605 (N_46605,N_46100,N_46497);
and U46606 (N_46606,N_46287,N_46080);
nor U46607 (N_46607,N_46273,N_46137);
and U46608 (N_46608,N_46160,N_46191);
or U46609 (N_46609,N_46127,N_46291);
and U46610 (N_46610,N_46478,N_46483);
and U46611 (N_46611,N_46491,N_46207);
nand U46612 (N_46612,N_46311,N_46256);
or U46613 (N_46613,N_46157,N_46044);
and U46614 (N_46614,N_46186,N_46331);
or U46615 (N_46615,N_46321,N_46076);
nor U46616 (N_46616,N_46053,N_46189);
nor U46617 (N_46617,N_46212,N_46036);
nand U46618 (N_46618,N_46384,N_46410);
nand U46619 (N_46619,N_46405,N_46024);
nand U46620 (N_46620,N_46066,N_46417);
or U46621 (N_46621,N_46245,N_46166);
or U46622 (N_46622,N_46240,N_46472);
and U46623 (N_46623,N_46012,N_46179);
nand U46624 (N_46624,N_46412,N_46244);
or U46625 (N_46625,N_46193,N_46479);
or U46626 (N_46626,N_46167,N_46215);
nand U46627 (N_46627,N_46089,N_46339);
or U46628 (N_46628,N_46062,N_46258);
and U46629 (N_46629,N_46040,N_46155);
xnor U46630 (N_46630,N_46221,N_46208);
nor U46631 (N_46631,N_46004,N_46025);
or U46632 (N_46632,N_46283,N_46368);
or U46633 (N_46633,N_46205,N_46357);
and U46634 (N_46634,N_46099,N_46134);
or U46635 (N_46635,N_46383,N_46413);
xnor U46636 (N_46636,N_46067,N_46418);
nor U46637 (N_46637,N_46116,N_46430);
nor U46638 (N_46638,N_46013,N_46109);
nor U46639 (N_46639,N_46228,N_46254);
nor U46640 (N_46640,N_46060,N_46278);
and U46641 (N_46641,N_46394,N_46169);
nor U46642 (N_46642,N_46095,N_46153);
or U46643 (N_46643,N_46388,N_46420);
xor U46644 (N_46644,N_46069,N_46404);
nor U46645 (N_46645,N_46103,N_46268);
nand U46646 (N_46646,N_46075,N_46407);
xnor U46647 (N_46647,N_46063,N_46493);
xnor U46648 (N_46648,N_46049,N_46277);
and U46649 (N_46649,N_46362,N_46473);
nand U46650 (N_46650,N_46073,N_46380);
nor U46651 (N_46651,N_46232,N_46332);
nor U46652 (N_46652,N_46110,N_46301);
xor U46653 (N_46653,N_46016,N_46021);
and U46654 (N_46654,N_46282,N_46350);
and U46655 (N_46655,N_46308,N_46336);
nand U46656 (N_46656,N_46224,N_46390);
nand U46657 (N_46657,N_46093,N_46499);
nor U46658 (N_46658,N_46476,N_46387);
or U46659 (N_46659,N_46253,N_46159);
or U46660 (N_46660,N_46154,N_46317);
or U46661 (N_46661,N_46081,N_46124);
nor U46662 (N_46662,N_46072,N_46171);
nand U46663 (N_46663,N_46183,N_46366);
nand U46664 (N_46664,N_46202,N_46391);
or U46665 (N_46665,N_46443,N_46101);
nand U46666 (N_46666,N_46285,N_46057);
and U46667 (N_46667,N_46170,N_46129);
and U46668 (N_46668,N_46435,N_46425);
xor U46669 (N_46669,N_46037,N_46438);
nor U46670 (N_46670,N_46033,N_46345);
nand U46671 (N_46671,N_46377,N_46020);
and U46672 (N_46672,N_46453,N_46314);
or U46673 (N_46673,N_46098,N_46307);
or U46674 (N_46674,N_46121,N_46094);
and U46675 (N_46675,N_46009,N_46061);
or U46676 (N_46676,N_46018,N_46048);
nand U46677 (N_46677,N_46347,N_46082);
nand U46678 (N_46678,N_46441,N_46315);
nand U46679 (N_46679,N_46320,N_46264);
or U46680 (N_46680,N_46027,N_46023);
nand U46681 (N_46681,N_46329,N_46003);
nor U46682 (N_46682,N_46477,N_46455);
and U46683 (N_46683,N_46265,N_46452);
and U46684 (N_46684,N_46141,N_46227);
and U46685 (N_46685,N_46190,N_46424);
nand U46686 (N_46686,N_46178,N_46113);
and U46687 (N_46687,N_46298,N_46419);
nand U46688 (N_46688,N_46487,N_46338);
or U46689 (N_46689,N_46220,N_46257);
or U46690 (N_46690,N_46026,N_46485);
nand U46691 (N_46691,N_46090,N_46046);
nand U46692 (N_46692,N_46042,N_46454);
nor U46693 (N_46693,N_46213,N_46369);
nand U46694 (N_46694,N_46204,N_46102);
and U46695 (N_46695,N_46156,N_46484);
and U46696 (N_46696,N_46447,N_46163);
and U46697 (N_46697,N_46238,N_46058);
or U46698 (N_46698,N_46488,N_46398);
and U46699 (N_46699,N_46172,N_46444);
or U46700 (N_46700,N_46459,N_46335);
nor U46701 (N_46701,N_46126,N_46174);
nand U46702 (N_46702,N_46341,N_46421);
and U46703 (N_46703,N_46087,N_46005);
nand U46704 (N_46704,N_46119,N_46367);
nand U46705 (N_46705,N_46327,N_46354);
nand U46706 (N_46706,N_46226,N_46112);
or U46707 (N_46707,N_46052,N_46386);
nand U46708 (N_46708,N_46032,N_46029);
nand U46709 (N_46709,N_46475,N_46356);
nor U46710 (N_46710,N_46343,N_46381);
nand U46711 (N_46711,N_46349,N_46416);
nor U46712 (N_46712,N_46464,N_46372);
xnor U46713 (N_46713,N_46122,N_46440);
and U46714 (N_46714,N_46246,N_46008);
nand U46715 (N_46715,N_46086,N_46296);
nand U46716 (N_46716,N_46295,N_46313);
and U46717 (N_46717,N_46271,N_46456);
and U46718 (N_46718,N_46019,N_46217);
nor U46719 (N_46719,N_46409,N_46325);
and U46720 (N_46720,N_46059,N_46279);
or U46721 (N_46721,N_46077,N_46469);
nand U46722 (N_46722,N_46239,N_46437);
xor U46723 (N_46723,N_46281,N_46324);
or U46724 (N_46724,N_46233,N_46397);
nor U46725 (N_46725,N_46136,N_46114);
nor U46726 (N_46726,N_46323,N_46352);
nand U46727 (N_46727,N_46302,N_46306);
nor U46728 (N_46728,N_46206,N_46248);
xnor U46729 (N_46729,N_46195,N_46305);
and U46730 (N_46730,N_46428,N_46068);
nor U46731 (N_46731,N_46168,N_46142);
and U46732 (N_46732,N_46131,N_46432);
or U46733 (N_46733,N_46312,N_46303);
or U46734 (N_46734,N_46097,N_46139);
nand U46735 (N_46735,N_46333,N_46111);
and U46736 (N_46736,N_46158,N_46294);
nand U46737 (N_46737,N_46038,N_46385);
nor U46738 (N_46738,N_46125,N_46448);
or U46739 (N_46739,N_46050,N_46187);
or U46740 (N_46740,N_46147,N_46468);
or U46741 (N_46741,N_46465,N_46498);
nor U46742 (N_46742,N_46280,N_46235);
nor U46743 (N_46743,N_46319,N_46353);
nor U46744 (N_46744,N_46200,N_46286);
and U46745 (N_46745,N_46337,N_46234);
nand U46746 (N_46746,N_46242,N_46297);
and U46747 (N_46747,N_46000,N_46463);
and U46748 (N_46748,N_46494,N_46218);
or U46749 (N_46749,N_46375,N_46045);
and U46750 (N_46750,N_46212,N_46013);
nand U46751 (N_46751,N_46280,N_46301);
and U46752 (N_46752,N_46297,N_46472);
xor U46753 (N_46753,N_46122,N_46004);
xnor U46754 (N_46754,N_46083,N_46401);
or U46755 (N_46755,N_46128,N_46432);
nand U46756 (N_46756,N_46027,N_46375);
nand U46757 (N_46757,N_46255,N_46189);
nand U46758 (N_46758,N_46301,N_46349);
and U46759 (N_46759,N_46086,N_46308);
nand U46760 (N_46760,N_46204,N_46277);
and U46761 (N_46761,N_46139,N_46413);
or U46762 (N_46762,N_46100,N_46088);
nand U46763 (N_46763,N_46268,N_46301);
nand U46764 (N_46764,N_46393,N_46279);
and U46765 (N_46765,N_46391,N_46408);
nand U46766 (N_46766,N_46295,N_46165);
xnor U46767 (N_46767,N_46468,N_46455);
nor U46768 (N_46768,N_46440,N_46134);
and U46769 (N_46769,N_46280,N_46333);
or U46770 (N_46770,N_46218,N_46030);
xnor U46771 (N_46771,N_46407,N_46260);
or U46772 (N_46772,N_46188,N_46291);
nor U46773 (N_46773,N_46134,N_46359);
nand U46774 (N_46774,N_46222,N_46130);
and U46775 (N_46775,N_46017,N_46217);
nand U46776 (N_46776,N_46216,N_46167);
or U46777 (N_46777,N_46472,N_46287);
nand U46778 (N_46778,N_46075,N_46472);
xor U46779 (N_46779,N_46079,N_46233);
xor U46780 (N_46780,N_46450,N_46099);
and U46781 (N_46781,N_46135,N_46336);
and U46782 (N_46782,N_46071,N_46203);
nand U46783 (N_46783,N_46132,N_46161);
or U46784 (N_46784,N_46174,N_46244);
nand U46785 (N_46785,N_46388,N_46498);
and U46786 (N_46786,N_46212,N_46087);
nor U46787 (N_46787,N_46181,N_46260);
xor U46788 (N_46788,N_46421,N_46149);
nor U46789 (N_46789,N_46138,N_46122);
or U46790 (N_46790,N_46318,N_46132);
nand U46791 (N_46791,N_46453,N_46228);
nor U46792 (N_46792,N_46029,N_46127);
nand U46793 (N_46793,N_46349,N_46386);
and U46794 (N_46794,N_46365,N_46449);
or U46795 (N_46795,N_46306,N_46220);
nand U46796 (N_46796,N_46063,N_46081);
nor U46797 (N_46797,N_46497,N_46128);
nand U46798 (N_46798,N_46152,N_46293);
or U46799 (N_46799,N_46089,N_46233);
nor U46800 (N_46800,N_46482,N_46399);
or U46801 (N_46801,N_46262,N_46165);
or U46802 (N_46802,N_46038,N_46421);
xor U46803 (N_46803,N_46342,N_46030);
nand U46804 (N_46804,N_46197,N_46458);
or U46805 (N_46805,N_46162,N_46462);
nand U46806 (N_46806,N_46017,N_46456);
or U46807 (N_46807,N_46412,N_46448);
xnor U46808 (N_46808,N_46462,N_46067);
nand U46809 (N_46809,N_46224,N_46455);
nand U46810 (N_46810,N_46230,N_46052);
nand U46811 (N_46811,N_46033,N_46340);
nor U46812 (N_46812,N_46345,N_46296);
nor U46813 (N_46813,N_46228,N_46183);
xnor U46814 (N_46814,N_46046,N_46129);
nand U46815 (N_46815,N_46135,N_46392);
nor U46816 (N_46816,N_46434,N_46093);
xor U46817 (N_46817,N_46038,N_46459);
nor U46818 (N_46818,N_46052,N_46271);
and U46819 (N_46819,N_46286,N_46223);
nor U46820 (N_46820,N_46325,N_46214);
nand U46821 (N_46821,N_46286,N_46107);
nor U46822 (N_46822,N_46320,N_46387);
and U46823 (N_46823,N_46281,N_46411);
nand U46824 (N_46824,N_46446,N_46419);
and U46825 (N_46825,N_46144,N_46150);
xnor U46826 (N_46826,N_46296,N_46275);
nand U46827 (N_46827,N_46131,N_46112);
or U46828 (N_46828,N_46277,N_46253);
nor U46829 (N_46829,N_46375,N_46080);
and U46830 (N_46830,N_46158,N_46103);
nor U46831 (N_46831,N_46302,N_46073);
nand U46832 (N_46832,N_46265,N_46118);
or U46833 (N_46833,N_46457,N_46451);
or U46834 (N_46834,N_46370,N_46171);
and U46835 (N_46835,N_46292,N_46012);
and U46836 (N_46836,N_46452,N_46405);
or U46837 (N_46837,N_46219,N_46359);
or U46838 (N_46838,N_46011,N_46075);
xnor U46839 (N_46839,N_46007,N_46240);
or U46840 (N_46840,N_46292,N_46219);
and U46841 (N_46841,N_46100,N_46286);
nor U46842 (N_46842,N_46391,N_46411);
nor U46843 (N_46843,N_46462,N_46107);
and U46844 (N_46844,N_46215,N_46413);
nor U46845 (N_46845,N_46323,N_46061);
and U46846 (N_46846,N_46202,N_46056);
and U46847 (N_46847,N_46386,N_46406);
nor U46848 (N_46848,N_46491,N_46060);
xor U46849 (N_46849,N_46141,N_46132);
xor U46850 (N_46850,N_46436,N_46214);
nand U46851 (N_46851,N_46138,N_46357);
or U46852 (N_46852,N_46408,N_46184);
and U46853 (N_46853,N_46276,N_46430);
or U46854 (N_46854,N_46236,N_46341);
or U46855 (N_46855,N_46362,N_46133);
and U46856 (N_46856,N_46453,N_46386);
nand U46857 (N_46857,N_46337,N_46414);
nor U46858 (N_46858,N_46339,N_46001);
and U46859 (N_46859,N_46165,N_46137);
or U46860 (N_46860,N_46406,N_46049);
nand U46861 (N_46861,N_46235,N_46404);
nand U46862 (N_46862,N_46357,N_46304);
nand U46863 (N_46863,N_46423,N_46130);
xnor U46864 (N_46864,N_46405,N_46281);
or U46865 (N_46865,N_46211,N_46045);
nand U46866 (N_46866,N_46124,N_46357);
or U46867 (N_46867,N_46035,N_46125);
and U46868 (N_46868,N_46436,N_46250);
and U46869 (N_46869,N_46299,N_46302);
nand U46870 (N_46870,N_46433,N_46217);
nand U46871 (N_46871,N_46167,N_46245);
nor U46872 (N_46872,N_46327,N_46182);
nand U46873 (N_46873,N_46467,N_46308);
nand U46874 (N_46874,N_46350,N_46133);
nand U46875 (N_46875,N_46331,N_46466);
xor U46876 (N_46876,N_46499,N_46158);
xnor U46877 (N_46877,N_46410,N_46378);
or U46878 (N_46878,N_46272,N_46498);
and U46879 (N_46879,N_46311,N_46195);
nand U46880 (N_46880,N_46445,N_46131);
xor U46881 (N_46881,N_46144,N_46275);
nor U46882 (N_46882,N_46177,N_46010);
and U46883 (N_46883,N_46301,N_46271);
nor U46884 (N_46884,N_46220,N_46468);
xnor U46885 (N_46885,N_46494,N_46180);
nor U46886 (N_46886,N_46425,N_46200);
nor U46887 (N_46887,N_46464,N_46364);
or U46888 (N_46888,N_46499,N_46279);
or U46889 (N_46889,N_46242,N_46389);
and U46890 (N_46890,N_46457,N_46299);
nand U46891 (N_46891,N_46028,N_46160);
or U46892 (N_46892,N_46209,N_46250);
or U46893 (N_46893,N_46230,N_46297);
nor U46894 (N_46894,N_46337,N_46043);
or U46895 (N_46895,N_46109,N_46263);
nand U46896 (N_46896,N_46371,N_46057);
nor U46897 (N_46897,N_46345,N_46391);
or U46898 (N_46898,N_46163,N_46428);
nand U46899 (N_46899,N_46056,N_46182);
nand U46900 (N_46900,N_46117,N_46025);
nand U46901 (N_46901,N_46288,N_46032);
and U46902 (N_46902,N_46196,N_46107);
nor U46903 (N_46903,N_46352,N_46225);
and U46904 (N_46904,N_46354,N_46380);
and U46905 (N_46905,N_46394,N_46243);
or U46906 (N_46906,N_46286,N_46068);
or U46907 (N_46907,N_46159,N_46488);
nor U46908 (N_46908,N_46254,N_46065);
or U46909 (N_46909,N_46202,N_46441);
xnor U46910 (N_46910,N_46430,N_46280);
nand U46911 (N_46911,N_46050,N_46474);
xnor U46912 (N_46912,N_46012,N_46155);
nor U46913 (N_46913,N_46481,N_46112);
nor U46914 (N_46914,N_46349,N_46288);
or U46915 (N_46915,N_46038,N_46415);
nand U46916 (N_46916,N_46271,N_46090);
and U46917 (N_46917,N_46074,N_46124);
or U46918 (N_46918,N_46313,N_46028);
nor U46919 (N_46919,N_46093,N_46401);
nor U46920 (N_46920,N_46165,N_46021);
and U46921 (N_46921,N_46119,N_46326);
and U46922 (N_46922,N_46188,N_46386);
and U46923 (N_46923,N_46384,N_46318);
or U46924 (N_46924,N_46459,N_46483);
nand U46925 (N_46925,N_46312,N_46488);
or U46926 (N_46926,N_46231,N_46233);
nor U46927 (N_46927,N_46266,N_46060);
and U46928 (N_46928,N_46200,N_46311);
xor U46929 (N_46929,N_46016,N_46145);
and U46930 (N_46930,N_46463,N_46461);
nor U46931 (N_46931,N_46343,N_46432);
nand U46932 (N_46932,N_46099,N_46064);
or U46933 (N_46933,N_46284,N_46034);
xnor U46934 (N_46934,N_46020,N_46071);
and U46935 (N_46935,N_46330,N_46461);
nor U46936 (N_46936,N_46103,N_46428);
nor U46937 (N_46937,N_46259,N_46113);
xor U46938 (N_46938,N_46276,N_46216);
and U46939 (N_46939,N_46376,N_46174);
and U46940 (N_46940,N_46357,N_46380);
nand U46941 (N_46941,N_46089,N_46174);
and U46942 (N_46942,N_46476,N_46380);
and U46943 (N_46943,N_46358,N_46429);
xnor U46944 (N_46944,N_46431,N_46216);
xor U46945 (N_46945,N_46414,N_46221);
and U46946 (N_46946,N_46068,N_46329);
and U46947 (N_46947,N_46099,N_46416);
xnor U46948 (N_46948,N_46483,N_46358);
or U46949 (N_46949,N_46104,N_46246);
nand U46950 (N_46950,N_46063,N_46011);
xnor U46951 (N_46951,N_46415,N_46161);
and U46952 (N_46952,N_46229,N_46336);
or U46953 (N_46953,N_46391,N_46297);
and U46954 (N_46954,N_46135,N_46341);
or U46955 (N_46955,N_46260,N_46383);
and U46956 (N_46956,N_46396,N_46102);
nand U46957 (N_46957,N_46176,N_46212);
nor U46958 (N_46958,N_46468,N_46162);
nor U46959 (N_46959,N_46196,N_46204);
nand U46960 (N_46960,N_46393,N_46444);
nand U46961 (N_46961,N_46482,N_46354);
or U46962 (N_46962,N_46379,N_46145);
nor U46963 (N_46963,N_46290,N_46110);
and U46964 (N_46964,N_46483,N_46124);
nand U46965 (N_46965,N_46284,N_46157);
or U46966 (N_46966,N_46391,N_46033);
nor U46967 (N_46967,N_46395,N_46484);
nor U46968 (N_46968,N_46449,N_46158);
xor U46969 (N_46969,N_46119,N_46015);
and U46970 (N_46970,N_46101,N_46130);
nand U46971 (N_46971,N_46324,N_46177);
nand U46972 (N_46972,N_46210,N_46010);
nand U46973 (N_46973,N_46198,N_46123);
xnor U46974 (N_46974,N_46138,N_46160);
or U46975 (N_46975,N_46430,N_46439);
and U46976 (N_46976,N_46258,N_46116);
nand U46977 (N_46977,N_46350,N_46174);
and U46978 (N_46978,N_46484,N_46372);
nand U46979 (N_46979,N_46280,N_46419);
nand U46980 (N_46980,N_46140,N_46299);
nor U46981 (N_46981,N_46415,N_46254);
nand U46982 (N_46982,N_46131,N_46160);
and U46983 (N_46983,N_46152,N_46305);
nand U46984 (N_46984,N_46000,N_46297);
nor U46985 (N_46985,N_46286,N_46332);
or U46986 (N_46986,N_46103,N_46420);
and U46987 (N_46987,N_46301,N_46385);
or U46988 (N_46988,N_46192,N_46166);
or U46989 (N_46989,N_46238,N_46262);
nor U46990 (N_46990,N_46321,N_46331);
xnor U46991 (N_46991,N_46145,N_46463);
or U46992 (N_46992,N_46060,N_46207);
and U46993 (N_46993,N_46470,N_46320);
and U46994 (N_46994,N_46310,N_46345);
nor U46995 (N_46995,N_46277,N_46152);
and U46996 (N_46996,N_46318,N_46123);
nor U46997 (N_46997,N_46228,N_46186);
or U46998 (N_46998,N_46322,N_46318);
xor U46999 (N_46999,N_46299,N_46031);
nand U47000 (N_47000,N_46629,N_46870);
nand U47001 (N_47001,N_46945,N_46669);
or U47002 (N_47002,N_46983,N_46982);
or U47003 (N_47003,N_46840,N_46925);
nand U47004 (N_47004,N_46697,N_46984);
or U47005 (N_47005,N_46685,N_46847);
and U47006 (N_47006,N_46689,N_46839);
nand U47007 (N_47007,N_46572,N_46949);
or U47008 (N_47008,N_46814,N_46961);
xor U47009 (N_47009,N_46594,N_46642);
and U47010 (N_47010,N_46536,N_46844);
nor U47011 (N_47011,N_46716,N_46987);
and U47012 (N_47012,N_46862,N_46765);
and U47013 (N_47013,N_46729,N_46922);
nand U47014 (N_47014,N_46653,N_46526);
or U47015 (N_47015,N_46905,N_46745);
nor U47016 (N_47016,N_46752,N_46662);
nor U47017 (N_47017,N_46767,N_46746);
and U47018 (N_47018,N_46970,N_46943);
and U47019 (N_47019,N_46728,N_46613);
nor U47020 (N_47020,N_46780,N_46656);
nor U47021 (N_47021,N_46515,N_46712);
or U47022 (N_47022,N_46644,N_46545);
nand U47023 (N_47023,N_46991,N_46963);
nand U47024 (N_47024,N_46919,N_46518);
nor U47025 (N_47025,N_46665,N_46530);
and U47026 (N_47026,N_46574,N_46514);
and U47027 (N_47027,N_46828,N_46869);
or U47028 (N_47028,N_46579,N_46565);
or U47029 (N_47029,N_46886,N_46956);
nor U47030 (N_47030,N_46528,N_46820);
and U47031 (N_47031,N_46638,N_46819);
nor U47032 (N_47032,N_46757,N_46842);
nand U47033 (N_47033,N_46798,N_46512);
nor U47034 (N_47034,N_46965,N_46584);
or U47035 (N_47035,N_46604,N_46951);
nand U47036 (N_47036,N_46749,N_46960);
nand U47037 (N_47037,N_46535,N_46880);
nand U47038 (N_47038,N_46845,N_46836);
nor U47039 (N_47039,N_46873,N_46702);
nand U47040 (N_47040,N_46748,N_46505);
or U47041 (N_47041,N_46585,N_46760);
or U47042 (N_47042,N_46599,N_46672);
or U47043 (N_47043,N_46529,N_46999);
or U47044 (N_47044,N_46639,N_46687);
nand U47045 (N_47045,N_46776,N_46795);
and U47046 (N_47046,N_46583,N_46944);
or U47047 (N_47047,N_46540,N_46829);
or U47048 (N_47048,N_46722,N_46877);
xor U47049 (N_47049,N_46813,N_46502);
nor U47050 (N_47050,N_46582,N_46854);
xor U47051 (N_47051,N_46668,N_46994);
or U47052 (N_47052,N_46710,N_46695);
and U47053 (N_47053,N_46513,N_46742);
and U47054 (N_47054,N_46903,N_46622);
nand U47055 (N_47055,N_46802,N_46974);
nand U47056 (N_47056,N_46577,N_46875);
and U47057 (N_47057,N_46643,N_46589);
nand U47058 (N_47058,N_46511,N_46785);
nor U47059 (N_47059,N_46831,N_46586);
nor U47060 (N_47060,N_46867,N_46857);
and U47061 (N_47061,N_46849,N_46773);
or U47062 (N_47062,N_46976,N_46504);
and U47063 (N_47063,N_46835,N_46939);
nor U47064 (N_47064,N_46830,N_46608);
nand U47065 (N_47065,N_46959,N_46507);
and U47066 (N_47066,N_46704,N_46995);
nand U47067 (N_47067,N_46630,N_46544);
nand U47068 (N_47068,N_46894,N_46985);
nand U47069 (N_47069,N_46954,N_46726);
nand U47070 (N_47070,N_46524,N_46966);
nor U47071 (N_47071,N_46759,N_46724);
or U47072 (N_47072,N_46821,N_46861);
or U47073 (N_47073,N_46611,N_46986);
or U47074 (N_47074,N_46764,N_46996);
or U47075 (N_47075,N_46688,N_46874);
nand U47076 (N_47076,N_46800,N_46901);
and U47077 (N_47077,N_46787,N_46631);
or U47078 (N_47078,N_46603,N_46698);
xor U47079 (N_47079,N_46834,N_46678);
xor U47080 (N_47080,N_46932,N_46935);
xnor U47081 (N_47081,N_46768,N_46595);
and U47082 (N_47082,N_46897,N_46917);
nand U47083 (N_47083,N_46560,N_46633);
or U47084 (N_47084,N_46715,N_46937);
nand U47085 (N_47085,N_46872,N_46906);
or U47086 (N_47086,N_46988,N_46805);
and U47087 (N_47087,N_46660,N_46924);
or U47088 (N_47088,N_46566,N_46509);
or U47089 (N_47089,N_46676,N_46626);
and U47090 (N_47090,N_46717,N_46900);
or U47091 (N_47091,N_46896,N_46812);
and U47092 (N_47092,N_46868,N_46910);
nand U47093 (N_47093,N_46701,N_46827);
or U47094 (N_47094,N_46538,N_46789);
nand U47095 (N_47095,N_46694,N_46720);
and U47096 (N_47096,N_46684,N_46997);
nand U47097 (N_47097,N_46573,N_46967);
nor U47098 (N_47098,N_46761,N_46989);
nand U47099 (N_47099,N_46731,N_46593);
and U47100 (N_47100,N_46636,N_46667);
and U47101 (N_47101,N_46580,N_46592);
or U47102 (N_47102,N_46686,N_46755);
nand U47103 (N_47103,N_46774,N_46568);
nand U47104 (N_47104,N_46576,N_46531);
or U47105 (N_47105,N_46751,N_46602);
nand U47106 (N_47106,N_46693,N_46898);
and U47107 (N_47107,N_46794,N_46570);
or U47108 (N_47108,N_46930,N_46516);
nand U47109 (N_47109,N_46915,N_46882);
or U47110 (N_47110,N_46851,N_46889);
and U47111 (N_47111,N_46973,N_46623);
nor U47112 (N_47112,N_46750,N_46635);
xnor U47113 (N_47113,N_46615,N_46581);
nor U47114 (N_47114,N_46806,N_46777);
and U47115 (N_47115,N_46914,N_46858);
nor U47116 (N_47116,N_46918,N_46879);
and U47117 (N_47117,N_46853,N_46534);
nor U47118 (N_47118,N_46838,N_46904);
or U47119 (N_47119,N_46876,N_46571);
and U47120 (N_47120,N_46620,N_46519);
nand U47121 (N_47121,N_46679,N_46542);
or U47122 (N_47122,N_46654,N_46981);
and U47123 (N_47123,N_46552,N_46683);
or U47124 (N_47124,N_46744,N_46508);
and U47125 (N_47125,N_46895,N_46887);
nor U47126 (N_47126,N_46646,N_46523);
nor U47127 (N_47127,N_46779,N_46899);
xnor U47128 (N_47128,N_46569,N_46992);
nand U47129 (N_47129,N_46527,N_46969);
or U47130 (N_47130,N_46826,N_46975);
xor U47131 (N_47131,N_46559,N_46625);
nor U47132 (N_47132,N_46561,N_46650);
nor U47133 (N_47133,N_46766,N_46664);
xnor U47134 (N_47134,N_46929,N_46637);
and U47135 (N_47135,N_46763,N_46549);
or U47136 (N_47136,N_46605,N_46815);
or U47137 (N_47137,N_46558,N_46762);
or U47138 (N_47138,N_46968,N_46737);
nor U47139 (N_47139,N_46972,N_46675);
and U47140 (N_47140,N_46856,N_46553);
nor U47141 (N_47141,N_46804,N_46707);
or U47142 (N_47142,N_46657,N_46883);
nand U47143 (N_47143,N_46913,N_46781);
and U47144 (N_47144,N_46543,N_46567);
nand U47145 (N_47145,N_46947,N_46733);
and U47146 (N_47146,N_46998,N_46866);
nand U47147 (N_47147,N_46993,N_46647);
nor U47148 (N_47148,N_46634,N_46713);
and U47149 (N_47149,N_46846,N_46628);
and U47150 (N_47150,N_46788,N_46546);
nor U47151 (N_47151,N_46618,N_46539);
xnor U47152 (N_47152,N_46841,N_46727);
nand U47153 (N_47153,N_46597,N_46934);
nand U47154 (N_47154,N_46933,N_46769);
nand U47155 (N_47155,N_46817,N_46740);
or U47156 (N_47156,N_46962,N_46770);
xor U47157 (N_47157,N_46865,N_46738);
or U47158 (N_47158,N_46714,N_46557);
or U47159 (N_47159,N_46892,N_46923);
nand U47160 (N_47160,N_46578,N_46554);
or U47161 (N_47161,N_46703,N_46940);
nand U47162 (N_47162,N_46550,N_46601);
nand U47163 (N_47163,N_46790,N_46734);
xnor U47164 (N_47164,N_46736,N_46772);
nand U47165 (N_47165,N_46670,N_46721);
and U47166 (N_47166,N_46801,N_46616);
nand U47167 (N_47167,N_46600,N_46786);
and U47168 (N_47168,N_46797,N_46941);
nor U47169 (N_47169,N_46718,N_46907);
and U47170 (N_47170,N_46500,N_46658);
nor U47171 (N_47171,N_46852,N_46690);
nor U47172 (N_47172,N_46556,N_46663);
or U47173 (N_47173,N_46659,N_46708);
nand U47174 (N_47174,N_46803,N_46958);
or U47175 (N_47175,N_46885,N_46501);
nand U47176 (N_47176,N_46575,N_46799);
xnor U47177 (N_47177,N_46950,N_46606);
nand U47178 (N_47178,N_46607,N_46893);
and U47179 (N_47179,N_46506,N_46735);
nand U47180 (N_47180,N_46522,N_46541);
nor U47181 (N_47181,N_46902,N_46548);
nand U47182 (N_47182,N_46909,N_46624);
nand U47183 (N_47183,N_46822,N_46564);
nand U47184 (N_47184,N_46723,N_46725);
xnor U47185 (N_47185,N_46691,N_46948);
nor U47186 (N_47186,N_46871,N_46641);
and U47187 (N_47187,N_46833,N_46588);
nor U47188 (N_47188,N_46640,N_46942);
nand U47189 (N_47189,N_46916,N_46673);
nor U47190 (N_47190,N_46621,N_46741);
nor U47191 (N_47191,N_46955,N_46730);
nand U47192 (N_47192,N_46587,N_46562);
nor U47193 (N_47193,N_46807,N_46520);
and U47194 (N_47194,N_46931,N_46783);
nand U47195 (N_47195,N_46911,N_46980);
nand U47196 (N_47196,N_46610,N_46758);
or U47197 (N_47197,N_46743,N_46649);
or U47198 (N_47198,N_46732,N_46719);
nand U47199 (N_47199,N_46920,N_46705);
nand U47200 (N_47200,N_46699,N_46936);
or U47201 (N_47201,N_46946,N_46859);
nor U47202 (N_47202,N_46928,N_46843);
or U47203 (N_47203,N_46775,N_46816);
xnor U47204 (N_47204,N_46739,N_46661);
nor U47205 (N_47205,N_46824,N_46677);
and U47206 (N_47206,N_46537,N_46927);
nor U47207 (N_47207,N_46778,N_46706);
and U47208 (N_47208,N_46614,N_46525);
xnor U47209 (N_47209,N_46696,N_46666);
nand U47210 (N_47210,N_46890,N_46979);
nand U47211 (N_47211,N_46837,N_46521);
or U47212 (N_47212,N_46503,N_46848);
and U47213 (N_47213,N_46971,N_46860);
nor U47214 (N_47214,N_46793,N_46754);
nand U47215 (N_47215,N_46555,N_46655);
nor U47216 (N_47216,N_46791,N_46964);
and U47217 (N_47217,N_46632,N_46792);
or U47218 (N_47218,N_46921,N_46957);
and U47219 (N_47219,N_46609,N_46912);
and U47220 (N_47220,N_46590,N_46818);
nand U47221 (N_47221,N_46612,N_46598);
and U47222 (N_47222,N_46711,N_46952);
or U47223 (N_47223,N_46864,N_46532);
nand U47224 (N_47224,N_46888,N_46510);
nand U47225 (N_47225,N_46619,N_46850);
nand U47226 (N_47226,N_46908,N_46878);
nor U47227 (N_47227,N_46809,N_46617);
nand U47228 (N_47228,N_46674,N_46978);
or U47229 (N_47229,N_46591,N_46596);
and U47230 (N_47230,N_46648,N_46753);
or U47231 (N_47231,N_46682,N_46680);
nor U47232 (N_47232,N_46855,N_46796);
and U47233 (N_47233,N_46784,N_46782);
or U47234 (N_47234,N_46891,N_46771);
nand U47235 (N_47235,N_46563,N_46671);
nand U47236 (N_47236,N_46681,N_46926);
xor U47237 (N_47237,N_46700,N_46533);
nor U47238 (N_47238,N_46547,N_46517);
nand U47239 (N_47239,N_46810,N_46977);
nand U47240 (N_47240,N_46881,N_46811);
and U47241 (N_47241,N_46884,N_46645);
and U47242 (N_47242,N_46938,N_46953);
or U47243 (N_47243,N_46692,N_46823);
and U47244 (N_47244,N_46627,N_46825);
nand U47245 (N_47245,N_46651,N_46756);
or U47246 (N_47246,N_46709,N_46832);
nand U47247 (N_47247,N_46747,N_46863);
nand U47248 (N_47248,N_46990,N_46551);
nand U47249 (N_47249,N_46808,N_46652);
nand U47250 (N_47250,N_46756,N_46753);
and U47251 (N_47251,N_46610,N_46624);
xnor U47252 (N_47252,N_46673,N_46503);
or U47253 (N_47253,N_46730,N_46795);
and U47254 (N_47254,N_46663,N_46959);
nand U47255 (N_47255,N_46775,N_46774);
and U47256 (N_47256,N_46698,N_46983);
or U47257 (N_47257,N_46962,N_46778);
nor U47258 (N_47258,N_46852,N_46771);
nor U47259 (N_47259,N_46955,N_46669);
nand U47260 (N_47260,N_46952,N_46590);
or U47261 (N_47261,N_46627,N_46936);
nor U47262 (N_47262,N_46933,N_46910);
or U47263 (N_47263,N_46954,N_46995);
or U47264 (N_47264,N_46919,N_46560);
and U47265 (N_47265,N_46626,N_46624);
nor U47266 (N_47266,N_46999,N_46863);
nand U47267 (N_47267,N_46914,N_46868);
and U47268 (N_47268,N_46961,N_46957);
and U47269 (N_47269,N_46768,N_46566);
xnor U47270 (N_47270,N_46646,N_46569);
xor U47271 (N_47271,N_46902,N_46585);
or U47272 (N_47272,N_46937,N_46943);
and U47273 (N_47273,N_46596,N_46557);
nand U47274 (N_47274,N_46775,N_46524);
and U47275 (N_47275,N_46710,N_46561);
nand U47276 (N_47276,N_46915,N_46590);
or U47277 (N_47277,N_46625,N_46921);
or U47278 (N_47278,N_46556,N_46884);
nand U47279 (N_47279,N_46771,N_46915);
or U47280 (N_47280,N_46958,N_46768);
and U47281 (N_47281,N_46844,N_46859);
or U47282 (N_47282,N_46852,N_46663);
nor U47283 (N_47283,N_46836,N_46975);
nand U47284 (N_47284,N_46720,N_46843);
nor U47285 (N_47285,N_46953,N_46527);
nor U47286 (N_47286,N_46615,N_46889);
or U47287 (N_47287,N_46659,N_46669);
and U47288 (N_47288,N_46778,N_46900);
and U47289 (N_47289,N_46957,N_46666);
nor U47290 (N_47290,N_46735,N_46624);
xnor U47291 (N_47291,N_46843,N_46966);
xor U47292 (N_47292,N_46559,N_46549);
nand U47293 (N_47293,N_46763,N_46684);
or U47294 (N_47294,N_46913,N_46581);
or U47295 (N_47295,N_46564,N_46526);
or U47296 (N_47296,N_46918,N_46969);
nand U47297 (N_47297,N_46975,N_46814);
or U47298 (N_47298,N_46585,N_46730);
nor U47299 (N_47299,N_46885,N_46984);
nor U47300 (N_47300,N_46622,N_46718);
and U47301 (N_47301,N_46790,N_46627);
nor U47302 (N_47302,N_46965,N_46524);
nor U47303 (N_47303,N_46548,N_46573);
and U47304 (N_47304,N_46785,N_46548);
nand U47305 (N_47305,N_46701,N_46824);
nor U47306 (N_47306,N_46746,N_46819);
and U47307 (N_47307,N_46880,N_46626);
and U47308 (N_47308,N_46662,N_46900);
and U47309 (N_47309,N_46852,N_46748);
nand U47310 (N_47310,N_46715,N_46924);
nand U47311 (N_47311,N_46752,N_46955);
nor U47312 (N_47312,N_46925,N_46976);
or U47313 (N_47313,N_46735,N_46689);
nand U47314 (N_47314,N_46643,N_46732);
nor U47315 (N_47315,N_46983,N_46835);
and U47316 (N_47316,N_46650,N_46858);
nor U47317 (N_47317,N_46633,N_46792);
nand U47318 (N_47318,N_46707,N_46622);
or U47319 (N_47319,N_46573,N_46976);
xor U47320 (N_47320,N_46557,N_46547);
and U47321 (N_47321,N_46686,N_46744);
and U47322 (N_47322,N_46800,N_46838);
and U47323 (N_47323,N_46608,N_46639);
or U47324 (N_47324,N_46649,N_46606);
nor U47325 (N_47325,N_46707,N_46544);
nor U47326 (N_47326,N_46944,N_46980);
or U47327 (N_47327,N_46667,N_46567);
or U47328 (N_47328,N_46514,N_46756);
nand U47329 (N_47329,N_46883,N_46691);
xor U47330 (N_47330,N_46954,N_46563);
and U47331 (N_47331,N_46951,N_46852);
nand U47332 (N_47332,N_46910,N_46640);
or U47333 (N_47333,N_46879,N_46735);
nor U47334 (N_47334,N_46773,N_46910);
and U47335 (N_47335,N_46811,N_46529);
and U47336 (N_47336,N_46552,N_46798);
or U47337 (N_47337,N_46925,N_46594);
nand U47338 (N_47338,N_46944,N_46639);
nor U47339 (N_47339,N_46523,N_46712);
and U47340 (N_47340,N_46884,N_46712);
nand U47341 (N_47341,N_46615,N_46771);
nor U47342 (N_47342,N_46961,N_46866);
nand U47343 (N_47343,N_46730,N_46866);
nor U47344 (N_47344,N_46930,N_46725);
or U47345 (N_47345,N_46533,N_46977);
and U47346 (N_47346,N_46798,N_46882);
or U47347 (N_47347,N_46624,N_46611);
and U47348 (N_47348,N_46619,N_46724);
or U47349 (N_47349,N_46718,N_46599);
or U47350 (N_47350,N_46794,N_46843);
nand U47351 (N_47351,N_46940,N_46960);
nor U47352 (N_47352,N_46818,N_46525);
or U47353 (N_47353,N_46754,N_46813);
nand U47354 (N_47354,N_46617,N_46868);
nor U47355 (N_47355,N_46810,N_46759);
or U47356 (N_47356,N_46800,N_46886);
nor U47357 (N_47357,N_46701,N_46705);
and U47358 (N_47358,N_46970,N_46621);
xnor U47359 (N_47359,N_46574,N_46677);
or U47360 (N_47360,N_46542,N_46792);
nand U47361 (N_47361,N_46757,N_46930);
nor U47362 (N_47362,N_46754,N_46539);
nor U47363 (N_47363,N_46953,N_46815);
or U47364 (N_47364,N_46580,N_46893);
nor U47365 (N_47365,N_46777,N_46690);
nor U47366 (N_47366,N_46677,N_46842);
or U47367 (N_47367,N_46998,N_46673);
and U47368 (N_47368,N_46575,N_46536);
or U47369 (N_47369,N_46548,N_46696);
nor U47370 (N_47370,N_46703,N_46556);
nand U47371 (N_47371,N_46984,N_46875);
nand U47372 (N_47372,N_46847,N_46989);
nor U47373 (N_47373,N_46726,N_46695);
xnor U47374 (N_47374,N_46745,N_46670);
nand U47375 (N_47375,N_46909,N_46933);
or U47376 (N_47376,N_46548,N_46603);
xnor U47377 (N_47377,N_46845,N_46721);
nor U47378 (N_47378,N_46847,N_46661);
or U47379 (N_47379,N_46540,N_46934);
nand U47380 (N_47380,N_46792,N_46851);
and U47381 (N_47381,N_46680,N_46754);
and U47382 (N_47382,N_46918,N_46810);
and U47383 (N_47383,N_46853,N_46575);
or U47384 (N_47384,N_46825,N_46670);
nor U47385 (N_47385,N_46833,N_46856);
and U47386 (N_47386,N_46527,N_46751);
or U47387 (N_47387,N_46604,N_46734);
and U47388 (N_47388,N_46717,N_46589);
nand U47389 (N_47389,N_46633,N_46810);
nor U47390 (N_47390,N_46699,N_46706);
nand U47391 (N_47391,N_46926,N_46830);
and U47392 (N_47392,N_46709,N_46684);
and U47393 (N_47393,N_46929,N_46764);
nand U47394 (N_47394,N_46563,N_46904);
and U47395 (N_47395,N_46510,N_46853);
or U47396 (N_47396,N_46959,N_46737);
nand U47397 (N_47397,N_46945,N_46705);
or U47398 (N_47398,N_46996,N_46651);
xnor U47399 (N_47399,N_46617,N_46950);
nand U47400 (N_47400,N_46604,N_46528);
nor U47401 (N_47401,N_46955,N_46811);
nand U47402 (N_47402,N_46645,N_46916);
nor U47403 (N_47403,N_46858,N_46802);
nor U47404 (N_47404,N_46590,N_46691);
nand U47405 (N_47405,N_46821,N_46551);
nand U47406 (N_47406,N_46588,N_46881);
nor U47407 (N_47407,N_46788,N_46935);
xor U47408 (N_47408,N_46551,N_46537);
nand U47409 (N_47409,N_46567,N_46844);
nand U47410 (N_47410,N_46566,N_46999);
and U47411 (N_47411,N_46918,N_46780);
or U47412 (N_47412,N_46635,N_46818);
xor U47413 (N_47413,N_46765,N_46700);
or U47414 (N_47414,N_46991,N_46565);
nor U47415 (N_47415,N_46685,N_46691);
and U47416 (N_47416,N_46765,N_46515);
nand U47417 (N_47417,N_46754,N_46887);
or U47418 (N_47418,N_46717,N_46547);
xnor U47419 (N_47419,N_46797,N_46695);
and U47420 (N_47420,N_46748,N_46612);
nor U47421 (N_47421,N_46931,N_46503);
or U47422 (N_47422,N_46873,N_46907);
nor U47423 (N_47423,N_46813,N_46785);
xnor U47424 (N_47424,N_46920,N_46926);
nand U47425 (N_47425,N_46816,N_46555);
xor U47426 (N_47426,N_46719,N_46661);
nor U47427 (N_47427,N_46742,N_46723);
xor U47428 (N_47428,N_46803,N_46973);
or U47429 (N_47429,N_46743,N_46769);
nand U47430 (N_47430,N_46957,N_46553);
nor U47431 (N_47431,N_46515,N_46811);
nand U47432 (N_47432,N_46980,N_46643);
and U47433 (N_47433,N_46874,N_46716);
or U47434 (N_47434,N_46628,N_46763);
nand U47435 (N_47435,N_46804,N_46812);
nand U47436 (N_47436,N_46666,N_46817);
or U47437 (N_47437,N_46577,N_46688);
nand U47438 (N_47438,N_46550,N_46986);
nand U47439 (N_47439,N_46929,N_46543);
nor U47440 (N_47440,N_46909,N_46628);
nand U47441 (N_47441,N_46950,N_46762);
or U47442 (N_47442,N_46837,N_46529);
nand U47443 (N_47443,N_46578,N_46926);
or U47444 (N_47444,N_46885,N_46502);
nor U47445 (N_47445,N_46949,N_46948);
nand U47446 (N_47446,N_46619,N_46912);
and U47447 (N_47447,N_46692,N_46565);
and U47448 (N_47448,N_46659,N_46755);
nor U47449 (N_47449,N_46951,N_46673);
and U47450 (N_47450,N_46565,N_46773);
xor U47451 (N_47451,N_46656,N_46511);
nand U47452 (N_47452,N_46986,N_46896);
or U47453 (N_47453,N_46511,N_46882);
nor U47454 (N_47454,N_46740,N_46812);
xor U47455 (N_47455,N_46763,N_46522);
and U47456 (N_47456,N_46850,N_46683);
xnor U47457 (N_47457,N_46530,N_46919);
or U47458 (N_47458,N_46583,N_46514);
and U47459 (N_47459,N_46684,N_46692);
nor U47460 (N_47460,N_46980,N_46774);
or U47461 (N_47461,N_46688,N_46782);
or U47462 (N_47462,N_46572,N_46716);
nor U47463 (N_47463,N_46835,N_46793);
nand U47464 (N_47464,N_46992,N_46972);
and U47465 (N_47465,N_46669,N_46831);
nor U47466 (N_47466,N_46889,N_46697);
and U47467 (N_47467,N_46969,N_46875);
and U47468 (N_47468,N_46621,N_46725);
nand U47469 (N_47469,N_46540,N_46958);
xor U47470 (N_47470,N_46930,N_46584);
or U47471 (N_47471,N_46580,N_46904);
or U47472 (N_47472,N_46746,N_46764);
or U47473 (N_47473,N_46611,N_46995);
nand U47474 (N_47474,N_46731,N_46517);
xor U47475 (N_47475,N_46745,N_46914);
nand U47476 (N_47476,N_46605,N_46672);
or U47477 (N_47477,N_46901,N_46672);
nand U47478 (N_47478,N_46507,N_46906);
and U47479 (N_47479,N_46844,N_46977);
xor U47480 (N_47480,N_46894,N_46591);
nor U47481 (N_47481,N_46545,N_46560);
or U47482 (N_47482,N_46979,N_46784);
and U47483 (N_47483,N_46530,N_46702);
nand U47484 (N_47484,N_46588,N_46572);
nor U47485 (N_47485,N_46795,N_46908);
and U47486 (N_47486,N_46959,N_46693);
and U47487 (N_47487,N_46931,N_46720);
or U47488 (N_47488,N_46937,N_46525);
nand U47489 (N_47489,N_46521,N_46707);
nor U47490 (N_47490,N_46713,N_46675);
and U47491 (N_47491,N_46762,N_46832);
nor U47492 (N_47492,N_46801,N_46837);
nor U47493 (N_47493,N_46898,N_46977);
nand U47494 (N_47494,N_46586,N_46528);
or U47495 (N_47495,N_46968,N_46742);
nand U47496 (N_47496,N_46558,N_46501);
xor U47497 (N_47497,N_46770,N_46542);
or U47498 (N_47498,N_46901,N_46745);
nand U47499 (N_47499,N_46640,N_46554);
and U47500 (N_47500,N_47066,N_47315);
nand U47501 (N_47501,N_47223,N_47329);
xor U47502 (N_47502,N_47033,N_47252);
nand U47503 (N_47503,N_47455,N_47103);
nor U47504 (N_47504,N_47399,N_47101);
or U47505 (N_47505,N_47105,N_47124);
nand U47506 (N_47506,N_47338,N_47367);
nor U47507 (N_47507,N_47487,N_47100);
and U47508 (N_47508,N_47218,N_47012);
nand U47509 (N_47509,N_47092,N_47258);
or U47510 (N_47510,N_47490,N_47387);
or U47511 (N_47511,N_47467,N_47028);
or U47512 (N_47512,N_47266,N_47286);
nand U47513 (N_47513,N_47144,N_47323);
or U47514 (N_47514,N_47169,N_47190);
or U47515 (N_47515,N_47165,N_47217);
or U47516 (N_47516,N_47001,N_47304);
nand U47517 (N_47517,N_47435,N_47000);
or U47518 (N_47518,N_47226,N_47061);
or U47519 (N_47519,N_47275,N_47204);
nand U47520 (N_47520,N_47088,N_47018);
and U47521 (N_47521,N_47414,N_47240);
or U47522 (N_47522,N_47307,N_47216);
xnor U47523 (N_47523,N_47401,N_47276);
nand U47524 (N_47524,N_47043,N_47071);
and U47525 (N_47525,N_47324,N_47040);
or U47526 (N_47526,N_47164,N_47462);
or U47527 (N_47527,N_47354,N_47433);
nand U47528 (N_47528,N_47412,N_47316);
nand U47529 (N_47529,N_47042,N_47384);
nor U47530 (N_47530,N_47446,N_47023);
xor U47531 (N_47531,N_47402,N_47129);
and U47532 (N_47532,N_47491,N_47182);
nor U47533 (N_47533,N_47256,N_47498);
and U47534 (N_47534,N_47158,N_47044);
nor U47535 (N_47535,N_47097,N_47121);
nor U47536 (N_47536,N_47213,N_47283);
nor U47537 (N_47537,N_47377,N_47478);
nor U47538 (N_47538,N_47034,N_47448);
nor U47539 (N_47539,N_47476,N_47429);
or U47540 (N_47540,N_47398,N_47020);
and U47541 (N_47541,N_47473,N_47149);
nor U47542 (N_47542,N_47115,N_47472);
or U47543 (N_47543,N_47015,N_47123);
xnor U47544 (N_47544,N_47450,N_47239);
nor U47545 (N_47545,N_47395,N_47362);
nor U47546 (N_47546,N_47055,N_47209);
nand U47547 (N_47547,N_47137,N_47425);
and U47548 (N_47548,N_47003,N_47198);
nor U47549 (N_47549,N_47379,N_47150);
or U47550 (N_47550,N_47375,N_47094);
nor U47551 (N_47551,N_47328,N_47480);
or U47552 (N_47552,N_47152,N_47441);
and U47553 (N_47553,N_47408,N_47278);
nor U47554 (N_47554,N_47026,N_47053);
nand U47555 (N_47555,N_47070,N_47037);
or U47556 (N_47556,N_47447,N_47471);
or U47557 (N_47557,N_47443,N_47393);
and U47558 (N_47558,N_47048,N_47288);
nand U47559 (N_47559,N_47267,N_47006);
nand U47560 (N_47560,N_47325,N_47093);
or U47561 (N_47561,N_47135,N_47078);
nor U47562 (N_47562,N_47493,N_47394);
nor U47563 (N_47563,N_47131,N_47380);
nor U47564 (N_47564,N_47067,N_47069);
or U47565 (N_47565,N_47259,N_47013);
nor U47566 (N_47566,N_47306,N_47424);
nor U47567 (N_47567,N_47335,N_47475);
or U47568 (N_47568,N_47326,N_47434);
and U47569 (N_47569,N_47214,N_47389);
xnor U47570 (N_47570,N_47457,N_47073);
xor U47571 (N_47571,N_47219,N_47481);
and U47572 (N_47572,N_47297,N_47438);
and U47573 (N_47573,N_47489,N_47064);
nor U47574 (N_47574,N_47268,N_47157);
and U47575 (N_47575,N_47415,N_47247);
nor U47576 (N_47576,N_47059,N_47386);
or U47577 (N_47577,N_47045,N_47253);
and U47578 (N_47578,N_47255,N_47177);
nor U47579 (N_47579,N_47349,N_47086);
nor U47580 (N_47580,N_47459,N_47179);
or U47581 (N_47581,N_47230,N_47180);
and U47582 (N_47582,N_47257,N_47147);
nor U47583 (N_47583,N_47280,N_47080);
or U47584 (N_47584,N_47461,N_47321);
or U47585 (N_47585,N_47336,N_47156);
or U47586 (N_47586,N_47451,N_47248);
or U47587 (N_47587,N_47373,N_47482);
xnor U47588 (N_47588,N_47337,N_47126);
and U47589 (N_47589,N_47273,N_47263);
nor U47590 (N_47590,N_47250,N_47232);
or U47591 (N_47591,N_47151,N_47363);
nor U47592 (N_47592,N_47351,N_47109);
or U47593 (N_47593,N_47272,N_47162);
or U47594 (N_47594,N_47465,N_47102);
nand U47595 (N_47595,N_47021,N_47167);
nor U47596 (N_47596,N_47153,N_47269);
nand U47597 (N_47597,N_47423,N_47111);
or U47598 (N_47598,N_47422,N_47206);
and U47599 (N_47599,N_47056,N_47293);
nand U47600 (N_47600,N_47175,N_47385);
nand U47601 (N_47601,N_47074,N_47041);
nand U47602 (N_47602,N_47492,N_47166);
and U47603 (N_47603,N_47350,N_47205);
and U47604 (N_47604,N_47388,N_47227);
nand U47605 (N_47605,N_47311,N_47090);
nand U47606 (N_47606,N_47188,N_47127);
nor U47607 (N_47607,N_47265,N_47348);
nor U47608 (N_47608,N_47495,N_47108);
nand U47609 (N_47609,N_47104,N_47212);
or U47610 (N_47610,N_47468,N_47030);
and U47611 (N_47611,N_47322,N_47346);
and U47612 (N_47612,N_47072,N_47353);
nor U47613 (N_47613,N_47284,N_47183);
nand U47614 (N_47614,N_47031,N_47008);
and U47615 (N_47615,N_47222,N_47305);
nand U47616 (N_47616,N_47174,N_47430);
nor U47617 (N_47617,N_47159,N_47303);
nor U47618 (N_47618,N_47317,N_47211);
nand U47619 (N_47619,N_47196,N_47413);
nor U47620 (N_47620,N_47087,N_47359);
xnor U47621 (N_47621,N_47002,N_47197);
nor U47622 (N_47622,N_47371,N_47405);
or U47623 (N_47623,N_47397,N_47428);
nor U47624 (N_47624,N_47215,N_47300);
nand U47625 (N_47625,N_47485,N_47095);
nand U47626 (N_47626,N_47107,N_47187);
nand U47627 (N_47627,N_47199,N_47208);
nor U47628 (N_47628,N_47075,N_47302);
nor U47629 (N_47629,N_47310,N_47005);
nor U47630 (N_47630,N_47084,N_47235);
nor U47631 (N_47631,N_47486,N_47010);
or U47632 (N_47632,N_47444,N_47301);
or U47633 (N_47633,N_47148,N_47463);
and U47634 (N_47634,N_47277,N_47185);
or U47635 (N_47635,N_47085,N_47421);
or U47636 (N_47636,N_47130,N_47029);
nand U47637 (N_47637,N_47391,N_47369);
nor U47638 (N_47638,N_47281,N_47051);
nand U47639 (N_47639,N_47117,N_47155);
nor U47640 (N_47640,N_47309,N_47125);
nor U47641 (N_47641,N_47356,N_47036);
xnor U47642 (N_47642,N_47192,N_47173);
nor U47643 (N_47643,N_47054,N_47396);
and U47644 (N_47644,N_47499,N_47091);
or U47645 (N_47645,N_47096,N_47243);
and U47646 (N_47646,N_47469,N_47342);
or U47647 (N_47647,N_47017,N_47110);
and U47648 (N_47648,N_47494,N_47210);
and U47649 (N_47649,N_47296,N_47334);
and U47650 (N_47650,N_47260,N_47294);
or U47651 (N_47651,N_47254,N_47083);
or U47652 (N_47652,N_47050,N_47418);
xor U47653 (N_47653,N_47186,N_47119);
and U47654 (N_47654,N_47345,N_47470);
nor U47655 (N_47655,N_47058,N_47202);
nor U47656 (N_47656,N_47079,N_47314);
xor U47657 (N_47657,N_47057,N_47238);
or U47658 (N_47658,N_47406,N_47496);
xnor U47659 (N_47659,N_47331,N_47392);
or U47660 (N_47660,N_47292,N_47466);
nor U47661 (N_47661,N_47047,N_47274);
xnor U47662 (N_47662,N_47114,N_47483);
and U47663 (N_47663,N_47228,N_47403);
and U47664 (N_47664,N_47138,N_47365);
nor U47665 (N_47665,N_47207,N_47178);
nor U47666 (N_47666,N_47464,N_47344);
or U47667 (N_47667,N_47060,N_47407);
or U47668 (N_47668,N_47333,N_47172);
nand U47669 (N_47669,N_47411,N_47065);
nand U47670 (N_47670,N_47452,N_47193);
nor U47671 (N_47671,N_47308,N_47035);
nand U47672 (N_47672,N_47390,N_47236);
or U47673 (N_47673,N_47132,N_47246);
and U47674 (N_47674,N_47383,N_47370);
or U47675 (N_47675,N_47376,N_47231);
or U47676 (N_47676,N_47319,N_47357);
xnor U47677 (N_47677,N_47437,N_47409);
nor U47678 (N_47678,N_47161,N_47032);
nand U47679 (N_47679,N_47460,N_47264);
or U47680 (N_47680,N_47019,N_47237);
nor U47681 (N_47681,N_47171,N_47025);
or U47682 (N_47682,N_47427,N_47458);
nor U47683 (N_47683,N_47416,N_47378);
xor U47684 (N_47684,N_47241,N_47176);
nand U47685 (N_47685,N_47453,N_47233);
xnor U47686 (N_47686,N_47251,N_47244);
and U47687 (N_47687,N_47442,N_47089);
or U47688 (N_47688,N_47439,N_47191);
and U47689 (N_47689,N_47113,N_47189);
nand U47690 (N_47690,N_47364,N_47400);
and U47691 (N_47691,N_47488,N_47068);
and U47692 (N_47692,N_47339,N_47221);
or U47693 (N_47693,N_47249,N_47295);
or U47694 (N_47694,N_47082,N_47320);
xor U47695 (N_47695,N_47194,N_47099);
and U47696 (N_47696,N_47360,N_47220);
nor U47697 (N_47697,N_47184,N_47039);
nand U47698 (N_47698,N_47122,N_47352);
and U47699 (N_47699,N_47229,N_47106);
and U47700 (N_47700,N_47134,N_47361);
and U47701 (N_47701,N_47046,N_47477);
nand U47702 (N_47702,N_47142,N_47168);
xor U47703 (N_47703,N_47062,N_47340);
and U47704 (N_47704,N_47016,N_47063);
nand U47705 (N_47705,N_47456,N_47245);
nor U47706 (N_47706,N_47140,N_47291);
or U47707 (N_47707,N_47382,N_47143);
nor U47708 (N_47708,N_47234,N_47436);
or U47709 (N_47709,N_47312,N_47410);
nor U47710 (N_47710,N_47454,N_47009);
and U47711 (N_47711,N_47139,N_47497);
or U47712 (N_47712,N_47195,N_47170);
and U47713 (N_47713,N_47038,N_47022);
nand U47714 (N_47714,N_47118,N_47474);
and U47715 (N_47715,N_47154,N_47076);
nor U47716 (N_47716,N_47136,N_47327);
nand U47717 (N_47717,N_47014,N_47440);
nand U47718 (N_47718,N_47287,N_47270);
nand U47719 (N_47719,N_47049,N_47372);
or U47720 (N_47720,N_47479,N_47330);
or U47721 (N_47721,N_47160,N_47011);
and U47722 (N_47722,N_47116,N_47381);
nand U47723 (N_47723,N_47081,N_47431);
xnor U47724 (N_47724,N_47449,N_47366);
nor U47725 (N_47725,N_47289,N_47261);
nand U47726 (N_47726,N_47298,N_47484);
nor U47727 (N_47727,N_47313,N_47358);
nand U47728 (N_47728,N_47343,N_47290);
or U47729 (N_47729,N_47098,N_47341);
nand U47730 (N_47730,N_47445,N_47432);
nor U47731 (N_47731,N_47024,N_47112);
and U47732 (N_47732,N_47355,N_47133);
and U47733 (N_47733,N_47285,N_47120);
nand U47734 (N_47734,N_47420,N_47200);
nor U47735 (N_47735,N_47368,N_47262);
and U47736 (N_47736,N_47282,N_47225);
and U47737 (N_47737,N_47299,N_47077);
or U47738 (N_47738,N_47201,N_47332);
nand U47739 (N_47739,N_47027,N_47145);
nand U47740 (N_47740,N_47146,N_47419);
or U47741 (N_47741,N_47271,N_47141);
nor U47742 (N_47742,N_47203,N_47347);
nand U47743 (N_47743,N_47374,N_47426);
and U47744 (N_47744,N_47417,N_47163);
nor U47745 (N_47745,N_47007,N_47004);
nor U47746 (N_47746,N_47181,N_47404);
or U47747 (N_47747,N_47318,N_47242);
nor U47748 (N_47748,N_47279,N_47224);
or U47749 (N_47749,N_47128,N_47052);
and U47750 (N_47750,N_47357,N_47193);
xor U47751 (N_47751,N_47348,N_47061);
and U47752 (N_47752,N_47258,N_47298);
and U47753 (N_47753,N_47058,N_47035);
nand U47754 (N_47754,N_47317,N_47202);
or U47755 (N_47755,N_47221,N_47338);
and U47756 (N_47756,N_47289,N_47104);
nand U47757 (N_47757,N_47074,N_47047);
or U47758 (N_47758,N_47036,N_47375);
and U47759 (N_47759,N_47062,N_47449);
nor U47760 (N_47760,N_47256,N_47274);
or U47761 (N_47761,N_47255,N_47276);
or U47762 (N_47762,N_47371,N_47079);
and U47763 (N_47763,N_47421,N_47492);
and U47764 (N_47764,N_47427,N_47286);
or U47765 (N_47765,N_47153,N_47407);
nor U47766 (N_47766,N_47471,N_47466);
nand U47767 (N_47767,N_47155,N_47351);
and U47768 (N_47768,N_47026,N_47456);
nand U47769 (N_47769,N_47342,N_47258);
or U47770 (N_47770,N_47121,N_47163);
or U47771 (N_47771,N_47429,N_47415);
xor U47772 (N_47772,N_47223,N_47272);
xor U47773 (N_47773,N_47117,N_47281);
nor U47774 (N_47774,N_47469,N_47472);
nand U47775 (N_47775,N_47364,N_47100);
nor U47776 (N_47776,N_47374,N_47246);
nor U47777 (N_47777,N_47201,N_47191);
or U47778 (N_47778,N_47085,N_47492);
nand U47779 (N_47779,N_47110,N_47294);
or U47780 (N_47780,N_47254,N_47356);
nor U47781 (N_47781,N_47109,N_47274);
nand U47782 (N_47782,N_47355,N_47010);
nand U47783 (N_47783,N_47423,N_47312);
nand U47784 (N_47784,N_47472,N_47203);
or U47785 (N_47785,N_47107,N_47291);
or U47786 (N_47786,N_47021,N_47288);
nor U47787 (N_47787,N_47184,N_47139);
nor U47788 (N_47788,N_47206,N_47339);
nand U47789 (N_47789,N_47344,N_47067);
nor U47790 (N_47790,N_47306,N_47294);
or U47791 (N_47791,N_47060,N_47117);
xnor U47792 (N_47792,N_47181,N_47496);
nand U47793 (N_47793,N_47416,N_47084);
or U47794 (N_47794,N_47063,N_47321);
xor U47795 (N_47795,N_47354,N_47248);
nor U47796 (N_47796,N_47207,N_47395);
nor U47797 (N_47797,N_47337,N_47095);
nand U47798 (N_47798,N_47012,N_47034);
nor U47799 (N_47799,N_47190,N_47307);
nand U47800 (N_47800,N_47247,N_47229);
or U47801 (N_47801,N_47491,N_47126);
nand U47802 (N_47802,N_47408,N_47158);
nand U47803 (N_47803,N_47438,N_47317);
nand U47804 (N_47804,N_47131,N_47268);
nor U47805 (N_47805,N_47438,N_47455);
nor U47806 (N_47806,N_47215,N_47410);
nand U47807 (N_47807,N_47095,N_47060);
or U47808 (N_47808,N_47131,N_47221);
xor U47809 (N_47809,N_47128,N_47304);
or U47810 (N_47810,N_47188,N_47285);
or U47811 (N_47811,N_47126,N_47108);
and U47812 (N_47812,N_47458,N_47132);
nor U47813 (N_47813,N_47184,N_47150);
nor U47814 (N_47814,N_47326,N_47070);
nand U47815 (N_47815,N_47025,N_47493);
and U47816 (N_47816,N_47405,N_47433);
or U47817 (N_47817,N_47080,N_47023);
and U47818 (N_47818,N_47466,N_47293);
xor U47819 (N_47819,N_47442,N_47335);
and U47820 (N_47820,N_47386,N_47274);
xor U47821 (N_47821,N_47489,N_47079);
nor U47822 (N_47822,N_47226,N_47433);
nor U47823 (N_47823,N_47027,N_47434);
or U47824 (N_47824,N_47237,N_47078);
nand U47825 (N_47825,N_47429,N_47056);
and U47826 (N_47826,N_47288,N_47059);
nand U47827 (N_47827,N_47174,N_47168);
or U47828 (N_47828,N_47095,N_47027);
or U47829 (N_47829,N_47014,N_47217);
or U47830 (N_47830,N_47022,N_47212);
or U47831 (N_47831,N_47270,N_47156);
nand U47832 (N_47832,N_47368,N_47143);
nor U47833 (N_47833,N_47130,N_47079);
nor U47834 (N_47834,N_47066,N_47280);
or U47835 (N_47835,N_47355,N_47482);
or U47836 (N_47836,N_47309,N_47410);
nor U47837 (N_47837,N_47443,N_47372);
and U47838 (N_47838,N_47458,N_47002);
or U47839 (N_47839,N_47353,N_47334);
and U47840 (N_47840,N_47343,N_47137);
nand U47841 (N_47841,N_47301,N_47136);
xor U47842 (N_47842,N_47141,N_47034);
and U47843 (N_47843,N_47404,N_47068);
nor U47844 (N_47844,N_47154,N_47394);
or U47845 (N_47845,N_47067,N_47342);
and U47846 (N_47846,N_47140,N_47278);
and U47847 (N_47847,N_47156,N_47230);
nor U47848 (N_47848,N_47328,N_47403);
and U47849 (N_47849,N_47296,N_47011);
nor U47850 (N_47850,N_47461,N_47139);
and U47851 (N_47851,N_47113,N_47358);
and U47852 (N_47852,N_47452,N_47409);
nand U47853 (N_47853,N_47057,N_47254);
and U47854 (N_47854,N_47237,N_47176);
nand U47855 (N_47855,N_47128,N_47031);
and U47856 (N_47856,N_47023,N_47056);
nor U47857 (N_47857,N_47039,N_47289);
or U47858 (N_47858,N_47331,N_47180);
and U47859 (N_47859,N_47407,N_47189);
or U47860 (N_47860,N_47486,N_47374);
or U47861 (N_47861,N_47388,N_47140);
xnor U47862 (N_47862,N_47234,N_47137);
nand U47863 (N_47863,N_47357,N_47299);
and U47864 (N_47864,N_47388,N_47193);
xor U47865 (N_47865,N_47302,N_47372);
nor U47866 (N_47866,N_47375,N_47132);
nor U47867 (N_47867,N_47447,N_47062);
and U47868 (N_47868,N_47421,N_47445);
and U47869 (N_47869,N_47294,N_47230);
nand U47870 (N_47870,N_47057,N_47417);
or U47871 (N_47871,N_47475,N_47261);
nand U47872 (N_47872,N_47355,N_47360);
and U47873 (N_47873,N_47150,N_47039);
nand U47874 (N_47874,N_47150,N_47143);
and U47875 (N_47875,N_47150,N_47297);
nand U47876 (N_47876,N_47371,N_47066);
and U47877 (N_47877,N_47466,N_47188);
and U47878 (N_47878,N_47454,N_47326);
nor U47879 (N_47879,N_47410,N_47375);
nand U47880 (N_47880,N_47458,N_47182);
and U47881 (N_47881,N_47026,N_47248);
or U47882 (N_47882,N_47464,N_47440);
or U47883 (N_47883,N_47388,N_47195);
or U47884 (N_47884,N_47054,N_47248);
nand U47885 (N_47885,N_47273,N_47281);
nand U47886 (N_47886,N_47318,N_47108);
nor U47887 (N_47887,N_47139,N_47087);
nor U47888 (N_47888,N_47225,N_47429);
xnor U47889 (N_47889,N_47322,N_47288);
or U47890 (N_47890,N_47289,N_47334);
nor U47891 (N_47891,N_47351,N_47144);
nor U47892 (N_47892,N_47257,N_47345);
nor U47893 (N_47893,N_47006,N_47247);
nor U47894 (N_47894,N_47323,N_47197);
nor U47895 (N_47895,N_47403,N_47368);
nor U47896 (N_47896,N_47457,N_47433);
nand U47897 (N_47897,N_47061,N_47214);
or U47898 (N_47898,N_47293,N_47095);
or U47899 (N_47899,N_47206,N_47128);
nor U47900 (N_47900,N_47263,N_47459);
or U47901 (N_47901,N_47127,N_47160);
and U47902 (N_47902,N_47191,N_47052);
or U47903 (N_47903,N_47127,N_47281);
nand U47904 (N_47904,N_47308,N_47429);
nand U47905 (N_47905,N_47224,N_47498);
nor U47906 (N_47906,N_47400,N_47249);
and U47907 (N_47907,N_47270,N_47491);
nand U47908 (N_47908,N_47428,N_47339);
nor U47909 (N_47909,N_47299,N_47356);
or U47910 (N_47910,N_47344,N_47493);
nor U47911 (N_47911,N_47384,N_47323);
nand U47912 (N_47912,N_47223,N_47200);
or U47913 (N_47913,N_47370,N_47325);
or U47914 (N_47914,N_47139,N_47108);
and U47915 (N_47915,N_47398,N_47035);
or U47916 (N_47916,N_47407,N_47000);
nor U47917 (N_47917,N_47443,N_47203);
and U47918 (N_47918,N_47446,N_47309);
nor U47919 (N_47919,N_47264,N_47411);
nor U47920 (N_47920,N_47143,N_47342);
or U47921 (N_47921,N_47485,N_47425);
nand U47922 (N_47922,N_47133,N_47054);
nand U47923 (N_47923,N_47246,N_47461);
nor U47924 (N_47924,N_47358,N_47047);
nor U47925 (N_47925,N_47498,N_47051);
or U47926 (N_47926,N_47217,N_47184);
and U47927 (N_47927,N_47420,N_47379);
nor U47928 (N_47928,N_47387,N_47474);
nor U47929 (N_47929,N_47099,N_47092);
nand U47930 (N_47930,N_47324,N_47426);
nor U47931 (N_47931,N_47236,N_47113);
nor U47932 (N_47932,N_47361,N_47318);
or U47933 (N_47933,N_47190,N_47255);
nand U47934 (N_47934,N_47161,N_47014);
nand U47935 (N_47935,N_47278,N_47067);
nand U47936 (N_47936,N_47014,N_47407);
or U47937 (N_47937,N_47349,N_47433);
nand U47938 (N_47938,N_47494,N_47144);
nor U47939 (N_47939,N_47435,N_47439);
or U47940 (N_47940,N_47259,N_47053);
nor U47941 (N_47941,N_47377,N_47179);
or U47942 (N_47942,N_47153,N_47333);
or U47943 (N_47943,N_47098,N_47392);
or U47944 (N_47944,N_47287,N_47175);
nor U47945 (N_47945,N_47251,N_47091);
xor U47946 (N_47946,N_47173,N_47368);
and U47947 (N_47947,N_47243,N_47006);
or U47948 (N_47948,N_47224,N_47238);
nand U47949 (N_47949,N_47068,N_47107);
nor U47950 (N_47950,N_47080,N_47051);
or U47951 (N_47951,N_47227,N_47130);
or U47952 (N_47952,N_47332,N_47231);
or U47953 (N_47953,N_47425,N_47256);
nor U47954 (N_47954,N_47456,N_47007);
or U47955 (N_47955,N_47475,N_47351);
and U47956 (N_47956,N_47044,N_47375);
and U47957 (N_47957,N_47073,N_47016);
nand U47958 (N_47958,N_47275,N_47464);
and U47959 (N_47959,N_47252,N_47262);
or U47960 (N_47960,N_47370,N_47126);
or U47961 (N_47961,N_47432,N_47353);
or U47962 (N_47962,N_47068,N_47102);
nand U47963 (N_47963,N_47301,N_47144);
and U47964 (N_47964,N_47255,N_47458);
nand U47965 (N_47965,N_47141,N_47042);
or U47966 (N_47966,N_47060,N_47444);
or U47967 (N_47967,N_47296,N_47386);
nor U47968 (N_47968,N_47212,N_47103);
nand U47969 (N_47969,N_47087,N_47177);
or U47970 (N_47970,N_47287,N_47173);
nand U47971 (N_47971,N_47476,N_47402);
nand U47972 (N_47972,N_47222,N_47100);
and U47973 (N_47973,N_47032,N_47245);
nand U47974 (N_47974,N_47161,N_47184);
nand U47975 (N_47975,N_47167,N_47293);
nor U47976 (N_47976,N_47218,N_47246);
and U47977 (N_47977,N_47145,N_47443);
and U47978 (N_47978,N_47155,N_47165);
nand U47979 (N_47979,N_47333,N_47291);
nor U47980 (N_47980,N_47179,N_47118);
or U47981 (N_47981,N_47435,N_47154);
nand U47982 (N_47982,N_47152,N_47370);
xor U47983 (N_47983,N_47123,N_47446);
nor U47984 (N_47984,N_47320,N_47259);
nand U47985 (N_47985,N_47060,N_47363);
nand U47986 (N_47986,N_47038,N_47350);
nand U47987 (N_47987,N_47210,N_47275);
and U47988 (N_47988,N_47076,N_47060);
and U47989 (N_47989,N_47227,N_47105);
and U47990 (N_47990,N_47151,N_47306);
nor U47991 (N_47991,N_47026,N_47415);
nand U47992 (N_47992,N_47279,N_47296);
nand U47993 (N_47993,N_47238,N_47399);
and U47994 (N_47994,N_47396,N_47209);
or U47995 (N_47995,N_47020,N_47306);
and U47996 (N_47996,N_47312,N_47445);
and U47997 (N_47997,N_47045,N_47327);
nor U47998 (N_47998,N_47075,N_47187);
and U47999 (N_47999,N_47388,N_47407);
and U48000 (N_48000,N_47954,N_47635);
or U48001 (N_48001,N_47883,N_47513);
and U48002 (N_48002,N_47609,N_47777);
xnor U48003 (N_48003,N_47903,N_47727);
nor U48004 (N_48004,N_47991,N_47873);
nand U48005 (N_48005,N_47530,N_47826);
and U48006 (N_48006,N_47669,N_47736);
nor U48007 (N_48007,N_47834,N_47960);
nand U48008 (N_48008,N_47706,N_47857);
nor U48009 (N_48009,N_47810,N_47629);
nand U48010 (N_48010,N_47798,N_47648);
nand U48011 (N_48011,N_47713,N_47579);
or U48012 (N_48012,N_47967,N_47818);
nor U48013 (N_48013,N_47658,N_47984);
nand U48014 (N_48014,N_47731,N_47760);
nand U48015 (N_48015,N_47677,N_47787);
and U48016 (N_48016,N_47679,N_47612);
nor U48017 (N_48017,N_47910,N_47567);
nor U48018 (N_48018,N_47718,N_47772);
nand U48019 (N_48019,N_47992,N_47801);
nor U48020 (N_48020,N_47889,N_47596);
nor U48021 (N_48021,N_47781,N_47861);
nand U48022 (N_48022,N_47649,N_47887);
or U48023 (N_48023,N_47585,N_47763);
and U48024 (N_48024,N_47599,N_47837);
nand U48025 (N_48025,N_47730,N_47848);
and U48026 (N_48026,N_47556,N_47886);
nor U48027 (N_48027,N_47979,N_47690);
nor U48028 (N_48028,N_47842,N_47581);
nor U48029 (N_48029,N_47877,N_47605);
nor U48030 (N_48030,N_47944,N_47621);
nand U48031 (N_48031,N_47930,N_47571);
xor U48032 (N_48032,N_47866,N_47878);
nor U48033 (N_48033,N_47533,N_47687);
or U48034 (N_48034,N_47500,N_47568);
or U48035 (N_48035,N_47570,N_47696);
nand U48036 (N_48036,N_47720,N_47558);
or U48037 (N_48037,N_47752,N_47935);
or U48038 (N_48038,N_47539,N_47574);
or U48039 (N_48039,N_47789,N_47526);
nand U48040 (N_48040,N_47983,N_47628);
and U48041 (N_48041,N_47775,N_47901);
and U48042 (N_48042,N_47667,N_47729);
nand U48043 (N_48043,N_47817,N_47521);
and U48044 (N_48044,N_47623,N_47745);
or U48045 (N_48045,N_47898,N_47961);
and U48046 (N_48046,N_47823,N_47734);
and U48047 (N_48047,N_47660,N_47950);
or U48048 (N_48048,N_47917,N_47894);
and U48049 (N_48049,N_47754,N_47561);
and U48050 (N_48050,N_47790,N_47595);
xnor U48051 (N_48051,N_47590,N_47647);
and U48052 (N_48052,N_47914,N_47966);
and U48053 (N_48053,N_47562,N_47937);
or U48054 (N_48054,N_47583,N_47728);
nand U48055 (N_48055,N_47761,N_47924);
nand U48056 (N_48056,N_47929,N_47814);
nand U48057 (N_48057,N_47947,N_47618);
xnor U48058 (N_48058,N_47791,N_47515);
and U48059 (N_48059,N_47504,N_47938);
and U48060 (N_48060,N_47662,N_47698);
nand U48061 (N_48061,N_47815,N_47619);
nand U48062 (N_48062,N_47637,N_47587);
and U48063 (N_48063,N_47809,N_47964);
xnor U48064 (N_48064,N_47836,N_47970);
or U48065 (N_48065,N_47812,N_47594);
nand U48066 (N_48066,N_47650,N_47890);
nor U48067 (N_48067,N_47829,N_47719);
nand U48068 (N_48068,N_47525,N_47534);
or U48069 (N_48069,N_47514,N_47737);
nand U48070 (N_48070,N_47673,N_47545);
and U48071 (N_48071,N_47840,N_47926);
and U48072 (N_48072,N_47620,N_47633);
nand U48073 (N_48073,N_47502,N_47973);
and U48074 (N_48074,N_47614,N_47505);
xnor U48075 (N_48075,N_47674,N_47529);
nand U48076 (N_48076,N_47512,N_47601);
xor U48077 (N_48077,N_47990,N_47757);
xnor U48078 (N_48078,N_47661,N_47655);
or U48079 (N_48079,N_47506,N_47783);
nand U48080 (N_48080,N_47758,N_47700);
nand U48081 (N_48081,N_47535,N_47531);
nor U48082 (N_48082,N_47830,N_47805);
nor U48083 (N_48083,N_47880,N_47912);
and U48084 (N_48084,N_47527,N_47749);
and U48085 (N_48085,N_47824,N_47592);
nand U48086 (N_48086,N_47792,N_47785);
and U48087 (N_48087,N_47588,N_47872);
nor U48088 (N_48088,N_47904,N_47895);
nand U48089 (N_48089,N_47721,N_47780);
nor U48090 (N_48090,N_47600,N_47946);
nor U48091 (N_48091,N_47675,N_47831);
nor U48092 (N_48092,N_47701,N_47784);
xnor U48093 (N_48093,N_47897,N_47668);
or U48094 (N_48094,N_47551,N_47639);
or U48095 (N_48095,N_47825,N_47537);
or U48096 (N_48096,N_47835,N_47580);
nand U48097 (N_48097,N_47827,N_47766);
nand U48098 (N_48098,N_47578,N_47663);
or U48099 (N_48099,N_47833,N_47688);
nand U48100 (N_48100,N_47610,N_47799);
and U48101 (N_48101,N_47630,N_47975);
or U48102 (N_48102,N_47908,N_47987);
and U48103 (N_48103,N_47916,N_47750);
nor U48104 (N_48104,N_47869,N_47645);
or U48105 (N_48105,N_47516,N_47656);
nor U48106 (N_48106,N_47626,N_47849);
nor U48107 (N_48107,N_47949,N_47723);
nor U48108 (N_48108,N_47941,N_47747);
and U48109 (N_48109,N_47733,N_47510);
and U48110 (N_48110,N_47939,N_47786);
or U48111 (N_48111,N_47557,N_47739);
nor U48112 (N_48112,N_47998,N_47715);
and U48113 (N_48113,N_47816,N_47841);
nand U48114 (N_48114,N_47559,N_47968);
nor U48115 (N_48115,N_47928,N_47607);
and U48116 (N_48116,N_47552,N_47586);
nor U48117 (N_48117,N_47847,N_47519);
or U48118 (N_48118,N_47532,N_47523);
and U48119 (N_48119,N_47900,N_47804);
nand U48120 (N_48120,N_47778,N_47882);
nor U48121 (N_48121,N_47795,N_47803);
or U48122 (N_48122,N_47951,N_47572);
or U48123 (N_48123,N_47800,N_47710);
or U48124 (N_48124,N_47993,N_47683);
xor U48125 (N_48125,N_47615,N_47940);
nor U48126 (N_48126,N_47867,N_47691);
nor U48127 (N_48127,N_47909,N_47651);
nand U48128 (N_48128,N_47746,N_47709);
and U48129 (N_48129,N_47845,N_47714);
or U48130 (N_48130,N_47982,N_47971);
and U48131 (N_48131,N_47832,N_47918);
nand U48132 (N_48132,N_47874,N_47627);
or U48133 (N_48133,N_47759,N_47606);
or U48134 (N_48134,N_47591,N_47767);
or U48135 (N_48135,N_47722,N_47546);
or U48136 (N_48136,N_47755,N_47875);
or U48137 (N_48137,N_47896,N_47797);
and U48138 (N_48138,N_47931,N_47925);
nand U48139 (N_48139,N_47879,N_47554);
nor U48140 (N_48140,N_47892,N_47977);
or U48141 (N_48141,N_47576,N_47888);
and U48142 (N_48142,N_47646,N_47988);
nor U48143 (N_48143,N_47756,N_47996);
and U48144 (N_48144,N_47509,N_47632);
nor U48145 (N_48145,N_47779,N_47743);
nand U48146 (N_48146,N_47764,N_47828);
nand U48147 (N_48147,N_47859,N_47684);
or U48148 (N_48148,N_47744,N_47689);
nand U48149 (N_48149,N_47920,N_47997);
or U48150 (N_48150,N_47952,N_47616);
or U48151 (N_48151,N_47666,N_47905);
and U48152 (N_48152,N_47642,N_47943);
or U48153 (N_48153,N_47507,N_47582);
nor U48154 (N_48154,N_47770,N_47972);
nand U48155 (N_48155,N_47962,N_47547);
or U48156 (N_48156,N_47680,N_47707);
nand U48157 (N_48157,N_47697,N_47638);
or U48158 (N_48158,N_47520,N_47870);
nand U48159 (N_48159,N_47553,N_47643);
nor U48160 (N_48160,N_47564,N_47907);
and U48161 (N_48161,N_47994,N_47508);
nor U48162 (N_48162,N_47664,N_47919);
nor U48163 (N_48163,N_47604,N_47773);
nor U48164 (N_48164,N_47565,N_47819);
and U48165 (N_48165,N_47672,N_47838);
xor U48166 (N_48166,N_47902,N_47942);
and U48167 (N_48167,N_47732,N_47974);
xor U48168 (N_48168,N_47913,N_47569);
nor U48169 (N_48169,N_47884,N_47522);
or U48170 (N_48170,N_47589,N_47922);
and U48171 (N_48171,N_47858,N_47685);
nor U48172 (N_48172,N_47808,N_47712);
xnor U48173 (N_48173,N_47981,N_47774);
xor U48174 (N_48174,N_47566,N_47822);
and U48175 (N_48175,N_47573,N_47765);
nand U48176 (N_48176,N_47694,N_47654);
nand U48177 (N_48177,N_47915,N_47641);
or U48178 (N_48178,N_47598,N_47978);
or U48179 (N_48179,N_47724,N_47549);
nand U48180 (N_48180,N_47540,N_47548);
nand U48181 (N_48181,N_47665,N_47524);
nor U48182 (N_48182,N_47839,N_47936);
nor U48183 (N_48183,N_47813,N_47821);
or U48184 (N_48184,N_47652,N_47602);
nand U48185 (N_48185,N_47871,N_47986);
and U48186 (N_48186,N_47948,N_47699);
nor U48187 (N_48187,N_47906,N_47891);
xnor U48188 (N_48188,N_47934,N_47850);
nand U48189 (N_48189,N_47544,N_47608);
and U48190 (N_48190,N_47741,N_47711);
nand U48191 (N_48191,N_47692,N_47682);
and U48192 (N_48192,N_47538,N_47686);
and U48193 (N_48193,N_47807,N_47503);
nor U48194 (N_48194,N_47703,N_47885);
nor U48195 (N_48195,N_47852,N_47868);
and U48196 (N_48196,N_47853,N_47542);
xnor U48197 (N_48197,N_47577,N_47927);
nand U48198 (N_48198,N_47959,N_47613);
or U48199 (N_48199,N_47517,N_47881);
and U48200 (N_48200,N_47536,N_47980);
nor U48201 (N_48201,N_47989,N_47851);
nor U48202 (N_48202,N_47956,N_47725);
or U48203 (N_48203,N_47768,N_47541);
and U48204 (N_48204,N_47657,N_47911);
nand U48205 (N_48205,N_47933,N_47863);
or U48206 (N_48206,N_47622,N_47854);
nand U48207 (N_48207,N_47705,N_47528);
nor U48208 (N_48208,N_47862,N_47788);
or U48209 (N_48209,N_47678,N_47625);
nand U48210 (N_48210,N_47670,N_47796);
and U48211 (N_48211,N_47624,N_47958);
or U48212 (N_48212,N_47846,N_47738);
xor U48213 (N_48213,N_47511,N_47593);
or U48214 (N_48214,N_47969,N_47702);
nor U48215 (N_48215,N_47999,N_47976);
or U48216 (N_48216,N_47793,N_47735);
or U48217 (N_48217,N_47995,N_47603);
xor U48218 (N_48218,N_47865,N_47611);
or U48219 (N_48219,N_47676,N_47597);
and U48220 (N_48220,N_47636,N_47802);
and U48221 (N_48221,N_47634,N_47501);
nand U48222 (N_48222,N_47932,N_47681);
nor U48223 (N_48223,N_47751,N_47794);
nand U48224 (N_48224,N_47844,N_47923);
or U48225 (N_48225,N_47893,N_47716);
nand U48226 (N_48226,N_47776,N_47563);
and U48227 (N_48227,N_47695,N_47762);
nor U48228 (N_48228,N_47644,N_47575);
nor U48229 (N_48229,N_47945,N_47985);
or U48230 (N_48230,N_47806,N_47771);
nor U48231 (N_48231,N_47782,N_47717);
nor U48232 (N_48232,N_47659,N_47860);
and U48233 (N_48233,N_47708,N_47653);
and U48234 (N_48234,N_47560,N_47631);
or U48235 (N_48235,N_47671,N_47640);
or U48236 (N_48236,N_47965,N_47693);
xor U48237 (N_48237,N_47899,N_47753);
nor U48238 (N_48238,N_47748,N_47543);
nand U48239 (N_48239,N_47855,N_47518);
or U48240 (N_48240,N_47726,N_47843);
and U48241 (N_48241,N_47921,N_47555);
and U48242 (N_48242,N_47876,N_47820);
or U48243 (N_48243,N_47704,N_47856);
nor U48244 (N_48244,N_47811,N_47769);
nor U48245 (N_48245,N_47957,N_47953);
nor U48246 (N_48246,N_47963,N_47955);
nand U48247 (N_48247,N_47617,N_47742);
nor U48248 (N_48248,N_47550,N_47584);
nor U48249 (N_48249,N_47864,N_47740);
and U48250 (N_48250,N_47833,N_47587);
or U48251 (N_48251,N_47545,N_47911);
or U48252 (N_48252,N_47861,N_47606);
and U48253 (N_48253,N_47925,N_47914);
and U48254 (N_48254,N_47918,N_47966);
nand U48255 (N_48255,N_47944,N_47666);
nor U48256 (N_48256,N_47515,N_47912);
and U48257 (N_48257,N_47882,N_47962);
and U48258 (N_48258,N_47571,N_47968);
or U48259 (N_48259,N_47651,N_47701);
or U48260 (N_48260,N_47741,N_47607);
nor U48261 (N_48261,N_47789,N_47764);
nand U48262 (N_48262,N_47696,N_47885);
and U48263 (N_48263,N_47576,N_47890);
and U48264 (N_48264,N_47596,N_47805);
or U48265 (N_48265,N_47890,N_47928);
and U48266 (N_48266,N_47632,N_47828);
or U48267 (N_48267,N_47508,N_47699);
nor U48268 (N_48268,N_47731,N_47648);
xnor U48269 (N_48269,N_47761,N_47732);
and U48270 (N_48270,N_47543,N_47866);
xor U48271 (N_48271,N_47929,N_47664);
or U48272 (N_48272,N_47524,N_47523);
nand U48273 (N_48273,N_47658,N_47806);
and U48274 (N_48274,N_47916,N_47628);
nor U48275 (N_48275,N_47595,N_47581);
and U48276 (N_48276,N_47626,N_47547);
or U48277 (N_48277,N_47764,N_47993);
and U48278 (N_48278,N_47543,N_47580);
xor U48279 (N_48279,N_47576,N_47905);
nand U48280 (N_48280,N_47510,N_47785);
or U48281 (N_48281,N_47892,N_47922);
nor U48282 (N_48282,N_47989,N_47978);
or U48283 (N_48283,N_47522,N_47896);
and U48284 (N_48284,N_47670,N_47759);
nand U48285 (N_48285,N_47643,N_47611);
nor U48286 (N_48286,N_47652,N_47962);
or U48287 (N_48287,N_47949,N_47919);
nand U48288 (N_48288,N_47796,N_47557);
and U48289 (N_48289,N_47876,N_47625);
nand U48290 (N_48290,N_47972,N_47889);
nand U48291 (N_48291,N_47568,N_47561);
nor U48292 (N_48292,N_47607,N_47535);
nand U48293 (N_48293,N_47610,N_47895);
nor U48294 (N_48294,N_47867,N_47709);
or U48295 (N_48295,N_47626,N_47709);
or U48296 (N_48296,N_47983,N_47746);
or U48297 (N_48297,N_47855,N_47954);
or U48298 (N_48298,N_47791,N_47805);
and U48299 (N_48299,N_47667,N_47813);
nand U48300 (N_48300,N_47521,N_47550);
or U48301 (N_48301,N_47671,N_47827);
nand U48302 (N_48302,N_47666,N_47923);
and U48303 (N_48303,N_47837,N_47621);
nand U48304 (N_48304,N_47819,N_47632);
or U48305 (N_48305,N_47993,N_47954);
and U48306 (N_48306,N_47590,N_47796);
nor U48307 (N_48307,N_47981,N_47995);
or U48308 (N_48308,N_47517,N_47681);
nor U48309 (N_48309,N_47504,N_47627);
nor U48310 (N_48310,N_47762,N_47760);
and U48311 (N_48311,N_47591,N_47836);
nor U48312 (N_48312,N_47983,N_47669);
nor U48313 (N_48313,N_47657,N_47974);
nand U48314 (N_48314,N_47513,N_47947);
and U48315 (N_48315,N_47689,N_47690);
nand U48316 (N_48316,N_47622,N_47658);
nor U48317 (N_48317,N_47808,N_47914);
and U48318 (N_48318,N_47596,N_47684);
and U48319 (N_48319,N_47998,N_47924);
nand U48320 (N_48320,N_47692,N_47902);
nand U48321 (N_48321,N_47795,N_47664);
or U48322 (N_48322,N_47546,N_47640);
and U48323 (N_48323,N_47741,N_47680);
and U48324 (N_48324,N_47808,N_47880);
nor U48325 (N_48325,N_47771,N_47678);
nor U48326 (N_48326,N_47539,N_47898);
nor U48327 (N_48327,N_47645,N_47526);
or U48328 (N_48328,N_47818,N_47843);
xor U48329 (N_48329,N_47701,N_47829);
or U48330 (N_48330,N_47623,N_47790);
or U48331 (N_48331,N_47518,N_47960);
or U48332 (N_48332,N_47618,N_47847);
xor U48333 (N_48333,N_47565,N_47697);
nor U48334 (N_48334,N_47516,N_47799);
or U48335 (N_48335,N_47972,N_47967);
or U48336 (N_48336,N_47737,N_47963);
nor U48337 (N_48337,N_47886,N_47719);
and U48338 (N_48338,N_47628,N_47843);
nand U48339 (N_48339,N_47975,N_47922);
nor U48340 (N_48340,N_47990,N_47833);
and U48341 (N_48341,N_47902,N_47805);
or U48342 (N_48342,N_47592,N_47858);
xnor U48343 (N_48343,N_47550,N_47969);
or U48344 (N_48344,N_47926,N_47675);
nand U48345 (N_48345,N_47562,N_47657);
nor U48346 (N_48346,N_47794,N_47796);
and U48347 (N_48347,N_47699,N_47899);
nor U48348 (N_48348,N_47840,N_47830);
nor U48349 (N_48349,N_47807,N_47828);
and U48350 (N_48350,N_47841,N_47880);
and U48351 (N_48351,N_47797,N_47785);
or U48352 (N_48352,N_47892,N_47559);
and U48353 (N_48353,N_47833,N_47933);
nand U48354 (N_48354,N_47913,N_47640);
nand U48355 (N_48355,N_47792,N_47925);
nand U48356 (N_48356,N_47745,N_47545);
nor U48357 (N_48357,N_47573,N_47834);
and U48358 (N_48358,N_47581,N_47904);
nor U48359 (N_48359,N_47601,N_47870);
and U48360 (N_48360,N_47868,N_47726);
and U48361 (N_48361,N_47626,N_47944);
nand U48362 (N_48362,N_47909,N_47881);
nor U48363 (N_48363,N_47555,N_47563);
nand U48364 (N_48364,N_47834,N_47741);
nand U48365 (N_48365,N_47788,N_47604);
nor U48366 (N_48366,N_47642,N_47842);
nor U48367 (N_48367,N_47576,N_47573);
nor U48368 (N_48368,N_47963,N_47992);
and U48369 (N_48369,N_47826,N_47741);
nor U48370 (N_48370,N_47569,N_47559);
and U48371 (N_48371,N_47892,N_47709);
nor U48372 (N_48372,N_47910,N_47653);
xnor U48373 (N_48373,N_47716,N_47991);
nand U48374 (N_48374,N_47794,N_47840);
nand U48375 (N_48375,N_47873,N_47586);
or U48376 (N_48376,N_47744,N_47684);
or U48377 (N_48377,N_47660,N_47959);
or U48378 (N_48378,N_47645,N_47792);
nor U48379 (N_48379,N_47729,N_47883);
and U48380 (N_48380,N_47608,N_47859);
or U48381 (N_48381,N_47693,N_47964);
or U48382 (N_48382,N_47587,N_47604);
or U48383 (N_48383,N_47631,N_47585);
and U48384 (N_48384,N_47804,N_47641);
nor U48385 (N_48385,N_47757,N_47690);
nand U48386 (N_48386,N_47566,N_47577);
xnor U48387 (N_48387,N_47857,N_47804);
or U48388 (N_48388,N_47752,N_47619);
and U48389 (N_48389,N_47837,N_47582);
or U48390 (N_48390,N_47556,N_47923);
or U48391 (N_48391,N_47606,N_47654);
or U48392 (N_48392,N_47931,N_47880);
nor U48393 (N_48393,N_47578,N_47652);
nand U48394 (N_48394,N_47772,N_47688);
nand U48395 (N_48395,N_47617,N_47894);
or U48396 (N_48396,N_47649,N_47845);
xnor U48397 (N_48397,N_47684,N_47565);
or U48398 (N_48398,N_47560,N_47810);
xor U48399 (N_48399,N_47821,N_47770);
or U48400 (N_48400,N_47701,N_47723);
nor U48401 (N_48401,N_47703,N_47591);
or U48402 (N_48402,N_47530,N_47791);
nand U48403 (N_48403,N_47691,N_47543);
nor U48404 (N_48404,N_47852,N_47914);
and U48405 (N_48405,N_47852,N_47675);
nand U48406 (N_48406,N_47731,N_47756);
nand U48407 (N_48407,N_47700,N_47944);
and U48408 (N_48408,N_47574,N_47955);
nand U48409 (N_48409,N_47790,N_47943);
nor U48410 (N_48410,N_47567,N_47729);
and U48411 (N_48411,N_47505,N_47633);
nand U48412 (N_48412,N_47638,N_47754);
nand U48413 (N_48413,N_47737,N_47637);
nand U48414 (N_48414,N_47551,N_47818);
nand U48415 (N_48415,N_47566,N_47667);
nor U48416 (N_48416,N_47713,N_47677);
or U48417 (N_48417,N_47833,N_47541);
and U48418 (N_48418,N_47871,N_47654);
nor U48419 (N_48419,N_47999,N_47595);
or U48420 (N_48420,N_47771,N_47819);
or U48421 (N_48421,N_47596,N_47825);
or U48422 (N_48422,N_47727,N_47802);
nand U48423 (N_48423,N_47960,N_47525);
and U48424 (N_48424,N_47508,N_47501);
and U48425 (N_48425,N_47871,N_47591);
nor U48426 (N_48426,N_47972,N_47916);
or U48427 (N_48427,N_47953,N_47571);
nand U48428 (N_48428,N_47812,N_47637);
nor U48429 (N_48429,N_47540,N_47920);
and U48430 (N_48430,N_47967,N_47875);
xnor U48431 (N_48431,N_47897,N_47672);
nor U48432 (N_48432,N_47647,N_47954);
and U48433 (N_48433,N_47588,N_47623);
or U48434 (N_48434,N_47741,N_47800);
xnor U48435 (N_48435,N_47626,N_47605);
or U48436 (N_48436,N_47785,N_47608);
nand U48437 (N_48437,N_47845,N_47529);
and U48438 (N_48438,N_47712,N_47661);
nor U48439 (N_48439,N_47757,N_47730);
or U48440 (N_48440,N_47875,N_47807);
nand U48441 (N_48441,N_47563,N_47796);
and U48442 (N_48442,N_47515,N_47634);
and U48443 (N_48443,N_47888,N_47928);
nor U48444 (N_48444,N_47663,N_47964);
nand U48445 (N_48445,N_47853,N_47846);
and U48446 (N_48446,N_47801,N_47906);
nand U48447 (N_48447,N_47914,N_47985);
and U48448 (N_48448,N_47625,N_47825);
nor U48449 (N_48449,N_47870,N_47677);
nand U48450 (N_48450,N_47972,N_47942);
nand U48451 (N_48451,N_47847,N_47922);
and U48452 (N_48452,N_47834,N_47677);
or U48453 (N_48453,N_47909,N_47753);
or U48454 (N_48454,N_47697,N_47788);
and U48455 (N_48455,N_47628,N_47768);
and U48456 (N_48456,N_47575,N_47563);
or U48457 (N_48457,N_47621,N_47722);
and U48458 (N_48458,N_47741,N_47876);
nand U48459 (N_48459,N_47939,N_47711);
and U48460 (N_48460,N_47936,N_47808);
xnor U48461 (N_48461,N_47963,N_47886);
nand U48462 (N_48462,N_47839,N_47617);
or U48463 (N_48463,N_47590,N_47611);
and U48464 (N_48464,N_47542,N_47812);
or U48465 (N_48465,N_47637,N_47991);
nor U48466 (N_48466,N_47559,N_47804);
nand U48467 (N_48467,N_47628,N_47862);
nor U48468 (N_48468,N_47896,N_47610);
nand U48469 (N_48469,N_47954,N_47668);
nand U48470 (N_48470,N_47893,N_47534);
or U48471 (N_48471,N_47771,N_47561);
xor U48472 (N_48472,N_47684,N_47865);
and U48473 (N_48473,N_47727,N_47753);
and U48474 (N_48474,N_47856,N_47759);
nand U48475 (N_48475,N_47726,N_47526);
nor U48476 (N_48476,N_47544,N_47836);
and U48477 (N_48477,N_47702,N_47572);
nor U48478 (N_48478,N_47976,N_47751);
and U48479 (N_48479,N_47969,N_47576);
and U48480 (N_48480,N_47987,N_47588);
nor U48481 (N_48481,N_47529,N_47615);
nand U48482 (N_48482,N_47697,N_47679);
nand U48483 (N_48483,N_47575,N_47519);
or U48484 (N_48484,N_47781,N_47556);
xor U48485 (N_48485,N_47785,N_47942);
nand U48486 (N_48486,N_47649,N_47689);
or U48487 (N_48487,N_47577,N_47537);
nand U48488 (N_48488,N_47977,N_47675);
xnor U48489 (N_48489,N_47707,N_47802);
and U48490 (N_48490,N_47695,N_47717);
nand U48491 (N_48491,N_47565,N_47701);
and U48492 (N_48492,N_47670,N_47669);
and U48493 (N_48493,N_47661,N_47801);
nand U48494 (N_48494,N_47909,N_47951);
nor U48495 (N_48495,N_47670,N_47813);
or U48496 (N_48496,N_47991,N_47937);
nor U48497 (N_48497,N_47998,N_47832);
and U48498 (N_48498,N_47644,N_47611);
and U48499 (N_48499,N_47885,N_47746);
or U48500 (N_48500,N_48169,N_48363);
nor U48501 (N_48501,N_48215,N_48037);
or U48502 (N_48502,N_48456,N_48444);
nand U48503 (N_48503,N_48297,N_48217);
and U48504 (N_48504,N_48030,N_48402);
nand U48505 (N_48505,N_48151,N_48435);
nor U48506 (N_48506,N_48290,N_48374);
and U48507 (N_48507,N_48276,N_48117);
nor U48508 (N_48508,N_48116,N_48181);
or U48509 (N_48509,N_48162,N_48430);
nor U48510 (N_48510,N_48343,N_48112);
or U48511 (N_48511,N_48106,N_48242);
nor U48512 (N_48512,N_48475,N_48462);
and U48513 (N_48513,N_48328,N_48197);
and U48514 (N_48514,N_48043,N_48263);
nand U48515 (N_48515,N_48377,N_48452);
nor U48516 (N_48516,N_48153,N_48454);
and U48517 (N_48517,N_48257,N_48023);
xor U48518 (N_48518,N_48413,N_48400);
nand U48519 (N_48519,N_48029,N_48253);
and U48520 (N_48520,N_48451,N_48237);
xor U48521 (N_48521,N_48414,N_48418);
and U48522 (N_48522,N_48318,N_48099);
or U48523 (N_48523,N_48009,N_48333);
and U48524 (N_48524,N_48062,N_48348);
or U48525 (N_48525,N_48330,N_48178);
or U48526 (N_48526,N_48235,N_48026);
nand U48527 (N_48527,N_48423,N_48130);
and U48528 (N_48528,N_48119,N_48264);
nand U48529 (N_48529,N_48344,N_48381);
xor U48530 (N_48530,N_48221,N_48284);
and U48531 (N_48531,N_48079,N_48110);
nor U48532 (N_48532,N_48187,N_48408);
or U48533 (N_48533,N_48411,N_48025);
nor U48534 (N_48534,N_48380,N_48142);
nor U48535 (N_48535,N_48273,N_48222);
and U48536 (N_48536,N_48440,N_48319);
and U48537 (N_48537,N_48450,N_48096);
and U48538 (N_48538,N_48189,N_48464);
and U48539 (N_48539,N_48275,N_48077);
nor U48540 (N_48540,N_48059,N_48072);
nor U48541 (N_48541,N_48383,N_48461);
xor U48542 (N_48542,N_48240,N_48457);
nand U48543 (N_48543,N_48011,N_48499);
and U48544 (N_48544,N_48442,N_48172);
and U48545 (N_48545,N_48047,N_48213);
and U48546 (N_48546,N_48075,N_48107);
nand U48547 (N_48547,N_48313,N_48299);
and U48548 (N_48548,N_48433,N_48326);
nand U48549 (N_48549,N_48448,N_48366);
nor U48550 (N_48550,N_48355,N_48340);
or U48551 (N_48551,N_48122,N_48298);
nor U48552 (N_48552,N_48485,N_48310);
nor U48553 (N_48553,N_48155,N_48102);
xnor U48554 (N_48554,N_48300,N_48397);
and U48555 (N_48555,N_48312,N_48125);
xor U48556 (N_48556,N_48458,N_48289);
nand U48557 (N_48557,N_48426,N_48252);
or U48558 (N_48558,N_48233,N_48286);
and U48559 (N_48559,N_48419,N_48295);
and U48560 (N_48560,N_48357,N_48164);
and U48561 (N_48561,N_48323,N_48111);
nor U48562 (N_48562,N_48376,N_48018);
xnor U48563 (N_48563,N_48347,N_48439);
xor U48564 (N_48564,N_48453,N_48051);
and U48565 (N_48565,N_48209,N_48204);
or U48566 (N_48566,N_48086,N_48385);
nand U48567 (N_48567,N_48294,N_48128);
nand U48568 (N_48568,N_48049,N_48466);
nor U48569 (N_48569,N_48489,N_48285);
nor U48570 (N_48570,N_48195,N_48492);
nor U48571 (N_48571,N_48250,N_48185);
nor U48572 (N_48572,N_48027,N_48415);
nand U48573 (N_48573,N_48177,N_48341);
nor U48574 (N_48574,N_48071,N_48021);
nand U48575 (N_48575,N_48490,N_48005);
or U48576 (N_48576,N_48254,N_48293);
and U48577 (N_48577,N_48024,N_48074);
nor U48578 (N_48578,N_48068,N_48272);
and U48579 (N_48579,N_48126,N_48244);
xor U48580 (N_48580,N_48156,N_48329);
or U48581 (N_48581,N_48225,N_48494);
and U48582 (N_48582,N_48139,N_48095);
or U48583 (N_48583,N_48283,N_48199);
nand U48584 (N_48584,N_48212,N_48054);
nor U48585 (N_48585,N_48133,N_48045);
or U48586 (N_48586,N_48032,N_48201);
nand U48587 (N_48587,N_48168,N_48473);
and U48588 (N_48588,N_48417,N_48281);
xnor U48589 (N_48589,N_48144,N_48196);
xor U48590 (N_48590,N_48375,N_48065);
or U48591 (N_48591,N_48121,N_48279);
xnor U48592 (N_48592,N_48371,N_48069);
or U48593 (N_48593,N_48152,N_48131);
or U48594 (N_48594,N_48409,N_48339);
nor U48595 (N_48595,N_48113,N_48484);
or U48596 (N_48596,N_48114,N_48472);
xor U48597 (N_48597,N_48309,N_48039);
nand U48598 (N_48598,N_48488,N_48470);
nor U48599 (N_48599,N_48124,N_48186);
nor U48600 (N_48600,N_48365,N_48447);
or U48601 (N_48601,N_48307,N_48245);
nor U48602 (N_48602,N_48493,N_48007);
nand U48603 (N_48603,N_48277,N_48287);
or U48604 (N_48604,N_48033,N_48481);
and U48605 (N_48605,N_48350,N_48308);
and U48606 (N_48606,N_48266,N_48120);
or U48607 (N_48607,N_48478,N_48282);
and U48608 (N_48608,N_48449,N_48459);
nor U48609 (N_48609,N_48429,N_48268);
xor U48610 (N_48610,N_48378,N_48424);
or U48611 (N_48611,N_48425,N_48081);
and U48612 (N_48612,N_48150,N_48082);
nand U48613 (N_48613,N_48104,N_48249);
nand U48614 (N_48614,N_48042,N_48198);
nor U48615 (N_48615,N_48392,N_48191);
nand U48616 (N_48616,N_48076,N_48256);
or U48617 (N_48617,N_48336,N_48428);
and U48618 (N_48618,N_48384,N_48161);
or U48619 (N_48619,N_48231,N_48483);
nor U48620 (N_48620,N_48006,N_48353);
xnor U48621 (N_48621,N_48265,N_48141);
nand U48622 (N_48622,N_48427,N_48214);
xnor U48623 (N_48623,N_48239,N_48302);
or U48624 (N_48624,N_48108,N_48261);
and U48625 (N_48625,N_48129,N_48008);
or U48626 (N_48626,N_48498,N_48248);
and U48627 (N_48627,N_48432,N_48109);
or U48628 (N_48628,N_48057,N_48325);
nor U48629 (N_48629,N_48190,N_48480);
or U48630 (N_48630,N_48159,N_48438);
nand U48631 (N_48631,N_48016,N_48017);
or U48632 (N_48632,N_48145,N_48013);
nand U48633 (N_48633,N_48183,N_48166);
nand U48634 (N_48634,N_48398,N_48140);
nand U48635 (N_48635,N_48404,N_48137);
nand U48636 (N_48636,N_48000,N_48474);
nand U48637 (N_48637,N_48089,N_48291);
or U48638 (N_48638,N_48223,N_48497);
and U48639 (N_48639,N_48094,N_48200);
and U48640 (N_48640,N_48251,N_48052);
and U48641 (N_48641,N_48446,N_48314);
nand U48642 (N_48642,N_48046,N_48136);
and U48643 (N_48643,N_48403,N_48331);
nand U48644 (N_48644,N_48028,N_48192);
or U48645 (N_48645,N_48345,N_48334);
nor U48646 (N_48646,N_48203,N_48078);
nor U48647 (N_48647,N_48002,N_48361);
or U48648 (N_48648,N_48154,N_48445);
or U48649 (N_48649,N_48210,N_48389);
nand U48650 (N_48650,N_48218,N_48486);
nand U48651 (N_48651,N_48247,N_48055);
and U48652 (N_48652,N_48170,N_48066);
nand U48653 (N_48653,N_48269,N_48394);
and U48654 (N_48654,N_48320,N_48422);
nor U48655 (N_48655,N_48146,N_48360);
and U48656 (N_48656,N_48138,N_48056);
and U48657 (N_48657,N_48160,N_48471);
xnor U48658 (N_48658,N_48048,N_48399);
and U48659 (N_48659,N_48227,N_48167);
nor U48660 (N_48660,N_48182,N_48158);
nor U48661 (N_48661,N_48338,N_48479);
nand U48662 (N_48662,N_48332,N_48349);
or U48663 (N_48663,N_48238,N_48220);
nor U48664 (N_48664,N_48356,N_48020);
or U48665 (N_48665,N_48469,N_48219);
and U48666 (N_48666,N_48091,N_48386);
xnor U48667 (N_48667,N_48004,N_48335);
and U48668 (N_48668,N_48070,N_48436);
nand U48669 (N_48669,N_48019,N_48093);
or U48670 (N_48670,N_48373,N_48393);
nor U48671 (N_48671,N_48379,N_48229);
and U48672 (N_48672,N_48487,N_48034);
and U48673 (N_48673,N_48080,N_48206);
nand U48674 (N_48674,N_48064,N_48270);
nand U48675 (N_48675,N_48262,N_48135);
nor U48676 (N_48676,N_48001,N_48097);
nor U48677 (N_48677,N_48387,N_48053);
nand U48678 (N_48678,N_48304,N_48255);
xor U48679 (N_48679,N_48084,N_48370);
and U48680 (N_48680,N_48038,N_48036);
and U48681 (N_48681,N_48098,N_48259);
nor U48682 (N_48682,N_48022,N_48143);
and U48683 (N_48683,N_48073,N_48207);
nor U48684 (N_48684,N_48342,N_48316);
nand U48685 (N_48685,N_48226,N_48202);
nor U48686 (N_48686,N_48437,N_48205);
or U48687 (N_48687,N_48224,N_48115);
and U48688 (N_48688,N_48063,N_48044);
or U48689 (N_48689,N_48067,N_48321);
or U48690 (N_48690,N_48118,N_48061);
nor U48691 (N_48691,N_48179,N_48431);
nor U48692 (N_48692,N_48088,N_48406);
or U48693 (N_48693,N_48232,N_48463);
or U48694 (N_48694,N_48467,N_48041);
xor U48695 (N_48695,N_48100,N_48010);
or U48696 (N_48696,N_48176,N_48003);
and U48697 (N_48697,N_48180,N_48317);
nor U48698 (N_48698,N_48230,N_48496);
or U48699 (N_48699,N_48271,N_48157);
or U48700 (N_48700,N_48040,N_48188);
xnor U48701 (N_48701,N_48364,N_48491);
and U48702 (N_48702,N_48274,N_48288);
nand U48703 (N_48703,N_48482,N_48184);
nor U48704 (N_48704,N_48258,N_48083);
nor U48705 (N_48705,N_48301,N_48085);
nor U48706 (N_48706,N_48337,N_48455);
nand U48707 (N_48707,N_48148,N_48015);
nor U48708 (N_48708,N_48292,N_48372);
nor U48709 (N_48709,N_48346,N_48127);
nand U48710 (N_48710,N_48246,N_48228);
nand U48711 (N_48711,N_48477,N_48367);
and U48712 (N_48712,N_48211,N_48407);
nand U48713 (N_48713,N_48171,N_48322);
or U48714 (N_48714,N_48165,N_48443);
and U48715 (N_48715,N_48410,N_48058);
and U48716 (N_48716,N_48362,N_48175);
or U48717 (N_48717,N_48090,N_48382);
nand U48718 (N_48718,N_48311,N_48050);
xnor U48719 (N_48719,N_48354,N_48193);
nand U48720 (N_48720,N_48267,N_48306);
nand U48721 (N_48721,N_48234,N_48087);
nor U48722 (N_48722,N_48105,N_48278);
nand U48723 (N_48723,N_48420,N_48012);
xnor U48724 (N_48724,N_48351,N_48315);
nor U48725 (N_48725,N_48147,N_48412);
xnor U48726 (N_48726,N_48236,N_48123);
nand U48727 (N_48727,N_48305,N_48369);
xor U48728 (N_48728,N_48173,N_48103);
nor U48729 (N_48729,N_48391,N_48243);
nor U48730 (N_48730,N_48401,N_48390);
and U48731 (N_48731,N_48303,N_48416);
or U48732 (N_48732,N_48208,N_48421);
or U48733 (N_48733,N_48101,N_48260);
or U48734 (N_48734,N_48352,N_48241);
nand U48735 (N_48735,N_48327,N_48134);
or U48736 (N_48736,N_48296,N_48194);
nand U48737 (N_48737,N_48359,N_48368);
nor U48738 (N_48738,N_48476,N_48149);
or U48739 (N_48739,N_48163,N_48441);
and U48740 (N_48740,N_48280,N_48035);
nand U48741 (N_48741,N_48460,N_48014);
nand U48742 (N_48742,N_48324,N_48465);
nand U48743 (N_48743,N_48031,N_48388);
and U48744 (N_48744,N_48132,N_48060);
xor U48745 (N_48745,N_48358,N_48495);
nand U48746 (N_48746,N_48216,N_48092);
nand U48747 (N_48747,N_48405,N_48174);
and U48748 (N_48748,N_48396,N_48434);
xnor U48749 (N_48749,N_48468,N_48395);
nand U48750 (N_48750,N_48243,N_48354);
and U48751 (N_48751,N_48394,N_48005);
nor U48752 (N_48752,N_48093,N_48172);
and U48753 (N_48753,N_48435,N_48062);
xor U48754 (N_48754,N_48238,N_48367);
nor U48755 (N_48755,N_48022,N_48383);
nand U48756 (N_48756,N_48261,N_48026);
and U48757 (N_48757,N_48010,N_48495);
nor U48758 (N_48758,N_48072,N_48447);
xor U48759 (N_48759,N_48365,N_48198);
or U48760 (N_48760,N_48013,N_48093);
and U48761 (N_48761,N_48065,N_48285);
nand U48762 (N_48762,N_48191,N_48391);
and U48763 (N_48763,N_48094,N_48321);
or U48764 (N_48764,N_48207,N_48087);
and U48765 (N_48765,N_48115,N_48088);
nor U48766 (N_48766,N_48131,N_48085);
or U48767 (N_48767,N_48466,N_48434);
nand U48768 (N_48768,N_48270,N_48235);
xor U48769 (N_48769,N_48059,N_48050);
or U48770 (N_48770,N_48321,N_48464);
nand U48771 (N_48771,N_48173,N_48281);
or U48772 (N_48772,N_48419,N_48266);
or U48773 (N_48773,N_48193,N_48248);
nor U48774 (N_48774,N_48294,N_48298);
xnor U48775 (N_48775,N_48371,N_48325);
and U48776 (N_48776,N_48276,N_48253);
xor U48777 (N_48777,N_48490,N_48353);
and U48778 (N_48778,N_48261,N_48080);
or U48779 (N_48779,N_48168,N_48494);
and U48780 (N_48780,N_48409,N_48288);
nor U48781 (N_48781,N_48093,N_48125);
or U48782 (N_48782,N_48125,N_48077);
nor U48783 (N_48783,N_48434,N_48433);
nand U48784 (N_48784,N_48486,N_48411);
and U48785 (N_48785,N_48246,N_48069);
nor U48786 (N_48786,N_48386,N_48220);
and U48787 (N_48787,N_48177,N_48381);
and U48788 (N_48788,N_48131,N_48490);
nor U48789 (N_48789,N_48017,N_48477);
and U48790 (N_48790,N_48454,N_48486);
and U48791 (N_48791,N_48048,N_48320);
or U48792 (N_48792,N_48068,N_48368);
or U48793 (N_48793,N_48344,N_48112);
nor U48794 (N_48794,N_48280,N_48428);
xnor U48795 (N_48795,N_48118,N_48169);
and U48796 (N_48796,N_48367,N_48033);
and U48797 (N_48797,N_48370,N_48218);
or U48798 (N_48798,N_48232,N_48171);
or U48799 (N_48799,N_48260,N_48312);
nor U48800 (N_48800,N_48453,N_48036);
nand U48801 (N_48801,N_48380,N_48426);
and U48802 (N_48802,N_48421,N_48001);
or U48803 (N_48803,N_48435,N_48382);
nor U48804 (N_48804,N_48375,N_48293);
and U48805 (N_48805,N_48330,N_48357);
nand U48806 (N_48806,N_48067,N_48363);
nand U48807 (N_48807,N_48019,N_48314);
xor U48808 (N_48808,N_48194,N_48285);
nand U48809 (N_48809,N_48405,N_48298);
nor U48810 (N_48810,N_48409,N_48255);
xor U48811 (N_48811,N_48060,N_48133);
nand U48812 (N_48812,N_48138,N_48249);
nor U48813 (N_48813,N_48002,N_48090);
nand U48814 (N_48814,N_48097,N_48370);
nand U48815 (N_48815,N_48185,N_48019);
or U48816 (N_48816,N_48293,N_48486);
xnor U48817 (N_48817,N_48380,N_48027);
and U48818 (N_48818,N_48157,N_48420);
and U48819 (N_48819,N_48200,N_48301);
nor U48820 (N_48820,N_48214,N_48185);
nor U48821 (N_48821,N_48397,N_48416);
nor U48822 (N_48822,N_48011,N_48250);
nand U48823 (N_48823,N_48062,N_48491);
or U48824 (N_48824,N_48219,N_48360);
xnor U48825 (N_48825,N_48167,N_48317);
nor U48826 (N_48826,N_48174,N_48454);
nor U48827 (N_48827,N_48355,N_48488);
nand U48828 (N_48828,N_48138,N_48488);
nand U48829 (N_48829,N_48296,N_48013);
xnor U48830 (N_48830,N_48330,N_48070);
and U48831 (N_48831,N_48064,N_48170);
nor U48832 (N_48832,N_48246,N_48371);
xnor U48833 (N_48833,N_48223,N_48409);
or U48834 (N_48834,N_48034,N_48361);
or U48835 (N_48835,N_48250,N_48245);
and U48836 (N_48836,N_48086,N_48115);
and U48837 (N_48837,N_48201,N_48452);
nand U48838 (N_48838,N_48326,N_48217);
nand U48839 (N_48839,N_48498,N_48087);
and U48840 (N_48840,N_48423,N_48194);
and U48841 (N_48841,N_48057,N_48250);
nand U48842 (N_48842,N_48278,N_48392);
nor U48843 (N_48843,N_48302,N_48159);
nor U48844 (N_48844,N_48270,N_48182);
nor U48845 (N_48845,N_48369,N_48342);
or U48846 (N_48846,N_48312,N_48100);
or U48847 (N_48847,N_48411,N_48321);
nand U48848 (N_48848,N_48344,N_48353);
nand U48849 (N_48849,N_48445,N_48055);
and U48850 (N_48850,N_48169,N_48347);
and U48851 (N_48851,N_48235,N_48283);
nand U48852 (N_48852,N_48161,N_48463);
nand U48853 (N_48853,N_48143,N_48209);
nand U48854 (N_48854,N_48076,N_48038);
and U48855 (N_48855,N_48364,N_48211);
nor U48856 (N_48856,N_48022,N_48196);
nor U48857 (N_48857,N_48349,N_48382);
nand U48858 (N_48858,N_48001,N_48122);
nand U48859 (N_48859,N_48340,N_48305);
nand U48860 (N_48860,N_48326,N_48233);
or U48861 (N_48861,N_48487,N_48348);
nand U48862 (N_48862,N_48445,N_48157);
and U48863 (N_48863,N_48014,N_48183);
nand U48864 (N_48864,N_48341,N_48466);
and U48865 (N_48865,N_48446,N_48062);
nor U48866 (N_48866,N_48314,N_48107);
nor U48867 (N_48867,N_48478,N_48393);
nand U48868 (N_48868,N_48250,N_48397);
nor U48869 (N_48869,N_48006,N_48296);
and U48870 (N_48870,N_48217,N_48335);
nor U48871 (N_48871,N_48381,N_48308);
nor U48872 (N_48872,N_48323,N_48097);
and U48873 (N_48873,N_48428,N_48465);
nand U48874 (N_48874,N_48351,N_48167);
nor U48875 (N_48875,N_48244,N_48488);
nor U48876 (N_48876,N_48125,N_48232);
xnor U48877 (N_48877,N_48270,N_48152);
xor U48878 (N_48878,N_48247,N_48410);
nor U48879 (N_48879,N_48245,N_48093);
nand U48880 (N_48880,N_48120,N_48006);
xnor U48881 (N_48881,N_48154,N_48129);
xor U48882 (N_48882,N_48150,N_48046);
nor U48883 (N_48883,N_48191,N_48040);
and U48884 (N_48884,N_48300,N_48147);
or U48885 (N_48885,N_48086,N_48059);
nand U48886 (N_48886,N_48107,N_48025);
xnor U48887 (N_48887,N_48116,N_48255);
or U48888 (N_48888,N_48173,N_48019);
nand U48889 (N_48889,N_48269,N_48238);
or U48890 (N_48890,N_48291,N_48467);
nand U48891 (N_48891,N_48372,N_48329);
and U48892 (N_48892,N_48089,N_48230);
nand U48893 (N_48893,N_48022,N_48329);
xor U48894 (N_48894,N_48432,N_48441);
nand U48895 (N_48895,N_48221,N_48323);
or U48896 (N_48896,N_48382,N_48136);
or U48897 (N_48897,N_48176,N_48164);
or U48898 (N_48898,N_48472,N_48143);
xnor U48899 (N_48899,N_48186,N_48119);
and U48900 (N_48900,N_48287,N_48062);
nor U48901 (N_48901,N_48192,N_48376);
or U48902 (N_48902,N_48496,N_48319);
and U48903 (N_48903,N_48179,N_48261);
nor U48904 (N_48904,N_48016,N_48169);
nand U48905 (N_48905,N_48310,N_48074);
nor U48906 (N_48906,N_48490,N_48480);
and U48907 (N_48907,N_48456,N_48472);
or U48908 (N_48908,N_48055,N_48341);
nor U48909 (N_48909,N_48421,N_48278);
and U48910 (N_48910,N_48464,N_48128);
xor U48911 (N_48911,N_48055,N_48175);
xnor U48912 (N_48912,N_48092,N_48263);
or U48913 (N_48913,N_48014,N_48389);
and U48914 (N_48914,N_48315,N_48020);
xor U48915 (N_48915,N_48165,N_48416);
and U48916 (N_48916,N_48422,N_48082);
nor U48917 (N_48917,N_48076,N_48393);
or U48918 (N_48918,N_48450,N_48433);
nor U48919 (N_48919,N_48439,N_48370);
or U48920 (N_48920,N_48129,N_48143);
and U48921 (N_48921,N_48088,N_48423);
and U48922 (N_48922,N_48267,N_48110);
nand U48923 (N_48923,N_48343,N_48017);
and U48924 (N_48924,N_48040,N_48472);
or U48925 (N_48925,N_48046,N_48182);
nand U48926 (N_48926,N_48005,N_48245);
or U48927 (N_48927,N_48019,N_48311);
xor U48928 (N_48928,N_48343,N_48051);
and U48929 (N_48929,N_48210,N_48067);
xnor U48930 (N_48930,N_48382,N_48301);
nor U48931 (N_48931,N_48005,N_48195);
nand U48932 (N_48932,N_48112,N_48020);
and U48933 (N_48933,N_48379,N_48303);
and U48934 (N_48934,N_48457,N_48306);
and U48935 (N_48935,N_48243,N_48480);
or U48936 (N_48936,N_48237,N_48481);
or U48937 (N_48937,N_48371,N_48472);
nor U48938 (N_48938,N_48162,N_48403);
nor U48939 (N_48939,N_48067,N_48270);
nor U48940 (N_48940,N_48211,N_48068);
xor U48941 (N_48941,N_48117,N_48082);
nor U48942 (N_48942,N_48207,N_48169);
nor U48943 (N_48943,N_48240,N_48287);
nor U48944 (N_48944,N_48382,N_48388);
nand U48945 (N_48945,N_48000,N_48006);
and U48946 (N_48946,N_48437,N_48365);
and U48947 (N_48947,N_48098,N_48315);
nor U48948 (N_48948,N_48393,N_48286);
and U48949 (N_48949,N_48289,N_48408);
nand U48950 (N_48950,N_48268,N_48386);
nand U48951 (N_48951,N_48403,N_48110);
nor U48952 (N_48952,N_48290,N_48134);
nand U48953 (N_48953,N_48321,N_48049);
or U48954 (N_48954,N_48439,N_48048);
nor U48955 (N_48955,N_48135,N_48454);
nor U48956 (N_48956,N_48333,N_48102);
or U48957 (N_48957,N_48401,N_48358);
nor U48958 (N_48958,N_48495,N_48180);
and U48959 (N_48959,N_48214,N_48365);
or U48960 (N_48960,N_48201,N_48017);
or U48961 (N_48961,N_48443,N_48293);
nand U48962 (N_48962,N_48257,N_48042);
nand U48963 (N_48963,N_48387,N_48289);
or U48964 (N_48964,N_48328,N_48103);
xor U48965 (N_48965,N_48462,N_48081);
xnor U48966 (N_48966,N_48078,N_48371);
nor U48967 (N_48967,N_48306,N_48358);
nor U48968 (N_48968,N_48400,N_48184);
nand U48969 (N_48969,N_48018,N_48081);
nor U48970 (N_48970,N_48241,N_48465);
nand U48971 (N_48971,N_48489,N_48335);
and U48972 (N_48972,N_48236,N_48208);
or U48973 (N_48973,N_48244,N_48054);
nand U48974 (N_48974,N_48483,N_48005);
and U48975 (N_48975,N_48419,N_48490);
and U48976 (N_48976,N_48345,N_48365);
or U48977 (N_48977,N_48340,N_48326);
nand U48978 (N_48978,N_48454,N_48151);
nand U48979 (N_48979,N_48385,N_48129);
or U48980 (N_48980,N_48332,N_48494);
or U48981 (N_48981,N_48461,N_48497);
nand U48982 (N_48982,N_48128,N_48330);
nand U48983 (N_48983,N_48278,N_48405);
nor U48984 (N_48984,N_48429,N_48423);
or U48985 (N_48985,N_48156,N_48185);
or U48986 (N_48986,N_48108,N_48366);
nor U48987 (N_48987,N_48206,N_48115);
nand U48988 (N_48988,N_48134,N_48219);
nand U48989 (N_48989,N_48144,N_48316);
nor U48990 (N_48990,N_48221,N_48349);
nand U48991 (N_48991,N_48045,N_48277);
nor U48992 (N_48992,N_48237,N_48068);
nand U48993 (N_48993,N_48436,N_48215);
nand U48994 (N_48994,N_48192,N_48328);
or U48995 (N_48995,N_48134,N_48008);
or U48996 (N_48996,N_48436,N_48261);
nor U48997 (N_48997,N_48160,N_48240);
nor U48998 (N_48998,N_48116,N_48426);
and U48999 (N_48999,N_48419,N_48379);
xor U49000 (N_49000,N_48675,N_48876);
nor U49001 (N_49001,N_48757,N_48955);
nand U49002 (N_49002,N_48559,N_48682);
or U49003 (N_49003,N_48859,N_48670);
nand U49004 (N_49004,N_48945,N_48927);
and U49005 (N_49005,N_48525,N_48771);
xor U49006 (N_49006,N_48936,N_48884);
nor U49007 (N_49007,N_48779,N_48941);
or U49008 (N_49008,N_48838,N_48685);
nand U49009 (N_49009,N_48904,N_48697);
nor U49010 (N_49010,N_48960,N_48813);
or U49011 (N_49011,N_48580,N_48714);
and U49012 (N_49012,N_48734,N_48750);
nor U49013 (N_49013,N_48817,N_48637);
and U49014 (N_49014,N_48988,N_48998);
and U49015 (N_49015,N_48668,N_48792);
nor U49016 (N_49016,N_48852,N_48585);
or U49017 (N_49017,N_48641,N_48732);
nand U49018 (N_49018,N_48934,N_48550);
nand U49019 (N_49019,N_48969,N_48623);
and U49020 (N_49020,N_48849,N_48797);
nand U49021 (N_49021,N_48747,N_48579);
or U49022 (N_49022,N_48723,N_48707);
and U49023 (N_49023,N_48776,N_48592);
and U49024 (N_49024,N_48693,N_48967);
nor U49025 (N_49025,N_48501,N_48522);
and U49026 (N_49026,N_48658,N_48773);
xor U49027 (N_49027,N_48566,N_48701);
nand U49028 (N_49028,N_48725,N_48547);
xnor U49029 (N_49029,N_48573,N_48749);
nor U49030 (N_49030,N_48694,N_48890);
nand U49031 (N_49031,N_48856,N_48843);
or U49032 (N_49032,N_48931,N_48917);
nor U49033 (N_49033,N_48735,N_48646);
nor U49034 (N_49034,N_48978,N_48982);
and U49035 (N_49035,N_48791,N_48558);
nor U49036 (N_49036,N_48502,N_48834);
nor U49037 (N_49037,N_48516,N_48989);
xor U49038 (N_49038,N_48795,N_48906);
nand U49039 (N_49039,N_48862,N_48690);
nand U49040 (N_49040,N_48833,N_48878);
nor U49041 (N_49041,N_48542,N_48663);
xnor U49042 (N_49042,N_48865,N_48796);
nor U49043 (N_49043,N_48899,N_48526);
or U49044 (N_49044,N_48587,N_48742);
and U49045 (N_49045,N_48786,N_48996);
nor U49046 (N_49046,N_48745,N_48816);
and U49047 (N_49047,N_48778,N_48640);
and U49048 (N_49048,N_48660,N_48861);
nand U49049 (N_49049,N_48973,N_48851);
nor U49050 (N_49050,N_48507,N_48942);
or U49051 (N_49051,N_48599,N_48958);
xnor U49052 (N_49052,N_48536,N_48828);
nor U49053 (N_49053,N_48667,N_48777);
or U49054 (N_49054,N_48544,N_48897);
nor U49055 (N_49055,N_48709,N_48823);
or U49056 (N_49056,N_48885,N_48543);
xor U49057 (N_49057,N_48681,N_48821);
nor U49058 (N_49058,N_48606,N_48551);
or U49059 (N_49059,N_48560,N_48972);
and U49060 (N_49060,N_48744,N_48647);
and U49061 (N_49061,N_48586,N_48625);
and U49062 (N_49062,N_48844,N_48620);
nor U49063 (N_49063,N_48517,N_48824);
and U49064 (N_49064,N_48617,N_48503);
and U49065 (N_49065,N_48621,N_48649);
or U49066 (N_49066,N_48918,N_48879);
or U49067 (N_49067,N_48948,N_48807);
nand U49068 (N_49068,N_48650,N_48896);
nor U49069 (N_49069,N_48928,N_48787);
and U49070 (N_49070,N_48588,N_48537);
and U49071 (N_49071,N_48780,N_48842);
nor U49072 (N_49072,N_48546,N_48983);
or U49073 (N_49073,N_48577,N_48557);
or U49074 (N_49074,N_48811,N_48812);
nor U49075 (N_49075,N_48863,N_48894);
nand U49076 (N_49076,N_48582,N_48611);
nor U49077 (N_49077,N_48881,N_48565);
and U49078 (N_49078,N_48979,N_48561);
or U49079 (N_49079,N_48968,N_48788);
xnor U49080 (N_49080,N_48549,N_48596);
nor U49081 (N_49081,N_48704,N_48528);
xor U49082 (N_49082,N_48840,N_48769);
nor U49083 (N_49083,N_48743,N_48784);
xor U49084 (N_49084,N_48850,N_48509);
or U49085 (N_49085,N_48916,N_48990);
and U49086 (N_49086,N_48804,N_48766);
and U49087 (N_49087,N_48963,N_48614);
and U49088 (N_49088,N_48531,N_48871);
and U49089 (N_49089,N_48654,N_48728);
nand U49090 (N_49090,N_48853,N_48688);
and U49091 (N_49091,N_48913,N_48980);
or U49092 (N_49092,N_48790,N_48775);
nor U49093 (N_49093,N_48576,N_48892);
nand U49094 (N_49094,N_48671,N_48657);
nor U49095 (N_49095,N_48827,N_48594);
nand U49096 (N_49096,N_48866,N_48883);
nand U49097 (N_49097,N_48541,N_48947);
or U49098 (N_49098,N_48706,N_48864);
xor U49099 (N_49099,N_48635,N_48652);
or U49100 (N_49100,N_48765,N_48629);
nor U49101 (N_49101,N_48943,N_48506);
nand U49102 (N_49102,N_48539,N_48902);
nor U49103 (N_49103,N_48532,N_48691);
xnor U49104 (N_49104,N_48970,N_48710);
nand U49105 (N_49105,N_48781,N_48738);
xnor U49106 (N_49106,N_48814,N_48951);
nor U49107 (N_49107,N_48589,N_48932);
or U49108 (N_49108,N_48985,N_48793);
nor U49109 (N_49109,N_48605,N_48914);
nand U49110 (N_49110,N_48767,N_48661);
nand U49111 (N_49111,N_48504,N_48680);
nand U49112 (N_49112,N_48760,N_48957);
and U49113 (N_49113,N_48854,N_48949);
nor U49114 (N_49114,N_48774,N_48518);
nor U49115 (N_49115,N_48672,N_48722);
or U49116 (N_49116,N_48692,N_48527);
nor U49117 (N_49117,N_48900,N_48583);
and U49118 (N_49118,N_48855,N_48826);
nand U49119 (N_49119,N_48829,N_48648);
nor U49120 (N_49120,N_48993,N_48505);
nor U49121 (N_49121,N_48868,N_48719);
nand U49122 (N_49122,N_48705,N_48636);
or U49123 (N_49123,N_48977,N_48848);
or U49124 (N_49124,N_48739,N_48674);
nor U49125 (N_49125,N_48665,N_48572);
nand U49126 (N_49126,N_48940,N_48889);
nand U49127 (N_49127,N_48919,N_48656);
nor U49128 (N_49128,N_48836,N_48761);
or U49129 (N_49129,N_48802,N_48820);
xnor U49130 (N_49130,N_48593,N_48893);
or U49131 (N_49131,N_48961,N_48514);
nand U49132 (N_49132,N_48603,N_48831);
nand U49133 (N_49133,N_48712,N_48800);
nand U49134 (N_49134,N_48677,N_48591);
and U49135 (N_49135,N_48903,N_48651);
and U49136 (N_49136,N_48756,N_48875);
nand U49137 (N_49137,N_48555,N_48740);
and U49138 (N_49138,N_48999,N_48717);
and U49139 (N_49139,N_48590,N_48830);
or U49140 (N_49140,N_48644,N_48624);
nor U49141 (N_49141,N_48616,N_48930);
or U49142 (N_49142,N_48939,N_48570);
xor U49143 (N_49143,N_48638,N_48995);
nor U49144 (N_49144,N_48708,N_48911);
nor U49145 (N_49145,N_48716,N_48751);
and U49146 (N_49146,N_48713,N_48870);
nand U49147 (N_49147,N_48803,N_48581);
nor U49148 (N_49148,N_48923,N_48954);
and U49149 (N_49149,N_48642,N_48615);
nand U49150 (N_49150,N_48782,N_48630);
xnor U49151 (N_49151,N_48521,N_48772);
or U49152 (N_49152,N_48634,N_48633);
and U49153 (N_49153,N_48976,N_48835);
and U49154 (N_49154,N_48729,N_48763);
nand U49155 (N_49155,N_48724,N_48741);
or U49156 (N_49156,N_48818,N_48815);
nor U49157 (N_49157,N_48695,N_48511);
nand U49158 (N_49158,N_48698,N_48845);
xnor U49159 (N_49159,N_48891,N_48832);
nand U49160 (N_49160,N_48676,N_48915);
and U49161 (N_49161,N_48987,N_48910);
and U49162 (N_49162,N_48748,N_48628);
nand U49163 (N_49163,N_48898,N_48627);
nand U49164 (N_49164,N_48515,N_48584);
nand U49165 (N_49165,N_48877,N_48562);
nor U49166 (N_49166,N_48520,N_48500);
xor U49167 (N_49167,N_48512,N_48554);
or U49168 (N_49168,N_48598,N_48612);
nand U49169 (N_49169,N_48703,N_48726);
nor U49170 (N_49170,N_48924,N_48510);
nand U49171 (N_49171,N_48847,N_48762);
xor U49172 (N_49172,N_48600,N_48770);
or U49173 (N_49173,N_48901,N_48737);
xnor U49174 (N_49174,N_48758,N_48965);
and U49175 (N_49175,N_48991,N_48673);
or U49176 (N_49176,N_48822,N_48632);
or U49177 (N_49177,N_48643,N_48720);
nor U49178 (N_49178,N_48545,N_48922);
nand U49179 (N_49179,N_48857,N_48626);
nor U49180 (N_49180,N_48597,N_48622);
nand U49181 (N_49181,N_48711,N_48926);
nand U49182 (N_49182,N_48768,N_48935);
or U49183 (N_49183,N_48604,N_48994);
or U49184 (N_49184,N_48873,N_48944);
or U49185 (N_49185,N_48921,N_48696);
or U49186 (N_49186,N_48721,N_48874);
nand U49187 (N_49187,N_48538,N_48755);
or U49188 (N_49188,N_48810,N_48574);
nand U49189 (N_49189,N_48533,N_48887);
or U49190 (N_49190,N_48882,N_48801);
nand U49191 (N_49191,N_48846,N_48952);
and U49192 (N_49192,N_48752,N_48799);
and U49193 (N_49193,N_48568,N_48553);
nor U49194 (N_49194,N_48575,N_48548);
and U49195 (N_49195,N_48933,N_48684);
and U49196 (N_49196,N_48872,N_48908);
nand U49197 (N_49197,N_48825,N_48764);
nand U49198 (N_49198,N_48805,N_48731);
nor U49199 (N_49199,N_48595,N_48997);
or U49200 (N_49200,N_48905,N_48608);
and U49201 (N_49201,N_48733,N_48886);
or U49202 (N_49202,N_48888,N_48956);
xnor U49203 (N_49203,N_48607,N_48530);
nor U49204 (N_49204,N_48513,N_48699);
nor U49205 (N_49205,N_48981,N_48938);
nand U49206 (N_49206,N_48662,N_48986);
or U49207 (N_49207,N_48571,N_48754);
and U49208 (N_49208,N_48678,N_48867);
or U49209 (N_49209,N_48962,N_48534);
or U49210 (N_49210,N_48610,N_48727);
nand U49211 (N_49211,N_48659,N_48789);
nor U49212 (N_49212,N_48759,N_48798);
nand U49213 (N_49213,N_48552,N_48702);
nor U49214 (N_49214,N_48860,N_48959);
and U49215 (N_49215,N_48839,N_48809);
nor U49216 (N_49216,N_48895,N_48687);
or U49217 (N_49217,N_48966,N_48601);
or U49218 (N_49218,N_48535,N_48974);
xnor U49219 (N_49219,N_48669,N_48794);
nor U49220 (N_49220,N_48564,N_48556);
and U49221 (N_49221,N_48819,N_48666);
nor U49222 (N_49222,N_48569,N_48946);
nor U49223 (N_49223,N_48683,N_48953);
nor U49224 (N_49224,N_48619,N_48715);
or U49225 (N_49225,N_48992,N_48508);
or U49226 (N_49226,N_48907,N_48950);
or U49227 (N_49227,N_48655,N_48524);
or U49228 (N_49228,N_48613,N_48964);
or U49229 (N_49229,N_48880,N_48567);
or U49230 (N_49230,N_48686,N_48645);
nor U49231 (N_49231,N_48563,N_48523);
nor U49232 (N_49232,N_48700,N_48783);
and U49233 (N_49233,N_48653,N_48718);
or U49234 (N_49234,N_48540,N_48971);
xor U49235 (N_49235,N_48529,N_48664);
and U49236 (N_49236,N_48912,N_48806);
nor U49237 (N_49237,N_48679,N_48519);
or U49238 (N_49238,N_48631,N_48730);
nor U49239 (N_49239,N_48920,N_48785);
and U49240 (N_49240,N_48689,N_48639);
and U49241 (N_49241,N_48736,N_48975);
xnor U49242 (N_49242,N_48937,N_48578);
and U49243 (N_49243,N_48808,N_48984);
or U49244 (N_49244,N_48837,N_48858);
and U49245 (N_49245,N_48618,N_48909);
nor U49246 (N_49246,N_48753,N_48869);
or U49247 (N_49247,N_48609,N_48602);
or U49248 (N_49248,N_48746,N_48929);
and U49249 (N_49249,N_48841,N_48925);
nand U49250 (N_49250,N_48904,N_48919);
nand U49251 (N_49251,N_48984,N_48989);
xor U49252 (N_49252,N_48837,N_48940);
nor U49253 (N_49253,N_48747,N_48709);
nand U49254 (N_49254,N_48527,N_48649);
or U49255 (N_49255,N_48680,N_48621);
and U49256 (N_49256,N_48746,N_48636);
nor U49257 (N_49257,N_48505,N_48705);
nand U49258 (N_49258,N_48733,N_48945);
nor U49259 (N_49259,N_48934,N_48837);
or U49260 (N_49260,N_48760,N_48926);
xnor U49261 (N_49261,N_48643,N_48694);
nor U49262 (N_49262,N_48987,N_48610);
or U49263 (N_49263,N_48750,N_48661);
nor U49264 (N_49264,N_48641,N_48954);
nand U49265 (N_49265,N_48663,N_48793);
nor U49266 (N_49266,N_48754,N_48745);
nor U49267 (N_49267,N_48633,N_48670);
nor U49268 (N_49268,N_48816,N_48901);
or U49269 (N_49269,N_48730,N_48999);
and U49270 (N_49270,N_48916,N_48798);
xor U49271 (N_49271,N_48635,N_48566);
nor U49272 (N_49272,N_48936,N_48842);
and U49273 (N_49273,N_48541,N_48890);
and U49274 (N_49274,N_48805,N_48944);
xnor U49275 (N_49275,N_48505,N_48714);
nand U49276 (N_49276,N_48884,N_48917);
xor U49277 (N_49277,N_48658,N_48581);
and U49278 (N_49278,N_48939,N_48872);
nand U49279 (N_49279,N_48644,N_48733);
and U49280 (N_49280,N_48769,N_48865);
and U49281 (N_49281,N_48886,N_48525);
or U49282 (N_49282,N_48879,N_48787);
and U49283 (N_49283,N_48914,N_48948);
nand U49284 (N_49284,N_48610,N_48768);
nand U49285 (N_49285,N_48842,N_48920);
and U49286 (N_49286,N_48894,N_48666);
xnor U49287 (N_49287,N_48976,N_48813);
nor U49288 (N_49288,N_48818,N_48798);
or U49289 (N_49289,N_48976,N_48936);
nor U49290 (N_49290,N_48964,N_48837);
and U49291 (N_49291,N_48753,N_48881);
or U49292 (N_49292,N_48640,N_48945);
nor U49293 (N_49293,N_48840,N_48738);
and U49294 (N_49294,N_48920,N_48848);
nand U49295 (N_49295,N_48980,N_48701);
and U49296 (N_49296,N_48721,N_48678);
or U49297 (N_49297,N_48661,N_48673);
and U49298 (N_49298,N_48506,N_48925);
nor U49299 (N_49299,N_48684,N_48858);
nand U49300 (N_49300,N_48846,N_48822);
or U49301 (N_49301,N_48821,N_48669);
xnor U49302 (N_49302,N_48909,N_48695);
nand U49303 (N_49303,N_48540,N_48938);
and U49304 (N_49304,N_48552,N_48741);
or U49305 (N_49305,N_48649,N_48770);
nand U49306 (N_49306,N_48744,N_48668);
nor U49307 (N_49307,N_48765,N_48722);
or U49308 (N_49308,N_48690,N_48767);
xor U49309 (N_49309,N_48736,N_48900);
nor U49310 (N_49310,N_48554,N_48737);
and U49311 (N_49311,N_48718,N_48893);
nor U49312 (N_49312,N_48512,N_48535);
and U49313 (N_49313,N_48932,N_48536);
nor U49314 (N_49314,N_48694,N_48513);
xor U49315 (N_49315,N_48847,N_48969);
and U49316 (N_49316,N_48531,N_48525);
nor U49317 (N_49317,N_48934,N_48561);
nor U49318 (N_49318,N_48614,N_48973);
nand U49319 (N_49319,N_48965,N_48567);
xnor U49320 (N_49320,N_48644,N_48970);
and U49321 (N_49321,N_48784,N_48639);
nor U49322 (N_49322,N_48729,N_48751);
nor U49323 (N_49323,N_48688,N_48919);
or U49324 (N_49324,N_48748,N_48729);
or U49325 (N_49325,N_48669,N_48756);
nand U49326 (N_49326,N_48843,N_48898);
nand U49327 (N_49327,N_48990,N_48723);
or U49328 (N_49328,N_48900,N_48803);
and U49329 (N_49329,N_48776,N_48847);
and U49330 (N_49330,N_48959,N_48660);
nand U49331 (N_49331,N_48972,N_48686);
and U49332 (N_49332,N_48738,N_48548);
nor U49333 (N_49333,N_48659,N_48850);
xor U49334 (N_49334,N_48590,N_48540);
or U49335 (N_49335,N_48571,N_48941);
nand U49336 (N_49336,N_48505,N_48713);
nand U49337 (N_49337,N_48905,N_48892);
nand U49338 (N_49338,N_48851,N_48506);
or U49339 (N_49339,N_48784,N_48548);
and U49340 (N_49340,N_48921,N_48908);
or U49341 (N_49341,N_48864,N_48574);
and U49342 (N_49342,N_48717,N_48805);
nor U49343 (N_49343,N_48804,N_48685);
nand U49344 (N_49344,N_48828,N_48723);
or U49345 (N_49345,N_48996,N_48601);
nand U49346 (N_49346,N_48744,N_48643);
xnor U49347 (N_49347,N_48524,N_48768);
nand U49348 (N_49348,N_48750,N_48635);
nand U49349 (N_49349,N_48722,N_48693);
or U49350 (N_49350,N_48660,N_48804);
nor U49351 (N_49351,N_48906,N_48580);
and U49352 (N_49352,N_48639,N_48722);
or U49353 (N_49353,N_48722,N_48867);
or U49354 (N_49354,N_48983,N_48780);
and U49355 (N_49355,N_48696,N_48632);
nand U49356 (N_49356,N_48777,N_48973);
nand U49357 (N_49357,N_48956,N_48831);
nor U49358 (N_49358,N_48512,N_48653);
or U49359 (N_49359,N_48704,N_48518);
nand U49360 (N_49360,N_48679,N_48775);
and U49361 (N_49361,N_48726,N_48737);
nor U49362 (N_49362,N_48570,N_48803);
and U49363 (N_49363,N_48951,N_48940);
nand U49364 (N_49364,N_48681,N_48861);
or U49365 (N_49365,N_48929,N_48939);
or U49366 (N_49366,N_48601,N_48719);
and U49367 (N_49367,N_48825,N_48573);
nor U49368 (N_49368,N_48915,N_48998);
nor U49369 (N_49369,N_48597,N_48509);
or U49370 (N_49370,N_48562,N_48611);
xor U49371 (N_49371,N_48948,N_48572);
or U49372 (N_49372,N_48758,N_48714);
and U49373 (N_49373,N_48856,N_48785);
xor U49374 (N_49374,N_48845,N_48938);
nand U49375 (N_49375,N_48795,N_48750);
and U49376 (N_49376,N_48691,N_48565);
and U49377 (N_49377,N_48851,N_48555);
and U49378 (N_49378,N_48978,N_48993);
and U49379 (N_49379,N_48714,N_48902);
or U49380 (N_49380,N_48985,N_48748);
and U49381 (N_49381,N_48651,N_48818);
or U49382 (N_49382,N_48962,N_48817);
xor U49383 (N_49383,N_48512,N_48796);
or U49384 (N_49384,N_48746,N_48552);
or U49385 (N_49385,N_48719,N_48757);
nand U49386 (N_49386,N_48715,N_48878);
or U49387 (N_49387,N_48942,N_48634);
or U49388 (N_49388,N_48564,N_48848);
and U49389 (N_49389,N_48669,N_48898);
or U49390 (N_49390,N_48751,N_48978);
and U49391 (N_49391,N_48526,N_48730);
and U49392 (N_49392,N_48570,N_48761);
or U49393 (N_49393,N_48588,N_48681);
xnor U49394 (N_49394,N_48933,N_48533);
xor U49395 (N_49395,N_48722,N_48813);
nand U49396 (N_49396,N_48794,N_48781);
and U49397 (N_49397,N_48808,N_48675);
nand U49398 (N_49398,N_48931,N_48685);
or U49399 (N_49399,N_48519,N_48646);
and U49400 (N_49400,N_48537,N_48947);
nor U49401 (N_49401,N_48800,N_48656);
or U49402 (N_49402,N_48585,N_48695);
xor U49403 (N_49403,N_48973,N_48935);
or U49404 (N_49404,N_48599,N_48573);
and U49405 (N_49405,N_48511,N_48685);
nand U49406 (N_49406,N_48936,N_48557);
nor U49407 (N_49407,N_48797,N_48980);
nor U49408 (N_49408,N_48627,N_48933);
nand U49409 (N_49409,N_48883,N_48899);
nand U49410 (N_49410,N_48938,N_48800);
nand U49411 (N_49411,N_48941,N_48717);
or U49412 (N_49412,N_48757,N_48581);
or U49413 (N_49413,N_48687,N_48868);
or U49414 (N_49414,N_48981,N_48667);
nand U49415 (N_49415,N_48996,N_48815);
and U49416 (N_49416,N_48804,N_48577);
and U49417 (N_49417,N_48982,N_48554);
xnor U49418 (N_49418,N_48549,N_48652);
nor U49419 (N_49419,N_48836,N_48915);
nor U49420 (N_49420,N_48792,N_48659);
xor U49421 (N_49421,N_48811,N_48850);
and U49422 (N_49422,N_48659,N_48730);
nand U49423 (N_49423,N_48661,N_48660);
nand U49424 (N_49424,N_48501,N_48879);
nor U49425 (N_49425,N_48654,N_48863);
nor U49426 (N_49426,N_48525,N_48508);
and U49427 (N_49427,N_48982,N_48886);
or U49428 (N_49428,N_48812,N_48857);
or U49429 (N_49429,N_48689,N_48596);
or U49430 (N_49430,N_48849,N_48501);
and U49431 (N_49431,N_48647,N_48675);
nand U49432 (N_49432,N_48824,N_48969);
nor U49433 (N_49433,N_48911,N_48795);
and U49434 (N_49434,N_48804,N_48993);
nand U49435 (N_49435,N_48967,N_48845);
xor U49436 (N_49436,N_48840,N_48788);
xor U49437 (N_49437,N_48749,N_48750);
and U49438 (N_49438,N_48560,N_48631);
nor U49439 (N_49439,N_48961,N_48620);
or U49440 (N_49440,N_48813,N_48628);
or U49441 (N_49441,N_48733,N_48838);
nor U49442 (N_49442,N_48548,N_48552);
and U49443 (N_49443,N_48818,N_48863);
nor U49444 (N_49444,N_48949,N_48982);
and U49445 (N_49445,N_48985,N_48575);
xor U49446 (N_49446,N_48855,N_48796);
or U49447 (N_49447,N_48758,N_48890);
nand U49448 (N_49448,N_48552,N_48770);
nand U49449 (N_49449,N_48669,N_48607);
xnor U49450 (N_49450,N_48590,N_48564);
nand U49451 (N_49451,N_48798,N_48769);
nor U49452 (N_49452,N_48951,N_48685);
nand U49453 (N_49453,N_48896,N_48544);
nor U49454 (N_49454,N_48559,N_48623);
and U49455 (N_49455,N_48784,N_48706);
and U49456 (N_49456,N_48521,N_48529);
or U49457 (N_49457,N_48517,N_48901);
nor U49458 (N_49458,N_48612,N_48870);
xor U49459 (N_49459,N_48592,N_48948);
and U49460 (N_49460,N_48868,N_48677);
nor U49461 (N_49461,N_48884,N_48517);
and U49462 (N_49462,N_48875,N_48914);
and U49463 (N_49463,N_48839,N_48585);
xnor U49464 (N_49464,N_48987,N_48646);
nor U49465 (N_49465,N_48900,N_48844);
and U49466 (N_49466,N_48527,N_48964);
and U49467 (N_49467,N_48824,N_48770);
and U49468 (N_49468,N_48922,N_48837);
nor U49469 (N_49469,N_48838,N_48925);
or U49470 (N_49470,N_48685,N_48802);
nor U49471 (N_49471,N_48933,N_48693);
and U49472 (N_49472,N_48963,N_48881);
or U49473 (N_49473,N_48767,N_48515);
and U49474 (N_49474,N_48787,N_48930);
nand U49475 (N_49475,N_48501,N_48888);
nor U49476 (N_49476,N_48910,N_48768);
nand U49477 (N_49477,N_48569,N_48653);
or U49478 (N_49478,N_48795,N_48566);
nor U49479 (N_49479,N_48820,N_48979);
and U49480 (N_49480,N_48909,N_48522);
nand U49481 (N_49481,N_48823,N_48913);
and U49482 (N_49482,N_48732,N_48764);
or U49483 (N_49483,N_48514,N_48883);
nand U49484 (N_49484,N_48631,N_48724);
and U49485 (N_49485,N_48920,N_48579);
nor U49486 (N_49486,N_48621,N_48623);
nand U49487 (N_49487,N_48602,N_48962);
and U49488 (N_49488,N_48729,N_48657);
and U49489 (N_49489,N_48776,N_48533);
nor U49490 (N_49490,N_48954,N_48746);
or U49491 (N_49491,N_48552,N_48868);
nand U49492 (N_49492,N_48966,N_48665);
or U49493 (N_49493,N_48719,N_48861);
or U49494 (N_49494,N_48546,N_48570);
nor U49495 (N_49495,N_48631,N_48706);
nor U49496 (N_49496,N_48828,N_48766);
and U49497 (N_49497,N_48742,N_48779);
xnor U49498 (N_49498,N_48552,N_48613);
xnor U49499 (N_49499,N_48751,N_48689);
xor U49500 (N_49500,N_49252,N_49256);
or U49501 (N_49501,N_49019,N_49209);
nand U49502 (N_49502,N_49216,N_49100);
nor U49503 (N_49503,N_49284,N_49345);
xor U49504 (N_49504,N_49364,N_49208);
and U49505 (N_49505,N_49101,N_49144);
nor U49506 (N_49506,N_49304,N_49108);
nor U49507 (N_49507,N_49259,N_49131);
and U49508 (N_49508,N_49330,N_49343);
nand U49509 (N_49509,N_49319,N_49480);
or U49510 (N_49510,N_49188,N_49384);
and U49511 (N_49511,N_49309,N_49196);
or U49512 (N_49512,N_49268,N_49288);
and U49513 (N_49513,N_49102,N_49221);
nand U49514 (N_49514,N_49332,N_49064);
or U49515 (N_49515,N_49308,N_49126);
or U49516 (N_49516,N_49392,N_49408);
nand U49517 (N_49517,N_49241,N_49041);
nand U49518 (N_49518,N_49334,N_49464);
or U49519 (N_49519,N_49470,N_49119);
and U49520 (N_49520,N_49182,N_49389);
and U49521 (N_49521,N_49289,N_49206);
and U49522 (N_49522,N_49032,N_49331);
and U49523 (N_49523,N_49140,N_49461);
nand U49524 (N_49524,N_49025,N_49129);
or U49525 (N_49525,N_49281,N_49254);
or U49526 (N_49526,N_49454,N_49077);
xnor U49527 (N_49527,N_49061,N_49214);
nand U49528 (N_49528,N_49431,N_49350);
nor U49529 (N_49529,N_49085,N_49072);
and U49530 (N_49530,N_49133,N_49448);
or U49531 (N_49531,N_49030,N_49462);
nand U49532 (N_49532,N_49486,N_49298);
and U49533 (N_49533,N_49482,N_49321);
nor U49534 (N_49534,N_49029,N_49436);
nand U49535 (N_49535,N_49409,N_49283);
nand U49536 (N_49536,N_49338,N_49230);
nor U49537 (N_49537,N_49406,N_49478);
xor U49538 (N_49538,N_49477,N_49494);
nand U49539 (N_49539,N_49179,N_49273);
and U49540 (N_49540,N_49247,N_49390);
or U49541 (N_49541,N_49191,N_49336);
or U49542 (N_49542,N_49178,N_49271);
nor U49543 (N_49543,N_49052,N_49489);
nand U49544 (N_49544,N_49099,N_49377);
nor U49545 (N_49545,N_49050,N_49204);
or U49546 (N_49546,N_49347,N_49376);
and U49547 (N_49547,N_49155,N_49495);
xor U49548 (N_49548,N_49276,N_49493);
nand U49549 (N_49549,N_49156,N_49311);
nor U49550 (N_49550,N_49388,N_49199);
nor U49551 (N_49551,N_49357,N_49459);
nor U49552 (N_49552,N_49250,N_49112);
or U49553 (N_49553,N_49143,N_49103);
and U49554 (N_49554,N_49068,N_49255);
and U49555 (N_49555,N_49344,N_49387);
nor U49556 (N_49556,N_49487,N_49246);
nand U49557 (N_49557,N_49303,N_49257);
nor U49558 (N_49558,N_49456,N_49203);
or U49559 (N_49559,N_49318,N_49240);
or U49560 (N_49560,N_49003,N_49417);
and U49561 (N_49561,N_49114,N_49346);
nor U49562 (N_49562,N_49323,N_49136);
nor U49563 (N_49563,N_49186,N_49149);
nand U49564 (N_49564,N_49253,N_49135);
nor U49565 (N_49565,N_49429,N_49139);
or U49566 (N_49566,N_49169,N_49094);
nor U49567 (N_49567,N_49123,N_49227);
and U49568 (N_49568,N_49127,N_49484);
and U49569 (N_49569,N_49235,N_49095);
nor U49570 (N_49570,N_49457,N_49010);
or U49571 (N_49571,N_49258,N_49084);
or U49572 (N_49572,N_49016,N_49471);
nand U49573 (N_49573,N_49231,N_49385);
nor U49574 (N_49574,N_49349,N_49411);
nand U49575 (N_49575,N_49372,N_49195);
and U49576 (N_49576,N_49212,N_49382);
nor U49577 (N_49577,N_49189,N_49292);
nand U49578 (N_49578,N_49138,N_49491);
or U49579 (N_49579,N_49415,N_49176);
nor U49580 (N_49580,N_49205,N_49055);
and U49581 (N_49581,N_49090,N_49224);
and U49582 (N_49582,N_49442,N_49481);
nand U49583 (N_49583,N_49180,N_49402);
nor U49584 (N_49584,N_49437,N_49162);
xor U49585 (N_49585,N_49386,N_49369);
nand U49586 (N_49586,N_49215,N_49071);
xnor U49587 (N_49587,N_49297,N_49210);
and U49588 (N_49588,N_49360,N_49065);
nand U49589 (N_49589,N_49428,N_49058);
nor U49590 (N_49590,N_49383,N_49109);
or U49591 (N_49591,N_49416,N_49479);
nand U49592 (N_49592,N_49042,N_49053);
and U49593 (N_49593,N_49290,N_49165);
nor U49594 (N_49594,N_49317,N_49286);
xor U49595 (N_49595,N_49399,N_49089);
and U49596 (N_49596,N_49020,N_49096);
or U49597 (N_49597,N_49453,N_49353);
nand U49598 (N_49598,N_49397,N_49274);
xor U49599 (N_49599,N_49130,N_49352);
nor U49600 (N_49600,N_49356,N_49467);
nor U49601 (N_49601,N_49031,N_49223);
and U49602 (N_49602,N_49418,N_49026);
or U49603 (N_49603,N_49435,N_49159);
nand U49604 (N_49604,N_49270,N_49358);
nor U49605 (N_49605,N_49219,N_49440);
nand U49606 (N_49606,N_49426,N_49266);
and U49607 (N_49607,N_49451,N_49198);
nand U49608 (N_49608,N_49007,N_49009);
nor U49609 (N_49609,N_49312,N_49296);
xnor U49610 (N_49610,N_49264,N_49217);
nor U49611 (N_49611,N_49306,N_49115);
xor U49612 (N_49612,N_49122,N_49335);
and U49613 (N_49613,N_49245,N_49022);
or U49614 (N_49614,N_49151,N_49174);
nor U49615 (N_49615,N_49474,N_49063);
nor U49616 (N_49616,N_49412,N_49171);
nor U49617 (N_49617,N_49237,N_49234);
or U49618 (N_49618,N_49425,N_49326);
or U49619 (N_49619,N_49472,N_49076);
nor U49620 (N_49620,N_49152,N_49260);
and U49621 (N_49621,N_49083,N_49476);
or U49622 (N_49622,N_49314,N_49341);
or U49623 (N_49623,N_49396,N_49157);
nand U49624 (N_49624,N_49069,N_49267);
or U49625 (N_49625,N_49299,N_49348);
xor U49626 (N_49626,N_49465,N_49438);
xor U49627 (N_49627,N_49407,N_49012);
nor U49628 (N_49628,N_49499,N_49430);
nand U49629 (N_49629,N_49351,N_49413);
and U49630 (N_49630,N_49036,N_49327);
nor U49631 (N_49631,N_49125,N_49378);
or U49632 (N_49632,N_49124,N_49024);
nor U49633 (N_49633,N_49229,N_49232);
or U49634 (N_49634,N_49164,N_49211);
or U49635 (N_49635,N_49488,N_49458);
and U49636 (N_49636,N_49166,N_49177);
and U49637 (N_49637,N_49294,N_49490);
xnor U49638 (N_49638,N_49104,N_49265);
nor U49639 (N_49639,N_49170,N_49371);
nand U49640 (N_49640,N_49339,N_49080);
nor U49641 (N_49641,N_49316,N_49074);
nand U49642 (N_49642,N_49220,N_49280);
and U49643 (N_49643,N_49066,N_49048);
nor U49644 (N_49644,N_49365,N_49106);
nor U49645 (N_49645,N_49410,N_49146);
or U49646 (N_49646,N_49051,N_49118);
nand U49647 (N_49647,N_49008,N_49049);
or U49648 (N_49648,N_49374,N_49168);
nand U49649 (N_49649,N_49173,N_49006);
or U49650 (N_49650,N_49145,N_49087);
or U49651 (N_49651,N_49185,N_49263);
nand U49652 (N_49652,N_49450,N_49107);
nor U49653 (N_49653,N_49251,N_49302);
or U49654 (N_49654,N_49455,N_49277);
or U49655 (N_49655,N_49466,N_49313);
nor U49656 (N_49656,N_49027,N_49307);
xnor U49657 (N_49657,N_49393,N_49422);
nand U49658 (N_49658,N_49395,N_49305);
or U49659 (N_49659,N_49391,N_49197);
or U49660 (N_49660,N_49282,N_49405);
nor U49661 (N_49661,N_49021,N_49043);
nor U49662 (N_49662,N_49207,N_49213);
nand U49663 (N_49663,N_49278,N_49359);
nor U49664 (N_49664,N_49034,N_49194);
nand U49665 (N_49665,N_49449,N_49400);
or U49666 (N_49666,N_49329,N_49293);
nor U49667 (N_49667,N_49483,N_49023);
or U49668 (N_49668,N_49243,N_49242);
nor U49669 (N_49669,N_49128,N_49423);
and U49670 (N_49670,N_49262,N_49161);
or U49671 (N_49671,N_49047,N_49301);
nand U49672 (N_49672,N_49088,N_49040);
or U49673 (N_49673,N_49498,N_49175);
nand U49674 (N_49674,N_49355,N_49419);
nor U49675 (N_49675,N_49045,N_49249);
nor U49676 (N_49676,N_49018,N_49086);
nor U49677 (N_49677,N_49398,N_49075);
or U49678 (N_49678,N_49366,N_49005);
or U49679 (N_49679,N_49037,N_49379);
nand U49680 (N_49680,N_49000,N_49187);
nor U49681 (N_49681,N_49137,N_49113);
nor U49682 (N_49682,N_49433,N_49272);
nor U49683 (N_49683,N_49078,N_49233);
or U49684 (N_49684,N_49193,N_49097);
nand U49685 (N_49685,N_49081,N_49424);
nor U49686 (N_49686,N_49443,N_49062);
nand U49687 (N_49687,N_49291,N_49147);
or U49688 (N_49688,N_49117,N_49222);
or U49689 (N_49689,N_49035,N_49340);
and U49690 (N_49690,N_49060,N_49445);
xor U49691 (N_49691,N_49160,N_49275);
or U49692 (N_49692,N_49322,N_49333);
or U49693 (N_49693,N_49141,N_49401);
xnor U49694 (N_49694,N_49226,N_49046);
and U49695 (N_49695,N_49015,N_49218);
xnor U49696 (N_49696,N_49201,N_49380);
nand U49697 (N_49697,N_49142,N_49192);
or U49698 (N_49698,N_49287,N_49497);
nand U49699 (N_49699,N_49093,N_49367);
and U49700 (N_49700,N_49056,N_49420);
and U49701 (N_49701,N_49121,N_49202);
nor U49702 (N_49702,N_49342,N_49325);
nand U49703 (N_49703,N_49167,N_49070);
nor U49704 (N_49704,N_49446,N_49238);
nor U49705 (N_49705,N_49116,N_49375);
nor U49706 (N_49706,N_49285,N_49039);
and U49707 (N_49707,N_49363,N_49044);
nor U49708 (N_49708,N_49183,N_49427);
or U49709 (N_49709,N_49381,N_49404);
nor U49710 (N_49710,N_49134,N_49485);
xnor U49711 (N_49711,N_49315,N_49432);
and U49712 (N_49712,N_49200,N_49496);
and U49713 (N_49713,N_49261,N_49225);
and U49714 (N_49714,N_49033,N_49434);
and U49715 (N_49715,N_49001,N_49011);
and U49716 (N_49716,N_49236,N_49362);
and U49717 (N_49717,N_49414,N_49150);
and U49718 (N_49718,N_49463,N_49004);
or U49719 (N_49719,N_49067,N_49190);
nor U49720 (N_49720,N_49468,N_49054);
xnor U49721 (N_49721,N_49337,N_49403);
nor U49722 (N_49722,N_49073,N_49300);
nor U49723 (N_49723,N_49228,N_49017);
xnor U49724 (N_49724,N_49269,N_49370);
nand U49725 (N_49725,N_49394,N_49013);
or U49726 (N_49726,N_49244,N_49132);
and U49727 (N_49727,N_49098,N_49091);
or U49728 (N_49728,N_49059,N_49248);
or U49729 (N_49729,N_49361,N_49368);
nand U49730 (N_49730,N_49239,N_49002);
and U49731 (N_49731,N_49328,N_49492);
nand U49732 (N_49732,N_49158,N_49460);
xor U49733 (N_49733,N_49057,N_49439);
and U49734 (N_49734,N_49441,N_49110);
or U49735 (N_49735,N_49105,N_49444);
or U49736 (N_49736,N_49310,N_49092);
xnor U49737 (N_49737,N_49421,N_49038);
nor U49738 (N_49738,N_49373,N_49111);
xnor U49739 (N_49739,N_49324,N_49447);
nor U49740 (N_49740,N_49475,N_49354);
nor U49741 (N_49741,N_49163,N_49082);
or U49742 (N_49742,N_49172,N_49181);
nor U49743 (N_49743,N_49120,N_49028);
nand U49744 (N_49744,N_49154,N_49473);
and U49745 (N_49745,N_49469,N_49279);
nand U49746 (N_49746,N_49184,N_49320);
nor U49747 (N_49747,N_49148,N_49079);
or U49748 (N_49748,N_49153,N_49295);
nor U49749 (N_49749,N_49014,N_49452);
and U49750 (N_49750,N_49012,N_49280);
nand U49751 (N_49751,N_49425,N_49296);
xnor U49752 (N_49752,N_49362,N_49244);
and U49753 (N_49753,N_49004,N_49456);
nand U49754 (N_49754,N_49253,N_49374);
nor U49755 (N_49755,N_49473,N_49243);
xor U49756 (N_49756,N_49355,N_49428);
and U49757 (N_49757,N_49211,N_49028);
and U49758 (N_49758,N_49123,N_49005);
nor U49759 (N_49759,N_49180,N_49484);
and U49760 (N_49760,N_49184,N_49013);
nor U49761 (N_49761,N_49279,N_49243);
nor U49762 (N_49762,N_49324,N_49437);
nand U49763 (N_49763,N_49384,N_49204);
xnor U49764 (N_49764,N_49493,N_49366);
xnor U49765 (N_49765,N_49226,N_49402);
nor U49766 (N_49766,N_49447,N_49486);
nor U49767 (N_49767,N_49410,N_49326);
and U49768 (N_49768,N_49401,N_49176);
nor U49769 (N_49769,N_49017,N_49412);
nor U49770 (N_49770,N_49234,N_49301);
or U49771 (N_49771,N_49218,N_49029);
and U49772 (N_49772,N_49442,N_49428);
nor U49773 (N_49773,N_49125,N_49240);
xnor U49774 (N_49774,N_49265,N_49215);
nor U49775 (N_49775,N_49303,N_49375);
and U49776 (N_49776,N_49439,N_49277);
nand U49777 (N_49777,N_49345,N_49212);
nand U49778 (N_49778,N_49059,N_49082);
nand U49779 (N_49779,N_49205,N_49350);
nand U49780 (N_49780,N_49140,N_49207);
nand U49781 (N_49781,N_49032,N_49220);
and U49782 (N_49782,N_49274,N_49364);
nand U49783 (N_49783,N_49498,N_49004);
or U49784 (N_49784,N_49043,N_49266);
nand U49785 (N_49785,N_49110,N_49117);
nor U49786 (N_49786,N_49367,N_49331);
nor U49787 (N_49787,N_49280,N_49216);
xnor U49788 (N_49788,N_49024,N_49453);
nand U49789 (N_49789,N_49017,N_49322);
or U49790 (N_49790,N_49177,N_49463);
and U49791 (N_49791,N_49353,N_49418);
nand U49792 (N_49792,N_49329,N_49051);
or U49793 (N_49793,N_49117,N_49353);
nor U49794 (N_49794,N_49052,N_49419);
nor U49795 (N_49795,N_49049,N_49304);
or U49796 (N_49796,N_49114,N_49255);
nor U49797 (N_49797,N_49180,N_49187);
or U49798 (N_49798,N_49453,N_49418);
nor U49799 (N_49799,N_49374,N_49075);
or U49800 (N_49800,N_49179,N_49264);
nand U49801 (N_49801,N_49048,N_49253);
nand U49802 (N_49802,N_49496,N_49484);
and U49803 (N_49803,N_49415,N_49075);
xnor U49804 (N_49804,N_49492,N_49414);
or U49805 (N_49805,N_49127,N_49216);
or U49806 (N_49806,N_49039,N_49437);
and U49807 (N_49807,N_49026,N_49129);
nor U49808 (N_49808,N_49187,N_49071);
nand U49809 (N_49809,N_49265,N_49342);
nand U49810 (N_49810,N_49412,N_49193);
nand U49811 (N_49811,N_49135,N_49295);
nand U49812 (N_49812,N_49486,N_49070);
and U49813 (N_49813,N_49215,N_49047);
nand U49814 (N_49814,N_49120,N_49135);
nor U49815 (N_49815,N_49302,N_49430);
nor U49816 (N_49816,N_49246,N_49147);
nor U49817 (N_49817,N_49126,N_49277);
nor U49818 (N_49818,N_49113,N_49173);
nor U49819 (N_49819,N_49005,N_49092);
nor U49820 (N_49820,N_49390,N_49455);
xnor U49821 (N_49821,N_49075,N_49191);
or U49822 (N_49822,N_49262,N_49341);
or U49823 (N_49823,N_49031,N_49498);
nor U49824 (N_49824,N_49361,N_49212);
xor U49825 (N_49825,N_49332,N_49212);
and U49826 (N_49826,N_49234,N_49019);
nor U49827 (N_49827,N_49286,N_49216);
and U49828 (N_49828,N_49329,N_49338);
or U49829 (N_49829,N_49185,N_49124);
xnor U49830 (N_49830,N_49029,N_49406);
nor U49831 (N_49831,N_49403,N_49019);
nor U49832 (N_49832,N_49360,N_49000);
nand U49833 (N_49833,N_49347,N_49212);
or U49834 (N_49834,N_49492,N_49145);
and U49835 (N_49835,N_49266,N_49019);
and U49836 (N_49836,N_49160,N_49038);
nor U49837 (N_49837,N_49358,N_49400);
or U49838 (N_49838,N_49403,N_49346);
nand U49839 (N_49839,N_49466,N_49078);
xnor U49840 (N_49840,N_49328,N_49102);
nor U49841 (N_49841,N_49008,N_49075);
or U49842 (N_49842,N_49464,N_49475);
or U49843 (N_49843,N_49390,N_49105);
and U49844 (N_49844,N_49373,N_49155);
and U49845 (N_49845,N_49130,N_49409);
nand U49846 (N_49846,N_49241,N_49181);
nand U49847 (N_49847,N_49405,N_49453);
nand U49848 (N_49848,N_49224,N_49322);
nand U49849 (N_49849,N_49450,N_49394);
nand U49850 (N_49850,N_49085,N_49043);
nand U49851 (N_49851,N_49317,N_49235);
and U49852 (N_49852,N_49188,N_49007);
nand U49853 (N_49853,N_49461,N_49229);
nand U49854 (N_49854,N_49248,N_49276);
and U49855 (N_49855,N_49444,N_49121);
or U49856 (N_49856,N_49202,N_49254);
and U49857 (N_49857,N_49383,N_49000);
xnor U49858 (N_49858,N_49455,N_49027);
nand U49859 (N_49859,N_49346,N_49395);
nand U49860 (N_49860,N_49381,N_49397);
nand U49861 (N_49861,N_49214,N_49292);
nand U49862 (N_49862,N_49023,N_49121);
nand U49863 (N_49863,N_49335,N_49049);
or U49864 (N_49864,N_49465,N_49236);
nor U49865 (N_49865,N_49325,N_49475);
nor U49866 (N_49866,N_49425,N_49178);
nor U49867 (N_49867,N_49229,N_49142);
nor U49868 (N_49868,N_49225,N_49004);
nand U49869 (N_49869,N_49348,N_49042);
nor U49870 (N_49870,N_49259,N_49411);
nor U49871 (N_49871,N_49320,N_49029);
and U49872 (N_49872,N_49352,N_49092);
xnor U49873 (N_49873,N_49133,N_49180);
and U49874 (N_49874,N_49417,N_49042);
or U49875 (N_49875,N_49457,N_49325);
nor U49876 (N_49876,N_49266,N_49346);
or U49877 (N_49877,N_49358,N_49285);
and U49878 (N_49878,N_49466,N_49373);
nand U49879 (N_49879,N_49174,N_49002);
or U49880 (N_49880,N_49310,N_49322);
xor U49881 (N_49881,N_49470,N_49458);
xnor U49882 (N_49882,N_49294,N_49348);
nor U49883 (N_49883,N_49308,N_49194);
or U49884 (N_49884,N_49143,N_49098);
nand U49885 (N_49885,N_49461,N_49183);
and U49886 (N_49886,N_49258,N_49324);
nor U49887 (N_49887,N_49345,N_49052);
and U49888 (N_49888,N_49179,N_49436);
and U49889 (N_49889,N_49376,N_49193);
nand U49890 (N_49890,N_49451,N_49387);
nand U49891 (N_49891,N_49066,N_49430);
or U49892 (N_49892,N_49222,N_49287);
and U49893 (N_49893,N_49166,N_49114);
nor U49894 (N_49894,N_49494,N_49163);
or U49895 (N_49895,N_49095,N_49387);
nor U49896 (N_49896,N_49282,N_49459);
nand U49897 (N_49897,N_49244,N_49489);
xor U49898 (N_49898,N_49449,N_49448);
xor U49899 (N_49899,N_49072,N_49474);
and U49900 (N_49900,N_49136,N_49299);
nand U49901 (N_49901,N_49425,N_49075);
and U49902 (N_49902,N_49230,N_49173);
nor U49903 (N_49903,N_49343,N_49368);
or U49904 (N_49904,N_49280,N_49486);
or U49905 (N_49905,N_49028,N_49254);
or U49906 (N_49906,N_49183,N_49388);
xor U49907 (N_49907,N_49150,N_49488);
nand U49908 (N_49908,N_49046,N_49053);
or U49909 (N_49909,N_49123,N_49207);
nor U49910 (N_49910,N_49280,N_49169);
nor U49911 (N_49911,N_49142,N_49473);
nand U49912 (N_49912,N_49130,N_49358);
nor U49913 (N_49913,N_49165,N_49277);
and U49914 (N_49914,N_49345,N_49089);
nor U49915 (N_49915,N_49328,N_49286);
and U49916 (N_49916,N_49412,N_49037);
nand U49917 (N_49917,N_49056,N_49190);
and U49918 (N_49918,N_49018,N_49399);
nor U49919 (N_49919,N_49184,N_49492);
or U49920 (N_49920,N_49264,N_49181);
nor U49921 (N_49921,N_49476,N_49372);
nand U49922 (N_49922,N_49144,N_49089);
nand U49923 (N_49923,N_49211,N_49017);
and U49924 (N_49924,N_49286,N_49200);
and U49925 (N_49925,N_49228,N_49434);
nand U49926 (N_49926,N_49165,N_49088);
nor U49927 (N_49927,N_49271,N_49160);
and U49928 (N_49928,N_49323,N_49029);
nor U49929 (N_49929,N_49281,N_49150);
or U49930 (N_49930,N_49204,N_49299);
xor U49931 (N_49931,N_49076,N_49144);
and U49932 (N_49932,N_49149,N_49010);
and U49933 (N_49933,N_49075,N_49201);
nor U49934 (N_49934,N_49321,N_49262);
and U49935 (N_49935,N_49478,N_49080);
and U49936 (N_49936,N_49171,N_49061);
or U49937 (N_49937,N_49273,N_49157);
nand U49938 (N_49938,N_49117,N_49448);
or U49939 (N_49939,N_49316,N_49278);
nand U49940 (N_49940,N_49243,N_49374);
or U49941 (N_49941,N_49333,N_49496);
nor U49942 (N_49942,N_49261,N_49112);
or U49943 (N_49943,N_49004,N_49193);
nor U49944 (N_49944,N_49439,N_49023);
or U49945 (N_49945,N_49369,N_49080);
nand U49946 (N_49946,N_49033,N_49220);
or U49947 (N_49947,N_49256,N_49462);
or U49948 (N_49948,N_49105,N_49246);
nor U49949 (N_49949,N_49481,N_49359);
or U49950 (N_49950,N_49069,N_49238);
and U49951 (N_49951,N_49446,N_49448);
and U49952 (N_49952,N_49419,N_49474);
and U49953 (N_49953,N_49308,N_49367);
and U49954 (N_49954,N_49336,N_49376);
nor U49955 (N_49955,N_49194,N_49190);
or U49956 (N_49956,N_49407,N_49139);
or U49957 (N_49957,N_49153,N_49234);
nand U49958 (N_49958,N_49092,N_49426);
and U49959 (N_49959,N_49455,N_49466);
or U49960 (N_49960,N_49171,N_49021);
and U49961 (N_49961,N_49209,N_49336);
or U49962 (N_49962,N_49211,N_49388);
nor U49963 (N_49963,N_49416,N_49075);
or U49964 (N_49964,N_49401,N_49116);
and U49965 (N_49965,N_49088,N_49243);
nor U49966 (N_49966,N_49391,N_49037);
nor U49967 (N_49967,N_49481,N_49317);
xor U49968 (N_49968,N_49372,N_49239);
nand U49969 (N_49969,N_49130,N_49337);
xnor U49970 (N_49970,N_49009,N_49409);
and U49971 (N_49971,N_49151,N_49218);
and U49972 (N_49972,N_49332,N_49256);
or U49973 (N_49973,N_49493,N_49468);
or U49974 (N_49974,N_49129,N_49259);
or U49975 (N_49975,N_49157,N_49297);
nand U49976 (N_49976,N_49396,N_49071);
and U49977 (N_49977,N_49257,N_49263);
nor U49978 (N_49978,N_49348,N_49327);
nor U49979 (N_49979,N_49066,N_49473);
nand U49980 (N_49980,N_49282,N_49434);
or U49981 (N_49981,N_49144,N_49340);
and U49982 (N_49982,N_49091,N_49376);
and U49983 (N_49983,N_49162,N_49371);
nor U49984 (N_49984,N_49391,N_49097);
nor U49985 (N_49985,N_49083,N_49305);
xor U49986 (N_49986,N_49216,N_49066);
nor U49987 (N_49987,N_49064,N_49353);
nor U49988 (N_49988,N_49180,N_49493);
nand U49989 (N_49989,N_49392,N_49316);
or U49990 (N_49990,N_49191,N_49028);
and U49991 (N_49991,N_49348,N_49324);
nor U49992 (N_49992,N_49462,N_49307);
and U49993 (N_49993,N_49467,N_49086);
nand U49994 (N_49994,N_49485,N_49179);
or U49995 (N_49995,N_49334,N_49042);
nor U49996 (N_49996,N_49424,N_49005);
or U49997 (N_49997,N_49076,N_49131);
and U49998 (N_49998,N_49178,N_49295);
and U49999 (N_49999,N_49351,N_49323);
xnor UO_0 (O_0,N_49686,N_49739);
nor UO_1 (O_1,N_49526,N_49761);
nor UO_2 (O_2,N_49816,N_49942);
or UO_3 (O_3,N_49852,N_49784);
nor UO_4 (O_4,N_49898,N_49648);
xor UO_5 (O_5,N_49675,N_49943);
nor UO_6 (O_6,N_49862,N_49902);
xor UO_7 (O_7,N_49732,N_49996);
nand UO_8 (O_8,N_49820,N_49983);
nor UO_9 (O_9,N_49651,N_49554);
or UO_10 (O_10,N_49661,N_49896);
nand UO_11 (O_11,N_49581,N_49792);
and UO_12 (O_12,N_49873,N_49745);
or UO_13 (O_13,N_49850,N_49580);
and UO_14 (O_14,N_49855,N_49975);
nand UO_15 (O_15,N_49876,N_49595);
nand UO_16 (O_16,N_49821,N_49640);
nand UO_17 (O_17,N_49625,N_49921);
nor UO_18 (O_18,N_49712,N_49796);
and UO_19 (O_19,N_49813,N_49513);
or UO_20 (O_20,N_49673,N_49683);
xnor UO_21 (O_21,N_49729,N_49946);
nand UO_22 (O_22,N_49711,N_49805);
nand UO_23 (O_23,N_49629,N_49658);
xor UO_24 (O_24,N_49609,N_49924);
or UO_25 (O_25,N_49841,N_49857);
or UO_26 (O_26,N_49970,N_49905);
or UO_27 (O_27,N_49716,N_49984);
xnor UO_28 (O_28,N_49824,N_49529);
xnor UO_29 (O_29,N_49897,N_49669);
nand UO_30 (O_30,N_49659,N_49626);
nor UO_31 (O_31,N_49551,N_49537);
nand UO_32 (O_32,N_49746,N_49516);
nor UO_33 (O_33,N_49934,N_49822);
or UO_34 (O_34,N_49586,N_49724);
nor UO_35 (O_35,N_49919,N_49999);
or UO_36 (O_36,N_49622,N_49961);
xor UO_37 (O_37,N_49515,N_49639);
and UO_38 (O_38,N_49915,N_49688);
and UO_39 (O_39,N_49657,N_49735);
or UO_40 (O_40,N_49869,N_49979);
and UO_41 (O_41,N_49684,N_49590);
nand UO_42 (O_42,N_49974,N_49593);
nand UO_43 (O_43,N_49742,N_49570);
xor UO_44 (O_44,N_49730,N_49765);
nor UO_45 (O_45,N_49604,N_49885);
and UO_46 (O_46,N_49705,N_49619);
nor UO_47 (O_47,N_49932,N_49553);
and UO_48 (O_48,N_49685,N_49965);
nand UO_49 (O_49,N_49632,N_49534);
nor UO_50 (O_50,N_49879,N_49546);
and UO_51 (O_51,N_49752,N_49717);
nor UO_52 (O_52,N_49738,N_49891);
and UO_53 (O_53,N_49702,N_49759);
nand UO_54 (O_54,N_49678,N_49696);
or UO_55 (O_55,N_49720,N_49571);
and UO_56 (O_56,N_49769,N_49789);
or UO_57 (O_57,N_49587,N_49680);
nor UO_58 (O_58,N_49670,N_49950);
nand UO_59 (O_59,N_49653,N_49887);
and UO_60 (O_60,N_49621,N_49874);
nand UO_61 (O_61,N_49788,N_49505);
and UO_62 (O_62,N_49731,N_49888);
xor UO_63 (O_63,N_49875,N_49848);
or UO_64 (O_64,N_49517,N_49886);
nand UO_65 (O_65,N_49694,N_49592);
nor UO_66 (O_66,N_49695,N_49901);
or UO_67 (O_67,N_49851,N_49804);
or UO_68 (O_68,N_49504,N_49636);
nor UO_69 (O_69,N_49785,N_49995);
or UO_70 (O_70,N_49584,N_49960);
xnor UO_71 (O_71,N_49849,N_49906);
or UO_72 (O_72,N_49650,N_49681);
or UO_73 (O_73,N_49531,N_49642);
or UO_74 (O_74,N_49550,N_49925);
or UO_75 (O_75,N_49547,N_49687);
or UO_76 (O_76,N_49986,N_49613);
and UO_77 (O_77,N_49579,N_49972);
nand UO_78 (O_78,N_49677,N_49598);
and UO_79 (O_79,N_49741,N_49819);
xor UO_80 (O_80,N_49519,N_49956);
xor UO_81 (O_81,N_49935,N_49698);
nand UO_82 (O_82,N_49842,N_49647);
nor UO_83 (O_83,N_49985,N_49889);
nor UO_84 (O_84,N_49556,N_49962);
or UO_85 (O_85,N_49572,N_49542);
nand UO_86 (O_86,N_49706,N_49558);
nor UO_87 (O_87,N_49544,N_49603);
nand UO_88 (O_88,N_49564,N_49952);
or UO_89 (O_89,N_49778,N_49917);
nor UO_90 (O_90,N_49583,N_49870);
or UO_91 (O_91,N_49908,N_49797);
or UO_92 (O_92,N_49700,N_49839);
nor UO_93 (O_93,N_49866,N_49922);
nor UO_94 (O_94,N_49633,N_49576);
nand UO_95 (O_95,N_49528,N_49777);
or UO_96 (O_96,N_49566,N_49682);
or UO_97 (O_97,N_49998,N_49944);
and UO_98 (O_98,N_49780,N_49760);
or UO_99 (O_99,N_49913,N_49541);
and UO_100 (O_100,N_49568,N_49545);
and UO_101 (O_101,N_49988,N_49623);
nor UO_102 (O_102,N_49693,N_49617);
and UO_103 (O_103,N_49666,N_49817);
and UO_104 (O_104,N_49563,N_49993);
and UO_105 (O_105,N_49614,N_49881);
and UO_106 (O_106,N_49606,N_49781);
nand UO_107 (O_107,N_49751,N_49691);
nand UO_108 (O_108,N_49854,N_49522);
or UO_109 (O_109,N_49802,N_49575);
nor UO_110 (O_110,N_49722,N_49864);
nor UO_111 (O_111,N_49643,N_49527);
nor UO_112 (O_112,N_49912,N_49937);
or UO_113 (O_113,N_49540,N_49747);
nor UO_114 (O_114,N_49939,N_49786);
nand UO_115 (O_115,N_49882,N_49872);
and UO_116 (O_116,N_49818,N_49782);
and UO_117 (O_117,N_49708,N_49612);
or UO_118 (O_118,N_49749,N_49790);
or UO_119 (O_119,N_49968,N_49811);
nor UO_120 (O_120,N_49800,N_49689);
nor UO_121 (O_121,N_49883,N_49903);
xor UO_122 (O_122,N_49667,N_49524);
nor UO_123 (O_123,N_49721,N_49826);
and UO_124 (O_124,N_49941,N_49899);
and UO_125 (O_125,N_49930,N_49837);
xnor UO_126 (O_126,N_49649,N_49577);
and UO_127 (O_127,N_49798,N_49674);
nand UO_128 (O_128,N_49668,N_49753);
and UO_129 (O_129,N_49871,N_49562);
nor UO_130 (O_130,N_49940,N_49947);
nand UO_131 (O_131,N_49815,N_49585);
nor UO_132 (O_132,N_49861,N_49763);
nand UO_133 (O_133,N_49825,N_49949);
xnor UO_134 (O_134,N_49840,N_49920);
nand UO_135 (O_135,N_49884,N_49699);
xnor UO_136 (O_136,N_49665,N_49980);
xor UO_137 (O_137,N_49801,N_49518);
nand UO_138 (O_138,N_49863,N_49890);
nor UO_139 (O_139,N_49756,N_49503);
nor UO_140 (O_140,N_49757,N_49823);
or UO_141 (O_141,N_49827,N_49836);
nand UO_142 (O_142,N_49601,N_49966);
nand UO_143 (O_143,N_49954,N_49525);
and UO_144 (O_144,N_49953,N_49904);
and UO_145 (O_145,N_49914,N_49624);
or UO_146 (O_146,N_49588,N_49548);
nor UO_147 (O_147,N_49755,N_49536);
or UO_148 (O_148,N_49710,N_49832);
nand UO_149 (O_149,N_49814,N_49559);
and UO_150 (O_150,N_49725,N_49766);
and UO_151 (O_151,N_49707,N_49557);
nand UO_152 (O_152,N_49654,N_49877);
xor UO_153 (O_153,N_49918,N_49631);
or UO_154 (O_154,N_49641,N_49715);
and UO_155 (O_155,N_49634,N_49690);
and UO_156 (O_156,N_49552,N_49646);
or UO_157 (O_157,N_49977,N_49560);
nor UO_158 (O_158,N_49845,N_49701);
nand UO_159 (O_159,N_49771,N_49533);
or UO_160 (O_160,N_49971,N_49511);
nand UO_161 (O_161,N_49602,N_49521);
or UO_162 (O_162,N_49847,N_49795);
or UO_163 (O_163,N_49713,N_49997);
or UO_164 (O_164,N_49726,N_49867);
or UO_165 (O_165,N_49990,N_49958);
nor UO_166 (O_166,N_49762,N_49933);
nor UO_167 (O_167,N_49500,N_49768);
or UO_168 (O_168,N_49793,N_49714);
nand UO_169 (O_169,N_49514,N_49978);
and UO_170 (O_170,N_49509,N_49502);
and UO_171 (O_171,N_49736,N_49697);
and UO_172 (O_172,N_49645,N_49573);
nand UO_173 (O_173,N_49892,N_49574);
nand UO_174 (O_174,N_49600,N_49737);
or UO_175 (O_175,N_49565,N_49843);
and UO_176 (O_176,N_49754,N_49868);
and UO_177 (O_177,N_49994,N_49909);
nand UO_178 (O_178,N_49549,N_49808);
and UO_179 (O_179,N_49963,N_49964);
nor UO_180 (O_180,N_49679,N_49703);
nor UO_181 (O_181,N_49894,N_49638);
and UO_182 (O_182,N_49510,N_49567);
xnor UO_183 (O_183,N_49628,N_49858);
or UO_184 (O_184,N_49607,N_49829);
nand UO_185 (O_185,N_49671,N_49779);
or UO_186 (O_186,N_49676,N_49809);
and UO_187 (O_187,N_49794,N_49938);
xor UO_188 (O_188,N_49538,N_49927);
nor UO_189 (O_189,N_49926,N_49608);
and UO_190 (O_190,N_49856,N_49512);
nor UO_191 (O_191,N_49589,N_49611);
nor UO_192 (O_192,N_49728,N_49615);
nor UO_193 (O_193,N_49652,N_49991);
or UO_194 (O_194,N_49507,N_49539);
nor UO_195 (O_195,N_49893,N_49772);
nor UO_196 (O_196,N_49764,N_49773);
xor UO_197 (O_197,N_49969,N_49535);
nor UO_198 (O_198,N_49561,N_49791);
nor UO_199 (O_199,N_49618,N_49846);
nand UO_200 (O_200,N_49709,N_49929);
xnor UO_201 (O_201,N_49838,N_49506);
nor UO_202 (O_202,N_49835,N_49959);
nor UO_203 (O_203,N_49627,N_49767);
nand UO_204 (O_204,N_49770,N_49532);
nor UO_205 (O_205,N_49758,N_49931);
nand UO_206 (O_206,N_49723,N_49644);
and UO_207 (O_207,N_49594,N_49981);
nand UO_208 (O_208,N_49973,N_49923);
and UO_209 (O_209,N_49704,N_49555);
and UO_210 (O_210,N_49945,N_49895);
xnor UO_211 (O_211,N_49880,N_49637);
nor UO_212 (O_212,N_49989,N_49812);
nor UO_213 (O_213,N_49803,N_49967);
or UO_214 (O_214,N_49834,N_49630);
nor UO_215 (O_215,N_49976,N_49810);
or UO_216 (O_216,N_49692,N_49597);
and UO_217 (O_217,N_49663,N_49900);
and UO_218 (O_218,N_49774,N_49596);
nand UO_219 (O_219,N_49928,N_49740);
and UO_220 (O_220,N_49748,N_49907);
or UO_221 (O_221,N_49936,N_49955);
nor UO_222 (O_222,N_49806,N_49616);
nor UO_223 (O_223,N_49656,N_49520);
nor UO_224 (O_224,N_49582,N_49733);
nand UO_225 (O_225,N_49775,N_49718);
and UO_226 (O_226,N_49578,N_49865);
or UO_227 (O_227,N_49992,N_49776);
nand UO_228 (O_228,N_49635,N_49655);
nand UO_229 (O_229,N_49844,N_49916);
and UO_230 (O_230,N_49591,N_49599);
and UO_231 (O_231,N_49951,N_49830);
and UO_232 (O_232,N_49987,N_49605);
nor UO_233 (O_233,N_49727,N_49744);
or UO_234 (O_234,N_49982,N_49543);
nor UO_235 (O_235,N_49660,N_49828);
xnor UO_236 (O_236,N_49787,N_49878);
and UO_237 (O_237,N_49853,N_49833);
and UO_238 (O_238,N_49750,N_49664);
and UO_239 (O_239,N_49569,N_49743);
or UO_240 (O_240,N_49807,N_49719);
or UO_241 (O_241,N_49610,N_49799);
or UO_242 (O_242,N_49530,N_49948);
and UO_243 (O_243,N_49831,N_49783);
nor UO_244 (O_244,N_49910,N_49911);
or UO_245 (O_245,N_49672,N_49860);
xnor UO_246 (O_246,N_49662,N_49508);
and UO_247 (O_247,N_49523,N_49734);
or UO_248 (O_248,N_49859,N_49957);
and UO_249 (O_249,N_49501,N_49620);
nand UO_250 (O_250,N_49755,N_49613);
nor UO_251 (O_251,N_49829,N_49765);
or UO_252 (O_252,N_49561,N_49511);
and UO_253 (O_253,N_49786,N_49782);
nand UO_254 (O_254,N_49614,N_49739);
and UO_255 (O_255,N_49809,N_49743);
or UO_256 (O_256,N_49656,N_49914);
or UO_257 (O_257,N_49695,N_49871);
xor UO_258 (O_258,N_49574,N_49968);
nor UO_259 (O_259,N_49697,N_49533);
nor UO_260 (O_260,N_49925,N_49830);
or UO_261 (O_261,N_49669,N_49691);
nand UO_262 (O_262,N_49886,N_49898);
or UO_263 (O_263,N_49831,N_49515);
nor UO_264 (O_264,N_49961,N_49656);
nand UO_265 (O_265,N_49862,N_49810);
xnor UO_266 (O_266,N_49935,N_49778);
or UO_267 (O_267,N_49692,N_49655);
nor UO_268 (O_268,N_49521,N_49804);
or UO_269 (O_269,N_49500,N_49621);
nor UO_270 (O_270,N_49543,N_49569);
nor UO_271 (O_271,N_49826,N_49529);
nor UO_272 (O_272,N_49734,N_49639);
nand UO_273 (O_273,N_49911,N_49979);
xor UO_274 (O_274,N_49677,N_49881);
nand UO_275 (O_275,N_49987,N_49917);
nor UO_276 (O_276,N_49720,N_49603);
and UO_277 (O_277,N_49976,N_49670);
xor UO_278 (O_278,N_49879,N_49774);
or UO_279 (O_279,N_49521,N_49588);
or UO_280 (O_280,N_49950,N_49730);
or UO_281 (O_281,N_49942,N_49660);
or UO_282 (O_282,N_49744,N_49510);
or UO_283 (O_283,N_49578,N_49689);
nand UO_284 (O_284,N_49672,N_49798);
and UO_285 (O_285,N_49956,N_49827);
xnor UO_286 (O_286,N_49627,N_49788);
nor UO_287 (O_287,N_49947,N_49859);
nor UO_288 (O_288,N_49689,N_49946);
nor UO_289 (O_289,N_49637,N_49825);
nand UO_290 (O_290,N_49815,N_49616);
and UO_291 (O_291,N_49714,N_49859);
or UO_292 (O_292,N_49836,N_49859);
nand UO_293 (O_293,N_49906,N_49613);
nand UO_294 (O_294,N_49827,N_49579);
xor UO_295 (O_295,N_49916,N_49843);
nor UO_296 (O_296,N_49760,N_49746);
or UO_297 (O_297,N_49751,N_49657);
nor UO_298 (O_298,N_49939,N_49971);
nand UO_299 (O_299,N_49759,N_49692);
nand UO_300 (O_300,N_49606,N_49753);
nand UO_301 (O_301,N_49809,N_49841);
and UO_302 (O_302,N_49708,N_49663);
or UO_303 (O_303,N_49888,N_49622);
or UO_304 (O_304,N_49809,N_49501);
and UO_305 (O_305,N_49735,N_49995);
nand UO_306 (O_306,N_49951,N_49869);
xor UO_307 (O_307,N_49660,N_49744);
nand UO_308 (O_308,N_49914,N_49661);
and UO_309 (O_309,N_49775,N_49724);
and UO_310 (O_310,N_49995,N_49923);
and UO_311 (O_311,N_49941,N_49980);
or UO_312 (O_312,N_49859,N_49619);
nor UO_313 (O_313,N_49604,N_49948);
xnor UO_314 (O_314,N_49677,N_49581);
or UO_315 (O_315,N_49939,N_49914);
nor UO_316 (O_316,N_49815,N_49572);
xnor UO_317 (O_317,N_49540,N_49953);
nor UO_318 (O_318,N_49738,N_49639);
nand UO_319 (O_319,N_49510,N_49787);
and UO_320 (O_320,N_49522,N_49784);
nor UO_321 (O_321,N_49724,N_49739);
or UO_322 (O_322,N_49682,N_49802);
or UO_323 (O_323,N_49519,N_49670);
nand UO_324 (O_324,N_49796,N_49551);
nand UO_325 (O_325,N_49913,N_49801);
nor UO_326 (O_326,N_49595,N_49970);
and UO_327 (O_327,N_49706,N_49634);
or UO_328 (O_328,N_49770,N_49801);
and UO_329 (O_329,N_49825,N_49686);
and UO_330 (O_330,N_49705,N_49874);
or UO_331 (O_331,N_49686,N_49922);
xor UO_332 (O_332,N_49563,N_49768);
and UO_333 (O_333,N_49708,N_49807);
and UO_334 (O_334,N_49640,N_49552);
or UO_335 (O_335,N_49706,N_49575);
or UO_336 (O_336,N_49507,N_49710);
nand UO_337 (O_337,N_49630,N_49843);
or UO_338 (O_338,N_49731,N_49590);
nor UO_339 (O_339,N_49727,N_49643);
and UO_340 (O_340,N_49519,N_49936);
or UO_341 (O_341,N_49935,N_49879);
nand UO_342 (O_342,N_49810,N_49540);
and UO_343 (O_343,N_49558,N_49571);
nand UO_344 (O_344,N_49655,N_49511);
and UO_345 (O_345,N_49594,N_49921);
and UO_346 (O_346,N_49965,N_49834);
or UO_347 (O_347,N_49918,N_49687);
xnor UO_348 (O_348,N_49973,N_49843);
and UO_349 (O_349,N_49701,N_49702);
nand UO_350 (O_350,N_49752,N_49694);
or UO_351 (O_351,N_49564,N_49735);
nor UO_352 (O_352,N_49841,N_49991);
nor UO_353 (O_353,N_49686,N_49845);
xor UO_354 (O_354,N_49704,N_49518);
nand UO_355 (O_355,N_49718,N_49561);
and UO_356 (O_356,N_49637,N_49561);
nand UO_357 (O_357,N_49741,N_49822);
or UO_358 (O_358,N_49871,N_49687);
nand UO_359 (O_359,N_49679,N_49678);
or UO_360 (O_360,N_49552,N_49970);
or UO_361 (O_361,N_49973,N_49665);
nand UO_362 (O_362,N_49673,N_49640);
nand UO_363 (O_363,N_49946,N_49645);
and UO_364 (O_364,N_49686,N_49694);
nand UO_365 (O_365,N_49738,N_49588);
or UO_366 (O_366,N_49647,N_49765);
or UO_367 (O_367,N_49527,N_49869);
nand UO_368 (O_368,N_49818,N_49669);
nand UO_369 (O_369,N_49631,N_49500);
nand UO_370 (O_370,N_49514,N_49857);
and UO_371 (O_371,N_49530,N_49588);
nor UO_372 (O_372,N_49833,N_49917);
nor UO_373 (O_373,N_49808,N_49636);
nor UO_374 (O_374,N_49908,N_49508);
and UO_375 (O_375,N_49840,N_49570);
or UO_376 (O_376,N_49945,N_49707);
or UO_377 (O_377,N_49876,N_49603);
and UO_378 (O_378,N_49599,N_49909);
nand UO_379 (O_379,N_49907,N_49970);
nand UO_380 (O_380,N_49834,N_49918);
and UO_381 (O_381,N_49551,N_49744);
or UO_382 (O_382,N_49642,N_49814);
nor UO_383 (O_383,N_49678,N_49756);
or UO_384 (O_384,N_49762,N_49819);
or UO_385 (O_385,N_49836,N_49595);
or UO_386 (O_386,N_49622,N_49545);
or UO_387 (O_387,N_49895,N_49642);
nand UO_388 (O_388,N_49737,N_49955);
or UO_389 (O_389,N_49510,N_49866);
or UO_390 (O_390,N_49925,N_49670);
nand UO_391 (O_391,N_49850,N_49886);
and UO_392 (O_392,N_49664,N_49566);
or UO_393 (O_393,N_49905,N_49793);
and UO_394 (O_394,N_49605,N_49573);
xor UO_395 (O_395,N_49897,N_49558);
or UO_396 (O_396,N_49696,N_49764);
nor UO_397 (O_397,N_49949,N_49942);
nand UO_398 (O_398,N_49518,N_49515);
and UO_399 (O_399,N_49905,N_49610);
or UO_400 (O_400,N_49691,N_49775);
xnor UO_401 (O_401,N_49933,N_49895);
nor UO_402 (O_402,N_49573,N_49600);
or UO_403 (O_403,N_49813,N_49832);
nor UO_404 (O_404,N_49632,N_49561);
nor UO_405 (O_405,N_49621,N_49632);
nand UO_406 (O_406,N_49593,N_49738);
or UO_407 (O_407,N_49794,N_49733);
and UO_408 (O_408,N_49823,N_49993);
or UO_409 (O_409,N_49611,N_49576);
or UO_410 (O_410,N_49652,N_49752);
nor UO_411 (O_411,N_49513,N_49805);
xor UO_412 (O_412,N_49577,N_49835);
or UO_413 (O_413,N_49928,N_49723);
nor UO_414 (O_414,N_49553,N_49587);
nand UO_415 (O_415,N_49638,N_49566);
nor UO_416 (O_416,N_49694,N_49504);
or UO_417 (O_417,N_49500,N_49706);
nor UO_418 (O_418,N_49964,N_49981);
nand UO_419 (O_419,N_49971,N_49567);
nor UO_420 (O_420,N_49778,N_49775);
and UO_421 (O_421,N_49530,N_49965);
nor UO_422 (O_422,N_49537,N_49657);
nor UO_423 (O_423,N_49797,N_49696);
nand UO_424 (O_424,N_49981,N_49986);
xor UO_425 (O_425,N_49970,N_49715);
or UO_426 (O_426,N_49578,N_49875);
nand UO_427 (O_427,N_49839,N_49879);
and UO_428 (O_428,N_49584,N_49700);
nor UO_429 (O_429,N_49576,N_49910);
nor UO_430 (O_430,N_49912,N_49538);
and UO_431 (O_431,N_49885,N_49982);
nor UO_432 (O_432,N_49519,N_49827);
and UO_433 (O_433,N_49697,N_49584);
or UO_434 (O_434,N_49745,N_49741);
or UO_435 (O_435,N_49749,N_49761);
nor UO_436 (O_436,N_49560,N_49799);
xor UO_437 (O_437,N_49575,N_49646);
xnor UO_438 (O_438,N_49652,N_49548);
nand UO_439 (O_439,N_49763,N_49715);
xor UO_440 (O_440,N_49929,N_49504);
nand UO_441 (O_441,N_49611,N_49503);
or UO_442 (O_442,N_49722,N_49845);
xor UO_443 (O_443,N_49888,N_49738);
or UO_444 (O_444,N_49580,N_49513);
or UO_445 (O_445,N_49753,N_49927);
and UO_446 (O_446,N_49853,N_49882);
or UO_447 (O_447,N_49809,N_49854);
nor UO_448 (O_448,N_49510,N_49583);
nand UO_449 (O_449,N_49956,N_49515);
nor UO_450 (O_450,N_49591,N_49797);
and UO_451 (O_451,N_49752,N_49936);
nand UO_452 (O_452,N_49819,N_49715);
nor UO_453 (O_453,N_49992,N_49699);
nand UO_454 (O_454,N_49869,N_49728);
or UO_455 (O_455,N_49724,N_49879);
nor UO_456 (O_456,N_49979,N_49784);
nand UO_457 (O_457,N_49955,N_49689);
nor UO_458 (O_458,N_49595,N_49797);
and UO_459 (O_459,N_49776,N_49822);
nand UO_460 (O_460,N_49947,N_49952);
nor UO_461 (O_461,N_49715,N_49638);
and UO_462 (O_462,N_49896,N_49698);
or UO_463 (O_463,N_49711,N_49674);
nand UO_464 (O_464,N_49966,N_49746);
nor UO_465 (O_465,N_49632,N_49826);
or UO_466 (O_466,N_49536,N_49998);
nand UO_467 (O_467,N_49521,N_49552);
nand UO_468 (O_468,N_49921,N_49909);
nor UO_469 (O_469,N_49978,N_49525);
nand UO_470 (O_470,N_49687,N_49998);
nand UO_471 (O_471,N_49754,N_49629);
nand UO_472 (O_472,N_49900,N_49810);
nor UO_473 (O_473,N_49540,N_49668);
nor UO_474 (O_474,N_49666,N_49807);
and UO_475 (O_475,N_49760,N_49789);
nor UO_476 (O_476,N_49597,N_49795);
nand UO_477 (O_477,N_49686,N_49695);
nand UO_478 (O_478,N_49773,N_49871);
or UO_479 (O_479,N_49917,N_49895);
nor UO_480 (O_480,N_49649,N_49501);
nand UO_481 (O_481,N_49642,N_49691);
nor UO_482 (O_482,N_49817,N_49598);
or UO_483 (O_483,N_49619,N_49900);
and UO_484 (O_484,N_49763,N_49981);
or UO_485 (O_485,N_49543,N_49984);
nor UO_486 (O_486,N_49522,N_49729);
and UO_487 (O_487,N_49786,N_49716);
nand UO_488 (O_488,N_49807,N_49846);
and UO_489 (O_489,N_49931,N_49774);
xor UO_490 (O_490,N_49602,N_49901);
nor UO_491 (O_491,N_49951,N_49870);
nand UO_492 (O_492,N_49991,N_49889);
and UO_493 (O_493,N_49827,N_49784);
nand UO_494 (O_494,N_49900,N_49517);
and UO_495 (O_495,N_49906,N_49945);
or UO_496 (O_496,N_49825,N_49533);
or UO_497 (O_497,N_49983,N_49773);
xnor UO_498 (O_498,N_49595,N_49968);
and UO_499 (O_499,N_49837,N_49980);
nand UO_500 (O_500,N_49791,N_49622);
nand UO_501 (O_501,N_49564,N_49986);
and UO_502 (O_502,N_49843,N_49831);
or UO_503 (O_503,N_49885,N_49892);
nor UO_504 (O_504,N_49959,N_49661);
nand UO_505 (O_505,N_49799,N_49875);
or UO_506 (O_506,N_49771,N_49913);
xor UO_507 (O_507,N_49553,N_49541);
nand UO_508 (O_508,N_49889,N_49970);
and UO_509 (O_509,N_49822,N_49989);
and UO_510 (O_510,N_49651,N_49650);
and UO_511 (O_511,N_49926,N_49839);
or UO_512 (O_512,N_49530,N_49904);
nor UO_513 (O_513,N_49804,N_49545);
or UO_514 (O_514,N_49870,N_49721);
and UO_515 (O_515,N_49850,N_49767);
or UO_516 (O_516,N_49762,N_49735);
nor UO_517 (O_517,N_49782,N_49769);
nand UO_518 (O_518,N_49720,N_49751);
xor UO_519 (O_519,N_49520,N_49650);
nor UO_520 (O_520,N_49706,N_49893);
nor UO_521 (O_521,N_49537,N_49815);
xnor UO_522 (O_522,N_49748,N_49729);
and UO_523 (O_523,N_49866,N_49544);
and UO_524 (O_524,N_49541,N_49642);
nand UO_525 (O_525,N_49746,N_49588);
and UO_526 (O_526,N_49950,N_49741);
nand UO_527 (O_527,N_49502,N_49946);
nand UO_528 (O_528,N_49873,N_49697);
nor UO_529 (O_529,N_49730,N_49760);
or UO_530 (O_530,N_49747,N_49767);
xor UO_531 (O_531,N_49788,N_49513);
xor UO_532 (O_532,N_49597,N_49814);
and UO_533 (O_533,N_49935,N_49838);
nand UO_534 (O_534,N_49898,N_49759);
and UO_535 (O_535,N_49668,N_49617);
xnor UO_536 (O_536,N_49924,N_49828);
or UO_537 (O_537,N_49877,N_49758);
nand UO_538 (O_538,N_49901,N_49821);
and UO_539 (O_539,N_49777,N_49597);
or UO_540 (O_540,N_49579,N_49782);
or UO_541 (O_541,N_49695,N_49739);
nand UO_542 (O_542,N_49528,N_49815);
nand UO_543 (O_543,N_49816,N_49675);
nand UO_544 (O_544,N_49919,N_49712);
xnor UO_545 (O_545,N_49776,N_49560);
nand UO_546 (O_546,N_49694,N_49501);
and UO_547 (O_547,N_49716,N_49919);
and UO_548 (O_548,N_49848,N_49701);
and UO_549 (O_549,N_49900,N_49826);
and UO_550 (O_550,N_49730,N_49957);
nor UO_551 (O_551,N_49756,N_49696);
nor UO_552 (O_552,N_49754,N_49526);
nor UO_553 (O_553,N_49798,N_49665);
nand UO_554 (O_554,N_49579,N_49973);
or UO_555 (O_555,N_49796,N_49841);
xor UO_556 (O_556,N_49672,N_49974);
or UO_557 (O_557,N_49548,N_49741);
and UO_558 (O_558,N_49832,N_49903);
or UO_559 (O_559,N_49650,N_49707);
and UO_560 (O_560,N_49738,N_49992);
xor UO_561 (O_561,N_49556,N_49533);
or UO_562 (O_562,N_49832,N_49932);
nand UO_563 (O_563,N_49790,N_49584);
and UO_564 (O_564,N_49726,N_49743);
xnor UO_565 (O_565,N_49749,N_49843);
nor UO_566 (O_566,N_49841,N_49675);
and UO_567 (O_567,N_49957,N_49793);
nor UO_568 (O_568,N_49547,N_49919);
nand UO_569 (O_569,N_49828,N_49948);
xor UO_570 (O_570,N_49984,N_49757);
nor UO_571 (O_571,N_49761,N_49759);
and UO_572 (O_572,N_49663,N_49510);
nand UO_573 (O_573,N_49673,N_49601);
or UO_574 (O_574,N_49723,N_49523);
nand UO_575 (O_575,N_49756,N_49670);
and UO_576 (O_576,N_49508,N_49625);
and UO_577 (O_577,N_49596,N_49783);
and UO_578 (O_578,N_49857,N_49744);
or UO_579 (O_579,N_49515,N_49767);
nand UO_580 (O_580,N_49796,N_49768);
nor UO_581 (O_581,N_49959,N_49632);
nand UO_582 (O_582,N_49508,N_49527);
and UO_583 (O_583,N_49586,N_49585);
and UO_584 (O_584,N_49504,N_49785);
nand UO_585 (O_585,N_49850,N_49650);
nand UO_586 (O_586,N_49502,N_49912);
or UO_587 (O_587,N_49669,N_49511);
nor UO_588 (O_588,N_49757,N_49873);
nor UO_589 (O_589,N_49753,N_49892);
nand UO_590 (O_590,N_49657,N_49578);
or UO_591 (O_591,N_49829,N_49548);
and UO_592 (O_592,N_49762,N_49752);
nand UO_593 (O_593,N_49971,N_49877);
and UO_594 (O_594,N_49641,N_49663);
or UO_595 (O_595,N_49701,N_49834);
or UO_596 (O_596,N_49585,N_49985);
nor UO_597 (O_597,N_49921,N_49723);
nor UO_598 (O_598,N_49865,N_49846);
or UO_599 (O_599,N_49666,N_49716);
nor UO_600 (O_600,N_49589,N_49691);
xor UO_601 (O_601,N_49972,N_49757);
nand UO_602 (O_602,N_49886,N_49935);
nand UO_603 (O_603,N_49970,N_49657);
xor UO_604 (O_604,N_49523,N_49757);
or UO_605 (O_605,N_49838,N_49954);
nand UO_606 (O_606,N_49502,N_49723);
nand UO_607 (O_607,N_49942,N_49502);
and UO_608 (O_608,N_49775,N_49797);
nor UO_609 (O_609,N_49742,N_49540);
and UO_610 (O_610,N_49872,N_49965);
and UO_611 (O_611,N_49592,N_49945);
and UO_612 (O_612,N_49830,N_49676);
and UO_613 (O_613,N_49651,N_49586);
or UO_614 (O_614,N_49529,N_49815);
or UO_615 (O_615,N_49644,N_49788);
nor UO_616 (O_616,N_49637,N_49762);
nand UO_617 (O_617,N_49994,N_49778);
nor UO_618 (O_618,N_49993,N_49739);
nand UO_619 (O_619,N_49524,N_49784);
or UO_620 (O_620,N_49709,N_49991);
or UO_621 (O_621,N_49866,N_49610);
or UO_622 (O_622,N_49990,N_49544);
and UO_623 (O_623,N_49936,N_49520);
or UO_624 (O_624,N_49996,N_49507);
and UO_625 (O_625,N_49765,N_49534);
or UO_626 (O_626,N_49797,N_49964);
nor UO_627 (O_627,N_49928,N_49555);
nor UO_628 (O_628,N_49934,N_49520);
nor UO_629 (O_629,N_49893,N_49607);
nor UO_630 (O_630,N_49878,N_49672);
or UO_631 (O_631,N_49980,N_49591);
or UO_632 (O_632,N_49895,N_49708);
nor UO_633 (O_633,N_49628,N_49692);
or UO_634 (O_634,N_49747,N_49500);
nand UO_635 (O_635,N_49836,N_49750);
nand UO_636 (O_636,N_49940,N_49920);
xnor UO_637 (O_637,N_49688,N_49508);
or UO_638 (O_638,N_49794,N_49536);
xor UO_639 (O_639,N_49525,N_49849);
nand UO_640 (O_640,N_49876,N_49723);
nand UO_641 (O_641,N_49605,N_49859);
nand UO_642 (O_642,N_49921,N_49934);
and UO_643 (O_643,N_49817,N_49738);
nor UO_644 (O_644,N_49643,N_49713);
xnor UO_645 (O_645,N_49537,N_49744);
nand UO_646 (O_646,N_49781,N_49789);
or UO_647 (O_647,N_49850,N_49768);
nor UO_648 (O_648,N_49617,N_49548);
and UO_649 (O_649,N_49523,N_49726);
or UO_650 (O_650,N_49545,N_49712);
nand UO_651 (O_651,N_49914,N_49590);
nor UO_652 (O_652,N_49773,N_49933);
nand UO_653 (O_653,N_49651,N_49735);
nand UO_654 (O_654,N_49731,N_49724);
xor UO_655 (O_655,N_49544,N_49719);
and UO_656 (O_656,N_49580,N_49889);
xor UO_657 (O_657,N_49788,N_49821);
or UO_658 (O_658,N_49803,N_49915);
or UO_659 (O_659,N_49999,N_49853);
xor UO_660 (O_660,N_49505,N_49792);
nand UO_661 (O_661,N_49731,N_49885);
xnor UO_662 (O_662,N_49877,N_49521);
xnor UO_663 (O_663,N_49655,N_49529);
or UO_664 (O_664,N_49588,N_49890);
nand UO_665 (O_665,N_49547,N_49715);
nor UO_666 (O_666,N_49636,N_49791);
and UO_667 (O_667,N_49945,N_49931);
nand UO_668 (O_668,N_49750,N_49570);
and UO_669 (O_669,N_49567,N_49765);
and UO_670 (O_670,N_49516,N_49694);
nor UO_671 (O_671,N_49697,N_49838);
xnor UO_672 (O_672,N_49877,N_49635);
nand UO_673 (O_673,N_49703,N_49894);
nor UO_674 (O_674,N_49842,N_49800);
nand UO_675 (O_675,N_49922,N_49649);
nand UO_676 (O_676,N_49756,N_49961);
or UO_677 (O_677,N_49884,N_49915);
and UO_678 (O_678,N_49922,N_49764);
nand UO_679 (O_679,N_49525,N_49698);
and UO_680 (O_680,N_49537,N_49675);
nor UO_681 (O_681,N_49928,N_49704);
nand UO_682 (O_682,N_49628,N_49637);
xnor UO_683 (O_683,N_49989,N_49582);
xor UO_684 (O_684,N_49837,N_49701);
and UO_685 (O_685,N_49984,N_49566);
nand UO_686 (O_686,N_49911,N_49908);
nor UO_687 (O_687,N_49731,N_49857);
or UO_688 (O_688,N_49556,N_49985);
and UO_689 (O_689,N_49528,N_49651);
nand UO_690 (O_690,N_49966,N_49689);
or UO_691 (O_691,N_49633,N_49630);
nand UO_692 (O_692,N_49774,N_49593);
nand UO_693 (O_693,N_49529,N_49962);
or UO_694 (O_694,N_49639,N_49896);
nor UO_695 (O_695,N_49657,N_49992);
or UO_696 (O_696,N_49790,N_49859);
nor UO_697 (O_697,N_49684,N_49717);
xnor UO_698 (O_698,N_49947,N_49904);
nand UO_699 (O_699,N_49816,N_49912);
and UO_700 (O_700,N_49694,N_49524);
or UO_701 (O_701,N_49686,N_49593);
xor UO_702 (O_702,N_49609,N_49741);
nand UO_703 (O_703,N_49874,N_49793);
or UO_704 (O_704,N_49537,N_49979);
and UO_705 (O_705,N_49895,N_49657);
xnor UO_706 (O_706,N_49981,N_49739);
or UO_707 (O_707,N_49801,N_49950);
nand UO_708 (O_708,N_49579,N_49736);
or UO_709 (O_709,N_49629,N_49748);
nor UO_710 (O_710,N_49920,N_49792);
nand UO_711 (O_711,N_49667,N_49851);
nor UO_712 (O_712,N_49705,N_49697);
nor UO_713 (O_713,N_49682,N_49724);
and UO_714 (O_714,N_49548,N_49914);
nor UO_715 (O_715,N_49921,N_49966);
and UO_716 (O_716,N_49865,N_49602);
and UO_717 (O_717,N_49788,N_49797);
and UO_718 (O_718,N_49770,N_49970);
nor UO_719 (O_719,N_49857,N_49920);
and UO_720 (O_720,N_49892,N_49842);
nor UO_721 (O_721,N_49906,N_49766);
xnor UO_722 (O_722,N_49759,N_49907);
nand UO_723 (O_723,N_49859,N_49939);
nor UO_724 (O_724,N_49761,N_49692);
nor UO_725 (O_725,N_49953,N_49893);
and UO_726 (O_726,N_49570,N_49715);
nor UO_727 (O_727,N_49862,N_49505);
or UO_728 (O_728,N_49548,N_49506);
xor UO_729 (O_729,N_49879,N_49756);
nand UO_730 (O_730,N_49946,N_49603);
xor UO_731 (O_731,N_49827,N_49568);
nand UO_732 (O_732,N_49616,N_49634);
and UO_733 (O_733,N_49803,N_49596);
nor UO_734 (O_734,N_49561,N_49776);
and UO_735 (O_735,N_49817,N_49990);
or UO_736 (O_736,N_49829,N_49902);
nor UO_737 (O_737,N_49579,N_49862);
nor UO_738 (O_738,N_49833,N_49712);
nand UO_739 (O_739,N_49949,N_49607);
nand UO_740 (O_740,N_49525,N_49798);
nand UO_741 (O_741,N_49657,N_49590);
xor UO_742 (O_742,N_49812,N_49821);
and UO_743 (O_743,N_49796,N_49759);
and UO_744 (O_744,N_49707,N_49673);
or UO_745 (O_745,N_49893,N_49982);
xor UO_746 (O_746,N_49912,N_49531);
or UO_747 (O_747,N_49987,N_49637);
nor UO_748 (O_748,N_49711,N_49826);
nand UO_749 (O_749,N_49826,N_49857);
nor UO_750 (O_750,N_49614,N_49697);
nand UO_751 (O_751,N_49740,N_49668);
xor UO_752 (O_752,N_49609,N_49509);
and UO_753 (O_753,N_49600,N_49548);
and UO_754 (O_754,N_49958,N_49857);
or UO_755 (O_755,N_49768,N_49946);
nand UO_756 (O_756,N_49766,N_49767);
or UO_757 (O_757,N_49608,N_49911);
or UO_758 (O_758,N_49715,N_49596);
and UO_759 (O_759,N_49654,N_49503);
nor UO_760 (O_760,N_49972,N_49787);
nor UO_761 (O_761,N_49507,N_49960);
or UO_762 (O_762,N_49988,N_49912);
nand UO_763 (O_763,N_49990,N_49512);
and UO_764 (O_764,N_49807,N_49631);
or UO_765 (O_765,N_49930,N_49650);
nor UO_766 (O_766,N_49930,N_49881);
and UO_767 (O_767,N_49683,N_49771);
and UO_768 (O_768,N_49852,N_49965);
or UO_769 (O_769,N_49549,N_49748);
or UO_770 (O_770,N_49688,N_49913);
and UO_771 (O_771,N_49836,N_49603);
and UO_772 (O_772,N_49580,N_49680);
and UO_773 (O_773,N_49628,N_49899);
nor UO_774 (O_774,N_49877,N_49712);
nand UO_775 (O_775,N_49659,N_49672);
nand UO_776 (O_776,N_49751,N_49514);
nand UO_777 (O_777,N_49719,N_49885);
or UO_778 (O_778,N_49518,N_49956);
or UO_779 (O_779,N_49537,N_49521);
or UO_780 (O_780,N_49892,N_49858);
xnor UO_781 (O_781,N_49930,N_49879);
nor UO_782 (O_782,N_49745,N_49803);
or UO_783 (O_783,N_49581,N_49684);
nand UO_784 (O_784,N_49825,N_49924);
nor UO_785 (O_785,N_49662,N_49781);
nor UO_786 (O_786,N_49989,N_49969);
nand UO_787 (O_787,N_49987,N_49527);
or UO_788 (O_788,N_49786,N_49915);
and UO_789 (O_789,N_49542,N_49768);
nor UO_790 (O_790,N_49840,N_49548);
or UO_791 (O_791,N_49522,N_49960);
xnor UO_792 (O_792,N_49614,N_49908);
or UO_793 (O_793,N_49563,N_49699);
nand UO_794 (O_794,N_49525,N_49925);
xor UO_795 (O_795,N_49523,N_49930);
nand UO_796 (O_796,N_49923,N_49823);
and UO_797 (O_797,N_49581,N_49759);
or UO_798 (O_798,N_49642,N_49799);
nand UO_799 (O_799,N_49675,N_49936);
nor UO_800 (O_800,N_49512,N_49964);
xor UO_801 (O_801,N_49967,N_49631);
nand UO_802 (O_802,N_49562,N_49591);
nor UO_803 (O_803,N_49517,N_49946);
nand UO_804 (O_804,N_49755,N_49736);
or UO_805 (O_805,N_49753,N_49561);
xnor UO_806 (O_806,N_49994,N_49644);
nor UO_807 (O_807,N_49573,N_49929);
and UO_808 (O_808,N_49750,N_49706);
and UO_809 (O_809,N_49980,N_49664);
and UO_810 (O_810,N_49602,N_49884);
and UO_811 (O_811,N_49895,N_49610);
or UO_812 (O_812,N_49740,N_49771);
and UO_813 (O_813,N_49743,N_49762);
nor UO_814 (O_814,N_49647,N_49741);
nand UO_815 (O_815,N_49862,N_49845);
nor UO_816 (O_816,N_49983,N_49978);
nor UO_817 (O_817,N_49806,N_49660);
nor UO_818 (O_818,N_49523,N_49978);
xor UO_819 (O_819,N_49579,N_49927);
and UO_820 (O_820,N_49640,N_49761);
nand UO_821 (O_821,N_49605,N_49510);
and UO_822 (O_822,N_49549,N_49645);
nand UO_823 (O_823,N_49802,N_49612);
nand UO_824 (O_824,N_49701,N_49822);
nor UO_825 (O_825,N_49710,N_49524);
and UO_826 (O_826,N_49664,N_49671);
nor UO_827 (O_827,N_49699,N_49839);
nand UO_828 (O_828,N_49920,N_49754);
or UO_829 (O_829,N_49517,N_49785);
and UO_830 (O_830,N_49971,N_49574);
nand UO_831 (O_831,N_49518,N_49973);
nor UO_832 (O_832,N_49625,N_49925);
nand UO_833 (O_833,N_49728,N_49519);
and UO_834 (O_834,N_49890,N_49990);
or UO_835 (O_835,N_49603,N_49771);
and UO_836 (O_836,N_49674,N_49856);
xnor UO_837 (O_837,N_49554,N_49514);
nand UO_838 (O_838,N_49775,N_49855);
nor UO_839 (O_839,N_49581,N_49608);
nor UO_840 (O_840,N_49750,N_49900);
and UO_841 (O_841,N_49680,N_49716);
nor UO_842 (O_842,N_49875,N_49914);
and UO_843 (O_843,N_49743,N_49869);
and UO_844 (O_844,N_49967,N_49843);
or UO_845 (O_845,N_49528,N_49753);
or UO_846 (O_846,N_49657,N_49614);
nor UO_847 (O_847,N_49508,N_49953);
nand UO_848 (O_848,N_49702,N_49917);
and UO_849 (O_849,N_49754,N_49819);
xor UO_850 (O_850,N_49566,N_49759);
or UO_851 (O_851,N_49517,N_49990);
nand UO_852 (O_852,N_49560,N_49556);
xnor UO_853 (O_853,N_49994,N_49895);
nand UO_854 (O_854,N_49857,N_49650);
nor UO_855 (O_855,N_49935,N_49614);
and UO_856 (O_856,N_49977,N_49739);
xnor UO_857 (O_857,N_49767,N_49828);
and UO_858 (O_858,N_49560,N_49686);
or UO_859 (O_859,N_49526,N_49619);
or UO_860 (O_860,N_49910,N_49754);
nand UO_861 (O_861,N_49668,N_49989);
nor UO_862 (O_862,N_49518,N_49785);
nor UO_863 (O_863,N_49541,N_49975);
and UO_864 (O_864,N_49643,N_49521);
nor UO_865 (O_865,N_49607,N_49694);
nand UO_866 (O_866,N_49843,N_49604);
or UO_867 (O_867,N_49894,N_49787);
nor UO_868 (O_868,N_49720,N_49775);
or UO_869 (O_869,N_49806,N_49713);
nand UO_870 (O_870,N_49700,N_49807);
and UO_871 (O_871,N_49544,N_49523);
or UO_872 (O_872,N_49512,N_49903);
and UO_873 (O_873,N_49861,N_49583);
or UO_874 (O_874,N_49752,N_49521);
or UO_875 (O_875,N_49771,N_49668);
nand UO_876 (O_876,N_49995,N_49764);
nand UO_877 (O_877,N_49591,N_49594);
or UO_878 (O_878,N_49521,N_49671);
nand UO_879 (O_879,N_49719,N_49682);
nor UO_880 (O_880,N_49939,N_49984);
nor UO_881 (O_881,N_49610,N_49875);
nand UO_882 (O_882,N_49974,N_49628);
xor UO_883 (O_883,N_49956,N_49887);
nor UO_884 (O_884,N_49865,N_49633);
nand UO_885 (O_885,N_49703,N_49607);
or UO_886 (O_886,N_49886,N_49960);
nor UO_887 (O_887,N_49729,N_49862);
or UO_888 (O_888,N_49749,N_49943);
nand UO_889 (O_889,N_49787,N_49893);
nand UO_890 (O_890,N_49784,N_49901);
and UO_891 (O_891,N_49637,N_49919);
xor UO_892 (O_892,N_49506,N_49538);
or UO_893 (O_893,N_49645,N_49698);
and UO_894 (O_894,N_49994,N_49983);
or UO_895 (O_895,N_49832,N_49850);
nor UO_896 (O_896,N_49570,N_49753);
nand UO_897 (O_897,N_49574,N_49895);
nand UO_898 (O_898,N_49803,N_49954);
or UO_899 (O_899,N_49910,N_49602);
nand UO_900 (O_900,N_49666,N_49594);
nand UO_901 (O_901,N_49642,N_49780);
and UO_902 (O_902,N_49838,N_49597);
and UO_903 (O_903,N_49898,N_49732);
nand UO_904 (O_904,N_49593,N_49941);
and UO_905 (O_905,N_49852,N_49500);
nor UO_906 (O_906,N_49633,N_49726);
nand UO_907 (O_907,N_49500,N_49851);
xor UO_908 (O_908,N_49627,N_49951);
nor UO_909 (O_909,N_49581,N_49821);
nor UO_910 (O_910,N_49831,N_49569);
nand UO_911 (O_911,N_49534,N_49842);
and UO_912 (O_912,N_49561,N_49572);
or UO_913 (O_913,N_49818,N_49800);
and UO_914 (O_914,N_49688,N_49639);
and UO_915 (O_915,N_49673,N_49716);
nand UO_916 (O_916,N_49800,N_49951);
or UO_917 (O_917,N_49990,N_49511);
or UO_918 (O_918,N_49569,N_49511);
and UO_919 (O_919,N_49671,N_49783);
nand UO_920 (O_920,N_49595,N_49503);
and UO_921 (O_921,N_49809,N_49786);
or UO_922 (O_922,N_49858,N_49651);
nor UO_923 (O_923,N_49781,N_49945);
or UO_924 (O_924,N_49801,N_49807);
nand UO_925 (O_925,N_49941,N_49509);
nor UO_926 (O_926,N_49822,N_49751);
nor UO_927 (O_927,N_49704,N_49650);
nor UO_928 (O_928,N_49546,N_49628);
and UO_929 (O_929,N_49552,N_49814);
nor UO_930 (O_930,N_49712,N_49636);
and UO_931 (O_931,N_49564,N_49655);
xnor UO_932 (O_932,N_49732,N_49686);
or UO_933 (O_933,N_49941,N_49530);
or UO_934 (O_934,N_49728,N_49745);
xor UO_935 (O_935,N_49757,N_49746);
nor UO_936 (O_936,N_49764,N_49972);
nand UO_937 (O_937,N_49658,N_49993);
and UO_938 (O_938,N_49917,N_49981);
nand UO_939 (O_939,N_49856,N_49943);
or UO_940 (O_940,N_49609,N_49923);
or UO_941 (O_941,N_49870,N_49907);
nor UO_942 (O_942,N_49813,N_49683);
or UO_943 (O_943,N_49772,N_49557);
and UO_944 (O_944,N_49507,N_49814);
or UO_945 (O_945,N_49872,N_49745);
nor UO_946 (O_946,N_49570,N_49695);
and UO_947 (O_947,N_49963,N_49520);
xor UO_948 (O_948,N_49779,N_49829);
nor UO_949 (O_949,N_49939,N_49641);
and UO_950 (O_950,N_49668,N_49978);
xnor UO_951 (O_951,N_49510,N_49548);
xnor UO_952 (O_952,N_49897,N_49704);
nor UO_953 (O_953,N_49874,N_49582);
and UO_954 (O_954,N_49847,N_49972);
or UO_955 (O_955,N_49658,N_49724);
xnor UO_956 (O_956,N_49916,N_49901);
and UO_957 (O_957,N_49797,N_49637);
and UO_958 (O_958,N_49911,N_49737);
xnor UO_959 (O_959,N_49529,N_49970);
or UO_960 (O_960,N_49888,N_49615);
and UO_961 (O_961,N_49913,N_49575);
xor UO_962 (O_962,N_49858,N_49685);
nand UO_963 (O_963,N_49799,N_49574);
nor UO_964 (O_964,N_49819,N_49880);
or UO_965 (O_965,N_49810,N_49623);
nor UO_966 (O_966,N_49877,N_49529);
nor UO_967 (O_967,N_49574,N_49996);
and UO_968 (O_968,N_49533,N_49593);
nor UO_969 (O_969,N_49661,N_49591);
and UO_970 (O_970,N_49727,N_49533);
nand UO_971 (O_971,N_49524,N_49666);
or UO_972 (O_972,N_49814,N_49960);
nor UO_973 (O_973,N_49691,N_49629);
nor UO_974 (O_974,N_49835,N_49585);
and UO_975 (O_975,N_49592,N_49735);
and UO_976 (O_976,N_49779,N_49672);
nor UO_977 (O_977,N_49518,N_49790);
nor UO_978 (O_978,N_49597,N_49686);
nand UO_979 (O_979,N_49834,N_49679);
nor UO_980 (O_980,N_49702,N_49994);
nor UO_981 (O_981,N_49831,N_49928);
and UO_982 (O_982,N_49857,N_49836);
nor UO_983 (O_983,N_49706,N_49871);
and UO_984 (O_984,N_49758,N_49896);
or UO_985 (O_985,N_49585,N_49915);
nor UO_986 (O_986,N_49595,N_49767);
or UO_987 (O_987,N_49740,N_49617);
and UO_988 (O_988,N_49647,N_49909);
xnor UO_989 (O_989,N_49712,N_49931);
and UO_990 (O_990,N_49673,N_49724);
or UO_991 (O_991,N_49592,N_49985);
and UO_992 (O_992,N_49787,N_49846);
xnor UO_993 (O_993,N_49514,N_49517);
and UO_994 (O_994,N_49688,N_49654);
or UO_995 (O_995,N_49962,N_49543);
or UO_996 (O_996,N_49723,N_49996);
and UO_997 (O_997,N_49977,N_49652);
nand UO_998 (O_998,N_49841,N_49859);
nor UO_999 (O_999,N_49703,N_49989);
and UO_1000 (O_1000,N_49819,N_49699);
or UO_1001 (O_1001,N_49835,N_49688);
nand UO_1002 (O_1002,N_49711,N_49515);
nand UO_1003 (O_1003,N_49836,N_49520);
or UO_1004 (O_1004,N_49590,N_49863);
nand UO_1005 (O_1005,N_49626,N_49657);
nand UO_1006 (O_1006,N_49568,N_49535);
nand UO_1007 (O_1007,N_49785,N_49721);
nor UO_1008 (O_1008,N_49638,N_49549);
or UO_1009 (O_1009,N_49945,N_49623);
nand UO_1010 (O_1010,N_49588,N_49994);
and UO_1011 (O_1011,N_49987,N_49569);
or UO_1012 (O_1012,N_49835,N_49549);
nor UO_1013 (O_1013,N_49704,N_49896);
nand UO_1014 (O_1014,N_49903,N_49738);
or UO_1015 (O_1015,N_49701,N_49880);
and UO_1016 (O_1016,N_49960,N_49948);
or UO_1017 (O_1017,N_49550,N_49721);
nor UO_1018 (O_1018,N_49523,N_49578);
xor UO_1019 (O_1019,N_49732,N_49986);
or UO_1020 (O_1020,N_49764,N_49864);
or UO_1021 (O_1021,N_49507,N_49694);
nand UO_1022 (O_1022,N_49814,N_49862);
nor UO_1023 (O_1023,N_49854,N_49979);
nand UO_1024 (O_1024,N_49781,N_49600);
nor UO_1025 (O_1025,N_49916,N_49913);
or UO_1026 (O_1026,N_49774,N_49949);
or UO_1027 (O_1027,N_49858,N_49976);
nor UO_1028 (O_1028,N_49639,N_49815);
nand UO_1029 (O_1029,N_49993,N_49793);
nor UO_1030 (O_1030,N_49754,N_49858);
or UO_1031 (O_1031,N_49839,N_49673);
nand UO_1032 (O_1032,N_49838,N_49689);
or UO_1033 (O_1033,N_49972,N_49935);
or UO_1034 (O_1034,N_49950,N_49558);
nand UO_1035 (O_1035,N_49843,N_49632);
nor UO_1036 (O_1036,N_49722,N_49872);
or UO_1037 (O_1037,N_49602,N_49674);
and UO_1038 (O_1038,N_49505,N_49582);
nand UO_1039 (O_1039,N_49685,N_49747);
nand UO_1040 (O_1040,N_49601,N_49571);
nor UO_1041 (O_1041,N_49606,N_49769);
or UO_1042 (O_1042,N_49765,N_49791);
nand UO_1043 (O_1043,N_49922,N_49565);
nand UO_1044 (O_1044,N_49767,N_49707);
or UO_1045 (O_1045,N_49777,N_49946);
nor UO_1046 (O_1046,N_49526,N_49736);
xnor UO_1047 (O_1047,N_49827,N_49879);
nand UO_1048 (O_1048,N_49662,N_49989);
and UO_1049 (O_1049,N_49772,N_49612);
nor UO_1050 (O_1050,N_49734,N_49597);
nand UO_1051 (O_1051,N_49735,N_49663);
or UO_1052 (O_1052,N_49636,N_49889);
nand UO_1053 (O_1053,N_49906,N_49544);
nor UO_1054 (O_1054,N_49765,N_49702);
or UO_1055 (O_1055,N_49725,N_49997);
and UO_1056 (O_1056,N_49651,N_49996);
and UO_1057 (O_1057,N_49989,N_49809);
and UO_1058 (O_1058,N_49895,N_49825);
and UO_1059 (O_1059,N_49714,N_49526);
or UO_1060 (O_1060,N_49968,N_49779);
nand UO_1061 (O_1061,N_49618,N_49663);
or UO_1062 (O_1062,N_49823,N_49794);
and UO_1063 (O_1063,N_49824,N_49920);
nor UO_1064 (O_1064,N_49880,N_49794);
or UO_1065 (O_1065,N_49930,N_49506);
or UO_1066 (O_1066,N_49799,N_49525);
nand UO_1067 (O_1067,N_49956,N_49536);
xnor UO_1068 (O_1068,N_49615,N_49519);
nor UO_1069 (O_1069,N_49636,N_49891);
xor UO_1070 (O_1070,N_49632,N_49662);
or UO_1071 (O_1071,N_49636,N_49562);
or UO_1072 (O_1072,N_49745,N_49639);
and UO_1073 (O_1073,N_49993,N_49629);
xor UO_1074 (O_1074,N_49760,N_49526);
and UO_1075 (O_1075,N_49721,N_49579);
and UO_1076 (O_1076,N_49881,N_49739);
and UO_1077 (O_1077,N_49886,N_49821);
nand UO_1078 (O_1078,N_49543,N_49801);
nand UO_1079 (O_1079,N_49651,N_49518);
and UO_1080 (O_1080,N_49519,N_49752);
nor UO_1081 (O_1081,N_49750,N_49798);
nor UO_1082 (O_1082,N_49583,N_49586);
or UO_1083 (O_1083,N_49719,N_49734);
and UO_1084 (O_1084,N_49837,N_49722);
or UO_1085 (O_1085,N_49979,N_49783);
or UO_1086 (O_1086,N_49661,N_49575);
xnor UO_1087 (O_1087,N_49503,N_49934);
and UO_1088 (O_1088,N_49765,N_49742);
or UO_1089 (O_1089,N_49732,N_49977);
or UO_1090 (O_1090,N_49911,N_49639);
xnor UO_1091 (O_1091,N_49594,N_49841);
nor UO_1092 (O_1092,N_49593,N_49860);
and UO_1093 (O_1093,N_49742,N_49906);
or UO_1094 (O_1094,N_49858,N_49666);
xnor UO_1095 (O_1095,N_49834,N_49723);
or UO_1096 (O_1096,N_49892,N_49625);
nand UO_1097 (O_1097,N_49919,N_49987);
nand UO_1098 (O_1098,N_49973,N_49986);
nor UO_1099 (O_1099,N_49663,N_49620);
or UO_1100 (O_1100,N_49545,N_49506);
or UO_1101 (O_1101,N_49808,N_49836);
and UO_1102 (O_1102,N_49639,N_49561);
xor UO_1103 (O_1103,N_49633,N_49563);
nor UO_1104 (O_1104,N_49713,N_49618);
nor UO_1105 (O_1105,N_49902,N_49630);
nand UO_1106 (O_1106,N_49618,N_49840);
nor UO_1107 (O_1107,N_49610,N_49697);
nor UO_1108 (O_1108,N_49991,N_49878);
nor UO_1109 (O_1109,N_49747,N_49817);
nor UO_1110 (O_1110,N_49985,N_49823);
xor UO_1111 (O_1111,N_49957,N_49833);
or UO_1112 (O_1112,N_49987,N_49790);
nor UO_1113 (O_1113,N_49615,N_49876);
or UO_1114 (O_1114,N_49886,N_49510);
nor UO_1115 (O_1115,N_49524,N_49901);
or UO_1116 (O_1116,N_49571,N_49777);
nand UO_1117 (O_1117,N_49509,N_49696);
and UO_1118 (O_1118,N_49661,N_49643);
and UO_1119 (O_1119,N_49677,N_49678);
xnor UO_1120 (O_1120,N_49609,N_49926);
and UO_1121 (O_1121,N_49662,N_49730);
and UO_1122 (O_1122,N_49730,N_49893);
and UO_1123 (O_1123,N_49686,N_49664);
nor UO_1124 (O_1124,N_49561,N_49565);
and UO_1125 (O_1125,N_49859,N_49895);
or UO_1126 (O_1126,N_49872,N_49632);
nand UO_1127 (O_1127,N_49600,N_49653);
nand UO_1128 (O_1128,N_49912,N_49716);
or UO_1129 (O_1129,N_49740,N_49545);
nand UO_1130 (O_1130,N_49740,N_49697);
nand UO_1131 (O_1131,N_49960,N_49800);
xor UO_1132 (O_1132,N_49976,N_49929);
nor UO_1133 (O_1133,N_49922,N_49852);
nor UO_1134 (O_1134,N_49870,N_49633);
or UO_1135 (O_1135,N_49532,N_49517);
or UO_1136 (O_1136,N_49697,N_49941);
or UO_1137 (O_1137,N_49719,N_49577);
nor UO_1138 (O_1138,N_49884,N_49516);
and UO_1139 (O_1139,N_49726,N_49591);
nor UO_1140 (O_1140,N_49684,N_49598);
nor UO_1141 (O_1141,N_49907,N_49523);
nand UO_1142 (O_1142,N_49965,N_49650);
or UO_1143 (O_1143,N_49673,N_49869);
nor UO_1144 (O_1144,N_49622,N_49821);
nor UO_1145 (O_1145,N_49564,N_49630);
or UO_1146 (O_1146,N_49746,N_49542);
and UO_1147 (O_1147,N_49591,N_49606);
or UO_1148 (O_1148,N_49836,N_49793);
or UO_1149 (O_1149,N_49697,N_49680);
and UO_1150 (O_1150,N_49745,N_49548);
nor UO_1151 (O_1151,N_49750,N_49661);
nand UO_1152 (O_1152,N_49739,N_49563);
and UO_1153 (O_1153,N_49818,N_49918);
nand UO_1154 (O_1154,N_49702,N_49686);
nor UO_1155 (O_1155,N_49791,N_49524);
or UO_1156 (O_1156,N_49756,N_49884);
nor UO_1157 (O_1157,N_49911,N_49957);
nand UO_1158 (O_1158,N_49901,N_49700);
nand UO_1159 (O_1159,N_49611,N_49568);
and UO_1160 (O_1160,N_49531,N_49608);
xnor UO_1161 (O_1161,N_49905,N_49657);
nand UO_1162 (O_1162,N_49880,N_49859);
and UO_1163 (O_1163,N_49507,N_49994);
nor UO_1164 (O_1164,N_49744,N_49887);
or UO_1165 (O_1165,N_49912,N_49785);
nand UO_1166 (O_1166,N_49627,N_49573);
nor UO_1167 (O_1167,N_49814,N_49619);
and UO_1168 (O_1168,N_49639,N_49602);
and UO_1169 (O_1169,N_49581,N_49711);
nor UO_1170 (O_1170,N_49623,N_49609);
nor UO_1171 (O_1171,N_49842,N_49934);
nor UO_1172 (O_1172,N_49613,N_49808);
xor UO_1173 (O_1173,N_49554,N_49628);
and UO_1174 (O_1174,N_49599,N_49590);
nor UO_1175 (O_1175,N_49870,N_49639);
and UO_1176 (O_1176,N_49626,N_49604);
nor UO_1177 (O_1177,N_49944,N_49743);
nor UO_1178 (O_1178,N_49949,N_49786);
and UO_1179 (O_1179,N_49556,N_49906);
nand UO_1180 (O_1180,N_49802,N_49759);
or UO_1181 (O_1181,N_49854,N_49807);
and UO_1182 (O_1182,N_49966,N_49564);
nor UO_1183 (O_1183,N_49907,N_49834);
nor UO_1184 (O_1184,N_49579,N_49617);
nor UO_1185 (O_1185,N_49814,N_49690);
nor UO_1186 (O_1186,N_49918,N_49709);
nor UO_1187 (O_1187,N_49732,N_49696);
nor UO_1188 (O_1188,N_49737,N_49550);
or UO_1189 (O_1189,N_49524,N_49763);
xor UO_1190 (O_1190,N_49943,N_49947);
or UO_1191 (O_1191,N_49996,N_49898);
nand UO_1192 (O_1192,N_49872,N_49559);
nor UO_1193 (O_1193,N_49648,N_49960);
nor UO_1194 (O_1194,N_49982,N_49797);
or UO_1195 (O_1195,N_49684,N_49955);
nor UO_1196 (O_1196,N_49762,N_49931);
or UO_1197 (O_1197,N_49810,N_49627);
xor UO_1198 (O_1198,N_49975,N_49907);
xnor UO_1199 (O_1199,N_49507,N_49706);
xor UO_1200 (O_1200,N_49819,N_49777);
and UO_1201 (O_1201,N_49772,N_49933);
nand UO_1202 (O_1202,N_49999,N_49743);
nor UO_1203 (O_1203,N_49714,N_49803);
nand UO_1204 (O_1204,N_49802,N_49580);
and UO_1205 (O_1205,N_49627,N_49843);
nand UO_1206 (O_1206,N_49646,N_49966);
nand UO_1207 (O_1207,N_49706,N_49822);
or UO_1208 (O_1208,N_49592,N_49941);
or UO_1209 (O_1209,N_49596,N_49695);
nor UO_1210 (O_1210,N_49551,N_49504);
nor UO_1211 (O_1211,N_49691,N_49941);
nand UO_1212 (O_1212,N_49516,N_49779);
or UO_1213 (O_1213,N_49922,N_49598);
and UO_1214 (O_1214,N_49982,N_49723);
and UO_1215 (O_1215,N_49605,N_49944);
and UO_1216 (O_1216,N_49801,N_49918);
or UO_1217 (O_1217,N_49526,N_49622);
and UO_1218 (O_1218,N_49801,N_49729);
and UO_1219 (O_1219,N_49601,N_49849);
xor UO_1220 (O_1220,N_49577,N_49879);
and UO_1221 (O_1221,N_49781,N_49625);
and UO_1222 (O_1222,N_49682,N_49922);
nor UO_1223 (O_1223,N_49539,N_49621);
or UO_1224 (O_1224,N_49600,N_49827);
nand UO_1225 (O_1225,N_49991,N_49582);
nor UO_1226 (O_1226,N_49969,N_49783);
nand UO_1227 (O_1227,N_49563,N_49670);
or UO_1228 (O_1228,N_49559,N_49873);
nor UO_1229 (O_1229,N_49538,N_49962);
and UO_1230 (O_1230,N_49545,N_49704);
or UO_1231 (O_1231,N_49683,N_49873);
and UO_1232 (O_1232,N_49720,N_49517);
or UO_1233 (O_1233,N_49952,N_49517);
nand UO_1234 (O_1234,N_49859,N_49532);
or UO_1235 (O_1235,N_49805,N_49523);
nand UO_1236 (O_1236,N_49679,N_49566);
and UO_1237 (O_1237,N_49810,N_49638);
xor UO_1238 (O_1238,N_49992,N_49683);
xor UO_1239 (O_1239,N_49695,N_49882);
nor UO_1240 (O_1240,N_49561,N_49545);
nor UO_1241 (O_1241,N_49946,N_49759);
nand UO_1242 (O_1242,N_49706,N_49767);
or UO_1243 (O_1243,N_49822,N_49560);
xnor UO_1244 (O_1244,N_49837,N_49686);
and UO_1245 (O_1245,N_49522,N_49605);
nand UO_1246 (O_1246,N_49727,N_49666);
and UO_1247 (O_1247,N_49874,N_49720);
nor UO_1248 (O_1248,N_49580,N_49946);
or UO_1249 (O_1249,N_49780,N_49733);
nor UO_1250 (O_1250,N_49612,N_49583);
or UO_1251 (O_1251,N_49831,N_49735);
and UO_1252 (O_1252,N_49572,N_49621);
and UO_1253 (O_1253,N_49856,N_49638);
nor UO_1254 (O_1254,N_49587,N_49709);
or UO_1255 (O_1255,N_49668,N_49645);
or UO_1256 (O_1256,N_49814,N_49518);
nor UO_1257 (O_1257,N_49952,N_49996);
or UO_1258 (O_1258,N_49893,N_49988);
nand UO_1259 (O_1259,N_49925,N_49720);
xnor UO_1260 (O_1260,N_49555,N_49643);
nand UO_1261 (O_1261,N_49821,N_49983);
and UO_1262 (O_1262,N_49685,N_49991);
and UO_1263 (O_1263,N_49761,N_49915);
or UO_1264 (O_1264,N_49738,N_49729);
or UO_1265 (O_1265,N_49509,N_49561);
and UO_1266 (O_1266,N_49674,N_49685);
nor UO_1267 (O_1267,N_49859,N_49873);
nand UO_1268 (O_1268,N_49692,N_49906);
nand UO_1269 (O_1269,N_49723,N_49513);
nor UO_1270 (O_1270,N_49653,N_49640);
or UO_1271 (O_1271,N_49904,N_49542);
and UO_1272 (O_1272,N_49504,N_49702);
or UO_1273 (O_1273,N_49564,N_49578);
nand UO_1274 (O_1274,N_49754,N_49900);
and UO_1275 (O_1275,N_49893,N_49589);
nand UO_1276 (O_1276,N_49799,N_49622);
nand UO_1277 (O_1277,N_49995,N_49877);
nand UO_1278 (O_1278,N_49530,N_49854);
nand UO_1279 (O_1279,N_49557,N_49603);
nand UO_1280 (O_1280,N_49988,N_49766);
nor UO_1281 (O_1281,N_49683,N_49796);
and UO_1282 (O_1282,N_49595,N_49886);
and UO_1283 (O_1283,N_49968,N_49628);
nor UO_1284 (O_1284,N_49797,N_49557);
and UO_1285 (O_1285,N_49768,N_49841);
and UO_1286 (O_1286,N_49700,N_49624);
xor UO_1287 (O_1287,N_49732,N_49652);
nand UO_1288 (O_1288,N_49630,N_49809);
and UO_1289 (O_1289,N_49895,N_49581);
nor UO_1290 (O_1290,N_49523,N_49906);
nand UO_1291 (O_1291,N_49693,N_49746);
and UO_1292 (O_1292,N_49668,N_49868);
nand UO_1293 (O_1293,N_49594,N_49508);
xnor UO_1294 (O_1294,N_49622,N_49646);
or UO_1295 (O_1295,N_49662,N_49925);
or UO_1296 (O_1296,N_49703,N_49609);
nand UO_1297 (O_1297,N_49936,N_49758);
nand UO_1298 (O_1298,N_49753,N_49738);
nor UO_1299 (O_1299,N_49652,N_49700);
or UO_1300 (O_1300,N_49780,N_49873);
or UO_1301 (O_1301,N_49930,N_49859);
xor UO_1302 (O_1302,N_49560,N_49926);
or UO_1303 (O_1303,N_49883,N_49639);
nand UO_1304 (O_1304,N_49688,N_49614);
nand UO_1305 (O_1305,N_49822,N_49892);
nor UO_1306 (O_1306,N_49942,N_49945);
or UO_1307 (O_1307,N_49629,N_49887);
and UO_1308 (O_1308,N_49684,N_49617);
or UO_1309 (O_1309,N_49565,N_49717);
and UO_1310 (O_1310,N_49548,N_49718);
nor UO_1311 (O_1311,N_49592,N_49673);
nor UO_1312 (O_1312,N_49888,N_49582);
nand UO_1313 (O_1313,N_49619,N_49748);
nand UO_1314 (O_1314,N_49955,N_49657);
or UO_1315 (O_1315,N_49755,N_49770);
and UO_1316 (O_1316,N_49982,N_49517);
nor UO_1317 (O_1317,N_49755,N_49813);
nor UO_1318 (O_1318,N_49571,N_49646);
or UO_1319 (O_1319,N_49572,N_49502);
nor UO_1320 (O_1320,N_49900,N_49719);
nor UO_1321 (O_1321,N_49864,N_49956);
and UO_1322 (O_1322,N_49810,N_49778);
nor UO_1323 (O_1323,N_49846,N_49569);
and UO_1324 (O_1324,N_49920,N_49634);
nor UO_1325 (O_1325,N_49701,N_49968);
or UO_1326 (O_1326,N_49756,N_49929);
and UO_1327 (O_1327,N_49541,N_49576);
nand UO_1328 (O_1328,N_49525,N_49804);
or UO_1329 (O_1329,N_49552,N_49603);
nor UO_1330 (O_1330,N_49779,N_49774);
xnor UO_1331 (O_1331,N_49850,N_49706);
nor UO_1332 (O_1332,N_49723,N_49701);
or UO_1333 (O_1333,N_49946,N_49694);
and UO_1334 (O_1334,N_49670,N_49534);
nand UO_1335 (O_1335,N_49761,N_49509);
and UO_1336 (O_1336,N_49761,N_49707);
xor UO_1337 (O_1337,N_49890,N_49953);
xor UO_1338 (O_1338,N_49685,N_49540);
and UO_1339 (O_1339,N_49627,N_49679);
and UO_1340 (O_1340,N_49809,N_49891);
nor UO_1341 (O_1341,N_49533,N_49641);
or UO_1342 (O_1342,N_49702,N_49603);
nand UO_1343 (O_1343,N_49647,N_49843);
nand UO_1344 (O_1344,N_49586,N_49986);
nor UO_1345 (O_1345,N_49926,N_49776);
or UO_1346 (O_1346,N_49799,N_49725);
nor UO_1347 (O_1347,N_49799,N_49587);
and UO_1348 (O_1348,N_49975,N_49882);
nor UO_1349 (O_1349,N_49595,N_49603);
and UO_1350 (O_1350,N_49519,N_49855);
and UO_1351 (O_1351,N_49842,N_49714);
or UO_1352 (O_1352,N_49557,N_49831);
nor UO_1353 (O_1353,N_49587,N_49522);
xnor UO_1354 (O_1354,N_49596,N_49921);
or UO_1355 (O_1355,N_49925,N_49501);
or UO_1356 (O_1356,N_49636,N_49624);
nor UO_1357 (O_1357,N_49532,N_49961);
xor UO_1358 (O_1358,N_49575,N_49593);
nand UO_1359 (O_1359,N_49561,N_49972);
nor UO_1360 (O_1360,N_49510,N_49737);
or UO_1361 (O_1361,N_49602,N_49591);
nand UO_1362 (O_1362,N_49668,N_49506);
nand UO_1363 (O_1363,N_49705,N_49661);
xor UO_1364 (O_1364,N_49606,N_49949);
nand UO_1365 (O_1365,N_49695,N_49865);
or UO_1366 (O_1366,N_49839,N_49730);
and UO_1367 (O_1367,N_49934,N_49897);
nor UO_1368 (O_1368,N_49631,N_49540);
nand UO_1369 (O_1369,N_49915,N_49735);
nand UO_1370 (O_1370,N_49900,N_49632);
nor UO_1371 (O_1371,N_49915,N_49796);
nor UO_1372 (O_1372,N_49847,N_49613);
nand UO_1373 (O_1373,N_49762,N_49997);
nor UO_1374 (O_1374,N_49956,N_49819);
nor UO_1375 (O_1375,N_49974,N_49917);
and UO_1376 (O_1376,N_49721,N_49875);
nand UO_1377 (O_1377,N_49833,N_49842);
or UO_1378 (O_1378,N_49523,N_49584);
nand UO_1379 (O_1379,N_49857,N_49917);
xnor UO_1380 (O_1380,N_49953,N_49616);
nor UO_1381 (O_1381,N_49609,N_49567);
nand UO_1382 (O_1382,N_49918,N_49582);
and UO_1383 (O_1383,N_49778,N_49634);
or UO_1384 (O_1384,N_49858,N_49705);
nor UO_1385 (O_1385,N_49594,N_49864);
nor UO_1386 (O_1386,N_49647,N_49806);
nor UO_1387 (O_1387,N_49948,N_49527);
nand UO_1388 (O_1388,N_49898,N_49838);
nand UO_1389 (O_1389,N_49520,N_49767);
nand UO_1390 (O_1390,N_49652,N_49829);
nor UO_1391 (O_1391,N_49713,N_49758);
and UO_1392 (O_1392,N_49503,N_49714);
nor UO_1393 (O_1393,N_49928,N_49732);
or UO_1394 (O_1394,N_49688,N_49963);
nand UO_1395 (O_1395,N_49572,N_49923);
nor UO_1396 (O_1396,N_49795,N_49536);
nor UO_1397 (O_1397,N_49909,N_49924);
nand UO_1398 (O_1398,N_49959,N_49957);
nor UO_1399 (O_1399,N_49630,N_49766);
nor UO_1400 (O_1400,N_49745,N_49902);
nand UO_1401 (O_1401,N_49625,N_49535);
nand UO_1402 (O_1402,N_49513,N_49874);
nand UO_1403 (O_1403,N_49939,N_49785);
nand UO_1404 (O_1404,N_49829,N_49738);
or UO_1405 (O_1405,N_49550,N_49781);
or UO_1406 (O_1406,N_49986,N_49623);
nor UO_1407 (O_1407,N_49591,N_49614);
or UO_1408 (O_1408,N_49924,N_49815);
xor UO_1409 (O_1409,N_49565,N_49695);
xnor UO_1410 (O_1410,N_49929,N_49935);
and UO_1411 (O_1411,N_49920,N_49873);
nand UO_1412 (O_1412,N_49802,N_49537);
or UO_1413 (O_1413,N_49793,N_49617);
nor UO_1414 (O_1414,N_49987,N_49754);
or UO_1415 (O_1415,N_49746,N_49947);
xor UO_1416 (O_1416,N_49844,N_49600);
nor UO_1417 (O_1417,N_49712,N_49756);
nor UO_1418 (O_1418,N_49918,N_49774);
and UO_1419 (O_1419,N_49615,N_49610);
and UO_1420 (O_1420,N_49559,N_49809);
nor UO_1421 (O_1421,N_49946,N_49722);
or UO_1422 (O_1422,N_49652,N_49571);
nor UO_1423 (O_1423,N_49845,N_49760);
nand UO_1424 (O_1424,N_49774,N_49920);
or UO_1425 (O_1425,N_49891,N_49978);
and UO_1426 (O_1426,N_49636,N_49841);
and UO_1427 (O_1427,N_49501,N_49553);
nand UO_1428 (O_1428,N_49744,N_49817);
nand UO_1429 (O_1429,N_49575,N_49711);
nor UO_1430 (O_1430,N_49598,N_49506);
xor UO_1431 (O_1431,N_49931,N_49589);
xnor UO_1432 (O_1432,N_49786,N_49726);
nor UO_1433 (O_1433,N_49781,N_49964);
nand UO_1434 (O_1434,N_49680,N_49631);
or UO_1435 (O_1435,N_49719,N_49809);
or UO_1436 (O_1436,N_49641,N_49756);
nor UO_1437 (O_1437,N_49539,N_49809);
nor UO_1438 (O_1438,N_49735,N_49552);
and UO_1439 (O_1439,N_49527,N_49788);
nor UO_1440 (O_1440,N_49875,N_49606);
and UO_1441 (O_1441,N_49910,N_49876);
nand UO_1442 (O_1442,N_49954,N_49714);
nand UO_1443 (O_1443,N_49805,N_49646);
or UO_1444 (O_1444,N_49833,N_49513);
nand UO_1445 (O_1445,N_49756,N_49970);
or UO_1446 (O_1446,N_49507,N_49632);
and UO_1447 (O_1447,N_49859,N_49845);
nand UO_1448 (O_1448,N_49683,N_49680);
or UO_1449 (O_1449,N_49554,N_49734);
nor UO_1450 (O_1450,N_49989,N_49776);
nor UO_1451 (O_1451,N_49536,N_49593);
and UO_1452 (O_1452,N_49834,N_49831);
nand UO_1453 (O_1453,N_49665,N_49954);
nand UO_1454 (O_1454,N_49502,N_49922);
or UO_1455 (O_1455,N_49618,N_49800);
xnor UO_1456 (O_1456,N_49582,N_49983);
or UO_1457 (O_1457,N_49599,N_49884);
nand UO_1458 (O_1458,N_49746,N_49713);
or UO_1459 (O_1459,N_49994,N_49782);
nand UO_1460 (O_1460,N_49588,N_49560);
nand UO_1461 (O_1461,N_49637,N_49641);
or UO_1462 (O_1462,N_49519,N_49845);
nand UO_1463 (O_1463,N_49597,N_49522);
and UO_1464 (O_1464,N_49738,N_49735);
xor UO_1465 (O_1465,N_49651,N_49725);
and UO_1466 (O_1466,N_49715,N_49552);
nand UO_1467 (O_1467,N_49506,N_49585);
nand UO_1468 (O_1468,N_49964,N_49670);
or UO_1469 (O_1469,N_49959,N_49964);
nand UO_1470 (O_1470,N_49832,N_49879);
and UO_1471 (O_1471,N_49934,N_49862);
xnor UO_1472 (O_1472,N_49777,N_49967);
or UO_1473 (O_1473,N_49593,N_49736);
and UO_1474 (O_1474,N_49638,N_49802);
nand UO_1475 (O_1475,N_49977,N_49704);
nor UO_1476 (O_1476,N_49726,N_49858);
nand UO_1477 (O_1477,N_49907,N_49680);
xnor UO_1478 (O_1478,N_49685,N_49638);
and UO_1479 (O_1479,N_49783,N_49773);
nor UO_1480 (O_1480,N_49560,N_49604);
or UO_1481 (O_1481,N_49632,N_49822);
nor UO_1482 (O_1482,N_49519,N_49644);
nor UO_1483 (O_1483,N_49906,N_49515);
nor UO_1484 (O_1484,N_49816,N_49518);
and UO_1485 (O_1485,N_49634,N_49558);
nand UO_1486 (O_1486,N_49665,N_49739);
and UO_1487 (O_1487,N_49825,N_49683);
xnor UO_1488 (O_1488,N_49851,N_49932);
or UO_1489 (O_1489,N_49771,N_49595);
nand UO_1490 (O_1490,N_49988,N_49510);
nand UO_1491 (O_1491,N_49746,N_49573);
xor UO_1492 (O_1492,N_49593,N_49664);
nand UO_1493 (O_1493,N_49661,N_49793);
and UO_1494 (O_1494,N_49700,N_49562);
and UO_1495 (O_1495,N_49774,N_49562);
or UO_1496 (O_1496,N_49896,N_49805);
or UO_1497 (O_1497,N_49930,N_49557);
nor UO_1498 (O_1498,N_49905,N_49561);
nor UO_1499 (O_1499,N_49941,N_49773);
nor UO_1500 (O_1500,N_49629,N_49974);
and UO_1501 (O_1501,N_49862,N_49596);
nand UO_1502 (O_1502,N_49701,N_49673);
xor UO_1503 (O_1503,N_49781,N_49556);
or UO_1504 (O_1504,N_49892,N_49672);
xnor UO_1505 (O_1505,N_49850,N_49849);
or UO_1506 (O_1506,N_49755,N_49932);
nand UO_1507 (O_1507,N_49574,N_49995);
and UO_1508 (O_1508,N_49546,N_49722);
nor UO_1509 (O_1509,N_49997,N_49509);
nand UO_1510 (O_1510,N_49760,N_49901);
nor UO_1511 (O_1511,N_49851,N_49745);
or UO_1512 (O_1512,N_49954,N_49741);
nor UO_1513 (O_1513,N_49874,N_49676);
nor UO_1514 (O_1514,N_49710,N_49619);
nor UO_1515 (O_1515,N_49646,N_49997);
or UO_1516 (O_1516,N_49636,N_49667);
nor UO_1517 (O_1517,N_49667,N_49501);
nor UO_1518 (O_1518,N_49972,N_49925);
or UO_1519 (O_1519,N_49777,N_49992);
nor UO_1520 (O_1520,N_49619,N_49817);
nor UO_1521 (O_1521,N_49535,N_49605);
or UO_1522 (O_1522,N_49705,N_49581);
nand UO_1523 (O_1523,N_49771,N_49612);
or UO_1524 (O_1524,N_49768,N_49707);
nor UO_1525 (O_1525,N_49752,N_49804);
nand UO_1526 (O_1526,N_49539,N_49797);
and UO_1527 (O_1527,N_49972,N_49980);
and UO_1528 (O_1528,N_49856,N_49835);
nand UO_1529 (O_1529,N_49956,N_49869);
or UO_1530 (O_1530,N_49729,N_49958);
and UO_1531 (O_1531,N_49827,N_49634);
xnor UO_1532 (O_1532,N_49517,N_49950);
nor UO_1533 (O_1533,N_49908,N_49859);
or UO_1534 (O_1534,N_49502,N_49734);
or UO_1535 (O_1535,N_49734,N_49891);
and UO_1536 (O_1536,N_49720,N_49937);
nor UO_1537 (O_1537,N_49619,N_49818);
or UO_1538 (O_1538,N_49971,N_49683);
xor UO_1539 (O_1539,N_49961,N_49933);
nand UO_1540 (O_1540,N_49963,N_49919);
nand UO_1541 (O_1541,N_49741,N_49594);
or UO_1542 (O_1542,N_49555,N_49827);
and UO_1543 (O_1543,N_49895,N_49664);
nand UO_1544 (O_1544,N_49773,N_49866);
and UO_1545 (O_1545,N_49999,N_49898);
xnor UO_1546 (O_1546,N_49513,N_49588);
and UO_1547 (O_1547,N_49605,N_49685);
nand UO_1548 (O_1548,N_49970,N_49710);
xnor UO_1549 (O_1549,N_49822,N_49966);
or UO_1550 (O_1550,N_49901,N_49515);
nand UO_1551 (O_1551,N_49872,N_49925);
nand UO_1552 (O_1552,N_49948,N_49560);
and UO_1553 (O_1553,N_49993,N_49603);
and UO_1554 (O_1554,N_49520,N_49809);
and UO_1555 (O_1555,N_49835,N_49831);
nand UO_1556 (O_1556,N_49669,N_49616);
and UO_1557 (O_1557,N_49575,N_49955);
and UO_1558 (O_1558,N_49576,N_49739);
nand UO_1559 (O_1559,N_49877,N_49746);
or UO_1560 (O_1560,N_49638,N_49897);
nand UO_1561 (O_1561,N_49572,N_49859);
or UO_1562 (O_1562,N_49609,N_49986);
nor UO_1563 (O_1563,N_49635,N_49954);
or UO_1564 (O_1564,N_49939,N_49935);
xnor UO_1565 (O_1565,N_49970,N_49973);
and UO_1566 (O_1566,N_49632,N_49592);
or UO_1567 (O_1567,N_49737,N_49697);
nor UO_1568 (O_1568,N_49989,N_49756);
or UO_1569 (O_1569,N_49832,N_49501);
nand UO_1570 (O_1570,N_49698,N_49975);
nand UO_1571 (O_1571,N_49637,N_49750);
and UO_1572 (O_1572,N_49844,N_49964);
or UO_1573 (O_1573,N_49605,N_49608);
and UO_1574 (O_1574,N_49509,N_49575);
or UO_1575 (O_1575,N_49819,N_49788);
xor UO_1576 (O_1576,N_49526,N_49872);
or UO_1577 (O_1577,N_49553,N_49717);
nand UO_1578 (O_1578,N_49990,N_49828);
nand UO_1579 (O_1579,N_49685,N_49892);
nor UO_1580 (O_1580,N_49521,N_49959);
nor UO_1581 (O_1581,N_49970,N_49584);
and UO_1582 (O_1582,N_49912,N_49978);
and UO_1583 (O_1583,N_49996,N_49600);
nor UO_1584 (O_1584,N_49878,N_49747);
or UO_1585 (O_1585,N_49954,N_49692);
xnor UO_1586 (O_1586,N_49627,N_49631);
and UO_1587 (O_1587,N_49769,N_49947);
xor UO_1588 (O_1588,N_49624,N_49949);
nand UO_1589 (O_1589,N_49643,N_49723);
or UO_1590 (O_1590,N_49911,N_49864);
or UO_1591 (O_1591,N_49789,N_49699);
nand UO_1592 (O_1592,N_49752,N_49807);
nor UO_1593 (O_1593,N_49972,N_49968);
xnor UO_1594 (O_1594,N_49642,N_49563);
nor UO_1595 (O_1595,N_49938,N_49511);
and UO_1596 (O_1596,N_49763,N_49731);
and UO_1597 (O_1597,N_49598,N_49901);
xnor UO_1598 (O_1598,N_49727,N_49991);
nand UO_1599 (O_1599,N_49565,N_49968);
nand UO_1600 (O_1600,N_49849,N_49702);
nor UO_1601 (O_1601,N_49550,N_49718);
nor UO_1602 (O_1602,N_49562,N_49537);
nor UO_1603 (O_1603,N_49987,N_49903);
and UO_1604 (O_1604,N_49979,N_49645);
nor UO_1605 (O_1605,N_49596,N_49898);
or UO_1606 (O_1606,N_49642,N_49721);
nand UO_1607 (O_1607,N_49594,N_49710);
nor UO_1608 (O_1608,N_49989,N_49632);
nand UO_1609 (O_1609,N_49737,N_49883);
nor UO_1610 (O_1610,N_49892,N_49829);
nor UO_1611 (O_1611,N_49990,N_49751);
nor UO_1612 (O_1612,N_49900,N_49588);
xnor UO_1613 (O_1613,N_49593,N_49968);
and UO_1614 (O_1614,N_49916,N_49942);
nor UO_1615 (O_1615,N_49898,N_49727);
nor UO_1616 (O_1616,N_49910,N_49957);
and UO_1617 (O_1617,N_49504,N_49695);
xnor UO_1618 (O_1618,N_49902,N_49760);
nor UO_1619 (O_1619,N_49580,N_49543);
nand UO_1620 (O_1620,N_49804,N_49785);
nand UO_1621 (O_1621,N_49833,N_49802);
and UO_1622 (O_1622,N_49751,N_49967);
nor UO_1623 (O_1623,N_49517,N_49576);
and UO_1624 (O_1624,N_49936,N_49745);
nand UO_1625 (O_1625,N_49673,N_49750);
nand UO_1626 (O_1626,N_49844,N_49547);
nand UO_1627 (O_1627,N_49920,N_49709);
and UO_1628 (O_1628,N_49635,N_49864);
nor UO_1629 (O_1629,N_49693,N_49758);
xor UO_1630 (O_1630,N_49668,N_49821);
nor UO_1631 (O_1631,N_49534,N_49565);
nor UO_1632 (O_1632,N_49876,N_49885);
nor UO_1633 (O_1633,N_49974,N_49811);
nand UO_1634 (O_1634,N_49656,N_49958);
nand UO_1635 (O_1635,N_49723,N_49503);
nor UO_1636 (O_1636,N_49720,N_49651);
nand UO_1637 (O_1637,N_49537,N_49661);
nor UO_1638 (O_1638,N_49812,N_49872);
or UO_1639 (O_1639,N_49553,N_49791);
or UO_1640 (O_1640,N_49755,N_49587);
or UO_1641 (O_1641,N_49637,N_49677);
nand UO_1642 (O_1642,N_49586,N_49900);
and UO_1643 (O_1643,N_49697,N_49681);
nor UO_1644 (O_1644,N_49894,N_49899);
nor UO_1645 (O_1645,N_49864,N_49768);
nand UO_1646 (O_1646,N_49569,N_49666);
xor UO_1647 (O_1647,N_49639,N_49997);
nand UO_1648 (O_1648,N_49899,N_49922);
or UO_1649 (O_1649,N_49990,N_49618);
nor UO_1650 (O_1650,N_49573,N_49517);
nand UO_1651 (O_1651,N_49636,N_49581);
and UO_1652 (O_1652,N_49515,N_49514);
or UO_1653 (O_1653,N_49895,N_49750);
nor UO_1654 (O_1654,N_49653,N_49605);
and UO_1655 (O_1655,N_49626,N_49654);
and UO_1656 (O_1656,N_49978,N_49799);
nand UO_1657 (O_1657,N_49681,N_49881);
nand UO_1658 (O_1658,N_49951,N_49881);
and UO_1659 (O_1659,N_49615,N_49853);
xnor UO_1660 (O_1660,N_49642,N_49754);
and UO_1661 (O_1661,N_49553,N_49528);
and UO_1662 (O_1662,N_49889,N_49865);
and UO_1663 (O_1663,N_49677,N_49718);
nand UO_1664 (O_1664,N_49748,N_49752);
nor UO_1665 (O_1665,N_49642,N_49553);
and UO_1666 (O_1666,N_49812,N_49602);
nor UO_1667 (O_1667,N_49790,N_49702);
nor UO_1668 (O_1668,N_49846,N_49908);
nand UO_1669 (O_1669,N_49913,N_49720);
or UO_1670 (O_1670,N_49710,N_49783);
nand UO_1671 (O_1671,N_49882,N_49766);
nor UO_1672 (O_1672,N_49988,N_49610);
nand UO_1673 (O_1673,N_49703,N_49694);
or UO_1674 (O_1674,N_49579,N_49722);
nor UO_1675 (O_1675,N_49840,N_49653);
and UO_1676 (O_1676,N_49956,N_49985);
xnor UO_1677 (O_1677,N_49791,N_49550);
nand UO_1678 (O_1678,N_49749,N_49630);
xnor UO_1679 (O_1679,N_49883,N_49712);
nor UO_1680 (O_1680,N_49709,N_49571);
nand UO_1681 (O_1681,N_49729,N_49629);
and UO_1682 (O_1682,N_49898,N_49782);
xor UO_1683 (O_1683,N_49808,N_49868);
or UO_1684 (O_1684,N_49662,N_49523);
nor UO_1685 (O_1685,N_49669,N_49958);
xor UO_1686 (O_1686,N_49655,N_49865);
and UO_1687 (O_1687,N_49584,N_49784);
or UO_1688 (O_1688,N_49676,N_49832);
nand UO_1689 (O_1689,N_49655,N_49656);
nor UO_1690 (O_1690,N_49502,N_49888);
nor UO_1691 (O_1691,N_49885,N_49545);
nand UO_1692 (O_1692,N_49922,N_49772);
or UO_1693 (O_1693,N_49888,N_49864);
nand UO_1694 (O_1694,N_49908,N_49627);
or UO_1695 (O_1695,N_49926,N_49851);
and UO_1696 (O_1696,N_49990,N_49662);
or UO_1697 (O_1697,N_49870,N_49786);
nor UO_1698 (O_1698,N_49581,N_49996);
or UO_1699 (O_1699,N_49841,N_49998);
and UO_1700 (O_1700,N_49777,N_49956);
nand UO_1701 (O_1701,N_49963,N_49948);
and UO_1702 (O_1702,N_49621,N_49823);
nand UO_1703 (O_1703,N_49747,N_49965);
or UO_1704 (O_1704,N_49798,N_49643);
or UO_1705 (O_1705,N_49873,N_49964);
or UO_1706 (O_1706,N_49810,N_49858);
nor UO_1707 (O_1707,N_49834,N_49880);
and UO_1708 (O_1708,N_49528,N_49861);
and UO_1709 (O_1709,N_49652,N_49889);
and UO_1710 (O_1710,N_49918,N_49912);
and UO_1711 (O_1711,N_49588,N_49790);
nor UO_1712 (O_1712,N_49993,N_49998);
xnor UO_1713 (O_1713,N_49659,N_49546);
nand UO_1714 (O_1714,N_49565,N_49671);
xnor UO_1715 (O_1715,N_49768,N_49620);
and UO_1716 (O_1716,N_49777,N_49548);
nor UO_1717 (O_1717,N_49703,N_49598);
or UO_1718 (O_1718,N_49869,N_49824);
nand UO_1719 (O_1719,N_49976,N_49877);
and UO_1720 (O_1720,N_49585,N_49845);
or UO_1721 (O_1721,N_49577,N_49864);
nor UO_1722 (O_1722,N_49908,N_49895);
and UO_1723 (O_1723,N_49654,N_49577);
or UO_1724 (O_1724,N_49880,N_49800);
and UO_1725 (O_1725,N_49772,N_49646);
or UO_1726 (O_1726,N_49567,N_49691);
and UO_1727 (O_1727,N_49812,N_49794);
nand UO_1728 (O_1728,N_49723,N_49544);
nand UO_1729 (O_1729,N_49644,N_49594);
xnor UO_1730 (O_1730,N_49959,N_49713);
nor UO_1731 (O_1731,N_49752,N_49772);
nor UO_1732 (O_1732,N_49827,N_49929);
and UO_1733 (O_1733,N_49624,N_49612);
nor UO_1734 (O_1734,N_49714,N_49505);
nand UO_1735 (O_1735,N_49523,N_49863);
and UO_1736 (O_1736,N_49728,N_49618);
or UO_1737 (O_1737,N_49798,N_49511);
and UO_1738 (O_1738,N_49504,N_49553);
or UO_1739 (O_1739,N_49800,N_49994);
or UO_1740 (O_1740,N_49880,N_49664);
or UO_1741 (O_1741,N_49905,N_49892);
nand UO_1742 (O_1742,N_49824,N_49795);
or UO_1743 (O_1743,N_49927,N_49583);
xnor UO_1744 (O_1744,N_49786,N_49659);
and UO_1745 (O_1745,N_49576,N_49761);
nor UO_1746 (O_1746,N_49997,N_49603);
xor UO_1747 (O_1747,N_49830,N_49843);
or UO_1748 (O_1748,N_49545,N_49546);
nor UO_1749 (O_1749,N_49826,N_49753);
or UO_1750 (O_1750,N_49640,N_49568);
or UO_1751 (O_1751,N_49775,N_49936);
and UO_1752 (O_1752,N_49768,N_49528);
nor UO_1753 (O_1753,N_49713,N_49593);
nand UO_1754 (O_1754,N_49758,N_49502);
or UO_1755 (O_1755,N_49579,N_49952);
or UO_1756 (O_1756,N_49905,N_49779);
and UO_1757 (O_1757,N_49949,N_49583);
and UO_1758 (O_1758,N_49967,N_49635);
nand UO_1759 (O_1759,N_49811,N_49694);
xor UO_1760 (O_1760,N_49584,N_49845);
nand UO_1761 (O_1761,N_49846,N_49880);
and UO_1762 (O_1762,N_49737,N_49771);
nor UO_1763 (O_1763,N_49561,N_49892);
xor UO_1764 (O_1764,N_49511,N_49527);
and UO_1765 (O_1765,N_49802,N_49505);
nand UO_1766 (O_1766,N_49881,N_49805);
nor UO_1767 (O_1767,N_49511,N_49550);
nor UO_1768 (O_1768,N_49563,N_49585);
and UO_1769 (O_1769,N_49827,N_49638);
or UO_1770 (O_1770,N_49829,N_49880);
nor UO_1771 (O_1771,N_49557,N_49933);
or UO_1772 (O_1772,N_49658,N_49956);
or UO_1773 (O_1773,N_49826,N_49971);
nand UO_1774 (O_1774,N_49845,N_49659);
and UO_1775 (O_1775,N_49685,N_49705);
xor UO_1776 (O_1776,N_49592,N_49708);
or UO_1777 (O_1777,N_49866,N_49778);
or UO_1778 (O_1778,N_49788,N_49738);
and UO_1779 (O_1779,N_49558,N_49785);
and UO_1780 (O_1780,N_49545,N_49855);
nor UO_1781 (O_1781,N_49624,N_49653);
nor UO_1782 (O_1782,N_49920,N_49731);
and UO_1783 (O_1783,N_49630,N_49836);
nand UO_1784 (O_1784,N_49579,N_49662);
and UO_1785 (O_1785,N_49875,N_49831);
nand UO_1786 (O_1786,N_49514,N_49693);
or UO_1787 (O_1787,N_49799,N_49790);
and UO_1788 (O_1788,N_49899,N_49956);
or UO_1789 (O_1789,N_49963,N_49956);
or UO_1790 (O_1790,N_49843,N_49515);
nor UO_1791 (O_1791,N_49717,N_49587);
nor UO_1792 (O_1792,N_49567,N_49814);
and UO_1793 (O_1793,N_49992,N_49765);
nand UO_1794 (O_1794,N_49601,N_49773);
nand UO_1795 (O_1795,N_49783,N_49873);
nor UO_1796 (O_1796,N_49693,N_49554);
and UO_1797 (O_1797,N_49943,N_49597);
and UO_1798 (O_1798,N_49705,N_49837);
nand UO_1799 (O_1799,N_49525,N_49590);
nand UO_1800 (O_1800,N_49811,N_49576);
nor UO_1801 (O_1801,N_49951,N_49661);
xor UO_1802 (O_1802,N_49670,N_49555);
or UO_1803 (O_1803,N_49871,N_49941);
and UO_1804 (O_1804,N_49599,N_49694);
and UO_1805 (O_1805,N_49743,N_49861);
nand UO_1806 (O_1806,N_49563,N_49531);
or UO_1807 (O_1807,N_49919,N_49901);
and UO_1808 (O_1808,N_49661,N_49523);
xor UO_1809 (O_1809,N_49896,N_49916);
nand UO_1810 (O_1810,N_49947,N_49808);
nand UO_1811 (O_1811,N_49714,N_49884);
nor UO_1812 (O_1812,N_49554,N_49667);
nand UO_1813 (O_1813,N_49510,N_49588);
nor UO_1814 (O_1814,N_49660,N_49889);
xnor UO_1815 (O_1815,N_49615,N_49779);
xor UO_1816 (O_1816,N_49857,N_49874);
nand UO_1817 (O_1817,N_49823,N_49802);
nand UO_1818 (O_1818,N_49507,N_49697);
and UO_1819 (O_1819,N_49540,N_49504);
nor UO_1820 (O_1820,N_49689,N_49712);
nand UO_1821 (O_1821,N_49585,N_49709);
xor UO_1822 (O_1822,N_49529,N_49744);
nor UO_1823 (O_1823,N_49979,N_49787);
nand UO_1824 (O_1824,N_49857,N_49711);
and UO_1825 (O_1825,N_49967,N_49904);
and UO_1826 (O_1826,N_49780,N_49603);
or UO_1827 (O_1827,N_49697,N_49587);
and UO_1828 (O_1828,N_49902,N_49716);
xnor UO_1829 (O_1829,N_49866,N_49691);
nor UO_1830 (O_1830,N_49963,N_49842);
and UO_1831 (O_1831,N_49953,N_49744);
nand UO_1832 (O_1832,N_49564,N_49940);
nor UO_1833 (O_1833,N_49513,N_49739);
or UO_1834 (O_1834,N_49780,N_49810);
nand UO_1835 (O_1835,N_49845,N_49640);
and UO_1836 (O_1836,N_49711,N_49712);
nor UO_1837 (O_1837,N_49708,N_49808);
nor UO_1838 (O_1838,N_49881,N_49566);
or UO_1839 (O_1839,N_49649,N_49576);
nand UO_1840 (O_1840,N_49904,N_49991);
nor UO_1841 (O_1841,N_49581,N_49503);
and UO_1842 (O_1842,N_49604,N_49887);
nand UO_1843 (O_1843,N_49974,N_49576);
or UO_1844 (O_1844,N_49543,N_49872);
or UO_1845 (O_1845,N_49876,N_49589);
or UO_1846 (O_1846,N_49909,N_49517);
nand UO_1847 (O_1847,N_49571,N_49694);
xnor UO_1848 (O_1848,N_49823,N_49575);
nor UO_1849 (O_1849,N_49773,N_49915);
and UO_1850 (O_1850,N_49928,N_49899);
and UO_1851 (O_1851,N_49693,N_49725);
xor UO_1852 (O_1852,N_49506,N_49993);
nor UO_1853 (O_1853,N_49993,N_49754);
or UO_1854 (O_1854,N_49735,N_49792);
nor UO_1855 (O_1855,N_49546,N_49528);
or UO_1856 (O_1856,N_49849,N_49512);
and UO_1857 (O_1857,N_49891,N_49910);
nor UO_1858 (O_1858,N_49678,N_49703);
nand UO_1859 (O_1859,N_49624,N_49855);
xnor UO_1860 (O_1860,N_49896,N_49884);
nand UO_1861 (O_1861,N_49672,N_49835);
nor UO_1862 (O_1862,N_49897,N_49693);
xor UO_1863 (O_1863,N_49654,N_49598);
and UO_1864 (O_1864,N_49868,N_49709);
nand UO_1865 (O_1865,N_49571,N_49977);
nor UO_1866 (O_1866,N_49771,N_49999);
nor UO_1867 (O_1867,N_49684,N_49797);
nor UO_1868 (O_1868,N_49788,N_49920);
and UO_1869 (O_1869,N_49522,N_49695);
nand UO_1870 (O_1870,N_49916,N_49768);
and UO_1871 (O_1871,N_49884,N_49844);
nand UO_1872 (O_1872,N_49626,N_49974);
and UO_1873 (O_1873,N_49803,N_49567);
nand UO_1874 (O_1874,N_49501,N_49906);
and UO_1875 (O_1875,N_49624,N_49760);
or UO_1876 (O_1876,N_49708,N_49876);
or UO_1877 (O_1877,N_49930,N_49798);
nand UO_1878 (O_1878,N_49891,N_49698);
and UO_1879 (O_1879,N_49508,N_49909);
nand UO_1880 (O_1880,N_49774,N_49882);
nand UO_1881 (O_1881,N_49915,N_49808);
nor UO_1882 (O_1882,N_49604,N_49620);
or UO_1883 (O_1883,N_49919,N_49611);
and UO_1884 (O_1884,N_49679,N_49780);
and UO_1885 (O_1885,N_49560,N_49550);
nand UO_1886 (O_1886,N_49961,N_49734);
nor UO_1887 (O_1887,N_49857,N_49805);
nand UO_1888 (O_1888,N_49715,N_49676);
nor UO_1889 (O_1889,N_49808,N_49568);
nand UO_1890 (O_1890,N_49944,N_49690);
or UO_1891 (O_1891,N_49627,N_49899);
and UO_1892 (O_1892,N_49776,N_49809);
xor UO_1893 (O_1893,N_49567,N_49707);
and UO_1894 (O_1894,N_49501,N_49577);
nand UO_1895 (O_1895,N_49899,N_49592);
nor UO_1896 (O_1896,N_49838,N_49716);
and UO_1897 (O_1897,N_49634,N_49933);
or UO_1898 (O_1898,N_49956,N_49828);
or UO_1899 (O_1899,N_49768,N_49638);
and UO_1900 (O_1900,N_49670,N_49906);
and UO_1901 (O_1901,N_49718,N_49816);
and UO_1902 (O_1902,N_49774,N_49840);
nor UO_1903 (O_1903,N_49881,N_49904);
or UO_1904 (O_1904,N_49530,N_49699);
and UO_1905 (O_1905,N_49576,N_49663);
nor UO_1906 (O_1906,N_49667,N_49618);
and UO_1907 (O_1907,N_49734,N_49527);
nand UO_1908 (O_1908,N_49599,N_49646);
or UO_1909 (O_1909,N_49511,N_49548);
nor UO_1910 (O_1910,N_49774,N_49990);
nor UO_1911 (O_1911,N_49721,N_49746);
nor UO_1912 (O_1912,N_49752,N_49955);
and UO_1913 (O_1913,N_49594,N_49527);
and UO_1914 (O_1914,N_49542,N_49620);
xor UO_1915 (O_1915,N_49509,N_49592);
nor UO_1916 (O_1916,N_49866,N_49538);
nor UO_1917 (O_1917,N_49976,N_49558);
or UO_1918 (O_1918,N_49702,N_49514);
and UO_1919 (O_1919,N_49577,N_49560);
and UO_1920 (O_1920,N_49646,N_49869);
nand UO_1921 (O_1921,N_49901,N_49912);
nand UO_1922 (O_1922,N_49580,N_49746);
and UO_1923 (O_1923,N_49506,N_49508);
nand UO_1924 (O_1924,N_49740,N_49809);
nand UO_1925 (O_1925,N_49793,N_49871);
or UO_1926 (O_1926,N_49603,N_49582);
nand UO_1927 (O_1927,N_49702,N_49929);
or UO_1928 (O_1928,N_49761,N_49507);
or UO_1929 (O_1929,N_49741,N_49962);
nand UO_1930 (O_1930,N_49830,N_49647);
xnor UO_1931 (O_1931,N_49911,N_49924);
nand UO_1932 (O_1932,N_49971,N_49913);
or UO_1933 (O_1933,N_49872,N_49609);
or UO_1934 (O_1934,N_49783,N_49829);
or UO_1935 (O_1935,N_49859,N_49778);
and UO_1936 (O_1936,N_49608,N_49808);
or UO_1937 (O_1937,N_49677,N_49574);
xor UO_1938 (O_1938,N_49714,N_49810);
xor UO_1939 (O_1939,N_49986,N_49798);
nor UO_1940 (O_1940,N_49590,N_49889);
and UO_1941 (O_1941,N_49937,N_49816);
or UO_1942 (O_1942,N_49999,N_49623);
nand UO_1943 (O_1943,N_49854,N_49620);
nand UO_1944 (O_1944,N_49957,N_49605);
nor UO_1945 (O_1945,N_49557,N_49663);
nor UO_1946 (O_1946,N_49880,N_49815);
and UO_1947 (O_1947,N_49550,N_49512);
nand UO_1948 (O_1948,N_49698,N_49728);
nor UO_1949 (O_1949,N_49864,N_49897);
nor UO_1950 (O_1950,N_49501,N_49903);
and UO_1951 (O_1951,N_49650,N_49770);
and UO_1952 (O_1952,N_49714,N_49608);
nand UO_1953 (O_1953,N_49991,N_49875);
nand UO_1954 (O_1954,N_49742,N_49617);
nand UO_1955 (O_1955,N_49813,N_49908);
and UO_1956 (O_1956,N_49889,N_49572);
xnor UO_1957 (O_1957,N_49868,N_49748);
or UO_1958 (O_1958,N_49571,N_49555);
or UO_1959 (O_1959,N_49625,N_49676);
and UO_1960 (O_1960,N_49534,N_49726);
and UO_1961 (O_1961,N_49604,N_49614);
nand UO_1962 (O_1962,N_49708,N_49745);
or UO_1963 (O_1963,N_49789,N_49994);
nor UO_1964 (O_1964,N_49820,N_49583);
or UO_1965 (O_1965,N_49937,N_49858);
nand UO_1966 (O_1966,N_49504,N_49813);
nor UO_1967 (O_1967,N_49852,N_49569);
and UO_1968 (O_1968,N_49815,N_49962);
or UO_1969 (O_1969,N_49662,N_49529);
nor UO_1970 (O_1970,N_49920,N_49957);
nand UO_1971 (O_1971,N_49761,N_49892);
or UO_1972 (O_1972,N_49961,N_49845);
nor UO_1973 (O_1973,N_49806,N_49675);
nand UO_1974 (O_1974,N_49514,N_49655);
nor UO_1975 (O_1975,N_49849,N_49648);
and UO_1976 (O_1976,N_49951,N_49561);
nand UO_1977 (O_1977,N_49754,N_49658);
or UO_1978 (O_1978,N_49906,N_49966);
nor UO_1979 (O_1979,N_49665,N_49920);
or UO_1980 (O_1980,N_49756,N_49746);
nand UO_1981 (O_1981,N_49788,N_49598);
nand UO_1982 (O_1982,N_49802,N_49714);
or UO_1983 (O_1983,N_49899,N_49693);
or UO_1984 (O_1984,N_49889,N_49935);
nand UO_1985 (O_1985,N_49983,N_49940);
nor UO_1986 (O_1986,N_49739,N_49515);
or UO_1987 (O_1987,N_49569,N_49792);
or UO_1988 (O_1988,N_49616,N_49718);
xnor UO_1989 (O_1989,N_49506,N_49910);
nor UO_1990 (O_1990,N_49815,N_49809);
or UO_1991 (O_1991,N_49633,N_49821);
nor UO_1992 (O_1992,N_49743,N_49631);
nor UO_1993 (O_1993,N_49967,N_49604);
xnor UO_1994 (O_1994,N_49944,N_49810);
nand UO_1995 (O_1995,N_49586,N_49705);
or UO_1996 (O_1996,N_49685,N_49822);
or UO_1997 (O_1997,N_49981,N_49823);
xor UO_1998 (O_1998,N_49743,N_49751);
nand UO_1999 (O_1999,N_49976,N_49741);
nand UO_2000 (O_2000,N_49676,N_49926);
or UO_2001 (O_2001,N_49521,N_49813);
and UO_2002 (O_2002,N_49693,N_49569);
nand UO_2003 (O_2003,N_49623,N_49773);
or UO_2004 (O_2004,N_49963,N_49670);
and UO_2005 (O_2005,N_49523,N_49611);
nor UO_2006 (O_2006,N_49688,N_49964);
nand UO_2007 (O_2007,N_49868,N_49718);
nand UO_2008 (O_2008,N_49971,N_49978);
and UO_2009 (O_2009,N_49646,N_49566);
nor UO_2010 (O_2010,N_49964,N_49565);
nor UO_2011 (O_2011,N_49826,N_49996);
nor UO_2012 (O_2012,N_49780,N_49533);
nand UO_2013 (O_2013,N_49764,N_49802);
xnor UO_2014 (O_2014,N_49971,N_49690);
and UO_2015 (O_2015,N_49954,N_49782);
or UO_2016 (O_2016,N_49823,N_49613);
and UO_2017 (O_2017,N_49647,N_49606);
xor UO_2018 (O_2018,N_49903,N_49510);
and UO_2019 (O_2019,N_49857,N_49815);
nand UO_2020 (O_2020,N_49896,N_49748);
or UO_2021 (O_2021,N_49934,N_49654);
nor UO_2022 (O_2022,N_49783,N_49741);
nor UO_2023 (O_2023,N_49624,N_49851);
or UO_2024 (O_2024,N_49844,N_49891);
or UO_2025 (O_2025,N_49573,N_49966);
nand UO_2026 (O_2026,N_49899,N_49779);
nand UO_2027 (O_2027,N_49991,N_49536);
and UO_2028 (O_2028,N_49999,N_49821);
or UO_2029 (O_2029,N_49819,N_49853);
and UO_2030 (O_2030,N_49836,N_49958);
and UO_2031 (O_2031,N_49828,N_49565);
nand UO_2032 (O_2032,N_49954,N_49754);
or UO_2033 (O_2033,N_49522,N_49815);
nor UO_2034 (O_2034,N_49761,N_49986);
and UO_2035 (O_2035,N_49953,N_49807);
and UO_2036 (O_2036,N_49505,N_49856);
and UO_2037 (O_2037,N_49911,N_49728);
nand UO_2038 (O_2038,N_49694,N_49576);
and UO_2039 (O_2039,N_49529,N_49730);
and UO_2040 (O_2040,N_49717,N_49815);
and UO_2041 (O_2041,N_49568,N_49918);
nand UO_2042 (O_2042,N_49632,N_49830);
or UO_2043 (O_2043,N_49566,N_49834);
and UO_2044 (O_2044,N_49851,N_49612);
xor UO_2045 (O_2045,N_49932,N_49522);
and UO_2046 (O_2046,N_49917,N_49737);
nand UO_2047 (O_2047,N_49838,N_49967);
and UO_2048 (O_2048,N_49718,N_49839);
nand UO_2049 (O_2049,N_49916,N_49904);
and UO_2050 (O_2050,N_49625,N_49567);
xor UO_2051 (O_2051,N_49553,N_49610);
nor UO_2052 (O_2052,N_49736,N_49747);
xor UO_2053 (O_2053,N_49706,N_49783);
and UO_2054 (O_2054,N_49874,N_49862);
or UO_2055 (O_2055,N_49859,N_49560);
xor UO_2056 (O_2056,N_49560,N_49716);
nand UO_2057 (O_2057,N_49995,N_49606);
and UO_2058 (O_2058,N_49590,N_49990);
nand UO_2059 (O_2059,N_49926,N_49618);
and UO_2060 (O_2060,N_49755,N_49697);
or UO_2061 (O_2061,N_49554,N_49856);
nand UO_2062 (O_2062,N_49696,N_49586);
nand UO_2063 (O_2063,N_49533,N_49785);
nand UO_2064 (O_2064,N_49906,N_49691);
nor UO_2065 (O_2065,N_49708,N_49962);
and UO_2066 (O_2066,N_49629,N_49843);
nand UO_2067 (O_2067,N_49640,N_49977);
nor UO_2068 (O_2068,N_49945,N_49965);
or UO_2069 (O_2069,N_49699,N_49559);
xor UO_2070 (O_2070,N_49516,N_49628);
xnor UO_2071 (O_2071,N_49855,N_49725);
nand UO_2072 (O_2072,N_49975,N_49787);
and UO_2073 (O_2073,N_49811,N_49670);
or UO_2074 (O_2074,N_49844,N_49848);
xor UO_2075 (O_2075,N_49891,N_49601);
nor UO_2076 (O_2076,N_49699,N_49920);
nand UO_2077 (O_2077,N_49731,N_49859);
nor UO_2078 (O_2078,N_49687,N_49510);
nor UO_2079 (O_2079,N_49909,N_49557);
nor UO_2080 (O_2080,N_49650,N_49542);
and UO_2081 (O_2081,N_49671,N_49610);
nand UO_2082 (O_2082,N_49907,N_49797);
nor UO_2083 (O_2083,N_49797,N_49803);
nand UO_2084 (O_2084,N_49809,N_49817);
and UO_2085 (O_2085,N_49539,N_49713);
nand UO_2086 (O_2086,N_49656,N_49845);
xor UO_2087 (O_2087,N_49794,N_49575);
and UO_2088 (O_2088,N_49609,N_49989);
nor UO_2089 (O_2089,N_49865,N_49507);
or UO_2090 (O_2090,N_49599,N_49794);
nor UO_2091 (O_2091,N_49641,N_49751);
xor UO_2092 (O_2092,N_49996,N_49956);
or UO_2093 (O_2093,N_49858,N_49918);
xnor UO_2094 (O_2094,N_49956,N_49910);
nand UO_2095 (O_2095,N_49818,N_49554);
nand UO_2096 (O_2096,N_49632,N_49586);
nor UO_2097 (O_2097,N_49741,N_49804);
or UO_2098 (O_2098,N_49756,N_49904);
nor UO_2099 (O_2099,N_49652,N_49970);
or UO_2100 (O_2100,N_49735,N_49947);
nor UO_2101 (O_2101,N_49771,N_49959);
nor UO_2102 (O_2102,N_49632,N_49929);
nor UO_2103 (O_2103,N_49624,N_49806);
or UO_2104 (O_2104,N_49651,N_49633);
and UO_2105 (O_2105,N_49529,N_49548);
nor UO_2106 (O_2106,N_49994,N_49877);
nand UO_2107 (O_2107,N_49571,N_49516);
nor UO_2108 (O_2108,N_49982,N_49891);
and UO_2109 (O_2109,N_49977,N_49678);
and UO_2110 (O_2110,N_49596,N_49584);
or UO_2111 (O_2111,N_49765,N_49870);
and UO_2112 (O_2112,N_49828,N_49500);
xor UO_2113 (O_2113,N_49759,N_49862);
nor UO_2114 (O_2114,N_49893,N_49596);
xor UO_2115 (O_2115,N_49787,N_49908);
or UO_2116 (O_2116,N_49787,N_49731);
nor UO_2117 (O_2117,N_49949,N_49909);
nand UO_2118 (O_2118,N_49534,N_49500);
and UO_2119 (O_2119,N_49966,N_49804);
xnor UO_2120 (O_2120,N_49886,N_49819);
xnor UO_2121 (O_2121,N_49728,N_49929);
nor UO_2122 (O_2122,N_49541,N_49744);
or UO_2123 (O_2123,N_49962,N_49630);
or UO_2124 (O_2124,N_49601,N_49863);
nor UO_2125 (O_2125,N_49571,N_49692);
nor UO_2126 (O_2126,N_49916,N_49562);
and UO_2127 (O_2127,N_49665,N_49764);
nand UO_2128 (O_2128,N_49870,N_49954);
nor UO_2129 (O_2129,N_49775,N_49520);
nor UO_2130 (O_2130,N_49861,N_49549);
xor UO_2131 (O_2131,N_49827,N_49695);
xnor UO_2132 (O_2132,N_49654,N_49658);
nand UO_2133 (O_2133,N_49999,N_49631);
nand UO_2134 (O_2134,N_49884,N_49957);
or UO_2135 (O_2135,N_49938,N_49959);
nor UO_2136 (O_2136,N_49911,N_49695);
and UO_2137 (O_2137,N_49891,N_49997);
or UO_2138 (O_2138,N_49970,N_49668);
nand UO_2139 (O_2139,N_49993,N_49698);
and UO_2140 (O_2140,N_49538,N_49664);
and UO_2141 (O_2141,N_49996,N_49857);
nand UO_2142 (O_2142,N_49767,N_49609);
or UO_2143 (O_2143,N_49924,N_49806);
nand UO_2144 (O_2144,N_49609,N_49612);
nor UO_2145 (O_2145,N_49867,N_49802);
nor UO_2146 (O_2146,N_49675,N_49955);
or UO_2147 (O_2147,N_49895,N_49694);
or UO_2148 (O_2148,N_49563,N_49779);
nor UO_2149 (O_2149,N_49837,N_49960);
nor UO_2150 (O_2150,N_49716,N_49822);
nand UO_2151 (O_2151,N_49566,N_49572);
nand UO_2152 (O_2152,N_49759,N_49888);
nand UO_2153 (O_2153,N_49723,N_49654);
or UO_2154 (O_2154,N_49978,N_49899);
or UO_2155 (O_2155,N_49882,N_49731);
nor UO_2156 (O_2156,N_49770,N_49670);
and UO_2157 (O_2157,N_49703,N_49665);
and UO_2158 (O_2158,N_49762,N_49809);
and UO_2159 (O_2159,N_49875,N_49932);
nor UO_2160 (O_2160,N_49877,N_49658);
nor UO_2161 (O_2161,N_49783,N_49701);
or UO_2162 (O_2162,N_49929,N_49813);
nor UO_2163 (O_2163,N_49765,N_49733);
xnor UO_2164 (O_2164,N_49968,N_49791);
and UO_2165 (O_2165,N_49875,N_49709);
xnor UO_2166 (O_2166,N_49727,N_49819);
xor UO_2167 (O_2167,N_49605,N_49826);
nor UO_2168 (O_2168,N_49541,N_49568);
and UO_2169 (O_2169,N_49987,N_49850);
xnor UO_2170 (O_2170,N_49630,N_49819);
nor UO_2171 (O_2171,N_49654,N_49735);
nor UO_2172 (O_2172,N_49876,N_49896);
nor UO_2173 (O_2173,N_49829,N_49885);
nor UO_2174 (O_2174,N_49790,N_49845);
nor UO_2175 (O_2175,N_49574,N_49774);
or UO_2176 (O_2176,N_49791,N_49812);
nand UO_2177 (O_2177,N_49767,N_49603);
nor UO_2178 (O_2178,N_49983,N_49593);
and UO_2179 (O_2179,N_49746,N_49867);
nor UO_2180 (O_2180,N_49555,N_49867);
or UO_2181 (O_2181,N_49540,N_49828);
and UO_2182 (O_2182,N_49822,N_49734);
nor UO_2183 (O_2183,N_49867,N_49609);
nand UO_2184 (O_2184,N_49544,N_49976);
nand UO_2185 (O_2185,N_49640,N_49535);
nor UO_2186 (O_2186,N_49839,N_49535);
xor UO_2187 (O_2187,N_49501,N_49507);
nand UO_2188 (O_2188,N_49779,N_49657);
nor UO_2189 (O_2189,N_49903,N_49620);
nor UO_2190 (O_2190,N_49843,N_49834);
or UO_2191 (O_2191,N_49649,N_49779);
nor UO_2192 (O_2192,N_49520,N_49671);
nor UO_2193 (O_2193,N_49884,N_49980);
xor UO_2194 (O_2194,N_49603,N_49635);
nor UO_2195 (O_2195,N_49841,N_49754);
nand UO_2196 (O_2196,N_49753,N_49759);
and UO_2197 (O_2197,N_49754,N_49992);
and UO_2198 (O_2198,N_49984,N_49962);
nand UO_2199 (O_2199,N_49859,N_49926);
or UO_2200 (O_2200,N_49804,N_49601);
or UO_2201 (O_2201,N_49532,N_49548);
xnor UO_2202 (O_2202,N_49561,N_49638);
nand UO_2203 (O_2203,N_49799,N_49900);
nor UO_2204 (O_2204,N_49522,N_49684);
nor UO_2205 (O_2205,N_49750,N_49773);
nor UO_2206 (O_2206,N_49501,N_49828);
nor UO_2207 (O_2207,N_49735,N_49533);
or UO_2208 (O_2208,N_49860,N_49517);
nand UO_2209 (O_2209,N_49974,N_49985);
xor UO_2210 (O_2210,N_49643,N_49796);
nand UO_2211 (O_2211,N_49972,N_49778);
xnor UO_2212 (O_2212,N_49757,N_49554);
xnor UO_2213 (O_2213,N_49799,N_49869);
nor UO_2214 (O_2214,N_49589,N_49501);
nand UO_2215 (O_2215,N_49919,N_49550);
xor UO_2216 (O_2216,N_49799,N_49865);
and UO_2217 (O_2217,N_49925,N_49591);
and UO_2218 (O_2218,N_49927,N_49684);
nor UO_2219 (O_2219,N_49660,N_49815);
nand UO_2220 (O_2220,N_49547,N_49992);
or UO_2221 (O_2221,N_49612,N_49852);
xnor UO_2222 (O_2222,N_49564,N_49936);
nand UO_2223 (O_2223,N_49570,N_49603);
nor UO_2224 (O_2224,N_49586,N_49859);
and UO_2225 (O_2225,N_49738,N_49830);
and UO_2226 (O_2226,N_49998,N_49923);
xor UO_2227 (O_2227,N_49988,N_49838);
nand UO_2228 (O_2228,N_49917,N_49951);
nand UO_2229 (O_2229,N_49806,N_49534);
nand UO_2230 (O_2230,N_49823,N_49733);
nand UO_2231 (O_2231,N_49535,N_49670);
nor UO_2232 (O_2232,N_49531,N_49796);
nand UO_2233 (O_2233,N_49872,N_49765);
or UO_2234 (O_2234,N_49893,N_49744);
and UO_2235 (O_2235,N_49733,N_49840);
or UO_2236 (O_2236,N_49798,N_49849);
nor UO_2237 (O_2237,N_49878,N_49939);
nand UO_2238 (O_2238,N_49660,N_49547);
and UO_2239 (O_2239,N_49956,N_49600);
or UO_2240 (O_2240,N_49998,N_49983);
nor UO_2241 (O_2241,N_49691,N_49795);
nand UO_2242 (O_2242,N_49945,N_49967);
nand UO_2243 (O_2243,N_49982,N_49835);
nand UO_2244 (O_2244,N_49697,N_49634);
xnor UO_2245 (O_2245,N_49877,N_49850);
nand UO_2246 (O_2246,N_49686,N_49693);
or UO_2247 (O_2247,N_49968,N_49867);
and UO_2248 (O_2248,N_49536,N_49939);
nor UO_2249 (O_2249,N_49996,N_49644);
nand UO_2250 (O_2250,N_49567,N_49824);
nor UO_2251 (O_2251,N_49503,N_49705);
or UO_2252 (O_2252,N_49574,N_49638);
or UO_2253 (O_2253,N_49815,N_49541);
xor UO_2254 (O_2254,N_49877,N_49807);
nand UO_2255 (O_2255,N_49836,N_49544);
nor UO_2256 (O_2256,N_49658,N_49595);
nand UO_2257 (O_2257,N_49646,N_49513);
nand UO_2258 (O_2258,N_49827,N_49592);
nand UO_2259 (O_2259,N_49790,N_49890);
nor UO_2260 (O_2260,N_49800,N_49779);
or UO_2261 (O_2261,N_49876,N_49871);
or UO_2262 (O_2262,N_49588,N_49976);
nor UO_2263 (O_2263,N_49683,N_49978);
and UO_2264 (O_2264,N_49780,N_49540);
or UO_2265 (O_2265,N_49510,N_49953);
nand UO_2266 (O_2266,N_49758,N_49889);
xnor UO_2267 (O_2267,N_49524,N_49827);
nand UO_2268 (O_2268,N_49986,N_49675);
or UO_2269 (O_2269,N_49542,N_49929);
or UO_2270 (O_2270,N_49618,N_49702);
nor UO_2271 (O_2271,N_49745,N_49989);
nand UO_2272 (O_2272,N_49870,N_49715);
nor UO_2273 (O_2273,N_49723,N_49674);
nor UO_2274 (O_2274,N_49600,N_49842);
or UO_2275 (O_2275,N_49580,N_49657);
nand UO_2276 (O_2276,N_49651,N_49770);
or UO_2277 (O_2277,N_49762,N_49561);
nor UO_2278 (O_2278,N_49529,N_49990);
nor UO_2279 (O_2279,N_49894,N_49694);
xnor UO_2280 (O_2280,N_49957,N_49544);
nor UO_2281 (O_2281,N_49873,N_49773);
or UO_2282 (O_2282,N_49813,N_49827);
nor UO_2283 (O_2283,N_49812,N_49575);
or UO_2284 (O_2284,N_49571,N_49985);
nand UO_2285 (O_2285,N_49830,N_49674);
nand UO_2286 (O_2286,N_49797,N_49616);
xnor UO_2287 (O_2287,N_49757,N_49939);
or UO_2288 (O_2288,N_49901,N_49615);
and UO_2289 (O_2289,N_49709,N_49678);
nor UO_2290 (O_2290,N_49565,N_49756);
or UO_2291 (O_2291,N_49952,N_49951);
and UO_2292 (O_2292,N_49719,N_49777);
nand UO_2293 (O_2293,N_49881,N_49741);
or UO_2294 (O_2294,N_49761,N_49684);
nand UO_2295 (O_2295,N_49795,N_49841);
xor UO_2296 (O_2296,N_49711,N_49615);
and UO_2297 (O_2297,N_49518,N_49677);
and UO_2298 (O_2298,N_49743,N_49904);
nor UO_2299 (O_2299,N_49958,N_49644);
nor UO_2300 (O_2300,N_49681,N_49963);
nor UO_2301 (O_2301,N_49633,N_49577);
and UO_2302 (O_2302,N_49546,N_49509);
nand UO_2303 (O_2303,N_49972,N_49737);
nor UO_2304 (O_2304,N_49986,N_49836);
nand UO_2305 (O_2305,N_49751,N_49798);
nand UO_2306 (O_2306,N_49579,N_49823);
nor UO_2307 (O_2307,N_49607,N_49548);
and UO_2308 (O_2308,N_49713,N_49566);
xor UO_2309 (O_2309,N_49742,N_49787);
or UO_2310 (O_2310,N_49828,N_49877);
xnor UO_2311 (O_2311,N_49857,N_49859);
nand UO_2312 (O_2312,N_49694,N_49665);
or UO_2313 (O_2313,N_49724,N_49794);
nor UO_2314 (O_2314,N_49593,N_49541);
nor UO_2315 (O_2315,N_49883,N_49946);
nand UO_2316 (O_2316,N_49914,N_49814);
xor UO_2317 (O_2317,N_49772,N_49561);
nor UO_2318 (O_2318,N_49830,N_49858);
and UO_2319 (O_2319,N_49841,N_49595);
or UO_2320 (O_2320,N_49552,N_49726);
and UO_2321 (O_2321,N_49936,N_49647);
and UO_2322 (O_2322,N_49501,N_49835);
and UO_2323 (O_2323,N_49783,N_49846);
and UO_2324 (O_2324,N_49647,N_49584);
or UO_2325 (O_2325,N_49754,N_49945);
nand UO_2326 (O_2326,N_49994,N_49639);
or UO_2327 (O_2327,N_49636,N_49597);
xnor UO_2328 (O_2328,N_49692,N_49842);
xnor UO_2329 (O_2329,N_49936,N_49957);
or UO_2330 (O_2330,N_49852,N_49596);
xnor UO_2331 (O_2331,N_49914,N_49633);
nand UO_2332 (O_2332,N_49755,N_49945);
nand UO_2333 (O_2333,N_49928,N_49836);
or UO_2334 (O_2334,N_49904,N_49636);
or UO_2335 (O_2335,N_49589,N_49987);
nor UO_2336 (O_2336,N_49518,N_49827);
or UO_2337 (O_2337,N_49532,N_49666);
nor UO_2338 (O_2338,N_49689,N_49772);
or UO_2339 (O_2339,N_49589,N_49650);
nor UO_2340 (O_2340,N_49635,N_49602);
and UO_2341 (O_2341,N_49777,N_49576);
xor UO_2342 (O_2342,N_49941,N_49875);
nor UO_2343 (O_2343,N_49904,N_49683);
nor UO_2344 (O_2344,N_49512,N_49908);
nor UO_2345 (O_2345,N_49837,N_49624);
and UO_2346 (O_2346,N_49814,N_49524);
nand UO_2347 (O_2347,N_49973,N_49514);
nand UO_2348 (O_2348,N_49587,N_49750);
and UO_2349 (O_2349,N_49543,N_49756);
or UO_2350 (O_2350,N_49945,N_49757);
or UO_2351 (O_2351,N_49671,N_49925);
xnor UO_2352 (O_2352,N_49750,N_49540);
or UO_2353 (O_2353,N_49541,N_49797);
nand UO_2354 (O_2354,N_49884,N_49600);
or UO_2355 (O_2355,N_49775,N_49843);
or UO_2356 (O_2356,N_49701,N_49562);
nand UO_2357 (O_2357,N_49753,N_49889);
xor UO_2358 (O_2358,N_49805,N_49633);
or UO_2359 (O_2359,N_49915,N_49659);
nand UO_2360 (O_2360,N_49694,N_49611);
or UO_2361 (O_2361,N_49893,N_49547);
nand UO_2362 (O_2362,N_49976,N_49542);
and UO_2363 (O_2363,N_49927,N_49966);
and UO_2364 (O_2364,N_49670,N_49550);
nor UO_2365 (O_2365,N_49934,N_49831);
nor UO_2366 (O_2366,N_49936,N_49873);
or UO_2367 (O_2367,N_49677,N_49623);
or UO_2368 (O_2368,N_49656,N_49637);
nand UO_2369 (O_2369,N_49644,N_49930);
nor UO_2370 (O_2370,N_49726,N_49960);
nor UO_2371 (O_2371,N_49624,N_49981);
and UO_2372 (O_2372,N_49827,N_49581);
xor UO_2373 (O_2373,N_49705,N_49960);
or UO_2374 (O_2374,N_49974,N_49994);
and UO_2375 (O_2375,N_49702,N_49531);
and UO_2376 (O_2376,N_49586,N_49752);
and UO_2377 (O_2377,N_49776,N_49639);
and UO_2378 (O_2378,N_49840,N_49982);
nor UO_2379 (O_2379,N_49772,N_49513);
and UO_2380 (O_2380,N_49719,N_49995);
and UO_2381 (O_2381,N_49625,N_49556);
nand UO_2382 (O_2382,N_49512,N_49984);
nor UO_2383 (O_2383,N_49711,N_49837);
xnor UO_2384 (O_2384,N_49875,N_49776);
nand UO_2385 (O_2385,N_49539,N_49803);
or UO_2386 (O_2386,N_49985,N_49862);
and UO_2387 (O_2387,N_49877,N_49977);
nand UO_2388 (O_2388,N_49819,N_49602);
nand UO_2389 (O_2389,N_49774,N_49989);
or UO_2390 (O_2390,N_49500,N_49783);
nor UO_2391 (O_2391,N_49522,N_49863);
nor UO_2392 (O_2392,N_49541,N_49944);
or UO_2393 (O_2393,N_49783,N_49751);
and UO_2394 (O_2394,N_49795,N_49677);
and UO_2395 (O_2395,N_49984,N_49592);
nand UO_2396 (O_2396,N_49621,N_49702);
nor UO_2397 (O_2397,N_49987,N_49801);
nor UO_2398 (O_2398,N_49770,N_49641);
nor UO_2399 (O_2399,N_49931,N_49818);
and UO_2400 (O_2400,N_49825,N_49793);
or UO_2401 (O_2401,N_49894,N_49634);
nand UO_2402 (O_2402,N_49693,N_49715);
or UO_2403 (O_2403,N_49681,N_49771);
xnor UO_2404 (O_2404,N_49826,N_49755);
and UO_2405 (O_2405,N_49698,N_49979);
and UO_2406 (O_2406,N_49726,N_49911);
nor UO_2407 (O_2407,N_49668,N_49542);
and UO_2408 (O_2408,N_49830,N_49888);
nor UO_2409 (O_2409,N_49833,N_49804);
nand UO_2410 (O_2410,N_49769,N_49873);
nand UO_2411 (O_2411,N_49836,N_49682);
nand UO_2412 (O_2412,N_49999,N_49767);
nor UO_2413 (O_2413,N_49860,N_49696);
or UO_2414 (O_2414,N_49710,N_49556);
or UO_2415 (O_2415,N_49563,N_49845);
nor UO_2416 (O_2416,N_49567,N_49637);
nor UO_2417 (O_2417,N_49915,N_49637);
or UO_2418 (O_2418,N_49993,N_49602);
nand UO_2419 (O_2419,N_49506,N_49792);
xor UO_2420 (O_2420,N_49883,N_49690);
and UO_2421 (O_2421,N_49977,N_49956);
and UO_2422 (O_2422,N_49853,N_49906);
or UO_2423 (O_2423,N_49695,N_49754);
or UO_2424 (O_2424,N_49510,N_49569);
xnor UO_2425 (O_2425,N_49609,N_49878);
and UO_2426 (O_2426,N_49524,N_49731);
nor UO_2427 (O_2427,N_49704,N_49884);
xnor UO_2428 (O_2428,N_49576,N_49949);
nor UO_2429 (O_2429,N_49834,N_49527);
nor UO_2430 (O_2430,N_49898,N_49994);
or UO_2431 (O_2431,N_49682,N_49648);
and UO_2432 (O_2432,N_49983,N_49710);
and UO_2433 (O_2433,N_49791,N_49695);
nand UO_2434 (O_2434,N_49526,N_49627);
or UO_2435 (O_2435,N_49782,N_49834);
and UO_2436 (O_2436,N_49738,N_49939);
nand UO_2437 (O_2437,N_49736,N_49548);
and UO_2438 (O_2438,N_49750,N_49735);
nor UO_2439 (O_2439,N_49681,N_49651);
nor UO_2440 (O_2440,N_49781,N_49565);
nand UO_2441 (O_2441,N_49744,N_49859);
nor UO_2442 (O_2442,N_49942,N_49595);
nor UO_2443 (O_2443,N_49771,N_49677);
xnor UO_2444 (O_2444,N_49531,N_49652);
and UO_2445 (O_2445,N_49754,N_49726);
and UO_2446 (O_2446,N_49825,N_49936);
nand UO_2447 (O_2447,N_49813,N_49779);
and UO_2448 (O_2448,N_49839,N_49734);
or UO_2449 (O_2449,N_49880,N_49876);
nand UO_2450 (O_2450,N_49534,N_49751);
nand UO_2451 (O_2451,N_49923,N_49582);
and UO_2452 (O_2452,N_49650,N_49962);
or UO_2453 (O_2453,N_49648,N_49802);
and UO_2454 (O_2454,N_49716,N_49650);
or UO_2455 (O_2455,N_49910,N_49782);
or UO_2456 (O_2456,N_49931,N_49833);
nor UO_2457 (O_2457,N_49749,N_49950);
and UO_2458 (O_2458,N_49869,N_49928);
nand UO_2459 (O_2459,N_49559,N_49867);
nor UO_2460 (O_2460,N_49946,N_49708);
or UO_2461 (O_2461,N_49740,N_49765);
nand UO_2462 (O_2462,N_49606,N_49696);
nand UO_2463 (O_2463,N_49623,N_49847);
and UO_2464 (O_2464,N_49682,N_49893);
or UO_2465 (O_2465,N_49545,N_49714);
xnor UO_2466 (O_2466,N_49724,N_49967);
nand UO_2467 (O_2467,N_49770,N_49986);
and UO_2468 (O_2468,N_49849,N_49645);
nor UO_2469 (O_2469,N_49526,N_49994);
and UO_2470 (O_2470,N_49857,N_49933);
nor UO_2471 (O_2471,N_49591,N_49702);
and UO_2472 (O_2472,N_49511,N_49999);
or UO_2473 (O_2473,N_49620,N_49910);
or UO_2474 (O_2474,N_49615,N_49687);
or UO_2475 (O_2475,N_49706,N_49642);
nor UO_2476 (O_2476,N_49667,N_49519);
and UO_2477 (O_2477,N_49906,N_49648);
nand UO_2478 (O_2478,N_49758,N_49532);
nand UO_2479 (O_2479,N_49728,N_49619);
or UO_2480 (O_2480,N_49992,N_49605);
or UO_2481 (O_2481,N_49809,N_49832);
xor UO_2482 (O_2482,N_49764,N_49777);
nor UO_2483 (O_2483,N_49814,N_49833);
nor UO_2484 (O_2484,N_49993,N_49821);
and UO_2485 (O_2485,N_49612,N_49868);
or UO_2486 (O_2486,N_49812,N_49915);
xnor UO_2487 (O_2487,N_49832,N_49668);
xnor UO_2488 (O_2488,N_49637,N_49947);
xnor UO_2489 (O_2489,N_49582,N_49982);
nand UO_2490 (O_2490,N_49796,N_49963);
and UO_2491 (O_2491,N_49819,N_49617);
and UO_2492 (O_2492,N_49523,N_49877);
nand UO_2493 (O_2493,N_49505,N_49949);
nand UO_2494 (O_2494,N_49918,N_49739);
nor UO_2495 (O_2495,N_49820,N_49669);
nand UO_2496 (O_2496,N_49732,N_49740);
and UO_2497 (O_2497,N_49711,N_49533);
nand UO_2498 (O_2498,N_49514,N_49781);
nand UO_2499 (O_2499,N_49919,N_49784);
or UO_2500 (O_2500,N_49860,N_49825);
nor UO_2501 (O_2501,N_49535,N_49924);
and UO_2502 (O_2502,N_49944,N_49870);
and UO_2503 (O_2503,N_49541,N_49700);
and UO_2504 (O_2504,N_49894,N_49584);
and UO_2505 (O_2505,N_49738,N_49548);
and UO_2506 (O_2506,N_49655,N_49937);
or UO_2507 (O_2507,N_49805,N_49990);
nand UO_2508 (O_2508,N_49806,N_49670);
nand UO_2509 (O_2509,N_49864,N_49642);
nand UO_2510 (O_2510,N_49649,N_49562);
or UO_2511 (O_2511,N_49800,N_49964);
or UO_2512 (O_2512,N_49926,N_49823);
nor UO_2513 (O_2513,N_49760,N_49523);
and UO_2514 (O_2514,N_49964,N_49566);
nor UO_2515 (O_2515,N_49673,N_49935);
nor UO_2516 (O_2516,N_49717,N_49991);
nand UO_2517 (O_2517,N_49942,N_49776);
and UO_2518 (O_2518,N_49512,N_49705);
nor UO_2519 (O_2519,N_49787,N_49542);
nor UO_2520 (O_2520,N_49773,N_49682);
and UO_2521 (O_2521,N_49633,N_49907);
nor UO_2522 (O_2522,N_49932,N_49616);
and UO_2523 (O_2523,N_49706,N_49914);
xnor UO_2524 (O_2524,N_49541,N_49505);
xor UO_2525 (O_2525,N_49584,N_49818);
nor UO_2526 (O_2526,N_49600,N_49992);
nor UO_2527 (O_2527,N_49922,N_49611);
or UO_2528 (O_2528,N_49584,N_49750);
or UO_2529 (O_2529,N_49730,N_49732);
xnor UO_2530 (O_2530,N_49793,N_49810);
nor UO_2531 (O_2531,N_49526,N_49803);
or UO_2532 (O_2532,N_49731,N_49865);
or UO_2533 (O_2533,N_49796,N_49770);
nand UO_2534 (O_2534,N_49987,N_49761);
nor UO_2535 (O_2535,N_49911,N_49780);
nand UO_2536 (O_2536,N_49661,N_49734);
or UO_2537 (O_2537,N_49701,N_49706);
nor UO_2538 (O_2538,N_49511,N_49812);
nand UO_2539 (O_2539,N_49600,N_49877);
and UO_2540 (O_2540,N_49525,N_49884);
or UO_2541 (O_2541,N_49707,N_49772);
and UO_2542 (O_2542,N_49960,N_49792);
or UO_2543 (O_2543,N_49827,N_49781);
nand UO_2544 (O_2544,N_49766,N_49814);
nor UO_2545 (O_2545,N_49948,N_49783);
or UO_2546 (O_2546,N_49731,N_49532);
and UO_2547 (O_2547,N_49729,N_49541);
or UO_2548 (O_2548,N_49673,N_49949);
nor UO_2549 (O_2549,N_49954,N_49922);
nand UO_2550 (O_2550,N_49681,N_49941);
or UO_2551 (O_2551,N_49684,N_49605);
and UO_2552 (O_2552,N_49955,N_49963);
nand UO_2553 (O_2553,N_49654,N_49724);
nor UO_2554 (O_2554,N_49909,N_49604);
nand UO_2555 (O_2555,N_49773,N_49566);
nand UO_2556 (O_2556,N_49898,N_49545);
and UO_2557 (O_2557,N_49921,N_49700);
or UO_2558 (O_2558,N_49876,N_49579);
nand UO_2559 (O_2559,N_49741,N_49714);
and UO_2560 (O_2560,N_49535,N_49953);
xnor UO_2561 (O_2561,N_49823,N_49890);
and UO_2562 (O_2562,N_49596,N_49869);
or UO_2563 (O_2563,N_49760,N_49566);
or UO_2564 (O_2564,N_49987,N_49871);
and UO_2565 (O_2565,N_49743,N_49754);
and UO_2566 (O_2566,N_49915,N_49531);
xor UO_2567 (O_2567,N_49644,N_49630);
nor UO_2568 (O_2568,N_49814,N_49924);
and UO_2569 (O_2569,N_49985,N_49576);
nand UO_2570 (O_2570,N_49732,N_49981);
or UO_2571 (O_2571,N_49818,N_49524);
nor UO_2572 (O_2572,N_49929,N_49540);
or UO_2573 (O_2573,N_49864,N_49787);
or UO_2574 (O_2574,N_49924,N_49766);
nand UO_2575 (O_2575,N_49678,N_49536);
nand UO_2576 (O_2576,N_49781,N_49515);
or UO_2577 (O_2577,N_49980,N_49885);
xor UO_2578 (O_2578,N_49674,N_49823);
xnor UO_2579 (O_2579,N_49997,N_49850);
and UO_2580 (O_2580,N_49867,N_49963);
nand UO_2581 (O_2581,N_49648,N_49782);
nor UO_2582 (O_2582,N_49863,N_49846);
nand UO_2583 (O_2583,N_49646,N_49959);
and UO_2584 (O_2584,N_49677,N_49880);
xnor UO_2585 (O_2585,N_49881,N_49908);
or UO_2586 (O_2586,N_49883,N_49791);
and UO_2587 (O_2587,N_49885,N_49748);
and UO_2588 (O_2588,N_49676,N_49795);
nand UO_2589 (O_2589,N_49689,N_49591);
nor UO_2590 (O_2590,N_49569,N_49798);
or UO_2591 (O_2591,N_49848,N_49882);
nand UO_2592 (O_2592,N_49826,N_49585);
and UO_2593 (O_2593,N_49995,N_49718);
nand UO_2594 (O_2594,N_49739,N_49929);
or UO_2595 (O_2595,N_49772,N_49964);
nor UO_2596 (O_2596,N_49799,N_49886);
nand UO_2597 (O_2597,N_49853,N_49773);
and UO_2598 (O_2598,N_49956,N_49676);
nor UO_2599 (O_2599,N_49796,N_49578);
xnor UO_2600 (O_2600,N_49701,N_49804);
or UO_2601 (O_2601,N_49905,N_49926);
nor UO_2602 (O_2602,N_49618,N_49621);
or UO_2603 (O_2603,N_49664,N_49808);
or UO_2604 (O_2604,N_49972,N_49872);
or UO_2605 (O_2605,N_49645,N_49752);
nor UO_2606 (O_2606,N_49686,N_49643);
or UO_2607 (O_2607,N_49708,N_49944);
or UO_2608 (O_2608,N_49525,N_49632);
or UO_2609 (O_2609,N_49976,N_49649);
or UO_2610 (O_2610,N_49856,N_49584);
nand UO_2611 (O_2611,N_49673,N_49589);
nand UO_2612 (O_2612,N_49955,N_49805);
nand UO_2613 (O_2613,N_49659,N_49925);
or UO_2614 (O_2614,N_49802,N_49771);
or UO_2615 (O_2615,N_49915,N_49886);
nor UO_2616 (O_2616,N_49837,N_49831);
xnor UO_2617 (O_2617,N_49645,N_49681);
and UO_2618 (O_2618,N_49515,N_49714);
xor UO_2619 (O_2619,N_49982,N_49530);
and UO_2620 (O_2620,N_49661,N_49695);
and UO_2621 (O_2621,N_49663,N_49502);
or UO_2622 (O_2622,N_49568,N_49759);
or UO_2623 (O_2623,N_49794,N_49786);
nand UO_2624 (O_2624,N_49610,N_49774);
xor UO_2625 (O_2625,N_49693,N_49866);
nand UO_2626 (O_2626,N_49563,N_49997);
and UO_2627 (O_2627,N_49652,N_49879);
nand UO_2628 (O_2628,N_49624,N_49927);
nand UO_2629 (O_2629,N_49515,N_49785);
nand UO_2630 (O_2630,N_49892,N_49676);
xor UO_2631 (O_2631,N_49950,N_49854);
or UO_2632 (O_2632,N_49667,N_49862);
xnor UO_2633 (O_2633,N_49914,N_49828);
xor UO_2634 (O_2634,N_49765,N_49952);
xor UO_2635 (O_2635,N_49805,N_49947);
or UO_2636 (O_2636,N_49762,N_49649);
and UO_2637 (O_2637,N_49511,N_49904);
nor UO_2638 (O_2638,N_49573,N_49769);
or UO_2639 (O_2639,N_49881,N_49539);
and UO_2640 (O_2640,N_49776,N_49857);
nand UO_2641 (O_2641,N_49767,N_49943);
and UO_2642 (O_2642,N_49585,N_49683);
xor UO_2643 (O_2643,N_49510,N_49796);
or UO_2644 (O_2644,N_49658,N_49605);
nand UO_2645 (O_2645,N_49947,N_49912);
nand UO_2646 (O_2646,N_49744,N_49780);
nor UO_2647 (O_2647,N_49525,N_49762);
or UO_2648 (O_2648,N_49788,N_49825);
nand UO_2649 (O_2649,N_49954,N_49785);
or UO_2650 (O_2650,N_49642,N_49798);
and UO_2651 (O_2651,N_49836,N_49914);
xor UO_2652 (O_2652,N_49554,N_49822);
xnor UO_2653 (O_2653,N_49562,N_49527);
nand UO_2654 (O_2654,N_49551,N_49688);
nand UO_2655 (O_2655,N_49621,N_49985);
nor UO_2656 (O_2656,N_49982,N_49825);
and UO_2657 (O_2657,N_49624,N_49877);
and UO_2658 (O_2658,N_49592,N_49634);
and UO_2659 (O_2659,N_49569,N_49533);
or UO_2660 (O_2660,N_49839,N_49903);
xor UO_2661 (O_2661,N_49504,N_49853);
and UO_2662 (O_2662,N_49745,N_49793);
or UO_2663 (O_2663,N_49916,N_49884);
and UO_2664 (O_2664,N_49878,N_49960);
and UO_2665 (O_2665,N_49740,N_49795);
nor UO_2666 (O_2666,N_49546,N_49944);
nand UO_2667 (O_2667,N_49535,N_49586);
nand UO_2668 (O_2668,N_49658,N_49581);
nand UO_2669 (O_2669,N_49730,N_49518);
nor UO_2670 (O_2670,N_49978,N_49596);
and UO_2671 (O_2671,N_49576,N_49767);
or UO_2672 (O_2672,N_49706,N_49977);
or UO_2673 (O_2673,N_49900,N_49952);
nor UO_2674 (O_2674,N_49644,N_49614);
and UO_2675 (O_2675,N_49849,N_49931);
nand UO_2676 (O_2676,N_49571,N_49915);
or UO_2677 (O_2677,N_49997,N_49735);
or UO_2678 (O_2678,N_49577,N_49524);
nor UO_2679 (O_2679,N_49884,N_49914);
and UO_2680 (O_2680,N_49782,N_49887);
and UO_2681 (O_2681,N_49660,N_49636);
or UO_2682 (O_2682,N_49789,N_49616);
or UO_2683 (O_2683,N_49635,N_49888);
and UO_2684 (O_2684,N_49888,N_49716);
and UO_2685 (O_2685,N_49659,N_49933);
or UO_2686 (O_2686,N_49833,N_49679);
xor UO_2687 (O_2687,N_49685,N_49900);
and UO_2688 (O_2688,N_49548,N_49886);
xor UO_2689 (O_2689,N_49742,N_49914);
nand UO_2690 (O_2690,N_49944,N_49622);
and UO_2691 (O_2691,N_49691,N_49714);
nor UO_2692 (O_2692,N_49901,N_49856);
or UO_2693 (O_2693,N_49684,N_49652);
and UO_2694 (O_2694,N_49905,N_49934);
or UO_2695 (O_2695,N_49747,N_49911);
nor UO_2696 (O_2696,N_49835,N_49896);
nor UO_2697 (O_2697,N_49594,N_49689);
nor UO_2698 (O_2698,N_49831,N_49779);
nor UO_2699 (O_2699,N_49666,N_49580);
and UO_2700 (O_2700,N_49725,N_49739);
nor UO_2701 (O_2701,N_49942,N_49860);
or UO_2702 (O_2702,N_49728,N_49933);
nor UO_2703 (O_2703,N_49754,N_49918);
xnor UO_2704 (O_2704,N_49749,N_49782);
nand UO_2705 (O_2705,N_49645,N_49959);
nand UO_2706 (O_2706,N_49770,N_49768);
nor UO_2707 (O_2707,N_49788,N_49565);
xor UO_2708 (O_2708,N_49768,N_49664);
nand UO_2709 (O_2709,N_49817,N_49672);
nand UO_2710 (O_2710,N_49678,N_49882);
and UO_2711 (O_2711,N_49892,N_49801);
nor UO_2712 (O_2712,N_49966,N_49611);
and UO_2713 (O_2713,N_49555,N_49554);
nor UO_2714 (O_2714,N_49580,N_49561);
or UO_2715 (O_2715,N_49721,N_49838);
and UO_2716 (O_2716,N_49714,N_49910);
nand UO_2717 (O_2717,N_49930,N_49730);
nor UO_2718 (O_2718,N_49643,N_49733);
nor UO_2719 (O_2719,N_49809,N_49732);
or UO_2720 (O_2720,N_49715,N_49735);
and UO_2721 (O_2721,N_49638,N_49550);
or UO_2722 (O_2722,N_49549,N_49592);
and UO_2723 (O_2723,N_49914,N_49637);
nor UO_2724 (O_2724,N_49823,N_49864);
nor UO_2725 (O_2725,N_49511,N_49782);
and UO_2726 (O_2726,N_49943,N_49505);
nand UO_2727 (O_2727,N_49682,N_49976);
nor UO_2728 (O_2728,N_49530,N_49570);
or UO_2729 (O_2729,N_49818,N_49968);
nand UO_2730 (O_2730,N_49888,N_49815);
and UO_2731 (O_2731,N_49650,N_49731);
or UO_2732 (O_2732,N_49768,N_49754);
or UO_2733 (O_2733,N_49855,N_49591);
nor UO_2734 (O_2734,N_49541,N_49545);
nand UO_2735 (O_2735,N_49752,N_49873);
nor UO_2736 (O_2736,N_49667,N_49514);
and UO_2737 (O_2737,N_49821,N_49782);
and UO_2738 (O_2738,N_49778,N_49969);
nor UO_2739 (O_2739,N_49824,N_49611);
or UO_2740 (O_2740,N_49989,N_49928);
or UO_2741 (O_2741,N_49700,N_49608);
and UO_2742 (O_2742,N_49973,N_49768);
nor UO_2743 (O_2743,N_49664,N_49921);
and UO_2744 (O_2744,N_49960,N_49675);
or UO_2745 (O_2745,N_49876,N_49520);
xnor UO_2746 (O_2746,N_49666,N_49539);
xor UO_2747 (O_2747,N_49842,N_49941);
and UO_2748 (O_2748,N_49505,N_49930);
xor UO_2749 (O_2749,N_49989,N_49539);
or UO_2750 (O_2750,N_49636,N_49659);
and UO_2751 (O_2751,N_49736,N_49960);
nand UO_2752 (O_2752,N_49566,N_49676);
nor UO_2753 (O_2753,N_49617,N_49972);
nand UO_2754 (O_2754,N_49861,N_49888);
or UO_2755 (O_2755,N_49744,N_49583);
and UO_2756 (O_2756,N_49881,N_49887);
or UO_2757 (O_2757,N_49678,N_49938);
nand UO_2758 (O_2758,N_49542,N_49854);
nor UO_2759 (O_2759,N_49772,N_49751);
nand UO_2760 (O_2760,N_49931,N_49829);
or UO_2761 (O_2761,N_49636,N_49922);
xnor UO_2762 (O_2762,N_49852,N_49736);
nor UO_2763 (O_2763,N_49628,N_49502);
nor UO_2764 (O_2764,N_49989,N_49984);
nor UO_2765 (O_2765,N_49811,N_49537);
and UO_2766 (O_2766,N_49799,N_49910);
and UO_2767 (O_2767,N_49669,N_49541);
or UO_2768 (O_2768,N_49877,N_49986);
xnor UO_2769 (O_2769,N_49675,N_49805);
nor UO_2770 (O_2770,N_49543,N_49767);
and UO_2771 (O_2771,N_49796,N_49635);
and UO_2772 (O_2772,N_49997,N_49890);
or UO_2773 (O_2773,N_49880,N_49723);
nand UO_2774 (O_2774,N_49639,N_49920);
nand UO_2775 (O_2775,N_49696,N_49834);
or UO_2776 (O_2776,N_49923,N_49643);
or UO_2777 (O_2777,N_49572,N_49772);
xnor UO_2778 (O_2778,N_49505,N_49561);
or UO_2779 (O_2779,N_49656,N_49862);
nor UO_2780 (O_2780,N_49865,N_49957);
and UO_2781 (O_2781,N_49528,N_49637);
nor UO_2782 (O_2782,N_49611,N_49900);
nand UO_2783 (O_2783,N_49947,N_49848);
and UO_2784 (O_2784,N_49905,N_49853);
nor UO_2785 (O_2785,N_49739,N_49668);
or UO_2786 (O_2786,N_49581,N_49524);
nor UO_2787 (O_2787,N_49898,N_49579);
nand UO_2788 (O_2788,N_49510,N_49650);
xnor UO_2789 (O_2789,N_49586,N_49634);
nand UO_2790 (O_2790,N_49768,N_49884);
nor UO_2791 (O_2791,N_49789,N_49540);
nor UO_2792 (O_2792,N_49883,N_49963);
and UO_2793 (O_2793,N_49887,N_49816);
and UO_2794 (O_2794,N_49742,N_49818);
or UO_2795 (O_2795,N_49853,N_49811);
and UO_2796 (O_2796,N_49948,N_49953);
or UO_2797 (O_2797,N_49759,N_49690);
and UO_2798 (O_2798,N_49857,N_49902);
and UO_2799 (O_2799,N_49715,N_49571);
or UO_2800 (O_2800,N_49652,N_49822);
or UO_2801 (O_2801,N_49543,N_49562);
and UO_2802 (O_2802,N_49724,N_49564);
or UO_2803 (O_2803,N_49617,N_49927);
or UO_2804 (O_2804,N_49759,N_49877);
and UO_2805 (O_2805,N_49934,N_49788);
or UO_2806 (O_2806,N_49959,N_49517);
nor UO_2807 (O_2807,N_49879,N_49996);
or UO_2808 (O_2808,N_49889,N_49622);
and UO_2809 (O_2809,N_49686,N_49878);
or UO_2810 (O_2810,N_49917,N_49875);
nand UO_2811 (O_2811,N_49793,N_49622);
nand UO_2812 (O_2812,N_49682,N_49500);
nor UO_2813 (O_2813,N_49525,N_49792);
and UO_2814 (O_2814,N_49800,N_49909);
xnor UO_2815 (O_2815,N_49558,N_49913);
or UO_2816 (O_2816,N_49546,N_49544);
nor UO_2817 (O_2817,N_49593,N_49515);
and UO_2818 (O_2818,N_49829,N_49739);
and UO_2819 (O_2819,N_49925,N_49593);
or UO_2820 (O_2820,N_49736,N_49868);
nand UO_2821 (O_2821,N_49522,N_49666);
nand UO_2822 (O_2822,N_49809,N_49710);
or UO_2823 (O_2823,N_49605,N_49607);
nand UO_2824 (O_2824,N_49817,N_49736);
nand UO_2825 (O_2825,N_49803,N_49566);
nor UO_2826 (O_2826,N_49579,N_49944);
xor UO_2827 (O_2827,N_49639,N_49897);
xnor UO_2828 (O_2828,N_49856,N_49530);
nand UO_2829 (O_2829,N_49628,N_49876);
and UO_2830 (O_2830,N_49968,N_49589);
or UO_2831 (O_2831,N_49936,N_49678);
or UO_2832 (O_2832,N_49588,N_49592);
and UO_2833 (O_2833,N_49663,N_49513);
nand UO_2834 (O_2834,N_49922,N_49608);
and UO_2835 (O_2835,N_49824,N_49843);
or UO_2836 (O_2836,N_49820,N_49738);
or UO_2837 (O_2837,N_49849,N_49783);
or UO_2838 (O_2838,N_49779,N_49691);
and UO_2839 (O_2839,N_49629,N_49823);
nor UO_2840 (O_2840,N_49820,N_49676);
xnor UO_2841 (O_2841,N_49600,N_49837);
nor UO_2842 (O_2842,N_49890,N_49926);
or UO_2843 (O_2843,N_49700,N_49924);
nand UO_2844 (O_2844,N_49607,N_49622);
and UO_2845 (O_2845,N_49879,N_49950);
nand UO_2846 (O_2846,N_49810,N_49984);
xor UO_2847 (O_2847,N_49801,N_49691);
and UO_2848 (O_2848,N_49627,N_49684);
and UO_2849 (O_2849,N_49846,N_49918);
nand UO_2850 (O_2850,N_49616,N_49620);
or UO_2851 (O_2851,N_49949,N_49758);
or UO_2852 (O_2852,N_49959,N_49510);
and UO_2853 (O_2853,N_49781,N_49905);
xnor UO_2854 (O_2854,N_49600,N_49976);
or UO_2855 (O_2855,N_49580,N_49812);
xor UO_2856 (O_2856,N_49759,N_49646);
xnor UO_2857 (O_2857,N_49818,N_49627);
and UO_2858 (O_2858,N_49733,N_49777);
xnor UO_2859 (O_2859,N_49884,N_49651);
nor UO_2860 (O_2860,N_49920,N_49706);
nand UO_2861 (O_2861,N_49881,N_49626);
nor UO_2862 (O_2862,N_49555,N_49950);
nand UO_2863 (O_2863,N_49906,N_49697);
nand UO_2864 (O_2864,N_49867,N_49720);
and UO_2865 (O_2865,N_49981,N_49519);
nor UO_2866 (O_2866,N_49964,N_49660);
or UO_2867 (O_2867,N_49503,N_49919);
nand UO_2868 (O_2868,N_49931,N_49915);
and UO_2869 (O_2869,N_49880,N_49650);
nor UO_2870 (O_2870,N_49797,N_49692);
or UO_2871 (O_2871,N_49537,N_49797);
nand UO_2872 (O_2872,N_49851,N_49507);
and UO_2873 (O_2873,N_49762,N_49994);
and UO_2874 (O_2874,N_49809,N_49685);
xor UO_2875 (O_2875,N_49677,N_49586);
nand UO_2876 (O_2876,N_49746,N_49553);
nand UO_2877 (O_2877,N_49632,N_49585);
nor UO_2878 (O_2878,N_49924,N_49941);
nand UO_2879 (O_2879,N_49787,N_49639);
or UO_2880 (O_2880,N_49673,N_49900);
nand UO_2881 (O_2881,N_49537,N_49786);
or UO_2882 (O_2882,N_49704,N_49705);
nand UO_2883 (O_2883,N_49734,N_49510);
nand UO_2884 (O_2884,N_49885,N_49508);
nor UO_2885 (O_2885,N_49958,N_49755);
and UO_2886 (O_2886,N_49543,N_49858);
or UO_2887 (O_2887,N_49836,N_49802);
nand UO_2888 (O_2888,N_49753,N_49601);
and UO_2889 (O_2889,N_49530,N_49561);
nor UO_2890 (O_2890,N_49528,N_49710);
and UO_2891 (O_2891,N_49620,N_49897);
or UO_2892 (O_2892,N_49537,N_49854);
nand UO_2893 (O_2893,N_49987,N_49806);
and UO_2894 (O_2894,N_49719,N_49653);
or UO_2895 (O_2895,N_49920,N_49601);
and UO_2896 (O_2896,N_49753,N_49944);
nor UO_2897 (O_2897,N_49690,N_49685);
and UO_2898 (O_2898,N_49509,N_49885);
and UO_2899 (O_2899,N_49657,N_49791);
or UO_2900 (O_2900,N_49853,N_49987);
or UO_2901 (O_2901,N_49758,N_49632);
and UO_2902 (O_2902,N_49617,N_49947);
or UO_2903 (O_2903,N_49636,N_49524);
or UO_2904 (O_2904,N_49712,N_49618);
and UO_2905 (O_2905,N_49856,N_49756);
nor UO_2906 (O_2906,N_49985,N_49702);
xnor UO_2907 (O_2907,N_49670,N_49619);
nor UO_2908 (O_2908,N_49631,N_49790);
nor UO_2909 (O_2909,N_49878,N_49602);
nor UO_2910 (O_2910,N_49739,N_49522);
nand UO_2911 (O_2911,N_49518,N_49842);
and UO_2912 (O_2912,N_49886,N_49622);
and UO_2913 (O_2913,N_49697,N_49591);
nor UO_2914 (O_2914,N_49670,N_49813);
nand UO_2915 (O_2915,N_49607,N_49766);
xnor UO_2916 (O_2916,N_49588,N_49892);
or UO_2917 (O_2917,N_49855,N_49927);
nand UO_2918 (O_2918,N_49977,N_49708);
nor UO_2919 (O_2919,N_49501,N_49939);
and UO_2920 (O_2920,N_49884,N_49609);
nand UO_2921 (O_2921,N_49699,N_49681);
and UO_2922 (O_2922,N_49912,N_49574);
or UO_2923 (O_2923,N_49737,N_49872);
and UO_2924 (O_2924,N_49603,N_49932);
or UO_2925 (O_2925,N_49589,N_49550);
nand UO_2926 (O_2926,N_49768,N_49779);
nor UO_2927 (O_2927,N_49690,N_49886);
or UO_2928 (O_2928,N_49565,N_49612);
or UO_2929 (O_2929,N_49660,N_49667);
or UO_2930 (O_2930,N_49678,N_49874);
xnor UO_2931 (O_2931,N_49770,N_49948);
xnor UO_2932 (O_2932,N_49520,N_49950);
nand UO_2933 (O_2933,N_49753,N_49958);
nand UO_2934 (O_2934,N_49791,N_49985);
nor UO_2935 (O_2935,N_49705,N_49742);
or UO_2936 (O_2936,N_49948,N_49931);
and UO_2937 (O_2937,N_49616,N_49776);
and UO_2938 (O_2938,N_49699,N_49565);
or UO_2939 (O_2939,N_49554,N_49918);
or UO_2940 (O_2940,N_49737,N_49779);
xor UO_2941 (O_2941,N_49937,N_49661);
nor UO_2942 (O_2942,N_49556,N_49922);
or UO_2943 (O_2943,N_49784,N_49518);
nor UO_2944 (O_2944,N_49993,N_49666);
and UO_2945 (O_2945,N_49593,N_49964);
xnor UO_2946 (O_2946,N_49833,N_49952);
or UO_2947 (O_2947,N_49984,N_49945);
nor UO_2948 (O_2948,N_49699,N_49628);
and UO_2949 (O_2949,N_49753,N_49505);
or UO_2950 (O_2950,N_49599,N_49967);
xor UO_2951 (O_2951,N_49922,N_49902);
or UO_2952 (O_2952,N_49667,N_49725);
or UO_2953 (O_2953,N_49900,N_49585);
or UO_2954 (O_2954,N_49759,N_49930);
nor UO_2955 (O_2955,N_49809,N_49800);
or UO_2956 (O_2956,N_49906,N_49819);
nand UO_2957 (O_2957,N_49638,N_49774);
nand UO_2958 (O_2958,N_49987,N_49655);
nor UO_2959 (O_2959,N_49753,N_49834);
or UO_2960 (O_2960,N_49692,N_49998);
or UO_2961 (O_2961,N_49767,N_49751);
and UO_2962 (O_2962,N_49626,N_49644);
nor UO_2963 (O_2963,N_49920,N_49776);
xnor UO_2964 (O_2964,N_49606,N_49616);
or UO_2965 (O_2965,N_49849,N_49576);
nand UO_2966 (O_2966,N_49993,N_49542);
and UO_2967 (O_2967,N_49735,N_49658);
or UO_2968 (O_2968,N_49877,N_49525);
xnor UO_2969 (O_2969,N_49847,N_49715);
and UO_2970 (O_2970,N_49924,N_49851);
or UO_2971 (O_2971,N_49749,N_49709);
or UO_2972 (O_2972,N_49810,N_49690);
or UO_2973 (O_2973,N_49753,N_49524);
and UO_2974 (O_2974,N_49574,N_49965);
or UO_2975 (O_2975,N_49909,N_49569);
or UO_2976 (O_2976,N_49822,N_49578);
nor UO_2977 (O_2977,N_49821,N_49606);
or UO_2978 (O_2978,N_49545,N_49585);
nand UO_2979 (O_2979,N_49528,N_49915);
nand UO_2980 (O_2980,N_49727,N_49654);
and UO_2981 (O_2981,N_49671,N_49600);
nand UO_2982 (O_2982,N_49759,N_49678);
xor UO_2983 (O_2983,N_49808,N_49571);
xnor UO_2984 (O_2984,N_49803,N_49926);
and UO_2985 (O_2985,N_49956,N_49920);
and UO_2986 (O_2986,N_49677,N_49742);
xnor UO_2987 (O_2987,N_49779,N_49746);
nand UO_2988 (O_2988,N_49711,N_49644);
nand UO_2989 (O_2989,N_49610,N_49802);
and UO_2990 (O_2990,N_49843,N_49816);
or UO_2991 (O_2991,N_49881,N_49553);
nor UO_2992 (O_2992,N_49670,N_49575);
or UO_2993 (O_2993,N_49739,N_49774);
nor UO_2994 (O_2994,N_49801,N_49615);
or UO_2995 (O_2995,N_49912,N_49955);
xnor UO_2996 (O_2996,N_49899,N_49700);
and UO_2997 (O_2997,N_49760,N_49870);
nand UO_2998 (O_2998,N_49691,N_49662);
or UO_2999 (O_2999,N_49560,N_49566);
and UO_3000 (O_3000,N_49635,N_49814);
and UO_3001 (O_3001,N_49571,N_49569);
and UO_3002 (O_3002,N_49685,N_49525);
nand UO_3003 (O_3003,N_49592,N_49886);
or UO_3004 (O_3004,N_49595,N_49770);
nand UO_3005 (O_3005,N_49580,N_49959);
nand UO_3006 (O_3006,N_49785,N_49791);
and UO_3007 (O_3007,N_49508,N_49529);
and UO_3008 (O_3008,N_49723,N_49660);
nor UO_3009 (O_3009,N_49692,N_49774);
nor UO_3010 (O_3010,N_49638,N_49658);
nand UO_3011 (O_3011,N_49920,N_49684);
or UO_3012 (O_3012,N_49702,N_49875);
and UO_3013 (O_3013,N_49536,N_49722);
nand UO_3014 (O_3014,N_49533,N_49752);
and UO_3015 (O_3015,N_49875,N_49928);
nand UO_3016 (O_3016,N_49538,N_49698);
nor UO_3017 (O_3017,N_49984,N_49692);
nand UO_3018 (O_3018,N_49813,N_49948);
nor UO_3019 (O_3019,N_49532,N_49796);
nand UO_3020 (O_3020,N_49967,N_49891);
nand UO_3021 (O_3021,N_49658,N_49968);
xor UO_3022 (O_3022,N_49671,N_49540);
nor UO_3023 (O_3023,N_49897,N_49946);
xor UO_3024 (O_3024,N_49867,N_49619);
nand UO_3025 (O_3025,N_49771,N_49703);
and UO_3026 (O_3026,N_49623,N_49800);
and UO_3027 (O_3027,N_49871,N_49521);
and UO_3028 (O_3028,N_49795,N_49682);
nand UO_3029 (O_3029,N_49638,N_49910);
or UO_3030 (O_3030,N_49709,N_49688);
nor UO_3031 (O_3031,N_49737,N_49778);
xnor UO_3032 (O_3032,N_49500,N_49916);
nand UO_3033 (O_3033,N_49513,N_49522);
nand UO_3034 (O_3034,N_49503,N_49667);
and UO_3035 (O_3035,N_49527,N_49622);
nor UO_3036 (O_3036,N_49582,N_49550);
and UO_3037 (O_3037,N_49805,N_49758);
nor UO_3038 (O_3038,N_49580,N_49973);
and UO_3039 (O_3039,N_49869,N_49524);
nor UO_3040 (O_3040,N_49674,N_49576);
or UO_3041 (O_3041,N_49648,N_49663);
and UO_3042 (O_3042,N_49773,N_49863);
or UO_3043 (O_3043,N_49625,N_49714);
and UO_3044 (O_3044,N_49607,N_49970);
nor UO_3045 (O_3045,N_49829,N_49791);
and UO_3046 (O_3046,N_49529,N_49631);
nand UO_3047 (O_3047,N_49982,N_49996);
or UO_3048 (O_3048,N_49659,N_49998);
nand UO_3049 (O_3049,N_49796,N_49540);
xnor UO_3050 (O_3050,N_49986,N_49550);
xnor UO_3051 (O_3051,N_49589,N_49623);
or UO_3052 (O_3052,N_49904,N_49574);
nand UO_3053 (O_3053,N_49665,N_49551);
or UO_3054 (O_3054,N_49954,N_49958);
nand UO_3055 (O_3055,N_49523,N_49985);
and UO_3056 (O_3056,N_49535,N_49913);
or UO_3057 (O_3057,N_49572,N_49660);
nand UO_3058 (O_3058,N_49778,N_49765);
or UO_3059 (O_3059,N_49703,N_49925);
nor UO_3060 (O_3060,N_49832,N_49680);
nand UO_3061 (O_3061,N_49781,N_49557);
and UO_3062 (O_3062,N_49724,N_49536);
and UO_3063 (O_3063,N_49927,N_49777);
nand UO_3064 (O_3064,N_49562,N_49970);
and UO_3065 (O_3065,N_49891,N_49951);
nand UO_3066 (O_3066,N_49590,N_49956);
or UO_3067 (O_3067,N_49969,N_49513);
nand UO_3068 (O_3068,N_49526,N_49513);
nand UO_3069 (O_3069,N_49671,N_49793);
nor UO_3070 (O_3070,N_49726,N_49924);
xnor UO_3071 (O_3071,N_49666,N_49754);
nor UO_3072 (O_3072,N_49836,N_49909);
or UO_3073 (O_3073,N_49958,N_49842);
or UO_3074 (O_3074,N_49738,N_49538);
and UO_3075 (O_3075,N_49803,N_49551);
and UO_3076 (O_3076,N_49665,N_49519);
nor UO_3077 (O_3077,N_49729,N_49758);
or UO_3078 (O_3078,N_49847,N_49693);
xor UO_3079 (O_3079,N_49685,N_49981);
nand UO_3080 (O_3080,N_49689,N_49929);
and UO_3081 (O_3081,N_49724,N_49991);
or UO_3082 (O_3082,N_49761,N_49604);
or UO_3083 (O_3083,N_49514,N_49793);
or UO_3084 (O_3084,N_49976,N_49632);
nor UO_3085 (O_3085,N_49869,N_49549);
and UO_3086 (O_3086,N_49710,N_49758);
nor UO_3087 (O_3087,N_49919,N_49595);
nor UO_3088 (O_3088,N_49543,N_49941);
or UO_3089 (O_3089,N_49830,N_49643);
and UO_3090 (O_3090,N_49608,N_49839);
xor UO_3091 (O_3091,N_49776,N_49768);
nor UO_3092 (O_3092,N_49796,N_49678);
or UO_3093 (O_3093,N_49537,N_49858);
nand UO_3094 (O_3094,N_49752,N_49513);
nand UO_3095 (O_3095,N_49564,N_49891);
nand UO_3096 (O_3096,N_49894,N_49521);
nor UO_3097 (O_3097,N_49989,N_49653);
nor UO_3098 (O_3098,N_49699,N_49720);
and UO_3099 (O_3099,N_49613,N_49827);
xnor UO_3100 (O_3100,N_49778,N_49652);
nand UO_3101 (O_3101,N_49910,N_49611);
nor UO_3102 (O_3102,N_49896,N_49928);
nand UO_3103 (O_3103,N_49815,N_49836);
xnor UO_3104 (O_3104,N_49624,N_49794);
nand UO_3105 (O_3105,N_49719,N_49890);
nor UO_3106 (O_3106,N_49968,N_49894);
nor UO_3107 (O_3107,N_49938,N_49883);
nand UO_3108 (O_3108,N_49576,N_49511);
and UO_3109 (O_3109,N_49963,N_49906);
nor UO_3110 (O_3110,N_49640,N_49608);
nor UO_3111 (O_3111,N_49755,N_49930);
and UO_3112 (O_3112,N_49670,N_49597);
nand UO_3113 (O_3113,N_49746,N_49642);
and UO_3114 (O_3114,N_49711,N_49654);
nand UO_3115 (O_3115,N_49602,N_49840);
and UO_3116 (O_3116,N_49522,N_49717);
xor UO_3117 (O_3117,N_49673,N_49969);
and UO_3118 (O_3118,N_49685,N_49920);
nor UO_3119 (O_3119,N_49999,N_49658);
and UO_3120 (O_3120,N_49968,N_49569);
nand UO_3121 (O_3121,N_49940,N_49979);
nor UO_3122 (O_3122,N_49617,N_49871);
nand UO_3123 (O_3123,N_49759,N_49922);
or UO_3124 (O_3124,N_49717,N_49554);
or UO_3125 (O_3125,N_49789,N_49787);
or UO_3126 (O_3126,N_49503,N_49989);
nand UO_3127 (O_3127,N_49933,N_49622);
or UO_3128 (O_3128,N_49601,N_49896);
nor UO_3129 (O_3129,N_49540,N_49936);
and UO_3130 (O_3130,N_49625,N_49684);
nand UO_3131 (O_3131,N_49592,N_49758);
or UO_3132 (O_3132,N_49884,N_49523);
nor UO_3133 (O_3133,N_49545,N_49668);
nor UO_3134 (O_3134,N_49845,N_49610);
or UO_3135 (O_3135,N_49533,N_49696);
or UO_3136 (O_3136,N_49554,N_49858);
or UO_3137 (O_3137,N_49567,N_49792);
and UO_3138 (O_3138,N_49597,N_49960);
or UO_3139 (O_3139,N_49787,N_49827);
nor UO_3140 (O_3140,N_49803,N_49598);
and UO_3141 (O_3141,N_49869,N_49905);
and UO_3142 (O_3142,N_49745,N_49946);
nand UO_3143 (O_3143,N_49857,N_49796);
nand UO_3144 (O_3144,N_49978,N_49853);
xor UO_3145 (O_3145,N_49958,N_49704);
nor UO_3146 (O_3146,N_49614,N_49884);
nand UO_3147 (O_3147,N_49659,N_49950);
or UO_3148 (O_3148,N_49874,N_49514);
nor UO_3149 (O_3149,N_49884,N_49866);
and UO_3150 (O_3150,N_49799,N_49940);
xor UO_3151 (O_3151,N_49529,N_49953);
nand UO_3152 (O_3152,N_49984,N_49627);
nand UO_3153 (O_3153,N_49957,N_49994);
and UO_3154 (O_3154,N_49890,N_49991);
nand UO_3155 (O_3155,N_49970,N_49724);
nor UO_3156 (O_3156,N_49560,N_49900);
xnor UO_3157 (O_3157,N_49501,N_49587);
and UO_3158 (O_3158,N_49706,N_49574);
nand UO_3159 (O_3159,N_49588,N_49584);
nand UO_3160 (O_3160,N_49876,N_49566);
and UO_3161 (O_3161,N_49781,N_49675);
and UO_3162 (O_3162,N_49795,N_49778);
nand UO_3163 (O_3163,N_49970,N_49532);
nand UO_3164 (O_3164,N_49668,N_49627);
and UO_3165 (O_3165,N_49796,N_49979);
or UO_3166 (O_3166,N_49584,N_49916);
and UO_3167 (O_3167,N_49729,N_49680);
nand UO_3168 (O_3168,N_49749,N_49592);
xnor UO_3169 (O_3169,N_49531,N_49569);
and UO_3170 (O_3170,N_49917,N_49806);
and UO_3171 (O_3171,N_49991,N_49830);
nor UO_3172 (O_3172,N_49705,N_49683);
and UO_3173 (O_3173,N_49523,N_49937);
or UO_3174 (O_3174,N_49846,N_49739);
nand UO_3175 (O_3175,N_49822,N_49829);
xnor UO_3176 (O_3176,N_49821,N_49557);
nor UO_3177 (O_3177,N_49553,N_49688);
or UO_3178 (O_3178,N_49739,N_49650);
or UO_3179 (O_3179,N_49727,N_49638);
nor UO_3180 (O_3180,N_49738,N_49535);
or UO_3181 (O_3181,N_49623,N_49848);
and UO_3182 (O_3182,N_49776,N_49514);
or UO_3183 (O_3183,N_49535,N_49558);
nor UO_3184 (O_3184,N_49730,N_49586);
or UO_3185 (O_3185,N_49696,N_49664);
nor UO_3186 (O_3186,N_49528,N_49720);
nor UO_3187 (O_3187,N_49523,N_49649);
nand UO_3188 (O_3188,N_49764,N_49734);
nand UO_3189 (O_3189,N_49828,N_49512);
and UO_3190 (O_3190,N_49976,N_49680);
nand UO_3191 (O_3191,N_49574,N_49723);
nand UO_3192 (O_3192,N_49622,N_49959);
or UO_3193 (O_3193,N_49911,N_49680);
nor UO_3194 (O_3194,N_49770,N_49847);
and UO_3195 (O_3195,N_49826,N_49507);
nand UO_3196 (O_3196,N_49831,N_49807);
nand UO_3197 (O_3197,N_49964,N_49672);
xor UO_3198 (O_3198,N_49774,N_49555);
or UO_3199 (O_3199,N_49671,N_49505);
nor UO_3200 (O_3200,N_49574,N_49735);
nor UO_3201 (O_3201,N_49602,N_49586);
and UO_3202 (O_3202,N_49864,N_49849);
nand UO_3203 (O_3203,N_49507,N_49779);
and UO_3204 (O_3204,N_49776,N_49661);
xnor UO_3205 (O_3205,N_49908,N_49586);
or UO_3206 (O_3206,N_49939,N_49674);
xor UO_3207 (O_3207,N_49870,N_49582);
nor UO_3208 (O_3208,N_49691,N_49672);
or UO_3209 (O_3209,N_49779,N_49918);
nand UO_3210 (O_3210,N_49612,N_49775);
and UO_3211 (O_3211,N_49823,N_49592);
nand UO_3212 (O_3212,N_49823,N_49737);
nand UO_3213 (O_3213,N_49863,N_49916);
and UO_3214 (O_3214,N_49896,N_49759);
or UO_3215 (O_3215,N_49911,N_49628);
xnor UO_3216 (O_3216,N_49553,N_49544);
nor UO_3217 (O_3217,N_49864,N_49553);
nand UO_3218 (O_3218,N_49517,N_49876);
nor UO_3219 (O_3219,N_49557,N_49780);
or UO_3220 (O_3220,N_49692,N_49889);
nor UO_3221 (O_3221,N_49694,N_49628);
and UO_3222 (O_3222,N_49635,N_49627);
nor UO_3223 (O_3223,N_49678,N_49669);
nand UO_3224 (O_3224,N_49779,N_49628);
nand UO_3225 (O_3225,N_49910,N_49959);
xor UO_3226 (O_3226,N_49537,N_49831);
xor UO_3227 (O_3227,N_49852,N_49928);
or UO_3228 (O_3228,N_49898,N_49806);
or UO_3229 (O_3229,N_49819,N_49807);
nor UO_3230 (O_3230,N_49946,N_49875);
nor UO_3231 (O_3231,N_49793,N_49644);
and UO_3232 (O_3232,N_49736,N_49883);
and UO_3233 (O_3233,N_49609,N_49691);
and UO_3234 (O_3234,N_49563,N_49931);
and UO_3235 (O_3235,N_49578,N_49616);
xnor UO_3236 (O_3236,N_49922,N_49929);
nor UO_3237 (O_3237,N_49990,N_49853);
or UO_3238 (O_3238,N_49992,N_49929);
nor UO_3239 (O_3239,N_49606,N_49565);
and UO_3240 (O_3240,N_49794,N_49593);
or UO_3241 (O_3241,N_49799,N_49948);
xor UO_3242 (O_3242,N_49796,N_49563);
nand UO_3243 (O_3243,N_49657,N_49752);
or UO_3244 (O_3244,N_49527,N_49729);
nand UO_3245 (O_3245,N_49508,N_49852);
and UO_3246 (O_3246,N_49588,N_49711);
nand UO_3247 (O_3247,N_49531,N_49821);
nand UO_3248 (O_3248,N_49701,N_49643);
or UO_3249 (O_3249,N_49654,N_49963);
or UO_3250 (O_3250,N_49687,N_49539);
nand UO_3251 (O_3251,N_49966,N_49954);
xnor UO_3252 (O_3252,N_49592,N_49787);
nor UO_3253 (O_3253,N_49956,N_49861);
nor UO_3254 (O_3254,N_49718,N_49741);
nor UO_3255 (O_3255,N_49953,N_49873);
nand UO_3256 (O_3256,N_49627,N_49592);
nor UO_3257 (O_3257,N_49996,N_49970);
nand UO_3258 (O_3258,N_49759,N_49924);
nor UO_3259 (O_3259,N_49741,N_49938);
or UO_3260 (O_3260,N_49723,N_49737);
xor UO_3261 (O_3261,N_49666,N_49644);
nand UO_3262 (O_3262,N_49739,N_49710);
xnor UO_3263 (O_3263,N_49656,N_49969);
xor UO_3264 (O_3264,N_49821,N_49712);
or UO_3265 (O_3265,N_49893,N_49715);
nor UO_3266 (O_3266,N_49788,N_49822);
and UO_3267 (O_3267,N_49930,N_49925);
xnor UO_3268 (O_3268,N_49756,N_49821);
nor UO_3269 (O_3269,N_49709,N_49739);
nor UO_3270 (O_3270,N_49813,N_49829);
nor UO_3271 (O_3271,N_49662,N_49721);
and UO_3272 (O_3272,N_49541,N_49511);
nor UO_3273 (O_3273,N_49991,N_49968);
and UO_3274 (O_3274,N_49778,N_49685);
and UO_3275 (O_3275,N_49971,N_49561);
and UO_3276 (O_3276,N_49704,N_49718);
nand UO_3277 (O_3277,N_49862,N_49556);
nor UO_3278 (O_3278,N_49517,N_49897);
nor UO_3279 (O_3279,N_49621,N_49773);
nor UO_3280 (O_3280,N_49888,N_49642);
xnor UO_3281 (O_3281,N_49988,N_49676);
nand UO_3282 (O_3282,N_49634,N_49691);
and UO_3283 (O_3283,N_49822,N_49513);
or UO_3284 (O_3284,N_49784,N_49544);
nand UO_3285 (O_3285,N_49508,N_49748);
and UO_3286 (O_3286,N_49540,N_49975);
and UO_3287 (O_3287,N_49697,N_49897);
nand UO_3288 (O_3288,N_49615,N_49898);
and UO_3289 (O_3289,N_49902,N_49948);
nor UO_3290 (O_3290,N_49959,N_49720);
or UO_3291 (O_3291,N_49990,N_49744);
xor UO_3292 (O_3292,N_49602,N_49911);
xor UO_3293 (O_3293,N_49895,N_49878);
and UO_3294 (O_3294,N_49764,N_49594);
nand UO_3295 (O_3295,N_49609,N_49836);
nand UO_3296 (O_3296,N_49947,N_49888);
or UO_3297 (O_3297,N_49937,N_49880);
or UO_3298 (O_3298,N_49974,N_49612);
or UO_3299 (O_3299,N_49960,N_49645);
nor UO_3300 (O_3300,N_49846,N_49823);
and UO_3301 (O_3301,N_49960,N_49810);
or UO_3302 (O_3302,N_49782,N_49886);
nor UO_3303 (O_3303,N_49805,N_49661);
xor UO_3304 (O_3304,N_49930,N_49860);
nor UO_3305 (O_3305,N_49560,N_49570);
xor UO_3306 (O_3306,N_49699,N_49652);
nor UO_3307 (O_3307,N_49657,N_49937);
or UO_3308 (O_3308,N_49636,N_49852);
nor UO_3309 (O_3309,N_49958,N_49864);
and UO_3310 (O_3310,N_49913,N_49649);
and UO_3311 (O_3311,N_49683,N_49776);
and UO_3312 (O_3312,N_49941,N_49894);
or UO_3313 (O_3313,N_49675,N_49618);
nand UO_3314 (O_3314,N_49622,N_49673);
and UO_3315 (O_3315,N_49576,N_49979);
xnor UO_3316 (O_3316,N_49952,N_49500);
nor UO_3317 (O_3317,N_49739,N_49945);
xor UO_3318 (O_3318,N_49962,N_49975);
xor UO_3319 (O_3319,N_49671,N_49923);
and UO_3320 (O_3320,N_49988,N_49820);
or UO_3321 (O_3321,N_49705,N_49528);
nand UO_3322 (O_3322,N_49924,N_49527);
nor UO_3323 (O_3323,N_49510,N_49643);
or UO_3324 (O_3324,N_49725,N_49656);
nand UO_3325 (O_3325,N_49707,N_49900);
xnor UO_3326 (O_3326,N_49900,N_49816);
nand UO_3327 (O_3327,N_49749,N_49783);
nor UO_3328 (O_3328,N_49787,N_49909);
nand UO_3329 (O_3329,N_49518,N_49667);
or UO_3330 (O_3330,N_49943,N_49993);
nor UO_3331 (O_3331,N_49636,N_49725);
and UO_3332 (O_3332,N_49674,N_49937);
nand UO_3333 (O_3333,N_49600,N_49983);
nor UO_3334 (O_3334,N_49621,N_49503);
nor UO_3335 (O_3335,N_49908,N_49868);
or UO_3336 (O_3336,N_49633,N_49642);
and UO_3337 (O_3337,N_49915,N_49942);
or UO_3338 (O_3338,N_49863,N_49588);
xnor UO_3339 (O_3339,N_49972,N_49708);
or UO_3340 (O_3340,N_49814,N_49901);
nand UO_3341 (O_3341,N_49909,N_49703);
xor UO_3342 (O_3342,N_49959,N_49575);
and UO_3343 (O_3343,N_49994,N_49861);
nor UO_3344 (O_3344,N_49589,N_49781);
nor UO_3345 (O_3345,N_49775,N_49505);
nor UO_3346 (O_3346,N_49776,N_49559);
and UO_3347 (O_3347,N_49809,N_49877);
xnor UO_3348 (O_3348,N_49680,N_49782);
and UO_3349 (O_3349,N_49520,N_49609);
xor UO_3350 (O_3350,N_49590,N_49904);
or UO_3351 (O_3351,N_49506,N_49988);
nor UO_3352 (O_3352,N_49832,N_49682);
nand UO_3353 (O_3353,N_49559,N_49832);
or UO_3354 (O_3354,N_49983,N_49909);
and UO_3355 (O_3355,N_49701,N_49758);
or UO_3356 (O_3356,N_49869,N_49965);
and UO_3357 (O_3357,N_49651,N_49631);
or UO_3358 (O_3358,N_49763,N_49783);
nor UO_3359 (O_3359,N_49724,N_49528);
xnor UO_3360 (O_3360,N_49921,N_49844);
nand UO_3361 (O_3361,N_49981,N_49707);
nand UO_3362 (O_3362,N_49551,N_49943);
nor UO_3363 (O_3363,N_49882,N_49537);
or UO_3364 (O_3364,N_49937,N_49623);
or UO_3365 (O_3365,N_49646,N_49827);
and UO_3366 (O_3366,N_49642,N_49686);
nor UO_3367 (O_3367,N_49530,N_49827);
nand UO_3368 (O_3368,N_49886,N_49978);
or UO_3369 (O_3369,N_49990,N_49524);
and UO_3370 (O_3370,N_49727,N_49548);
xnor UO_3371 (O_3371,N_49765,N_49976);
or UO_3372 (O_3372,N_49779,N_49524);
nand UO_3373 (O_3373,N_49860,N_49518);
nand UO_3374 (O_3374,N_49768,N_49855);
xor UO_3375 (O_3375,N_49911,N_49702);
nor UO_3376 (O_3376,N_49750,N_49934);
nand UO_3377 (O_3377,N_49746,N_49737);
or UO_3378 (O_3378,N_49609,N_49811);
nand UO_3379 (O_3379,N_49502,N_49963);
and UO_3380 (O_3380,N_49521,N_49918);
nor UO_3381 (O_3381,N_49855,N_49973);
nand UO_3382 (O_3382,N_49883,N_49623);
nand UO_3383 (O_3383,N_49610,N_49531);
nor UO_3384 (O_3384,N_49615,N_49767);
xnor UO_3385 (O_3385,N_49519,N_49524);
nand UO_3386 (O_3386,N_49679,N_49941);
and UO_3387 (O_3387,N_49649,N_49706);
and UO_3388 (O_3388,N_49930,N_49767);
and UO_3389 (O_3389,N_49990,N_49686);
or UO_3390 (O_3390,N_49723,N_49779);
nand UO_3391 (O_3391,N_49714,N_49665);
nor UO_3392 (O_3392,N_49566,N_49906);
or UO_3393 (O_3393,N_49593,N_49817);
and UO_3394 (O_3394,N_49724,N_49762);
and UO_3395 (O_3395,N_49891,N_49590);
and UO_3396 (O_3396,N_49920,N_49832);
nor UO_3397 (O_3397,N_49925,N_49523);
nand UO_3398 (O_3398,N_49694,N_49560);
nor UO_3399 (O_3399,N_49916,N_49726);
and UO_3400 (O_3400,N_49644,N_49715);
nor UO_3401 (O_3401,N_49661,N_49645);
nor UO_3402 (O_3402,N_49805,N_49622);
or UO_3403 (O_3403,N_49703,N_49701);
nor UO_3404 (O_3404,N_49661,N_49500);
nor UO_3405 (O_3405,N_49632,N_49789);
nor UO_3406 (O_3406,N_49553,N_49630);
nand UO_3407 (O_3407,N_49750,N_49909);
nand UO_3408 (O_3408,N_49509,N_49623);
nand UO_3409 (O_3409,N_49778,N_49873);
nand UO_3410 (O_3410,N_49739,N_49911);
nor UO_3411 (O_3411,N_49708,N_49536);
nand UO_3412 (O_3412,N_49745,N_49948);
nor UO_3413 (O_3413,N_49828,N_49707);
nand UO_3414 (O_3414,N_49761,N_49686);
nand UO_3415 (O_3415,N_49517,N_49873);
nand UO_3416 (O_3416,N_49627,N_49665);
nand UO_3417 (O_3417,N_49867,N_49715);
and UO_3418 (O_3418,N_49596,N_49661);
and UO_3419 (O_3419,N_49701,N_49914);
and UO_3420 (O_3420,N_49874,N_49940);
and UO_3421 (O_3421,N_49515,N_49652);
and UO_3422 (O_3422,N_49512,N_49801);
nand UO_3423 (O_3423,N_49988,N_49830);
nor UO_3424 (O_3424,N_49550,N_49673);
nor UO_3425 (O_3425,N_49764,N_49977);
nand UO_3426 (O_3426,N_49744,N_49697);
nor UO_3427 (O_3427,N_49804,N_49538);
nand UO_3428 (O_3428,N_49786,N_49808);
and UO_3429 (O_3429,N_49862,N_49712);
and UO_3430 (O_3430,N_49925,N_49807);
or UO_3431 (O_3431,N_49950,N_49534);
or UO_3432 (O_3432,N_49749,N_49823);
or UO_3433 (O_3433,N_49816,N_49864);
nor UO_3434 (O_3434,N_49526,N_49786);
nand UO_3435 (O_3435,N_49701,N_49782);
nand UO_3436 (O_3436,N_49956,N_49683);
or UO_3437 (O_3437,N_49779,N_49634);
nand UO_3438 (O_3438,N_49627,N_49964);
or UO_3439 (O_3439,N_49901,N_49983);
nor UO_3440 (O_3440,N_49963,N_49981);
or UO_3441 (O_3441,N_49961,N_49901);
nor UO_3442 (O_3442,N_49763,N_49752);
and UO_3443 (O_3443,N_49721,N_49853);
and UO_3444 (O_3444,N_49713,N_49722);
xor UO_3445 (O_3445,N_49700,N_49792);
nor UO_3446 (O_3446,N_49565,N_49879);
or UO_3447 (O_3447,N_49573,N_49520);
or UO_3448 (O_3448,N_49533,N_49792);
or UO_3449 (O_3449,N_49644,N_49628);
nand UO_3450 (O_3450,N_49761,N_49541);
and UO_3451 (O_3451,N_49529,N_49750);
and UO_3452 (O_3452,N_49689,N_49524);
and UO_3453 (O_3453,N_49849,N_49878);
xor UO_3454 (O_3454,N_49558,N_49609);
nor UO_3455 (O_3455,N_49948,N_49774);
or UO_3456 (O_3456,N_49757,N_49624);
nor UO_3457 (O_3457,N_49557,N_49974);
xnor UO_3458 (O_3458,N_49978,N_49882);
or UO_3459 (O_3459,N_49916,N_49833);
or UO_3460 (O_3460,N_49601,N_49993);
nand UO_3461 (O_3461,N_49736,N_49922);
nand UO_3462 (O_3462,N_49619,N_49552);
nand UO_3463 (O_3463,N_49677,N_49960);
nand UO_3464 (O_3464,N_49534,N_49981);
nand UO_3465 (O_3465,N_49879,N_49513);
and UO_3466 (O_3466,N_49863,N_49855);
and UO_3467 (O_3467,N_49523,N_49644);
nand UO_3468 (O_3468,N_49818,N_49654);
nor UO_3469 (O_3469,N_49695,N_49756);
and UO_3470 (O_3470,N_49811,N_49936);
or UO_3471 (O_3471,N_49822,N_49906);
and UO_3472 (O_3472,N_49804,N_49812);
nand UO_3473 (O_3473,N_49854,N_49871);
nor UO_3474 (O_3474,N_49894,N_49858);
nand UO_3475 (O_3475,N_49992,N_49766);
nand UO_3476 (O_3476,N_49674,N_49973);
and UO_3477 (O_3477,N_49560,N_49547);
nor UO_3478 (O_3478,N_49851,N_49889);
or UO_3479 (O_3479,N_49795,N_49714);
nand UO_3480 (O_3480,N_49645,N_49733);
and UO_3481 (O_3481,N_49810,N_49761);
nor UO_3482 (O_3482,N_49856,N_49697);
and UO_3483 (O_3483,N_49575,N_49897);
and UO_3484 (O_3484,N_49755,N_49706);
and UO_3485 (O_3485,N_49580,N_49526);
or UO_3486 (O_3486,N_49636,N_49616);
nor UO_3487 (O_3487,N_49769,N_49790);
xnor UO_3488 (O_3488,N_49539,N_49979);
or UO_3489 (O_3489,N_49825,N_49720);
nor UO_3490 (O_3490,N_49986,N_49891);
xor UO_3491 (O_3491,N_49951,N_49770);
nand UO_3492 (O_3492,N_49965,N_49669);
nor UO_3493 (O_3493,N_49722,N_49883);
nand UO_3494 (O_3494,N_49661,N_49994);
xnor UO_3495 (O_3495,N_49554,N_49817);
nor UO_3496 (O_3496,N_49792,N_49917);
or UO_3497 (O_3497,N_49955,N_49519);
nor UO_3498 (O_3498,N_49515,N_49915);
or UO_3499 (O_3499,N_49754,N_49566);
or UO_3500 (O_3500,N_49595,N_49900);
and UO_3501 (O_3501,N_49740,N_49678);
or UO_3502 (O_3502,N_49935,N_49919);
nor UO_3503 (O_3503,N_49520,N_49553);
nor UO_3504 (O_3504,N_49531,N_49712);
and UO_3505 (O_3505,N_49744,N_49812);
and UO_3506 (O_3506,N_49615,N_49701);
or UO_3507 (O_3507,N_49527,N_49739);
or UO_3508 (O_3508,N_49538,N_49653);
or UO_3509 (O_3509,N_49665,N_49921);
nor UO_3510 (O_3510,N_49895,N_49871);
or UO_3511 (O_3511,N_49724,N_49968);
xor UO_3512 (O_3512,N_49930,N_49885);
nor UO_3513 (O_3513,N_49653,N_49561);
nor UO_3514 (O_3514,N_49838,N_49539);
or UO_3515 (O_3515,N_49566,N_49896);
nor UO_3516 (O_3516,N_49634,N_49511);
and UO_3517 (O_3517,N_49574,N_49627);
or UO_3518 (O_3518,N_49567,N_49632);
or UO_3519 (O_3519,N_49769,N_49772);
and UO_3520 (O_3520,N_49563,N_49587);
nand UO_3521 (O_3521,N_49657,N_49708);
nand UO_3522 (O_3522,N_49608,N_49642);
or UO_3523 (O_3523,N_49588,N_49786);
nor UO_3524 (O_3524,N_49670,N_49702);
or UO_3525 (O_3525,N_49729,N_49613);
and UO_3526 (O_3526,N_49584,N_49555);
or UO_3527 (O_3527,N_49527,N_49621);
nand UO_3528 (O_3528,N_49686,N_49548);
or UO_3529 (O_3529,N_49832,N_49965);
or UO_3530 (O_3530,N_49718,N_49869);
or UO_3531 (O_3531,N_49658,N_49832);
nor UO_3532 (O_3532,N_49751,N_49527);
or UO_3533 (O_3533,N_49500,N_49754);
or UO_3534 (O_3534,N_49951,N_49505);
and UO_3535 (O_3535,N_49761,N_49504);
and UO_3536 (O_3536,N_49840,N_49954);
xor UO_3537 (O_3537,N_49671,N_49544);
and UO_3538 (O_3538,N_49758,N_49596);
or UO_3539 (O_3539,N_49829,N_49569);
and UO_3540 (O_3540,N_49988,N_49790);
or UO_3541 (O_3541,N_49577,N_49757);
or UO_3542 (O_3542,N_49904,N_49739);
and UO_3543 (O_3543,N_49727,N_49963);
xnor UO_3544 (O_3544,N_49728,N_49749);
nor UO_3545 (O_3545,N_49621,N_49828);
and UO_3546 (O_3546,N_49538,N_49557);
nand UO_3547 (O_3547,N_49717,N_49954);
nand UO_3548 (O_3548,N_49590,N_49735);
and UO_3549 (O_3549,N_49577,N_49668);
xor UO_3550 (O_3550,N_49976,N_49856);
nand UO_3551 (O_3551,N_49799,N_49557);
and UO_3552 (O_3552,N_49671,N_49709);
nor UO_3553 (O_3553,N_49521,N_49787);
or UO_3554 (O_3554,N_49605,N_49971);
and UO_3555 (O_3555,N_49858,N_49755);
nand UO_3556 (O_3556,N_49818,N_49890);
nand UO_3557 (O_3557,N_49664,N_49937);
nor UO_3558 (O_3558,N_49894,N_49909);
and UO_3559 (O_3559,N_49575,N_49898);
nor UO_3560 (O_3560,N_49708,N_49682);
nor UO_3561 (O_3561,N_49916,N_49727);
nand UO_3562 (O_3562,N_49774,N_49666);
nand UO_3563 (O_3563,N_49998,N_49939);
nor UO_3564 (O_3564,N_49944,N_49843);
nand UO_3565 (O_3565,N_49809,N_49869);
nor UO_3566 (O_3566,N_49742,N_49899);
and UO_3567 (O_3567,N_49968,N_49664);
nor UO_3568 (O_3568,N_49692,N_49638);
and UO_3569 (O_3569,N_49606,N_49597);
and UO_3570 (O_3570,N_49949,N_49868);
xnor UO_3571 (O_3571,N_49743,N_49958);
nor UO_3572 (O_3572,N_49998,N_49507);
nor UO_3573 (O_3573,N_49790,N_49656);
nor UO_3574 (O_3574,N_49730,N_49784);
or UO_3575 (O_3575,N_49654,N_49999);
and UO_3576 (O_3576,N_49950,N_49583);
and UO_3577 (O_3577,N_49847,N_49979);
xnor UO_3578 (O_3578,N_49966,N_49685);
nand UO_3579 (O_3579,N_49599,N_49547);
nor UO_3580 (O_3580,N_49872,N_49946);
nand UO_3581 (O_3581,N_49765,N_49911);
and UO_3582 (O_3582,N_49646,N_49905);
nor UO_3583 (O_3583,N_49503,N_49857);
or UO_3584 (O_3584,N_49526,N_49966);
and UO_3585 (O_3585,N_49762,N_49968);
and UO_3586 (O_3586,N_49968,N_49579);
nor UO_3587 (O_3587,N_49958,N_49642);
nor UO_3588 (O_3588,N_49517,N_49704);
nand UO_3589 (O_3589,N_49849,N_49886);
nor UO_3590 (O_3590,N_49883,N_49856);
nand UO_3591 (O_3591,N_49555,N_49561);
or UO_3592 (O_3592,N_49639,N_49980);
or UO_3593 (O_3593,N_49669,N_49571);
or UO_3594 (O_3594,N_49586,N_49870);
or UO_3595 (O_3595,N_49997,N_49789);
nor UO_3596 (O_3596,N_49974,N_49702);
or UO_3597 (O_3597,N_49618,N_49532);
or UO_3598 (O_3598,N_49707,N_49691);
nand UO_3599 (O_3599,N_49819,N_49828);
xnor UO_3600 (O_3600,N_49907,N_49893);
xnor UO_3601 (O_3601,N_49976,N_49786);
nand UO_3602 (O_3602,N_49629,N_49844);
or UO_3603 (O_3603,N_49827,N_49981);
xor UO_3604 (O_3604,N_49896,N_49547);
or UO_3605 (O_3605,N_49589,N_49937);
or UO_3606 (O_3606,N_49735,N_49779);
and UO_3607 (O_3607,N_49586,N_49825);
xnor UO_3608 (O_3608,N_49733,N_49824);
xnor UO_3609 (O_3609,N_49883,N_49780);
nor UO_3610 (O_3610,N_49775,N_49543);
nand UO_3611 (O_3611,N_49609,N_49958);
nand UO_3612 (O_3612,N_49925,N_49559);
nor UO_3613 (O_3613,N_49704,N_49741);
and UO_3614 (O_3614,N_49656,N_49632);
xor UO_3615 (O_3615,N_49763,N_49616);
and UO_3616 (O_3616,N_49672,N_49877);
nand UO_3617 (O_3617,N_49770,N_49517);
xnor UO_3618 (O_3618,N_49647,N_49798);
and UO_3619 (O_3619,N_49506,N_49578);
and UO_3620 (O_3620,N_49504,N_49981);
and UO_3621 (O_3621,N_49753,N_49769);
and UO_3622 (O_3622,N_49982,N_49633);
and UO_3623 (O_3623,N_49733,N_49647);
or UO_3624 (O_3624,N_49924,N_49703);
nor UO_3625 (O_3625,N_49849,N_49711);
or UO_3626 (O_3626,N_49715,N_49565);
nand UO_3627 (O_3627,N_49685,N_49864);
nor UO_3628 (O_3628,N_49831,N_49993);
and UO_3629 (O_3629,N_49920,N_49799);
nand UO_3630 (O_3630,N_49558,N_49627);
nand UO_3631 (O_3631,N_49609,N_49605);
nor UO_3632 (O_3632,N_49614,N_49791);
xnor UO_3633 (O_3633,N_49880,N_49600);
or UO_3634 (O_3634,N_49937,N_49784);
xnor UO_3635 (O_3635,N_49626,N_49543);
nor UO_3636 (O_3636,N_49852,N_49723);
nand UO_3637 (O_3637,N_49657,N_49509);
or UO_3638 (O_3638,N_49722,N_49638);
nor UO_3639 (O_3639,N_49541,N_49843);
and UO_3640 (O_3640,N_49917,N_49940);
nor UO_3641 (O_3641,N_49969,N_49681);
nor UO_3642 (O_3642,N_49715,N_49848);
or UO_3643 (O_3643,N_49500,N_49586);
and UO_3644 (O_3644,N_49949,N_49772);
or UO_3645 (O_3645,N_49863,N_49500);
and UO_3646 (O_3646,N_49538,N_49618);
or UO_3647 (O_3647,N_49752,N_49603);
and UO_3648 (O_3648,N_49811,N_49747);
xor UO_3649 (O_3649,N_49533,N_49539);
and UO_3650 (O_3650,N_49644,N_49911);
and UO_3651 (O_3651,N_49835,N_49855);
and UO_3652 (O_3652,N_49936,N_49826);
or UO_3653 (O_3653,N_49724,N_49623);
or UO_3654 (O_3654,N_49770,N_49994);
nor UO_3655 (O_3655,N_49597,N_49641);
nor UO_3656 (O_3656,N_49783,N_49988);
or UO_3657 (O_3657,N_49757,N_49890);
nor UO_3658 (O_3658,N_49951,N_49726);
nand UO_3659 (O_3659,N_49998,N_49895);
nor UO_3660 (O_3660,N_49578,N_49990);
or UO_3661 (O_3661,N_49969,N_49892);
nand UO_3662 (O_3662,N_49890,N_49771);
or UO_3663 (O_3663,N_49751,N_49509);
xor UO_3664 (O_3664,N_49640,N_49939);
xnor UO_3665 (O_3665,N_49811,N_49997);
nor UO_3666 (O_3666,N_49531,N_49688);
and UO_3667 (O_3667,N_49870,N_49958);
or UO_3668 (O_3668,N_49843,N_49737);
or UO_3669 (O_3669,N_49900,N_49851);
nand UO_3670 (O_3670,N_49506,N_49953);
nand UO_3671 (O_3671,N_49545,N_49768);
nor UO_3672 (O_3672,N_49910,N_49818);
and UO_3673 (O_3673,N_49953,N_49536);
nor UO_3674 (O_3674,N_49534,N_49901);
and UO_3675 (O_3675,N_49690,N_49809);
or UO_3676 (O_3676,N_49810,N_49559);
nor UO_3677 (O_3677,N_49753,N_49514);
and UO_3678 (O_3678,N_49574,N_49974);
or UO_3679 (O_3679,N_49802,N_49784);
xnor UO_3680 (O_3680,N_49983,N_49705);
nor UO_3681 (O_3681,N_49596,N_49837);
nor UO_3682 (O_3682,N_49908,N_49527);
nor UO_3683 (O_3683,N_49858,N_49908);
nand UO_3684 (O_3684,N_49586,N_49727);
xnor UO_3685 (O_3685,N_49995,N_49852);
nand UO_3686 (O_3686,N_49605,N_49814);
nor UO_3687 (O_3687,N_49826,N_49729);
nand UO_3688 (O_3688,N_49831,N_49982);
and UO_3689 (O_3689,N_49613,N_49661);
xor UO_3690 (O_3690,N_49821,N_49827);
and UO_3691 (O_3691,N_49899,N_49938);
or UO_3692 (O_3692,N_49742,N_49582);
and UO_3693 (O_3693,N_49734,N_49927);
and UO_3694 (O_3694,N_49903,N_49707);
nor UO_3695 (O_3695,N_49724,N_49960);
or UO_3696 (O_3696,N_49939,N_49725);
nor UO_3697 (O_3697,N_49635,N_49810);
nor UO_3698 (O_3698,N_49526,N_49650);
and UO_3699 (O_3699,N_49527,N_49602);
xor UO_3700 (O_3700,N_49937,N_49669);
nor UO_3701 (O_3701,N_49596,N_49957);
nor UO_3702 (O_3702,N_49533,N_49945);
nor UO_3703 (O_3703,N_49881,N_49947);
nand UO_3704 (O_3704,N_49943,N_49559);
or UO_3705 (O_3705,N_49621,N_49734);
or UO_3706 (O_3706,N_49703,N_49760);
and UO_3707 (O_3707,N_49798,N_49865);
or UO_3708 (O_3708,N_49514,N_49868);
or UO_3709 (O_3709,N_49606,N_49613);
and UO_3710 (O_3710,N_49620,N_49943);
nand UO_3711 (O_3711,N_49650,N_49853);
nand UO_3712 (O_3712,N_49627,N_49708);
xor UO_3713 (O_3713,N_49995,N_49543);
and UO_3714 (O_3714,N_49877,N_49818);
nand UO_3715 (O_3715,N_49539,N_49907);
and UO_3716 (O_3716,N_49611,N_49624);
nor UO_3717 (O_3717,N_49785,N_49758);
and UO_3718 (O_3718,N_49857,N_49609);
and UO_3719 (O_3719,N_49897,N_49789);
nor UO_3720 (O_3720,N_49624,N_49571);
nand UO_3721 (O_3721,N_49946,N_49723);
and UO_3722 (O_3722,N_49534,N_49703);
and UO_3723 (O_3723,N_49661,N_49846);
nand UO_3724 (O_3724,N_49740,N_49892);
or UO_3725 (O_3725,N_49733,N_49549);
nand UO_3726 (O_3726,N_49937,N_49860);
and UO_3727 (O_3727,N_49920,N_49695);
nand UO_3728 (O_3728,N_49934,N_49665);
xnor UO_3729 (O_3729,N_49592,N_49826);
nand UO_3730 (O_3730,N_49690,N_49974);
xor UO_3731 (O_3731,N_49622,N_49640);
nand UO_3732 (O_3732,N_49754,N_49890);
xnor UO_3733 (O_3733,N_49625,N_49655);
xor UO_3734 (O_3734,N_49589,N_49756);
xnor UO_3735 (O_3735,N_49872,N_49915);
or UO_3736 (O_3736,N_49896,N_49781);
and UO_3737 (O_3737,N_49772,N_49942);
nand UO_3738 (O_3738,N_49798,N_49781);
nor UO_3739 (O_3739,N_49931,N_49853);
nor UO_3740 (O_3740,N_49586,N_49729);
or UO_3741 (O_3741,N_49582,N_49713);
nor UO_3742 (O_3742,N_49689,N_49879);
and UO_3743 (O_3743,N_49799,N_49986);
nor UO_3744 (O_3744,N_49897,N_49850);
nor UO_3745 (O_3745,N_49851,N_49951);
nor UO_3746 (O_3746,N_49584,N_49744);
and UO_3747 (O_3747,N_49917,N_49830);
and UO_3748 (O_3748,N_49567,N_49797);
or UO_3749 (O_3749,N_49751,N_49854);
xnor UO_3750 (O_3750,N_49790,N_49754);
nor UO_3751 (O_3751,N_49951,N_49575);
nand UO_3752 (O_3752,N_49776,N_49909);
nor UO_3753 (O_3753,N_49762,N_49506);
nor UO_3754 (O_3754,N_49680,N_49954);
xor UO_3755 (O_3755,N_49616,N_49538);
and UO_3756 (O_3756,N_49980,N_49864);
xor UO_3757 (O_3757,N_49540,N_49895);
or UO_3758 (O_3758,N_49595,N_49765);
nand UO_3759 (O_3759,N_49851,N_49741);
and UO_3760 (O_3760,N_49627,N_49656);
or UO_3761 (O_3761,N_49783,N_49828);
or UO_3762 (O_3762,N_49966,N_49790);
xor UO_3763 (O_3763,N_49834,N_49589);
nor UO_3764 (O_3764,N_49720,N_49681);
or UO_3765 (O_3765,N_49805,N_49512);
and UO_3766 (O_3766,N_49618,N_49665);
and UO_3767 (O_3767,N_49531,N_49852);
and UO_3768 (O_3768,N_49930,N_49595);
and UO_3769 (O_3769,N_49678,N_49586);
and UO_3770 (O_3770,N_49687,N_49857);
xnor UO_3771 (O_3771,N_49621,N_49677);
or UO_3772 (O_3772,N_49839,N_49988);
nand UO_3773 (O_3773,N_49560,N_49912);
or UO_3774 (O_3774,N_49770,N_49937);
or UO_3775 (O_3775,N_49755,N_49822);
or UO_3776 (O_3776,N_49680,N_49913);
nor UO_3777 (O_3777,N_49551,N_49614);
or UO_3778 (O_3778,N_49721,N_49998);
nor UO_3779 (O_3779,N_49749,N_49873);
nor UO_3780 (O_3780,N_49844,N_49749);
nor UO_3781 (O_3781,N_49757,N_49616);
or UO_3782 (O_3782,N_49839,N_49803);
nor UO_3783 (O_3783,N_49552,N_49939);
or UO_3784 (O_3784,N_49808,N_49983);
nor UO_3785 (O_3785,N_49562,N_49900);
and UO_3786 (O_3786,N_49709,N_49631);
and UO_3787 (O_3787,N_49541,N_49529);
and UO_3788 (O_3788,N_49840,N_49734);
or UO_3789 (O_3789,N_49649,N_49713);
nand UO_3790 (O_3790,N_49995,N_49955);
xor UO_3791 (O_3791,N_49555,N_49736);
or UO_3792 (O_3792,N_49553,N_49612);
or UO_3793 (O_3793,N_49619,N_49787);
nor UO_3794 (O_3794,N_49828,N_49694);
nand UO_3795 (O_3795,N_49710,N_49728);
nor UO_3796 (O_3796,N_49906,N_49846);
or UO_3797 (O_3797,N_49883,N_49904);
nor UO_3798 (O_3798,N_49768,N_49510);
and UO_3799 (O_3799,N_49840,N_49765);
and UO_3800 (O_3800,N_49682,N_49963);
nor UO_3801 (O_3801,N_49634,N_49996);
nand UO_3802 (O_3802,N_49790,N_49805);
xor UO_3803 (O_3803,N_49900,N_49942);
nand UO_3804 (O_3804,N_49541,N_49746);
nand UO_3805 (O_3805,N_49937,N_49908);
nand UO_3806 (O_3806,N_49846,N_49627);
nand UO_3807 (O_3807,N_49571,N_49695);
and UO_3808 (O_3808,N_49552,N_49870);
and UO_3809 (O_3809,N_49620,N_49532);
nand UO_3810 (O_3810,N_49604,N_49744);
and UO_3811 (O_3811,N_49731,N_49790);
nand UO_3812 (O_3812,N_49553,N_49629);
and UO_3813 (O_3813,N_49810,N_49633);
nand UO_3814 (O_3814,N_49699,N_49697);
nand UO_3815 (O_3815,N_49544,N_49650);
nand UO_3816 (O_3816,N_49770,N_49912);
nor UO_3817 (O_3817,N_49561,N_49674);
or UO_3818 (O_3818,N_49841,N_49776);
and UO_3819 (O_3819,N_49855,N_49907);
nand UO_3820 (O_3820,N_49728,N_49748);
nor UO_3821 (O_3821,N_49959,N_49877);
or UO_3822 (O_3822,N_49991,N_49811);
nand UO_3823 (O_3823,N_49740,N_49745);
nand UO_3824 (O_3824,N_49682,N_49978);
nand UO_3825 (O_3825,N_49803,N_49807);
nor UO_3826 (O_3826,N_49912,N_49515);
nor UO_3827 (O_3827,N_49563,N_49549);
xnor UO_3828 (O_3828,N_49618,N_49597);
nor UO_3829 (O_3829,N_49714,N_49662);
or UO_3830 (O_3830,N_49585,N_49813);
nor UO_3831 (O_3831,N_49764,N_49857);
and UO_3832 (O_3832,N_49765,N_49670);
and UO_3833 (O_3833,N_49775,N_49553);
or UO_3834 (O_3834,N_49996,N_49796);
and UO_3835 (O_3835,N_49650,N_49769);
nor UO_3836 (O_3836,N_49592,N_49890);
nor UO_3837 (O_3837,N_49609,N_49750);
or UO_3838 (O_3838,N_49846,N_49521);
nor UO_3839 (O_3839,N_49505,N_49735);
nor UO_3840 (O_3840,N_49705,N_49541);
and UO_3841 (O_3841,N_49513,N_49970);
nand UO_3842 (O_3842,N_49725,N_49826);
and UO_3843 (O_3843,N_49856,N_49721);
or UO_3844 (O_3844,N_49750,N_49826);
or UO_3845 (O_3845,N_49833,N_49592);
nor UO_3846 (O_3846,N_49894,N_49917);
xnor UO_3847 (O_3847,N_49929,N_49905);
nand UO_3848 (O_3848,N_49903,N_49581);
nand UO_3849 (O_3849,N_49840,N_49824);
nor UO_3850 (O_3850,N_49665,N_49882);
nor UO_3851 (O_3851,N_49669,N_49759);
or UO_3852 (O_3852,N_49978,N_49724);
and UO_3853 (O_3853,N_49897,N_49580);
or UO_3854 (O_3854,N_49983,N_49891);
xor UO_3855 (O_3855,N_49959,N_49719);
and UO_3856 (O_3856,N_49571,N_49590);
nand UO_3857 (O_3857,N_49803,N_49589);
nor UO_3858 (O_3858,N_49594,N_49610);
or UO_3859 (O_3859,N_49643,N_49548);
or UO_3860 (O_3860,N_49942,N_49592);
and UO_3861 (O_3861,N_49900,N_49558);
or UO_3862 (O_3862,N_49785,N_49760);
nand UO_3863 (O_3863,N_49793,N_49685);
or UO_3864 (O_3864,N_49512,N_49515);
or UO_3865 (O_3865,N_49507,N_49972);
or UO_3866 (O_3866,N_49542,N_49648);
and UO_3867 (O_3867,N_49532,N_49643);
nor UO_3868 (O_3868,N_49935,N_49871);
xnor UO_3869 (O_3869,N_49588,N_49531);
or UO_3870 (O_3870,N_49737,N_49671);
nor UO_3871 (O_3871,N_49519,N_49590);
nand UO_3872 (O_3872,N_49514,N_49668);
and UO_3873 (O_3873,N_49923,N_49716);
nand UO_3874 (O_3874,N_49620,N_49537);
nand UO_3875 (O_3875,N_49772,N_49830);
and UO_3876 (O_3876,N_49680,N_49726);
nor UO_3877 (O_3877,N_49863,N_49751);
or UO_3878 (O_3878,N_49594,N_49920);
or UO_3879 (O_3879,N_49679,N_49696);
or UO_3880 (O_3880,N_49751,N_49683);
and UO_3881 (O_3881,N_49524,N_49872);
nand UO_3882 (O_3882,N_49561,N_49694);
or UO_3883 (O_3883,N_49534,N_49533);
and UO_3884 (O_3884,N_49654,N_49746);
nor UO_3885 (O_3885,N_49963,N_49673);
nand UO_3886 (O_3886,N_49893,N_49995);
and UO_3887 (O_3887,N_49934,N_49755);
nand UO_3888 (O_3888,N_49557,N_49708);
nor UO_3889 (O_3889,N_49672,N_49631);
nor UO_3890 (O_3890,N_49617,N_49749);
and UO_3891 (O_3891,N_49582,N_49843);
xnor UO_3892 (O_3892,N_49777,N_49529);
or UO_3893 (O_3893,N_49675,N_49676);
xor UO_3894 (O_3894,N_49964,N_49658);
xor UO_3895 (O_3895,N_49973,N_49999);
xnor UO_3896 (O_3896,N_49832,N_49788);
or UO_3897 (O_3897,N_49914,N_49948);
nand UO_3898 (O_3898,N_49643,N_49995);
xor UO_3899 (O_3899,N_49806,N_49860);
nand UO_3900 (O_3900,N_49767,N_49611);
or UO_3901 (O_3901,N_49752,N_49624);
nand UO_3902 (O_3902,N_49796,N_49593);
or UO_3903 (O_3903,N_49998,N_49546);
and UO_3904 (O_3904,N_49689,N_49786);
and UO_3905 (O_3905,N_49763,N_49739);
nor UO_3906 (O_3906,N_49639,N_49677);
nor UO_3907 (O_3907,N_49518,N_49832);
or UO_3908 (O_3908,N_49832,N_49754);
xor UO_3909 (O_3909,N_49920,N_49600);
xnor UO_3910 (O_3910,N_49930,N_49842);
nand UO_3911 (O_3911,N_49611,N_49921);
and UO_3912 (O_3912,N_49914,N_49659);
or UO_3913 (O_3913,N_49667,N_49700);
and UO_3914 (O_3914,N_49636,N_49971);
and UO_3915 (O_3915,N_49878,N_49516);
and UO_3916 (O_3916,N_49616,N_49986);
nor UO_3917 (O_3917,N_49741,N_49627);
and UO_3918 (O_3918,N_49584,N_49605);
nor UO_3919 (O_3919,N_49680,N_49884);
or UO_3920 (O_3920,N_49913,N_49547);
and UO_3921 (O_3921,N_49740,N_49592);
nand UO_3922 (O_3922,N_49714,N_49947);
nor UO_3923 (O_3923,N_49813,N_49649);
nor UO_3924 (O_3924,N_49985,N_49505);
xor UO_3925 (O_3925,N_49644,N_49813);
and UO_3926 (O_3926,N_49897,N_49889);
xnor UO_3927 (O_3927,N_49860,N_49623);
xor UO_3928 (O_3928,N_49970,N_49818);
nand UO_3929 (O_3929,N_49713,N_49571);
nor UO_3930 (O_3930,N_49879,N_49708);
nand UO_3931 (O_3931,N_49688,N_49671);
xor UO_3932 (O_3932,N_49860,N_49611);
or UO_3933 (O_3933,N_49926,N_49769);
or UO_3934 (O_3934,N_49686,N_49579);
xor UO_3935 (O_3935,N_49560,N_49636);
or UO_3936 (O_3936,N_49867,N_49742);
xnor UO_3937 (O_3937,N_49509,N_49812);
or UO_3938 (O_3938,N_49622,N_49735);
or UO_3939 (O_3939,N_49505,N_49879);
and UO_3940 (O_3940,N_49801,N_49850);
or UO_3941 (O_3941,N_49658,N_49521);
nor UO_3942 (O_3942,N_49617,N_49626);
nand UO_3943 (O_3943,N_49760,N_49643);
nand UO_3944 (O_3944,N_49896,N_49608);
nor UO_3945 (O_3945,N_49631,N_49740);
nand UO_3946 (O_3946,N_49908,N_49697);
nor UO_3947 (O_3947,N_49757,N_49858);
and UO_3948 (O_3948,N_49601,N_49917);
and UO_3949 (O_3949,N_49630,N_49627);
nand UO_3950 (O_3950,N_49835,N_49663);
or UO_3951 (O_3951,N_49831,N_49803);
nand UO_3952 (O_3952,N_49658,N_49580);
or UO_3953 (O_3953,N_49829,N_49859);
and UO_3954 (O_3954,N_49756,N_49739);
or UO_3955 (O_3955,N_49772,N_49858);
xnor UO_3956 (O_3956,N_49504,N_49977);
or UO_3957 (O_3957,N_49845,N_49581);
or UO_3958 (O_3958,N_49558,N_49935);
nor UO_3959 (O_3959,N_49751,N_49738);
or UO_3960 (O_3960,N_49549,N_49565);
nand UO_3961 (O_3961,N_49733,N_49618);
or UO_3962 (O_3962,N_49784,N_49911);
xor UO_3963 (O_3963,N_49871,N_49868);
or UO_3964 (O_3964,N_49789,N_49806);
and UO_3965 (O_3965,N_49856,N_49809);
nor UO_3966 (O_3966,N_49921,N_49805);
and UO_3967 (O_3967,N_49659,N_49767);
nand UO_3968 (O_3968,N_49836,N_49878);
or UO_3969 (O_3969,N_49705,N_49889);
or UO_3970 (O_3970,N_49818,N_49958);
nand UO_3971 (O_3971,N_49856,N_49845);
or UO_3972 (O_3972,N_49888,N_49984);
nor UO_3973 (O_3973,N_49864,N_49604);
nor UO_3974 (O_3974,N_49773,N_49553);
nor UO_3975 (O_3975,N_49755,N_49921);
nor UO_3976 (O_3976,N_49503,N_49910);
nor UO_3977 (O_3977,N_49722,N_49771);
or UO_3978 (O_3978,N_49734,N_49887);
and UO_3979 (O_3979,N_49985,N_49722);
and UO_3980 (O_3980,N_49827,N_49629);
nor UO_3981 (O_3981,N_49615,N_49825);
nand UO_3982 (O_3982,N_49519,N_49880);
nor UO_3983 (O_3983,N_49962,N_49551);
nor UO_3984 (O_3984,N_49869,N_49633);
nor UO_3985 (O_3985,N_49646,N_49633);
or UO_3986 (O_3986,N_49911,N_49757);
and UO_3987 (O_3987,N_49738,N_49872);
xnor UO_3988 (O_3988,N_49567,N_49846);
or UO_3989 (O_3989,N_49639,N_49610);
nand UO_3990 (O_3990,N_49587,N_49934);
or UO_3991 (O_3991,N_49523,N_49992);
and UO_3992 (O_3992,N_49772,N_49521);
nor UO_3993 (O_3993,N_49715,N_49973);
xnor UO_3994 (O_3994,N_49947,N_49718);
nand UO_3995 (O_3995,N_49741,N_49916);
and UO_3996 (O_3996,N_49660,N_49510);
nor UO_3997 (O_3997,N_49813,N_49510);
nand UO_3998 (O_3998,N_49723,N_49885);
or UO_3999 (O_3999,N_49573,N_49764);
nand UO_4000 (O_4000,N_49522,N_49747);
nor UO_4001 (O_4001,N_49713,N_49641);
and UO_4002 (O_4002,N_49551,N_49980);
and UO_4003 (O_4003,N_49527,N_49871);
or UO_4004 (O_4004,N_49554,N_49894);
nand UO_4005 (O_4005,N_49939,N_49699);
or UO_4006 (O_4006,N_49991,N_49791);
nor UO_4007 (O_4007,N_49879,N_49693);
nand UO_4008 (O_4008,N_49574,N_49764);
nor UO_4009 (O_4009,N_49873,N_49639);
xnor UO_4010 (O_4010,N_49746,N_49705);
and UO_4011 (O_4011,N_49794,N_49661);
and UO_4012 (O_4012,N_49860,N_49548);
nand UO_4013 (O_4013,N_49724,N_49710);
nor UO_4014 (O_4014,N_49632,N_49879);
or UO_4015 (O_4015,N_49839,N_49591);
and UO_4016 (O_4016,N_49607,N_49925);
nand UO_4017 (O_4017,N_49855,N_49838);
nand UO_4018 (O_4018,N_49517,N_49721);
and UO_4019 (O_4019,N_49539,N_49908);
and UO_4020 (O_4020,N_49515,N_49672);
xor UO_4021 (O_4021,N_49952,N_49985);
and UO_4022 (O_4022,N_49913,N_49701);
nor UO_4023 (O_4023,N_49592,N_49905);
nand UO_4024 (O_4024,N_49532,N_49944);
nand UO_4025 (O_4025,N_49686,N_49569);
and UO_4026 (O_4026,N_49725,N_49956);
xnor UO_4027 (O_4027,N_49850,N_49799);
xor UO_4028 (O_4028,N_49930,N_49500);
nand UO_4029 (O_4029,N_49697,N_49564);
nor UO_4030 (O_4030,N_49623,N_49956);
nor UO_4031 (O_4031,N_49800,N_49696);
and UO_4032 (O_4032,N_49917,N_49919);
xnor UO_4033 (O_4033,N_49507,N_49536);
or UO_4034 (O_4034,N_49509,N_49701);
or UO_4035 (O_4035,N_49778,N_49752);
nand UO_4036 (O_4036,N_49800,N_49892);
nand UO_4037 (O_4037,N_49700,N_49912);
or UO_4038 (O_4038,N_49504,N_49934);
or UO_4039 (O_4039,N_49756,N_49837);
nand UO_4040 (O_4040,N_49725,N_49663);
and UO_4041 (O_4041,N_49778,N_49674);
nor UO_4042 (O_4042,N_49632,N_49722);
nor UO_4043 (O_4043,N_49881,N_49883);
and UO_4044 (O_4044,N_49853,N_49788);
and UO_4045 (O_4045,N_49774,N_49544);
or UO_4046 (O_4046,N_49735,N_49906);
and UO_4047 (O_4047,N_49635,N_49703);
nand UO_4048 (O_4048,N_49819,N_49674);
and UO_4049 (O_4049,N_49858,N_49588);
or UO_4050 (O_4050,N_49739,N_49748);
or UO_4051 (O_4051,N_49974,N_49859);
xnor UO_4052 (O_4052,N_49514,N_49745);
nor UO_4053 (O_4053,N_49917,N_49816);
and UO_4054 (O_4054,N_49562,N_49890);
and UO_4055 (O_4055,N_49805,N_49578);
nor UO_4056 (O_4056,N_49718,N_49797);
and UO_4057 (O_4057,N_49944,N_49542);
or UO_4058 (O_4058,N_49559,N_49823);
nor UO_4059 (O_4059,N_49641,N_49651);
and UO_4060 (O_4060,N_49828,N_49774);
or UO_4061 (O_4061,N_49840,N_49621);
and UO_4062 (O_4062,N_49835,N_49625);
xor UO_4063 (O_4063,N_49706,N_49991);
or UO_4064 (O_4064,N_49538,N_49717);
nand UO_4065 (O_4065,N_49723,N_49664);
xor UO_4066 (O_4066,N_49902,N_49975);
nor UO_4067 (O_4067,N_49831,N_49791);
and UO_4068 (O_4068,N_49570,N_49510);
and UO_4069 (O_4069,N_49781,N_49707);
nor UO_4070 (O_4070,N_49951,N_49862);
nand UO_4071 (O_4071,N_49547,N_49592);
nor UO_4072 (O_4072,N_49673,N_49838);
and UO_4073 (O_4073,N_49860,N_49610);
and UO_4074 (O_4074,N_49779,N_49504);
nand UO_4075 (O_4075,N_49601,N_49685);
and UO_4076 (O_4076,N_49647,N_49528);
nand UO_4077 (O_4077,N_49672,N_49561);
nand UO_4078 (O_4078,N_49884,N_49827);
or UO_4079 (O_4079,N_49586,N_49824);
or UO_4080 (O_4080,N_49600,N_49581);
and UO_4081 (O_4081,N_49670,N_49817);
and UO_4082 (O_4082,N_49526,N_49992);
nand UO_4083 (O_4083,N_49758,N_49803);
xnor UO_4084 (O_4084,N_49614,N_49819);
nand UO_4085 (O_4085,N_49506,N_49985);
or UO_4086 (O_4086,N_49592,N_49657);
and UO_4087 (O_4087,N_49936,N_49634);
nor UO_4088 (O_4088,N_49815,N_49656);
or UO_4089 (O_4089,N_49537,N_49788);
nand UO_4090 (O_4090,N_49731,N_49704);
nor UO_4091 (O_4091,N_49636,N_49523);
nor UO_4092 (O_4092,N_49650,N_49967);
or UO_4093 (O_4093,N_49818,N_49921);
nor UO_4094 (O_4094,N_49936,N_49753);
and UO_4095 (O_4095,N_49896,N_49595);
or UO_4096 (O_4096,N_49987,N_49555);
or UO_4097 (O_4097,N_49891,N_49985);
or UO_4098 (O_4098,N_49706,N_49668);
xor UO_4099 (O_4099,N_49821,N_49655);
or UO_4100 (O_4100,N_49930,N_49747);
xnor UO_4101 (O_4101,N_49758,N_49910);
nand UO_4102 (O_4102,N_49555,N_49659);
nor UO_4103 (O_4103,N_49815,N_49562);
nor UO_4104 (O_4104,N_49845,N_49724);
or UO_4105 (O_4105,N_49635,N_49550);
nand UO_4106 (O_4106,N_49989,N_49588);
nand UO_4107 (O_4107,N_49596,N_49823);
or UO_4108 (O_4108,N_49591,N_49946);
or UO_4109 (O_4109,N_49748,N_49599);
and UO_4110 (O_4110,N_49851,N_49511);
nor UO_4111 (O_4111,N_49860,N_49862);
nor UO_4112 (O_4112,N_49747,N_49525);
nand UO_4113 (O_4113,N_49815,N_49768);
and UO_4114 (O_4114,N_49882,N_49551);
and UO_4115 (O_4115,N_49594,N_49834);
nand UO_4116 (O_4116,N_49951,N_49774);
xnor UO_4117 (O_4117,N_49607,N_49939);
and UO_4118 (O_4118,N_49871,N_49909);
nor UO_4119 (O_4119,N_49604,N_49603);
or UO_4120 (O_4120,N_49900,N_49656);
and UO_4121 (O_4121,N_49555,N_49985);
and UO_4122 (O_4122,N_49806,N_49550);
nand UO_4123 (O_4123,N_49603,N_49935);
or UO_4124 (O_4124,N_49590,N_49988);
or UO_4125 (O_4125,N_49609,N_49997);
and UO_4126 (O_4126,N_49551,N_49513);
xnor UO_4127 (O_4127,N_49552,N_49516);
and UO_4128 (O_4128,N_49813,N_49641);
or UO_4129 (O_4129,N_49718,N_49780);
or UO_4130 (O_4130,N_49634,N_49559);
xnor UO_4131 (O_4131,N_49840,N_49808);
or UO_4132 (O_4132,N_49503,N_49906);
nor UO_4133 (O_4133,N_49878,N_49579);
nor UO_4134 (O_4134,N_49527,N_49577);
nand UO_4135 (O_4135,N_49648,N_49796);
and UO_4136 (O_4136,N_49580,N_49963);
nand UO_4137 (O_4137,N_49502,N_49597);
or UO_4138 (O_4138,N_49853,N_49508);
nor UO_4139 (O_4139,N_49803,N_49703);
nand UO_4140 (O_4140,N_49602,N_49784);
or UO_4141 (O_4141,N_49698,N_49875);
nor UO_4142 (O_4142,N_49568,N_49744);
nand UO_4143 (O_4143,N_49604,N_49898);
nand UO_4144 (O_4144,N_49727,N_49867);
nor UO_4145 (O_4145,N_49767,N_49692);
and UO_4146 (O_4146,N_49656,N_49585);
nand UO_4147 (O_4147,N_49920,N_49741);
and UO_4148 (O_4148,N_49607,N_49777);
nand UO_4149 (O_4149,N_49927,N_49735);
nand UO_4150 (O_4150,N_49767,N_49819);
and UO_4151 (O_4151,N_49749,N_49559);
and UO_4152 (O_4152,N_49872,N_49774);
and UO_4153 (O_4153,N_49964,N_49574);
nor UO_4154 (O_4154,N_49853,N_49610);
nand UO_4155 (O_4155,N_49783,N_49970);
or UO_4156 (O_4156,N_49754,N_49662);
nand UO_4157 (O_4157,N_49537,N_49697);
nor UO_4158 (O_4158,N_49582,N_49686);
or UO_4159 (O_4159,N_49652,N_49775);
and UO_4160 (O_4160,N_49658,N_49929);
nand UO_4161 (O_4161,N_49967,N_49956);
nor UO_4162 (O_4162,N_49559,N_49816);
nor UO_4163 (O_4163,N_49546,N_49645);
and UO_4164 (O_4164,N_49714,N_49549);
or UO_4165 (O_4165,N_49519,N_49538);
xor UO_4166 (O_4166,N_49941,N_49551);
nor UO_4167 (O_4167,N_49871,N_49914);
or UO_4168 (O_4168,N_49791,N_49692);
nor UO_4169 (O_4169,N_49815,N_49597);
nor UO_4170 (O_4170,N_49809,N_49619);
nand UO_4171 (O_4171,N_49876,N_49503);
nand UO_4172 (O_4172,N_49815,N_49606);
and UO_4173 (O_4173,N_49946,N_49595);
xnor UO_4174 (O_4174,N_49750,N_49683);
or UO_4175 (O_4175,N_49692,N_49710);
and UO_4176 (O_4176,N_49718,N_49748);
xnor UO_4177 (O_4177,N_49906,N_49507);
or UO_4178 (O_4178,N_49782,N_49973);
and UO_4179 (O_4179,N_49738,N_49730);
nand UO_4180 (O_4180,N_49562,N_49590);
or UO_4181 (O_4181,N_49978,N_49806);
nor UO_4182 (O_4182,N_49694,N_49520);
nand UO_4183 (O_4183,N_49825,N_49785);
xnor UO_4184 (O_4184,N_49651,N_49938);
nand UO_4185 (O_4185,N_49992,N_49874);
and UO_4186 (O_4186,N_49988,N_49552);
and UO_4187 (O_4187,N_49632,N_49808);
nor UO_4188 (O_4188,N_49889,N_49850);
nand UO_4189 (O_4189,N_49945,N_49744);
nand UO_4190 (O_4190,N_49518,N_49866);
xor UO_4191 (O_4191,N_49729,N_49733);
or UO_4192 (O_4192,N_49597,N_49997);
or UO_4193 (O_4193,N_49900,N_49905);
and UO_4194 (O_4194,N_49826,N_49841);
or UO_4195 (O_4195,N_49915,N_49747);
nor UO_4196 (O_4196,N_49816,N_49848);
nor UO_4197 (O_4197,N_49572,N_49588);
nand UO_4198 (O_4198,N_49551,N_49584);
and UO_4199 (O_4199,N_49864,N_49820);
nor UO_4200 (O_4200,N_49861,N_49566);
or UO_4201 (O_4201,N_49969,N_49676);
and UO_4202 (O_4202,N_49641,N_49733);
and UO_4203 (O_4203,N_49787,N_49621);
xnor UO_4204 (O_4204,N_49584,N_49560);
and UO_4205 (O_4205,N_49886,N_49671);
or UO_4206 (O_4206,N_49897,N_49607);
nand UO_4207 (O_4207,N_49966,N_49962);
and UO_4208 (O_4208,N_49684,N_49936);
or UO_4209 (O_4209,N_49539,N_49990);
nand UO_4210 (O_4210,N_49525,N_49726);
nor UO_4211 (O_4211,N_49926,N_49562);
xnor UO_4212 (O_4212,N_49719,N_49988);
and UO_4213 (O_4213,N_49758,N_49646);
or UO_4214 (O_4214,N_49982,N_49691);
or UO_4215 (O_4215,N_49533,N_49629);
or UO_4216 (O_4216,N_49554,N_49827);
nand UO_4217 (O_4217,N_49805,N_49547);
and UO_4218 (O_4218,N_49758,N_49744);
nor UO_4219 (O_4219,N_49646,N_49608);
or UO_4220 (O_4220,N_49577,N_49680);
nor UO_4221 (O_4221,N_49826,N_49879);
nand UO_4222 (O_4222,N_49949,N_49765);
and UO_4223 (O_4223,N_49985,N_49529);
nand UO_4224 (O_4224,N_49914,N_49919);
nand UO_4225 (O_4225,N_49610,N_49645);
and UO_4226 (O_4226,N_49985,N_49560);
or UO_4227 (O_4227,N_49834,N_49878);
and UO_4228 (O_4228,N_49585,N_49878);
xor UO_4229 (O_4229,N_49790,N_49900);
nand UO_4230 (O_4230,N_49656,N_49883);
nand UO_4231 (O_4231,N_49893,N_49708);
nand UO_4232 (O_4232,N_49800,N_49593);
nand UO_4233 (O_4233,N_49561,N_49643);
nand UO_4234 (O_4234,N_49853,N_49693);
nand UO_4235 (O_4235,N_49931,N_49857);
or UO_4236 (O_4236,N_49692,N_49881);
and UO_4237 (O_4237,N_49691,N_49884);
or UO_4238 (O_4238,N_49868,N_49817);
or UO_4239 (O_4239,N_49816,N_49923);
nand UO_4240 (O_4240,N_49645,N_49665);
xor UO_4241 (O_4241,N_49523,N_49718);
nor UO_4242 (O_4242,N_49745,N_49621);
nand UO_4243 (O_4243,N_49580,N_49760);
and UO_4244 (O_4244,N_49918,N_49891);
nand UO_4245 (O_4245,N_49767,N_49708);
nand UO_4246 (O_4246,N_49852,N_49682);
and UO_4247 (O_4247,N_49733,N_49672);
and UO_4248 (O_4248,N_49791,N_49939);
or UO_4249 (O_4249,N_49623,N_49513);
xnor UO_4250 (O_4250,N_49723,N_49973);
nand UO_4251 (O_4251,N_49711,N_49852);
nand UO_4252 (O_4252,N_49759,N_49709);
nor UO_4253 (O_4253,N_49981,N_49840);
or UO_4254 (O_4254,N_49562,N_49957);
nor UO_4255 (O_4255,N_49844,N_49578);
nor UO_4256 (O_4256,N_49881,N_49700);
nand UO_4257 (O_4257,N_49815,N_49666);
or UO_4258 (O_4258,N_49730,N_49764);
nand UO_4259 (O_4259,N_49730,N_49872);
and UO_4260 (O_4260,N_49848,N_49821);
or UO_4261 (O_4261,N_49965,N_49661);
nand UO_4262 (O_4262,N_49979,N_49582);
nand UO_4263 (O_4263,N_49942,N_49578);
and UO_4264 (O_4264,N_49638,N_49548);
or UO_4265 (O_4265,N_49743,N_49534);
nor UO_4266 (O_4266,N_49686,N_49793);
nor UO_4267 (O_4267,N_49661,N_49735);
nand UO_4268 (O_4268,N_49508,N_49519);
xnor UO_4269 (O_4269,N_49821,N_49515);
nor UO_4270 (O_4270,N_49673,N_49505);
nand UO_4271 (O_4271,N_49990,N_49905);
and UO_4272 (O_4272,N_49754,N_49877);
nand UO_4273 (O_4273,N_49600,N_49756);
nand UO_4274 (O_4274,N_49538,N_49637);
nor UO_4275 (O_4275,N_49595,N_49548);
nor UO_4276 (O_4276,N_49612,N_49993);
nor UO_4277 (O_4277,N_49500,N_49878);
or UO_4278 (O_4278,N_49883,N_49758);
xnor UO_4279 (O_4279,N_49758,N_49623);
nand UO_4280 (O_4280,N_49532,N_49956);
nor UO_4281 (O_4281,N_49739,N_49590);
nand UO_4282 (O_4282,N_49731,N_49836);
nand UO_4283 (O_4283,N_49809,N_49657);
and UO_4284 (O_4284,N_49812,N_49999);
nor UO_4285 (O_4285,N_49747,N_49822);
and UO_4286 (O_4286,N_49541,N_49906);
and UO_4287 (O_4287,N_49688,N_49935);
nand UO_4288 (O_4288,N_49681,N_49831);
xnor UO_4289 (O_4289,N_49764,N_49781);
and UO_4290 (O_4290,N_49661,N_49612);
and UO_4291 (O_4291,N_49900,N_49717);
or UO_4292 (O_4292,N_49655,N_49830);
or UO_4293 (O_4293,N_49707,N_49558);
nand UO_4294 (O_4294,N_49570,N_49854);
and UO_4295 (O_4295,N_49798,N_49733);
and UO_4296 (O_4296,N_49984,N_49980);
and UO_4297 (O_4297,N_49594,N_49661);
or UO_4298 (O_4298,N_49871,N_49824);
nand UO_4299 (O_4299,N_49606,N_49799);
or UO_4300 (O_4300,N_49655,N_49569);
nor UO_4301 (O_4301,N_49810,N_49812);
or UO_4302 (O_4302,N_49731,N_49918);
nand UO_4303 (O_4303,N_49960,N_49593);
and UO_4304 (O_4304,N_49984,N_49850);
or UO_4305 (O_4305,N_49630,N_49688);
and UO_4306 (O_4306,N_49787,N_49900);
or UO_4307 (O_4307,N_49556,N_49729);
nor UO_4308 (O_4308,N_49780,N_49700);
nand UO_4309 (O_4309,N_49520,N_49940);
and UO_4310 (O_4310,N_49908,N_49748);
and UO_4311 (O_4311,N_49512,N_49798);
and UO_4312 (O_4312,N_49886,N_49878);
or UO_4313 (O_4313,N_49678,N_49562);
and UO_4314 (O_4314,N_49762,N_49901);
or UO_4315 (O_4315,N_49914,N_49655);
nand UO_4316 (O_4316,N_49785,N_49929);
nand UO_4317 (O_4317,N_49899,N_49961);
and UO_4318 (O_4318,N_49687,N_49692);
nand UO_4319 (O_4319,N_49854,N_49775);
nor UO_4320 (O_4320,N_49543,N_49667);
nor UO_4321 (O_4321,N_49604,N_49930);
and UO_4322 (O_4322,N_49856,N_49867);
and UO_4323 (O_4323,N_49954,N_49544);
or UO_4324 (O_4324,N_49549,N_49532);
and UO_4325 (O_4325,N_49604,N_49613);
nor UO_4326 (O_4326,N_49852,N_49765);
or UO_4327 (O_4327,N_49633,N_49531);
nand UO_4328 (O_4328,N_49752,N_49775);
nor UO_4329 (O_4329,N_49975,N_49927);
or UO_4330 (O_4330,N_49784,N_49890);
and UO_4331 (O_4331,N_49864,N_49880);
nand UO_4332 (O_4332,N_49555,N_49905);
nand UO_4333 (O_4333,N_49513,N_49894);
or UO_4334 (O_4334,N_49838,N_49794);
xnor UO_4335 (O_4335,N_49925,N_49789);
or UO_4336 (O_4336,N_49564,N_49618);
and UO_4337 (O_4337,N_49551,N_49984);
nor UO_4338 (O_4338,N_49975,N_49587);
xor UO_4339 (O_4339,N_49559,N_49713);
and UO_4340 (O_4340,N_49694,N_49582);
and UO_4341 (O_4341,N_49835,N_49516);
nand UO_4342 (O_4342,N_49574,N_49935);
nor UO_4343 (O_4343,N_49851,N_49863);
nor UO_4344 (O_4344,N_49649,N_49751);
xor UO_4345 (O_4345,N_49624,N_49857);
and UO_4346 (O_4346,N_49527,N_49813);
and UO_4347 (O_4347,N_49626,N_49655);
or UO_4348 (O_4348,N_49548,N_49724);
nand UO_4349 (O_4349,N_49509,N_49747);
nor UO_4350 (O_4350,N_49955,N_49871);
nor UO_4351 (O_4351,N_49826,N_49980);
nor UO_4352 (O_4352,N_49769,N_49503);
or UO_4353 (O_4353,N_49740,N_49776);
nor UO_4354 (O_4354,N_49732,N_49743);
and UO_4355 (O_4355,N_49800,N_49955);
or UO_4356 (O_4356,N_49545,N_49509);
or UO_4357 (O_4357,N_49814,N_49698);
xor UO_4358 (O_4358,N_49875,N_49805);
or UO_4359 (O_4359,N_49526,N_49811);
or UO_4360 (O_4360,N_49631,N_49959);
xor UO_4361 (O_4361,N_49932,N_49515);
nor UO_4362 (O_4362,N_49614,N_49654);
or UO_4363 (O_4363,N_49805,N_49636);
nand UO_4364 (O_4364,N_49548,N_49525);
nor UO_4365 (O_4365,N_49505,N_49871);
nand UO_4366 (O_4366,N_49582,N_49736);
nor UO_4367 (O_4367,N_49616,N_49596);
or UO_4368 (O_4368,N_49787,N_49616);
or UO_4369 (O_4369,N_49530,N_49691);
and UO_4370 (O_4370,N_49882,N_49838);
nand UO_4371 (O_4371,N_49934,N_49682);
or UO_4372 (O_4372,N_49823,N_49589);
or UO_4373 (O_4373,N_49568,N_49709);
or UO_4374 (O_4374,N_49532,N_49870);
nor UO_4375 (O_4375,N_49675,N_49922);
or UO_4376 (O_4376,N_49950,N_49771);
nor UO_4377 (O_4377,N_49879,N_49564);
and UO_4378 (O_4378,N_49616,N_49805);
nand UO_4379 (O_4379,N_49936,N_49870);
nor UO_4380 (O_4380,N_49622,N_49988);
nor UO_4381 (O_4381,N_49501,N_49638);
nor UO_4382 (O_4382,N_49699,N_49539);
nand UO_4383 (O_4383,N_49985,N_49896);
and UO_4384 (O_4384,N_49833,N_49896);
or UO_4385 (O_4385,N_49607,N_49830);
and UO_4386 (O_4386,N_49657,N_49577);
or UO_4387 (O_4387,N_49985,N_49513);
nor UO_4388 (O_4388,N_49651,N_49908);
or UO_4389 (O_4389,N_49989,N_49794);
nand UO_4390 (O_4390,N_49774,N_49816);
and UO_4391 (O_4391,N_49653,N_49500);
or UO_4392 (O_4392,N_49942,N_49545);
nor UO_4393 (O_4393,N_49714,N_49593);
nand UO_4394 (O_4394,N_49833,N_49593);
nand UO_4395 (O_4395,N_49768,N_49764);
nand UO_4396 (O_4396,N_49504,N_49657);
or UO_4397 (O_4397,N_49533,N_49609);
or UO_4398 (O_4398,N_49809,N_49681);
nand UO_4399 (O_4399,N_49812,N_49873);
and UO_4400 (O_4400,N_49572,N_49731);
and UO_4401 (O_4401,N_49965,N_49532);
or UO_4402 (O_4402,N_49750,N_49814);
and UO_4403 (O_4403,N_49562,N_49745);
xnor UO_4404 (O_4404,N_49950,N_49668);
xor UO_4405 (O_4405,N_49724,N_49722);
and UO_4406 (O_4406,N_49679,N_49795);
xnor UO_4407 (O_4407,N_49847,N_49912);
nor UO_4408 (O_4408,N_49665,N_49847);
or UO_4409 (O_4409,N_49701,N_49625);
xnor UO_4410 (O_4410,N_49840,N_49756);
or UO_4411 (O_4411,N_49531,N_49574);
or UO_4412 (O_4412,N_49834,N_49697);
nand UO_4413 (O_4413,N_49905,N_49632);
xnor UO_4414 (O_4414,N_49565,N_49901);
and UO_4415 (O_4415,N_49920,N_49871);
xor UO_4416 (O_4416,N_49503,N_49767);
xor UO_4417 (O_4417,N_49772,N_49753);
nand UO_4418 (O_4418,N_49539,N_49986);
and UO_4419 (O_4419,N_49961,N_49530);
xnor UO_4420 (O_4420,N_49632,N_49852);
and UO_4421 (O_4421,N_49696,N_49803);
nand UO_4422 (O_4422,N_49937,N_49508);
xnor UO_4423 (O_4423,N_49772,N_49833);
and UO_4424 (O_4424,N_49873,N_49576);
or UO_4425 (O_4425,N_49753,N_49735);
and UO_4426 (O_4426,N_49880,N_49682);
or UO_4427 (O_4427,N_49755,N_49788);
or UO_4428 (O_4428,N_49677,N_49700);
and UO_4429 (O_4429,N_49915,N_49560);
xor UO_4430 (O_4430,N_49636,N_49858);
nor UO_4431 (O_4431,N_49605,N_49927);
nand UO_4432 (O_4432,N_49649,N_49695);
or UO_4433 (O_4433,N_49690,N_49941);
nor UO_4434 (O_4434,N_49604,N_49673);
nand UO_4435 (O_4435,N_49609,N_49800);
and UO_4436 (O_4436,N_49935,N_49896);
nand UO_4437 (O_4437,N_49810,N_49977);
and UO_4438 (O_4438,N_49626,N_49964);
and UO_4439 (O_4439,N_49843,N_49513);
nand UO_4440 (O_4440,N_49650,N_49525);
nor UO_4441 (O_4441,N_49794,N_49891);
nor UO_4442 (O_4442,N_49690,N_49602);
and UO_4443 (O_4443,N_49594,N_49898);
xnor UO_4444 (O_4444,N_49544,N_49645);
nor UO_4445 (O_4445,N_49522,N_49812);
or UO_4446 (O_4446,N_49779,N_49670);
or UO_4447 (O_4447,N_49524,N_49580);
nor UO_4448 (O_4448,N_49841,N_49778);
nor UO_4449 (O_4449,N_49655,N_49687);
nor UO_4450 (O_4450,N_49640,N_49912);
and UO_4451 (O_4451,N_49625,N_49886);
nand UO_4452 (O_4452,N_49778,N_49507);
nor UO_4453 (O_4453,N_49775,N_49546);
and UO_4454 (O_4454,N_49973,N_49643);
and UO_4455 (O_4455,N_49642,N_49997);
nor UO_4456 (O_4456,N_49907,N_49505);
and UO_4457 (O_4457,N_49937,N_49759);
xnor UO_4458 (O_4458,N_49806,N_49815);
and UO_4459 (O_4459,N_49507,N_49948);
and UO_4460 (O_4460,N_49682,N_49849);
or UO_4461 (O_4461,N_49626,N_49909);
nor UO_4462 (O_4462,N_49533,N_49950);
nor UO_4463 (O_4463,N_49505,N_49996);
or UO_4464 (O_4464,N_49827,N_49729);
and UO_4465 (O_4465,N_49875,N_49956);
and UO_4466 (O_4466,N_49655,N_49607);
and UO_4467 (O_4467,N_49665,N_49671);
or UO_4468 (O_4468,N_49753,N_49813);
and UO_4469 (O_4469,N_49745,N_49623);
and UO_4470 (O_4470,N_49746,N_49781);
and UO_4471 (O_4471,N_49782,N_49968);
or UO_4472 (O_4472,N_49926,N_49783);
nor UO_4473 (O_4473,N_49575,N_49516);
nand UO_4474 (O_4474,N_49797,N_49937);
or UO_4475 (O_4475,N_49875,N_49861);
nand UO_4476 (O_4476,N_49512,N_49943);
nor UO_4477 (O_4477,N_49838,N_49743);
or UO_4478 (O_4478,N_49628,N_49962);
or UO_4479 (O_4479,N_49572,N_49927);
and UO_4480 (O_4480,N_49956,N_49584);
or UO_4481 (O_4481,N_49687,N_49755);
or UO_4482 (O_4482,N_49714,N_49576);
nand UO_4483 (O_4483,N_49801,N_49722);
and UO_4484 (O_4484,N_49800,N_49548);
and UO_4485 (O_4485,N_49513,N_49718);
or UO_4486 (O_4486,N_49558,N_49689);
nand UO_4487 (O_4487,N_49904,N_49915);
or UO_4488 (O_4488,N_49697,N_49606);
nand UO_4489 (O_4489,N_49779,N_49678);
or UO_4490 (O_4490,N_49991,N_49777);
and UO_4491 (O_4491,N_49883,N_49813);
nor UO_4492 (O_4492,N_49526,N_49604);
or UO_4493 (O_4493,N_49536,N_49531);
and UO_4494 (O_4494,N_49555,N_49746);
and UO_4495 (O_4495,N_49991,N_49679);
nand UO_4496 (O_4496,N_49670,N_49815);
and UO_4497 (O_4497,N_49729,N_49591);
or UO_4498 (O_4498,N_49668,N_49799);
nor UO_4499 (O_4499,N_49764,N_49698);
or UO_4500 (O_4500,N_49826,N_49831);
nor UO_4501 (O_4501,N_49753,N_49799);
nand UO_4502 (O_4502,N_49507,N_49869);
or UO_4503 (O_4503,N_49846,N_49731);
nand UO_4504 (O_4504,N_49533,N_49633);
xnor UO_4505 (O_4505,N_49523,N_49940);
and UO_4506 (O_4506,N_49587,N_49859);
and UO_4507 (O_4507,N_49783,N_49739);
xor UO_4508 (O_4508,N_49937,N_49883);
nand UO_4509 (O_4509,N_49755,N_49548);
or UO_4510 (O_4510,N_49582,N_49948);
or UO_4511 (O_4511,N_49739,N_49618);
nand UO_4512 (O_4512,N_49673,N_49813);
and UO_4513 (O_4513,N_49692,N_49843);
xor UO_4514 (O_4514,N_49976,N_49612);
or UO_4515 (O_4515,N_49566,N_49611);
xnor UO_4516 (O_4516,N_49690,N_49954);
or UO_4517 (O_4517,N_49694,N_49518);
xnor UO_4518 (O_4518,N_49922,N_49966);
or UO_4519 (O_4519,N_49542,N_49704);
nand UO_4520 (O_4520,N_49900,N_49629);
nand UO_4521 (O_4521,N_49503,N_49556);
nor UO_4522 (O_4522,N_49572,N_49903);
nor UO_4523 (O_4523,N_49810,N_49841);
nor UO_4524 (O_4524,N_49600,N_49715);
or UO_4525 (O_4525,N_49811,N_49603);
and UO_4526 (O_4526,N_49731,N_49973);
xnor UO_4527 (O_4527,N_49777,N_49744);
and UO_4528 (O_4528,N_49609,N_49831);
nand UO_4529 (O_4529,N_49863,N_49889);
and UO_4530 (O_4530,N_49654,N_49835);
and UO_4531 (O_4531,N_49915,N_49582);
nand UO_4532 (O_4532,N_49891,N_49712);
nor UO_4533 (O_4533,N_49620,N_49741);
and UO_4534 (O_4534,N_49784,N_49771);
and UO_4535 (O_4535,N_49947,N_49880);
nor UO_4536 (O_4536,N_49531,N_49749);
nand UO_4537 (O_4537,N_49840,N_49651);
nand UO_4538 (O_4538,N_49865,N_49891);
or UO_4539 (O_4539,N_49528,N_49642);
and UO_4540 (O_4540,N_49861,N_49797);
nand UO_4541 (O_4541,N_49900,N_49842);
or UO_4542 (O_4542,N_49533,N_49978);
nand UO_4543 (O_4543,N_49948,N_49856);
nand UO_4544 (O_4544,N_49722,N_49908);
and UO_4545 (O_4545,N_49873,N_49958);
and UO_4546 (O_4546,N_49972,N_49913);
or UO_4547 (O_4547,N_49690,N_49547);
nand UO_4548 (O_4548,N_49767,N_49812);
nand UO_4549 (O_4549,N_49996,N_49907);
xor UO_4550 (O_4550,N_49868,N_49892);
nor UO_4551 (O_4551,N_49617,N_49517);
and UO_4552 (O_4552,N_49711,N_49788);
or UO_4553 (O_4553,N_49898,N_49700);
nand UO_4554 (O_4554,N_49662,N_49880);
and UO_4555 (O_4555,N_49999,N_49559);
nor UO_4556 (O_4556,N_49965,N_49579);
or UO_4557 (O_4557,N_49968,N_49505);
nand UO_4558 (O_4558,N_49791,N_49560);
nand UO_4559 (O_4559,N_49527,N_49880);
xnor UO_4560 (O_4560,N_49514,N_49951);
xor UO_4561 (O_4561,N_49613,N_49758);
nor UO_4562 (O_4562,N_49645,N_49704);
nor UO_4563 (O_4563,N_49847,N_49500);
nand UO_4564 (O_4564,N_49979,N_49781);
and UO_4565 (O_4565,N_49738,N_49574);
or UO_4566 (O_4566,N_49889,N_49971);
nand UO_4567 (O_4567,N_49536,N_49576);
nor UO_4568 (O_4568,N_49889,N_49959);
nor UO_4569 (O_4569,N_49595,N_49940);
or UO_4570 (O_4570,N_49595,N_49795);
nor UO_4571 (O_4571,N_49924,N_49531);
or UO_4572 (O_4572,N_49531,N_49653);
or UO_4573 (O_4573,N_49911,N_49839);
and UO_4574 (O_4574,N_49717,N_49666);
or UO_4575 (O_4575,N_49952,N_49732);
and UO_4576 (O_4576,N_49991,N_49704);
nor UO_4577 (O_4577,N_49710,N_49860);
nand UO_4578 (O_4578,N_49679,N_49873);
and UO_4579 (O_4579,N_49794,N_49969);
nand UO_4580 (O_4580,N_49843,N_49581);
or UO_4581 (O_4581,N_49774,N_49794);
and UO_4582 (O_4582,N_49566,N_49879);
xor UO_4583 (O_4583,N_49752,N_49930);
or UO_4584 (O_4584,N_49624,N_49533);
nand UO_4585 (O_4585,N_49944,N_49962);
or UO_4586 (O_4586,N_49552,N_49578);
or UO_4587 (O_4587,N_49992,N_49755);
or UO_4588 (O_4588,N_49756,N_49825);
and UO_4589 (O_4589,N_49633,N_49825);
or UO_4590 (O_4590,N_49794,N_49990);
nand UO_4591 (O_4591,N_49538,N_49960);
or UO_4592 (O_4592,N_49967,N_49728);
or UO_4593 (O_4593,N_49895,N_49864);
nor UO_4594 (O_4594,N_49585,N_49648);
nand UO_4595 (O_4595,N_49721,N_49571);
nand UO_4596 (O_4596,N_49805,N_49717);
and UO_4597 (O_4597,N_49630,N_49938);
nand UO_4598 (O_4598,N_49792,N_49606);
or UO_4599 (O_4599,N_49820,N_49964);
nor UO_4600 (O_4600,N_49519,N_49641);
and UO_4601 (O_4601,N_49795,N_49926);
xor UO_4602 (O_4602,N_49593,N_49803);
nor UO_4603 (O_4603,N_49625,N_49774);
and UO_4604 (O_4604,N_49755,N_49909);
and UO_4605 (O_4605,N_49835,N_49696);
xor UO_4606 (O_4606,N_49960,N_49772);
and UO_4607 (O_4607,N_49538,N_49555);
nand UO_4608 (O_4608,N_49601,N_49526);
or UO_4609 (O_4609,N_49671,N_49667);
or UO_4610 (O_4610,N_49947,N_49609);
or UO_4611 (O_4611,N_49867,N_49782);
and UO_4612 (O_4612,N_49866,N_49714);
or UO_4613 (O_4613,N_49892,N_49865);
and UO_4614 (O_4614,N_49731,N_49925);
and UO_4615 (O_4615,N_49623,N_49891);
or UO_4616 (O_4616,N_49994,N_49550);
nand UO_4617 (O_4617,N_49610,N_49623);
and UO_4618 (O_4618,N_49849,N_49922);
xor UO_4619 (O_4619,N_49989,N_49876);
xor UO_4620 (O_4620,N_49638,N_49565);
or UO_4621 (O_4621,N_49667,N_49980);
and UO_4622 (O_4622,N_49930,N_49792);
or UO_4623 (O_4623,N_49968,N_49820);
and UO_4624 (O_4624,N_49611,N_49602);
or UO_4625 (O_4625,N_49742,N_49996);
nand UO_4626 (O_4626,N_49867,N_49787);
xor UO_4627 (O_4627,N_49763,N_49817);
or UO_4628 (O_4628,N_49942,N_49913);
nor UO_4629 (O_4629,N_49681,N_49975);
nand UO_4630 (O_4630,N_49784,N_49975);
nand UO_4631 (O_4631,N_49965,N_49842);
nand UO_4632 (O_4632,N_49627,N_49613);
and UO_4633 (O_4633,N_49666,N_49513);
and UO_4634 (O_4634,N_49567,N_49845);
and UO_4635 (O_4635,N_49950,N_49973);
and UO_4636 (O_4636,N_49902,N_49578);
nand UO_4637 (O_4637,N_49559,N_49522);
xor UO_4638 (O_4638,N_49506,N_49798);
and UO_4639 (O_4639,N_49644,N_49819);
nor UO_4640 (O_4640,N_49863,N_49939);
nand UO_4641 (O_4641,N_49822,N_49749);
and UO_4642 (O_4642,N_49519,N_49639);
or UO_4643 (O_4643,N_49880,N_49906);
and UO_4644 (O_4644,N_49917,N_49564);
and UO_4645 (O_4645,N_49677,N_49662);
nand UO_4646 (O_4646,N_49537,N_49687);
and UO_4647 (O_4647,N_49532,N_49629);
and UO_4648 (O_4648,N_49868,N_49543);
and UO_4649 (O_4649,N_49636,N_49770);
and UO_4650 (O_4650,N_49695,N_49750);
nor UO_4651 (O_4651,N_49844,N_49684);
xnor UO_4652 (O_4652,N_49633,N_49684);
or UO_4653 (O_4653,N_49885,N_49981);
nor UO_4654 (O_4654,N_49759,N_49682);
or UO_4655 (O_4655,N_49593,N_49971);
nand UO_4656 (O_4656,N_49829,N_49658);
and UO_4657 (O_4657,N_49817,N_49798);
nand UO_4658 (O_4658,N_49634,N_49976);
nor UO_4659 (O_4659,N_49862,N_49670);
or UO_4660 (O_4660,N_49985,N_49694);
or UO_4661 (O_4661,N_49932,N_49938);
nor UO_4662 (O_4662,N_49592,N_49537);
nand UO_4663 (O_4663,N_49770,N_49761);
and UO_4664 (O_4664,N_49512,N_49583);
nor UO_4665 (O_4665,N_49778,N_49872);
xor UO_4666 (O_4666,N_49698,N_49628);
nor UO_4667 (O_4667,N_49910,N_49710);
nand UO_4668 (O_4668,N_49668,N_49568);
xor UO_4669 (O_4669,N_49574,N_49644);
xor UO_4670 (O_4670,N_49742,N_49621);
xnor UO_4671 (O_4671,N_49564,N_49857);
nand UO_4672 (O_4672,N_49804,N_49651);
nand UO_4673 (O_4673,N_49743,N_49527);
and UO_4674 (O_4674,N_49724,N_49588);
nor UO_4675 (O_4675,N_49951,N_49538);
nand UO_4676 (O_4676,N_49912,N_49550);
nand UO_4677 (O_4677,N_49963,N_49575);
nor UO_4678 (O_4678,N_49550,N_49823);
and UO_4679 (O_4679,N_49853,N_49818);
nand UO_4680 (O_4680,N_49521,N_49917);
and UO_4681 (O_4681,N_49729,N_49934);
nand UO_4682 (O_4682,N_49557,N_49580);
nand UO_4683 (O_4683,N_49501,N_49837);
nand UO_4684 (O_4684,N_49873,N_49803);
and UO_4685 (O_4685,N_49936,N_49992);
or UO_4686 (O_4686,N_49583,N_49533);
or UO_4687 (O_4687,N_49512,N_49546);
nand UO_4688 (O_4688,N_49581,N_49965);
or UO_4689 (O_4689,N_49889,N_49545);
nand UO_4690 (O_4690,N_49689,N_49532);
nand UO_4691 (O_4691,N_49865,N_49537);
and UO_4692 (O_4692,N_49704,N_49814);
or UO_4693 (O_4693,N_49826,N_49914);
or UO_4694 (O_4694,N_49724,N_49813);
nor UO_4695 (O_4695,N_49910,N_49621);
nand UO_4696 (O_4696,N_49649,N_49707);
nor UO_4697 (O_4697,N_49960,N_49816);
and UO_4698 (O_4698,N_49892,N_49956);
or UO_4699 (O_4699,N_49822,N_49978);
nand UO_4700 (O_4700,N_49731,N_49931);
or UO_4701 (O_4701,N_49870,N_49925);
nand UO_4702 (O_4702,N_49537,N_49868);
nor UO_4703 (O_4703,N_49762,N_49558);
and UO_4704 (O_4704,N_49628,N_49711);
and UO_4705 (O_4705,N_49820,N_49943);
nand UO_4706 (O_4706,N_49911,N_49744);
and UO_4707 (O_4707,N_49862,N_49789);
nor UO_4708 (O_4708,N_49920,N_49704);
and UO_4709 (O_4709,N_49740,N_49594);
nand UO_4710 (O_4710,N_49813,N_49643);
and UO_4711 (O_4711,N_49962,N_49954);
xor UO_4712 (O_4712,N_49712,N_49685);
nor UO_4713 (O_4713,N_49992,N_49925);
and UO_4714 (O_4714,N_49678,N_49976);
and UO_4715 (O_4715,N_49656,N_49575);
nand UO_4716 (O_4716,N_49941,N_49852);
or UO_4717 (O_4717,N_49643,N_49601);
nand UO_4718 (O_4718,N_49874,N_49891);
xnor UO_4719 (O_4719,N_49801,N_49519);
nor UO_4720 (O_4720,N_49560,N_49705);
and UO_4721 (O_4721,N_49717,N_49712);
nor UO_4722 (O_4722,N_49897,N_49548);
nand UO_4723 (O_4723,N_49788,N_49982);
xor UO_4724 (O_4724,N_49922,N_49756);
or UO_4725 (O_4725,N_49627,N_49935);
or UO_4726 (O_4726,N_49826,N_49603);
or UO_4727 (O_4727,N_49678,N_49896);
nor UO_4728 (O_4728,N_49785,N_49942);
or UO_4729 (O_4729,N_49930,N_49850);
nand UO_4730 (O_4730,N_49660,N_49595);
and UO_4731 (O_4731,N_49778,N_49589);
xor UO_4732 (O_4732,N_49993,N_49999);
nand UO_4733 (O_4733,N_49502,N_49521);
and UO_4734 (O_4734,N_49849,N_49537);
nor UO_4735 (O_4735,N_49657,N_49984);
and UO_4736 (O_4736,N_49598,N_49628);
or UO_4737 (O_4737,N_49648,N_49978);
or UO_4738 (O_4738,N_49549,N_49561);
nor UO_4739 (O_4739,N_49801,N_49796);
nand UO_4740 (O_4740,N_49704,N_49963);
and UO_4741 (O_4741,N_49681,N_49742);
or UO_4742 (O_4742,N_49786,N_49632);
and UO_4743 (O_4743,N_49606,N_49525);
nor UO_4744 (O_4744,N_49645,N_49682);
nand UO_4745 (O_4745,N_49807,N_49556);
nand UO_4746 (O_4746,N_49917,N_49960);
nand UO_4747 (O_4747,N_49700,N_49843);
nand UO_4748 (O_4748,N_49675,N_49892);
or UO_4749 (O_4749,N_49755,N_49972);
nor UO_4750 (O_4750,N_49532,N_49975);
nor UO_4751 (O_4751,N_49849,N_49577);
and UO_4752 (O_4752,N_49982,N_49780);
and UO_4753 (O_4753,N_49647,N_49622);
nand UO_4754 (O_4754,N_49847,N_49853);
or UO_4755 (O_4755,N_49801,N_49837);
or UO_4756 (O_4756,N_49724,N_49568);
and UO_4757 (O_4757,N_49921,N_49728);
nand UO_4758 (O_4758,N_49975,N_49542);
xor UO_4759 (O_4759,N_49964,N_49590);
nor UO_4760 (O_4760,N_49772,N_49764);
nand UO_4761 (O_4761,N_49692,N_49511);
nor UO_4762 (O_4762,N_49520,N_49735);
and UO_4763 (O_4763,N_49791,N_49593);
and UO_4764 (O_4764,N_49982,N_49644);
and UO_4765 (O_4765,N_49566,N_49637);
nand UO_4766 (O_4766,N_49625,N_49933);
nand UO_4767 (O_4767,N_49881,N_49561);
nand UO_4768 (O_4768,N_49648,N_49515);
nand UO_4769 (O_4769,N_49565,N_49837);
xor UO_4770 (O_4770,N_49618,N_49825);
nor UO_4771 (O_4771,N_49517,N_49857);
and UO_4772 (O_4772,N_49983,N_49670);
nor UO_4773 (O_4773,N_49856,N_49620);
or UO_4774 (O_4774,N_49665,N_49826);
and UO_4775 (O_4775,N_49976,N_49820);
or UO_4776 (O_4776,N_49561,N_49513);
and UO_4777 (O_4777,N_49872,N_49808);
nor UO_4778 (O_4778,N_49550,N_49572);
or UO_4779 (O_4779,N_49784,N_49870);
nor UO_4780 (O_4780,N_49827,N_49642);
nor UO_4781 (O_4781,N_49620,N_49723);
xor UO_4782 (O_4782,N_49865,N_49827);
and UO_4783 (O_4783,N_49940,N_49534);
and UO_4784 (O_4784,N_49701,N_49541);
nand UO_4785 (O_4785,N_49633,N_49618);
nor UO_4786 (O_4786,N_49858,N_49983);
or UO_4787 (O_4787,N_49534,N_49688);
and UO_4788 (O_4788,N_49985,N_49831);
nor UO_4789 (O_4789,N_49738,N_49796);
and UO_4790 (O_4790,N_49962,N_49956);
nor UO_4791 (O_4791,N_49594,N_49825);
nor UO_4792 (O_4792,N_49542,N_49754);
or UO_4793 (O_4793,N_49920,N_49925);
or UO_4794 (O_4794,N_49971,N_49685);
nand UO_4795 (O_4795,N_49864,N_49658);
or UO_4796 (O_4796,N_49587,N_49840);
and UO_4797 (O_4797,N_49653,N_49782);
and UO_4798 (O_4798,N_49722,N_49889);
nor UO_4799 (O_4799,N_49616,N_49517);
nor UO_4800 (O_4800,N_49761,N_49902);
nand UO_4801 (O_4801,N_49580,N_49811);
or UO_4802 (O_4802,N_49811,N_49820);
or UO_4803 (O_4803,N_49708,N_49863);
nand UO_4804 (O_4804,N_49961,N_49981);
nand UO_4805 (O_4805,N_49667,N_49556);
and UO_4806 (O_4806,N_49740,N_49691);
nand UO_4807 (O_4807,N_49982,N_49765);
nor UO_4808 (O_4808,N_49963,N_49816);
nand UO_4809 (O_4809,N_49776,N_49938);
nand UO_4810 (O_4810,N_49639,N_49960);
nor UO_4811 (O_4811,N_49689,N_49882);
nand UO_4812 (O_4812,N_49885,N_49998);
or UO_4813 (O_4813,N_49799,N_49968);
nor UO_4814 (O_4814,N_49766,N_49517);
nor UO_4815 (O_4815,N_49832,N_49899);
nor UO_4816 (O_4816,N_49576,N_49638);
nor UO_4817 (O_4817,N_49836,N_49564);
nor UO_4818 (O_4818,N_49870,N_49926);
nand UO_4819 (O_4819,N_49908,N_49744);
or UO_4820 (O_4820,N_49549,N_49721);
and UO_4821 (O_4821,N_49500,N_49750);
and UO_4822 (O_4822,N_49793,N_49533);
and UO_4823 (O_4823,N_49677,N_49592);
nor UO_4824 (O_4824,N_49751,N_49511);
or UO_4825 (O_4825,N_49818,N_49657);
nor UO_4826 (O_4826,N_49931,N_49944);
or UO_4827 (O_4827,N_49682,N_49830);
nor UO_4828 (O_4828,N_49620,N_49630);
or UO_4829 (O_4829,N_49670,N_49821);
nand UO_4830 (O_4830,N_49867,N_49564);
and UO_4831 (O_4831,N_49527,N_49803);
nand UO_4832 (O_4832,N_49893,N_49598);
nor UO_4833 (O_4833,N_49835,N_49939);
or UO_4834 (O_4834,N_49714,N_49931);
nand UO_4835 (O_4835,N_49946,N_49913);
and UO_4836 (O_4836,N_49644,N_49724);
and UO_4837 (O_4837,N_49656,N_49686);
nor UO_4838 (O_4838,N_49516,N_49515);
and UO_4839 (O_4839,N_49905,N_49901);
xnor UO_4840 (O_4840,N_49724,N_49609);
and UO_4841 (O_4841,N_49710,N_49892);
or UO_4842 (O_4842,N_49996,N_49890);
and UO_4843 (O_4843,N_49792,N_49911);
nand UO_4844 (O_4844,N_49532,N_49789);
nor UO_4845 (O_4845,N_49534,N_49798);
xnor UO_4846 (O_4846,N_49579,N_49740);
or UO_4847 (O_4847,N_49590,N_49634);
or UO_4848 (O_4848,N_49885,N_49812);
or UO_4849 (O_4849,N_49543,N_49780);
and UO_4850 (O_4850,N_49826,N_49932);
or UO_4851 (O_4851,N_49555,N_49862);
and UO_4852 (O_4852,N_49615,N_49537);
and UO_4853 (O_4853,N_49651,N_49680);
nand UO_4854 (O_4854,N_49782,N_49602);
and UO_4855 (O_4855,N_49535,N_49749);
nand UO_4856 (O_4856,N_49979,N_49742);
nand UO_4857 (O_4857,N_49596,N_49533);
or UO_4858 (O_4858,N_49596,N_49810);
and UO_4859 (O_4859,N_49884,N_49706);
or UO_4860 (O_4860,N_49760,N_49613);
nor UO_4861 (O_4861,N_49955,N_49676);
nor UO_4862 (O_4862,N_49669,N_49996);
nand UO_4863 (O_4863,N_49587,N_49567);
and UO_4864 (O_4864,N_49505,N_49831);
nor UO_4865 (O_4865,N_49901,N_49962);
and UO_4866 (O_4866,N_49715,N_49679);
xor UO_4867 (O_4867,N_49774,N_49718);
nor UO_4868 (O_4868,N_49516,N_49534);
and UO_4869 (O_4869,N_49982,N_49889);
xor UO_4870 (O_4870,N_49745,N_49671);
nor UO_4871 (O_4871,N_49958,N_49772);
nand UO_4872 (O_4872,N_49535,N_49710);
nand UO_4873 (O_4873,N_49650,N_49673);
nand UO_4874 (O_4874,N_49539,N_49633);
and UO_4875 (O_4875,N_49700,N_49528);
nand UO_4876 (O_4876,N_49613,N_49900);
or UO_4877 (O_4877,N_49923,N_49925);
or UO_4878 (O_4878,N_49661,N_49707);
or UO_4879 (O_4879,N_49542,N_49921);
and UO_4880 (O_4880,N_49710,N_49732);
nand UO_4881 (O_4881,N_49685,N_49943);
nand UO_4882 (O_4882,N_49621,N_49995);
nand UO_4883 (O_4883,N_49791,N_49769);
nand UO_4884 (O_4884,N_49775,N_49746);
nand UO_4885 (O_4885,N_49711,N_49590);
and UO_4886 (O_4886,N_49836,N_49780);
or UO_4887 (O_4887,N_49959,N_49513);
or UO_4888 (O_4888,N_49993,N_49878);
nand UO_4889 (O_4889,N_49573,N_49801);
xor UO_4890 (O_4890,N_49694,N_49981);
or UO_4891 (O_4891,N_49908,N_49843);
or UO_4892 (O_4892,N_49684,N_49512);
xnor UO_4893 (O_4893,N_49683,N_49734);
nand UO_4894 (O_4894,N_49684,N_49811);
and UO_4895 (O_4895,N_49611,N_49619);
and UO_4896 (O_4896,N_49899,N_49535);
and UO_4897 (O_4897,N_49743,N_49866);
or UO_4898 (O_4898,N_49536,N_49731);
nand UO_4899 (O_4899,N_49996,N_49523);
and UO_4900 (O_4900,N_49518,N_49546);
nor UO_4901 (O_4901,N_49676,N_49636);
or UO_4902 (O_4902,N_49744,N_49735);
nor UO_4903 (O_4903,N_49869,N_49929);
and UO_4904 (O_4904,N_49891,N_49731);
and UO_4905 (O_4905,N_49502,N_49595);
xor UO_4906 (O_4906,N_49848,N_49745);
nand UO_4907 (O_4907,N_49534,N_49938);
nand UO_4908 (O_4908,N_49921,N_49796);
nand UO_4909 (O_4909,N_49548,N_49739);
and UO_4910 (O_4910,N_49630,N_49694);
xnor UO_4911 (O_4911,N_49728,N_49839);
or UO_4912 (O_4912,N_49536,N_49649);
and UO_4913 (O_4913,N_49772,N_49705);
nand UO_4914 (O_4914,N_49904,N_49501);
or UO_4915 (O_4915,N_49903,N_49604);
or UO_4916 (O_4916,N_49849,N_49729);
nor UO_4917 (O_4917,N_49618,N_49560);
or UO_4918 (O_4918,N_49987,N_49737);
or UO_4919 (O_4919,N_49975,N_49850);
and UO_4920 (O_4920,N_49618,N_49924);
nand UO_4921 (O_4921,N_49541,N_49721);
or UO_4922 (O_4922,N_49702,N_49676);
nand UO_4923 (O_4923,N_49906,N_49799);
and UO_4924 (O_4924,N_49765,N_49603);
xnor UO_4925 (O_4925,N_49654,N_49701);
or UO_4926 (O_4926,N_49697,N_49903);
nor UO_4927 (O_4927,N_49910,N_49884);
nand UO_4928 (O_4928,N_49588,N_49747);
xnor UO_4929 (O_4929,N_49718,N_49972);
xor UO_4930 (O_4930,N_49772,N_49937);
nor UO_4931 (O_4931,N_49945,N_49949);
or UO_4932 (O_4932,N_49740,N_49861);
and UO_4933 (O_4933,N_49591,N_49901);
nor UO_4934 (O_4934,N_49844,N_49642);
xor UO_4935 (O_4935,N_49967,N_49686);
or UO_4936 (O_4936,N_49828,N_49979);
nor UO_4937 (O_4937,N_49816,N_49772);
nor UO_4938 (O_4938,N_49658,N_49784);
nand UO_4939 (O_4939,N_49509,N_49684);
nor UO_4940 (O_4940,N_49931,N_49975);
or UO_4941 (O_4941,N_49733,N_49908);
nand UO_4942 (O_4942,N_49635,N_49876);
or UO_4943 (O_4943,N_49878,N_49676);
nor UO_4944 (O_4944,N_49542,N_49667);
nand UO_4945 (O_4945,N_49757,N_49596);
nor UO_4946 (O_4946,N_49721,N_49506);
or UO_4947 (O_4947,N_49541,N_49503);
xor UO_4948 (O_4948,N_49864,N_49983);
nor UO_4949 (O_4949,N_49646,N_49795);
and UO_4950 (O_4950,N_49550,N_49988);
xnor UO_4951 (O_4951,N_49615,N_49630);
or UO_4952 (O_4952,N_49787,N_49753);
nand UO_4953 (O_4953,N_49830,N_49904);
nor UO_4954 (O_4954,N_49875,N_49907);
and UO_4955 (O_4955,N_49619,N_49590);
nand UO_4956 (O_4956,N_49584,N_49644);
nand UO_4957 (O_4957,N_49861,N_49975);
or UO_4958 (O_4958,N_49769,N_49835);
xor UO_4959 (O_4959,N_49563,N_49884);
nor UO_4960 (O_4960,N_49661,N_49931);
or UO_4961 (O_4961,N_49600,N_49614);
and UO_4962 (O_4962,N_49834,N_49505);
nor UO_4963 (O_4963,N_49940,N_49736);
or UO_4964 (O_4964,N_49725,N_49973);
nor UO_4965 (O_4965,N_49921,N_49957);
nand UO_4966 (O_4966,N_49945,N_49763);
and UO_4967 (O_4967,N_49523,N_49669);
or UO_4968 (O_4968,N_49816,N_49614);
and UO_4969 (O_4969,N_49720,N_49689);
or UO_4970 (O_4970,N_49846,N_49998);
nand UO_4971 (O_4971,N_49911,N_49614);
or UO_4972 (O_4972,N_49862,N_49554);
nor UO_4973 (O_4973,N_49902,N_49559);
and UO_4974 (O_4974,N_49999,N_49791);
nand UO_4975 (O_4975,N_49646,N_49637);
or UO_4976 (O_4976,N_49825,N_49942);
or UO_4977 (O_4977,N_49918,N_49606);
nor UO_4978 (O_4978,N_49724,N_49570);
and UO_4979 (O_4979,N_49759,N_49961);
and UO_4980 (O_4980,N_49970,N_49606);
nor UO_4981 (O_4981,N_49821,N_49519);
nand UO_4982 (O_4982,N_49761,N_49716);
nor UO_4983 (O_4983,N_49643,N_49577);
and UO_4984 (O_4984,N_49794,N_49574);
or UO_4985 (O_4985,N_49679,N_49934);
nand UO_4986 (O_4986,N_49971,N_49869);
nor UO_4987 (O_4987,N_49933,N_49607);
nor UO_4988 (O_4988,N_49688,N_49521);
nand UO_4989 (O_4989,N_49881,N_49577);
nor UO_4990 (O_4990,N_49773,N_49837);
and UO_4991 (O_4991,N_49858,N_49598);
nor UO_4992 (O_4992,N_49784,N_49819);
nand UO_4993 (O_4993,N_49525,N_49918);
nand UO_4994 (O_4994,N_49653,N_49676);
or UO_4995 (O_4995,N_49978,N_49553);
xnor UO_4996 (O_4996,N_49755,N_49644);
nand UO_4997 (O_4997,N_49834,N_49546);
and UO_4998 (O_4998,N_49743,N_49970);
nand UO_4999 (O_4999,N_49654,N_49743);
endmodule