module basic_1500_15000_2000_120_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_402,In_1220);
or U1 (N_1,In_120,In_168);
nor U2 (N_2,In_1192,In_740);
and U3 (N_3,In_1404,In_1265);
or U4 (N_4,In_279,In_735);
xnor U5 (N_5,In_1084,In_796);
or U6 (N_6,In_1390,In_963);
or U7 (N_7,In_603,In_1438);
nor U8 (N_8,In_378,In_868);
nor U9 (N_9,In_344,In_571);
or U10 (N_10,In_232,In_561);
or U11 (N_11,In_53,In_725);
or U12 (N_12,In_1454,In_58);
xnor U13 (N_13,In_1450,In_1446);
xor U14 (N_14,In_55,In_543);
or U15 (N_15,In_913,In_658);
xnor U16 (N_16,In_493,In_1180);
xnor U17 (N_17,In_395,In_1392);
xor U18 (N_18,In_1149,In_1313);
or U19 (N_19,In_770,In_905);
nor U20 (N_20,In_1421,In_252);
nand U21 (N_21,In_159,In_529);
nor U22 (N_22,In_429,In_1455);
xnor U23 (N_23,In_726,In_939);
nand U24 (N_24,In_0,In_472);
xnor U25 (N_25,In_455,In_910);
and U26 (N_26,In_1197,In_68);
nor U27 (N_27,In_1399,In_565);
xor U28 (N_28,In_1221,In_592);
or U29 (N_29,In_1321,In_164);
nor U30 (N_30,In_986,In_652);
and U31 (N_31,In_14,In_234);
and U32 (N_32,In_1267,In_530);
nand U33 (N_33,In_1495,In_508);
and U34 (N_34,In_433,In_778);
nand U35 (N_35,In_1338,In_32);
or U36 (N_36,In_266,In_1339);
nand U37 (N_37,In_144,In_1484);
xnor U38 (N_38,In_886,In_676);
nor U39 (N_39,In_497,In_1199);
nor U40 (N_40,In_115,In_121);
nand U41 (N_41,In_909,In_817);
nand U42 (N_42,In_462,In_1058);
nor U43 (N_43,In_889,In_31);
xor U44 (N_44,In_44,In_798);
and U45 (N_45,In_668,In_1116);
nand U46 (N_46,In_81,In_265);
nor U47 (N_47,In_1427,In_1017);
xor U48 (N_48,In_774,In_339);
and U49 (N_49,In_945,In_687);
nand U50 (N_50,In_517,In_789);
nand U51 (N_51,In_439,In_628);
and U52 (N_52,In_1452,In_1329);
xor U53 (N_53,In_1053,In_1070);
and U54 (N_54,In_1039,In_1066);
and U55 (N_55,In_1309,In_299);
nor U56 (N_56,In_1198,In_793);
and U57 (N_57,In_843,In_42);
nor U58 (N_58,In_406,In_548);
or U59 (N_59,In_539,In_442);
and U60 (N_60,In_270,In_1021);
and U61 (N_61,In_468,In_469);
and U62 (N_62,In_61,In_657);
xnor U63 (N_63,In_825,In_610);
xor U64 (N_64,In_874,In_692);
nor U65 (N_65,In_632,In_209);
or U66 (N_66,In_346,In_284);
or U67 (N_67,In_1469,In_471);
xor U68 (N_68,In_615,In_716);
and U69 (N_69,In_29,In_1237);
nor U70 (N_70,In_764,In_1317);
nor U71 (N_71,In_1476,In_875);
and U72 (N_72,In_408,In_1101);
and U73 (N_73,In_570,In_136);
or U74 (N_74,In_487,In_664);
xor U75 (N_75,In_695,In_227);
or U76 (N_76,In_576,In_1184);
and U77 (N_77,In_180,In_37);
nand U78 (N_78,In_634,In_73);
xnor U79 (N_79,In_907,In_1445);
nand U80 (N_80,In_1023,In_291);
nand U81 (N_81,In_1418,In_1249);
nor U82 (N_82,In_217,In_1076);
nand U83 (N_83,In_641,In_1359);
nand U84 (N_84,In_72,In_544);
and U85 (N_85,In_1323,In_48);
or U86 (N_86,In_512,In_940);
or U87 (N_87,In_1134,In_88);
nor U88 (N_88,In_86,In_853);
nand U89 (N_89,In_1040,In_122);
nor U90 (N_90,In_294,In_505);
and U91 (N_91,In_998,In_391);
nand U92 (N_92,In_1242,In_877);
or U93 (N_93,In_1414,In_1081);
nor U94 (N_94,In_354,In_308);
xnor U95 (N_95,In_590,In_744);
nor U96 (N_96,In_1379,In_239);
nor U97 (N_97,In_1448,In_204);
and U98 (N_98,In_1335,In_928);
or U99 (N_99,In_852,In_409);
and U100 (N_100,In_763,In_810);
and U101 (N_101,In_1316,In_331);
or U102 (N_102,In_146,In_297);
nand U103 (N_103,In_1124,In_161);
and U104 (N_104,In_167,In_1229);
or U105 (N_105,In_1481,In_151);
nand U106 (N_106,In_1201,In_1370);
nor U107 (N_107,In_779,In_523);
xor U108 (N_108,In_401,In_50);
or U109 (N_109,In_4,In_23);
or U110 (N_110,In_950,In_1104);
nand U111 (N_111,In_1422,In_683);
xnor U112 (N_112,In_654,In_385);
and U113 (N_113,In_559,In_1274);
or U114 (N_114,In_1496,In_693);
xnor U115 (N_115,In_1402,In_797);
nand U116 (N_116,In_959,In_972);
xor U117 (N_117,In_682,In_524);
xnor U118 (N_118,In_1380,In_644);
and U119 (N_119,In_241,In_1016);
nor U120 (N_120,In_436,In_896);
xor U121 (N_121,In_35,In_225);
and U122 (N_122,In_991,In_719);
xnor U123 (N_123,In_375,In_430);
nor U124 (N_124,In_390,In_1491);
xnor U125 (N_125,In_1156,N_110);
and U126 (N_126,In_783,In_330);
or U127 (N_127,In_1408,In_606);
nand U128 (N_128,N_40,In_101);
nand U129 (N_129,In_662,In_410);
xor U130 (N_130,N_93,In_193);
and U131 (N_131,In_1305,In_12);
nand U132 (N_132,In_13,In_938);
nand U133 (N_133,In_1352,In_1123);
nor U134 (N_134,In_1085,In_513);
xnor U135 (N_135,In_511,N_62);
and U136 (N_136,In_202,In_1291);
xor U137 (N_137,N_65,In_1003);
or U138 (N_138,In_1294,In_148);
and U139 (N_139,In_105,In_816);
and U140 (N_140,In_510,In_1031);
nor U141 (N_141,In_1474,In_1119);
xor U142 (N_142,In_317,In_835);
or U143 (N_143,In_884,In_699);
and U144 (N_144,In_1374,In_1262);
nand U145 (N_145,In_1145,In_944);
or U146 (N_146,In_1138,In_251);
or U147 (N_147,In_475,In_153);
xor U148 (N_148,In_1458,In_737);
and U149 (N_149,In_1412,In_960);
xnor U150 (N_150,N_54,In_1312);
nor U151 (N_151,N_47,In_132);
or U152 (N_152,N_97,In_451);
nor U153 (N_153,In_675,In_200);
xor U154 (N_154,In_679,In_1463);
or U155 (N_155,In_1257,In_271);
and U156 (N_156,N_23,In_152);
or U157 (N_157,In_946,In_1396);
xor U158 (N_158,In_996,In_280);
or U159 (N_159,In_1147,In_482);
nor U160 (N_160,In_1459,In_1336);
or U161 (N_161,In_876,In_382);
nand U162 (N_162,In_1494,In_374);
nand U163 (N_163,In_748,In_210);
nand U164 (N_164,In_326,In_1461);
xor U165 (N_165,In_33,In_1343);
or U166 (N_166,In_1144,In_1132);
nor U167 (N_167,In_1034,In_1099);
nor U168 (N_168,In_399,In_678);
xor U169 (N_169,In_869,In_1363);
or U170 (N_170,In_655,In_597);
nand U171 (N_171,In_1401,In_1310);
and U172 (N_172,In_614,In_553);
nand U173 (N_173,In_752,In_1243);
and U174 (N_174,N_16,In_163);
xnor U175 (N_175,In_1111,In_1178);
xnor U176 (N_176,In_671,N_33);
nor U177 (N_177,In_864,In_760);
or U178 (N_178,In_862,In_1430);
or U179 (N_179,In_900,In_1383);
nand U180 (N_180,In_1087,N_75);
or U181 (N_181,In_428,In_1239);
xor U182 (N_182,In_1286,In_638);
nand U183 (N_183,In_1497,N_123);
nand U184 (N_184,In_912,In_139);
and U185 (N_185,In_674,In_228);
or U186 (N_186,In_355,N_8);
or U187 (N_187,In_198,In_393);
and U188 (N_188,In_775,In_926);
or U189 (N_189,In_1473,In_995);
nor U190 (N_190,In_785,In_1037);
nor U191 (N_191,In_484,In_310);
or U192 (N_192,In_1029,In_1096);
xnor U193 (N_193,In_306,In_64);
or U194 (N_194,N_98,In_1032);
xor U195 (N_195,In_286,In_1424);
and U196 (N_196,In_973,In_882);
and U197 (N_197,In_214,In_992);
xor U198 (N_198,N_43,In_231);
nor U199 (N_199,In_1432,In_935);
and U200 (N_200,In_1389,In_1036);
nand U201 (N_201,In_1167,In_1079);
and U202 (N_202,In_460,In_84);
nor U203 (N_203,In_863,In_437);
and U204 (N_204,In_1193,In_457);
nand U205 (N_205,In_259,In_1045);
and U206 (N_206,In_715,In_477);
and U207 (N_207,N_105,In_203);
nand U208 (N_208,In_696,In_1028);
nor U209 (N_209,In_1183,In_933);
nand U210 (N_210,In_870,In_697);
nand U211 (N_211,In_318,In_28);
xor U212 (N_212,In_269,In_818);
xnor U213 (N_213,In_463,In_514);
and U214 (N_214,In_1207,In_961);
xor U215 (N_215,In_1170,In_507);
nand U216 (N_216,In_9,In_1314);
xnor U217 (N_217,In_397,In_751);
nand U218 (N_218,In_1010,In_3);
xnor U219 (N_219,In_1030,In_822);
xor U220 (N_220,In_780,In_1210);
and U221 (N_221,In_413,In_966);
xnor U222 (N_222,In_328,In_921);
or U223 (N_223,In_185,In_129);
xor U224 (N_224,In_552,In_694);
xor U225 (N_225,In_18,In_1453);
and U226 (N_226,In_283,N_57);
nand U227 (N_227,In_157,In_516);
or U228 (N_228,N_21,In_786);
nand U229 (N_229,In_823,In_22);
xor U230 (N_230,In_617,In_1102);
nor U231 (N_231,In_322,In_242);
nand U232 (N_232,In_901,In_1175);
and U233 (N_233,In_1152,In_1261);
nand U234 (N_234,In_356,In_1200);
or U235 (N_235,In_222,In_1054);
nand U236 (N_236,In_769,In_381);
and U237 (N_237,In_321,In_916);
or U238 (N_238,In_724,In_1130);
and U239 (N_239,In_1011,N_26);
nand U240 (N_240,In_1333,In_677);
nand U241 (N_241,In_476,In_112);
xnor U242 (N_242,In_1282,N_51);
xnor U243 (N_243,In_248,In_108);
and U244 (N_244,N_115,In_1121);
and U245 (N_245,N_42,In_738);
xor U246 (N_246,In_1415,In_1384);
and U247 (N_247,In_894,In_551);
nand U248 (N_248,In_196,In_5);
and U249 (N_249,In_432,In_1002);
nor U250 (N_250,In_1351,In_262);
nand U251 (N_251,In_589,In_661);
xnor U252 (N_252,N_59,In_1120);
or U253 (N_253,In_659,In_1241);
xnor U254 (N_254,In_1108,In_371);
nand U255 (N_255,In_534,In_799);
or U256 (N_256,In_1187,In_838);
and U257 (N_257,In_282,N_240);
xor U258 (N_258,In_880,In_1442);
xor U259 (N_259,In_421,In_93);
and U260 (N_260,In_1234,In_837);
nor U261 (N_261,N_209,N_11);
xor U262 (N_262,In_1209,In_71);
nand U263 (N_263,N_91,In_701);
or U264 (N_264,In_518,In_117);
nand U265 (N_265,In_1354,N_134);
nand U266 (N_266,In_856,In_611);
nand U267 (N_267,In_80,In_246);
and U268 (N_268,In_965,In_1001);
xnor U269 (N_269,In_212,In_1434);
xnor U270 (N_270,In_135,In_700);
xnor U271 (N_271,In_70,In_1441);
or U272 (N_272,In_1324,In_1067);
or U273 (N_273,N_10,N_30);
nand U274 (N_274,In_345,N_28);
xor U275 (N_275,In_370,In_118);
xnor U276 (N_276,N_1,N_76);
nor U277 (N_277,In_581,N_154);
nor U278 (N_278,In_647,In_1208);
or U279 (N_279,N_215,In_8);
and U280 (N_280,In_461,In_1340);
nor U281 (N_281,N_73,In_133);
xor U282 (N_282,In_178,In_94);
nand U283 (N_283,In_1465,In_541);
or U284 (N_284,In_602,In_215);
xnor U285 (N_285,In_969,In_1378);
and U286 (N_286,N_182,In_1191);
xor U287 (N_287,In_979,In_240);
and U288 (N_288,In_444,In_929);
xor U289 (N_289,In_688,N_143);
and U290 (N_290,N_46,In_1107);
or U291 (N_291,In_1381,In_1413);
or U292 (N_292,N_13,In_1044);
and U293 (N_293,In_337,In_82);
xor U294 (N_294,In_622,In_566);
and U295 (N_295,In_263,In_1077);
nand U296 (N_296,In_1217,N_173);
or U297 (N_297,In_1190,In_1482);
nor U298 (N_298,N_41,In_555);
or U299 (N_299,In_126,In_314);
or U300 (N_300,In_383,In_845);
or U301 (N_301,In_947,In_1177);
xor U302 (N_302,In_40,In_298);
xnor U303 (N_303,In_1472,In_578);
nor U304 (N_304,In_782,In_10);
xor U305 (N_305,In_464,In_1375);
and U306 (N_306,In_968,In_450);
and U307 (N_307,N_223,N_197);
xnor U308 (N_308,In_333,In_1431);
and U309 (N_309,In_181,In_558);
and U310 (N_310,In_1105,N_245);
and U311 (N_311,N_6,In_1281);
and U312 (N_312,In_1136,In_1326);
or U313 (N_313,In_1385,N_172);
and U314 (N_314,In_1376,In_188);
nand U315 (N_315,In_645,In_373);
or U316 (N_316,In_443,In_633);
xnor U317 (N_317,N_177,In_1462);
nor U318 (N_318,In_1174,In_1301);
xor U319 (N_319,N_121,In_1290);
nor U320 (N_320,In_130,In_836);
and U321 (N_321,In_1033,In_557);
or U322 (N_322,In_987,N_88);
nor U323 (N_323,In_540,In_1179);
or U324 (N_324,In_651,In_596);
nor U325 (N_325,In_709,In_224);
or U326 (N_326,N_35,N_52);
nor U327 (N_327,N_192,In_1127);
or U328 (N_328,In_712,In_142);
or U329 (N_329,In_860,In_943);
or U330 (N_330,N_132,N_141);
nand U331 (N_331,In_7,In_771);
nor U332 (N_332,In_1219,N_191);
nor U333 (N_333,In_208,N_229);
and U334 (N_334,In_1006,N_167);
xor U335 (N_335,In_504,In_1288);
nand U336 (N_336,In_1150,In_59);
and U337 (N_337,N_210,In_140);
nor U338 (N_338,N_69,In_446);
or U339 (N_339,N_225,N_179);
nor U340 (N_340,In_1371,In_902);
and U341 (N_341,In_245,In_1012);
and U342 (N_342,In_743,N_239);
and U343 (N_343,In_1449,In_640);
nand U344 (N_344,In_149,In_1059);
nor U345 (N_345,In_1244,N_189);
xor U346 (N_346,In_533,N_20);
or U347 (N_347,In_1364,In_1303);
nor U348 (N_348,In_1162,In_171);
or U349 (N_349,In_325,In_273);
and U350 (N_350,N_87,In_422);
xnor U351 (N_351,In_1306,In_795);
xor U352 (N_352,In_1360,In_601);
or U353 (N_353,In_859,In_1141);
or U354 (N_354,In_1485,In_1166);
nand U355 (N_355,In_827,In_123);
and U356 (N_356,N_102,N_44);
or U357 (N_357,In_904,N_126);
and U358 (N_358,In_1230,In_277);
nor U359 (N_359,In_119,In_1366);
and U360 (N_360,In_1318,In_978);
and U361 (N_361,In_911,N_144);
and U362 (N_362,In_285,In_941);
and U363 (N_363,In_1487,In_45);
or U364 (N_364,In_705,N_185);
or U365 (N_365,In_172,In_791);
or U366 (N_366,In_293,In_792);
nand U367 (N_367,In_1470,In_295);
nand U368 (N_368,In_841,In_808);
xor U369 (N_369,In_6,N_63);
nand U370 (N_370,In_43,In_1428);
xnor U371 (N_371,In_1315,In_630);
or U372 (N_372,N_222,N_146);
or U373 (N_373,In_1135,In_249);
and U374 (N_374,In_582,N_0);
nor U375 (N_375,In_957,In_1035);
nand U376 (N_376,In_109,In_1074);
or U377 (N_377,In_915,In_494);
and U378 (N_378,N_249,In_386);
nor U379 (N_379,In_583,In_1355);
or U380 (N_380,In_499,In_828);
xor U381 (N_381,In_1328,In_1086);
or U382 (N_382,In_106,N_366);
nor U383 (N_383,In_1222,In_25);
nand U384 (N_384,In_1092,In_352);
or U385 (N_385,In_515,N_293);
nand U386 (N_386,In_319,N_118);
nand U387 (N_387,In_648,In_1475);
xnor U388 (N_388,N_31,In_689);
or U389 (N_389,In_964,In_492);
xor U390 (N_390,In_440,In_528);
or U391 (N_391,N_17,In_447);
nand U392 (N_392,In_1477,In_1499);
xnor U393 (N_393,In_951,In_250);
or U394 (N_394,N_295,In_936);
and U395 (N_395,N_176,In_414);
nor U396 (N_396,In_895,N_324);
nand U397 (N_397,In_1420,In_1115);
xor U398 (N_398,In_448,In_1275);
nand U399 (N_399,In_980,In_729);
xnor U400 (N_400,In_1195,In_595);
or U401 (N_401,In_521,In_179);
nor U402 (N_402,In_1240,In_806);
nor U403 (N_403,In_1387,N_272);
nand U404 (N_404,In_1047,In_348);
xnor U405 (N_405,N_86,In_643);
or U406 (N_406,In_727,N_243);
xor U407 (N_407,In_1005,In_1214);
nor U408 (N_408,In_650,N_319);
nor U409 (N_409,In_1483,In_335);
or U410 (N_410,In_878,In_1272);
or U411 (N_411,In_1069,In_958);
or U412 (N_412,N_290,In_1196);
xor U413 (N_413,In_237,In_722);
nand U414 (N_414,In_102,N_32);
nand U415 (N_415,In_830,In_759);
nand U416 (N_416,N_165,N_234);
xnor U417 (N_417,N_37,N_287);
nor U418 (N_418,In_1013,In_1346);
or U419 (N_419,N_255,In_253);
nand U420 (N_420,N_163,In_1299);
nor U421 (N_421,In_1304,In_1046);
and U422 (N_422,In_754,In_1228);
xnor U423 (N_423,In_1330,In_997);
and U424 (N_424,N_55,In_1276);
nor U425 (N_425,N_304,In_1122);
nand U426 (N_426,N_276,In_1489);
or U427 (N_427,In_788,N_230);
nand U428 (N_428,In_934,In_1161);
and U429 (N_429,N_340,N_7);
nand U430 (N_430,In_1114,N_262);
or U431 (N_431,In_994,N_212);
or U432 (N_432,N_95,N_36);
nor U433 (N_433,In_1419,In_599);
nor U434 (N_434,N_345,N_312);
xnor U435 (N_435,In_124,In_924);
xnor U436 (N_436,In_431,N_314);
nor U437 (N_437,In_1246,In_1320);
nor U438 (N_438,N_248,In_1041);
nor U439 (N_439,In_197,In_720);
xnor U440 (N_440,In_999,In_625);
xor U441 (N_441,In_223,In_1368);
xnor U442 (N_442,In_635,In_459);
xor U443 (N_443,N_186,In_1373);
and U444 (N_444,In_920,In_1008);
nor U445 (N_445,In_1165,N_27);
xor U446 (N_446,N_15,In_89);
xnor U447 (N_447,In_873,In_594);
or U448 (N_448,In_623,In_47);
and U449 (N_449,N_283,N_347);
nand U450 (N_450,In_1279,In_988);
xnor U451 (N_451,In_195,In_731);
xnor U452 (N_452,In_488,N_260);
nand U453 (N_453,N_374,In_160);
nand U454 (N_454,In_26,In_1160);
nand U455 (N_455,N_2,In_932);
nor U456 (N_456,In_569,In_456);
and U457 (N_457,In_174,In_11);
or U458 (N_458,In_1284,N_193);
nor U459 (N_459,In_1055,In_732);
nand U460 (N_460,In_736,In_772);
nand U461 (N_461,In_537,N_19);
nor U462 (N_462,In_1334,In_62);
and U463 (N_463,N_246,In_226);
or U464 (N_464,In_1259,In_1159);
nand U465 (N_465,N_352,N_351);
nand U466 (N_466,N_96,In_340);
nor U467 (N_467,N_217,N_247);
xnor U468 (N_468,In_304,In_267);
and U469 (N_469,In_98,In_560);
xnor U470 (N_470,In_1194,In_170);
nor U471 (N_471,In_794,N_257);
and U472 (N_472,In_368,N_251);
or U473 (N_473,In_1403,N_218);
nor U474 (N_474,In_741,In_1268);
or U475 (N_475,In_1164,In_1226);
xor U476 (N_476,N_301,In_821);
or U477 (N_477,N_78,In_211);
and U478 (N_478,In_307,In_626);
nor U479 (N_479,In_434,In_24);
xor U480 (N_480,N_306,In_379);
nand U481 (N_481,In_556,N_81);
nand U482 (N_482,N_135,N_64);
nor U483 (N_483,In_357,N_359);
nor U484 (N_484,N_104,N_256);
nand U485 (N_485,In_254,In_1043);
or U486 (N_486,In_1235,In_1218);
or U487 (N_487,In_186,N_72);
xor U488 (N_488,In_685,N_68);
and U489 (N_489,In_189,In_914);
and U490 (N_490,In_1142,N_151);
xnor U491 (N_491,In_1157,In_1100);
and U492 (N_492,In_51,In_233);
nand U493 (N_493,In_85,N_241);
nand U494 (N_494,In_207,In_1245);
xnor U495 (N_495,In_927,In_338);
nor U496 (N_496,N_137,In_49);
nor U497 (N_497,In_820,In_642);
or U498 (N_498,In_315,In_1163);
xnor U499 (N_499,In_76,In_329);
or U500 (N_500,In_649,In_1258);
or U501 (N_501,N_449,In_812);
nand U502 (N_502,In_467,N_432);
xor U503 (N_503,In_1133,In_1498);
and U504 (N_504,In_1250,N_318);
nand U505 (N_505,N_82,N_269);
or U506 (N_506,In_1395,In_264);
nand U507 (N_507,In_69,In_888);
nand U508 (N_508,N_461,N_420);
xnor U509 (N_509,N_349,In_288);
or U510 (N_510,In_804,In_39);
nor U511 (N_511,N_194,In_438);
or U512 (N_512,N_213,N_440);
nand U513 (N_513,In_1050,In_74);
or U514 (N_514,In_535,N_360);
nand U515 (N_515,In_656,N_411);
nand U516 (N_516,N_363,In_971);
xnor U517 (N_517,In_1146,N_430);
nand U518 (N_518,In_478,In_470);
nand U519 (N_519,In_527,In_176);
nand U520 (N_520,N_297,N_308);
or U521 (N_521,In_1327,N_353);
nor U522 (N_522,In_525,In_1325);
nand U523 (N_523,N_448,N_214);
and U524 (N_524,In_272,In_155);
and U525 (N_525,In_1263,In_34);
or U526 (N_526,N_168,In_351);
xor U527 (N_527,N_117,N_221);
or U528 (N_528,In_1407,In_1398);
and U529 (N_529,N_83,In_781);
xor U530 (N_530,In_116,In_750);
nor U531 (N_531,In_454,In_952);
xor U532 (N_532,N_207,In_1185);
and U533 (N_533,N_25,In_1007);
nor U534 (N_534,In_403,In_268);
and U535 (N_535,In_545,In_347);
and U536 (N_536,In_205,In_496);
nand U537 (N_537,In_1068,N_331);
nand U538 (N_538,In_491,N_368);
and U539 (N_539,In_187,In_1131);
xnor U540 (N_540,N_317,In_1022);
and U541 (N_541,In_396,In_369);
or U542 (N_542,In_303,N_142);
or U543 (N_543,In_665,N_485);
nor U544 (N_544,In_542,N_433);
nand U545 (N_545,N_183,In_201);
nor U546 (N_546,N_170,N_196);
nor U547 (N_547,In_360,In_698);
nand U548 (N_548,In_423,In_890);
xor U549 (N_549,N_358,In_567);
nand U550 (N_550,N_323,N_22);
nor U551 (N_551,In_849,In_1298);
and U552 (N_552,In_1154,In_605);
and U553 (N_553,N_275,N_128);
or U554 (N_554,In_417,N_289);
nand U555 (N_555,N_258,In_1173);
xor U556 (N_556,In_733,In_532);
and U557 (N_557,In_128,N_468);
or U558 (N_558,In_1176,N_79);
nand U559 (N_559,In_1270,In_1451);
xnor U560 (N_560,In_653,N_300);
xnor U561 (N_561,In_681,In_1302);
and U562 (N_562,In_1433,In_871);
nand U563 (N_563,In_296,In_831);
and U564 (N_564,In_776,In_256);
nand U565 (N_565,In_127,In_962);
and U566 (N_566,In_302,In_1297);
xnor U567 (N_567,N_242,In_365);
and U568 (N_568,In_1143,In_145);
or U569 (N_569,In_826,N_92);
and U570 (N_570,N_111,In_1106);
and U571 (N_571,In_1285,In_803);
and U572 (N_572,In_908,N_108);
nor U573 (N_573,In_1295,N_268);
nand U574 (N_574,N_472,N_282);
xor U575 (N_575,N_475,N_467);
and U576 (N_576,In_289,In_485);
or U577 (N_577,N_107,In_536);
xor U578 (N_578,In_313,In_353);
or U579 (N_579,In_261,In_96);
or U580 (N_580,N_206,In_844);
nor U581 (N_581,N_327,In_99);
and U582 (N_582,In_538,N_56);
and U583 (N_583,N_428,In_608);
nand U584 (N_584,In_1203,In_1361);
nor U585 (N_585,N_338,N_61);
or U586 (N_586,In_183,In_1493);
or U587 (N_587,N_50,N_49);
nor U588 (N_588,In_19,N_479);
nand U589 (N_589,In_480,N_288);
nand U590 (N_590,N_178,In_1051);
and U591 (N_591,In_1400,In_46);
or U592 (N_592,In_1429,N_453);
nand U593 (N_593,In_66,In_713);
nand U594 (N_594,In_449,In_1109);
nand U595 (N_595,In_937,In_1260);
xor U596 (N_596,N_84,N_303);
nand U597 (N_597,In_1342,In_1113);
or U598 (N_598,N_379,In_660);
nand U599 (N_599,In_1019,In_1232);
and U600 (N_600,In_766,In_579);
nor U601 (N_601,In_441,N_153);
xnor U602 (N_602,N_418,In_1460);
or U603 (N_603,N_94,In_1009);
nor U604 (N_604,N_205,N_339);
and U605 (N_605,N_484,N_174);
nor U606 (N_606,In_747,N_390);
nand U607 (N_607,In_278,N_14);
or U608 (N_608,In_531,N_329);
nor U609 (N_609,In_229,In_1447);
xnor U610 (N_610,In_1273,N_226);
and U611 (N_611,In_666,N_114);
nand U612 (N_612,In_218,In_75);
and U613 (N_613,In_125,In_922);
nand U614 (N_614,In_506,N_285);
or U615 (N_615,In_1026,In_861);
and U616 (N_616,In_1410,N_299);
or U617 (N_617,In_1227,N_478);
xor U618 (N_618,N_89,In_336);
or U619 (N_619,In_349,In_300);
or U620 (N_620,In_1126,In_811);
nand U621 (N_621,N_231,N_136);
xnor U622 (N_622,N_148,N_101);
or U623 (N_623,In_91,In_192);
or U624 (N_624,In_1211,In_1488);
xnor U625 (N_625,In_190,In_1000);
nand U626 (N_626,N_394,In_490);
and U627 (N_627,N_381,N_495);
xor U628 (N_628,In_388,N_371);
nand U629 (N_629,N_496,N_147);
nand U630 (N_630,In_855,In_881);
or U631 (N_631,N_116,N_441);
or U632 (N_632,In_173,In_255);
xor U633 (N_633,In_730,N_469);
nor U634 (N_634,In_773,In_819);
nand U635 (N_635,In_137,In_57);
and U636 (N_636,N_532,In_1248);
xnor U637 (N_637,In_832,N_499);
nor U638 (N_638,N_518,N_419);
and U639 (N_639,In_1307,In_1457);
nor U640 (N_640,N_581,In_1128);
xor U641 (N_641,N_609,In_435);
nand U642 (N_642,N_280,In_387);
or U643 (N_643,In_364,N_570);
or U644 (N_644,In_955,In_466);
nor U645 (N_645,In_1186,N_557);
nor U646 (N_646,N_399,In_680);
nor U647 (N_647,N_203,In_114);
nand U648 (N_648,In_78,N_544);
nand U649 (N_649,N_361,N_378);
and U650 (N_650,N_594,N_224);
nand U651 (N_651,N_382,In_1468);
nor U652 (N_652,N_598,In_1224);
nand U653 (N_653,N_608,In_359);
nor U654 (N_654,In_1151,N_70);
nor U655 (N_655,In_1168,In_587);
nand U656 (N_656,In_258,N_578);
xor U657 (N_657,N_492,In_1125);
and U658 (N_658,N_284,N_383);
xnor U659 (N_659,In_824,In_138);
xor U660 (N_660,N_412,In_412);
xor U661 (N_661,In_483,N_539);
nor U662 (N_662,In_509,In_376);
and U663 (N_663,N_466,In_755);
nor U664 (N_664,N_402,N_447);
and U665 (N_665,In_143,In_342);
or U666 (N_666,In_107,In_702);
xnor U667 (N_667,N_9,N_267);
nand U668 (N_668,In_851,In_1110);
xor U669 (N_669,N_586,N_460);
and U670 (N_670,N_277,N_444);
or U671 (N_671,In_230,In_1238);
nor U672 (N_672,In_609,N_405);
nand U673 (N_673,N_410,In_324);
and U674 (N_674,In_343,In_562);
nand U675 (N_675,In_1181,N_396);
nor U676 (N_676,N_376,N_521);
xor U677 (N_677,In_1332,N_575);
nand U678 (N_678,N_476,N_350);
nor U679 (N_679,In_63,In_840);
nor U680 (N_680,In_244,In_332);
and U681 (N_681,In_989,In_721);
and U682 (N_682,In_1094,In_790);
nand U683 (N_683,N_120,N_526);
and U684 (N_684,In_1353,N_515);
and U685 (N_685,N_38,In_427);
nand U686 (N_686,N_456,In_1416);
nand U687 (N_687,N_384,In_465);
and U688 (N_688,N_592,N_523);
or U689 (N_689,In_1377,N_292);
nand U690 (N_690,In_372,In_1038);
and U691 (N_691,N_568,N_561);
nand U692 (N_692,N_509,In_777);
or U693 (N_693,In_103,N_591);
nor U694 (N_694,In_1202,In_613);
and U695 (N_695,N_562,N_296);
nor U696 (N_696,N_613,N_204);
or U697 (N_697,In_1444,In_814);
and U698 (N_698,In_221,In_1097);
or U699 (N_699,In_706,In_1048);
and U700 (N_700,N_503,N_119);
or U701 (N_701,In_419,In_522);
or U702 (N_702,In_206,N_530);
nand U703 (N_703,In_850,N_80);
xnor U704 (N_704,In_1425,In_982);
nor U705 (N_705,N_537,In_276);
xor U706 (N_706,In_134,N_618);
xnor U707 (N_707,In_1215,N_211);
nand U708 (N_708,In_708,In_768);
and U709 (N_709,In_833,In_1212);
and U710 (N_710,N_491,In_169);
and U711 (N_711,N_375,N_131);
nand U712 (N_712,N_563,N_400);
and U713 (N_713,N_279,In_305);
or U714 (N_714,N_533,In_767);
nor U715 (N_715,N_505,In_320);
nand U716 (N_716,N_536,In_993);
and U717 (N_717,In_30,N_389);
nand U718 (N_718,In_549,In_416);
nor U719 (N_719,N_122,In_199);
nand U720 (N_720,N_408,In_573);
xnor U721 (N_721,N_335,N_403);
and U722 (N_722,In_585,In_418);
xor U723 (N_723,N_514,In_805);
or U724 (N_724,In_1344,In_526);
or U725 (N_725,In_636,In_1278);
nand U726 (N_726,In_1464,N_316);
or U727 (N_727,N_181,In_976);
xnor U728 (N_728,N_611,N_597);
or U729 (N_729,N_599,In_1466);
or U730 (N_730,N_471,N_330);
nand U731 (N_731,N_541,In_1435);
xor U732 (N_732,In_1437,N_397);
xnor U733 (N_733,In_975,N_614);
or U734 (N_734,N_457,N_622);
nor U735 (N_735,N_577,N_459);
nand U736 (N_736,In_1456,N_502);
and U737 (N_737,N_326,N_236);
nor U738 (N_738,N_607,In_362);
and U739 (N_739,In_637,In_1287);
nor U740 (N_740,In_897,In_756);
nor U741 (N_741,N_554,In_334);
nor U742 (N_742,N_158,In_316);
and U743 (N_743,In_1394,N_233);
nand U744 (N_744,In_854,In_892);
nor U745 (N_745,N_520,N_548);
nand U746 (N_746,In_942,N_166);
nor U747 (N_747,N_497,In_1223);
xor U748 (N_748,N_567,In_983);
or U749 (N_749,In_1088,In_453);
and U750 (N_750,N_415,N_680);
or U751 (N_751,In_718,In_607);
or U752 (N_752,In_954,In_1486);
xor U753 (N_753,N_129,In_104);
nor U754 (N_754,In_301,N_507);
or U755 (N_755,N_454,In_758);
nor U756 (N_756,In_801,N_305);
and U757 (N_757,N_71,N_631);
xor U758 (N_758,N_393,N_294);
or U759 (N_759,In_411,In_1417);
nand U760 (N_760,In_1155,N_707);
or U761 (N_761,N_60,N_309);
nand U762 (N_762,N_501,In_489);
xnor U763 (N_763,N_508,In_663);
nor U764 (N_764,N_372,N_600);
nor U765 (N_765,In_624,In_815);
or U766 (N_766,In_1117,In_807);
or U767 (N_767,N_749,N_159);
xnor U768 (N_768,In_166,N_364);
nor U769 (N_769,N_727,N_671);
nor U770 (N_770,N_451,N_157);
xor U771 (N_771,In_404,In_1064);
nor U772 (N_772,N_657,N_579);
and U773 (N_773,N_227,N_332);
or U774 (N_774,In_312,N_705);
nor U775 (N_775,In_95,In_1140);
and U776 (N_776,N_74,N_616);
nand U777 (N_777,N_605,N_615);
xor U778 (N_778,In_1367,In_458);
nor U779 (N_779,N_407,In_1331);
or U780 (N_780,In_1369,In_1405);
or U781 (N_781,N_623,In_550);
nor U782 (N_782,N_348,N_525);
xnor U783 (N_783,In_1072,In_867);
and U784 (N_784,In_572,N_109);
nand U785 (N_785,In_739,N_99);
nand U786 (N_786,N_656,In_1443);
or U787 (N_787,In_394,N_261);
xnor U788 (N_788,N_620,N_545);
nand U789 (N_789,N_745,N_670);
xor U790 (N_790,N_741,N_341);
and U791 (N_791,N_138,N_315);
or U792 (N_792,N_564,N_747);
or U793 (N_793,N_731,N_528);
and U794 (N_794,N_238,In_787);
nand U795 (N_795,In_1158,N_423);
and U796 (N_796,N_674,N_336);
and U797 (N_797,N_259,N_681);
xnor U798 (N_798,N_718,N_488);
nand U799 (N_799,N_511,In_247);
and U800 (N_800,N_271,In_502);
and U801 (N_801,N_735,In_1056);
nand U802 (N_802,N_610,In_1052);
or U803 (N_803,N_650,In_260);
or U804 (N_804,N_653,N_582);
nor U805 (N_805,N_235,In_967);
xor U806 (N_806,In_974,In_426);
xor U807 (N_807,In_948,N_18);
and U808 (N_808,In_1300,In_17);
or U809 (N_809,In_1231,In_1409);
or U810 (N_810,In_1269,N_273);
or U811 (N_811,In_1436,In_309);
nor U812 (N_812,In_380,N_549);
xnor U813 (N_813,N_274,N_387);
and U814 (N_814,N_734,N_298);
or U815 (N_815,In_519,N_254);
nor U816 (N_816,N_175,N_125);
nand U817 (N_817,N_721,In_865);
xnor U818 (N_818,In_445,N_198);
xor U819 (N_819,In_919,N_377);
or U820 (N_820,In_872,N_140);
xnor U821 (N_821,In_710,In_1254);
nor U822 (N_822,N_362,N_489);
nand U823 (N_823,N_4,N_333);
nor U824 (N_824,In_686,N_649);
nand U825 (N_825,N_596,In_350);
or U826 (N_826,N_356,N_263);
nor U827 (N_827,N_342,In_1093);
xnor U828 (N_828,In_1004,N_416);
xnor U829 (N_829,N_24,N_542);
and U830 (N_830,In_486,In_1189);
and U831 (N_831,N_337,In_742);
and U832 (N_832,N_388,N_429);
xnor U833 (N_833,N_617,N_516);
nor U834 (N_834,N_45,N_161);
xnor U835 (N_835,In_809,N_551);
or U836 (N_836,N_687,In_415);
and U837 (N_837,N_647,N_635);
and U838 (N_838,In_627,In_588);
and U839 (N_839,In_879,N_691);
or U840 (N_840,In_1439,N_638);
and U841 (N_841,N_685,N_746);
and U842 (N_842,N_698,In_358);
xor U843 (N_843,In_887,In_377);
or U844 (N_844,In_1063,In_213);
nor U845 (N_845,In_92,In_1015);
nand U846 (N_846,In_546,N_455);
xnor U847 (N_847,In_684,N_644);
nor U848 (N_848,In_1073,In_620);
nor U849 (N_849,N_346,In_1292);
nand U850 (N_850,In_866,N_589);
nand U851 (N_851,In_420,N_688);
nor U852 (N_852,N_481,N_3);
nand U853 (N_853,N_628,N_714);
nor U854 (N_854,N_100,In_498);
nor U855 (N_855,N_524,N_547);
nand U856 (N_856,In_1362,In_389);
nand U857 (N_857,N_113,In_287);
or U858 (N_858,In_1365,N_658);
xor U859 (N_859,N_370,In_1112);
nand U860 (N_860,N_171,N_264);
and U861 (N_861,In_584,N_307);
nor U862 (N_862,In_1204,In_1397);
and U863 (N_863,In_292,In_495);
nand U864 (N_864,In_691,N_587);
or U865 (N_865,N_646,In_834);
nand U866 (N_866,In_1049,N_458);
or U867 (N_867,In_1233,N_184);
nor U868 (N_868,In_711,N_487);
and U869 (N_869,In_113,N_535);
or U870 (N_870,N_380,N_590);
or U871 (N_871,N_604,In_1027);
and U872 (N_872,N_313,N_686);
or U873 (N_873,In_154,N_676);
or U874 (N_874,N_130,In_616);
xnor U875 (N_875,N_827,N_278);
xor U876 (N_876,N_546,N_654);
and U877 (N_877,In_1025,N_812);
nor U878 (N_878,N_661,N_12);
xor U879 (N_879,N_804,In_629);
xor U880 (N_880,N_845,N_438);
nand U881 (N_881,In_1148,N_435);
xnor U882 (N_882,In_745,In_1255);
or U883 (N_883,In_425,N_436);
nand U884 (N_884,In_1103,N_682);
nor U885 (N_885,N_90,In_1171);
or U886 (N_886,N_145,In_1391);
and U887 (N_887,N_766,N_855);
and U888 (N_888,In_1137,In_829);
or U889 (N_889,N_566,N_652);
and U890 (N_890,N_602,N_716);
xnor U891 (N_891,N_619,N_738);
nor U892 (N_892,In_1492,In_97);
or U893 (N_893,N_808,In_1256);
nor U894 (N_894,In_236,In_1388);
or U895 (N_895,N_796,N_666);
nand U896 (N_896,In_156,N_490);
nand U897 (N_897,N_603,N_150);
nand U898 (N_898,In_1118,N_216);
xor U899 (N_899,N_593,N_655);
or U900 (N_900,In_883,In_839);
or U901 (N_901,N_34,N_683);
nand U902 (N_902,N_543,N_723);
and U903 (N_903,N_866,In_36);
nand U904 (N_904,In_1062,N_756);
xor U905 (N_905,N_787,N_700);
and U906 (N_906,N_837,N_504);
nor U907 (N_907,In_100,In_1350);
nand U908 (N_908,In_930,In_1089);
nor U909 (N_909,In_15,N_850);
or U910 (N_910,In_554,In_405);
xor U911 (N_911,N_719,N_849);
xnor U912 (N_912,In_398,N_699);
or U913 (N_913,N_552,N_709);
nand U914 (N_914,In_1061,N_494);
or U915 (N_915,N_470,N_662);
nor U916 (N_916,N_443,N_791);
or U917 (N_917,N_629,N_835);
or U918 (N_918,In_452,N_584);
and U919 (N_919,In_1169,In_898);
xor U920 (N_920,In_925,In_1337);
nor U921 (N_921,N_270,N_811);
xnor U922 (N_922,N_625,N_391);
nand U923 (N_923,In_481,N_824);
nand U924 (N_924,N_846,N_624);
xor U925 (N_925,N_445,N_659);
and U926 (N_926,In_846,In_77);
xnor U927 (N_927,In_1213,In_1358);
nand U928 (N_928,In_216,N_853);
and U929 (N_929,In_1423,N_493);
and U930 (N_930,N_463,In_670);
nor U931 (N_931,N_645,In_717);
xor U932 (N_932,In_361,N_281);
and U933 (N_933,N_439,N_717);
nand U934 (N_934,N_832,N_778);
and U935 (N_935,In_473,N_867);
xor U936 (N_936,In_1271,In_257);
nand U937 (N_937,In_219,In_1090);
nand U938 (N_938,In_1382,In_366);
and U939 (N_939,N_398,In_802);
nor U940 (N_940,In_1264,N_667);
and U941 (N_941,N_232,In_619);
nor U942 (N_942,N_106,N_854);
nand U943 (N_943,In_848,N_799);
nor U944 (N_944,N_406,N_725);
and U945 (N_945,N_763,N_828);
xnor U946 (N_946,N_860,In_1311);
nand U947 (N_947,In_1172,N_580);
nor U948 (N_948,N_743,N_826);
nor U949 (N_949,N_710,N_529);
nor U950 (N_950,N_701,In_842);
nor U951 (N_951,N_310,N_612);
and U952 (N_952,N_199,In_639);
nand U953 (N_953,In_1411,N_810);
or U954 (N_954,N_572,N_434);
xor U955 (N_955,N_558,N_869);
and U956 (N_956,In_981,N_697);
nand U957 (N_957,In_1280,N_601);
or U958 (N_958,N_800,In_646);
nand U959 (N_959,N_868,N_417);
or U960 (N_960,In_2,N_792);
nand U961 (N_961,N_844,In_182);
nand U962 (N_962,In_734,In_392);
nor U963 (N_963,N_695,N_556);
and U964 (N_964,N_872,N_782);
and U965 (N_965,In_1478,N_595);
xnor U966 (N_966,N_354,In_1251);
nor U967 (N_967,N_818,In_714);
or U968 (N_968,In_593,In_857);
nor U969 (N_969,In_1216,N_187);
and U970 (N_970,N_286,In_970);
xor U971 (N_971,In_1182,N_651);
and U972 (N_972,N_367,N_480);
nand U973 (N_973,N_838,In_1296);
nand U974 (N_974,N_409,In_500);
or U975 (N_975,In_1206,N_809);
or U976 (N_976,N_820,N_648);
or U977 (N_977,In_1057,N_498);
nand U978 (N_978,N_540,In_131);
nor U979 (N_979,In_728,N_757);
and U980 (N_980,N_559,In_87);
nor U981 (N_981,N_774,N_322);
and U982 (N_982,N_208,N_200);
and U983 (N_983,In_238,N_873);
and U984 (N_984,In_899,N_626);
nor U985 (N_985,N_565,N_668);
nand U986 (N_986,In_1283,N_786);
nor U987 (N_987,N_630,N_553);
nor U988 (N_988,N_571,In_1129);
or U989 (N_989,In_1205,N_477);
or U990 (N_990,N_806,N_862);
nand U991 (N_991,N_783,N_426);
or U992 (N_992,N_155,In_984);
or U993 (N_993,N_736,In_1308);
nand U994 (N_994,N_252,N_482);
and U995 (N_995,In_407,In_985);
nor U996 (N_996,N_5,N_767);
xnor U997 (N_997,In_1440,In_184);
and U998 (N_998,N_852,N_797);
nand U999 (N_999,N_843,N_805);
nand U1000 (N_1000,N_739,N_913);
nand U1001 (N_1001,N_770,In_60);
nor U1002 (N_1002,In_800,N_679);
nand U1003 (N_1003,N_452,N_978);
nand U1004 (N_1004,N_926,N_219);
or U1005 (N_1005,In_568,N_989);
and U1006 (N_1006,N_365,N_715);
xnor U1007 (N_1007,N_919,N_574);
nand U1008 (N_1008,In_1372,N_250);
and U1009 (N_1009,N_890,N_425);
and U1010 (N_1010,In_885,N_517);
or U1011 (N_1011,In_765,N_998);
or U1012 (N_1012,N_798,N_677);
nor U1013 (N_1013,N_947,N_253);
xor U1014 (N_1014,N_321,N_752);
and U1015 (N_1015,In_1426,In_749);
xor U1016 (N_1016,N_946,N_908);
nand U1017 (N_1017,N_124,N_987);
nor U1018 (N_1018,In_618,N_871);
and U1019 (N_1019,In_753,N_881);
or U1020 (N_1020,N_980,In_574);
xnor U1021 (N_1021,In_580,N_958);
xnor U1022 (N_1022,N_874,N_807);
nand U1023 (N_1023,In_1083,N_983);
nand U1024 (N_1024,In_598,In_275);
or U1025 (N_1025,In_673,N_929);
nor U1026 (N_1026,N_942,In_21);
nor U1027 (N_1027,N_744,N_931);
or U1028 (N_1028,N_762,N_195);
or U1029 (N_1029,N_328,N_127);
and U1030 (N_1030,N_864,N_967);
or U1031 (N_1031,In_220,In_38);
nand U1032 (N_1032,N_66,In_1252);
or U1033 (N_1033,In_707,N_58);
nand U1034 (N_1034,N_29,In_162);
nor U1035 (N_1035,N_801,N_971);
or U1036 (N_1036,N_959,N_464);
or U1037 (N_1037,N_414,N_920);
or U1038 (N_1038,N_413,N_664);
xnor U1039 (N_1039,N_640,N_585);
or U1040 (N_1040,N_910,In_1467);
nor U1041 (N_1041,N_802,N_769);
nor U1042 (N_1042,N_149,N_244);
nor U1043 (N_1043,In_311,In_65);
and U1044 (N_1044,In_1080,N_941);
and U1045 (N_1045,In_575,N_737);
nand U1046 (N_1046,N_932,N_923);
nand U1047 (N_1047,N_880,N_814);
nor U1048 (N_1048,N_865,In_1075);
and U1049 (N_1049,N_773,N_760);
nor U1050 (N_1050,N_724,N_424);
or U1051 (N_1051,In_83,N_955);
or U1052 (N_1052,N_202,N_935);
nand U1053 (N_1053,N_851,In_194);
xor U1054 (N_1054,N_833,N_939);
xnor U1055 (N_1055,In_1471,N_133);
xor U1056 (N_1056,N_754,In_1341);
xor U1057 (N_1057,N_693,N_912);
xor U1058 (N_1058,N_334,N_450);
or U1059 (N_1059,N_992,In_1490);
or U1060 (N_1060,In_175,N_85);
or U1061 (N_1061,In_1349,N_550);
xor U1062 (N_1062,N_675,N_794);
or U1063 (N_1063,N_302,In_1356);
or U1064 (N_1064,In_1319,N_373);
and U1065 (N_1065,In_667,N_819);
nand U1066 (N_1066,In_703,N_779);
xor U1067 (N_1067,N_988,N_560);
xnor U1068 (N_1068,N_934,N_909);
nand U1069 (N_1069,N_993,N_981);
xnor U1070 (N_1070,N_961,N_576);
or U1071 (N_1071,N_555,N_750);
xor U1072 (N_1072,N_641,N_928);
and U1073 (N_1073,In_41,N_887);
or U1074 (N_1074,N_969,N_751);
xor U1075 (N_1075,N_422,N_703);
nand U1076 (N_1076,N_722,In_704);
nand U1077 (N_1077,N_994,N_901);
or U1078 (N_1078,In_1345,In_1020);
xor U1079 (N_1079,N_898,N_678);
xnor U1080 (N_1080,N_985,In_1393);
nor U1081 (N_1081,N_903,In_90);
xnor U1082 (N_1082,N_500,N_945);
and U1083 (N_1083,N_742,N_896);
or U1084 (N_1084,N_813,N_990);
or U1085 (N_1085,N_431,N_968);
nand U1086 (N_1086,N_883,N_385);
xor U1087 (N_1087,N_977,N_465);
nor U1088 (N_1088,N_462,In_784);
or U1089 (N_1089,N_673,In_591);
nor U1090 (N_1090,N_949,In_1018);
or U1091 (N_1091,In_327,N_982);
and U1092 (N_1092,N_861,In_631);
xnor U1093 (N_1093,N_392,In_1071);
or U1094 (N_1094,In_918,In_813);
nand U1095 (N_1095,N_975,In_847);
and U1096 (N_1096,N_936,In_723);
xnor U1097 (N_1097,In_672,N_512);
or U1098 (N_1098,N_621,In_690);
and U1099 (N_1099,In_141,N_974);
nand U1100 (N_1100,N_437,In_150);
and U1101 (N_1101,In_906,N_803);
xor U1102 (N_1102,In_858,N_729);
or U1103 (N_1103,N_266,N_162);
and U1104 (N_1104,N_704,In_1289);
nor U1105 (N_1105,N_870,In_757);
xnor U1106 (N_1106,In_111,N_815);
xor U1107 (N_1107,N_642,In_1225);
or U1108 (N_1108,N_748,N_937);
and U1109 (N_1109,N_772,N_964);
or U1110 (N_1110,N_103,In_1348);
or U1111 (N_1111,N_510,N_973);
and U1112 (N_1112,In_931,In_56);
nand U1113 (N_1113,N_768,N_954);
or U1114 (N_1114,N_884,In_323);
nor U1115 (N_1115,N_965,In_1082);
and U1116 (N_1116,N_569,N_534);
nand U1117 (N_1117,N_921,N_997);
nor U1118 (N_1118,N_858,N_882);
or U1119 (N_1119,N_639,N_728);
xnor U1120 (N_1120,N_634,N_900);
nor U1121 (N_1121,N_996,In_1253);
nor U1122 (N_1122,In_67,N_897);
and U1123 (N_1123,N_970,In_564);
nand U1124 (N_1124,N_924,N_950);
and U1125 (N_1125,In_903,N_784);
xor U1126 (N_1126,N_1057,N_726);
or U1127 (N_1127,N_637,N_1008);
xor U1128 (N_1128,N_1106,N_1081);
nor U1129 (N_1129,N_1116,N_1028);
nand U1130 (N_1130,N_169,N_1003);
and U1131 (N_1131,N_1123,N_922);
and U1132 (N_1132,N_112,N_1031);
or U1133 (N_1133,N_446,In_479);
or U1134 (N_1134,N_1030,N_720);
xor U1135 (N_1135,N_712,N_944);
xnor U1136 (N_1136,N_904,N_1054);
or U1137 (N_1137,N_1010,N_758);
nor U1138 (N_1138,N_780,N_899);
xnor U1139 (N_1139,N_583,In_917);
xnor U1140 (N_1140,In_604,N_863);
and U1141 (N_1141,N_1091,N_1087);
xnor U1142 (N_1142,N_976,N_531);
nor U1143 (N_1143,N_972,N_1104);
and U1144 (N_1144,N_421,N_856);
or U1145 (N_1145,In_1293,In_949);
and U1146 (N_1146,N_320,N_573);
nor U1147 (N_1147,In_1247,N_486);
or U1148 (N_1148,N_764,N_1115);
nor U1149 (N_1149,N_180,N_1094);
xnor U1150 (N_1150,N_902,N_708);
nor U1151 (N_1151,N_606,N_1044);
or U1152 (N_1152,N_847,N_1064);
nand U1153 (N_1153,N_918,In_27);
nor U1154 (N_1154,N_943,N_1080);
or U1155 (N_1155,N_1033,N_190);
or U1156 (N_1156,In_110,N_1067);
xnor U1157 (N_1157,N_761,N_1118);
nor U1158 (N_1158,N_1097,N_395);
or U1159 (N_1159,N_627,In_147);
or U1160 (N_1160,N_696,In_1322);
nand U1161 (N_1161,N_355,N_427);
xnor U1162 (N_1162,N_1018,N_829);
xor U1163 (N_1163,N_1025,In_367);
and U1164 (N_1164,In_1266,In_1042);
nor U1165 (N_1165,N_785,N_588);
nor U1166 (N_1166,In_54,In_474);
and U1167 (N_1167,N_1015,N_1016);
nor U1168 (N_1168,N_986,N_892);
nor U1169 (N_1169,N_343,N_979);
nor U1170 (N_1170,N_1050,N_999);
nor U1171 (N_1171,In_243,N_519);
xnor U1172 (N_1172,N_907,In_400);
xnor U1173 (N_1173,N_1113,N_684);
nand U1174 (N_1174,N_357,N_1049);
xor U1175 (N_1175,In_290,In_1188);
or U1176 (N_1176,N_1055,N_894);
and U1177 (N_1177,N_201,N_1023);
or U1178 (N_1178,N_732,N_788);
nand U1179 (N_1179,N_1013,N_1062);
xor U1180 (N_1180,N_1070,In_1091);
or U1181 (N_1181,N_1095,N_139);
or U1182 (N_1182,N_840,N_538);
and U1183 (N_1183,In_1386,N_789);
nor U1184 (N_1184,N_957,N_793);
and U1185 (N_1185,N_821,N_442);
or U1186 (N_1186,In_586,N_522);
nand U1187 (N_1187,In_79,N_1034);
nand U1188 (N_1188,N_1020,N_1002);
or U1189 (N_1189,N_895,In_1139);
or U1190 (N_1190,N_879,N_1029);
or U1191 (N_1191,N_1058,In_1153);
or U1192 (N_1192,N_1022,N_1109);
and U1193 (N_1193,N_1052,N_963);
xnor U1194 (N_1194,In_1024,N_1096);
and U1195 (N_1195,N_877,N_817);
or U1196 (N_1196,N_1075,In_1236);
and U1197 (N_1197,In_281,N_1082);
nor U1198 (N_1198,N_841,N_916);
nor U1199 (N_1199,In_1357,In_158);
nor U1200 (N_1200,N_1039,N_1078);
and U1201 (N_1201,N_991,N_1001);
and U1202 (N_1202,N_1068,N_915);
and U1203 (N_1203,N_776,N_506);
nand U1204 (N_1204,N_891,N_1032);
and U1205 (N_1205,In_501,N_1021);
nor U1206 (N_1206,N_905,N_1060);
and U1207 (N_1207,N_325,N_713);
nand U1208 (N_1208,N_1085,In_1347);
and U1209 (N_1209,In_956,N_823);
nor U1210 (N_1210,N_755,N_39);
and U1211 (N_1211,N_875,N_848);
nand U1212 (N_1212,In_669,N_790);
or U1213 (N_1213,N_1069,In_341);
and U1214 (N_1214,N_1076,N_1107);
or U1215 (N_1215,N_1051,In_563);
nand U1216 (N_1216,N_156,N_706);
nand U1217 (N_1217,N_1004,N_369);
nand U1218 (N_1218,N_694,N_237);
and U1219 (N_1219,In_547,N_1110);
nor U1220 (N_1220,N_995,N_1093);
nand U1221 (N_1221,N_67,N_692);
nor U1222 (N_1222,In_762,N_876);
nor U1223 (N_1223,N_474,N_925);
and U1224 (N_1224,N_1045,N_771);
nand U1225 (N_1225,N_689,N_633);
nand U1226 (N_1226,N_966,In_1078);
nor U1227 (N_1227,In_52,N_822);
nand U1228 (N_1228,N_1041,N_220);
nand U1229 (N_1229,In_20,N_1019);
xor U1230 (N_1230,N_164,N_960);
nand U1231 (N_1231,N_1065,N_1047);
and U1232 (N_1232,N_940,N_906);
or U1233 (N_1233,N_1099,N_911);
nand U1234 (N_1234,N_663,N_160);
nor U1235 (N_1235,N_765,N_1105);
or U1236 (N_1236,In_761,N_1114);
and U1237 (N_1237,N_914,N_1102);
nand U1238 (N_1238,N_291,In_235);
nor U1239 (N_1239,N_878,In_191);
or U1240 (N_1240,N_951,N_152);
and U1241 (N_1241,N_702,In_577);
xor U1242 (N_1242,N_917,In_165);
and U1243 (N_1243,N_53,N_759);
and U1244 (N_1244,In_1014,N_1005);
xnor U1245 (N_1245,N_886,N_669);
xnor U1246 (N_1246,N_1120,N_1071);
xnor U1247 (N_1247,N_1017,N_188);
or U1248 (N_1248,N_825,N_527);
xnor U1249 (N_1249,N_404,N_672);
xnor U1250 (N_1250,N_1000,N_1158);
xnor U1251 (N_1251,In_16,N_1161);
and U1252 (N_1252,N_1132,N_781);
or U1253 (N_1253,N_1155,N_1048);
and U1254 (N_1254,N_1026,N_1159);
and U1255 (N_1255,N_730,In_977);
xor U1256 (N_1256,In_384,N_1190);
or U1257 (N_1257,N_1220,N_1150);
nor U1258 (N_1258,N_930,N_1131);
or U1259 (N_1259,N_265,N_1231);
nor U1260 (N_1260,N_1227,N_1248);
nor U1261 (N_1261,N_1179,N_1122);
or U1262 (N_1262,N_1240,N_1172);
or U1263 (N_1263,N_1199,In_893);
or U1264 (N_1264,N_1239,N_1244);
nor U1265 (N_1265,In_923,N_1042);
xor U1266 (N_1266,In_953,N_1125);
nor U1267 (N_1267,N_1089,N_1143);
xnor U1268 (N_1268,N_1037,N_1200);
nor U1269 (N_1269,N_1061,N_1178);
nand U1270 (N_1270,N_933,N_1140);
and U1271 (N_1271,N_1187,N_1127);
or U1272 (N_1272,N_1012,N_1006);
nor U1273 (N_1273,N_956,N_1126);
nand U1274 (N_1274,N_1171,N_228);
nor U1275 (N_1275,N_1234,N_1014);
and U1276 (N_1276,N_1135,N_386);
or U1277 (N_1277,N_1242,N_1084);
and U1278 (N_1278,N_665,N_1232);
xor U1279 (N_1279,N_1163,N_859);
or U1280 (N_1280,N_1035,N_816);
nand U1281 (N_1281,N_1149,N_893);
and U1282 (N_1282,In_990,N_1083);
nor U1283 (N_1283,N_1134,N_1139);
nor U1284 (N_1284,N_1073,N_1229);
nor U1285 (N_1285,N_1166,N_1213);
nand U1286 (N_1286,N_1157,N_1117);
nor U1287 (N_1287,In_612,N_1249);
nand U1288 (N_1288,N_938,N_1228);
and U1289 (N_1289,In_363,N_836);
nor U1290 (N_1290,N_1088,N_1111);
xnor U1291 (N_1291,N_1112,N_1027);
and U1292 (N_1292,N_948,N_1138);
nor U1293 (N_1293,N_1192,N_1074);
xnor U1294 (N_1294,N_1079,N_1009);
or U1295 (N_1295,N_830,N_1130);
nor U1296 (N_1296,In_1480,N_831);
nand U1297 (N_1297,In_424,N_1136);
or U1298 (N_1298,In_891,N_1038);
xnor U1299 (N_1299,N_48,N_1165);
nand U1300 (N_1300,N_1156,N_1180);
nor U1301 (N_1301,N_1182,N_1043);
nor U1302 (N_1302,N_1141,In_621);
or U1303 (N_1303,N_1216,N_952);
nand U1304 (N_1304,N_1053,N_1145);
nor U1305 (N_1305,N_1210,N_1195);
nand U1306 (N_1306,N_1186,N_1202);
and U1307 (N_1307,N_1103,In_177);
and U1308 (N_1308,N_1147,N_1197);
xor U1309 (N_1309,N_636,N_483);
xor U1310 (N_1310,N_1198,N_1077);
nor U1311 (N_1311,N_1208,N_1226);
xor U1312 (N_1312,In_1406,In_600);
nand U1313 (N_1313,N_311,N_1219);
nand U1314 (N_1314,N_1201,N_1154);
nand U1315 (N_1315,N_1151,N_1146);
nand U1316 (N_1316,N_1108,N_1086);
or U1317 (N_1317,N_1230,N_1191);
or U1318 (N_1318,N_1040,N_1189);
or U1319 (N_1319,N_711,N_857);
or U1320 (N_1320,N_1237,N_1153);
xor U1321 (N_1321,N_1243,N_1100);
nor U1322 (N_1322,N_1204,N_1221);
and U1323 (N_1323,N_1225,N_1211);
nand U1324 (N_1324,N_77,N_1175);
or U1325 (N_1325,N_1212,In_1060);
or U1326 (N_1326,N_753,N_513);
nand U1327 (N_1327,N_1183,N_1152);
xnor U1328 (N_1328,N_1046,N_1119);
or U1329 (N_1329,N_740,N_1142);
xor U1330 (N_1330,N_1133,N_1185);
or U1331 (N_1331,N_1218,N_1090);
xnor U1332 (N_1332,N_1214,N_1170);
nor U1333 (N_1333,In_1277,N_1176);
xnor U1334 (N_1334,N_344,N_1238);
nor U1335 (N_1335,N_885,N_1235);
or U1336 (N_1336,N_927,N_1174);
xor U1337 (N_1337,N_1241,N_1137);
nor U1338 (N_1338,N_888,In_1479);
and U1339 (N_1339,N_1245,N_1066);
or U1340 (N_1340,N_1209,N_1224);
xnor U1341 (N_1341,N_842,N_660);
or U1342 (N_1342,N_1206,In_1065);
xnor U1343 (N_1343,N_1247,N_1128);
nand U1344 (N_1344,In_520,N_1056);
nor U1345 (N_1345,N_1167,N_632);
xor U1346 (N_1346,N_1129,N_962);
and U1347 (N_1347,N_1193,N_775);
and U1348 (N_1348,N_1169,N_1072);
or U1349 (N_1349,In_503,N_1168);
or U1350 (N_1350,N_953,N_1124);
and U1351 (N_1351,N_690,N_795);
nand U1352 (N_1352,N_1215,N_1207);
nor U1353 (N_1353,N_1101,N_1223);
nor U1354 (N_1354,N_1160,N_1063);
nor U1355 (N_1355,N_1007,In_746);
and U1356 (N_1356,N_1236,N_1203);
nand U1357 (N_1357,N_1024,N_1188);
or U1358 (N_1358,N_777,N_1181);
xor U1359 (N_1359,N_733,N_1098);
nand U1360 (N_1360,In_274,In_1095);
and U1361 (N_1361,N_643,N_1092);
and U1362 (N_1362,N_1246,N_401);
nand U1363 (N_1363,N_1177,In_1098);
nor U1364 (N_1364,N_1233,N_1121);
nor U1365 (N_1365,N_889,N_1194);
or U1366 (N_1366,N_1184,N_1164);
nor U1367 (N_1367,N_1205,In_1);
nand U1368 (N_1368,N_473,N_1148);
or U1369 (N_1369,N_1059,N_984);
or U1370 (N_1370,N_1144,N_834);
nand U1371 (N_1371,N_1162,N_1173);
nor U1372 (N_1372,N_1011,N_1036);
or U1373 (N_1373,N_1217,N_1222);
xor U1374 (N_1374,N_1196,N_839);
nand U1375 (N_1375,N_1272,N_1369);
nor U1376 (N_1376,N_1322,N_1364);
nor U1377 (N_1377,N_1273,N_1316);
nand U1378 (N_1378,N_1373,N_1319);
nor U1379 (N_1379,N_1334,N_1343);
nor U1380 (N_1380,N_1366,N_1289);
nand U1381 (N_1381,N_1256,N_1362);
nor U1382 (N_1382,N_1314,N_1265);
or U1383 (N_1383,N_1318,N_1264);
and U1384 (N_1384,N_1338,N_1276);
nand U1385 (N_1385,N_1269,N_1257);
nor U1386 (N_1386,N_1294,N_1359);
xnor U1387 (N_1387,N_1310,N_1287);
nor U1388 (N_1388,N_1296,N_1258);
nor U1389 (N_1389,N_1363,N_1326);
xnor U1390 (N_1390,N_1331,N_1297);
xnor U1391 (N_1391,N_1360,N_1354);
xnor U1392 (N_1392,N_1335,N_1302);
or U1393 (N_1393,N_1267,N_1374);
xor U1394 (N_1394,N_1327,N_1277);
nand U1395 (N_1395,N_1250,N_1266);
and U1396 (N_1396,N_1340,N_1353);
nand U1397 (N_1397,N_1252,N_1309);
xor U1398 (N_1398,N_1370,N_1371);
or U1399 (N_1399,N_1323,N_1357);
xor U1400 (N_1400,N_1358,N_1332);
and U1401 (N_1401,N_1367,N_1303);
nor U1402 (N_1402,N_1270,N_1307);
nor U1403 (N_1403,N_1259,N_1292);
xor U1404 (N_1404,N_1305,N_1308);
nor U1405 (N_1405,N_1281,N_1251);
and U1406 (N_1406,N_1274,N_1325);
or U1407 (N_1407,N_1328,N_1300);
or U1408 (N_1408,N_1283,N_1304);
nand U1409 (N_1409,N_1333,N_1348);
or U1410 (N_1410,N_1282,N_1286);
and U1411 (N_1411,N_1368,N_1284);
and U1412 (N_1412,N_1315,N_1321);
nand U1413 (N_1413,N_1311,N_1290);
nand U1414 (N_1414,N_1271,N_1336);
and U1415 (N_1415,N_1355,N_1285);
nor U1416 (N_1416,N_1299,N_1324);
and U1417 (N_1417,N_1261,N_1313);
nand U1418 (N_1418,N_1275,N_1262);
xnor U1419 (N_1419,N_1339,N_1317);
nor U1420 (N_1420,N_1279,N_1293);
or U1421 (N_1421,N_1342,N_1345);
or U1422 (N_1422,N_1349,N_1295);
or U1423 (N_1423,N_1253,N_1268);
nor U1424 (N_1424,N_1320,N_1372);
nor U1425 (N_1425,N_1330,N_1306);
xnor U1426 (N_1426,N_1352,N_1280);
or U1427 (N_1427,N_1361,N_1346);
and U1428 (N_1428,N_1254,N_1298);
nand U1429 (N_1429,N_1288,N_1344);
or U1430 (N_1430,N_1337,N_1255);
nand U1431 (N_1431,N_1351,N_1329);
xor U1432 (N_1432,N_1301,N_1291);
and U1433 (N_1433,N_1263,N_1350);
xor U1434 (N_1434,N_1356,N_1260);
and U1435 (N_1435,N_1278,N_1347);
and U1436 (N_1436,N_1365,N_1312);
nor U1437 (N_1437,N_1341,N_1330);
or U1438 (N_1438,N_1357,N_1276);
nor U1439 (N_1439,N_1356,N_1326);
nand U1440 (N_1440,N_1367,N_1369);
xor U1441 (N_1441,N_1282,N_1363);
nor U1442 (N_1442,N_1366,N_1326);
or U1443 (N_1443,N_1324,N_1361);
and U1444 (N_1444,N_1268,N_1333);
xor U1445 (N_1445,N_1344,N_1349);
or U1446 (N_1446,N_1365,N_1309);
and U1447 (N_1447,N_1348,N_1336);
xnor U1448 (N_1448,N_1370,N_1274);
nand U1449 (N_1449,N_1313,N_1302);
nor U1450 (N_1450,N_1261,N_1350);
nor U1451 (N_1451,N_1265,N_1337);
xnor U1452 (N_1452,N_1358,N_1373);
nor U1453 (N_1453,N_1278,N_1367);
or U1454 (N_1454,N_1312,N_1309);
nand U1455 (N_1455,N_1272,N_1370);
nor U1456 (N_1456,N_1313,N_1324);
nor U1457 (N_1457,N_1318,N_1336);
or U1458 (N_1458,N_1326,N_1305);
nor U1459 (N_1459,N_1289,N_1326);
and U1460 (N_1460,N_1360,N_1302);
xnor U1461 (N_1461,N_1282,N_1332);
or U1462 (N_1462,N_1347,N_1366);
or U1463 (N_1463,N_1367,N_1363);
nor U1464 (N_1464,N_1254,N_1360);
nor U1465 (N_1465,N_1343,N_1268);
nor U1466 (N_1466,N_1258,N_1338);
or U1467 (N_1467,N_1274,N_1309);
or U1468 (N_1468,N_1374,N_1282);
and U1469 (N_1469,N_1266,N_1337);
xor U1470 (N_1470,N_1270,N_1326);
xor U1471 (N_1471,N_1251,N_1268);
or U1472 (N_1472,N_1304,N_1329);
nand U1473 (N_1473,N_1310,N_1339);
and U1474 (N_1474,N_1342,N_1322);
nor U1475 (N_1475,N_1364,N_1346);
and U1476 (N_1476,N_1250,N_1261);
and U1477 (N_1477,N_1294,N_1280);
or U1478 (N_1478,N_1263,N_1306);
and U1479 (N_1479,N_1327,N_1274);
nor U1480 (N_1480,N_1306,N_1346);
or U1481 (N_1481,N_1269,N_1273);
and U1482 (N_1482,N_1315,N_1275);
and U1483 (N_1483,N_1325,N_1309);
nand U1484 (N_1484,N_1272,N_1317);
and U1485 (N_1485,N_1286,N_1335);
xor U1486 (N_1486,N_1315,N_1345);
and U1487 (N_1487,N_1289,N_1272);
nor U1488 (N_1488,N_1357,N_1282);
nor U1489 (N_1489,N_1278,N_1341);
xor U1490 (N_1490,N_1340,N_1327);
or U1491 (N_1491,N_1261,N_1303);
and U1492 (N_1492,N_1330,N_1260);
nand U1493 (N_1493,N_1353,N_1310);
nor U1494 (N_1494,N_1272,N_1363);
and U1495 (N_1495,N_1295,N_1340);
xor U1496 (N_1496,N_1281,N_1253);
nand U1497 (N_1497,N_1352,N_1270);
and U1498 (N_1498,N_1258,N_1264);
or U1499 (N_1499,N_1308,N_1360);
nand U1500 (N_1500,N_1490,N_1465);
and U1501 (N_1501,N_1479,N_1449);
or U1502 (N_1502,N_1413,N_1440);
or U1503 (N_1503,N_1463,N_1459);
xor U1504 (N_1504,N_1464,N_1484);
nor U1505 (N_1505,N_1397,N_1435);
xor U1506 (N_1506,N_1478,N_1385);
and U1507 (N_1507,N_1388,N_1441);
and U1508 (N_1508,N_1461,N_1383);
and U1509 (N_1509,N_1475,N_1426);
nand U1510 (N_1510,N_1453,N_1411);
and U1511 (N_1511,N_1396,N_1470);
nand U1512 (N_1512,N_1395,N_1438);
or U1513 (N_1513,N_1482,N_1418);
nor U1514 (N_1514,N_1445,N_1422);
and U1515 (N_1515,N_1480,N_1468);
and U1516 (N_1516,N_1416,N_1430);
nor U1517 (N_1517,N_1402,N_1389);
xor U1518 (N_1518,N_1405,N_1429);
and U1519 (N_1519,N_1476,N_1434);
or U1520 (N_1520,N_1447,N_1499);
and U1521 (N_1521,N_1448,N_1380);
and U1522 (N_1522,N_1393,N_1471);
xnor U1523 (N_1523,N_1378,N_1487);
or U1524 (N_1524,N_1424,N_1406);
and U1525 (N_1525,N_1376,N_1451);
nand U1526 (N_1526,N_1392,N_1444);
nand U1527 (N_1527,N_1497,N_1462);
or U1528 (N_1528,N_1417,N_1375);
nor U1529 (N_1529,N_1428,N_1379);
and U1530 (N_1530,N_1391,N_1486);
and U1531 (N_1531,N_1399,N_1458);
nor U1532 (N_1532,N_1457,N_1387);
nand U1533 (N_1533,N_1420,N_1390);
nor U1534 (N_1534,N_1450,N_1386);
nand U1535 (N_1535,N_1432,N_1492);
xor U1536 (N_1536,N_1384,N_1446);
xnor U1537 (N_1537,N_1466,N_1382);
nand U1538 (N_1538,N_1421,N_1442);
nand U1539 (N_1539,N_1454,N_1409);
nor U1540 (N_1540,N_1403,N_1489);
and U1541 (N_1541,N_1493,N_1398);
and U1542 (N_1542,N_1433,N_1419);
xnor U1543 (N_1543,N_1483,N_1496);
nor U1544 (N_1544,N_1404,N_1423);
nand U1545 (N_1545,N_1377,N_1472);
nor U1546 (N_1546,N_1431,N_1412);
nand U1547 (N_1547,N_1495,N_1491);
xor U1548 (N_1548,N_1427,N_1456);
xor U1549 (N_1549,N_1474,N_1477);
and U1550 (N_1550,N_1415,N_1467);
nor U1551 (N_1551,N_1460,N_1407);
nand U1552 (N_1552,N_1443,N_1439);
or U1553 (N_1553,N_1485,N_1494);
and U1554 (N_1554,N_1408,N_1381);
xnor U1555 (N_1555,N_1436,N_1498);
and U1556 (N_1556,N_1400,N_1455);
or U1557 (N_1557,N_1414,N_1401);
or U1558 (N_1558,N_1394,N_1437);
or U1559 (N_1559,N_1473,N_1425);
nand U1560 (N_1560,N_1410,N_1452);
or U1561 (N_1561,N_1488,N_1481);
and U1562 (N_1562,N_1469,N_1428);
nor U1563 (N_1563,N_1418,N_1386);
or U1564 (N_1564,N_1452,N_1421);
and U1565 (N_1565,N_1421,N_1443);
xor U1566 (N_1566,N_1420,N_1498);
xnor U1567 (N_1567,N_1412,N_1389);
and U1568 (N_1568,N_1396,N_1426);
or U1569 (N_1569,N_1425,N_1492);
nor U1570 (N_1570,N_1382,N_1449);
nand U1571 (N_1571,N_1408,N_1488);
or U1572 (N_1572,N_1495,N_1376);
and U1573 (N_1573,N_1417,N_1463);
nand U1574 (N_1574,N_1450,N_1462);
and U1575 (N_1575,N_1388,N_1462);
xor U1576 (N_1576,N_1392,N_1493);
nand U1577 (N_1577,N_1458,N_1426);
nor U1578 (N_1578,N_1475,N_1429);
xnor U1579 (N_1579,N_1401,N_1422);
xor U1580 (N_1580,N_1459,N_1379);
nor U1581 (N_1581,N_1391,N_1497);
nand U1582 (N_1582,N_1413,N_1443);
or U1583 (N_1583,N_1380,N_1463);
nor U1584 (N_1584,N_1461,N_1424);
and U1585 (N_1585,N_1412,N_1415);
and U1586 (N_1586,N_1483,N_1462);
and U1587 (N_1587,N_1482,N_1379);
xnor U1588 (N_1588,N_1419,N_1478);
xnor U1589 (N_1589,N_1494,N_1466);
nand U1590 (N_1590,N_1450,N_1446);
nor U1591 (N_1591,N_1499,N_1388);
xor U1592 (N_1592,N_1392,N_1391);
and U1593 (N_1593,N_1404,N_1420);
or U1594 (N_1594,N_1492,N_1394);
or U1595 (N_1595,N_1484,N_1487);
xnor U1596 (N_1596,N_1447,N_1385);
nand U1597 (N_1597,N_1414,N_1425);
nor U1598 (N_1598,N_1465,N_1486);
or U1599 (N_1599,N_1383,N_1467);
nor U1600 (N_1600,N_1463,N_1493);
nand U1601 (N_1601,N_1382,N_1460);
and U1602 (N_1602,N_1458,N_1419);
nor U1603 (N_1603,N_1472,N_1461);
nor U1604 (N_1604,N_1489,N_1492);
nor U1605 (N_1605,N_1425,N_1459);
xnor U1606 (N_1606,N_1383,N_1415);
and U1607 (N_1607,N_1381,N_1402);
or U1608 (N_1608,N_1388,N_1409);
nor U1609 (N_1609,N_1442,N_1413);
nand U1610 (N_1610,N_1471,N_1496);
nor U1611 (N_1611,N_1384,N_1441);
xnor U1612 (N_1612,N_1454,N_1474);
xnor U1613 (N_1613,N_1426,N_1430);
nor U1614 (N_1614,N_1379,N_1489);
and U1615 (N_1615,N_1481,N_1452);
nand U1616 (N_1616,N_1465,N_1443);
xnor U1617 (N_1617,N_1416,N_1467);
and U1618 (N_1618,N_1429,N_1457);
xnor U1619 (N_1619,N_1400,N_1391);
xnor U1620 (N_1620,N_1477,N_1496);
or U1621 (N_1621,N_1405,N_1388);
or U1622 (N_1622,N_1473,N_1388);
or U1623 (N_1623,N_1430,N_1486);
or U1624 (N_1624,N_1407,N_1490);
nor U1625 (N_1625,N_1566,N_1592);
or U1626 (N_1626,N_1558,N_1532);
and U1627 (N_1627,N_1517,N_1617);
nand U1628 (N_1628,N_1514,N_1610);
nor U1629 (N_1629,N_1593,N_1587);
nor U1630 (N_1630,N_1551,N_1502);
and U1631 (N_1631,N_1546,N_1596);
nor U1632 (N_1632,N_1588,N_1565);
nor U1633 (N_1633,N_1562,N_1619);
nand U1634 (N_1634,N_1611,N_1599);
nand U1635 (N_1635,N_1561,N_1595);
or U1636 (N_1636,N_1525,N_1601);
nor U1637 (N_1637,N_1605,N_1543);
nand U1638 (N_1638,N_1575,N_1600);
or U1639 (N_1639,N_1623,N_1554);
nand U1640 (N_1640,N_1569,N_1537);
or U1641 (N_1641,N_1585,N_1550);
xor U1642 (N_1642,N_1539,N_1507);
and U1643 (N_1643,N_1533,N_1563);
or U1644 (N_1644,N_1509,N_1570);
or U1645 (N_1645,N_1573,N_1621);
xor U1646 (N_1646,N_1607,N_1541);
and U1647 (N_1647,N_1521,N_1518);
xnor U1648 (N_1648,N_1549,N_1597);
nand U1649 (N_1649,N_1545,N_1559);
nand U1650 (N_1650,N_1523,N_1574);
or U1651 (N_1651,N_1624,N_1552);
nand U1652 (N_1652,N_1547,N_1556);
xor U1653 (N_1653,N_1506,N_1584);
or U1654 (N_1654,N_1555,N_1571);
xnor U1655 (N_1655,N_1604,N_1515);
xnor U1656 (N_1656,N_1580,N_1503);
xnor U1657 (N_1657,N_1504,N_1579);
nand U1658 (N_1658,N_1608,N_1582);
and U1659 (N_1659,N_1548,N_1508);
and U1660 (N_1660,N_1538,N_1567);
xor U1661 (N_1661,N_1589,N_1564);
nand U1662 (N_1662,N_1591,N_1516);
and U1663 (N_1663,N_1618,N_1594);
nor U1664 (N_1664,N_1568,N_1529);
or U1665 (N_1665,N_1519,N_1590);
and U1666 (N_1666,N_1524,N_1560);
and U1667 (N_1667,N_1578,N_1540);
nand U1668 (N_1668,N_1602,N_1615);
and U1669 (N_1669,N_1534,N_1622);
nand U1670 (N_1670,N_1510,N_1553);
xnor U1671 (N_1671,N_1603,N_1609);
and U1672 (N_1672,N_1535,N_1613);
nand U1673 (N_1673,N_1616,N_1586);
nor U1674 (N_1674,N_1606,N_1577);
or U1675 (N_1675,N_1527,N_1544);
xor U1676 (N_1676,N_1572,N_1528);
xor U1677 (N_1677,N_1581,N_1620);
nand U1678 (N_1678,N_1505,N_1598);
nand U1679 (N_1679,N_1576,N_1522);
nor U1680 (N_1680,N_1536,N_1531);
or U1681 (N_1681,N_1614,N_1520);
xor U1682 (N_1682,N_1501,N_1542);
nor U1683 (N_1683,N_1557,N_1511);
or U1684 (N_1684,N_1512,N_1612);
or U1685 (N_1685,N_1526,N_1583);
and U1686 (N_1686,N_1530,N_1500);
nor U1687 (N_1687,N_1513,N_1622);
nand U1688 (N_1688,N_1613,N_1622);
and U1689 (N_1689,N_1517,N_1502);
and U1690 (N_1690,N_1579,N_1503);
xor U1691 (N_1691,N_1574,N_1573);
nor U1692 (N_1692,N_1506,N_1624);
and U1693 (N_1693,N_1515,N_1586);
and U1694 (N_1694,N_1502,N_1531);
nor U1695 (N_1695,N_1588,N_1559);
nor U1696 (N_1696,N_1593,N_1604);
xnor U1697 (N_1697,N_1531,N_1594);
or U1698 (N_1698,N_1592,N_1553);
or U1699 (N_1699,N_1601,N_1572);
xor U1700 (N_1700,N_1510,N_1612);
nor U1701 (N_1701,N_1587,N_1580);
or U1702 (N_1702,N_1615,N_1608);
nor U1703 (N_1703,N_1624,N_1576);
nor U1704 (N_1704,N_1544,N_1539);
nand U1705 (N_1705,N_1554,N_1567);
nand U1706 (N_1706,N_1528,N_1593);
nand U1707 (N_1707,N_1507,N_1531);
nand U1708 (N_1708,N_1514,N_1536);
nand U1709 (N_1709,N_1622,N_1549);
nor U1710 (N_1710,N_1509,N_1595);
and U1711 (N_1711,N_1568,N_1611);
and U1712 (N_1712,N_1513,N_1619);
nand U1713 (N_1713,N_1613,N_1581);
or U1714 (N_1714,N_1558,N_1582);
nor U1715 (N_1715,N_1596,N_1536);
nor U1716 (N_1716,N_1573,N_1555);
nor U1717 (N_1717,N_1616,N_1517);
nand U1718 (N_1718,N_1544,N_1581);
or U1719 (N_1719,N_1587,N_1515);
or U1720 (N_1720,N_1575,N_1590);
and U1721 (N_1721,N_1516,N_1542);
nor U1722 (N_1722,N_1571,N_1501);
xnor U1723 (N_1723,N_1565,N_1564);
and U1724 (N_1724,N_1509,N_1501);
and U1725 (N_1725,N_1545,N_1541);
nand U1726 (N_1726,N_1508,N_1563);
and U1727 (N_1727,N_1572,N_1529);
and U1728 (N_1728,N_1610,N_1542);
nand U1729 (N_1729,N_1566,N_1531);
nor U1730 (N_1730,N_1569,N_1539);
or U1731 (N_1731,N_1507,N_1562);
and U1732 (N_1732,N_1581,N_1606);
or U1733 (N_1733,N_1590,N_1596);
and U1734 (N_1734,N_1617,N_1580);
or U1735 (N_1735,N_1591,N_1622);
nand U1736 (N_1736,N_1593,N_1615);
xnor U1737 (N_1737,N_1617,N_1530);
or U1738 (N_1738,N_1614,N_1617);
nor U1739 (N_1739,N_1541,N_1544);
and U1740 (N_1740,N_1521,N_1610);
and U1741 (N_1741,N_1554,N_1564);
and U1742 (N_1742,N_1547,N_1517);
or U1743 (N_1743,N_1616,N_1508);
nor U1744 (N_1744,N_1599,N_1525);
nand U1745 (N_1745,N_1549,N_1517);
or U1746 (N_1746,N_1556,N_1504);
and U1747 (N_1747,N_1532,N_1584);
and U1748 (N_1748,N_1563,N_1580);
nor U1749 (N_1749,N_1610,N_1511);
nand U1750 (N_1750,N_1648,N_1737);
or U1751 (N_1751,N_1679,N_1655);
xor U1752 (N_1752,N_1741,N_1696);
or U1753 (N_1753,N_1712,N_1704);
nor U1754 (N_1754,N_1720,N_1645);
nand U1755 (N_1755,N_1730,N_1680);
and U1756 (N_1756,N_1642,N_1708);
xnor U1757 (N_1757,N_1698,N_1691);
nand U1758 (N_1758,N_1744,N_1724);
nand U1759 (N_1759,N_1742,N_1735);
xnor U1760 (N_1760,N_1699,N_1690);
and U1761 (N_1761,N_1644,N_1686);
or U1762 (N_1762,N_1664,N_1719);
nand U1763 (N_1763,N_1703,N_1625);
and U1764 (N_1764,N_1736,N_1669);
nor U1765 (N_1765,N_1722,N_1677);
nand U1766 (N_1766,N_1632,N_1636);
or U1767 (N_1767,N_1668,N_1674);
or U1768 (N_1768,N_1672,N_1723);
xor U1769 (N_1769,N_1653,N_1656);
nor U1770 (N_1770,N_1713,N_1746);
nor U1771 (N_1771,N_1732,N_1688);
or U1772 (N_1772,N_1738,N_1661);
nor U1773 (N_1773,N_1666,N_1671);
xnor U1774 (N_1774,N_1727,N_1747);
xnor U1775 (N_1775,N_1633,N_1695);
or U1776 (N_1776,N_1675,N_1650);
xnor U1777 (N_1777,N_1647,N_1640);
nand U1778 (N_1778,N_1687,N_1658);
nand U1779 (N_1779,N_1649,N_1706);
or U1780 (N_1780,N_1683,N_1729);
or U1781 (N_1781,N_1748,N_1749);
nor U1782 (N_1782,N_1684,N_1638);
xor U1783 (N_1783,N_1725,N_1657);
nor U1784 (N_1784,N_1629,N_1711);
nor U1785 (N_1785,N_1697,N_1663);
nor U1786 (N_1786,N_1692,N_1739);
nor U1787 (N_1787,N_1630,N_1693);
xor U1788 (N_1788,N_1673,N_1716);
or U1789 (N_1789,N_1682,N_1707);
or U1790 (N_1790,N_1643,N_1681);
or U1791 (N_1791,N_1670,N_1685);
or U1792 (N_1792,N_1641,N_1717);
nor U1793 (N_1793,N_1705,N_1745);
and U1794 (N_1794,N_1628,N_1646);
xnor U1795 (N_1795,N_1651,N_1634);
xor U1796 (N_1796,N_1694,N_1652);
nand U1797 (N_1797,N_1689,N_1700);
or U1798 (N_1798,N_1740,N_1659);
nand U1799 (N_1799,N_1678,N_1728);
nand U1800 (N_1800,N_1710,N_1715);
and U1801 (N_1801,N_1667,N_1702);
and U1802 (N_1802,N_1662,N_1714);
nand U1803 (N_1803,N_1676,N_1635);
nand U1804 (N_1804,N_1631,N_1665);
xor U1805 (N_1805,N_1709,N_1627);
or U1806 (N_1806,N_1637,N_1726);
nor U1807 (N_1807,N_1701,N_1654);
and U1808 (N_1808,N_1743,N_1660);
xor U1809 (N_1809,N_1734,N_1626);
or U1810 (N_1810,N_1731,N_1721);
or U1811 (N_1811,N_1639,N_1733);
or U1812 (N_1812,N_1718,N_1666);
and U1813 (N_1813,N_1695,N_1652);
and U1814 (N_1814,N_1682,N_1694);
xnor U1815 (N_1815,N_1731,N_1688);
nor U1816 (N_1816,N_1642,N_1695);
nand U1817 (N_1817,N_1643,N_1631);
nand U1818 (N_1818,N_1653,N_1663);
xor U1819 (N_1819,N_1635,N_1652);
xnor U1820 (N_1820,N_1713,N_1747);
xor U1821 (N_1821,N_1639,N_1629);
and U1822 (N_1822,N_1685,N_1705);
nor U1823 (N_1823,N_1642,N_1647);
xor U1824 (N_1824,N_1731,N_1650);
nor U1825 (N_1825,N_1677,N_1709);
and U1826 (N_1826,N_1631,N_1656);
or U1827 (N_1827,N_1633,N_1746);
nand U1828 (N_1828,N_1730,N_1692);
xnor U1829 (N_1829,N_1741,N_1712);
nor U1830 (N_1830,N_1652,N_1675);
or U1831 (N_1831,N_1724,N_1645);
and U1832 (N_1832,N_1695,N_1722);
nand U1833 (N_1833,N_1676,N_1721);
or U1834 (N_1834,N_1743,N_1654);
or U1835 (N_1835,N_1631,N_1682);
xor U1836 (N_1836,N_1682,N_1660);
nand U1837 (N_1837,N_1743,N_1672);
or U1838 (N_1838,N_1671,N_1650);
and U1839 (N_1839,N_1638,N_1697);
nor U1840 (N_1840,N_1629,N_1632);
nor U1841 (N_1841,N_1715,N_1697);
nor U1842 (N_1842,N_1632,N_1673);
nor U1843 (N_1843,N_1734,N_1739);
or U1844 (N_1844,N_1666,N_1698);
nor U1845 (N_1845,N_1674,N_1693);
nand U1846 (N_1846,N_1648,N_1730);
nor U1847 (N_1847,N_1673,N_1737);
xor U1848 (N_1848,N_1661,N_1747);
nand U1849 (N_1849,N_1739,N_1691);
nand U1850 (N_1850,N_1708,N_1715);
nor U1851 (N_1851,N_1745,N_1648);
or U1852 (N_1852,N_1690,N_1647);
and U1853 (N_1853,N_1738,N_1712);
or U1854 (N_1854,N_1747,N_1683);
or U1855 (N_1855,N_1735,N_1749);
nor U1856 (N_1856,N_1707,N_1680);
xor U1857 (N_1857,N_1634,N_1657);
nand U1858 (N_1858,N_1652,N_1627);
and U1859 (N_1859,N_1636,N_1701);
xor U1860 (N_1860,N_1700,N_1704);
xnor U1861 (N_1861,N_1655,N_1647);
xor U1862 (N_1862,N_1711,N_1733);
and U1863 (N_1863,N_1696,N_1743);
nand U1864 (N_1864,N_1648,N_1650);
nor U1865 (N_1865,N_1745,N_1662);
nor U1866 (N_1866,N_1671,N_1693);
or U1867 (N_1867,N_1685,N_1677);
or U1868 (N_1868,N_1693,N_1691);
or U1869 (N_1869,N_1675,N_1727);
and U1870 (N_1870,N_1638,N_1661);
or U1871 (N_1871,N_1634,N_1749);
nor U1872 (N_1872,N_1681,N_1704);
and U1873 (N_1873,N_1748,N_1666);
xor U1874 (N_1874,N_1681,N_1725);
nand U1875 (N_1875,N_1817,N_1829);
nand U1876 (N_1876,N_1849,N_1762);
xnor U1877 (N_1877,N_1864,N_1768);
and U1878 (N_1878,N_1833,N_1750);
xnor U1879 (N_1879,N_1805,N_1795);
nand U1880 (N_1880,N_1764,N_1777);
and U1881 (N_1881,N_1774,N_1845);
nor U1882 (N_1882,N_1799,N_1760);
or U1883 (N_1883,N_1838,N_1779);
and U1884 (N_1884,N_1778,N_1852);
nand U1885 (N_1885,N_1843,N_1874);
nand U1886 (N_1886,N_1790,N_1786);
nand U1887 (N_1887,N_1844,N_1818);
nor U1888 (N_1888,N_1772,N_1847);
xor U1889 (N_1889,N_1751,N_1802);
and U1890 (N_1890,N_1857,N_1785);
nand U1891 (N_1891,N_1830,N_1822);
xnor U1892 (N_1892,N_1807,N_1811);
or U1893 (N_1893,N_1752,N_1765);
xnor U1894 (N_1894,N_1835,N_1859);
xnor U1895 (N_1895,N_1839,N_1831);
nand U1896 (N_1896,N_1826,N_1753);
nand U1897 (N_1897,N_1842,N_1856);
nor U1898 (N_1898,N_1797,N_1871);
nor U1899 (N_1899,N_1770,N_1793);
and U1900 (N_1900,N_1809,N_1781);
and U1901 (N_1901,N_1814,N_1780);
nand U1902 (N_1902,N_1800,N_1840);
nand U1903 (N_1903,N_1850,N_1754);
nand U1904 (N_1904,N_1815,N_1810);
nor U1905 (N_1905,N_1816,N_1819);
nor U1906 (N_1906,N_1769,N_1796);
nand U1907 (N_1907,N_1873,N_1862);
and U1908 (N_1908,N_1813,N_1855);
nand U1909 (N_1909,N_1771,N_1773);
and U1910 (N_1910,N_1821,N_1851);
nand U1911 (N_1911,N_1854,N_1755);
nor U1912 (N_1912,N_1792,N_1863);
nor U1913 (N_1913,N_1759,N_1823);
nand U1914 (N_1914,N_1758,N_1787);
or U1915 (N_1915,N_1834,N_1820);
nand U1916 (N_1916,N_1836,N_1782);
xnor U1917 (N_1917,N_1858,N_1798);
nor U1918 (N_1918,N_1824,N_1812);
nor U1919 (N_1919,N_1860,N_1756);
nand U1920 (N_1920,N_1868,N_1848);
xor U1921 (N_1921,N_1866,N_1861);
xor U1922 (N_1922,N_1783,N_1791);
xor U1923 (N_1923,N_1804,N_1763);
or U1924 (N_1924,N_1808,N_1767);
xnor U1925 (N_1925,N_1853,N_1827);
or U1926 (N_1926,N_1766,N_1846);
or U1927 (N_1927,N_1806,N_1867);
and U1928 (N_1928,N_1865,N_1869);
xor U1929 (N_1929,N_1837,N_1841);
nor U1930 (N_1930,N_1789,N_1761);
xnor U1931 (N_1931,N_1803,N_1776);
nand U1932 (N_1932,N_1775,N_1794);
and U1933 (N_1933,N_1784,N_1832);
or U1934 (N_1934,N_1870,N_1801);
xnor U1935 (N_1935,N_1872,N_1757);
and U1936 (N_1936,N_1828,N_1825);
and U1937 (N_1937,N_1788,N_1868);
xnor U1938 (N_1938,N_1763,N_1756);
nor U1939 (N_1939,N_1773,N_1756);
or U1940 (N_1940,N_1819,N_1787);
xnor U1941 (N_1941,N_1765,N_1827);
nor U1942 (N_1942,N_1781,N_1783);
and U1943 (N_1943,N_1856,N_1787);
nand U1944 (N_1944,N_1811,N_1857);
or U1945 (N_1945,N_1856,N_1765);
or U1946 (N_1946,N_1866,N_1765);
and U1947 (N_1947,N_1825,N_1759);
or U1948 (N_1948,N_1825,N_1768);
nor U1949 (N_1949,N_1788,N_1785);
nand U1950 (N_1950,N_1758,N_1781);
and U1951 (N_1951,N_1803,N_1869);
and U1952 (N_1952,N_1753,N_1861);
xnor U1953 (N_1953,N_1774,N_1849);
or U1954 (N_1954,N_1856,N_1753);
and U1955 (N_1955,N_1787,N_1869);
nor U1956 (N_1956,N_1764,N_1795);
nor U1957 (N_1957,N_1779,N_1828);
xor U1958 (N_1958,N_1801,N_1851);
nand U1959 (N_1959,N_1829,N_1770);
nor U1960 (N_1960,N_1846,N_1777);
nand U1961 (N_1961,N_1796,N_1803);
xor U1962 (N_1962,N_1810,N_1766);
xor U1963 (N_1963,N_1858,N_1790);
nor U1964 (N_1964,N_1837,N_1782);
xnor U1965 (N_1965,N_1823,N_1765);
nand U1966 (N_1966,N_1839,N_1808);
or U1967 (N_1967,N_1835,N_1830);
and U1968 (N_1968,N_1826,N_1835);
nand U1969 (N_1969,N_1807,N_1777);
or U1970 (N_1970,N_1767,N_1821);
and U1971 (N_1971,N_1806,N_1848);
nor U1972 (N_1972,N_1853,N_1839);
xor U1973 (N_1973,N_1834,N_1775);
nor U1974 (N_1974,N_1814,N_1822);
and U1975 (N_1975,N_1778,N_1858);
nand U1976 (N_1976,N_1833,N_1814);
xor U1977 (N_1977,N_1793,N_1771);
xor U1978 (N_1978,N_1771,N_1810);
or U1979 (N_1979,N_1857,N_1861);
nand U1980 (N_1980,N_1781,N_1777);
and U1981 (N_1981,N_1802,N_1847);
nor U1982 (N_1982,N_1794,N_1778);
nand U1983 (N_1983,N_1783,N_1810);
or U1984 (N_1984,N_1848,N_1776);
and U1985 (N_1985,N_1820,N_1783);
nand U1986 (N_1986,N_1774,N_1860);
and U1987 (N_1987,N_1841,N_1811);
and U1988 (N_1988,N_1793,N_1773);
nor U1989 (N_1989,N_1805,N_1778);
and U1990 (N_1990,N_1785,N_1845);
nand U1991 (N_1991,N_1768,N_1796);
nand U1992 (N_1992,N_1822,N_1811);
nand U1993 (N_1993,N_1804,N_1831);
nand U1994 (N_1994,N_1859,N_1826);
or U1995 (N_1995,N_1752,N_1851);
and U1996 (N_1996,N_1849,N_1770);
nand U1997 (N_1997,N_1843,N_1777);
or U1998 (N_1998,N_1752,N_1776);
nand U1999 (N_1999,N_1783,N_1853);
xnor U2000 (N_2000,N_1923,N_1942);
or U2001 (N_2001,N_1954,N_1890);
nand U2002 (N_2002,N_1995,N_1884);
and U2003 (N_2003,N_1902,N_1950);
and U2004 (N_2004,N_1883,N_1888);
and U2005 (N_2005,N_1933,N_1955);
xor U2006 (N_2006,N_1897,N_1951);
nor U2007 (N_2007,N_1878,N_1992);
nor U2008 (N_2008,N_1946,N_1931);
xnor U2009 (N_2009,N_1959,N_1948);
and U2010 (N_2010,N_1876,N_1961);
nand U2011 (N_2011,N_1970,N_1974);
nor U2012 (N_2012,N_1965,N_1964);
nand U2013 (N_2013,N_1885,N_1932);
nor U2014 (N_2014,N_1960,N_1994);
nand U2015 (N_2015,N_1913,N_1899);
or U2016 (N_2016,N_1953,N_1912);
nor U2017 (N_2017,N_1920,N_1985);
nor U2018 (N_2018,N_1898,N_1896);
and U2019 (N_2019,N_1988,N_1929);
nand U2020 (N_2020,N_1987,N_1937);
nand U2021 (N_2021,N_1893,N_1983);
or U2022 (N_2022,N_1900,N_1903);
and U2023 (N_2023,N_1962,N_1989);
nor U2024 (N_2024,N_1922,N_1926);
nor U2025 (N_2025,N_1982,N_1958);
nand U2026 (N_2026,N_1892,N_1947);
or U2027 (N_2027,N_1901,N_1921);
and U2028 (N_2028,N_1998,N_1945);
xnor U2029 (N_2029,N_1938,N_1963);
nand U2030 (N_2030,N_1887,N_1935);
and U2031 (N_2031,N_1911,N_1969);
nor U2032 (N_2032,N_1877,N_1977);
and U2033 (N_2033,N_1940,N_1915);
and U2034 (N_2034,N_1906,N_1975);
nand U2035 (N_2035,N_1918,N_1914);
and U2036 (N_2036,N_1928,N_1881);
nor U2037 (N_2037,N_1875,N_1981);
nand U2038 (N_2038,N_1882,N_1956);
xnor U2039 (N_2039,N_1991,N_1949);
xor U2040 (N_2040,N_1886,N_1909);
nor U2041 (N_2041,N_1957,N_1967);
and U2042 (N_2042,N_1891,N_1925);
nor U2043 (N_2043,N_1927,N_1910);
xor U2044 (N_2044,N_1895,N_1972);
nor U2045 (N_2045,N_1966,N_1984);
and U2046 (N_2046,N_1980,N_1979);
nor U2047 (N_2047,N_1936,N_1973);
or U2048 (N_2048,N_1904,N_1880);
nand U2049 (N_2049,N_1943,N_1997);
xnor U2050 (N_2050,N_1996,N_1919);
nor U2051 (N_2051,N_1907,N_1905);
xnor U2052 (N_2052,N_1894,N_1934);
or U2053 (N_2053,N_1968,N_1939);
nor U2054 (N_2054,N_1971,N_1924);
nor U2055 (N_2055,N_1993,N_1990);
xnor U2056 (N_2056,N_1930,N_1976);
nor U2057 (N_2057,N_1941,N_1917);
or U2058 (N_2058,N_1978,N_1944);
and U2059 (N_2059,N_1889,N_1908);
and U2060 (N_2060,N_1999,N_1986);
nand U2061 (N_2061,N_1952,N_1916);
or U2062 (N_2062,N_1879,N_1924);
nor U2063 (N_2063,N_1889,N_1898);
nor U2064 (N_2064,N_1937,N_1955);
nand U2065 (N_2065,N_1924,N_1929);
xor U2066 (N_2066,N_1971,N_1960);
or U2067 (N_2067,N_1903,N_1879);
nor U2068 (N_2068,N_1950,N_1878);
xnor U2069 (N_2069,N_1954,N_1932);
and U2070 (N_2070,N_1881,N_1901);
and U2071 (N_2071,N_1924,N_1941);
and U2072 (N_2072,N_1986,N_1982);
xor U2073 (N_2073,N_1948,N_1946);
nand U2074 (N_2074,N_1983,N_1918);
and U2075 (N_2075,N_1962,N_1966);
nor U2076 (N_2076,N_1938,N_1914);
or U2077 (N_2077,N_1981,N_1941);
and U2078 (N_2078,N_1957,N_1965);
nand U2079 (N_2079,N_1896,N_1901);
xnor U2080 (N_2080,N_1974,N_1907);
and U2081 (N_2081,N_1918,N_1943);
and U2082 (N_2082,N_1901,N_1903);
and U2083 (N_2083,N_1923,N_1925);
and U2084 (N_2084,N_1931,N_1903);
nor U2085 (N_2085,N_1948,N_1978);
nor U2086 (N_2086,N_1957,N_1979);
nand U2087 (N_2087,N_1954,N_1958);
and U2088 (N_2088,N_1992,N_1894);
xnor U2089 (N_2089,N_1908,N_1969);
or U2090 (N_2090,N_1970,N_1884);
nand U2091 (N_2091,N_1928,N_1943);
or U2092 (N_2092,N_1914,N_1950);
nand U2093 (N_2093,N_1913,N_1979);
nor U2094 (N_2094,N_1902,N_1922);
or U2095 (N_2095,N_1878,N_1900);
nand U2096 (N_2096,N_1938,N_1881);
nand U2097 (N_2097,N_1983,N_1958);
nand U2098 (N_2098,N_1941,N_1944);
xor U2099 (N_2099,N_1920,N_1955);
nand U2100 (N_2100,N_1977,N_1932);
and U2101 (N_2101,N_1923,N_1938);
or U2102 (N_2102,N_1913,N_1993);
nor U2103 (N_2103,N_1924,N_1895);
xnor U2104 (N_2104,N_1980,N_1888);
nand U2105 (N_2105,N_1981,N_1959);
or U2106 (N_2106,N_1965,N_1933);
nand U2107 (N_2107,N_1916,N_1960);
nand U2108 (N_2108,N_1916,N_1903);
xnor U2109 (N_2109,N_1973,N_1997);
nor U2110 (N_2110,N_1964,N_1895);
xnor U2111 (N_2111,N_1970,N_1930);
nand U2112 (N_2112,N_1987,N_1889);
nand U2113 (N_2113,N_1900,N_1911);
nand U2114 (N_2114,N_1997,N_1936);
and U2115 (N_2115,N_1955,N_1881);
or U2116 (N_2116,N_1882,N_1929);
nor U2117 (N_2117,N_1982,N_1972);
nor U2118 (N_2118,N_1989,N_1954);
nor U2119 (N_2119,N_1935,N_1946);
and U2120 (N_2120,N_1915,N_1996);
nand U2121 (N_2121,N_1911,N_1979);
nor U2122 (N_2122,N_1974,N_1949);
and U2123 (N_2123,N_1999,N_1893);
nand U2124 (N_2124,N_1938,N_1986);
nand U2125 (N_2125,N_2101,N_2000);
nor U2126 (N_2126,N_2094,N_2118);
and U2127 (N_2127,N_2107,N_2124);
or U2128 (N_2128,N_2114,N_2034);
and U2129 (N_2129,N_2057,N_2030);
and U2130 (N_2130,N_2042,N_2044);
or U2131 (N_2131,N_2008,N_2065);
nand U2132 (N_2132,N_2096,N_2012);
and U2133 (N_2133,N_2009,N_2120);
nand U2134 (N_2134,N_2004,N_2075);
xnor U2135 (N_2135,N_2122,N_2084);
nor U2136 (N_2136,N_2010,N_2046);
nand U2137 (N_2137,N_2028,N_2089);
and U2138 (N_2138,N_2091,N_2013);
xnor U2139 (N_2139,N_2056,N_2104);
nand U2140 (N_2140,N_2092,N_2006);
and U2141 (N_2141,N_2063,N_2053);
nand U2142 (N_2142,N_2025,N_2062);
nand U2143 (N_2143,N_2037,N_2069);
and U2144 (N_2144,N_2090,N_2111);
nor U2145 (N_2145,N_2060,N_2105);
nor U2146 (N_2146,N_2066,N_2020);
xor U2147 (N_2147,N_2074,N_2070);
xor U2148 (N_2148,N_2001,N_2061);
and U2149 (N_2149,N_2072,N_2102);
nand U2150 (N_2150,N_2049,N_2007);
xor U2151 (N_2151,N_2109,N_2005);
or U2152 (N_2152,N_2031,N_2050);
or U2153 (N_2153,N_2115,N_2011);
and U2154 (N_2154,N_2071,N_2018);
nand U2155 (N_2155,N_2059,N_2108);
and U2156 (N_2156,N_2058,N_2048);
and U2157 (N_2157,N_2117,N_2083);
or U2158 (N_2158,N_2045,N_2055);
nor U2159 (N_2159,N_2022,N_2015);
or U2160 (N_2160,N_2047,N_2024);
or U2161 (N_2161,N_2097,N_2032);
and U2162 (N_2162,N_2087,N_2113);
or U2163 (N_2163,N_2116,N_2021);
xnor U2164 (N_2164,N_2067,N_2014);
and U2165 (N_2165,N_2040,N_2019);
and U2166 (N_2166,N_2079,N_2099);
and U2167 (N_2167,N_2064,N_2054);
nand U2168 (N_2168,N_2016,N_2082);
and U2169 (N_2169,N_2100,N_2123);
xor U2170 (N_2170,N_2098,N_2026);
xnor U2171 (N_2171,N_2076,N_2095);
nor U2172 (N_2172,N_2038,N_2103);
xor U2173 (N_2173,N_2043,N_2035);
nor U2174 (N_2174,N_2080,N_2086);
nor U2175 (N_2175,N_2041,N_2077);
nand U2176 (N_2176,N_2002,N_2085);
nor U2177 (N_2177,N_2003,N_2121);
nand U2178 (N_2178,N_2081,N_2036);
nor U2179 (N_2179,N_2033,N_2088);
nor U2180 (N_2180,N_2110,N_2119);
or U2181 (N_2181,N_2052,N_2093);
xor U2182 (N_2182,N_2106,N_2039);
and U2183 (N_2183,N_2073,N_2027);
and U2184 (N_2184,N_2078,N_2112);
and U2185 (N_2185,N_2068,N_2029);
nor U2186 (N_2186,N_2017,N_2023);
or U2187 (N_2187,N_2051,N_2078);
nand U2188 (N_2188,N_2098,N_2095);
or U2189 (N_2189,N_2091,N_2118);
xnor U2190 (N_2190,N_2075,N_2018);
nor U2191 (N_2191,N_2022,N_2093);
or U2192 (N_2192,N_2065,N_2016);
and U2193 (N_2193,N_2037,N_2041);
xor U2194 (N_2194,N_2086,N_2047);
or U2195 (N_2195,N_2085,N_2123);
or U2196 (N_2196,N_2086,N_2052);
nor U2197 (N_2197,N_2003,N_2034);
nand U2198 (N_2198,N_2096,N_2080);
nand U2199 (N_2199,N_2095,N_2121);
xnor U2200 (N_2200,N_2097,N_2005);
xor U2201 (N_2201,N_2060,N_2087);
nor U2202 (N_2202,N_2113,N_2099);
or U2203 (N_2203,N_2062,N_2072);
xnor U2204 (N_2204,N_2014,N_2099);
nor U2205 (N_2205,N_2024,N_2080);
nor U2206 (N_2206,N_2095,N_2113);
nand U2207 (N_2207,N_2011,N_2029);
or U2208 (N_2208,N_2037,N_2039);
nand U2209 (N_2209,N_2073,N_2047);
or U2210 (N_2210,N_2049,N_2089);
nand U2211 (N_2211,N_2035,N_2098);
and U2212 (N_2212,N_2036,N_2060);
or U2213 (N_2213,N_2119,N_2005);
xnor U2214 (N_2214,N_2091,N_2019);
nand U2215 (N_2215,N_2052,N_2066);
or U2216 (N_2216,N_2075,N_2028);
or U2217 (N_2217,N_2048,N_2035);
xnor U2218 (N_2218,N_2070,N_2017);
nor U2219 (N_2219,N_2017,N_2008);
nand U2220 (N_2220,N_2085,N_2062);
nor U2221 (N_2221,N_2052,N_2065);
or U2222 (N_2222,N_2054,N_2044);
nand U2223 (N_2223,N_2056,N_2002);
xnor U2224 (N_2224,N_2114,N_2024);
nand U2225 (N_2225,N_2079,N_2117);
nand U2226 (N_2226,N_2033,N_2082);
nand U2227 (N_2227,N_2000,N_2097);
nand U2228 (N_2228,N_2104,N_2050);
or U2229 (N_2229,N_2016,N_2039);
and U2230 (N_2230,N_2112,N_2081);
xnor U2231 (N_2231,N_2099,N_2093);
or U2232 (N_2232,N_2003,N_2059);
nor U2233 (N_2233,N_2003,N_2057);
xnor U2234 (N_2234,N_2110,N_2116);
or U2235 (N_2235,N_2117,N_2120);
nand U2236 (N_2236,N_2067,N_2056);
nand U2237 (N_2237,N_2024,N_2020);
nand U2238 (N_2238,N_2034,N_2047);
xnor U2239 (N_2239,N_2004,N_2109);
or U2240 (N_2240,N_2006,N_2022);
nand U2241 (N_2241,N_2117,N_2115);
and U2242 (N_2242,N_2004,N_2121);
nor U2243 (N_2243,N_2096,N_2084);
nand U2244 (N_2244,N_2074,N_2031);
xnor U2245 (N_2245,N_2078,N_2022);
nand U2246 (N_2246,N_2051,N_2101);
xnor U2247 (N_2247,N_2095,N_2020);
or U2248 (N_2248,N_2111,N_2021);
and U2249 (N_2249,N_2005,N_2044);
xnor U2250 (N_2250,N_2240,N_2197);
nor U2251 (N_2251,N_2158,N_2205);
nand U2252 (N_2252,N_2146,N_2198);
and U2253 (N_2253,N_2248,N_2165);
xnor U2254 (N_2254,N_2208,N_2164);
nor U2255 (N_2255,N_2238,N_2142);
or U2256 (N_2256,N_2199,N_2176);
and U2257 (N_2257,N_2228,N_2174);
and U2258 (N_2258,N_2215,N_2173);
xor U2259 (N_2259,N_2128,N_2213);
nor U2260 (N_2260,N_2230,N_2217);
nand U2261 (N_2261,N_2239,N_2187);
or U2262 (N_2262,N_2138,N_2149);
nand U2263 (N_2263,N_2184,N_2135);
and U2264 (N_2264,N_2150,N_2237);
xor U2265 (N_2265,N_2136,N_2125);
and U2266 (N_2266,N_2185,N_2129);
nand U2267 (N_2267,N_2143,N_2233);
nor U2268 (N_2268,N_2211,N_2172);
and U2269 (N_2269,N_2157,N_2226);
nor U2270 (N_2270,N_2132,N_2231);
nor U2271 (N_2271,N_2227,N_2168);
xor U2272 (N_2272,N_2207,N_2148);
nand U2273 (N_2273,N_2234,N_2133);
or U2274 (N_2274,N_2181,N_2245);
or U2275 (N_2275,N_2242,N_2202);
and U2276 (N_2276,N_2201,N_2222);
nand U2277 (N_2277,N_2137,N_2126);
xnor U2278 (N_2278,N_2200,N_2166);
and U2279 (N_2279,N_2189,N_2195);
and U2280 (N_2280,N_2216,N_2139);
or U2281 (N_2281,N_2224,N_2221);
or U2282 (N_2282,N_2210,N_2183);
or U2283 (N_2283,N_2209,N_2163);
nor U2284 (N_2284,N_2127,N_2162);
or U2285 (N_2285,N_2167,N_2170);
and U2286 (N_2286,N_2175,N_2204);
nand U2287 (N_2287,N_2147,N_2193);
or U2288 (N_2288,N_2249,N_2241);
nor U2289 (N_2289,N_2196,N_2134);
and U2290 (N_2290,N_2179,N_2140);
or U2291 (N_2291,N_2206,N_2156);
xnor U2292 (N_2292,N_2153,N_2236);
and U2293 (N_2293,N_2130,N_2192);
nand U2294 (N_2294,N_2144,N_2177);
or U2295 (N_2295,N_2229,N_2246);
xor U2296 (N_2296,N_2219,N_2203);
nor U2297 (N_2297,N_2194,N_2244);
nand U2298 (N_2298,N_2212,N_2223);
xor U2299 (N_2299,N_2182,N_2171);
nand U2300 (N_2300,N_2235,N_2188);
xnor U2301 (N_2301,N_2161,N_2180);
nand U2302 (N_2302,N_2232,N_2160);
nor U2303 (N_2303,N_2190,N_2141);
nor U2304 (N_2304,N_2152,N_2247);
nand U2305 (N_2305,N_2191,N_2159);
nor U2306 (N_2306,N_2225,N_2131);
xnor U2307 (N_2307,N_2218,N_2214);
nand U2308 (N_2308,N_2154,N_2145);
xor U2309 (N_2309,N_2178,N_2151);
or U2310 (N_2310,N_2243,N_2155);
or U2311 (N_2311,N_2186,N_2169);
or U2312 (N_2312,N_2220,N_2171);
xnor U2313 (N_2313,N_2160,N_2162);
and U2314 (N_2314,N_2234,N_2197);
and U2315 (N_2315,N_2141,N_2147);
nand U2316 (N_2316,N_2170,N_2182);
nor U2317 (N_2317,N_2139,N_2211);
nor U2318 (N_2318,N_2245,N_2191);
nor U2319 (N_2319,N_2244,N_2188);
or U2320 (N_2320,N_2209,N_2235);
nand U2321 (N_2321,N_2180,N_2139);
or U2322 (N_2322,N_2191,N_2167);
and U2323 (N_2323,N_2183,N_2226);
and U2324 (N_2324,N_2236,N_2188);
or U2325 (N_2325,N_2204,N_2147);
nor U2326 (N_2326,N_2201,N_2196);
and U2327 (N_2327,N_2139,N_2168);
and U2328 (N_2328,N_2185,N_2144);
nand U2329 (N_2329,N_2159,N_2240);
xor U2330 (N_2330,N_2159,N_2141);
nand U2331 (N_2331,N_2247,N_2184);
or U2332 (N_2332,N_2222,N_2150);
nand U2333 (N_2333,N_2183,N_2177);
and U2334 (N_2334,N_2206,N_2242);
or U2335 (N_2335,N_2148,N_2162);
nor U2336 (N_2336,N_2219,N_2131);
nand U2337 (N_2337,N_2156,N_2183);
nand U2338 (N_2338,N_2241,N_2149);
or U2339 (N_2339,N_2242,N_2131);
nor U2340 (N_2340,N_2125,N_2188);
nor U2341 (N_2341,N_2163,N_2216);
and U2342 (N_2342,N_2171,N_2154);
xor U2343 (N_2343,N_2178,N_2134);
nor U2344 (N_2344,N_2152,N_2204);
or U2345 (N_2345,N_2156,N_2155);
or U2346 (N_2346,N_2233,N_2197);
and U2347 (N_2347,N_2152,N_2200);
nand U2348 (N_2348,N_2234,N_2211);
xor U2349 (N_2349,N_2130,N_2207);
xor U2350 (N_2350,N_2157,N_2233);
xor U2351 (N_2351,N_2212,N_2190);
nor U2352 (N_2352,N_2229,N_2233);
and U2353 (N_2353,N_2147,N_2238);
xor U2354 (N_2354,N_2193,N_2203);
nor U2355 (N_2355,N_2156,N_2199);
and U2356 (N_2356,N_2244,N_2234);
and U2357 (N_2357,N_2153,N_2246);
or U2358 (N_2358,N_2166,N_2137);
xor U2359 (N_2359,N_2169,N_2215);
or U2360 (N_2360,N_2145,N_2150);
or U2361 (N_2361,N_2238,N_2132);
nand U2362 (N_2362,N_2171,N_2214);
or U2363 (N_2363,N_2131,N_2192);
nor U2364 (N_2364,N_2226,N_2160);
xnor U2365 (N_2365,N_2130,N_2137);
or U2366 (N_2366,N_2186,N_2216);
and U2367 (N_2367,N_2191,N_2238);
xnor U2368 (N_2368,N_2224,N_2141);
and U2369 (N_2369,N_2225,N_2151);
nand U2370 (N_2370,N_2143,N_2179);
nor U2371 (N_2371,N_2153,N_2209);
or U2372 (N_2372,N_2237,N_2148);
nand U2373 (N_2373,N_2157,N_2189);
nor U2374 (N_2374,N_2143,N_2132);
or U2375 (N_2375,N_2306,N_2337);
or U2376 (N_2376,N_2360,N_2267);
xor U2377 (N_2377,N_2282,N_2280);
nor U2378 (N_2378,N_2349,N_2259);
xor U2379 (N_2379,N_2341,N_2355);
xor U2380 (N_2380,N_2340,N_2289);
and U2381 (N_2381,N_2262,N_2313);
and U2382 (N_2382,N_2298,N_2373);
or U2383 (N_2383,N_2351,N_2312);
nor U2384 (N_2384,N_2348,N_2332);
or U2385 (N_2385,N_2356,N_2270);
and U2386 (N_2386,N_2308,N_2350);
and U2387 (N_2387,N_2324,N_2319);
nand U2388 (N_2388,N_2305,N_2257);
nand U2389 (N_2389,N_2250,N_2374);
or U2390 (N_2390,N_2294,N_2309);
and U2391 (N_2391,N_2344,N_2307);
and U2392 (N_2392,N_2271,N_2327);
or U2393 (N_2393,N_2304,N_2335);
and U2394 (N_2394,N_2297,N_2264);
nor U2395 (N_2395,N_2368,N_2329);
xnor U2396 (N_2396,N_2261,N_2287);
nand U2397 (N_2397,N_2253,N_2302);
and U2398 (N_2398,N_2322,N_2275);
nor U2399 (N_2399,N_2310,N_2320);
nand U2400 (N_2400,N_2292,N_2254);
nand U2401 (N_2401,N_2252,N_2342);
nand U2402 (N_2402,N_2325,N_2359);
and U2403 (N_2403,N_2343,N_2326);
nor U2404 (N_2404,N_2290,N_2339);
xnor U2405 (N_2405,N_2272,N_2353);
nand U2406 (N_2406,N_2334,N_2278);
xor U2407 (N_2407,N_2362,N_2314);
xor U2408 (N_2408,N_2251,N_2285);
and U2409 (N_2409,N_2358,N_2315);
or U2410 (N_2410,N_2256,N_2372);
xor U2411 (N_2411,N_2345,N_2333);
and U2412 (N_2412,N_2352,N_2318);
or U2413 (N_2413,N_2331,N_2364);
nor U2414 (N_2414,N_2279,N_2366);
nor U2415 (N_2415,N_2301,N_2274);
xor U2416 (N_2416,N_2258,N_2269);
or U2417 (N_2417,N_2303,N_2370);
or U2418 (N_2418,N_2277,N_2328);
nor U2419 (N_2419,N_2260,N_2284);
and U2420 (N_2420,N_2354,N_2347);
and U2421 (N_2421,N_2317,N_2286);
xnor U2422 (N_2422,N_2265,N_2268);
nand U2423 (N_2423,N_2336,N_2369);
or U2424 (N_2424,N_2291,N_2293);
xnor U2425 (N_2425,N_2357,N_2323);
xnor U2426 (N_2426,N_2338,N_2311);
and U2427 (N_2427,N_2299,N_2365);
or U2428 (N_2428,N_2288,N_2371);
or U2429 (N_2429,N_2255,N_2263);
and U2430 (N_2430,N_2321,N_2361);
or U2431 (N_2431,N_2367,N_2266);
and U2432 (N_2432,N_2296,N_2300);
or U2433 (N_2433,N_2346,N_2281);
nand U2434 (N_2434,N_2330,N_2363);
and U2435 (N_2435,N_2273,N_2295);
or U2436 (N_2436,N_2316,N_2283);
and U2437 (N_2437,N_2276,N_2328);
nand U2438 (N_2438,N_2308,N_2251);
or U2439 (N_2439,N_2368,N_2271);
or U2440 (N_2440,N_2358,N_2290);
nor U2441 (N_2441,N_2281,N_2291);
and U2442 (N_2442,N_2295,N_2369);
nor U2443 (N_2443,N_2292,N_2326);
and U2444 (N_2444,N_2251,N_2330);
nor U2445 (N_2445,N_2304,N_2317);
nor U2446 (N_2446,N_2349,N_2365);
or U2447 (N_2447,N_2292,N_2267);
and U2448 (N_2448,N_2274,N_2302);
nor U2449 (N_2449,N_2335,N_2373);
xor U2450 (N_2450,N_2284,N_2371);
and U2451 (N_2451,N_2310,N_2252);
or U2452 (N_2452,N_2260,N_2364);
and U2453 (N_2453,N_2278,N_2269);
or U2454 (N_2454,N_2329,N_2343);
nor U2455 (N_2455,N_2267,N_2262);
nand U2456 (N_2456,N_2277,N_2261);
nand U2457 (N_2457,N_2322,N_2251);
nand U2458 (N_2458,N_2292,N_2296);
xnor U2459 (N_2459,N_2330,N_2333);
nand U2460 (N_2460,N_2334,N_2275);
xor U2461 (N_2461,N_2333,N_2353);
or U2462 (N_2462,N_2332,N_2259);
or U2463 (N_2463,N_2357,N_2259);
or U2464 (N_2464,N_2259,N_2269);
and U2465 (N_2465,N_2280,N_2309);
nor U2466 (N_2466,N_2315,N_2273);
and U2467 (N_2467,N_2371,N_2263);
xnor U2468 (N_2468,N_2252,N_2300);
xor U2469 (N_2469,N_2330,N_2341);
nand U2470 (N_2470,N_2357,N_2271);
and U2471 (N_2471,N_2283,N_2313);
nand U2472 (N_2472,N_2315,N_2258);
xnor U2473 (N_2473,N_2365,N_2295);
xor U2474 (N_2474,N_2264,N_2303);
nor U2475 (N_2475,N_2316,N_2331);
nor U2476 (N_2476,N_2374,N_2307);
nand U2477 (N_2477,N_2302,N_2281);
nor U2478 (N_2478,N_2278,N_2332);
nor U2479 (N_2479,N_2252,N_2360);
nor U2480 (N_2480,N_2337,N_2299);
xor U2481 (N_2481,N_2327,N_2319);
nand U2482 (N_2482,N_2279,N_2293);
and U2483 (N_2483,N_2251,N_2319);
xnor U2484 (N_2484,N_2269,N_2292);
nand U2485 (N_2485,N_2354,N_2255);
nand U2486 (N_2486,N_2266,N_2264);
or U2487 (N_2487,N_2291,N_2342);
or U2488 (N_2488,N_2317,N_2341);
xnor U2489 (N_2489,N_2368,N_2307);
xnor U2490 (N_2490,N_2274,N_2357);
xnor U2491 (N_2491,N_2255,N_2278);
and U2492 (N_2492,N_2362,N_2361);
nand U2493 (N_2493,N_2274,N_2295);
or U2494 (N_2494,N_2328,N_2337);
nand U2495 (N_2495,N_2295,N_2268);
nor U2496 (N_2496,N_2288,N_2271);
nor U2497 (N_2497,N_2351,N_2324);
xnor U2498 (N_2498,N_2370,N_2321);
and U2499 (N_2499,N_2368,N_2302);
and U2500 (N_2500,N_2426,N_2485);
or U2501 (N_2501,N_2440,N_2438);
nand U2502 (N_2502,N_2383,N_2483);
nand U2503 (N_2503,N_2476,N_2436);
xor U2504 (N_2504,N_2478,N_2393);
and U2505 (N_2505,N_2470,N_2451);
xor U2506 (N_2506,N_2437,N_2465);
or U2507 (N_2507,N_2379,N_2499);
nor U2508 (N_2508,N_2433,N_2460);
xnor U2509 (N_2509,N_2377,N_2475);
and U2510 (N_2510,N_2428,N_2402);
and U2511 (N_2511,N_2439,N_2411);
nor U2512 (N_2512,N_2445,N_2444);
nand U2513 (N_2513,N_2482,N_2490);
or U2514 (N_2514,N_2466,N_2446);
nor U2515 (N_2515,N_2409,N_2498);
or U2516 (N_2516,N_2415,N_2418);
nand U2517 (N_2517,N_2421,N_2486);
nand U2518 (N_2518,N_2403,N_2471);
nor U2519 (N_2519,N_2469,N_2462);
nand U2520 (N_2520,N_2396,N_2474);
nor U2521 (N_2521,N_2455,N_2427);
nor U2522 (N_2522,N_2449,N_2401);
nand U2523 (N_2523,N_2480,N_2399);
and U2524 (N_2524,N_2375,N_2441);
or U2525 (N_2525,N_2388,N_2420);
or U2526 (N_2526,N_2477,N_2468);
and U2527 (N_2527,N_2405,N_2452);
nor U2528 (N_2528,N_2395,N_2430);
and U2529 (N_2529,N_2412,N_2435);
xnor U2530 (N_2530,N_2472,N_2484);
nor U2531 (N_2531,N_2389,N_2416);
nor U2532 (N_2532,N_2424,N_2406);
and U2533 (N_2533,N_2419,N_2431);
or U2534 (N_2534,N_2385,N_2456);
nor U2535 (N_2535,N_2453,N_2479);
xnor U2536 (N_2536,N_2454,N_2387);
and U2537 (N_2537,N_2400,N_2378);
or U2538 (N_2538,N_2398,N_2493);
xnor U2539 (N_2539,N_2458,N_2414);
nor U2540 (N_2540,N_2423,N_2467);
nor U2541 (N_2541,N_2390,N_2457);
xnor U2542 (N_2542,N_2450,N_2392);
xnor U2543 (N_2543,N_2381,N_2404);
xor U2544 (N_2544,N_2386,N_2408);
or U2545 (N_2545,N_2487,N_2425);
xor U2546 (N_2546,N_2410,N_2397);
or U2547 (N_2547,N_2394,N_2461);
nor U2548 (N_2548,N_2382,N_2489);
xor U2549 (N_2549,N_2492,N_2407);
or U2550 (N_2550,N_2496,N_2448);
nor U2551 (N_2551,N_2380,N_2417);
xnor U2552 (N_2552,N_2443,N_2429);
or U2553 (N_2553,N_2491,N_2447);
nand U2554 (N_2554,N_2463,N_2481);
or U2555 (N_2555,N_2422,N_2413);
and U2556 (N_2556,N_2497,N_2391);
nand U2557 (N_2557,N_2473,N_2442);
xor U2558 (N_2558,N_2376,N_2432);
nor U2559 (N_2559,N_2494,N_2464);
or U2560 (N_2560,N_2384,N_2459);
and U2561 (N_2561,N_2434,N_2495);
and U2562 (N_2562,N_2488,N_2386);
and U2563 (N_2563,N_2445,N_2377);
nand U2564 (N_2564,N_2437,N_2462);
nor U2565 (N_2565,N_2490,N_2496);
nor U2566 (N_2566,N_2407,N_2382);
nor U2567 (N_2567,N_2499,N_2431);
xnor U2568 (N_2568,N_2414,N_2375);
nand U2569 (N_2569,N_2410,N_2395);
and U2570 (N_2570,N_2496,N_2433);
and U2571 (N_2571,N_2428,N_2396);
xor U2572 (N_2572,N_2450,N_2464);
or U2573 (N_2573,N_2449,N_2426);
or U2574 (N_2574,N_2402,N_2464);
and U2575 (N_2575,N_2388,N_2466);
or U2576 (N_2576,N_2445,N_2378);
nand U2577 (N_2577,N_2487,N_2395);
and U2578 (N_2578,N_2390,N_2441);
nand U2579 (N_2579,N_2386,N_2496);
or U2580 (N_2580,N_2477,N_2486);
nor U2581 (N_2581,N_2395,N_2483);
xor U2582 (N_2582,N_2433,N_2497);
and U2583 (N_2583,N_2481,N_2404);
and U2584 (N_2584,N_2438,N_2419);
nor U2585 (N_2585,N_2392,N_2490);
and U2586 (N_2586,N_2421,N_2464);
xor U2587 (N_2587,N_2478,N_2432);
or U2588 (N_2588,N_2431,N_2469);
or U2589 (N_2589,N_2423,N_2431);
nand U2590 (N_2590,N_2395,N_2432);
or U2591 (N_2591,N_2463,N_2493);
xor U2592 (N_2592,N_2437,N_2449);
or U2593 (N_2593,N_2398,N_2495);
nor U2594 (N_2594,N_2423,N_2384);
and U2595 (N_2595,N_2416,N_2402);
nand U2596 (N_2596,N_2421,N_2450);
xnor U2597 (N_2597,N_2437,N_2429);
nand U2598 (N_2598,N_2409,N_2437);
and U2599 (N_2599,N_2427,N_2385);
and U2600 (N_2600,N_2465,N_2474);
nand U2601 (N_2601,N_2431,N_2409);
nand U2602 (N_2602,N_2382,N_2437);
nor U2603 (N_2603,N_2458,N_2496);
and U2604 (N_2604,N_2459,N_2385);
nand U2605 (N_2605,N_2412,N_2484);
nor U2606 (N_2606,N_2408,N_2409);
or U2607 (N_2607,N_2412,N_2401);
nand U2608 (N_2608,N_2397,N_2496);
nor U2609 (N_2609,N_2438,N_2475);
xor U2610 (N_2610,N_2455,N_2435);
xnor U2611 (N_2611,N_2410,N_2452);
and U2612 (N_2612,N_2425,N_2420);
nand U2613 (N_2613,N_2487,N_2489);
xor U2614 (N_2614,N_2422,N_2407);
nor U2615 (N_2615,N_2428,N_2419);
nand U2616 (N_2616,N_2448,N_2421);
xor U2617 (N_2617,N_2488,N_2437);
nor U2618 (N_2618,N_2431,N_2459);
xnor U2619 (N_2619,N_2437,N_2492);
or U2620 (N_2620,N_2482,N_2403);
nand U2621 (N_2621,N_2385,N_2392);
xnor U2622 (N_2622,N_2453,N_2382);
nor U2623 (N_2623,N_2377,N_2386);
or U2624 (N_2624,N_2381,N_2397);
nand U2625 (N_2625,N_2508,N_2562);
and U2626 (N_2626,N_2545,N_2523);
or U2627 (N_2627,N_2614,N_2548);
and U2628 (N_2628,N_2518,N_2570);
xor U2629 (N_2629,N_2531,N_2500);
nand U2630 (N_2630,N_2506,N_2608);
and U2631 (N_2631,N_2547,N_2576);
nand U2632 (N_2632,N_2596,N_2538);
and U2633 (N_2633,N_2516,N_2615);
nor U2634 (N_2634,N_2619,N_2624);
or U2635 (N_2635,N_2505,N_2607);
nor U2636 (N_2636,N_2620,N_2546);
nand U2637 (N_2637,N_2600,N_2528);
xnor U2638 (N_2638,N_2514,N_2583);
xor U2639 (N_2639,N_2551,N_2550);
and U2640 (N_2640,N_2535,N_2575);
nor U2641 (N_2641,N_2590,N_2557);
xnor U2642 (N_2642,N_2571,N_2527);
and U2643 (N_2643,N_2605,N_2599);
and U2644 (N_2644,N_2542,N_2593);
xnor U2645 (N_2645,N_2517,N_2623);
nor U2646 (N_2646,N_2563,N_2616);
nor U2647 (N_2647,N_2604,N_2578);
nand U2648 (N_2648,N_2553,N_2592);
xor U2649 (N_2649,N_2606,N_2533);
and U2650 (N_2650,N_2552,N_2584);
and U2651 (N_2651,N_2532,N_2618);
nor U2652 (N_2652,N_2511,N_2539);
nor U2653 (N_2653,N_2567,N_2568);
xnor U2654 (N_2654,N_2591,N_2536);
and U2655 (N_2655,N_2502,N_2581);
xnor U2656 (N_2656,N_2587,N_2556);
nor U2657 (N_2657,N_2589,N_2549);
nor U2658 (N_2658,N_2555,N_2519);
and U2659 (N_2659,N_2507,N_2577);
nor U2660 (N_2660,N_2522,N_2530);
xnor U2661 (N_2661,N_2503,N_2534);
nand U2662 (N_2662,N_2595,N_2510);
or U2663 (N_2663,N_2515,N_2540);
nand U2664 (N_2664,N_2504,N_2585);
xnor U2665 (N_2665,N_2579,N_2611);
nor U2666 (N_2666,N_2586,N_2554);
nand U2667 (N_2667,N_2521,N_2565);
nand U2668 (N_2668,N_2512,N_2509);
or U2669 (N_2669,N_2525,N_2582);
xor U2670 (N_2670,N_2559,N_2543);
xor U2671 (N_2671,N_2524,N_2617);
nand U2672 (N_2672,N_2513,N_2602);
nor U2673 (N_2673,N_2613,N_2573);
or U2674 (N_2674,N_2603,N_2537);
xnor U2675 (N_2675,N_2588,N_2580);
or U2676 (N_2676,N_2572,N_2560);
xor U2677 (N_2677,N_2566,N_2501);
nand U2678 (N_2678,N_2544,N_2526);
or U2679 (N_2679,N_2541,N_2564);
and U2680 (N_2680,N_2622,N_2601);
or U2681 (N_2681,N_2574,N_2594);
nor U2682 (N_2682,N_2609,N_2597);
nor U2683 (N_2683,N_2558,N_2529);
xor U2684 (N_2684,N_2598,N_2612);
nor U2685 (N_2685,N_2520,N_2610);
or U2686 (N_2686,N_2569,N_2561);
or U2687 (N_2687,N_2621,N_2531);
or U2688 (N_2688,N_2543,N_2586);
nand U2689 (N_2689,N_2589,N_2618);
nand U2690 (N_2690,N_2570,N_2619);
or U2691 (N_2691,N_2511,N_2506);
and U2692 (N_2692,N_2594,N_2603);
nand U2693 (N_2693,N_2559,N_2508);
and U2694 (N_2694,N_2516,N_2506);
and U2695 (N_2695,N_2572,N_2542);
and U2696 (N_2696,N_2584,N_2542);
xnor U2697 (N_2697,N_2584,N_2530);
and U2698 (N_2698,N_2618,N_2521);
nor U2699 (N_2699,N_2587,N_2521);
or U2700 (N_2700,N_2509,N_2515);
and U2701 (N_2701,N_2566,N_2581);
and U2702 (N_2702,N_2595,N_2591);
and U2703 (N_2703,N_2574,N_2508);
or U2704 (N_2704,N_2519,N_2621);
nor U2705 (N_2705,N_2588,N_2574);
xor U2706 (N_2706,N_2519,N_2502);
and U2707 (N_2707,N_2557,N_2502);
and U2708 (N_2708,N_2582,N_2622);
nor U2709 (N_2709,N_2567,N_2604);
or U2710 (N_2710,N_2542,N_2575);
nand U2711 (N_2711,N_2547,N_2560);
nor U2712 (N_2712,N_2573,N_2557);
xnor U2713 (N_2713,N_2603,N_2619);
xor U2714 (N_2714,N_2564,N_2585);
or U2715 (N_2715,N_2508,N_2577);
xor U2716 (N_2716,N_2567,N_2617);
nor U2717 (N_2717,N_2552,N_2602);
and U2718 (N_2718,N_2552,N_2614);
and U2719 (N_2719,N_2533,N_2527);
nand U2720 (N_2720,N_2582,N_2521);
xor U2721 (N_2721,N_2586,N_2579);
xor U2722 (N_2722,N_2527,N_2509);
and U2723 (N_2723,N_2588,N_2603);
and U2724 (N_2724,N_2592,N_2563);
xnor U2725 (N_2725,N_2514,N_2584);
xnor U2726 (N_2726,N_2574,N_2580);
nand U2727 (N_2727,N_2536,N_2514);
nand U2728 (N_2728,N_2598,N_2543);
nor U2729 (N_2729,N_2526,N_2579);
xnor U2730 (N_2730,N_2616,N_2541);
and U2731 (N_2731,N_2556,N_2552);
nand U2732 (N_2732,N_2550,N_2561);
or U2733 (N_2733,N_2529,N_2578);
nor U2734 (N_2734,N_2500,N_2556);
nand U2735 (N_2735,N_2511,N_2611);
nor U2736 (N_2736,N_2511,N_2518);
xor U2737 (N_2737,N_2519,N_2583);
or U2738 (N_2738,N_2571,N_2555);
nand U2739 (N_2739,N_2610,N_2534);
nand U2740 (N_2740,N_2524,N_2577);
or U2741 (N_2741,N_2526,N_2561);
nor U2742 (N_2742,N_2601,N_2523);
and U2743 (N_2743,N_2506,N_2586);
nor U2744 (N_2744,N_2545,N_2539);
or U2745 (N_2745,N_2596,N_2551);
and U2746 (N_2746,N_2541,N_2531);
and U2747 (N_2747,N_2577,N_2568);
nand U2748 (N_2748,N_2598,N_2602);
nand U2749 (N_2749,N_2505,N_2581);
nor U2750 (N_2750,N_2677,N_2690);
and U2751 (N_2751,N_2682,N_2696);
nor U2752 (N_2752,N_2651,N_2638);
and U2753 (N_2753,N_2704,N_2691);
nand U2754 (N_2754,N_2632,N_2659);
or U2755 (N_2755,N_2683,N_2646);
or U2756 (N_2756,N_2729,N_2667);
and U2757 (N_2757,N_2711,N_2739);
xor U2758 (N_2758,N_2698,N_2745);
and U2759 (N_2759,N_2733,N_2653);
and U2760 (N_2760,N_2658,N_2678);
nand U2761 (N_2761,N_2634,N_2702);
and U2762 (N_2762,N_2717,N_2668);
or U2763 (N_2763,N_2643,N_2661);
nand U2764 (N_2764,N_2660,N_2710);
xor U2765 (N_2765,N_2675,N_2665);
nor U2766 (N_2766,N_2748,N_2712);
nor U2767 (N_2767,N_2656,N_2688);
nor U2768 (N_2768,N_2746,N_2666);
or U2769 (N_2769,N_2727,N_2686);
nand U2770 (N_2770,N_2640,N_2685);
xor U2771 (N_2771,N_2674,N_2743);
and U2772 (N_2772,N_2716,N_2635);
xnor U2773 (N_2773,N_2681,N_2655);
nor U2774 (N_2774,N_2719,N_2722);
nor U2775 (N_2775,N_2676,N_2639);
xnor U2776 (N_2776,N_2664,N_2636);
nor U2777 (N_2777,N_2679,N_2631);
nand U2778 (N_2778,N_2721,N_2709);
xor U2779 (N_2779,N_2648,N_2650);
and U2780 (N_2780,N_2693,N_2687);
xor U2781 (N_2781,N_2713,N_2749);
and U2782 (N_2782,N_2663,N_2708);
nand U2783 (N_2783,N_2652,N_2703);
nand U2784 (N_2784,N_2714,N_2626);
nor U2785 (N_2785,N_2747,N_2705);
or U2786 (N_2786,N_2706,N_2738);
xor U2787 (N_2787,N_2724,N_2697);
nand U2788 (N_2788,N_2673,N_2644);
xor U2789 (N_2789,N_2633,N_2737);
nor U2790 (N_2790,N_2736,N_2642);
xnor U2791 (N_2791,N_2741,N_2728);
nand U2792 (N_2792,N_2700,N_2689);
and U2793 (N_2793,N_2742,N_2699);
or U2794 (N_2794,N_2672,N_2671);
and U2795 (N_2795,N_2641,N_2740);
nand U2796 (N_2796,N_2734,N_2670);
and U2797 (N_2797,N_2630,N_2695);
and U2798 (N_2798,N_2731,N_2718);
nand U2799 (N_2799,N_2735,N_2625);
xnor U2800 (N_2800,N_2715,N_2645);
or U2801 (N_2801,N_2692,N_2725);
nor U2802 (N_2802,N_2628,N_2726);
xor U2803 (N_2803,N_2732,N_2701);
and U2804 (N_2804,N_2649,N_2723);
nand U2805 (N_2805,N_2669,N_2744);
or U2806 (N_2806,N_2720,N_2654);
and U2807 (N_2807,N_2707,N_2629);
or U2808 (N_2808,N_2694,N_2680);
xnor U2809 (N_2809,N_2684,N_2662);
nand U2810 (N_2810,N_2730,N_2627);
or U2811 (N_2811,N_2657,N_2637);
nand U2812 (N_2812,N_2647,N_2733);
or U2813 (N_2813,N_2646,N_2685);
nor U2814 (N_2814,N_2672,N_2652);
and U2815 (N_2815,N_2647,N_2701);
xor U2816 (N_2816,N_2705,N_2733);
xnor U2817 (N_2817,N_2664,N_2717);
and U2818 (N_2818,N_2643,N_2732);
and U2819 (N_2819,N_2667,N_2668);
nor U2820 (N_2820,N_2735,N_2723);
and U2821 (N_2821,N_2731,N_2722);
nand U2822 (N_2822,N_2639,N_2627);
nor U2823 (N_2823,N_2689,N_2675);
nand U2824 (N_2824,N_2706,N_2663);
nand U2825 (N_2825,N_2654,N_2668);
nand U2826 (N_2826,N_2698,N_2670);
nor U2827 (N_2827,N_2716,N_2630);
nor U2828 (N_2828,N_2702,N_2683);
and U2829 (N_2829,N_2745,N_2677);
xnor U2830 (N_2830,N_2705,N_2669);
nand U2831 (N_2831,N_2682,N_2706);
or U2832 (N_2832,N_2739,N_2681);
nand U2833 (N_2833,N_2692,N_2742);
nand U2834 (N_2834,N_2626,N_2648);
nand U2835 (N_2835,N_2668,N_2653);
nand U2836 (N_2836,N_2707,N_2668);
nor U2837 (N_2837,N_2654,N_2714);
and U2838 (N_2838,N_2687,N_2730);
nor U2839 (N_2839,N_2680,N_2683);
or U2840 (N_2840,N_2704,N_2703);
xnor U2841 (N_2841,N_2647,N_2694);
or U2842 (N_2842,N_2706,N_2686);
or U2843 (N_2843,N_2709,N_2656);
and U2844 (N_2844,N_2634,N_2648);
or U2845 (N_2845,N_2648,N_2698);
or U2846 (N_2846,N_2702,N_2649);
or U2847 (N_2847,N_2663,N_2735);
xnor U2848 (N_2848,N_2630,N_2667);
nand U2849 (N_2849,N_2721,N_2658);
xnor U2850 (N_2850,N_2645,N_2688);
and U2851 (N_2851,N_2646,N_2654);
xor U2852 (N_2852,N_2644,N_2639);
and U2853 (N_2853,N_2629,N_2743);
and U2854 (N_2854,N_2702,N_2654);
nand U2855 (N_2855,N_2703,N_2734);
or U2856 (N_2856,N_2646,N_2670);
xor U2857 (N_2857,N_2736,N_2634);
nand U2858 (N_2858,N_2703,N_2717);
nand U2859 (N_2859,N_2633,N_2728);
xnor U2860 (N_2860,N_2716,N_2726);
or U2861 (N_2861,N_2692,N_2696);
and U2862 (N_2862,N_2688,N_2672);
nor U2863 (N_2863,N_2717,N_2732);
and U2864 (N_2864,N_2725,N_2745);
nand U2865 (N_2865,N_2723,N_2715);
or U2866 (N_2866,N_2643,N_2747);
nor U2867 (N_2867,N_2626,N_2630);
or U2868 (N_2868,N_2737,N_2696);
xnor U2869 (N_2869,N_2673,N_2694);
nor U2870 (N_2870,N_2656,N_2633);
or U2871 (N_2871,N_2701,N_2666);
and U2872 (N_2872,N_2679,N_2721);
nor U2873 (N_2873,N_2673,N_2739);
or U2874 (N_2874,N_2659,N_2660);
nand U2875 (N_2875,N_2754,N_2804);
or U2876 (N_2876,N_2861,N_2782);
or U2877 (N_2877,N_2845,N_2850);
and U2878 (N_2878,N_2844,N_2751);
and U2879 (N_2879,N_2866,N_2795);
nand U2880 (N_2880,N_2839,N_2833);
nand U2881 (N_2881,N_2761,N_2788);
xnor U2882 (N_2882,N_2829,N_2811);
xnor U2883 (N_2883,N_2794,N_2780);
nor U2884 (N_2884,N_2825,N_2787);
nor U2885 (N_2885,N_2842,N_2752);
nand U2886 (N_2886,N_2873,N_2853);
xnor U2887 (N_2887,N_2816,N_2789);
or U2888 (N_2888,N_2810,N_2760);
or U2889 (N_2889,N_2874,N_2769);
xor U2890 (N_2890,N_2772,N_2823);
nand U2891 (N_2891,N_2831,N_2854);
and U2892 (N_2892,N_2792,N_2863);
nor U2893 (N_2893,N_2764,N_2791);
and U2894 (N_2894,N_2826,N_2757);
xor U2895 (N_2895,N_2770,N_2828);
nand U2896 (N_2896,N_2836,N_2774);
and U2897 (N_2897,N_2801,N_2835);
nand U2898 (N_2898,N_2777,N_2798);
xor U2899 (N_2899,N_2822,N_2805);
xor U2900 (N_2900,N_2786,N_2864);
nor U2901 (N_2901,N_2750,N_2830);
nor U2902 (N_2902,N_2824,N_2840);
or U2903 (N_2903,N_2753,N_2834);
nor U2904 (N_2904,N_2807,N_2779);
and U2905 (N_2905,N_2775,N_2758);
nand U2906 (N_2906,N_2759,N_2806);
xnor U2907 (N_2907,N_2756,N_2762);
and U2908 (N_2908,N_2859,N_2773);
and U2909 (N_2909,N_2800,N_2838);
nand U2910 (N_2910,N_2778,N_2849);
or U2911 (N_2911,N_2796,N_2808);
nand U2912 (N_2912,N_2776,N_2785);
and U2913 (N_2913,N_2793,N_2818);
xor U2914 (N_2914,N_2765,N_2812);
nand U2915 (N_2915,N_2862,N_2872);
nor U2916 (N_2916,N_2821,N_2848);
xnor U2917 (N_2917,N_2781,N_2809);
and U2918 (N_2918,N_2797,N_2832);
nand U2919 (N_2919,N_2846,N_2766);
nand U2920 (N_2920,N_2819,N_2851);
nor U2921 (N_2921,N_2869,N_2817);
nor U2922 (N_2922,N_2815,N_2870);
nand U2923 (N_2923,N_2820,N_2803);
and U2924 (N_2924,N_2784,N_2799);
xnor U2925 (N_2925,N_2763,N_2814);
or U2926 (N_2926,N_2767,N_2868);
nand U2927 (N_2927,N_2841,N_2813);
or U2928 (N_2928,N_2783,N_2860);
or U2929 (N_2929,N_2865,N_2858);
nand U2930 (N_2930,N_2855,N_2847);
nand U2931 (N_2931,N_2755,N_2768);
nor U2932 (N_2932,N_2856,N_2802);
xor U2933 (N_2933,N_2827,N_2843);
xor U2934 (N_2934,N_2790,N_2857);
and U2935 (N_2935,N_2852,N_2871);
xnor U2936 (N_2936,N_2867,N_2837);
or U2937 (N_2937,N_2771,N_2759);
nand U2938 (N_2938,N_2874,N_2755);
nor U2939 (N_2939,N_2810,N_2787);
xnor U2940 (N_2940,N_2858,N_2843);
nand U2941 (N_2941,N_2870,N_2864);
and U2942 (N_2942,N_2857,N_2812);
nand U2943 (N_2943,N_2858,N_2793);
nor U2944 (N_2944,N_2755,N_2818);
nor U2945 (N_2945,N_2849,N_2798);
nor U2946 (N_2946,N_2872,N_2809);
or U2947 (N_2947,N_2789,N_2874);
or U2948 (N_2948,N_2794,N_2867);
xnor U2949 (N_2949,N_2775,N_2836);
and U2950 (N_2950,N_2776,N_2766);
nor U2951 (N_2951,N_2793,N_2797);
nand U2952 (N_2952,N_2835,N_2757);
or U2953 (N_2953,N_2847,N_2758);
or U2954 (N_2954,N_2822,N_2811);
and U2955 (N_2955,N_2847,N_2816);
nor U2956 (N_2956,N_2762,N_2869);
nand U2957 (N_2957,N_2821,N_2771);
nand U2958 (N_2958,N_2786,N_2874);
nand U2959 (N_2959,N_2803,N_2855);
xnor U2960 (N_2960,N_2850,N_2840);
and U2961 (N_2961,N_2855,N_2817);
nor U2962 (N_2962,N_2818,N_2751);
xnor U2963 (N_2963,N_2811,N_2861);
xnor U2964 (N_2964,N_2778,N_2804);
nor U2965 (N_2965,N_2768,N_2854);
or U2966 (N_2966,N_2819,N_2780);
xnor U2967 (N_2967,N_2814,N_2803);
nand U2968 (N_2968,N_2760,N_2804);
xor U2969 (N_2969,N_2756,N_2830);
nand U2970 (N_2970,N_2824,N_2816);
nor U2971 (N_2971,N_2797,N_2848);
or U2972 (N_2972,N_2829,N_2752);
nor U2973 (N_2973,N_2835,N_2802);
nand U2974 (N_2974,N_2865,N_2768);
xnor U2975 (N_2975,N_2803,N_2848);
xnor U2976 (N_2976,N_2819,N_2778);
nand U2977 (N_2977,N_2763,N_2770);
xor U2978 (N_2978,N_2754,N_2794);
or U2979 (N_2979,N_2864,N_2773);
nor U2980 (N_2980,N_2873,N_2752);
xor U2981 (N_2981,N_2838,N_2794);
nand U2982 (N_2982,N_2774,N_2817);
nor U2983 (N_2983,N_2753,N_2751);
nand U2984 (N_2984,N_2782,N_2815);
xor U2985 (N_2985,N_2827,N_2750);
nor U2986 (N_2986,N_2859,N_2870);
nand U2987 (N_2987,N_2861,N_2844);
nor U2988 (N_2988,N_2839,N_2807);
or U2989 (N_2989,N_2866,N_2750);
and U2990 (N_2990,N_2801,N_2863);
or U2991 (N_2991,N_2771,N_2756);
xnor U2992 (N_2992,N_2757,N_2771);
or U2993 (N_2993,N_2873,N_2766);
xor U2994 (N_2994,N_2783,N_2789);
nor U2995 (N_2995,N_2803,N_2815);
nor U2996 (N_2996,N_2839,N_2789);
nor U2997 (N_2997,N_2843,N_2874);
nor U2998 (N_2998,N_2867,N_2871);
xor U2999 (N_2999,N_2817,N_2861);
xor U3000 (N_3000,N_2878,N_2931);
nor U3001 (N_3001,N_2921,N_2894);
and U3002 (N_3002,N_2987,N_2900);
and U3003 (N_3003,N_2940,N_2984);
nor U3004 (N_3004,N_2957,N_2893);
xor U3005 (N_3005,N_2920,N_2917);
nor U3006 (N_3006,N_2967,N_2899);
xor U3007 (N_3007,N_2929,N_2932);
nor U3008 (N_3008,N_2948,N_2960);
nor U3009 (N_3009,N_2946,N_2980);
nor U3010 (N_3010,N_2947,N_2989);
nand U3011 (N_3011,N_2964,N_2901);
or U3012 (N_3012,N_2965,N_2949);
nand U3013 (N_3013,N_2945,N_2936);
or U3014 (N_3014,N_2919,N_2950);
nand U3015 (N_3015,N_2876,N_2886);
xnor U3016 (N_3016,N_2885,N_2986);
nor U3017 (N_3017,N_2913,N_2963);
xor U3018 (N_3018,N_2959,N_2882);
xnor U3019 (N_3019,N_2978,N_2916);
and U3020 (N_3020,N_2981,N_2969);
or U3021 (N_3021,N_2970,N_2897);
and U3022 (N_3022,N_2937,N_2976);
nand U3023 (N_3023,N_2995,N_2880);
xor U3024 (N_3024,N_2889,N_2892);
or U3025 (N_3025,N_2962,N_2942);
nand U3026 (N_3026,N_2908,N_2982);
or U3027 (N_3027,N_2972,N_2915);
xor U3028 (N_3028,N_2879,N_2891);
or U3029 (N_3029,N_2961,N_2890);
or U3030 (N_3030,N_2906,N_2991);
nand U3031 (N_3031,N_2926,N_2924);
nor U3032 (N_3032,N_2910,N_2895);
nand U3033 (N_3033,N_2943,N_2994);
or U3034 (N_3034,N_2914,N_2912);
nor U3035 (N_3035,N_2934,N_2883);
xnor U3036 (N_3036,N_2938,N_2907);
or U3037 (N_3037,N_2977,N_2918);
xnor U3038 (N_3038,N_2998,N_2888);
xor U3039 (N_3039,N_2979,N_2958);
nand U3040 (N_3040,N_2898,N_2975);
nor U3041 (N_3041,N_2992,N_2930);
nand U3042 (N_3042,N_2935,N_2974);
xnor U3043 (N_3043,N_2996,N_2955);
nor U3044 (N_3044,N_2971,N_2922);
xor U3045 (N_3045,N_2884,N_2966);
nand U3046 (N_3046,N_2952,N_2983);
nor U3047 (N_3047,N_2896,N_2881);
nand U3048 (N_3048,N_2928,N_2904);
nor U3049 (N_3049,N_2956,N_2903);
nor U3050 (N_3050,N_2973,N_2990);
and U3051 (N_3051,N_2939,N_2911);
nand U3052 (N_3052,N_2951,N_2941);
nand U3053 (N_3053,N_2925,N_2988);
and U3054 (N_3054,N_2909,N_2902);
nor U3055 (N_3055,N_2999,N_2985);
and U3056 (N_3056,N_2877,N_2927);
xor U3057 (N_3057,N_2933,N_2905);
nand U3058 (N_3058,N_2944,N_2923);
or U3059 (N_3059,N_2887,N_2953);
nand U3060 (N_3060,N_2997,N_2968);
and U3061 (N_3061,N_2954,N_2993);
nand U3062 (N_3062,N_2875,N_2961);
nand U3063 (N_3063,N_2974,N_2890);
or U3064 (N_3064,N_2942,N_2907);
xnor U3065 (N_3065,N_2922,N_2997);
or U3066 (N_3066,N_2925,N_2975);
and U3067 (N_3067,N_2979,N_2899);
nand U3068 (N_3068,N_2958,N_2935);
xor U3069 (N_3069,N_2930,N_2978);
xnor U3070 (N_3070,N_2936,N_2926);
nor U3071 (N_3071,N_2982,N_2922);
nand U3072 (N_3072,N_2927,N_2876);
or U3073 (N_3073,N_2964,N_2929);
xor U3074 (N_3074,N_2917,N_2905);
xnor U3075 (N_3075,N_2959,N_2954);
and U3076 (N_3076,N_2920,N_2951);
xor U3077 (N_3077,N_2906,N_2929);
and U3078 (N_3078,N_2967,N_2905);
xnor U3079 (N_3079,N_2876,N_2972);
or U3080 (N_3080,N_2881,N_2966);
and U3081 (N_3081,N_2936,N_2928);
xnor U3082 (N_3082,N_2923,N_2920);
nand U3083 (N_3083,N_2924,N_2887);
nor U3084 (N_3084,N_2999,N_2879);
nor U3085 (N_3085,N_2876,N_2922);
xor U3086 (N_3086,N_2991,N_2968);
nand U3087 (N_3087,N_2998,N_2963);
xor U3088 (N_3088,N_2993,N_2989);
nand U3089 (N_3089,N_2899,N_2926);
nor U3090 (N_3090,N_2960,N_2888);
xor U3091 (N_3091,N_2927,N_2875);
nor U3092 (N_3092,N_2983,N_2964);
xnor U3093 (N_3093,N_2974,N_2960);
nor U3094 (N_3094,N_2880,N_2881);
or U3095 (N_3095,N_2946,N_2970);
or U3096 (N_3096,N_2955,N_2969);
or U3097 (N_3097,N_2880,N_2952);
nor U3098 (N_3098,N_2910,N_2974);
or U3099 (N_3099,N_2949,N_2907);
nor U3100 (N_3100,N_2901,N_2878);
and U3101 (N_3101,N_2911,N_2920);
nor U3102 (N_3102,N_2984,N_2986);
nand U3103 (N_3103,N_2948,N_2902);
or U3104 (N_3104,N_2912,N_2945);
nand U3105 (N_3105,N_2960,N_2966);
or U3106 (N_3106,N_2950,N_2905);
xor U3107 (N_3107,N_2966,N_2969);
xor U3108 (N_3108,N_2883,N_2937);
or U3109 (N_3109,N_2956,N_2997);
nor U3110 (N_3110,N_2987,N_2982);
nand U3111 (N_3111,N_2938,N_2875);
xor U3112 (N_3112,N_2957,N_2907);
nand U3113 (N_3113,N_2958,N_2999);
xor U3114 (N_3114,N_2891,N_2907);
nand U3115 (N_3115,N_2944,N_2913);
nand U3116 (N_3116,N_2895,N_2963);
xor U3117 (N_3117,N_2902,N_2934);
nor U3118 (N_3118,N_2926,N_2878);
or U3119 (N_3119,N_2897,N_2925);
xor U3120 (N_3120,N_2924,N_2984);
or U3121 (N_3121,N_2992,N_2929);
or U3122 (N_3122,N_2875,N_2934);
nor U3123 (N_3123,N_2875,N_2944);
xor U3124 (N_3124,N_2924,N_2946);
xor U3125 (N_3125,N_3091,N_3009);
or U3126 (N_3126,N_3064,N_3078);
nor U3127 (N_3127,N_3111,N_3006);
and U3128 (N_3128,N_3096,N_3025);
or U3129 (N_3129,N_3075,N_3116);
and U3130 (N_3130,N_3060,N_3080);
and U3131 (N_3131,N_3093,N_3123);
xnor U3132 (N_3132,N_3014,N_3110);
nand U3133 (N_3133,N_3054,N_3021);
or U3134 (N_3134,N_3092,N_3115);
or U3135 (N_3135,N_3073,N_3070);
nand U3136 (N_3136,N_3055,N_3047);
xnor U3137 (N_3137,N_3012,N_3121);
nor U3138 (N_3138,N_3068,N_3119);
nor U3139 (N_3139,N_3077,N_3035);
or U3140 (N_3140,N_3086,N_3007);
nand U3141 (N_3141,N_3005,N_3108);
xnor U3142 (N_3142,N_3113,N_3114);
or U3143 (N_3143,N_3087,N_3066);
and U3144 (N_3144,N_3106,N_3027);
and U3145 (N_3145,N_3122,N_3008);
or U3146 (N_3146,N_3024,N_3118);
or U3147 (N_3147,N_3028,N_3015);
or U3148 (N_3148,N_3090,N_3053);
nor U3149 (N_3149,N_3112,N_3098);
nor U3150 (N_3150,N_3022,N_3082);
and U3151 (N_3151,N_3065,N_3019);
and U3152 (N_3152,N_3020,N_3044);
xor U3153 (N_3153,N_3050,N_3029);
xnor U3154 (N_3154,N_3079,N_3051);
nand U3155 (N_3155,N_3059,N_3081);
or U3156 (N_3156,N_3036,N_3109);
xor U3157 (N_3157,N_3001,N_3084);
nand U3158 (N_3158,N_3107,N_3041);
nand U3159 (N_3159,N_3105,N_3103);
and U3160 (N_3160,N_3018,N_3076);
nor U3161 (N_3161,N_3061,N_3083);
xnor U3162 (N_3162,N_3045,N_3069);
xor U3163 (N_3163,N_3048,N_3101);
nand U3164 (N_3164,N_3004,N_3002);
nand U3165 (N_3165,N_3052,N_3095);
or U3166 (N_3166,N_3000,N_3039);
and U3167 (N_3167,N_3062,N_3037);
or U3168 (N_3168,N_3030,N_3034);
xor U3169 (N_3169,N_3031,N_3120);
xor U3170 (N_3170,N_3057,N_3011);
nand U3171 (N_3171,N_3074,N_3032);
or U3172 (N_3172,N_3058,N_3056);
and U3173 (N_3173,N_3072,N_3042);
nor U3174 (N_3174,N_3099,N_3016);
xnor U3175 (N_3175,N_3023,N_3063);
or U3176 (N_3176,N_3089,N_3043);
nor U3177 (N_3177,N_3038,N_3117);
nand U3178 (N_3178,N_3033,N_3071);
and U3179 (N_3179,N_3124,N_3049);
xnor U3180 (N_3180,N_3097,N_3013);
nor U3181 (N_3181,N_3040,N_3100);
or U3182 (N_3182,N_3088,N_3010);
xor U3183 (N_3183,N_3085,N_3094);
and U3184 (N_3184,N_3046,N_3102);
and U3185 (N_3185,N_3026,N_3067);
and U3186 (N_3186,N_3104,N_3017);
nor U3187 (N_3187,N_3003,N_3015);
and U3188 (N_3188,N_3093,N_3051);
and U3189 (N_3189,N_3080,N_3014);
or U3190 (N_3190,N_3079,N_3052);
xnor U3191 (N_3191,N_3061,N_3012);
or U3192 (N_3192,N_3069,N_3122);
xor U3193 (N_3193,N_3110,N_3056);
nand U3194 (N_3194,N_3079,N_3036);
and U3195 (N_3195,N_3109,N_3053);
and U3196 (N_3196,N_3092,N_3079);
nor U3197 (N_3197,N_3067,N_3096);
and U3198 (N_3198,N_3119,N_3046);
nor U3199 (N_3199,N_3058,N_3021);
or U3200 (N_3200,N_3055,N_3040);
xnor U3201 (N_3201,N_3092,N_3094);
nand U3202 (N_3202,N_3100,N_3008);
xnor U3203 (N_3203,N_3037,N_3097);
and U3204 (N_3204,N_3114,N_3076);
and U3205 (N_3205,N_3050,N_3120);
and U3206 (N_3206,N_3097,N_3066);
nand U3207 (N_3207,N_3116,N_3034);
nand U3208 (N_3208,N_3082,N_3105);
nand U3209 (N_3209,N_3053,N_3093);
xnor U3210 (N_3210,N_3075,N_3042);
or U3211 (N_3211,N_3113,N_3037);
or U3212 (N_3212,N_3090,N_3001);
nor U3213 (N_3213,N_3003,N_3028);
xnor U3214 (N_3214,N_3089,N_3039);
or U3215 (N_3215,N_3070,N_3029);
or U3216 (N_3216,N_3039,N_3074);
or U3217 (N_3217,N_3101,N_3002);
nand U3218 (N_3218,N_3043,N_3030);
and U3219 (N_3219,N_3015,N_3066);
or U3220 (N_3220,N_3081,N_3026);
and U3221 (N_3221,N_3111,N_3106);
or U3222 (N_3222,N_3074,N_3108);
nor U3223 (N_3223,N_3061,N_3009);
nor U3224 (N_3224,N_3080,N_3089);
or U3225 (N_3225,N_3019,N_3047);
or U3226 (N_3226,N_3120,N_3097);
xor U3227 (N_3227,N_3083,N_3114);
or U3228 (N_3228,N_3023,N_3120);
and U3229 (N_3229,N_3059,N_3087);
nand U3230 (N_3230,N_3002,N_3008);
xnor U3231 (N_3231,N_3082,N_3120);
nor U3232 (N_3232,N_3008,N_3048);
nor U3233 (N_3233,N_3043,N_3034);
and U3234 (N_3234,N_3071,N_3025);
nand U3235 (N_3235,N_3036,N_3083);
or U3236 (N_3236,N_3053,N_3051);
nor U3237 (N_3237,N_3012,N_3086);
nand U3238 (N_3238,N_3100,N_3006);
nor U3239 (N_3239,N_3111,N_3058);
nand U3240 (N_3240,N_3063,N_3067);
nand U3241 (N_3241,N_3072,N_3011);
xor U3242 (N_3242,N_3048,N_3024);
nand U3243 (N_3243,N_3091,N_3008);
and U3244 (N_3244,N_3106,N_3089);
xor U3245 (N_3245,N_3084,N_3058);
nand U3246 (N_3246,N_3003,N_3023);
nor U3247 (N_3247,N_3011,N_3036);
nand U3248 (N_3248,N_3109,N_3070);
xnor U3249 (N_3249,N_3033,N_3063);
and U3250 (N_3250,N_3146,N_3197);
nor U3251 (N_3251,N_3224,N_3211);
and U3252 (N_3252,N_3132,N_3154);
nand U3253 (N_3253,N_3246,N_3171);
xor U3254 (N_3254,N_3240,N_3173);
and U3255 (N_3255,N_3182,N_3198);
nand U3256 (N_3256,N_3205,N_3125);
nor U3257 (N_3257,N_3166,N_3190);
nand U3258 (N_3258,N_3201,N_3141);
nor U3259 (N_3259,N_3143,N_3175);
or U3260 (N_3260,N_3239,N_3229);
xor U3261 (N_3261,N_3207,N_3153);
or U3262 (N_3262,N_3161,N_3232);
or U3263 (N_3263,N_3218,N_3188);
and U3264 (N_3264,N_3204,N_3168);
xnor U3265 (N_3265,N_3227,N_3178);
xnor U3266 (N_3266,N_3128,N_3158);
nand U3267 (N_3267,N_3219,N_3160);
xnor U3268 (N_3268,N_3247,N_3234);
and U3269 (N_3269,N_3170,N_3223);
xor U3270 (N_3270,N_3163,N_3216);
nor U3271 (N_3271,N_3226,N_3186);
or U3272 (N_3272,N_3157,N_3194);
xnor U3273 (N_3273,N_3235,N_3209);
xor U3274 (N_3274,N_3195,N_3180);
and U3275 (N_3275,N_3133,N_3220);
nor U3276 (N_3276,N_3185,N_3245);
nand U3277 (N_3277,N_3184,N_3215);
or U3278 (N_3278,N_3203,N_3155);
xor U3279 (N_3279,N_3202,N_3244);
and U3280 (N_3280,N_3248,N_3151);
and U3281 (N_3281,N_3149,N_3127);
and U3282 (N_3282,N_3136,N_3243);
and U3283 (N_3283,N_3144,N_3200);
and U3284 (N_3284,N_3181,N_3213);
nor U3285 (N_3285,N_3162,N_3165);
nand U3286 (N_3286,N_3169,N_3238);
nand U3287 (N_3287,N_3130,N_3191);
nand U3288 (N_3288,N_3129,N_3152);
or U3289 (N_3289,N_3164,N_3176);
or U3290 (N_3290,N_3249,N_3131);
or U3291 (N_3291,N_3208,N_3199);
or U3292 (N_3292,N_3183,N_3138);
and U3293 (N_3293,N_3193,N_3189);
and U3294 (N_3294,N_3214,N_3135);
nor U3295 (N_3295,N_3196,N_3137);
and U3296 (N_3296,N_3126,N_3222);
and U3297 (N_3297,N_3221,N_3187);
xor U3298 (N_3298,N_3172,N_3241);
nor U3299 (N_3299,N_3167,N_3242);
nor U3300 (N_3300,N_3233,N_3142);
or U3301 (N_3301,N_3159,N_3236);
and U3302 (N_3302,N_3192,N_3148);
nand U3303 (N_3303,N_3179,N_3134);
xnor U3304 (N_3304,N_3210,N_3139);
or U3305 (N_3305,N_3212,N_3147);
nand U3306 (N_3306,N_3230,N_3156);
nor U3307 (N_3307,N_3174,N_3217);
nor U3308 (N_3308,N_3150,N_3237);
xnor U3309 (N_3309,N_3145,N_3231);
xor U3310 (N_3310,N_3228,N_3225);
nor U3311 (N_3311,N_3140,N_3177);
nor U3312 (N_3312,N_3206,N_3217);
nand U3313 (N_3313,N_3210,N_3166);
or U3314 (N_3314,N_3194,N_3161);
nand U3315 (N_3315,N_3142,N_3160);
nor U3316 (N_3316,N_3125,N_3221);
nand U3317 (N_3317,N_3210,N_3175);
nand U3318 (N_3318,N_3167,N_3237);
xor U3319 (N_3319,N_3185,N_3186);
nand U3320 (N_3320,N_3159,N_3129);
nor U3321 (N_3321,N_3225,N_3183);
nand U3322 (N_3322,N_3235,N_3185);
nor U3323 (N_3323,N_3125,N_3235);
and U3324 (N_3324,N_3194,N_3137);
and U3325 (N_3325,N_3161,N_3143);
nand U3326 (N_3326,N_3168,N_3218);
or U3327 (N_3327,N_3170,N_3235);
nor U3328 (N_3328,N_3132,N_3202);
xnor U3329 (N_3329,N_3200,N_3172);
and U3330 (N_3330,N_3184,N_3213);
xnor U3331 (N_3331,N_3139,N_3154);
nand U3332 (N_3332,N_3178,N_3161);
and U3333 (N_3333,N_3182,N_3223);
and U3334 (N_3334,N_3130,N_3159);
nand U3335 (N_3335,N_3166,N_3240);
nor U3336 (N_3336,N_3238,N_3186);
nand U3337 (N_3337,N_3246,N_3213);
nand U3338 (N_3338,N_3141,N_3166);
or U3339 (N_3339,N_3235,N_3202);
or U3340 (N_3340,N_3234,N_3192);
xnor U3341 (N_3341,N_3241,N_3240);
or U3342 (N_3342,N_3180,N_3196);
nand U3343 (N_3343,N_3153,N_3225);
xnor U3344 (N_3344,N_3170,N_3133);
xnor U3345 (N_3345,N_3158,N_3141);
or U3346 (N_3346,N_3203,N_3213);
xnor U3347 (N_3347,N_3180,N_3125);
nand U3348 (N_3348,N_3234,N_3175);
nand U3349 (N_3349,N_3161,N_3184);
nor U3350 (N_3350,N_3243,N_3138);
nand U3351 (N_3351,N_3241,N_3136);
nand U3352 (N_3352,N_3212,N_3235);
and U3353 (N_3353,N_3185,N_3136);
xor U3354 (N_3354,N_3167,N_3158);
nand U3355 (N_3355,N_3237,N_3134);
nand U3356 (N_3356,N_3232,N_3150);
nor U3357 (N_3357,N_3192,N_3161);
or U3358 (N_3358,N_3231,N_3244);
xor U3359 (N_3359,N_3170,N_3182);
or U3360 (N_3360,N_3198,N_3185);
nand U3361 (N_3361,N_3185,N_3240);
or U3362 (N_3362,N_3178,N_3209);
xnor U3363 (N_3363,N_3138,N_3141);
nor U3364 (N_3364,N_3176,N_3230);
or U3365 (N_3365,N_3192,N_3217);
nand U3366 (N_3366,N_3158,N_3191);
nand U3367 (N_3367,N_3209,N_3210);
or U3368 (N_3368,N_3234,N_3125);
xnor U3369 (N_3369,N_3213,N_3234);
xnor U3370 (N_3370,N_3226,N_3246);
nand U3371 (N_3371,N_3177,N_3126);
nand U3372 (N_3372,N_3231,N_3154);
nand U3373 (N_3373,N_3216,N_3147);
or U3374 (N_3374,N_3192,N_3238);
xnor U3375 (N_3375,N_3257,N_3253);
and U3376 (N_3376,N_3347,N_3298);
nand U3377 (N_3377,N_3269,N_3301);
and U3378 (N_3378,N_3280,N_3285);
nor U3379 (N_3379,N_3361,N_3288);
xnor U3380 (N_3380,N_3362,N_3329);
nand U3381 (N_3381,N_3279,N_3357);
nor U3382 (N_3382,N_3354,N_3311);
nand U3383 (N_3383,N_3322,N_3369);
and U3384 (N_3384,N_3368,N_3272);
nor U3385 (N_3385,N_3268,N_3295);
xor U3386 (N_3386,N_3303,N_3328);
or U3387 (N_3387,N_3313,N_3348);
xnor U3388 (N_3388,N_3330,N_3270);
nor U3389 (N_3389,N_3259,N_3349);
xor U3390 (N_3390,N_3296,N_3315);
nand U3391 (N_3391,N_3281,N_3343);
nor U3392 (N_3392,N_3340,N_3353);
xor U3393 (N_3393,N_3364,N_3317);
nor U3394 (N_3394,N_3358,N_3284);
nor U3395 (N_3395,N_3351,N_3250);
or U3396 (N_3396,N_3256,N_3338);
or U3397 (N_3397,N_3307,N_3318);
nor U3398 (N_3398,N_3350,N_3275);
nand U3399 (N_3399,N_3314,N_3255);
and U3400 (N_3400,N_3286,N_3297);
and U3401 (N_3401,N_3344,N_3370);
nor U3402 (N_3402,N_3302,N_3282);
xor U3403 (N_3403,N_3372,N_3291);
nor U3404 (N_3404,N_3326,N_3304);
nand U3405 (N_3405,N_3287,N_3316);
xor U3406 (N_3406,N_3345,N_3331);
nand U3407 (N_3407,N_3312,N_3262);
and U3408 (N_3408,N_3327,N_3320);
or U3409 (N_3409,N_3306,N_3373);
xnor U3410 (N_3410,N_3271,N_3360);
and U3411 (N_3411,N_3337,N_3352);
and U3412 (N_3412,N_3323,N_3371);
or U3413 (N_3413,N_3277,N_3254);
nor U3414 (N_3414,N_3265,N_3258);
and U3415 (N_3415,N_3273,N_3332);
nand U3416 (N_3416,N_3252,N_3283);
and U3417 (N_3417,N_3251,N_3319);
nor U3418 (N_3418,N_3335,N_3299);
nand U3419 (N_3419,N_3374,N_3276);
nor U3420 (N_3420,N_3324,N_3278);
or U3421 (N_3421,N_3359,N_3300);
nand U3422 (N_3422,N_3274,N_3321);
or U3423 (N_3423,N_3336,N_3305);
and U3424 (N_3424,N_3261,N_3310);
or U3425 (N_3425,N_3293,N_3341);
and U3426 (N_3426,N_3292,N_3325);
or U3427 (N_3427,N_3289,N_3366);
xor U3428 (N_3428,N_3266,N_3356);
and U3429 (N_3429,N_3290,N_3308);
nor U3430 (N_3430,N_3333,N_3264);
xnor U3431 (N_3431,N_3339,N_3355);
nand U3432 (N_3432,N_3334,N_3263);
nand U3433 (N_3433,N_3342,N_3367);
nand U3434 (N_3434,N_3346,N_3363);
nand U3435 (N_3435,N_3260,N_3267);
nand U3436 (N_3436,N_3294,N_3365);
and U3437 (N_3437,N_3309,N_3324);
and U3438 (N_3438,N_3312,N_3335);
nand U3439 (N_3439,N_3364,N_3360);
nand U3440 (N_3440,N_3353,N_3299);
and U3441 (N_3441,N_3273,N_3363);
or U3442 (N_3442,N_3265,N_3372);
and U3443 (N_3443,N_3318,N_3364);
or U3444 (N_3444,N_3323,N_3293);
nor U3445 (N_3445,N_3356,N_3343);
nand U3446 (N_3446,N_3274,N_3275);
xnor U3447 (N_3447,N_3326,N_3275);
nor U3448 (N_3448,N_3358,N_3257);
xor U3449 (N_3449,N_3354,N_3258);
nand U3450 (N_3450,N_3291,N_3363);
and U3451 (N_3451,N_3372,N_3293);
nor U3452 (N_3452,N_3264,N_3368);
xnor U3453 (N_3453,N_3373,N_3316);
nor U3454 (N_3454,N_3302,N_3265);
xnor U3455 (N_3455,N_3353,N_3294);
or U3456 (N_3456,N_3298,N_3344);
and U3457 (N_3457,N_3308,N_3363);
xnor U3458 (N_3458,N_3362,N_3330);
or U3459 (N_3459,N_3352,N_3280);
nor U3460 (N_3460,N_3352,N_3371);
nand U3461 (N_3461,N_3347,N_3327);
and U3462 (N_3462,N_3288,N_3312);
nor U3463 (N_3463,N_3334,N_3282);
and U3464 (N_3464,N_3352,N_3296);
and U3465 (N_3465,N_3330,N_3258);
xnor U3466 (N_3466,N_3311,N_3321);
nand U3467 (N_3467,N_3356,N_3310);
and U3468 (N_3468,N_3315,N_3348);
nand U3469 (N_3469,N_3340,N_3287);
nor U3470 (N_3470,N_3343,N_3292);
and U3471 (N_3471,N_3372,N_3281);
and U3472 (N_3472,N_3319,N_3264);
nor U3473 (N_3473,N_3293,N_3307);
and U3474 (N_3474,N_3253,N_3340);
nor U3475 (N_3475,N_3299,N_3268);
and U3476 (N_3476,N_3281,N_3254);
xnor U3477 (N_3477,N_3278,N_3334);
and U3478 (N_3478,N_3267,N_3359);
nor U3479 (N_3479,N_3346,N_3290);
xnor U3480 (N_3480,N_3295,N_3357);
xor U3481 (N_3481,N_3277,N_3252);
or U3482 (N_3482,N_3269,N_3274);
or U3483 (N_3483,N_3369,N_3329);
or U3484 (N_3484,N_3258,N_3305);
nand U3485 (N_3485,N_3329,N_3294);
xor U3486 (N_3486,N_3257,N_3342);
nor U3487 (N_3487,N_3315,N_3317);
xnor U3488 (N_3488,N_3368,N_3344);
and U3489 (N_3489,N_3321,N_3316);
or U3490 (N_3490,N_3343,N_3266);
nor U3491 (N_3491,N_3353,N_3281);
nor U3492 (N_3492,N_3309,N_3342);
nand U3493 (N_3493,N_3292,N_3271);
and U3494 (N_3494,N_3295,N_3335);
or U3495 (N_3495,N_3289,N_3267);
nand U3496 (N_3496,N_3319,N_3307);
nor U3497 (N_3497,N_3288,N_3348);
xor U3498 (N_3498,N_3355,N_3250);
and U3499 (N_3499,N_3370,N_3254);
and U3500 (N_3500,N_3481,N_3454);
and U3501 (N_3501,N_3487,N_3485);
and U3502 (N_3502,N_3443,N_3422);
xnor U3503 (N_3503,N_3465,N_3471);
and U3504 (N_3504,N_3382,N_3403);
and U3505 (N_3505,N_3461,N_3408);
and U3506 (N_3506,N_3464,N_3463);
xnor U3507 (N_3507,N_3375,N_3387);
nand U3508 (N_3508,N_3415,N_3386);
xnor U3509 (N_3509,N_3409,N_3429);
and U3510 (N_3510,N_3434,N_3383);
or U3511 (N_3511,N_3445,N_3446);
and U3512 (N_3512,N_3482,N_3380);
xnor U3513 (N_3513,N_3489,N_3458);
or U3514 (N_3514,N_3427,N_3433);
or U3515 (N_3515,N_3478,N_3448);
nand U3516 (N_3516,N_3394,N_3431);
and U3517 (N_3517,N_3395,N_3411);
nor U3518 (N_3518,N_3494,N_3412);
and U3519 (N_3519,N_3451,N_3444);
nand U3520 (N_3520,N_3417,N_3496);
nor U3521 (N_3521,N_3376,N_3447);
nand U3522 (N_3522,N_3384,N_3421);
nand U3523 (N_3523,N_3459,N_3406);
nor U3524 (N_3524,N_3484,N_3392);
nor U3525 (N_3525,N_3476,N_3390);
nand U3526 (N_3526,N_3493,N_3396);
or U3527 (N_3527,N_3450,N_3407);
xor U3528 (N_3528,N_3405,N_3460);
nand U3529 (N_3529,N_3470,N_3455);
xnor U3530 (N_3530,N_3379,N_3440);
xnor U3531 (N_3531,N_3400,N_3410);
and U3532 (N_3532,N_3377,N_3483);
nor U3533 (N_3533,N_3488,N_3449);
nor U3534 (N_3534,N_3420,N_3381);
and U3535 (N_3535,N_3438,N_3462);
nor U3536 (N_3536,N_3441,N_3495);
nand U3537 (N_3537,N_3436,N_3423);
xnor U3538 (N_3538,N_3418,N_3413);
or U3539 (N_3539,N_3479,N_3472);
or U3540 (N_3540,N_3442,N_3480);
nor U3541 (N_3541,N_3416,N_3498);
nor U3542 (N_3542,N_3397,N_3477);
nor U3543 (N_3543,N_3457,N_3486);
nor U3544 (N_3544,N_3492,N_3424);
xnor U3545 (N_3545,N_3389,N_3466);
nand U3546 (N_3546,N_3391,N_3414);
or U3547 (N_3547,N_3378,N_3419);
xor U3548 (N_3548,N_3393,N_3497);
nand U3549 (N_3549,N_3398,N_3467);
nor U3550 (N_3550,N_3435,N_3428);
xnor U3551 (N_3551,N_3453,N_3388);
xnor U3552 (N_3552,N_3437,N_3491);
nand U3553 (N_3553,N_3402,N_3404);
xnor U3554 (N_3554,N_3425,N_3468);
nor U3555 (N_3555,N_3499,N_3452);
nand U3556 (N_3556,N_3432,N_3473);
nor U3557 (N_3557,N_3385,N_3430);
and U3558 (N_3558,N_3456,N_3399);
and U3559 (N_3559,N_3490,N_3474);
nor U3560 (N_3560,N_3439,N_3475);
nor U3561 (N_3561,N_3469,N_3401);
nand U3562 (N_3562,N_3426,N_3448);
xor U3563 (N_3563,N_3382,N_3465);
nor U3564 (N_3564,N_3430,N_3401);
nand U3565 (N_3565,N_3429,N_3431);
or U3566 (N_3566,N_3441,N_3458);
nand U3567 (N_3567,N_3402,N_3467);
nor U3568 (N_3568,N_3481,N_3380);
xnor U3569 (N_3569,N_3483,N_3496);
or U3570 (N_3570,N_3473,N_3386);
xor U3571 (N_3571,N_3482,N_3477);
xnor U3572 (N_3572,N_3445,N_3429);
and U3573 (N_3573,N_3435,N_3489);
or U3574 (N_3574,N_3451,N_3462);
or U3575 (N_3575,N_3409,N_3441);
xnor U3576 (N_3576,N_3414,N_3380);
or U3577 (N_3577,N_3457,N_3463);
nand U3578 (N_3578,N_3381,N_3493);
nor U3579 (N_3579,N_3414,N_3431);
nand U3580 (N_3580,N_3383,N_3446);
and U3581 (N_3581,N_3470,N_3401);
nor U3582 (N_3582,N_3432,N_3472);
nand U3583 (N_3583,N_3385,N_3375);
nor U3584 (N_3584,N_3387,N_3384);
xor U3585 (N_3585,N_3495,N_3447);
or U3586 (N_3586,N_3479,N_3376);
xor U3587 (N_3587,N_3473,N_3472);
or U3588 (N_3588,N_3446,N_3416);
or U3589 (N_3589,N_3390,N_3440);
xnor U3590 (N_3590,N_3388,N_3481);
nor U3591 (N_3591,N_3458,N_3465);
and U3592 (N_3592,N_3459,N_3401);
nor U3593 (N_3593,N_3436,N_3457);
or U3594 (N_3594,N_3375,N_3443);
or U3595 (N_3595,N_3494,N_3442);
nand U3596 (N_3596,N_3425,N_3428);
xor U3597 (N_3597,N_3458,N_3494);
and U3598 (N_3598,N_3462,N_3489);
xor U3599 (N_3599,N_3406,N_3414);
and U3600 (N_3600,N_3387,N_3420);
and U3601 (N_3601,N_3398,N_3473);
nand U3602 (N_3602,N_3497,N_3462);
and U3603 (N_3603,N_3411,N_3416);
or U3604 (N_3604,N_3416,N_3439);
nor U3605 (N_3605,N_3460,N_3401);
nor U3606 (N_3606,N_3415,N_3413);
nor U3607 (N_3607,N_3375,N_3437);
and U3608 (N_3608,N_3395,N_3393);
or U3609 (N_3609,N_3461,N_3481);
xor U3610 (N_3610,N_3388,N_3450);
nor U3611 (N_3611,N_3475,N_3406);
xor U3612 (N_3612,N_3475,N_3409);
nand U3613 (N_3613,N_3430,N_3437);
nor U3614 (N_3614,N_3433,N_3443);
or U3615 (N_3615,N_3456,N_3439);
xnor U3616 (N_3616,N_3437,N_3472);
or U3617 (N_3617,N_3375,N_3410);
nor U3618 (N_3618,N_3461,N_3400);
nand U3619 (N_3619,N_3453,N_3467);
nor U3620 (N_3620,N_3398,N_3456);
nor U3621 (N_3621,N_3488,N_3406);
xnor U3622 (N_3622,N_3385,N_3417);
xor U3623 (N_3623,N_3381,N_3425);
nor U3624 (N_3624,N_3429,N_3439);
nand U3625 (N_3625,N_3622,N_3568);
xor U3626 (N_3626,N_3573,N_3606);
and U3627 (N_3627,N_3538,N_3555);
xnor U3628 (N_3628,N_3514,N_3536);
nand U3629 (N_3629,N_3578,N_3554);
or U3630 (N_3630,N_3520,N_3613);
nand U3631 (N_3631,N_3602,N_3582);
nor U3632 (N_3632,N_3614,N_3569);
nand U3633 (N_3633,N_3560,N_3524);
or U3634 (N_3634,N_3526,N_3551);
and U3635 (N_3635,N_3503,N_3597);
nand U3636 (N_3636,N_3604,N_3600);
nor U3637 (N_3637,N_3550,N_3599);
nor U3638 (N_3638,N_3505,N_3501);
or U3639 (N_3639,N_3615,N_3611);
nor U3640 (N_3640,N_3577,N_3541);
or U3641 (N_3641,N_3504,N_3570);
and U3642 (N_3642,N_3532,N_3587);
and U3643 (N_3643,N_3521,N_3556);
xor U3644 (N_3644,N_3512,N_3529);
nand U3645 (N_3645,N_3603,N_3547);
or U3646 (N_3646,N_3583,N_3588);
nor U3647 (N_3647,N_3579,N_3619);
nand U3648 (N_3648,N_3605,N_3539);
or U3649 (N_3649,N_3574,N_3517);
or U3650 (N_3650,N_3598,N_3562);
nor U3651 (N_3651,N_3516,N_3585);
xnor U3652 (N_3652,N_3540,N_3552);
xor U3653 (N_3653,N_3595,N_3527);
or U3654 (N_3654,N_3528,N_3565);
nand U3655 (N_3655,N_3559,N_3621);
xor U3656 (N_3656,N_3601,N_3572);
and U3657 (N_3657,N_3544,N_3612);
and U3658 (N_3658,N_3590,N_3563);
nor U3659 (N_3659,N_3542,N_3557);
nor U3660 (N_3660,N_3511,N_3518);
nand U3661 (N_3661,N_3593,N_3620);
nand U3662 (N_3662,N_3580,N_3519);
or U3663 (N_3663,N_3589,N_3531);
and U3664 (N_3664,N_3575,N_3533);
nor U3665 (N_3665,N_3607,N_3618);
and U3666 (N_3666,N_3510,N_3522);
nor U3667 (N_3667,N_3591,N_3515);
nand U3668 (N_3668,N_3525,N_3624);
or U3669 (N_3669,N_3610,N_3543);
xor U3670 (N_3670,N_3530,N_3500);
or U3671 (N_3671,N_3546,N_3608);
and U3672 (N_3672,N_3584,N_3509);
xnor U3673 (N_3673,N_3548,N_3596);
xnor U3674 (N_3674,N_3609,N_3507);
and U3675 (N_3675,N_3535,N_3564);
nand U3676 (N_3676,N_3586,N_3623);
and U3677 (N_3677,N_3616,N_3553);
or U3678 (N_3678,N_3571,N_3617);
or U3679 (N_3679,N_3534,N_3506);
nand U3680 (N_3680,N_3581,N_3537);
nand U3681 (N_3681,N_3561,N_3549);
and U3682 (N_3682,N_3558,N_3576);
nand U3683 (N_3683,N_3523,N_3592);
and U3684 (N_3684,N_3594,N_3502);
and U3685 (N_3685,N_3545,N_3513);
or U3686 (N_3686,N_3566,N_3508);
nor U3687 (N_3687,N_3567,N_3558);
and U3688 (N_3688,N_3551,N_3558);
and U3689 (N_3689,N_3501,N_3539);
and U3690 (N_3690,N_3607,N_3603);
xor U3691 (N_3691,N_3609,N_3514);
and U3692 (N_3692,N_3610,N_3595);
or U3693 (N_3693,N_3520,N_3531);
or U3694 (N_3694,N_3579,N_3597);
or U3695 (N_3695,N_3567,N_3603);
or U3696 (N_3696,N_3603,N_3503);
xor U3697 (N_3697,N_3595,N_3620);
or U3698 (N_3698,N_3617,N_3509);
nor U3699 (N_3699,N_3558,N_3543);
xnor U3700 (N_3700,N_3559,N_3509);
nand U3701 (N_3701,N_3612,N_3591);
and U3702 (N_3702,N_3566,N_3517);
nand U3703 (N_3703,N_3587,N_3547);
or U3704 (N_3704,N_3517,N_3593);
and U3705 (N_3705,N_3584,N_3603);
xnor U3706 (N_3706,N_3558,N_3532);
nand U3707 (N_3707,N_3610,N_3591);
xnor U3708 (N_3708,N_3603,N_3536);
nor U3709 (N_3709,N_3564,N_3552);
or U3710 (N_3710,N_3624,N_3622);
nor U3711 (N_3711,N_3585,N_3523);
nand U3712 (N_3712,N_3619,N_3507);
nand U3713 (N_3713,N_3534,N_3500);
nor U3714 (N_3714,N_3565,N_3577);
and U3715 (N_3715,N_3500,N_3552);
and U3716 (N_3716,N_3619,N_3610);
xnor U3717 (N_3717,N_3534,N_3624);
nor U3718 (N_3718,N_3505,N_3571);
nand U3719 (N_3719,N_3619,N_3542);
and U3720 (N_3720,N_3563,N_3534);
or U3721 (N_3721,N_3578,N_3551);
and U3722 (N_3722,N_3561,N_3579);
nand U3723 (N_3723,N_3508,N_3535);
or U3724 (N_3724,N_3603,N_3502);
nor U3725 (N_3725,N_3541,N_3550);
and U3726 (N_3726,N_3506,N_3596);
xor U3727 (N_3727,N_3612,N_3542);
nor U3728 (N_3728,N_3516,N_3598);
nand U3729 (N_3729,N_3569,N_3618);
nor U3730 (N_3730,N_3517,N_3538);
xor U3731 (N_3731,N_3544,N_3533);
xor U3732 (N_3732,N_3588,N_3549);
xnor U3733 (N_3733,N_3507,N_3584);
xnor U3734 (N_3734,N_3603,N_3509);
nor U3735 (N_3735,N_3567,N_3560);
and U3736 (N_3736,N_3584,N_3599);
or U3737 (N_3737,N_3508,N_3528);
nor U3738 (N_3738,N_3604,N_3622);
xnor U3739 (N_3739,N_3516,N_3569);
xor U3740 (N_3740,N_3507,N_3589);
nand U3741 (N_3741,N_3603,N_3554);
and U3742 (N_3742,N_3542,N_3525);
or U3743 (N_3743,N_3512,N_3623);
or U3744 (N_3744,N_3537,N_3542);
and U3745 (N_3745,N_3572,N_3557);
and U3746 (N_3746,N_3559,N_3615);
nor U3747 (N_3747,N_3520,N_3615);
or U3748 (N_3748,N_3509,N_3613);
and U3749 (N_3749,N_3623,N_3528);
xnor U3750 (N_3750,N_3691,N_3648);
or U3751 (N_3751,N_3702,N_3744);
xor U3752 (N_3752,N_3718,N_3717);
and U3753 (N_3753,N_3671,N_3683);
xor U3754 (N_3754,N_3741,N_3703);
nor U3755 (N_3755,N_3685,N_3738);
nor U3756 (N_3756,N_3666,N_3719);
nor U3757 (N_3757,N_3704,N_3707);
and U3758 (N_3758,N_3633,N_3734);
xnor U3759 (N_3759,N_3645,N_3700);
and U3760 (N_3760,N_3670,N_3661);
and U3761 (N_3761,N_3727,N_3667);
xor U3762 (N_3762,N_3743,N_3636);
and U3763 (N_3763,N_3684,N_3663);
or U3764 (N_3764,N_3669,N_3720);
nand U3765 (N_3765,N_3641,N_3640);
or U3766 (N_3766,N_3737,N_3639);
and U3767 (N_3767,N_3736,N_3735);
and U3768 (N_3768,N_3710,N_3635);
nand U3769 (N_3769,N_3730,N_3642);
nor U3770 (N_3770,N_3660,N_3726);
and U3771 (N_3771,N_3647,N_3729);
xnor U3772 (N_3772,N_3631,N_3644);
nand U3773 (N_3773,N_3628,N_3716);
or U3774 (N_3774,N_3712,N_3654);
and U3775 (N_3775,N_3652,N_3678);
nor U3776 (N_3776,N_3664,N_3698);
or U3777 (N_3777,N_3749,N_3714);
nand U3778 (N_3778,N_3655,N_3651);
nor U3779 (N_3779,N_3746,N_3689);
nor U3780 (N_3780,N_3662,N_3657);
nand U3781 (N_3781,N_3687,N_3626);
xnor U3782 (N_3782,N_3659,N_3688);
or U3783 (N_3783,N_3711,N_3679);
nor U3784 (N_3784,N_3747,N_3630);
xor U3785 (N_3785,N_3653,N_3637);
xnor U3786 (N_3786,N_3715,N_3681);
xor U3787 (N_3787,N_3680,N_3646);
nand U3788 (N_3788,N_3674,N_3643);
and U3789 (N_3789,N_3706,N_3625);
nand U3790 (N_3790,N_3733,N_3692);
nor U3791 (N_3791,N_3723,N_3725);
nand U3792 (N_3792,N_3696,N_3632);
and U3793 (N_3793,N_3629,N_3672);
nand U3794 (N_3794,N_3728,N_3699);
xnor U3795 (N_3795,N_3713,N_3722);
or U3796 (N_3796,N_3745,N_3690);
xnor U3797 (N_3797,N_3701,N_3656);
and U3798 (N_3798,N_3665,N_3650);
and U3799 (N_3799,N_3638,N_3705);
xor U3800 (N_3800,N_3739,N_3708);
nand U3801 (N_3801,N_3695,N_3709);
or U3802 (N_3802,N_3658,N_3721);
nor U3803 (N_3803,N_3682,N_3649);
nor U3804 (N_3804,N_3748,N_3668);
and U3805 (N_3805,N_3732,N_3724);
nand U3806 (N_3806,N_3673,N_3742);
nor U3807 (N_3807,N_3693,N_3694);
and U3808 (N_3808,N_3697,N_3686);
xor U3809 (N_3809,N_3627,N_3676);
xnor U3810 (N_3810,N_3675,N_3740);
nor U3811 (N_3811,N_3677,N_3731);
xnor U3812 (N_3812,N_3634,N_3638);
or U3813 (N_3813,N_3727,N_3644);
nand U3814 (N_3814,N_3704,N_3625);
or U3815 (N_3815,N_3692,N_3672);
xor U3816 (N_3816,N_3663,N_3708);
nor U3817 (N_3817,N_3721,N_3648);
or U3818 (N_3818,N_3699,N_3700);
or U3819 (N_3819,N_3646,N_3696);
xnor U3820 (N_3820,N_3745,N_3685);
or U3821 (N_3821,N_3678,N_3666);
nor U3822 (N_3822,N_3703,N_3638);
and U3823 (N_3823,N_3709,N_3705);
and U3824 (N_3824,N_3682,N_3745);
nand U3825 (N_3825,N_3631,N_3719);
nor U3826 (N_3826,N_3729,N_3741);
xnor U3827 (N_3827,N_3677,N_3745);
nand U3828 (N_3828,N_3675,N_3749);
or U3829 (N_3829,N_3745,N_3720);
nor U3830 (N_3830,N_3730,N_3668);
or U3831 (N_3831,N_3708,N_3678);
or U3832 (N_3832,N_3629,N_3677);
nand U3833 (N_3833,N_3719,N_3670);
and U3834 (N_3834,N_3745,N_3722);
nor U3835 (N_3835,N_3663,N_3670);
and U3836 (N_3836,N_3675,N_3641);
and U3837 (N_3837,N_3701,N_3685);
nor U3838 (N_3838,N_3730,N_3684);
nor U3839 (N_3839,N_3654,N_3658);
or U3840 (N_3840,N_3731,N_3687);
nor U3841 (N_3841,N_3716,N_3742);
nor U3842 (N_3842,N_3688,N_3626);
and U3843 (N_3843,N_3718,N_3633);
nor U3844 (N_3844,N_3746,N_3655);
xor U3845 (N_3845,N_3672,N_3746);
xor U3846 (N_3846,N_3662,N_3691);
nor U3847 (N_3847,N_3673,N_3726);
nor U3848 (N_3848,N_3635,N_3683);
and U3849 (N_3849,N_3735,N_3679);
nand U3850 (N_3850,N_3648,N_3671);
and U3851 (N_3851,N_3656,N_3715);
xnor U3852 (N_3852,N_3715,N_3682);
nand U3853 (N_3853,N_3637,N_3706);
or U3854 (N_3854,N_3707,N_3628);
xnor U3855 (N_3855,N_3660,N_3661);
nor U3856 (N_3856,N_3668,N_3646);
and U3857 (N_3857,N_3745,N_3633);
nor U3858 (N_3858,N_3728,N_3705);
nor U3859 (N_3859,N_3660,N_3717);
nand U3860 (N_3860,N_3652,N_3647);
nor U3861 (N_3861,N_3646,N_3721);
xnor U3862 (N_3862,N_3633,N_3686);
xor U3863 (N_3863,N_3730,N_3704);
nor U3864 (N_3864,N_3646,N_3636);
nor U3865 (N_3865,N_3634,N_3734);
xor U3866 (N_3866,N_3678,N_3644);
nand U3867 (N_3867,N_3719,N_3740);
or U3868 (N_3868,N_3639,N_3714);
nand U3869 (N_3869,N_3708,N_3649);
nor U3870 (N_3870,N_3641,N_3672);
and U3871 (N_3871,N_3680,N_3685);
nor U3872 (N_3872,N_3700,N_3709);
nor U3873 (N_3873,N_3702,N_3647);
or U3874 (N_3874,N_3639,N_3630);
or U3875 (N_3875,N_3803,N_3858);
nor U3876 (N_3876,N_3773,N_3855);
or U3877 (N_3877,N_3798,N_3809);
xnor U3878 (N_3878,N_3859,N_3864);
nor U3879 (N_3879,N_3761,N_3767);
nor U3880 (N_3880,N_3756,N_3825);
and U3881 (N_3881,N_3805,N_3837);
and U3882 (N_3882,N_3799,N_3784);
and U3883 (N_3883,N_3827,N_3786);
and U3884 (N_3884,N_3765,N_3819);
or U3885 (N_3885,N_3848,N_3793);
xor U3886 (N_3886,N_3755,N_3865);
xnor U3887 (N_3887,N_3833,N_3790);
nand U3888 (N_3888,N_3812,N_3842);
or U3889 (N_3889,N_3787,N_3838);
nand U3890 (N_3890,N_3792,N_3808);
and U3891 (N_3891,N_3832,N_3866);
or U3892 (N_3892,N_3785,N_3804);
nand U3893 (N_3893,N_3847,N_3759);
xnor U3894 (N_3894,N_3802,N_3769);
nand U3895 (N_3895,N_3826,N_3823);
nor U3896 (N_3896,N_3760,N_3778);
xnor U3897 (N_3897,N_3811,N_3852);
nand U3898 (N_3898,N_3830,N_3782);
and U3899 (N_3899,N_3816,N_3857);
nand U3900 (N_3900,N_3860,N_3750);
or U3901 (N_3901,N_3814,N_3783);
nand U3902 (N_3902,N_3817,N_3766);
nand U3903 (N_3903,N_3751,N_3774);
nand U3904 (N_3904,N_3763,N_3835);
and U3905 (N_3905,N_3821,N_3839);
and U3906 (N_3906,N_3795,N_3813);
nand U3907 (N_3907,N_3818,N_3849);
nor U3908 (N_3908,N_3781,N_3831);
and U3909 (N_3909,N_3753,N_3851);
nor U3910 (N_3910,N_3770,N_3867);
or U3911 (N_3911,N_3828,N_3868);
xnor U3912 (N_3912,N_3789,N_3788);
or U3913 (N_3913,N_3841,N_3872);
and U3914 (N_3914,N_3796,N_3764);
and U3915 (N_3915,N_3776,N_3807);
and U3916 (N_3916,N_3806,N_3797);
and U3917 (N_3917,N_3794,N_3752);
nor U3918 (N_3918,N_3854,N_3824);
and U3919 (N_3919,N_3810,N_3772);
or U3920 (N_3920,N_3844,N_3800);
or U3921 (N_3921,N_3873,N_3762);
xnor U3922 (N_3922,N_3815,N_3850);
nor U3923 (N_3923,N_3757,N_3829);
and U3924 (N_3924,N_3820,N_3862);
nor U3925 (N_3925,N_3840,N_3861);
nor U3926 (N_3926,N_3853,N_3822);
xor U3927 (N_3927,N_3869,N_3843);
nand U3928 (N_3928,N_3768,N_3754);
nand U3929 (N_3929,N_3777,N_3874);
and U3930 (N_3930,N_3846,N_3834);
or U3931 (N_3931,N_3791,N_3856);
or U3932 (N_3932,N_3779,N_3780);
xor U3933 (N_3933,N_3845,N_3836);
nand U3934 (N_3934,N_3870,N_3771);
or U3935 (N_3935,N_3801,N_3863);
xor U3936 (N_3936,N_3871,N_3758);
or U3937 (N_3937,N_3775,N_3859);
xor U3938 (N_3938,N_3819,N_3818);
or U3939 (N_3939,N_3832,N_3786);
nor U3940 (N_3940,N_3817,N_3764);
nand U3941 (N_3941,N_3803,N_3873);
and U3942 (N_3942,N_3769,N_3771);
or U3943 (N_3943,N_3781,N_3851);
and U3944 (N_3944,N_3841,N_3786);
nor U3945 (N_3945,N_3785,N_3796);
and U3946 (N_3946,N_3809,N_3806);
and U3947 (N_3947,N_3775,N_3810);
and U3948 (N_3948,N_3778,N_3805);
xor U3949 (N_3949,N_3833,N_3818);
xor U3950 (N_3950,N_3782,N_3802);
nand U3951 (N_3951,N_3791,N_3850);
or U3952 (N_3952,N_3775,N_3852);
nor U3953 (N_3953,N_3861,N_3841);
nor U3954 (N_3954,N_3769,N_3843);
or U3955 (N_3955,N_3801,N_3775);
nand U3956 (N_3956,N_3841,N_3858);
and U3957 (N_3957,N_3764,N_3871);
and U3958 (N_3958,N_3827,N_3781);
or U3959 (N_3959,N_3854,N_3860);
xor U3960 (N_3960,N_3844,N_3860);
nand U3961 (N_3961,N_3758,N_3843);
or U3962 (N_3962,N_3800,N_3798);
or U3963 (N_3963,N_3781,N_3812);
and U3964 (N_3964,N_3807,N_3866);
nand U3965 (N_3965,N_3827,N_3788);
xnor U3966 (N_3966,N_3846,N_3753);
and U3967 (N_3967,N_3763,N_3798);
nand U3968 (N_3968,N_3778,N_3848);
nand U3969 (N_3969,N_3784,N_3786);
xor U3970 (N_3970,N_3836,N_3804);
nand U3971 (N_3971,N_3808,N_3780);
xnor U3972 (N_3972,N_3848,N_3851);
nor U3973 (N_3973,N_3792,N_3800);
or U3974 (N_3974,N_3845,N_3806);
xnor U3975 (N_3975,N_3865,N_3799);
nor U3976 (N_3976,N_3784,N_3853);
and U3977 (N_3977,N_3775,N_3760);
nand U3978 (N_3978,N_3853,N_3790);
nand U3979 (N_3979,N_3803,N_3852);
xor U3980 (N_3980,N_3765,N_3766);
nand U3981 (N_3981,N_3784,N_3873);
or U3982 (N_3982,N_3818,N_3863);
or U3983 (N_3983,N_3835,N_3841);
or U3984 (N_3984,N_3781,N_3770);
nand U3985 (N_3985,N_3760,N_3762);
nand U3986 (N_3986,N_3776,N_3799);
nor U3987 (N_3987,N_3772,N_3847);
nand U3988 (N_3988,N_3797,N_3794);
nor U3989 (N_3989,N_3840,N_3868);
and U3990 (N_3990,N_3868,N_3869);
nor U3991 (N_3991,N_3793,N_3867);
nand U3992 (N_3992,N_3847,N_3827);
nand U3993 (N_3993,N_3791,N_3765);
and U3994 (N_3994,N_3766,N_3808);
and U3995 (N_3995,N_3785,N_3860);
xor U3996 (N_3996,N_3788,N_3856);
or U3997 (N_3997,N_3781,N_3778);
nand U3998 (N_3998,N_3767,N_3807);
nor U3999 (N_3999,N_3750,N_3855);
nor U4000 (N_4000,N_3948,N_3887);
nand U4001 (N_4001,N_3978,N_3935);
and U4002 (N_4002,N_3898,N_3920);
nor U4003 (N_4003,N_3928,N_3925);
nand U4004 (N_4004,N_3999,N_3956);
nor U4005 (N_4005,N_3955,N_3906);
xnor U4006 (N_4006,N_3913,N_3875);
xor U4007 (N_4007,N_3989,N_3900);
or U4008 (N_4008,N_3943,N_3903);
nor U4009 (N_4009,N_3924,N_3915);
nand U4010 (N_4010,N_3939,N_3946);
nand U4011 (N_4011,N_3967,N_3944);
and U4012 (N_4012,N_3910,N_3963);
and U4013 (N_4013,N_3973,N_3895);
or U4014 (N_4014,N_3986,N_3897);
or U4015 (N_4015,N_3996,N_3994);
xor U4016 (N_4016,N_3883,N_3917);
nor U4017 (N_4017,N_3893,N_3938);
or U4018 (N_4018,N_3899,N_3908);
xor U4019 (N_4019,N_3894,N_3905);
and U4020 (N_4020,N_3936,N_3968);
xor U4021 (N_4021,N_3988,N_3902);
nand U4022 (N_4022,N_3942,N_3987);
and U4023 (N_4023,N_3964,N_3975);
and U4024 (N_4024,N_3941,N_3927);
nor U4025 (N_4025,N_3951,N_3914);
or U4026 (N_4026,N_3977,N_3884);
xor U4027 (N_4027,N_3993,N_3947);
or U4028 (N_4028,N_3998,N_3958);
xnor U4029 (N_4029,N_3926,N_3892);
and U4030 (N_4030,N_3891,N_3981);
or U4031 (N_4031,N_3923,N_3904);
and U4032 (N_4032,N_3980,N_3990);
and U4033 (N_4033,N_3878,N_3952);
nand U4034 (N_4034,N_3881,N_3901);
nor U4035 (N_4035,N_3957,N_3916);
nor U4036 (N_4036,N_3896,N_3911);
nand U4037 (N_4037,N_3937,N_3921);
nor U4038 (N_4038,N_3953,N_3992);
nor U4039 (N_4039,N_3933,N_3888);
nand U4040 (N_4040,N_3960,N_3976);
nand U4041 (N_4041,N_3890,N_3991);
nor U4042 (N_4042,N_3995,N_3966);
xnor U4043 (N_4043,N_3962,N_3907);
nand U4044 (N_4044,N_3997,N_3961);
and U4045 (N_4045,N_3886,N_3970);
xor U4046 (N_4046,N_3922,N_3876);
and U4047 (N_4047,N_3877,N_3934);
xnor U4048 (N_4048,N_3950,N_3880);
nand U4049 (N_4049,N_3929,N_3945);
nand U4050 (N_4050,N_3965,N_3879);
or U4051 (N_4051,N_3889,N_3885);
xor U4052 (N_4052,N_3969,N_3954);
xnor U4053 (N_4053,N_3983,N_3882);
nor U4054 (N_4054,N_3930,N_3932);
xnor U4055 (N_4055,N_3909,N_3959);
or U4056 (N_4056,N_3931,N_3918);
and U4057 (N_4057,N_3949,N_3974);
nor U4058 (N_4058,N_3972,N_3985);
nand U4059 (N_4059,N_3971,N_3940);
nor U4060 (N_4060,N_3984,N_3982);
or U4061 (N_4061,N_3919,N_3979);
or U4062 (N_4062,N_3912,N_3952);
or U4063 (N_4063,N_3946,N_3881);
nor U4064 (N_4064,N_3899,N_3924);
or U4065 (N_4065,N_3976,N_3876);
and U4066 (N_4066,N_3910,N_3989);
nor U4067 (N_4067,N_3977,N_3912);
nor U4068 (N_4068,N_3949,N_3885);
or U4069 (N_4069,N_3937,N_3957);
xnor U4070 (N_4070,N_3952,N_3893);
xor U4071 (N_4071,N_3954,N_3881);
or U4072 (N_4072,N_3921,N_3965);
nor U4073 (N_4073,N_3960,N_3898);
or U4074 (N_4074,N_3993,N_3923);
xor U4075 (N_4075,N_3925,N_3927);
and U4076 (N_4076,N_3944,N_3905);
nand U4077 (N_4077,N_3984,N_3962);
nor U4078 (N_4078,N_3944,N_3896);
or U4079 (N_4079,N_3906,N_3933);
nor U4080 (N_4080,N_3942,N_3981);
nand U4081 (N_4081,N_3968,N_3965);
and U4082 (N_4082,N_3957,N_3983);
xor U4083 (N_4083,N_3978,N_3971);
and U4084 (N_4084,N_3883,N_3896);
and U4085 (N_4085,N_3885,N_3910);
xor U4086 (N_4086,N_3922,N_3878);
nand U4087 (N_4087,N_3921,N_3876);
nor U4088 (N_4088,N_3922,N_3976);
or U4089 (N_4089,N_3909,N_3877);
nor U4090 (N_4090,N_3945,N_3875);
xnor U4091 (N_4091,N_3909,N_3990);
nand U4092 (N_4092,N_3895,N_3933);
nand U4093 (N_4093,N_3916,N_3882);
xor U4094 (N_4094,N_3928,N_3901);
nand U4095 (N_4095,N_3897,N_3903);
and U4096 (N_4096,N_3985,N_3945);
xnor U4097 (N_4097,N_3961,N_3924);
nor U4098 (N_4098,N_3988,N_3931);
nor U4099 (N_4099,N_3991,N_3911);
xor U4100 (N_4100,N_3984,N_3880);
nand U4101 (N_4101,N_3897,N_3892);
or U4102 (N_4102,N_3959,N_3974);
or U4103 (N_4103,N_3945,N_3893);
nand U4104 (N_4104,N_3970,N_3903);
or U4105 (N_4105,N_3876,N_3878);
and U4106 (N_4106,N_3939,N_3998);
and U4107 (N_4107,N_3995,N_3932);
xor U4108 (N_4108,N_3911,N_3877);
nand U4109 (N_4109,N_3933,N_3964);
or U4110 (N_4110,N_3996,N_3923);
xnor U4111 (N_4111,N_3899,N_3925);
nand U4112 (N_4112,N_3875,N_3932);
nand U4113 (N_4113,N_3994,N_3897);
or U4114 (N_4114,N_3989,N_3967);
or U4115 (N_4115,N_3959,N_3991);
nor U4116 (N_4116,N_3959,N_3898);
or U4117 (N_4117,N_3954,N_3908);
or U4118 (N_4118,N_3968,N_3964);
and U4119 (N_4119,N_3969,N_3941);
xor U4120 (N_4120,N_3954,N_3984);
nand U4121 (N_4121,N_3999,N_3922);
nand U4122 (N_4122,N_3883,N_3984);
nand U4123 (N_4123,N_3901,N_3953);
nor U4124 (N_4124,N_3941,N_3934);
and U4125 (N_4125,N_4117,N_4084);
xnor U4126 (N_4126,N_4035,N_4068);
nand U4127 (N_4127,N_4115,N_4110);
nand U4128 (N_4128,N_4097,N_4099);
nor U4129 (N_4129,N_4015,N_4094);
nor U4130 (N_4130,N_4118,N_4091);
nor U4131 (N_4131,N_4029,N_4012);
or U4132 (N_4132,N_4053,N_4036);
and U4133 (N_4133,N_4000,N_4079);
nor U4134 (N_4134,N_4089,N_4070);
and U4135 (N_4135,N_4047,N_4098);
nand U4136 (N_4136,N_4083,N_4078);
xor U4137 (N_4137,N_4034,N_4121);
xor U4138 (N_4138,N_4027,N_4033);
nand U4139 (N_4139,N_4050,N_4093);
or U4140 (N_4140,N_4032,N_4011);
and U4141 (N_4141,N_4046,N_4082);
xnor U4142 (N_4142,N_4080,N_4122);
and U4143 (N_4143,N_4030,N_4076);
or U4144 (N_4144,N_4109,N_4003);
xnor U4145 (N_4145,N_4088,N_4111);
or U4146 (N_4146,N_4075,N_4096);
xor U4147 (N_4147,N_4037,N_4045);
nor U4148 (N_4148,N_4028,N_4042);
nor U4149 (N_4149,N_4025,N_4104);
nor U4150 (N_4150,N_4038,N_4064);
xnor U4151 (N_4151,N_4002,N_4018);
or U4152 (N_4152,N_4081,N_4017);
nand U4153 (N_4153,N_4040,N_4086);
and U4154 (N_4154,N_4065,N_4105);
nand U4155 (N_4155,N_4026,N_4061);
nor U4156 (N_4156,N_4077,N_4113);
xor U4157 (N_4157,N_4116,N_4072);
nand U4158 (N_4158,N_4013,N_4052);
and U4159 (N_4159,N_4023,N_4063);
nor U4160 (N_4160,N_4090,N_4020);
xnor U4161 (N_4161,N_4074,N_4006);
nand U4162 (N_4162,N_4041,N_4067);
and U4163 (N_4163,N_4048,N_4044);
and U4164 (N_4164,N_4057,N_4112);
xor U4165 (N_4165,N_4119,N_4107);
xor U4166 (N_4166,N_4106,N_4087);
nor U4167 (N_4167,N_4120,N_4014);
or U4168 (N_4168,N_4039,N_4066);
nand U4169 (N_4169,N_4021,N_4103);
and U4170 (N_4170,N_4059,N_4102);
nand U4171 (N_4171,N_4054,N_4124);
nand U4172 (N_4172,N_4043,N_4100);
nand U4173 (N_4173,N_4004,N_4049);
or U4174 (N_4174,N_4071,N_4008);
and U4175 (N_4175,N_4092,N_4062);
xnor U4176 (N_4176,N_4055,N_4085);
nand U4177 (N_4177,N_4009,N_4114);
nand U4178 (N_4178,N_4069,N_4095);
xnor U4179 (N_4179,N_4123,N_4051);
nand U4180 (N_4180,N_4101,N_4060);
and U4181 (N_4181,N_4005,N_4056);
xor U4182 (N_4182,N_4019,N_4073);
nor U4183 (N_4183,N_4058,N_4022);
or U4184 (N_4184,N_4010,N_4016);
and U4185 (N_4185,N_4007,N_4108);
nor U4186 (N_4186,N_4024,N_4031);
xor U4187 (N_4187,N_4001,N_4060);
nand U4188 (N_4188,N_4112,N_4011);
nor U4189 (N_4189,N_4017,N_4075);
and U4190 (N_4190,N_4054,N_4093);
or U4191 (N_4191,N_4122,N_4077);
nand U4192 (N_4192,N_4002,N_4086);
xnor U4193 (N_4193,N_4018,N_4098);
nor U4194 (N_4194,N_4036,N_4012);
nor U4195 (N_4195,N_4043,N_4044);
or U4196 (N_4196,N_4005,N_4042);
or U4197 (N_4197,N_4082,N_4121);
and U4198 (N_4198,N_4001,N_4053);
and U4199 (N_4199,N_4026,N_4086);
or U4200 (N_4200,N_4000,N_4071);
and U4201 (N_4201,N_4026,N_4029);
or U4202 (N_4202,N_4041,N_4116);
or U4203 (N_4203,N_4098,N_4067);
xor U4204 (N_4204,N_4003,N_4049);
xor U4205 (N_4205,N_4030,N_4018);
nor U4206 (N_4206,N_4007,N_4084);
and U4207 (N_4207,N_4075,N_4000);
or U4208 (N_4208,N_4026,N_4073);
or U4209 (N_4209,N_4083,N_4070);
nor U4210 (N_4210,N_4076,N_4015);
and U4211 (N_4211,N_4001,N_4111);
xnor U4212 (N_4212,N_4107,N_4053);
xnor U4213 (N_4213,N_4005,N_4055);
nand U4214 (N_4214,N_4124,N_4062);
nand U4215 (N_4215,N_4003,N_4020);
nand U4216 (N_4216,N_4066,N_4070);
xnor U4217 (N_4217,N_4110,N_4028);
or U4218 (N_4218,N_4087,N_4089);
nand U4219 (N_4219,N_4050,N_4077);
or U4220 (N_4220,N_4029,N_4015);
or U4221 (N_4221,N_4076,N_4001);
nand U4222 (N_4222,N_4001,N_4082);
nand U4223 (N_4223,N_4101,N_4109);
nor U4224 (N_4224,N_4001,N_4114);
or U4225 (N_4225,N_4086,N_4113);
nor U4226 (N_4226,N_4076,N_4093);
and U4227 (N_4227,N_4019,N_4091);
or U4228 (N_4228,N_4116,N_4115);
or U4229 (N_4229,N_4070,N_4028);
nand U4230 (N_4230,N_4075,N_4089);
nand U4231 (N_4231,N_4039,N_4105);
nand U4232 (N_4232,N_4102,N_4022);
nand U4233 (N_4233,N_4096,N_4060);
nor U4234 (N_4234,N_4036,N_4064);
nand U4235 (N_4235,N_4058,N_4078);
nor U4236 (N_4236,N_4095,N_4024);
nand U4237 (N_4237,N_4112,N_4107);
nand U4238 (N_4238,N_4074,N_4030);
nand U4239 (N_4239,N_4005,N_4085);
and U4240 (N_4240,N_4025,N_4067);
nand U4241 (N_4241,N_4009,N_4001);
or U4242 (N_4242,N_4040,N_4044);
xnor U4243 (N_4243,N_4065,N_4032);
nand U4244 (N_4244,N_4028,N_4044);
and U4245 (N_4245,N_4121,N_4070);
and U4246 (N_4246,N_4112,N_4048);
nand U4247 (N_4247,N_4061,N_4070);
nor U4248 (N_4248,N_4115,N_4088);
or U4249 (N_4249,N_4036,N_4080);
xnor U4250 (N_4250,N_4173,N_4162);
xnor U4251 (N_4251,N_4138,N_4210);
nor U4252 (N_4252,N_4144,N_4176);
or U4253 (N_4253,N_4148,N_4212);
xor U4254 (N_4254,N_4145,N_4228);
and U4255 (N_4255,N_4195,N_4218);
nand U4256 (N_4256,N_4225,N_4182);
nor U4257 (N_4257,N_4203,N_4244);
or U4258 (N_4258,N_4245,N_4169);
or U4259 (N_4259,N_4198,N_4231);
nand U4260 (N_4260,N_4134,N_4174);
nand U4261 (N_4261,N_4136,N_4154);
or U4262 (N_4262,N_4213,N_4215);
nor U4263 (N_4263,N_4164,N_4149);
nor U4264 (N_4264,N_4177,N_4196);
or U4265 (N_4265,N_4188,N_4223);
or U4266 (N_4266,N_4159,N_4157);
nand U4267 (N_4267,N_4161,N_4240);
or U4268 (N_4268,N_4192,N_4128);
nor U4269 (N_4269,N_4220,N_4202);
nand U4270 (N_4270,N_4249,N_4178);
nand U4271 (N_4271,N_4156,N_4126);
nor U4272 (N_4272,N_4175,N_4221);
xnor U4273 (N_4273,N_4242,N_4230);
or U4274 (N_4274,N_4236,N_4191);
nor U4275 (N_4275,N_4224,N_4247);
xor U4276 (N_4276,N_4235,N_4181);
xnor U4277 (N_4277,N_4189,N_4205);
xor U4278 (N_4278,N_4137,N_4170);
xor U4279 (N_4279,N_4211,N_4186);
or U4280 (N_4280,N_4172,N_4127);
nor U4281 (N_4281,N_4227,N_4153);
nor U4282 (N_4282,N_4216,N_4197);
nor U4283 (N_4283,N_4226,N_4229);
or U4284 (N_4284,N_4150,N_4139);
and U4285 (N_4285,N_4163,N_4142);
nand U4286 (N_4286,N_4160,N_4246);
and U4287 (N_4287,N_4135,N_4180);
xnor U4288 (N_4288,N_4155,N_4241);
or U4289 (N_4289,N_4201,N_4130);
nand U4290 (N_4290,N_4243,N_4183);
or U4291 (N_4291,N_4167,N_4187);
nor U4292 (N_4292,N_4143,N_4168);
nand U4293 (N_4293,N_4141,N_4129);
or U4294 (N_4294,N_4204,N_4179);
nor U4295 (N_4295,N_4184,N_4125);
nand U4296 (N_4296,N_4237,N_4209);
xnor U4297 (N_4297,N_4199,N_4152);
xor U4298 (N_4298,N_4217,N_4200);
and U4299 (N_4299,N_4248,N_4190);
xnor U4300 (N_4300,N_4214,N_4171);
nand U4301 (N_4301,N_4158,N_4146);
or U4302 (N_4302,N_4166,N_4239);
and U4303 (N_4303,N_4133,N_4132);
nand U4304 (N_4304,N_4219,N_4222);
nand U4305 (N_4305,N_4233,N_4208);
nor U4306 (N_4306,N_4165,N_4185);
xnor U4307 (N_4307,N_4206,N_4238);
nand U4308 (N_4308,N_4140,N_4234);
xor U4309 (N_4309,N_4193,N_4232);
nand U4310 (N_4310,N_4151,N_4207);
nand U4311 (N_4311,N_4131,N_4147);
nand U4312 (N_4312,N_4194,N_4207);
nand U4313 (N_4313,N_4242,N_4182);
xor U4314 (N_4314,N_4237,N_4207);
nand U4315 (N_4315,N_4209,N_4248);
and U4316 (N_4316,N_4177,N_4151);
or U4317 (N_4317,N_4234,N_4229);
nor U4318 (N_4318,N_4145,N_4237);
nor U4319 (N_4319,N_4128,N_4147);
or U4320 (N_4320,N_4178,N_4210);
and U4321 (N_4321,N_4210,N_4131);
xnor U4322 (N_4322,N_4142,N_4180);
nor U4323 (N_4323,N_4157,N_4205);
nand U4324 (N_4324,N_4137,N_4218);
xor U4325 (N_4325,N_4214,N_4193);
and U4326 (N_4326,N_4202,N_4216);
or U4327 (N_4327,N_4199,N_4145);
xor U4328 (N_4328,N_4189,N_4240);
nor U4329 (N_4329,N_4185,N_4172);
nor U4330 (N_4330,N_4151,N_4205);
xor U4331 (N_4331,N_4147,N_4144);
and U4332 (N_4332,N_4188,N_4213);
xor U4333 (N_4333,N_4189,N_4137);
nand U4334 (N_4334,N_4151,N_4139);
nor U4335 (N_4335,N_4236,N_4187);
nor U4336 (N_4336,N_4128,N_4143);
or U4337 (N_4337,N_4214,N_4169);
and U4338 (N_4338,N_4144,N_4244);
nand U4339 (N_4339,N_4196,N_4153);
nand U4340 (N_4340,N_4129,N_4155);
nand U4341 (N_4341,N_4151,N_4163);
and U4342 (N_4342,N_4139,N_4136);
nor U4343 (N_4343,N_4178,N_4189);
nor U4344 (N_4344,N_4213,N_4186);
nand U4345 (N_4345,N_4224,N_4155);
xor U4346 (N_4346,N_4132,N_4195);
nor U4347 (N_4347,N_4200,N_4138);
and U4348 (N_4348,N_4242,N_4151);
or U4349 (N_4349,N_4170,N_4164);
xnor U4350 (N_4350,N_4239,N_4204);
or U4351 (N_4351,N_4146,N_4173);
xor U4352 (N_4352,N_4192,N_4191);
or U4353 (N_4353,N_4232,N_4224);
nor U4354 (N_4354,N_4182,N_4240);
nand U4355 (N_4355,N_4215,N_4171);
or U4356 (N_4356,N_4198,N_4200);
or U4357 (N_4357,N_4131,N_4142);
nor U4358 (N_4358,N_4172,N_4244);
and U4359 (N_4359,N_4170,N_4195);
or U4360 (N_4360,N_4149,N_4144);
or U4361 (N_4361,N_4138,N_4157);
xnor U4362 (N_4362,N_4179,N_4185);
and U4363 (N_4363,N_4189,N_4138);
nand U4364 (N_4364,N_4198,N_4229);
or U4365 (N_4365,N_4138,N_4235);
nand U4366 (N_4366,N_4209,N_4132);
xnor U4367 (N_4367,N_4199,N_4231);
and U4368 (N_4368,N_4137,N_4151);
or U4369 (N_4369,N_4126,N_4151);
nand U4370 (N_4370,N_4145,N_4178);
and U4371 (N_4371,N_4133,N_4247);
nor U4372 (N_4372,N_4161,N_4191);
and U4373 (N_4373,N_4223,N_4246);
nand U4374 (N_4374,N_4204,N_4212);
xor U4375 (N_4375,N_4354,N_4338);
and U4376 (N_4376,N_4350,N_4341);
xor U4377 (N_4377,N_4331,N_4305);
or U4378 (N_4378,N_4348,N_4282);
xor U4379 (N_4379,N_4367,N_4294);
and U4380 (N_4380,N_4308,N_4273);
xor U4381 (N_4381,N_4276,N_4333);
nor U4382 (N_4382,N_4265,N_4297);
nor U4383 (N_4383,N_4323,N_4343);
nand U4384 (N_4384,N_4255,N_4256);
nor U4385 (N_4385,N_4303,N_4372);
nand U4386 (N_4386,N_4327,N_4285);
xor U4387 (N_4387,N_4309,N_4369);
and U4388 (N_4388,N_4317,N_4361);
nor U4389 (N_4389,N_4352,N_4342);
or U4390 (N_4390,N_4374,N_4292);
xnor U4391 (N_4391,N_4259,N_4290);
or U4392 (N_4392,N_4293,N_4275);
nand U4393 (N_4393,N_4349,N_4300);
nand U4394 (N_4394,N_4360,N_4268);
nor U4395 (N_4395,N_4298,N_4332);
xor U4396 (N_4396,N_4362,N_4336);
and U4397 (N_4397,N_4254,N_4281);
and U4398 (N_4398,N_4364,N_4301);
xnor U4399 (N_4399,N_4316,N_4264);
or U4400 (N_4400,N_4251,N_4344);
and U4401 (N_4401,N_4335,N_4337);
nor U4402 (N_4402,N_4289,N_4267);
nor U4403 (N_4403,N_4358,N_4258);
nand U4404 (N_4404,N_4257,N_4329);
nor U4405 (N_4405,N_4373,N_4271);
xor U4406 (N_4406,N_4287,N_4288);
nor U4407 (N_4407,N_4325,N_4299);
nand U4408 (N_4408,N_4311,N_4263);
nor U4409 (N_4409,N_4266,N_4353);
nand U4410 (N_4410,N_4359,N_4334);
or U4411 (N_4411,N_4260,N_4365);
xnor U4412 (N_4412,N_4357,N_4340);
nor U4413 (N_4413,N_4330,N_4370);
or U4414 (N_4414,N_4313,N_4253);
xor U4415 (N_4415,N_4278,N_4261);
nand U4416 (N_4416,N_4250,N_4328);
and U4417 (N_4417,N_4291,N_4269);
or U4418 (N_4418,N_4306,N_4347);
or U4419 (N_4419,N_4318,N_4363);
or U4420 (N_4420,N_4339,N_4326);
nand U4421 (N_4421,N_4296,N_4274);
xnor U4422 (N_4422,N_4280,N_4319);
nand U4423 (N_4423,N_4315,N_4286);
or U4424 (N_4424,N_4270,N_4356);
nand U4425 (N_4425,N_4371,N_4272);
nor U4426 (N_4426,N_4321,N_4279);
nor U4427 (N_4427,N_4277,N_4345);
xnor U4428 (N_4428,N_4346,N_4314);
xor U4429 (N_4429,N_4284,N_4355);
or U4430 (N_4430,N_4307,N_4322);
or U4431 (N_4431,N_4351,N_4368);
xor U4432 (N_4432,N_4366,N_4310);
nor U4433 (N_4433,N_4324,N_4283);
nor U4434 (N_4434,N_4295,N_4252);
nand U4435 (N_4435,N_4302,N_4262);
nand U4436 (N_4436,N_4304,N_4320);
nand U4437 (N_4437,N_4312,N_4284);
nor U4438 (N_4438,N_4260,N_4349);
and U4439 (N_4439,N_4318,N_4331);
and U4440 (N_4440,N_4321,N_4320);
nand U4441 (N_4441,N_4276,N_4341);
nor U4442 (N_4442,N_4261,N_4360);
nor U4443 (N_4443,N_4347,N_4338);
nand U4444 (N_4444,N_4324,N_4298);
nand U4445 (N_4445,N_4298,N_4368);
nand U4446 (N_4446,N_4316,N_4354);
xnor U4447 (N_4447,N_4273,N_4369);
nor U4448 (N_4448,N_4335,N_4327);
nor U4449 (N_4449,N_4314,N_4305);
nor U4450 (N_4450,N_4309,N_4320);
and U4451 (N_4451,N_4358,N_4270);
xor U4452 (N_4452,N_4311,N_4280);
or U4453 (N_4453,N_4307,N_4348);
nand U4454 (N_4454,N_4271,N_4343);
or U4455 (N_4455,N_4324,N_4346);
xnor U4456 (N_4456,N_4266,N_4357);
or U4457 (N_4457,N_4261,N_4263);
or U4458 (N_4458,N_4370,N_4326);
xnor U4459 (N_4459,N_4290,N_4284);
xor U4460 (N_4460,N_4256,N_4333);
and U4461 (N_4461,N_4253,N_4318);
nor U4462 (N_4462,N_4288,N_4335);
nand U4463 (N_4463,N_4365,N_4267);
or U4464 (N_4464,N_4371,N_4301);
and U4465 (N_4465,N_4314,N_4332);
nand U4466 (N_4466,N_4334,N_4316);
and U4467 (N_4467,N_4366,N_4298);
and U4468 (N_4468,N_4255,N_4349);
nand U4469 (N_4469,N_4355,N_4316);
nor U4470 (N_4470,N_4341,N_4274);
and U4471 (N_4471,N_4326,N_4267);
or U4472 (N_4472,N_4374,N_4328);
nor U4473 (N_4473,N_4254,N_4274);
or U4474 (N_4474,N_4332,N_4322);
and U4475 (N_4475,N_4260,N_4369);
xnor U4476 (N_4476,N_4279,N_4327);
nand U4477 (N_4477,N_4320,N_4354);
xnor U4478 (N_4478,N_4373,N_4374);
and U4479 (N_4479,N_4263,N_4331);
nor U4480 (N_4480,N_4356,N_4334);
or U4481 (N_4481,N_4266,N_4317);
or U4482 (N_4482,N_4320,N_4331);
and U4483 (N_4483,N_4266,N_4360);
nor U4484 (N_4484,N_4326,N_4368);
nand U4485 (N_4485,N_4263,N_4257);
or U4486 (N_4486,N_4305,N_4251);
nor U4487 (N_4487,N_4309,N_4335);
xor U4488 (N_4488,N_4371,N_4372);
and U4489 (N_4489,N_4334,N_4363);
nand U4490 (N_4490,N_4329,N_4321);
nor U4491 (N_4491,N_4313,N_4299);
or U4492 (N_4492,N_4352,N_4328);
or U4493 (N_4493,N_4341,N_4270);
nor U4494 (N_4494,N_4364,N_4348);
nor U4495 (N_4495,N_4255,N_4338);
and U4496 (N_4496,N_4362,N_4272);
or U4497 (N_4497,N_4367,N_4368);
or U4498 (N_4498,N_4325,N_4343);
and U4499 (N_4499,N_4259,N_4300);
nand U4500 (N_4500,N_4490,N_4458);
xor U4501 (N_4501,N_4404,N_4447);
nor U4502 (N_4502,N_4461,N_4464);
nor U4503 (N_4503,N_4474,N_4479);
or U4504 (N_4504,N_4389,N_4439);
or U4505 (N_4505,N_4489,N_4408);
and U4506 (N_4506,N_4432,N_4418);
and U4507 (N_4507,N_4440,N_4397);
xor U4508 (N_4508,N_4423,N_4495);
nand U4509 (N_4509,N_4394,N_4415);
xnor U4510 (N_4510,N_4409,N_4485);
nand U4511 (N_4511,N_4488,N_4421);
or U4512 (N_4512,N_4426,N_4417);
nand U4513 (N_4513,N_4497,N_4449);
or U4514 (N_4514,N_4414,N_4403);
nand U4515 (N_4515,N_4399,N_4400);
nor U4516 (N_4516,N_4377,N_4435);
nor U4517 (N_4517,N_4473,N_4407);
xor U4518 (N_4518,N_4442,N_4430);
nor U4519 (N_4519,N_4451,N_4422);
xnor U4520 (N_4520,N_4445,N_4446);
nor U4521 (N_4521,N_4454,N_4481);
nor U4522 (N_4522,N_4405,N_4390);
nand U4523 (N_4523,N_4386,N_4378);
nand U4524 (N_4524,N_4455,N_4427);
xnor U4525 (N_4525,N_4463,N_4385);
nor U4526 (N_4526,N_4460,N_4484);
nand U4527 (N_4527,N_4387,N_4483);
xnor U4528 (N_4528,N_4406,N_4482);
xnor U4529 (N_4529,N_4496,N_4491);
or U4530 (N_4530,N_4410,N_4382);
xor U4531 (N_4531,N_4487,N_4453);
nor U4532 (N_4532,N_4393,N_4467);
and U4533 (N_4533,N_4499,N_4469);
xor U4534 (N_4534,N_4416,N_4480);
nand U4535 (N_4535,N_4425,N_4420);
nand U4536 (N_4536,N_4424,N_4450);
nand U4537 (N_4537,N_4429,N_4438);
xor U4538 (N_4538,N_4478,N_4401);
xor U4539 (N_4539,N_4498,N_4457);
nand U4540 (N_4540,N_4470,N_4379);
and U4541 (N_4541,N_4402,N_4412);
xnor U4542 (N_4542,N_4441,N_4468);
xnor U4543 (N_4543,N_4392,N_4396);
and U4544 (N_4544,N_4471,N_4444);
or U4545 (N_4545,N_4398,N_4493);
nand U4546 (N_4546,N_4434,N_4465);
or U4547 (N_4547,N_4431,N_4383);
nand U4548 (N_4548,N_4436,N_4384);
nor U4549 (N_4549,N_4492,N_4437);
nor U4550 (N_4550,N_4475,N_4388);
nor U4551 (N_4551,N_4462,N_4433);
xor U4552 (N_4552,N_4376,N_4477);
nor U4553 (N_4553,N_4381,N_4428);
nor U4554 (N_4554,N_4459,N_4380);
xor U4555 (N_4555,N_4472,N_4448);
xnor U4556 (N_4556,N_4486,N_4476);
and U4557 (N_4557,N_4443,N_4494);
or U4558 (N_4558,N_4452,N_4466);
or U4559 (N_4559,N_4391,N_4419);
nand U4560 (N_4560,N_4395,N_4411);
nand U4561 (N_4561,N_4375,N_4413);
and U4562 (N_4562,N_4456,N_4479);
nor U4563 (N_4563,N_4450,N_4415);
and U4564 (N_4564,N_4435,N_4495);
nor U4565 (N_4565,N_4399,N_4402);
nand U4566 (N_4566,N_4390,N_4380);
and U4567 (N_4567,N_4499,N_4377);
or U4568 (N_4568,N_4396,N_4388);
nand U4569 (N_4569,N_4404,N_4446);
or U4570 (N_4570,N_4410,N_4396);
nand U4571 (N_4571,N_4481,N_4485);
xnor U4572 (N_4572,N_4426,N_4421);
xnor U4573 (N_4573,N_4437,N_4484);
or U4574 (N_4574,N_4466,N_4414);
nor U4575 (N_4575,N_4460,N_4487);
and U4576 (N_4576,N_4487,N_4416);
and U4577 (N_4577,N_4492,N_4377);
nand U4578 (N_4578,N_4445,N_4394);
or U4579 (N_4579,N_4439,N_4377);
nand U4580 (N_4580,N_4421,N_4394);
nand U4581 (N_4581,N_4498,N_4452);
or U4582 (N_4582,N_4466,N_4459);
xor U4583 (N_4583,N_4480,N_4499);
nand U4584 (N_4584,N_4437,N_4416);
or U4585 (N_4585,N_4382,N_4381);
nor U4586 (N_4586,N_4400,N_4421);
nand U4587 (N_4587,N_4404,N_4459);
and U4588 (N_4588,N_4434,N_4436);
nor U4589 (N_4589,N_4458,N_4422);
and U4590 (N_4590,N_4476,N_4442);
nand U4591 (N_4591,N_4426,N_4431);
nand U4592 (N_4592,N_4388,N_4418);
xor U4593 (N_4593,N_4391,N_4476);
nand U4594 (N_4594,N_4449,N_4420);
nand U4595 (N_4595,N_4376,N_4454);
nor U4596 (N_4596,N_4442,N_4402);
nor U4597 (N_4597,N_4466,N_4375);
or U4598 (N_4598,N_4386,N_4461);
nor U4599 (N_4599,N_4449,N_4463);
and U4600 (N_4600,N_4474,N_4401);
nand U4601 (N_4601,N_4406,N_4451);
xnor U4602 (N_4602,N_4387,N_4424);
and U4603 (N_4603,N_4388,N_4399);
nand U4604 (N_4604,N_4445,N_4487);
or U4605 (N_4605,N_4401,N_4441);
xnor U4606 (N_4606,N_4433,N_4394);
or U4607 (N_4607,N_4474,N_4399);
or U4608 (N_4608,N_4420,N_4415);
or U4609 (N_4609,N_4469,N_4460);
xor U4610 (N_4610,N_4429,N_4413);
nor U4611 (N_4611,N_4378,N_4443);
or U4612 (N_4612,N_4385,N_4429);
xor U4613 (N_4613,N_4433,N_4395);
or U4614 (N_4614,N_4437,N_4395);
nand U4615 (N_4615,N_4389,N_4450);
xnor U4616 (N_4616,N_4494,N_4391);
nand U4617 (N_4617,N_4446,N_4491);
and U4618 (N_4618,N_4476,N_4449);
and U4619 (N_4619,N_4428,N_4423);
or U4620 (N_4620,N_4483,N_4383);
nor U4621 (N_4621,N_4417,N_4433);
nor U4622 (N_4622,N_4393,N_4391);
nor U4623 (N_4623,N_4418,N_4395);
nand U4624 (N_4624,N_4470,N_4408);
xnor U4625 (N_4625,N_4580,N_4570);
and U4626 (N_4626,N_4562,N_4583);
or U4627 (N_4627,N_4572,N_4536);
and U4628 (N_4628,N_4526,N_4531);
xor U4629 (N_4629,N_4523,N_4578);
xor U4630 (N_4630,N_4524,N_4597);
nor U4631 (N_4631,N_4582,N_4588);
and U4632 (N_4632,N_4587,N_4603);
and U4633 (N_4633,N_4615,N_4514);
nand U4634 (N_4634,N_4528,N_4507);
nor U4635 (N_4635,N_4547,N_4569);
or U4636 (N_4636,N_4612,N_4533);
nor U4637 (N_4637,N_4609,N_4563);
nor U4638 (N_4638,N_4561,N_4596);
and U4639 (N_4639,N_4584,N_4558);
nor U4640 (N_4640,N_4599,N_4618);
nand U4641 (N_4641,N_4513,N_4503);
and U4642 (N_4642,N_4559,N_4517);
nor U4643 (N_4643,N_4568,N_4617);
or U4644 (N_4644,N_4532,N_4508);
xor U4645 (N_4645,N_4549,N_4548);
xnor U4646 (N_4646,N_4607,N_4519);
or U4647 (N_4647,N_4576,N_4571);
xnor U4648 (N_4648,N_4622,N_4520);
or U4649 (N_4649,N_4619,N_4606);
nand U4650 (N_4650,N_4598,N_4504);
nor U4651 (N_4651,N_4616,N_4539);
nor U4652 (N_4652,N_4610,N_4564);
or U4653 (N_4653,N_4541,N_4511);
nor U4654 (N_4654,N_4567,N_4574);
and U4655 (N_4655,N_4542,N_4518);
xnor U4656 (N_4656,N_4579,N_4577);
nand U4657 (N_4657,N_4509,N_4546);
xor U4658 (N_4658,N_4553,N_4543);
nand U4659 (N_4659,N_4534,N_4613);
nor U4660 (N_4660,N_4557,N_4620);
and U4661 (N_4661,N_4594,N_4611);
nand U4662 (N_4662,N_4510,N_4551);
or U4663 (N_4663,N_4555,N_4595);
xor U4664 (N_4664,N_4614,N_4565);
nand U4665 (N_4665,N_4601,N_4624);
or U4666 (N_4666,N_4527,N_4538);
nand U4667 (N_4667,N_4581,N_4589);
xnor U4668 (N_4668,N_4525,N_4545);
and U4669 (N_4669,N_4593,N_4590);
nor U4670 (N_4670,N_4586,N_4604);
xor U4671 (N_4671,N_4537,N_4522);
or U4672 (N_4672,N_4550,N_4575);
or U4673 (N_4673,N_4530,N_4556);
and U4674 (N_4674,N_4552,N_4623);
nand U4675 (N_4675,N_4592,N_4573);
and U4676 (N_4676,N_4560,N_4591);
or U4677 (N_4677,N_4535,N_4512);
and U4678 (N_4678,N_4501,N_4521);
or U4679 (N_4679,N_4515,N_4600);
xor U4680 (N_4680,N_4554,N_4544);
nor U4681 (N_4681,N_4605,N_4566);
nand U4682 (N_4682,N_4529,N_4608);
or U4683 (N_4683,N_4585,N_4602);
xnor U4684 (N_4684,N_4502,N_4506);
nor U4685 (N_4685,N_4540,N_4500);
and U4686 (N_4686,N_4505,N_4516);
xnor U4687 (N_4687,N_4621,N_4595);
or U4688 (N_4688,N_4587,N_4567);
or U4689 (N_4689,N_4537,N_4591);
nor U4690 (N_4690,N_4583,N_4507);
or U4691 (N_4691,N_4517,N_4624);
nand U4692 (N_4692,N_4511,N_4590);
xor U4693 (N_4693,N_4554,N_4531);
nand U4694 (N_4694,N_4538,N_4523);
nor U4695 (N_4695,N_4533,N_4592);
and U4696 (N_4696,N_4539,N_4526);
nor U4697 (N_4697,N_4525,N_4570);
xnor U4698 (N_4698,N_4510,N_4604);
or U4699 (N_4699,N_4612,N_4539);
and U4700 (N_4700,N_4537,N_4571);
xnor U4701 (N_4701,N_4559,N_4552);
and U4702 (N_4702,N_4561,N_4578);
nor U4703 (N_4703,N_4567,N_4591);
xnor U4704 (N_4704,N_4566,N_4571);
and U4705 (N_4705,N_4621,N_4527);
nand U4706 (N_4706,N_4592,N_4524);
nand U4707 (N_4707,N_4554,N_4514);
nor U4708 (N_4708,N_4521,N_4539);
nor U4709 (N_4709,N_4573,N_4514);
and U4710 (N_4710,N_4508,N_4520);
nor U4711 (N_4711,N_4508,N_4536);
nand U4712 (N_4712,N_4561,N_4502);
nand U4713 (N_4713,N_4617,N_4511);
nor U4714 (N_4714,N_4509,N_4576);
and U4715 (N_4715,N_4601,N_4565);
or U4716 (N_4716,N_4597,N_4595);
and U4717 (N_4717,N_4614,N_4518);
nand U4718 (N_4718,N_4534,N_4564);
or U4719 (N_4719,N_4583,N_4510);
and U4720 (N_4720,N_4600,N_4507);
and U4721 (N_4721,N_4614,N_4529);
nor U4722 (N_4722,N_4543,N_4621);
and U4723 (N_4723,N_4515,N_4562);
or U4724 (N_4724,N_4585,N_4553);
or U4725 (N_4725,N_4541,N_4549);
or U4726 (N_4726,N_4602,N_4555);
nand U4727 (N_4727,N_4608,N_4552);
xnor U4728 (N_4728,N_4623,N_4594);
nor U4729 (N_4729,N_4533,N_4504);
or U4730 (N_4730,N_4598,N_4537);
nor U4731 (N_4731,N_4501,N_4545);
xor U4732 (N_4732,N_4559,N_4570);
or U4733 (N_4733,N_4532,N_4528);
xor U4734 (N_4734,N_4526,N_4551);
or U4735 (N_4735,N_4523,N_4504);
nor U4736 (N_4736,N_4576,N_4534);
and U4737 (N_4737,N_4601,N_4599);
xor U4738 (N_4738,N_4541,N_4574);
or U4739 (N_4739,N_4561,N_4576);
or U4740 (N_4740,N_4543,N_4515);
xnor U4741 (N_4741,N_4621,N_4545);
xnor U4742 (N_4742,N_4518,N_4508);
or U4743 (N_4743,N_4554,N_4539);
nand U4744 (N_4744,N_4514,N_4526);
and U4745 (N_4745,N_4610,N_4566);
nand U4746 (N_4746,N_4597,N_4504);
nand U4747 (N_4747,N_4515,N_4511);
nor U4748 (N_4748,N_4547,N_4564);
nor U4749 (N_4749,N_4605,N_4587);
and U4750 (N_4750,N_4685,N_4671);
or U4751 (N_4751,N_4731,N_4662);
and U4752 (N_4752,N_4655,N_4735);
xor U4753 (N_4753,N_4670,N_4716);
nand U4754 (N_4754,N_4708,N_4626);
xnor U4755 (N_4755,N_4637,N_4741);
and U4756 (N_4756,N_4669,N_4684);
nor U4757 (N_4757,N_4678,N_4640);
and U4758 (N_4758,N_4635,N_4701);
xor U4759 (N_4759,N_4725,N_4694);
or U4760 (N_4760,N_4665,N_4718);
and U4761 (N_4761,N_4703,N_4729);
xor U4762 (N_4762,N_4642,N_4636);
xor U4763 (N_4763,N_4667,N_4742);
xor U4764 (N_4764,N_4668,N_4656);
xor U4765 (N_4765,N_4714,N_4720);
and U4766 (N_4766,N_4739,N_4747);
xnor U4767 (N_4767,N_4641,N_4664);
xor U4768 (N_4768,N_4730,N_4632);
nand U4769 (N_4769,N_4659,N_4650);
nand U4770 (N_4770,N_4709,N_4674);
nand U4771 (N_4771,N_4738,N_4746);
and U4772 (N_4772,N_4724,N_4692);
xnor U4773 (N_4773,N_4732,N_4745);
or U4774 (N_4774,N_4657,N_4629);
nor U4775 (N_4775,N_4712,N_4643);
or U4776 (N_4776,N_4706,N_4699);
or U4777 (N_4777,N_4689,N_4644);
xnor U4778 (N_4778,N_4722,N_4663);
or U4779 (N_4779,N_4700,N_4660);
or U4780 (N_4780,N_4680,N_4697);
xnor U4781 (N_4781,N_4649,N_4707);
and U4782 (N_4782,N_4717,N_4740);
nand U4783 (N_4783,N_4625,N_4744);
and U4784 (N_4784,N_4723,N_4683);
nor U4785 (N_4785,N_4726,N_4727);
or U4786 (N_4786,N_4628,N_4690);
nor U4787 (N_4787,N_4654,N_4666);
nand U4788 (N_4788,N_4695,N_4719);
or U4789 (N_4789,N_4711,N_4630);
xor U4790 (N_4790,N_4702,N_4710);
xor U4791 (N_4791,N_4715,N_4653);
and U4792 (N_4792,N_4652,N_4661);
nor U4793 (N_4793,N_4728,N_4639);
nor U4794 (N_4794,N_4672,N_4749);
or U4795 (N_4795,N_4658,N_4704);
nand U4796 (N_4796,N_4688,N_4638);
xnor U4797 (N_4797,N_4627,N_4691);
and U4798 (N_4798,N_4673,N_4698);
nand U4799 (N_4799,N_4648,N_4676);
and U4800 (N_4800,N_4693,N_4696);
and U4801 (N_4801,N_4736,N_4713);
nor U4802 (N_4802,N_4743,N_4647);
nand U4803 (N_4803,N_4733,N_4645);
nand U4804 (N_4804,N_4679,N_4634);
or U4805 (N_4805,N_4651,N_4705);
nand U4806 (N_4806,N_4737,N_4682);
nor U4807 (N_4807,N_4677,N_4721);
nor U4808 (N_4808,N_4633,N_4646);
xnor U4809 (N_4809,N_4631,N_4734);
nor U4810 (N_4810,N_4748,N_4687);
xnor U4811 (N_4811,N_4686,N_4681);
or U4812 (N_4812,N_4675,N_4726);
xor U4813 (N_4813,N_4662,N_4714);
nand U4814 (N_4814,N_4706,N_4740);
and U4815 (N_4815,N_4647,N_4673);
nor U4816 (N_4816,N_4681,N_4737);
xnor U4817 (N_4817,N_4733,N_4714);
xor U4818 (N_4818,N_4726,N_4719);
or U4819 (N_4819,N_4684,N_4632);
xnor U4820 (N_4820,N_4731,N_4692);
nor U4821 (N_4821,N_4701,N_4741);
nand U4822 (N_4822,N_4627,N_4651);
or U4823 (N_4823,N_4625,N_4722);
nor U4824 (N_4824,N_4645,N_4675);
nand U4825 (N_4825,N_4726,N_4664);
or U4826 (N_4826,N_4650,N_4635);
and U4827 (N_4827,N_4709,N_4728);
or U4828 (N_4828,N_4713,N_4678);
and U4829 (N_4829,N_4749,N_4715);
nand U4830 (N_4830,N_4680,N_4643);
nand U4831 (N_4831,N_4717,N_4695);
and U4832 (N_4832,N_4736,N_4687);
nand U4833 (N_4833,N_4701,N_4712);
and U4834 (N_4834,N_4625,N_4710);
nor U4835 (N_4835,N_4635,N_4689);
or U4836 (N_4836,N_4725,N_4628);
or U4837 (N_4837,N_4719,N_4690);
xnor U4838 (N_4838,N_4634,N_4693);
xnor U4839 (N_4839,N_4644,N_4641);
nand U4840 (N_4840,N_4683,N_4680);
or U4841 (N_4841,N_4698,N_4664);
nand U4842 (N_4842,N_4739,N_4730);
and U4843 (N_4843,N_4655,N_4635);
xnor U4844 (N_4844,N_4655,N_4689);
and U4845 (N_4845,N_4748,N_4725);
or U4846 (N_4846,N_4690,N_4657);
and U4847 (N_4847,N_4682,N_4742);
and U4848 (N_4848,N_4708,N_4633);
nand U4849 (N_4849,N_4658,N_4705);
or U4850 (N_4850,N_4650,N_4673);
xor U4851 (N_4851,N_4632,N_4627);
and U4852 (N_4852,N_4749,N_4713);
nor U4853 (N_4853,N_4734,N_4727);
and U4854 (N_4854,N_4735,N_4722);
nor U4855 (N_4855,N_4643,N_4727);
nor U4856 (N_4856,N_4709,N_4732);
nor U4857 (N_4857,N_4699,N_4710);
or U4858 (N_4858,N_4656,N_4632);
nor U4859 (N_4859,N_4711,N_4740);
or U4860 (N_4860,N_4702,N_4645);
nor U4861 (N_4861,N_4679,N_4652);
xor U4862 (N_4862,N_4726,N_4658);
nor U4863 (N_4863,N_4702,N_4697);
and U4864 (N_4864,N_4699,N_4748);
xnor U4865 (N_4865,N_4678,N_4734);
nor U4866 (N_4866,N_4660,N_4637);
xor U4867 (N_4867,N_4665,N_4676);
and U4868 (N_4868,N_4651,N_4644);
xor U4869 (N_4869,N_4643,N_4718);
nand U4870 (N_4870,N_4679,N_4675);
and U4871 (N_4871,N_4734,N_4724);
or U4872 (N_4872,N_4674,N_4710);
nand U4873 (N_4873,N_4708,N_4630);
xor U4874 (N_4874,N_4689,N_4629);
nand U4875 (N_4875,N_4776,N_4861);
or U4876 (N_4876,N_4765,N_4777);
xnor U4877 (N_4877,N_4780,N_4805);
xor U4878 (N_4878,N_4864,N_4751);
or U4879 (N_4879,N_4827,N_4796);
and U4880 (N_4880,N_4781,N_4753);
nor U4881 (N_4881,N_4823,N_4755);
xnor U4882 (N_4882,N_4820,N_4871);
and U4883 (N_4883,N_4803,N_4788);
nor U4884 (N_4884,N_4815,N_4854);
nor U4885 (N_4885,N_4873,N_4760);
nand U4886 (N_4886,N_4822,N_4817);
or U4887 (N_4887,N_4791,N_4858);
nor U4888 (N_4888,N_4774,N_4869);
xnor U4889 (N_4889,N_4834,N_4789);
xnor U4890 (N_4890,N_4838,N_4856);
or U4891 (N_4891,N_4830,N_4860);
nand U4892 (N_4892,N_4851,N_4779);
or U4893 (N_4893,N_4752,N_4802);
and U4894 (N_4894,N_4850,N_4835);
nand U4895 (N_4895,N_4841,N_4792);
nor U4896 (N_4896,N_4813,N_4800);
nor U4897 (N_4897,N_4868,N_4794);
nand U4898 (N_4898,N_4865,N_4846);
or U4899 (N_4899,N_4787,N_4872);
or U4900 (N_4900,N_4754,N_4855);
nor U4901 (N_4901,N_4811,N_4843);
and U4902 (N_4902,N_4784,N_4763);
or U4903 (N_4903,N_4766,N_4839);
or U4904 (N_4904,N_4769,N_4764);
or U4905 (N_4905,N_4842,N_4867);
nand U4906 (N_4906,N_4863,N_4825);
xor U4907 (N_4907,N_4808,N_4810);
nor U4908 (N_4908,N_4826,N_4819);
nand U4909 (N_4909,N_4828,N_4773);
nand U4910 (N_4910,N_4845,N_4804);
xnor U4911 (N_4911,N_4829,N_4833);
nor U4912 (N_4912,N_4785,N_4836);
and U4913 (N_4913,N_4853,N_4757);
nand U4914 (N_4914,N_4756,N_4807);
nand U4915 (N_4915,N_4852,N_4772);
nand U4916 (N_4916,N_4832,N_4783);
nand U4917 (N_4917,N_4775,N_4818);
nor U4918 (N_4918,N_4844,N_4768);
or U4919 (N_4919,N_4857,N_4801);
nor U4920 (N_4920,N_4874,N_4790);
and U4921 (N_4921,N_4859,N_4762);
nor U4922 (N_4922,N_4750,N_4816);
nor U4923 (N_4923,N_4795,N_4761);
nand U4924 (N_4924,N_4809,N_4782);
or U4925 (N_4925,N_4824,N_4831);
or U4926 (N_4926,N_4758,N_4821);
xnor U4927 (N_4927,N_4799,N_4798);
nor U4928 (N_4928,N_4849,N_4814);
and U4929 (N_4929,N_4866,N_4812);
and U4930 (N_4930,N_4862,N_4837);
and U4931 (N_4931,N_4806,N_4847);
xnor U4932 (N_4932,N_4840,N_4778);
and U4933 (N_4933,N_4848,N_4770);
xor U4934 (N_4934,N_4759,N_4771);
nor U4935 (N_4935,N_4767,N_4793);
nand U4936 (N_4936,N_4797,N_4786);
nand U4937 (N_4937,N_4870,N_4756);
nand U4938 (N_4938,N_4843,N_4832);
or U4939 (N_4939,N_4836,N_4792);
nand U4940 (N_4940,N_4816,N_4862);
nor U4941 (N_4941,N_4807,N_4864);
and U4942 (N_4942,N_4798,N_4858);
nor U4943 (N_4943,N_4769,N_4760);
nand U4944 (N_4944,N_4779,N_4801);
or U4945 (N_4945,N_4834,N_4858);
xnor U4946 (N_4946,N_4779,N_4759);
or U4947 (N_4947,N_4861,N_4791);
xnor U4948 (N_4948,N_4814,N_4752);
and U4949 (N_4949,N_4863,N_4807);
or U4950 (N_4950,N_4866,N_4859);
or U4951 (N_4951,N_4856,N_4761);
nand U4952 (N_4952,N_4862,N_4802);
nor U4953 (N_4953,N_4792,N_4774);
nor U4954 (N_4954,N_4787,N_4777);
nor U4955 (N_4955,N_4816,N_4780);
and U4956 (N_4956,N_4802,N_4869);
nor U4957 (N_4957,N_4851,N_4872);
or U4958 (N_4958,N_4795,N_4816);
or U4959 (N_4959,N_4859,N_4850);
nor U4960 (N_4960,N_4822,N_4752);
nand U4961 (N_4961,N_4812,N_4846);
nor U4962 (N_4962,N_4854,N_4774);
nand U4963 (N_4963,N_4852,N_4784);
or U4964 (N_4964,N_4765,N_4781);
and U4965 (N_4965,N_4819,N_4762);
xnor U4966 (N_4966,N_4791,N_4860);
or U4967 (N_4967,N_4756,N_4801);
or U4968 (N_4968,N_4824,N_4855);
or U4969 (N_4969,N_4802,N_4805);
nor U4970 (N_4970,N_4798,N_4829);
xor U4971 (N_4971,N_4829,N_4786);
nand U4972 (N_4972,N_4799,N_4762);
nand U4973 (N_4973,N_4782,N_4838);
nand U4974 (N_4974,N_4839,N_4764);
xnor U4975 (N_4975,N_4849,N_4805);
nand U4976 (N_4976,N_4863,N_4854);
nor U4977 (N_4977,N_4771,N_4751);
nand U4978 (N_4978,N_4853,N_4784);
or U4979 (N_4979,N_4770,N_4835);
nor U4980 (N_4980,N_4860,N_4852);
nor U4981 (N_4981,N_4757,N_4856);
and U4982 (N_4982,N_4787,N_4810);
xnor U4983 (N_4983,N_4815,N_4784);
or U4984 (N_4984,N_4751,N_4795);
nand U4985 (N_4985,N_4843,N_4790);
nor U4986 (N_4986,N_4782,N_4825);
nand U4987 (N_4987,N_4757,N_4800);
and U4988 (N_4988,N_4856,N_4841);
nor U4989 (N_4989,N_4815,N_4754);
nand U4990 (N_4990,N_4828,N_4752);
nand U4991 (N_4991,N_4775,N_4782);
and U4992 (N_4992,N_4790,N_4751);
or U4993 (N_4993,N_4861,N_4784);
and U4994 (N_4994,N_4864,N_4799);
or U4995 (N_4995,N_4863,N_4860);
xor U4996 (N_4996,N_4771,N_4866);
xnor U4997 (N_4997,N_4824,N_4854);
and U4998 (N_4998,N_4798,N_4824);
or U4999 (N_4999,N_4770,N_4808);
nand U5000 (N_5000,N_4992,N_4963);
xor U5001 (N_5001,N_4927,N_4991);
nor U5002 (N_5002,N_4977,N_4984);
nand U5003 (N_5003,N_4897,N_4983);
and U5004 (N_5004,N_4907,N_4911);
xnor U5005 (N_5005,N_4995,N_4885);
nand U5006 (N_5006,N_4890,N_4878);
xnor U5007 (N_5007,N_4945,N_4894);
and U5008 (N_5008,N_4950,N_4930);
nor U5009 (N_5009,N_4994,N_4981);
xnor U5010 (N_5010,N_4923,N_4875);
nand U5011 (N_5011,N_4975,N_4880);
or U5012 (N_5012,N_4958,N_4899);
nand U5013 (N_5013,N_4989,N_4957);
nand U5014 (N_5014,N_4956,N_4943);
xor U5015 (N_5015,N_4931,N_4969);
xnor U5016 (N_5016,N_4920,N_4908);
and U5017 (N_5017,N_4925,N_4881);
and U5018 (N_5018,N_4997,N_4948);
nand U5019 (N_5019,N_4993,N_4888);
xor U5020 (N_5020,N_4909,N_4936);
nor U5021 (N_5021,N_4966,N_4924);
nor U5022 (N_5022,N_4998,N_4971);
or U5023 (N_5023,N_4987,N_4941);
or U5024 (N_5024,N_4973,N_4976);
and U5025 (N_5025,N_4999,N_4882);
or U5026 (N_5026,N_4938,N_4972);
nor U5027 (N_5027,N_4900,N_4940);
xor U5028 (N_5028,N_4955,N_4944);
nand U5029 (N_5029,N_4921,N_4906);
nand U5030 (N_5030,N_4903,N_4961);
or U5031 (N_5031,N_4967,N_4954);
or U5032 (N_5032,N_4928,N_4946);
or U5033 (N_5033,N_4985,N_4883);
xnor U5034 (N_5034,N_4922,N_4951);
xor U5035 (N_5035,N_4902,N_4913);
and U5036 (N_5036,N_4926,N_4974);
nand U5037 (N_5037,N_4953,N_4935);
xor U5038 (N_5038,N_4978,N_4949);
or U5039 (N_5039,N_4996,N_4916);
nand U5040 (N_5040,N_4877,N_4889);
and U5041 (N_5041,N_4988,N_4947);
and U5042 (N_5042,N_4905,N_4917);
xor U5043 (N_5043,N_4915,N_4879);
or U5044 (N_5044,N_4970,N_4895);
or U5045 (N_5045,N_4968,N_4962);
nor U5046 (N_5046,N_4937,N_4964);
or U5047 (N_5047,N_4965,N_4904);
nor U5048 (N_5048,N_4918,N_4979);
nand U5049 (N_5049,N_4942,N_4896);
and U5050 (N_5050,N_4914,N_4898);
nor U5051 (N_5051,N_4910,N_4933);
nor U5052 (N_5052,N_4980,N_4892);
nor U5053 (N_5053,N_4982,N_4876);
or U5054 (N_5054,N_4893,N_4960);
nand U5055 (N_5055,N_4912,N_4929);
xnor U5056 (N_5056,N_4932,N_4886);
xnor U5057 (N_5057,N_4884,N_4901);
or U5058 (N_5058,N_4990,N_4986);
and U5059 (N_5059,N_4939,N_4934);
xor U5060 (N_5060,N_4919,N_4952);
or U5061 (N_5061,N_4887,N_4959);
or U5062 (N_5062,N_4891,N_4912);
nand U5063 (N_5063,N_4904,N_4993);
nand U5064 (N_5064,N_4935,N_4932);
xnor U5065 (N_5065,N_4996,N_4933);
nand U5066 (N_5066,N_4951,N_4902);
nor U5067 (N_5067,N_4979,N_4881);
and U5068 (N_5068,N_4889,N_4880);
and U5069 (N_5069,N_4959,N_4922);
xor U5070 (N_5070,N_4924,N_4887);
or U5071 (N_5071,N_4948,N_4913);
and U5072 (N_5072,N_4927,N_4887);
and U5073 (N_5073,N_4996,N_4958);
nor U5074 (N_5074,N_4967,N_4973);
nand U5075 (N_5075,N_4958,N_4897);
nand U5076 (N_5076,N_4944,N_4981);
xnor U5077 (N_5077,N_4896,N_4968);
or U5078 (N_5078,N_4968,N_4888);
xnor U5079 (N_5079,N_4925,N_4923);
xnor U5080 (N_5080,N_4968,N_4904);
nand U5081 (N_5081,N_4960,N_4938);
and U5082 (N_5082,N_4971,N_4941);
xnor U5083 (N_5083,N_4928,N_4959);
nor U5084 (N_5084,N_4936,N_4993);
xor U5085 (N_5085,N_4880,N_4901);
xor U5086 (N_5086,N_4985,N_4922);
nand U5087 (N_5087,N_4912,N_4979);
or U5088 (N_5088,N_4892,N_4927);
xnor U5089 (N_5089,N_4876,N_4992);
xnor U5090 (N_5090,N_4876,N_4980);
or U5091 (N_5091,N_4933,N_4891);
nor U5092 (N_5092,N_4926,N_4934);
xor U5093 (N_5093,N_4878,N_4978);
or U5094 (N_5094,N_4962,N_4929);
nor U5095 (N_5095,N_4915,N_4919);
and U5096 (N_5096,N_4876,N_4975);
nand U5097 (N_5097,N_4976,N_4885);
and U5098 (N_5098,N_4974,N_4885);
and U5099 (N_5099,N_4966,N_4974);
nor U5100 (N_5100,N_4886,N_4958);
or U5101 (N_5101,N_4883,N_4968);
xnor U5102 (N_5102,N_4973,N_4939);
and U5103 (N_5103,N_4936,N_4958);
nand U5104 (N_5104,N_4886,N_4920);
or U5105 (N_5105,N_4938,N_4965);
or U5106 (N_5106,N_4946,N_4885);
xnor U5107 (N_5107,N_4959,N_4895);
or U5108 (N_5108,N_4947,N_4904);
nor U5109 (N_5109,N_4999,N_4956);
xor U5110 (N_5110,N_4977,N_4904);
or U5111 (N_5111,N_4953,N_4973);
or U5112 (N_5112,N_4888,N_4990);
nor U5113 (N_5113,N_4952,N_4898);
or U5114 (N_5114,N_4940,N_4957);
or U5115 (N_5115,N_4912,N_4993);
and U5116 (N_5116,N_4942,N_4975);
or U5117 (N_5117,N_4883,N_4928);
nand U5118 (N_5118,N_4991,N_4894);
nand U5119 (N_5119,N_4961,N_4881);
nand U5120 (N_5120,N_4930,N_4878);
and U5121 (N_5121,N_4902,N_4884);
nor U5122 (N_5122,N_4952,N_4893);
nor U5123 (N_5123,N_4930,N_4934);
and U5124 (N_5124,N_4896,N_4969);
nand U5125 (N_5125,N_5038,N_5104);
and U5126 (N_5126,N_5082,N_5040);
nor U5127 (N_5127,N_5019,N_5045);
xnor U5128 (N_5128,N_5120,N_5003);
and U5129 (N_5129,N_5058,N_5077);
nand U5130 (N_5130,N_5026,N_5053);
and U5131 (N_5131,N_5081,N_5029);
nand U5132 (N_5132,N_5076,N_5094);
and U5133 (N_5133,N_5044,N_5123);
xnor U5134 (N_5134,N_5075,N_5013);
nand U5135 (N_5135,N_5032,N_5011);
nor U5136 (N_5136,N_5052,N_5031);
or U5137 (N_5137,N_5116,N_5014);
or U5138 (N_5138,N_5096,N_5064);
nand U5139 (N_5139,N_5004,N_5056);
xnor U5140 (N_5140,N_5102,N_5110);
xor U5141 (N_5141,N_5118,N_5095);
xor U5142 (N_5142,N_5054,N_5039);
nor U5143 (N_5143,N_5080,N_5068);
nor U5144 (N_5144,N_5018,N_5061);
nand U5145 (N_5145,N_5106,N_5103);
and U5146 (N_5146,N_5049,N_5017);
nor U5147 (N_5147,N_5041,N_5067);
nand U5148 (N_5148,N_5122,N_5105);
xnor U5149 (N_5149,N_5022,N_5083);
or U5150 (N_5150,N_5101,N_5030);
xor U5151 (N_5151,N_5078,N_5088);
xnor U5152 (N_5152,N_5009,N_5033);
nor U5153 (N_5153,N_5117,N_5050);
xor U5154 (N_5154,N_5001,N_5107);
nor U5155 (N_5155,N_5073,N_5070);
and U5156 (N_5156,N_5097,N_5113);
xor U5157 (N_5157,N_5059,N_5112);
xnor U5158 (N_5158,N_5035,N_5037);
and U5159 (N_5159,N_5006,N_5074);
xnor U5160 (N_5160,N_5066,N_5091);
nand U5161 (N_5161,N_5025,N_5002);
or U5162 (N_5162,N_5069,N_5109);
nand U5163 (N_5163,N_5089,N_5048);
and U5164 (N_5164,N_5098,N_5023);
xor U5165 (N_5165,N_5010,N_5021);
nand U5166 (N_5166,N_5020,N_5057);
or U5167 (N_5167,N_5008,N_5084);
xnor U5168 (N_5168,N_5047,N_5055);
or U5169 (N_5169,N_5119,N_5108);
nor U5170 (N_5170,N_5027,N_5036);
xnor U5171 (N_5171,N_5063,N_5079);
and U5172 (N_5172,N_5114,N_5111);
nor U5173 (N_5173,N_5072,N_5051);
or U5174 (N_5174,N_5034,N_5099);
xnor U5175 (N_5175,N_5100,N_5092);
nor U5176 (N_5176,N_5028,N_5046);
nor U5177 (N_5177,N_5115,N_5043);
nor U5178 (N_5178,N_5042,N_5065);
and U5179 (N_5179,N_5085,N_5024);
xor U5180 (N_5180,N_5016,N_5121);
nand U5181 (N_5181,N_5087,N_5093);
xor U5182 (N_5182,N_5000,N_5071);
and U5183 (N_5183,N_5124,N_5060);
nor U5184 (N_5184,N_5015,N_5090);
nand U5185 (N_5185,N_5005,N_5086);
and U5186 (N_5186,N_5062,N_5012);
and U5187 (N_5187,N_5007,N_5114);
nor U5188 (N_5188,N_5037,N_5105);
nand U5189 (N_5189,N_5055,N_5003);
nand U5190 (N_5190,N_5112,N_5074);
and U5191 (N_5191,N_5077,N_5065);
and U5192 (N_5192,N_5006,N_5047);
nor U5193 (N_5193,N_5010,N_5040);
and U5194 (N_5194,N_5112,N_5116);
nor U5195 (N_5195,N_5103,N_5094);
nand U5196 (N_5196,N_5114,N_5088);
nand U5197 (N_5197,N_5001,N_5073);
nand U5198 (N_5198,N_5083,N_5086);
xor U5199 (N_5199,N_5113,N_5064);
and U5200 (N_5200,N_5107,N_5115);
nor U5201 (N_5201,N_5078,N_5050);
or U5202 (N_5202,N_5042,N_5115);
and U5203 (N_5203,N_5100,N_5019);
nand U5204 (N_5204,N_5041,N_5058);
nor U5205 (N_5205,N_5019,N_5023);
nor U5206 (N_5206,N_5120,N_5099);
or U5207 (N_5207,N_5062,N_5112);
xor U5208 (N_5208,N_5086,N_5119);
nor U5209 (N_5209,N_5027,N_5002);
nand U5210 (N_5210,N_5004,N_5039);
xnor U5211 (N_5211,N_5061,N_5019);
nor U5212 (N_5212,N_5035,N_5095);
and U5213 (N_5213,N_5112,N_5092);
nor U5214 (N_5214,N_5026,N_5096);
and U5215 (N_5215,N_5044,N_5083);
nand U5216 (N_5216,N_5013,N_5048);
or U5217 (N_5217,N_5098,N_5039);
xnor U5218 (N_5218,N_5090,N_5068);
xor U5219 (N_5219,N_5064,N_5072);
and U5220 (N_5220,N_5076,N_5062);
xor U5221 (N_5221,N_5028,N_5103);
nand U5222 (N_5222,N_5069,N_5081);
and U5223 (N_5223,N_5067,N_5006);
and U5224 (N_5224,N_5073,N_5121);
nand U5225 (N_5225,N_5107,N_5108);
nand U5226 (N_5226,N_5028,N_5047);
nor U5227 (N_5227,N_5045,N_5054);
and U5228 (N_5228,N_5022,N_5107);
nand U5229 (N_5229,N_5085,N_5080);
nor U5230 (N_5230,N_5073,N_5057);
nand U5231 (N_5231,N_5059,N_5024);
xnor U5232 (N_5232,N_5084,N_5043);
nor U5233 (N_5233,N_5122,N_5092);
xor U5234 (N_5234,N_5091,N_5039);
nand U5235 (N_5235,N_5073,N_5023);
nor U5236 (N_5236,N_5010,N_5001);
or U5237 (N_5237,N_5011,N_5097);
or U5238 (N_5238,N_5016,N_5083);
or U5239 (N_5239,N_5023,N_5044);
nand U5240 (N_5240,N_5102,N_5004);
and U5241 (N_5241,N_5117,N_5097);
nor U5242 (N_5242,N_5057,N_5075);
nand U5243 (N_5243,N_5018,N_5087);
nor U5244 (N_5244,N_5022,N_5003);
and U5245 (N_5245,N_5043,N_5050);
nand U5246 (N_5246,N_5061,N_5033);
nor U5247 (N_5247,N_5024,N_5031);
and U5248 (N_5248,N_5052,N_5004);
and U5249 (N_5249,N_5068,N_5064);
xor U5250 (N_5250,N_5187,N_5138);
or U5251 (N_5251,N_5148,N_5128);
xnor U5252 (N_5252,N_5129,N_5243);
or U5253 (N_5253,N_5233,N_5158);
nor U5254 (N_5254,N_5212,N_5240);
nand U5255 (N_5255,N_5170,N_5226);
xnor U5256 (N_5256,N_5194,N_5225);
xnor U5257 (N_5257,N_5237,N_5159);
or U5258 (N_5258,N_5185,N_5204);
nor U5259 (N_5259,N_5244,N_5214);
nand U5260 (N_5260,N_5166,N_5169);
nor U5261 (N_5261,N_5199,N_5155);
or U5262 (N_5262,N_5189,N_5142);
and U5263 (N_5263,N_5147,N_5133);
or U5264 (N_5264,N_5134,N_5221);
and U5265 (N_5265,N_5248,N_5218);
or U5266 (N_5266,N_5247,N_5165);
and U5267 (N_5267,N_5198,N_5143);
xor U5268 (N_5268,N_5164,N_5130);
xor U5269 (N_5269,N_5172,N_5191);
xnor U5270 (N_5270,N_5127,N_5153);
and U5271 (N_5271,N_5245,N_5144);
nand U5272 (N_5272,N_5206,N_5203);
and U5273 (N_5273,N_5249,N_5180);
xnor U5274 (N_5274,N_5157,N_5241);
or U5275 (N_5275,N_5223,N_5131);
or U5276 (N_5276,N_5154,N_5176);
nand U5277 (N_5277,N_5238,N_5205);
xor U5278 (N_5278,N_5163,N_5208);
nand U5279 (N_5279,N_5232,N_5175);
nor U5280 (N_5280,N_5140,N_5246);
or U5281 (N_5281,N_5149,N_5211);
nand U5282 (N_5282,N_5196,N_5216);
nor U5283 (N_5283,N_5190,N_5227);
xnor U5284 (N_5284,N_5219,N_5224);
xor U5285 (N_5285,N_5230,N_5160);
nor U5286 (N_5286,N_5228,N_5183);
and U5287 (N_5287,N_5186,N_5222);
xor U5288 (N_5288,N_5152,N_5177);
nand U5289 (N_5289,N_5174,N_5231);
nor U5290 (N_5290,N_5178,N_5192);
nor U5291 (N_5291,N_5173,N_5146);
nand U5292 (N_5292,N_5156,N_5235);
xor U5293 (N_5293,N_5239,N_5229);
and U5294 (N_5294,N_5125,N_5236);
and U5295 (N_5295,N_5151,N_5126);
nand U5296 (N_5296,N_5184,N_5181);
nand U5297 (N_5297,N_5234,N_5193);
or U5298 (N_5298,N_5171,N_5207);
xnor U5299 (N_5299,N_5209,N_5195);
nor U5300 (N_5300,N_5202,N_5200);
or U5301 (N_5301,N_5161,N_5132);
and U5302 (N_5302,N_5141,N_5145);
and U5303 (N_5303,N_5162,N_5188);
nor U5304 (N_5304,N_5217,N_5182);
or U5305 (N_5305,N_5139,N_5201);
nand U5306 (N_5306,N_5220,N_5168);
or U5307 (N_5307,N_5242,N_5135);
or U5308 (N_5308,N_5167,N_5197);
or U5309 (N_5309,N_5179,N_5150);
nand U5310 (N_5310,N_5137,N_5210);
or U5311 (N_5311,N_5136,N_5215);
nand U5312 (N_5312,N_5213,N_5174);
and U5313 (N_5313,N_5237,N_5197);
xor U5314 (N_5314,N_5125,N_5242);
nand U5315 (N_5315,N_5226,N_5180);
xnor U5316 (N_5316,N_5178,N_5139);
nor U5317 (N_5317,N_5236,N_5160);
and U5318 (N_5318,N_5203,N_5126);
nor U5319 (N_5319,N_5175,N_5147);
xnor U5320 (N_5320,N_5233,N_5211);
or U5321 (N_5321,N_5218,N_5226);
or U5322 (N_5322,N_5161,N_5237);
xnor U5323 (N_5323,N_5155,N_5167);
nand U5324 (N_5324,N_5147,N_5161);
xnor U5325 (N_5325,N_5219,N_5168);
nor U5326 (N_5326,N_5187,N_5227);
nand U5327 (N_5327,N_5225,N_5196);
nand U5328 (N_5328,N_5224,N_5246);
nand U5329 (N_5329,N_5238,N_5178);
or U5330 (N_5330,N_5158,N_5224);
xor U5331 (N_5331,N_5157,N_5236);
xnor U5332 (N_5332,N_5231,N_5229);
or U5333 (N_5333,N_5240,N_5187);
nand U5334 (N_5334,N_5166,N_5237);
nor U5335 (N_5335,N_5137,N_5199);
and U5336 (N_5336,N_5243,N_5238);
nand U5337 (N_5337,N_5142,N_5216);
nand U5338 (N_5338,N_5151,N_5235);
xnor U5339 (N_5339,N_5242,N_5183);
nor U5340 (N_5340,N_5156,N_5167);
xnor U5341 (N_5341,N_5177,N_5249);
nor U5342 (N_5342,N_5211,N_5158);
or U5343 (N_5343,N_5221,N_5135);
xnor U5344 (N_5344,N_5225,N_5203);
xor U5345 (N_5345,N_5237,N_5238);
xor U5346 (N_5346,N_5179,N_5173);
nor U5347 (N_5347,N_5245,N_5219);
nand U5348 (N_5348,N_5227,N_5175);
and U5349 (N_5349,N_5224,N_5143);
nand U5350 (N_5350,N_5169,N_5175);
nor U5351 (N_5351,N_5210,N_5224);
nand U5352 (N_5352,N_5220,N_5166);
nor U5353 (N_5353,N_5150,N_5140);
nor U5354 (N_5354,N_5171,N_5189);
xnor U5355 (N_5355,N_5188,N_5209);
nor U5356 (N_5356,N_5140,N_5149);
xnor U5357 (N_5357,N_5156,N_5202);
or U5358 (N_5358,N_5217,N_5247);
xnor U5359 (N_5359,N_5125,N_5174);
xnor U5360 (N_5360,N_5218,N_5153);
or U5361 (N_5361,N_5233,N_5181);
xnor U5362 (N_5362,N_5161,N_5148);
or U5363 (N_5363,N_5223,N_5214);
or U5364 (N_5364,N_5157,N_5240);
and U5365 (N_5365,N_5203,N_5125);
and U5366 (N_5366,N_5249,N_5195);
and U5367 (N_5367,N_5213,N_5140);
xor U5368 (N_5368,N_5189,N_5197);
nand U5369 (N_5369,N_5132,N_5180);
or U5370 (N_5370,N_5165,N_5130);
xor U5371 (N_5371,N_5214,N_5196);
nor U5372 (N_5372,N_5214,N_5158);
nand U5373 (N_5373,N_5211,N_5217);
and U5374 (N_5374,N_5153,N_5132);
and U5375 (N_5375,N_5362,N_5253);
nor U5376 (N_5376,N_5281,N_5306);
and U5377 (N_5377,N_5256,N_5353);
nor U5378 (N_5378,N_5329,N_5273);
nor U5379 (N_5379,N_5322,N_5305);
or U5380 (N_5380,N_5252,N_5356);
nand U5381 (N_5381,N_5259,N_5286);
nor U5382 (N_5382,N_5254,N_5374);
and U5383 (N_5383,N_5317,N_5360);
nor U5384 (N_5384,N_5303,N_5316);
xnor U5385 (N_5385,N_5347,N_5278);
and U5386 (N_5386,N_5355,N_5351);
nand U5387 (N_5387,N_5296,N_5361);
or U5388 (N_5388,N_5269,N_5308);
or U5389 (N_5389,N_5369,N_5321);
or U5390 (N_5390,N_5338,N_5366);
and U5391 (N_5391,N_5345,N_5287);
nand U5392 (N_5392,N_5282,N_5370);
nor U5393 (N_5393,N_5260,N_5330);
nand U5394 (N_5394,N_5276,N_5365);
or U5395 (N_5395,N_5320,N_5346);
xor U5396 (N_5396,N_5325,N_5279);
nand U5397 (N_5397,N_5271,N_5290);
nor U5398 (N_5398,N_5364,N_5314);
xor U5399 (N_5399,N_5334,N_5265);
or U5400 (N_5400,N_5342,N_5367);
nand U5401 (N_5401,N_5285,N_5284);
and U5402 (N_5402,N_5310,N_5298);
nor U5403 (N_5403,N_5272,N_5293);
xnor U5404 (N_5404,N_5267,N_5300);
or U5405 (N_5405,N_5262,N_5280);
nand U5406 (N_5406,N_5333,N_5363);
or U5407 (N_5407,N_5266,N_5350);
nand U5408 (N_5408,N_5258,N_5302);
and U5409 (N_5409,N_5327,N_5344);
or U5410 (N_5410,N_5337,N_5250);
nand U5411 (N_5411,N_5307,N_5312);
xnor U5412 (N_5412,N_5348,N_5340);
nor U5413 (N_5413,N_5328,N_5357);
or U5414 (N_5414,N_5368,N_5319);
xnor U5415 (N_5415,N_5263,N_5371);
and U5416 (N_5416,N_5294,N_5315);
or U5417 (N_5417,N_5324,N_5277);
and U5418 (N_5418,N_5251,N_5349);
nand U5419 (N_5419,N_5318,N_5343);
nor U5420 (N_5420,N_5288,N_5275);
nor U5421 (N_5421,N_5274,N_5326);
xnor U5422 (N_5422,N_5257,N_5309);
and U5423 (N_5423,N_5291,N_5311);
nand U5424 (N_5424,N_5373,N_5332);
xor U5425 (N_5425,N_5336,N_5339);
nor U5426 (N_5426,N_5358,N_5261);
xor U5427 (N_5427,N_5289,N_5341);
nor U5428 (N_5428,N_5301,N_5372);
or U5429 (N_5429,N_5268,N_5304);
nand U5430 (N_5430,N_5359,N_5295);
and U5431 (N_5431,N_5331,N_5283);
or U5432 (N_5432,N_5297,N_5354);
nor U5433 (N_5433,N_5335,N_5299);
xor U5434 (N_5434,N_5352,N_5255);
and U5435 (N_5435,N_5264,N_5292);
nor U5436 (N_5436,N_5313,N_5323);
and U5437 (N_5437,N_5270,N_5263);
nand U5438 (N_5438,N_5345,N_5299);
nor U5439 (N_5439,N_5298,N_5288);
nor U5440 (N_5440,N_5308,N_5278);
and U5441 (N_5441,N_5267,N_5302);
nor U5442 (N_5442,N_5266,N_5300);
or U5443 (N_5443,N_5293,N_5342);
or U5444 (N_5444,N_5369,N_5270);
or U5445 (N_5445,N_5312,N_5302);
nand U5446 (N_5446,N_5254,N_5371);
nand U5447 (N_5447,N_5282,N_5348);
xor U5448 (N_5448,N_5354,N_5348);
nand U5449 (N_5449,N_5308,N_5270);
nor U5450 (N_5450,N_5266,N_5326);
or U5451 (N_5451,N_5280,N_5317);
xnor U5452 (N_5452,N_5287,N_5303);
xnor U5453 (N_5453,N_5314,N_5276);
and U5454 (N_5454,N_5343,N_5267);
or U5455 (N_5455,N_5314,N_5327);
nor U5456 (N_5456,N_5305,N_5297);
or U5457 (N_5457,N_5364,N_5297);
and U5458 (N_5458,N_5307,N_5267);
nand U5459 (N_5459,N_5325,N_5374);
xnor U5460 (N_5460,N_5348,N_5299);
and U5461 (N_5461,N_5259,N_5308);
nor U5462 (N_5462,N_5309,N_5255);
nand U5463 (N_5463,N_5299,N_5369);
or U5464 (N_5464,N_5347,N_5285);
nand U5465 (N_5465,N_5295,N_5265);
and U5466 (N_5466,N_5321,N_5279);
or U5467 (N_5467,N_5324,N_5323);
xnor U5468 (N_5468,N_5373,N_5316);
xor U5469 (N_5469,N_5251,N_5363);
nor U5470 (N_5470,N_5276,N_5329);
nor U5471 (N_5471,N_5323,N_5337);
and U5472 (N_5472,N_5270,N_5315);
nor U5473 (N_5473,N_5352,N_5313);
and U5474 (N_5474,N_5275,N_5356);
nand U5475 (N_5475,N_5282,N_5273);
or U5476 (N_5476,N_5284,N_5350);
nand U5477 (N_5477,N_5304,N_5331);
or U5478 (N_5478,N_5276,N_5255);
and U5479 (N_5479,N_5346,N_5267);
nand U5480 (N_5480,N_5284,N_5362);
nor U5481 (N_5481,N_5295,N_5348);
nand U5482 (N_5482,N_5314,N_5325);
nand U5483 (N_5483,N_5341,N_5263);
nand U5484 (N_5484,N_5255,N_5366);
and U5485 (N_5485,N_5359,N_5260);
or U5486 (N_5486,N_5295,N_5272);
nand U5487 (N_5487,N_5259,N_5288);
or U5488 (N_5488,N_5367,N_5346);
and U5489 (N_5489,N_5331,N_5368);
nand U5490 (N_5490,N_5363,N_5254);
or U5491 (N_5491,N_5303,N_5355);
xnor U5492 (N_5492,N_5358,N_5267);
and U5493 (N_5493,N_5362,N_5341);
xor U5494 (N_5494,N_5347,N_5252);
nor U5495 (N_5495,N_5324,N_5314);
and U5496 (N_5496,N_5352,N_5296);
and U5497 (N_5497,N_5276,N_5309);
xnor U5498 (N_5498,N_5291,N_5288);
xor U5499 (N_5499,N_5284,N_5328);
and U5500 (N_5500,N_5392,N_5429);
nand U5501 (N_5501,N_5498,N_5432);
nand U5502 (N_5502,N_5404,N_5474);
nor U5503 (N_5503,N_5430,N_5449);
and U5504 (N_5504,N_5494,N_5391);
xnor U5505 (N_5505,N_5478,N_5459);
and U5506 (N_5506,N_5415,N_5460);
xor U5507 (N_5507,N_5428,N_5470);
or U5508 (N_5508,N_5379,N_5469);
nor U5509 (N_5509,N_5390,N_5466);
nand U5510 (N_5510,N_5385,N_5465);
nor U5511 (N_5511,N_5485,N_5377);
or U5512 (N_5512,N_5422,N_5407);
or U5513 (N_5513,N_5477,N_5398);
and U5514 (N_5514,N_5473,N_5386);
xor U5515 (N_5515,N_5421,N_5417);
xnor U5516 (N_5516,N_5495,N_5457);
xor U5517 (N_5517,N_5409,N_5427);
and U5518 (N_5518,N_5475,N_5437);
or U5519 (N_5519,N_5463,N_5426);
xor U5520 (N_5520,N_5451,N_5378);
and U5521 (N_5521,N_5440,N_5425);
nand U5522 (N_5522,N_5448,N_5414);
nor U5523 (N_5523,N_5394,N_5453);
or U5524 (N_5524,N_5413,N_5497);
and U5525 (N_5525,N_5435,N_5444);
or U5526 (N_5526,N_5450,N_5441);
or U5527 (N_5527,N_5499,N_5420);
or U5528 (N_5528,N_5484,N_5431);
and U5529 (N_5529,N_5403,N_5452);
and U5530 (N_5530,N_5480,N_5424);
nand U5531 (N_5531,N_5380,N_5493);
nor U5532 (N_5532,N_5464,N_5399);
nand U5533 (N_5533,N_5445,N_5433);
nor U5534 (N_5534,N_5387,N_5412);
and U5535 (N_5535,N_5384,N_5481);
and U5536 (N_5536,N_5401,N_5406);
nor U5537 (N_5537,N_5471,N_5447);
or U5538 (N_5538,N_5397,N_5393);
xnor U5539 (N_5539,N_5439,N_5454);
xor U5540 (N_5540,N_5383,N_5461);
nand U5541 (N_5541,N_5434,N_5381);
nand U5542 (N_5542,N_5456,N_5436);
nand U5543 (N_5543,N_5476,N_5455);
nand U5544 (N_5544,N_5458,N_5405);
xnor U5545 (N_5545,N_5443,N_5376);
nand U5546 (N_5546,N_5446,N_5408);
and U5547 (N_5547,N_5411,N_5418);
nor U5548 (N_5548,N_5483,N_5487);
xnor U5549 (N_5549,N_5438,N_5419);
xor U5550 (N_5550,N_5402,N_5488);
nor U5551 (N_5551,N_5496,N_5389);
xor U5552 (N_5552,N_5375,N_5472);
or U5553 (N_5553,N_5423,N_5482);
or U5554 (N_5554,N_5396,N_5491);
nand U5555 (N_5555,N_5395,N_5486);
xnor U5556 (N_5556,N_5489,N_5400);
nand U5557 (N_5557,N_5442,N_5382);
nand U5558 (N_5558,N_5410,N_5388);
nand U5559 (N_5559,N_5490,N_5467);
nor U5560 (N_5560,N_5416,N_5479);
or U5561 (N_5561,N_5462,N_5468);
or U5562 (N_5562,N_5492,N_5393);
or U5563 (N_5563,N_5394,N_5378);
xnor U5564 (N_5564,N_5479,N_5462);
nand U5565 (N_5565,N_5410,N_5436);
or U5566 (N_5566,N_5406,N_5431);
nor U5567 (N_5567,N_5435,N_5498);
nor U5568 (N_5568,N_5470,N_5499);
xnor U5569 (N_5569,N_5402,N_5464);
or U5570 (N_5570,N_5482,N_5430);
nand U5571 (N_5571,N_5487,N_5465);
nand U5572 (N_5572,N_5476,N_5410);
nand U5573 (N_5573,N_5425,N_5478);
or U5574 (N_5574,N_5496,N_5479);
and U5575 (N_5575,N_5434,N_5484);
xor U5576 (N_5576,N_5439,N_5478);
nand U5577 (N_5577,N_5396,N_5466);
and U5578 (N_5578,N_5480,N_5472);
or U5579 (N_5579,N_5464,N_5460);
xnor U5580 (N_5580,N_5399,N_5488);
nor U5581 (N_5581,N_5382,N_5445);
xor U5582 (N_5582,N_5440,N_5436);
xnor U5583 (N_5583,N_5426,N_5410);
nor U5584 (N_5584,N_5488,N_5497);
or U5585 (N_5585,N_5456,N_5465);
nand U5586 (N_5586,N_5439,N_5480);
xor U5587 (N_5587,N_5468,N_5486);
nand U5588 (N_5588,N_5480,N_5448);
nand U5589 (N_5589,N_5483,N_5441);
or U5590 (N_5590,N_5445,N_5489);
and U5591 (N_5591,N_5432,N_5409);
nand U5592 (N_5592,N_5416,N_5455);
nor U5593 (N_5593,N_5376,N_5426);
or U5594 (N_5594,N_5443,N_5493);
and U5595 (N_5595,N_5470,N_5491);
xor U5596 (N_5596,N_5440,N_5470);
and U5597 (N_5597,N_5380,N_5448);
nand U5598 (N_5598,N_5410,N_5478);
nand U5599 (N_5599,N_5427,N_5415);
nand U5600 (N_5600,N_5387,N_5493);
nor U5601 (N_5601,N_5406,N_5429);
or U5602 (N_5602,N_5483,N_5472);
nand U5603 (N_5603,N_5494,N_5438);
or U5604 (N_5604,N_5470,N_5490);
nor U5605 (N_5605,N_5432,N_5451);
nand U5606 (N_5606,N_5461,N_5455);
and U5607 (N_5607,N_5415,N_5375);
nor U5608 (N_5608,N_5439,N_5421);
nand U5609 (N_5609,N_5499,N_5425);
nor U5610 (N_5610,N_5424,N_5405);
nand U5611 (N_5611,N_5375,N_5377);
xor U5612 (N_5612,N_5458,N_5423);
nor U5613 (N_5613,N_5395,N_5400);
or U5614 (N_5614,N_5433,N_5409);
and U5615 (N_5615,N_5466,N_5428);
xnor U5616 (N_5616,N_5396,N_5498);
or U5617 (N_5617,N_5442,N_5475);
nand U5618 (N_5618,N_5415,N_5468);
or U5619 (N_5619,N_5441,N_5409);
or U5620 (N_5620,N_5463,N_5393);
nor U5621 (N_5621,N_5398,N_5447);
nor U5622 (N_5622,N_5390,N_5379);
and U5623 (N_5623,N_5397,N_5413);
nand U5624 (N_5624,N_5452,N_5498);
nand U5625 (N_5625,N_5576,N_5554);
xor U5626 (N_5626,N_5609,N_5569);
or U5627 (N_5627,N_5589,N_5595);
xor U5628 (N_5628,N_5590,N_5622);
nand U5629 (N_5629,N_5521,N_5535);
or U5630 (N_5630,N_5547,N_5603);
xnor U5631 (N_5631,N_5610,N_5566);
or U5632 (N_5632,N_5567,N_5596);
xnor U5633 (N_5633,N_5504,N_5579);
nand U5634 (N_5634,N_5527,N_5509);
and U5635 (N_5635,N_5523,N_5586);
and U5636 (N_5636,N_5502,N_5507);
xnor U5637 (N_5637,N_5594,N_5544);
nor U5638 (N_5638,N_5575,N_5584);
nor U5639 (N_5639,N_5537,N_5549);
and U5640 (N_5640,N_5602,N_5570);
xor U5641 (N_5641,N_5506,N_5536);
nor U5642 (N_5642,N_5597,N_5518);
xor U5643 (N_5643,N_5592,N_5587);
or U5644 (N_5644,N_5534,N_5553);
xnor U5645 (N_5645,N_5560,N_5582);
and U5646 (N_5646,N_5613,N_5501);
nor U5647 (N_5647,N_5545,N_5503);
or U5648 (N_5648,N_5533,N_5561);
nor U5649 (N_5649,N_5600,N_5565);
nand U5650 (N_5650,N_5624,N_5524);
or U5651 (N_5651,N_5606,N_5525);
nor U5652 (N_5652,N_5529,N_5580);
nor U5653 (N_5653,N_5559,N_5530);
xnor U5654 (N_5654,N_5614,N_5607);
or U5655 (N_5655,N_5519,N_5574);
nand U5656 (N_5656,N_5577,N_5608);
nor U5657 (N_5657,N_5532,N_5623);
xor U5658 (N_5658,N_5621,N_5555);
xor U5659 (N_5659,N_5585,N_5604);
or U5660 (N_5660,N_5612,N_5540);
nand U5661 (N_5661,N_5505,N_5556);
xnor U5662 (N_5662,N_5573,N_5511);
nand U5663 (N_5663,N_5557,N_5611);
or U5664 (N_5664,N_5513,N_5562);
and U5665 (N_5665,N_5520,N_5543);
and U5666 (N_5666,N_5617,N_5571);
xnor U5667 (N_5667,N_5548,N_5620);
and U5668 (N_5668,N_5542,N_5526);
and U5669 (N_5669,N_5572,N_5528);
or U5670 (N_5670,N_5615,N_5558);
or U5671 (N_5671,N_5551,N_5616);
and U5672 (N_5672,N_5546,N_5581);
and U5673 (N_5673,N_5563,N_5552);
xnor U5674 (N_5674,N_5593,N_5598);
nor U5675 (N_5675,N_5591,N_5564);
nand U5676 (N_5676,N_5601,N_5531);
nor U5677 (N_5677,N_5619,N_5541);
nand U5678 (N_5678,N_5550,N_5516);
nand U5679 (N_5679,N_5514,N_5588);
nor U5680 (N_5680,N_5512,N_5508);
nor U5681 (N_5681,N_5515,N_5522);
nand U5682 (N_5682,N_5510,N_5618);
xnor U5683 (N_5683,N_5500,N_5583);
nand U5684 (N_5684,N_5605,N_5539);
xnor U5685 (N_5685,N_5578,N_5538);
or U5686 (N_5686,N_5568,N_5517);
or U5687 (N_5687,N_5599,N_5516);
or U5688 (N_5688,N_5526,N_5559);
or U5689 (N_5689,N_5608,N_5530);
and U5690 (N_5690,N_5505,N_5569);
nor U5691 (N_5691,N_5541,N_5620);
nor U5692 (N_5692,N_5509,N_5530);
xnor U5693 (N_5693,N_5584,N_5580);
nand U5694 (N_5694,N_5586,N_5508);
nor U5695 (N_5695,N_5615,N_5503);
xnor U5696 (N_5696,N_5548,N_5517);
nand U5697 (N_5697,N_5559,N_5542);
nand U5698 (N_5698,N_5593,N_5590);
or U5699 (N_5699,N_5575,N_5501);
nand U5700 (N_5700,N_5558,N_5590);
and U5701 (N_5701,N_5554,N_5525);
or U5702 (N_5702,N_5529,N_5597);
nand U5703 (N_5703,N_5570,N_5516);
xor U5704 (N_5704,N_5516,N_5533);
or U5705 (N_5705,N_5590,N_5591);
and U5706 (N_5706,N_5566,N_5617);
or U5707 (N_5707,N_5596,N_5548);
xnor U5708 (N_5708,N_5526,N_5520);
xnor U5709 (N_5709,N_5582,N_5589);
nand U5710 (N_5710,N_5621,N_5508);
nor U5711 (N_5711,N_5515,N_5621);
xor U5712 (N_5712,N_5562,N_5567);
and U5713 (N_5713,N_5552,N_5528);
nor U5714 (N_5714,N_5541,N_5506);
and U5715 (N_5715,N_5555,N_5617);
xnor U5716 (N_5716,N_5579,N_5516);
nor U5717 (N_5717,N_5505,N_5587);
nand U5718 (N_5718,N_5621,N_5550);
nand U5719 (N_5719,N_5619,N_5568);
and U5720 (N_5720,N_5607,N_5612);
and U5721 (N_5721,N_5611,N_5563);
xnor U5722 (N_5722,N_5604,N_5622);
xor U5723 (N_5723,N_5570,N_5522);
and U5724 (N_5724,N_5523,N_5581);
xnor U5725 (N_5725,N_5515,N_5543);
xnor U5726 (N_5726,N_5608,N_5612);
or U5727 (N_5727,N_5533,N_5624);
or U5728 (N_5728,N_5561,N_5615);
or U5729 (N_5729,N_5520,N_5585);
nor U5730 (N_5730,N_5587,N_5606);
nor U5731 (N_5731,N_5524,N_5597);
xor U5732 (N_5732,N_5622,N_5517);
nand U5733 (N_5733,N_5607,N_5583);
and U5734 (N_5734,N_5585,N_5578);
xnor U5735 (N_5735,N_5546,N_5612);
xor U5736 (N_5736,N_5570,N_5559);
nor U5737 (N_5737,N_5577,N_5522);
nand U5738 (N_5738,N_5621,N_5619);
or U5739 (N_5739,N_5549,N_5622);
xor U5740 (N_5740,N_5507,N_5520);
and U5741 (N_5741,N_5514,N_5590);
nand U5742 (N_5742,N_5605,N_5553);
nand U5743 (N_5743,N_5621,N_5584);
xor U5744 (N_5744,N_5598,N_5604);
xnor U5745 (N_5745,N_5603,N_5612);
nor U5746 (N_5746,N_5537,N_5607);
nor U5747 (N_5747,N_5593,N_5558);
or U5748 (N_5748,N_5528,N_5542);
nand U5749 (N_5749,N_5607,N_5603);
and U5750 (N_5750,N_5657,N_5743);
nand U5751 (N_5751,N_5651,N_5732);
nor U5752 (N_5752,N_5737,N_5638);
nand U5753 (N_5753,N_5728,N_5626);
xor U5754 (N_5754,N_5692,N_5719);
and U5755 (N_5755,N_5643,N_5693);
nor U5756 (N_5756,N_5704,N_5709);
nand U5757 (N_5757,N_5746,N_5644);
nor U5758 (N_5758,N_5749,N_5652);
nand U5759 (N_5759,N_5676,N_5669);
xor U5760 (N_5760,N_5641,N_5739);
or U5761 (N_5761,N_5744,N_5702);
and U5762 (N_5762,N_5637,N_5722);
xor U5763 (N_5763,N_5631,N_5649);
and U5764 (N_5764,N_5664,N_5672);
nor U5765 (N_5765,N_5736,N_5661);
nand U5766 (N_5766,N_5642,N_5650);
and U5767 (N_5767,N_5742,N_5691);
nor U5768 (N_5768,N_5721,N_5738);
nor U5769 (N_5769,N_5665,N_5681);
nor U5770 (N_5770,N_5690,N_5636);
nand U5771 (N_5771,N_5682,N_5674);
nor U5772 (N_5772,N_5727,N_5632);
nor U5773 (N_5773,N_5679,N_5668);
and U5774 (N_5774,N_5680,N_5716);
xor U5775 (N_5775,N_5627,N_5720);
nor U5776 (N_5776,N_5697,N_5726);
nand U5777 (N_5777,N_5698,N_5629);
or U5778 (N_5778,N_5683,N_5640);
or U5779 (N_5779,N_5653,N_5717);
nand U5780 (N_5780,N_5677,N_5670);
xor U5781 (N_5781,N_5699,N_5725);
xnor U5782 (N_5782,N_5662,N_5666);
xor U5783 (N_5783,N_5731,N_5645);
xor U5784 (N_5784,N_5705,N_5635);
and U5785 (N_5785,N_5686,N_5694);
nor U5786 (N_5786,N_5688,N_5639);
and U5787 (N_5787,N_5735,N_5748);
xnor U5788 (N_5788,N_5701,N_5625);
nand U5789 (N_5789,N_5655,N_5660);
xor U5790 (N_5790,N_5700,N_5745);
nor U5791 (N_5791,N_5648,N_5715);
xor U5792 (N_5792,N_5634,N_5707);
or U5793 (N_5793,N_5673,N_5647);
nand U5794 (N_5794,N_5740,N_5718);
nand U5795 (N_5795,N_5628,N_5724);
and U5796 (N_5796,N_5671,N_5741);
nor U5797 (N_5797,N_5714,N_5656);
nand U5798 (N_5798,N_5684,N_5729);
nor U5799 (N_5799,N_5712,N_5723);
or U5800 (N_5800,N_5689,N_5658);
or U5801 (N_5801,N_5659,N_5654);
xnor U5802 (N_5802,N_5667,N_5711);
nand U5803 (N_5803,N_5633,N_5675);
and U5804 (N_5804,N_5685,N_5695);
xnor U5805 (N_5805,N_5630,N_5734);
nand U5806 (N_5806,N_5678,N_5733);
nor U5807 (N_5807,N_5696,N_5710);
or U5808 (N_5808,N_5687,N_5747);
nand U5809 (N_5809,N_5703,N_5730);
or U5810 (N_5810,N_5646,N_5708);
or U5811 (N_5811,N_5706,N_5713);
nand U5812 (N_5812,N_5663,N_5637);
or U5813 (N_5813,N_5704,N_5636);
or U5814 (N_5814,N_5738,N_5662);
nor U5815 (N_5815,N_5667,N_5681);
xnor U5816 (N_5816,N_5676,N_5650);
nand U5817 (N_5817,N_5642,N_5730);
xnor U5818 (N_5818,N_5742,N_5661);
nand U5819 (N_5819,N_5658,N_5744);
nand U5820 (N_5820,N_5662,N_5743);
nor U5821 (N_5821,N_5748,N_5683);
and U5822 (N_5822,N_5710,N_5731);
or U5823 (N_5823,N_5656,N_5638);
or U5824 (N_5824,N_5682,N_5692);
nor U5825 (N_5825,N_5666,N_5711);
and U5826 (N_5826,N_5679,N_5749);
or U5827 (N_5827,N_5737,N_5643);
nor U5828 (N_5828,N_5632,N_5718);
nor U5829 (N_5829,N_5630,N_5719);
xor U5830 (N_5830,N_5708,N_5715);
nand U5831 (N_5831,N_5715,N_5703);
nand U5832 (N_5832,N_5645,N_5686);
and U5833 (N_5833,N_5690,N_5660);
xor U5834 (N_5834,N_5675,N_5718);
nor U5835 (N_5835,N_5707,N_5731);
or U5836 (N_5836,N_5686,N_5637);
or U5837 (N_5837,N_5726,N_5641);
xnor U5838 (N_5838,N_5711,N_5655);
or U5839 (N_5839,N_5679,N_5637);
nand U5840 (N_5840,N_5711,N_5739);
nor U5841 (N_5841,N_5720,N_5704);
nor U5842 (N_5842,N_5638,N_5710);
xnor U5843 (N_5843,N_5645,N_5648);
nor U5844 (N_5844,N_5643,N_5655);
nor U5845 (N_5845,N_5630,N_5640);
and U5846 (N_5846,N_5667,N_5725);
and U5847 (N_5847,N_5726,N_5749);
or U5848 (N_5848,N_5629,N_5695);
xnor U5849 (N_5849,N_5642,N_5664);
or U5850 (N_5850,N_5681,N_5713);
xor U5851 (N_5851,N_5723,N_5707);
or U5852 (N_5852,N_5675,N_5724);
or U5853 (N_5853,N_5693,N_5723);
or U5854 (N_5854,N_5645,N_5745);
or U5855 (N_5855,N_5635,N_5743);
nor U5856 (N_5856,N_5735,N_5649);
nand U5857 (N_5857,N_5660,N_5656);
nor U5858 (N_5858,N_5656,N_5626);
nand U5859 (N_5859,N_5712,N_5667);
nand U5860 (N_5860,N_5684,N_5634);
nor U5861 (N_5861,N_5660,N_5731);
nand U5862 (N_5862,N_5723,N_5718);
nor U5863 (N_5863,N_5738,N_5650);
and U5864 (N_5864,N_5711,N_5737);
nor U5865 (N_5865,N_5727,N_5635);
or U5866 (N_5866,N_5659,N_5666);
or U5867 (N_5867,N_5662,N_5726);
nor U5868 (N_5868,N_5667,N_5648);
nand U5869 (N_5869,N_5635,N_5715);
nand U5870 (N_5870,N_5695,N_5625);
xnor U5871 (N_5871,N_5725,N_5708);
nor U5872 (N_5872,N_5650,N_5655);
xor U5873 (N_5873,N_5732,N_5635);
nor U5874 (N_5874,N_5723,N_5678);
xor U5875 (N_5875,N_5834,N_5819);
nand U5876 (N_5876,N_5817,N_5867);
or U5877 (N_5877,N_5859,N_5770);
nand U5878 (N_5878,N_5837,N_5756);
xnor U5879 (N_5879,N_5855,N_5755);
xnor U5880 (N_5880,N_5754,N_5814);
or U5881 (N_5881,N_5772,N_5843);
or U5882 (N_5882,N_5750,N_5802);
nand U5883 (N_5883,N_5849,N_5799);
and U5884 (N_5884,N_5767,N_5761);
or U5885 (N_5885,N_5823,N_5848);
nor U5886 (N_5886,N_5791,N_5800);
nor U5887 (N_5887,N_5769,N_5759);
and U5888 (N_5888,N_5826,N_5760);
nor U5889 (N_5889,N_5807,N_5863);
nor U5890 (N_5890,N_5777,N_5874);
or U5891 (N_5891,N_5792,N_5758);
and U5892 (N_5892,N_5808,N_5872);
and U5893 (N_5893,N_5763,N_5816);
xnor U5894 (N_5894,N_5827,N_5873);
and U5895 (N_5895,N_5846,N_5821);
or U5896 (N_5896,N_5845,N_5786);
xor U5897 (N_5897,N_5774,N_5779);
xnor U5898 (N_5898,N_5778,N_5787);
nand U5899 (N_5899,N_5809,N_5868);
and U5900 (N_5900,N_5751,N_5815);
or U5901 (N_5901,N_5833,N_5762);
or U5902 (N_5902,N_5806,N_5781);
and U5903 (N_5903,N_5862,N_5798);
xnor U5904 (N_5904,N_5822,N_5836);
nor U5905 (N_5905,N_5857,N_5832);
nor U5906 (N_5906,N_5856,N_5794);
nor U5907 (N_5907,N_5776,N_5818);
and U5908 (N_5908,N_5847,N_5785);
and U5909 (N_5909,N_5851,N_5801);
nor U5910 (N_5910,N_5852,N_5813);
xor U5911 (N_5911,N_5773,N_5829);
nand U5912 (N_5912,N_5805,N_5789);
nand U5913 (N_5913,N_5842,N_5784);
or U5914 (N_5914,N_5830,N_5804);
and U5915 (N_5915,N_5752,N_5757);
and U5916 (N_5916,N_5782,N_5771);
or U5917 (N_5917,N_5870,N_5871);
and U5918 (N_5918,N_5839,N_5831);
or U5919 (N_5919,N_5793,N_5768);
nand U5920 (N_5920,N_5765,N_5753);
nand U5921 (N_5921,N_5780,N_5869);
nor U5922 (N_5922,N_5812,N_5795);
nor U5923 (N_5923,N_5865,N_5797);
nand U5924 (N_5924,N_5854,N_5790);
nand U5925 (N_5925,N_5835,N_5764);
and U5926 (N_5926,N_5824,N_5864);
or U5927 (N_5927,N_5866,N_5811);
xor U5928 (N_5928,N_5861,N_5828);
and U5929 (N_5929,N_5803,N_5841);
xnor U5930 (N_5930,N_5820,N_5840);
xor U5931 (N_5931,N_5860,N_5796);
or U5932 (N_5932,N_5838,N_5825);
nor U5933 (N_5933,N_5775,N_5853);
and U5934 (N_5934,N_5858,N_5850);
nor U5935 (N_5935,N_5783,N_5788);
nand U5936 (N_5936,N_5810,N_5844);
nand U5937 (N_5937,N_5766,N_5838);
nor U5938 (N_5938,N_5795,N_5767);
nor U5939 (N_5939,N_5826,N_5811);
nand U5940 (N_5940,N_5860,N_5869);
nor U5941 (N_5941,N_5856,N_5783);
nor U5942 (N_5942,N_5850,N_5851);
nand U5943 (N_5943,N_5758,N_5861);
or U5944 (N_5944,N_5803,N_5754);
nor U5945 (N_5945,N_5750,N_5790);
xor U5946 (N_5946,N_5755,N_5869);
xnor U5947 (N_5947,N_5786,N_5833);
or U5948 (N_5948,N_5859,N_5847);
or U5949 (N_5949,N_5867,N_5804);
and U5950 (N_5950,N_5830,N_5841);
xor U5951 (N_5951,N_5823,N_5764);
and U5952 (N_5952,N_5832,N_5751);
and U5953 (N_5953,N_5867,N_5779);
and U5954 (N_5954,N_5763,N_5784);
xnor U5955 (N_5955,N_5755,N_5826);
or U5956 (N_5956,N_5824,N_5831);
xnor U5957 (N_5957,N_5800,N_5789);
or U5958 (N_5958,N_5867,N_5826);
or U5959 (N_5959,N_5774,N_5777);
or U5960 (N_5960,N_5805,N_5847);
xor U5961 (N_5961,N_5869,N_5754);
or U5962 (N_5962,N_5822,N_5847);
xor U5963 (N_5963,N_5854,N_5832);
xor U5964 (N_5964,N_5844,N_5860);
or U5965 (N_5965,N_5860,N_5764);
nor U5966 (N_5966,N_5868,N_5817);
xnor U5967 (N_5967,N_5865,N_5850);
xnor U5968 (N_5968,N_5801,N_5792);
nor U5969 (N_5969,N_5869,N_5858);
nor U5970 (N_5970,N_5768,N_5757);
nand U5971 (N_5971,N_5760,N_5847);
nand U5972 (N_5972,N_5766,N_5848);
or U5973 (N_5973,N_5851,N_5848);
nand U5974 (N_5974,N_5807,N_5849);
and U5975 (N_5975,N_5754,N_5865);
xnor U5976 (N_5976,N_5861,N_5809);
or U5977 (N_5977,N_5752,N_5814);
xnor U5978 (N_5978,N_5851,N_5784);
nand U5979 (N_5979,N_5785,N_5798);
nor U5980 (N_5980,N_5771,N_5777);
and U5981 (N_5981,N_5837,N_5765);
and U5982 (N_5982,N_5787,N_5767);
and U5983 (N_5983,N_5874,N_5757);
or U5984 (N_5984,N_5754,N_5751);
or U5985 (N_5985,N_5804,N_5860);
and U5986 (N_5986,N_5757,N_5787);
nor U5987 (N_5987,N_5849,N_5822);
and U5988 (N_5988,N_5867,N_5873);
or U5989 (N_5989,N_5830,N_5835);
xor U5990 (N_5990,N_5767,N_5840);
and U5991 (N_5991,N_5850,N_5867);
nand U5992 (N_5992,N_5790,N_5800);
or U5993 (N_5993,N_5796,N_5851);
xor U5994 (N_5994,N_5792,N_5769);
xnor U5995 (N_5995,N_5756,N_5868);
xor U5996 (N_5996,N_5793,N_5847);
or U5997 (N_5997,N_5778,N_5811);
nor U5998 (N_5998,N_5833,N_5858);
nand U5999 (N_5999,N_5794,N_5849);
xnor U6000 (N_6000,N_5909,N_5875);
xnor U6001 (N_6001,N_5915,N_5951);
xnor U6002 (N_6002,N_5898,N_5941);
nor U6003 (N_6003,N_5964,N_5999);
or U6004 (N_6004,N_5905,N_5912);
nand U6005 (N_6005,N_5992,N_5975);
nand U6006 (N_6006,N_5973,N_5903);
xnor U6007 (N_6007,N_5893,N_5966);
and U6008 (N_6008,N_5879,N_5894);
xor U6009 (N_6009,N_5980,N_5919);
or U6010 (N_6010,N_5946,N_5886);
and U6011 (N_6011,N_5906,N_5901);
and U6012 (N_6012,N_5931,N_5904);
nand U6013 (N_6013,N_5953,N_5985);
nand U6014 (N_6014,N_5892,N_5920);
nor U6015 (N_6015,N_5889,N_5922);
nand U6016 (N_6016,N_5917,N_5902);
nand U6017 (N_6017,N_5952,N_5998);
nor U6018 (N_6018,N_5995,N_5895);
nand U6019 (N_6019,N_5994,N_5927);
and U6020 (N_6020,N_5974,N_5921);
nand U6021 (N_6021,N_5885,N_5929);
or U6022 (N_6022,N_5996,N_5949);
xor U6023 (N_6023,N_5988,N_5958);
or U6024 (N_6024,N_5950,N_5944);
or U6025 (N_6025,N_5930,N_5925);
and U6026 (N_6026,N_5897,N_5926);
nand U6027 (N_6027,N_5971,N_5884);
nor U6028 (N_6028,N_5936,N_5991);
and U6029 (N_6029,N_5888,N_5924);
or U6030 (N_6030,N_5918,N_5932);
or U6031 (N_6031,N_5965,N_5987);
xor U6032 (N_6032,N_5981,N_5989);
nor U6033 (N_6033,N_5969,N_5977);
nand U6034 (N_6034,N_5900,N_5957);
nor U6035 (N_6035,N_5896,N_5940);
and U6036 (N_6036,N_5890,N_5947);
and U6037 (N_6037,N_5887,N_5908);
xor U6038 (N_6038,N_5880,N_5955);
xor U6039 (N_6039,N_5914,N_5937);
and U6040 (N_6040,N_5962,N_5881);
or U6041 (N_6041,N_5997,N_5934);
nand U6042 (N_6042,N_5876,N_5935);
or U6043 (N_6043,N_5986,N_5978);
or U6044 (N_6044,N_5993,N_5972);
nand U6045 (N_6045,N_5933,N_5911);
and U6046 (N_6046,N_5899,N_5943);
xnor U6047 (N_6047,N_5913,N_5976);
nor U6048 (N_6048,N_5948,N_5877);
xnor U6049 (N_6049,N_5938,N_5959);
and U6050 (N_6050,N_5970,N_5963);
xnor U6051 (N_6051,N_5979,N_5983);
and U6052 (N_6052,N_5878,N_5910);
or U6053 (N_6053,N_5928,N_5968);
and U6054 (N_6054,N_5990,N_5923);
xnor U6055 (N_6055,N_5939,N_5891);
nor U6056 (N_6056,N_5954,N_5907);
nand U6057 (N_6057,N_5956,N_5961);
and U6058 (N_6058,N_5984,N_5945);
nand U6059 (N_6059,N_5883,N_5967);
or U6060 (N_6060,N_5942,N_5916);
nand U6061 (N_6061,N_5982,N_5882);
and U6062 (N_6062,N_5960,N_5904);
nor U6063 (N_6063,N_5990,N_5943);
or U6064 (N_6064,N_5974,N_5975);
and U6065 (N_6065,N_5991,N_5944);
and U6066 (N_6066,N_5938,N_5935);
nand U6067 (N_6067,N_5929,N_5911);
nand U6068 (N_6068,N_5902,N_5915);
and U6069 (N_6069,N_5999,N_5920);
xor U6070 (N_6070,N_5885,N_5880);
xor U6071 (N_6071,N_5976,N_5965);
nor U6072 (N_6072,N_5893,N_5991);
nand U6073 (N_6073,N_5909,N_5984);
or U6074 (N_6074,N_5973,N_5875);
or U6075 (N_6075,N_5996,N_5929);
nor U6076 (N_6076,N_5979,N_5927);
nor U6077 (N_6077,N_5907,N_5970);
xnor U6078 (N_6078,N_5920,N_5889);
xor U6079 (N_6079,N_5945,N_5908);
nor U6080 (N_6080,N_5943,N_5969);
xor U6081 (N_6081,N_5924,N_5955);
nor U6082 (N_6082,N_5897,N_5918);
nor U6083 (N_6083,N_5972,N_5901);
or U6084 (N_6084,N_5951,N_5977);
nand U6085 (N_6085,N_5982,N_5977);
xor U6086 (N_6086,N_5902,N_5942);
nor U6087 (N_6087,N_5916,N_5940);
nor U6088 (N_6088,N_5983,N_5927);
or U6089 (N_6089,N_5893,N_5904);
nor U6090 (N_6090,N_5887,N_5992);
nor U6091 (N_6091,N_5991,N_5880);
nand U6092 (N_6092,N_5920,N_5884);
and U6093 (N_6093,N_5969,N_5911);
nand U6094 (N_6094,N_5984,N_5905);
xnor U6095 (N_6095,N_5918,N_5885);
and U6096 (N_6096,N_5962,N_5915);
nand U6097 (N_6097,N_5949,N_5932);
nor U6098 (N_6098,N_5977,N_5989);
and U6099 (N_6099,N_5882,N_5911);
and U6100 (N_6100,N_5926,N_5960);
xor U6101 (N_6101,N_5962,N_5996);
nor U6102 (N_6102,N_5944,N_5982);
nor U6103 (N_6103,N_5997,N_5893);
nor U6104 (N_6104,N_5940,N_5978);
xor U6105 (N_6105,N_5961,N_5925);
nand U6106 (N_6106,N_5906,N_5993);
or U6107 (N_6107,N_5878,N_5903);
xor U6108 (N_6108,N_5947,N_5993);
and U6109 (N_6109,N_5929,N_5891);
nand U6110 (N_6110,N_5971,N_5881);
and U6111 (N_6111,N_5925,N_5934);
xnor U6112 (N_6112,N_5887,N_5932);
xor U6113 (N_6113,N_5978,N_5908);
nor U6114 (N_6114,N_5911,N_5997);
nand U6115 (N_6115,N_5891,N_5948);
xor U6116 (N_6116,N_5966,N_5934);
and U6117 (N_6117,N_5897,N_5888);
nand U6118 (N_6118,N_5899,N_5889);
nand U6119 (N_6119,N_5945,N_5897);
nor U6120 (N_6120,N_5943,N_5889);
xnor U6121 (N_6121,N_5940,N_5979);
nor U6122 (N_6122,N_5925,N_5926);
nor U6123 (N_6123,N_5895,N_5990);
or U6124 (N_6124,N_5946,N_5972);
or U6125 (N_6125,N_6020,N_6110);
nand U6126 (N_6126,N_6075,N_6023);
nor U6127 (N_6127,N_6119,N_6086);
nor U6128 (N_6128,N_6078,N_6089);
xnor U6129 (N_6129,N_6114,N_6076);
xor U6130 (N_6130,N_6059,N_6030);
nand U6131 (N_6131,N_6021,N_6025);
or U6132 (N_6132,N_6102,N_6108);
xor U6133 (N_6133,N_6055,N_6091);
nand U6134 (N_6134,N_6074,N_6037);
or U6135 (N_6135,N_6071,N_6095);
nor U6136 (N_6136,N_6022,N_6067);
nand U6137 (N_6137,N_6106,N_6070);
nor U6138 (N_6138,N_6079,N_6101);
nor U6139 (N_6139,N_6117,N_6027);
nor U6140 (N_6140,N_6016,N_6103);
or U6141 (N_6141,N_6082,N_6105);
nor U6142 (N_6142,N_6080,N_6015);
nor U6143 (N_6143,N_6061,N_6001);
or U6144 (N_6144,N_6120,N_6058);
or U6145 (N_6145,N_6111,N_6113);
xnor U6146 (N_6146,N_6083,N_6123);
xor U6147 (N_6147,N_6044,N_6104);
nand U6148 (N_6148,N_6039,N_6084);
or U6149 (N_6149,N_6097,N_6065);
and U6150 (N_6150,N_6118,N_6122);
and U6151 (N_6151,N_6046,N_6099);
or U6152 (N_6152,N_6034,N_6017);
nand U6153 (N_6153,N_6000,N_6073);
xnor U6154 (N_6154,N_6032,N_6047);
xor U6155 (N_6155,N_6042,N_6115);
nor U6156 (N_6156,N_6049,N_6033);
xor U6157 (N_6157,N_6031,N_6004);
xnor U6158 (N_6158,N_6038,N_6028);
and U6159 (N_6159,N_6092,N_6088);
and U6160 (N_6160,N_6087,N_6054);
nor U6161 (N_6161,N_6043,N_6002);
and U6162 (N_6162,N_6093,N_6006);
xnor U6163 (N_6163,N_6057,N_6012);
nor U6164 (N_6164,N_6041,N_6014);
and U6165 (N_6165,N_6085,N_6050);
xnor U6166 (N_6166,N_6040,N_6035);
nand U6167 (N_6167,N_6068,N_6107);
and U6168 (N_6168,N_6026,N_6124);
xnor U6169 (N_6169,N_6077,N_6008);
nor U6170 (N_6170,N_6060,N_6063);
or U6171 (N_6171,N_6090,N_6121);
and U6172 (N_6172,N_6066,N_6064);
xor U6173 (N_6173,N_6024,N_6112);
xnor U6174 (N_6174,N_6019,N_6056);
or U6175 (N_6175,N_6010,N_6013);
or U6176 (N_6176,N_6109,N_6048);
nand U6177 (N_6177,N_6005,N_6081);
or U6178 (N_6178,N_6003,N_6094);
nor U6179 (N_6179,N_6052,N_6098);
and U6180 (N_6180,N_6036,N_6045);
xor U6181 (N_6181,N_6009,N_6062);
nand U6182 (N_6182,N_6053,N_6051);
and U6183 (N_6183,N_6069,N_6100);
xnor U6184 (N_6184,N_6018,N_6007);
nand U6185 (N_6185,N_6072,N_6096);
or U6186 (N_6186,N_6011,N_6029);
nor U6187 (N_6187,N_6116,N_6109);
nand U6188 (N_6188,N_6034,N_6040);
nand U6189 (N_6189,N_6004,N_6069);
or U6190 (N_6190,N_6036,N_6101);
xnor U6191 (N_6191,N_6028,N_6073);
nor U6192 (N_6192,N_6097,N_6039);
nand U6193 (N_6193,N_6123,N_6097);
or U6194 (N_6194,N_6104,N_6071);
and U6195 (N_6195,N_6012,N_6017);
nor U6196 (N_6196,N_6007,N_6100);
and U6197 (N_6197,N_6119,N_6081);
xor U6198 (N_6198,N_6005,N_6092);
nand U6199 (N_6199,N_6092,N_6108);
xnor U6200 (N_6200,N_6069,N_6067);
and U6201 (N_6201,N_6075,N_6086);
xor U6202 (N_6202,N_6074,N_6034);
xor U6203 (N_6203,N_6115,N_6015);
and U6204 (N_6204,N_6095,N_6017);
nor U6205 (N_6205,N_6015,N_6008);
nand U6206 (N_6206,N_6041,N_6094);
and U6207 (N_6207,N_6038,N_6003);
or U6208 (N_6208,N_6020,N_6122);
and U6209 (N_6209,N_6074,N_6094);
nor U6210 (N_6210,N_6115,N_6098);
and U6211 (N_6211,N_6114,N_6031);
and U6212 (N_6212,N_6053,N_6038);
nor U6213 (N_6213,N_6069,N_6117);
and U6214 (N_6214,N_6072,N_6106);
nand U6215 (N_6215,N_6101,N_6123);
nand U6216 (N_6216,N_6115,N_6012);
or U6217 (N_6217,N_6057,N_6061);
nor U6218 (N_6218,N_6112,N_6118);
and U6219 (N_6219,N_6071,N_6009);
and U6220 (N_6220,N_6076,N_6084);
nor U6221 (N_6221,N_6054,N_6007);
nor U6222 (N_6222,N_6119,N_6094);
or U6223 (N_6223,N_6082,N_6036);
nand U6224 (N_6224,N_6066,N_6006);
and U6225 (N_6225,N_6013,N_6049);
and U6226 (N_6226,N_6040,N_6075);
or U6227 (N_6227,N_6001,N_6120);
and U6228 (N_6228,N_6086,N_6029);
nor U6229 (N_6229,N_6025,N_6097);
nand U6230 (N_6230,N_6004,N_6036);
nor U6231 (N_6231,N_6010,N_6019);
xnor U6232 (N_6232,N_6009,N_6004);
and U6233 (N_6233,N_6061,N_6029);
nand U6234 (N_6234,N_6050,N_6006);
xnor U6235 (N_6235,N_6117,N_6000);
nand U6236 (N_6236,N_6061,N_6047);
nand U6237 (N_6237,N_6036,N_6017);
and U6238 (N_6238,N_6124,N_6088);
nor U6239 (N_6239,N_6080,N_6039);
xnor U6240 (N_6240,N_6000,N_6087);
or U6241 (N_6241,N_6008,N_6075);
xor U6242 (N_6242,N_6031,N_6104);
xnor U6243 (N_6243,N_6004,N_6000);
nand U6244 (N_6244,N_6093,N_6095);
or U6245 (N_6245,N_6036,N_6083);
nor U6246 (N_6246,N_6066,N_6086);
nand U6247 (N_6247,N_6083,N_6052);
and U6248 (N_6248,N_6039,N_6112);
nor U6249 (N_6249,N_6120,N_6096);
and U6250 (N_6250,N_6140,N_6147);
nand U6251 (N_6251,N_6204,N_6156);
or U6252 (N_6252,N_6181,N_6155);
nand U6253 (N_6253,N_6143,N_6167);
xor U6254 (N_6254,N_6223,N_6221);
nor U6255 (N_6255,N_6174,N_6135);
and U6256 (N_6256,N_6212,N_6226);
nand U6257 (N_6257,N_6232,N_6131);
or U6258 (N_6258,N_6228,N_6241);
nor U6259 (N_6259,N_6187,N_6242);
and U6260 (N_6260,N_6125,N_6165);
xor U6261 (N_6261,N_6216,N_6200);
or U6262 (N_6262,N_6153,N_6206);
or U6263 (N_6263,N_6136,N_6133);
nor U6264 (N_6264,N_6126,N_6183);
or U6265 (N_6265,N_6130,N_6248);
nor U6266 (N_6266,N_6168,N_6154);
and U6267 (N_6267,N_6235,N_6182);
nor U6268 (N_6268,N_6246,N_6176);
and U6269 (N_6269,N_6243,N_6230);
nor U6270 (N_6270,N_6218,N_6207);
and U6271 (N_6271,N_6178,N_6198);
or U6272 (N_6272,N_6129,N_6161);
or U6273 (N_6273,N_6148,N_6146);
xnor U6274 (N_6274,N_6138,N_6215);
xor U6275 (N_6275,N_6247,N_6249);
xor U6276 (N_6276,N_6240,N_6175);
and U6277 (N_6277,N_6202,N_6211);
nand U6278 (N_6278,N_6185,N_6231);
xnor U6279 (N_6279,N_6137,N_6160);
nor U6280 (N_6280,N_6186,N_6225);
or U6281 (N_6281,N_6224,N_6166);
nand U6282 (N_6282,N_6162,N_6203);
xnor U6283 (N_6283,N_6149,N_6213);
nand U6284 (N_6284,N_6188,N_6141);
xnor U6285 (N_6285,N_6239,N_6194);
nand U6286 (N_6286,N_6134,N_6150);
nand U6287 (N_6287,N_6205,N_6157);
or U6288 (N_6288,N_6234,N_6192);
nand U6289 (N_6289,N_6171,N_6193);
and U6290 (N_6290,N_6236,N_6169);
or U6291 (N_6291,N_6163,N_6229);
nor U6292 (N_6292,N_6144,N_6173);
nand U6293 (N_6293,N_6158,N_6196);
nand U6294 (N_6294,N_6151,N_6245);
or U6295 (N_6295,N_6172,N_6217);
and U6296 (N_6296,N_6139,N_6238);
and U6297 (N_6297,N_6210,N_6177);
or U6298 (N_6298,N_6244,N_6179);
or U6299 (N_6299,N_6190,N_6197);
xor U6300 (N_6300,N_6127,N_6222);
and U6301 (N_6301,N_6220,N_6195);
nand U6302 (N_6302,N_6189,N_6208);
nand U6303 (N_6303,N_6227,N_6201);
nand U6304 (N_6304,N_6219,N_6142);
and U6305 (N_6305,N_6164,N_6214);
and U6306 (N_6306,N_6128,N_6132);
and U6307 (N_6307,N_6184,N_6159);
or U6308 (N_6308,N_6233,N_6170);
and U6309 (N_6309,N_6145,N_6237);
nand U6310 (N_6310,N_6199,N_6152);
xnor U6311 (N_6311,N_6209,N_6191);
or U6312 (N_6312,N_6180,N_6151);
and U6313 (N_6313,N_6224,N_6183);
or U6314 (N_6314,N_6186,N_6177);
nor U6315 (N_6315,N_6130,N_6215);
xnor U6316 (N_6316,N_6148,N_6150);
nor U6317 (N_6317,N_6237,N_6230);
or U6318 (N_6318,N_6204,N_6241);
nand U6319 (N_6319,N_6219,N_6205);
nor U6320 (N_6320,N_6218,N_6200);
and U6321 (N_6321,N_6244,N_6172);
nor U6322 (N_6322,N_6241,N_6183);
nand U6323 (N_6323,N_6191,N_6167);
xor U6324 (N_6324,N_6205,N_6211);
or U6325 (N_6325,N_6201,N_6240);
and U6326 (N_6326,N_6177,N_6194);
nor U6327 (N_6327,N_6158,N_6191);
nor U6328 (N_6328,N_6170,N_6174);
nor U6329 (N_6329,N_6219,N_6148);
nor U6330 (N_6330,N_6224,N_6142);
xor U6331 (N_6331,N_6165,N_6211);
nor U6332 (N_6332,N_6224,N_6204);
nand U6333 (N_6333,N_6148,N_6220);
and U6334 (N_6334,N_6239,N_6172);
nor U6335 (N_6335,N_6249,N_6184);
or U6336 (N_6336,N_6222,N_6230);
or U6337 (N_6337,N_6133,N_6218);
xor U6338 (N_6338,N_6178,N_6221);
and U6339 (N_6339,N_6176,N_6234);
or U6340 (N_6340,N_6133,N_6217);
and U6341 (N_6341,N_6190,N_6183);
or U6342 (N_6342,N_6185,N_6228);
nand U6343 (N_6343,N_6178,N_6214);
nand U6344 (N_6344,N_6142,N_6215);
and U6345 (N_6345,N_6167,N_6248);
nor U6346 (N_6346,N_6155,N_6236);
and U6347 (N_6347,N_6199,N_6211);
xnor U6348 (N_6348,N_6140,N_6150);
or U6349 (N_6349,N_6195,N_6128);
xor U6350 (N_6350,N_6179,N_6150);
xnor U6351 (N_6351,N_6142,N_6190);
xor U6352 (N_6352,N_6231,N_6203);
or U6353 (N_6353,N_6242,N_6233);
xnor U6354 (N_6354,N_6227,N_6244);
xor U6355 (N_6355,N_6137,N_6206);
xnor U6356 (N_6356,N_6225,N_6208);
nand U6357 (N_6357,N_6233,N_6187);
nor U6358 (N_6358,N_6168,N_6186);
and U6359 (N_6359,N_6230,N_6146);
and U6360 (N_6360,N_6150,N_6242);
or U6361 (N_6361,N_6190,N_6133);
and U6362 (N_6362,N_6191,N_6235);
and U6363 (N_6363,N_6215,N_6126);
xor U6364 (N_6364,N_6141,N_6182);
nand U6365 (N_6365,N_6202,N_6172);
nand U6366 (N_6366,N_6214,N_6140);
and U6367 (N_6367,N_6154,N_6175);
and U6368 (N_6368,N_6139,N_6133);
nor U6369 (N_6369,N_6158,N_6194);
or U6370 (N_6370,N_6204,N_6234);
or U6371 (N_6371,N_6170,N_6200);
xnor U6372 (N_6372,N_6169,N_6233);
and U6373 (N_6373,N_6171,N_6164);
nor U6374 (N_6374,N_6230,N_6134);
nor U6375 (N_6375,N_6310,N_6364);
nor U6376 (N_6376,N_6360,N_6257);
and U6377 (N_6377,N_6262,N_6327);
and U6378 (N_6378,N_6302,N_6279);
and U6379 (N_6379,N_6367,N_6368);
xnor U6380 (N_6380,N_6321,N_6260);
nand U6381 (N_6381,N_6306,N_6316);
or U6382 (N_6382,N_6251,N_6338);
or U6383 (N_6383,N_6303,N_6370);
xnor U6384 (N_6384,N_6344,N_6340);
or U6385 (N_6385,N_6274,N_6334);
or U6386 (N_6386,N_6280,N_6269);
nor U6387 (N_6387,N_6284,N_6304);
nand U6388 (N_6388,N_6352,N_6325);
xor U6389 (N_6389,N_6372,N_6319);
xnor U6390 (N_6390,N_6286,N_6362);
and U6391 (N_6391,N_6264,N_6265);
or U6392 (N_6392,N_6361,N_6293);
xor U6393 (N_6393,N_6369,N_6341);
or U6394 (N_6394,N_6353,N_6301);
and U6395 (N_6395,N_6343,N_6261);
nor U6396 (N_6396,N_6258,N_6282);
nor U6397 (N_6397,N_6328,N_6305);
or U6398 (N_6398,N_6339,N_6296);
nand U6399 (N_6399,N_6289,N_6326);
nand U6400 (N_6400,N_6288,N_6324);
and U6401 (N_6401,N_6287,N_6354);
nand U6402 (N_6402,N_6290,N_6278);
nand U6403 (N_6403,N_6281,N_6313);
nor U6404 (N_6404,N_6263,N_6355);
and U6405 (N_6405,N_6347,N_6317);
nor U6406 (N_6406,N_6314,N_6275);
nand U6407 (N_6407,N_6307,N_6253);
and U6408 (N_6408,N_6291,N_6358);
nor U6409 (N_6409,N_6331,N_6351);
nand U6410 (N_6410,N_6371,N_6270);
or U6411 (N_6411,N_6342,N_6273);
or U6412 (N_6412,N_6322,N_6346);
nand U6413 (N_6413,N_6299,N_6348);
and U6414 (N_6414,N_6276,N_6272);
nor U6415 (N_6415,N_6363,N_6277);
or U6416 (N_6416,N_6312,N_6374);
xor U6417 (N_6417,N_6349,N_6309);
nor U6418 (N_6418,N_6252,N_6356);
nor U6419 (N_6419,N_6336,N_6259);
nor U6420 (N_6420,N_6268,N_6335);
xnor U6421 (N_6421,N_6297,N_6250);
nor U6422 (N_6422,N_6298,N_6323);
nand U6423 (N_6423,N_6320,N_6266);
nor U6424 (N_6424,N_6318,N_6366);
and U6425 (N_6425,N_6359,N_6271);
nor U6426 (N_6426,N_6329,N_6333);
nand U6427 (N_6427,N_6373,N_6315);
xor U6428 (N_6428,N_6283,N_6308);
xor U6429 (N_6429,N_6300,N_6295);
and U6430 (N_6430,N_6332,N_6345);
xnor U6431 (N_6431,N_6311,N_6267);
nand U6432 (N_6432,N_6337,N_6256);
nor U6433 (N_6433,N_6255,N_6330);
or U6434 (N_6434,N_6365,N_6294);
nor U6435 (N_6435,N_6254,N_6285);
nor U6436 (N_6436,N_6292,N_6357);
or U6437 (N_6437,N_6350,N_6360);
nand U6438 (N_6438,N_6282,N_6359);
and U6439 (N_6439,N_6276,N_6303);
and U6440 (N_6440,N_6294,N_6268);
or U6441 (N_6441,N_6319,N_6272);
xor U6442 (N_6442,N_6358,N_6279);
nor U6443 (N_6443,N_6267,N_6357);
nand U6444 (N_6444,N_6371,N_6305);
and U6445 (N_6445,N_6264,N_6327);
or U6446 (N_6446,N_6272,N_6354);
xor U6447 (N_6447,N_6259,N_6312);
nand U6448 (N_6448,N_6294,N_6265);
nand U6449 (N_6449,N_6296,N_6312);
xor U6450 (N_6450,N_6283,N_6257);
nand U6451 (N_6451,N_6284,N_6297);
xnor U6452 (N_6452,N_6321,N_6342);
nor U6453 (N_6453,N_6343,N_6273);
nand U6454 (N_6454,N_6348,N_6292);
and U6455 (N_6455,N_6272,N_6326);
and U6456 (N_6456,N_6262,N_6285);
xnor U6457 (N_6457,N_6343,N_6326);
and U6458 (N_6458,N_6291,N_6271);
xnor U6459 (N_6459,N_6345,N_6333);
nand U6460 (N_6460,N_6279,N_6274);
and U6461 (N_6461,N_6281,N_6334);
and U6462 (N_6462,N_6349,N_6358);
nor U6463 (N_6463,N_6280,N_6314);
nor U6464 (N_6464,N_6290,N_6354);
xnor U6465 (N_6465,N_6369,N_6273);
and U6466 (N_6466,N_6286,N_6270);
xor U6467 (N_6467,N_6366,N_6278);
nand U6468 (N_6468,N_6251,N_6335);
xnor U6469 (N_6469,N_6324,N_6363);
or U6470 (N_6470,N_6319,N_6337);
xor U6471 (N_6471,N_6316,N_6303);
xnor U6472 (N_6472,N_6297,N_6276);
nor U6473 (N_6473,N_6368,N_6353);
or U6474 (N_6474,N_6329,N_6253);
nor U6475 (N_6475,N_6353,N_6262);
nor U6476 (N_6476,N_6299,N_6277);
xnor U6477 (N_6477,N_6333,N_6259);
nor U6478 (N_6478,N_6254,N_6278);
nor U6479 (N_6479,N_6368,N_6350);
or U6480 (N_6480,N_6370,N_6360);
nand U6481 (N_6481,N_6320,N_6374);
or U6482 (N_6482,N_6305,N_6319);
or U6483 (N_6483,N_6374,N_6287);
or U6484 (N_6484,N_6277,N_6321);
nor U6485 (N_6485,N_6275,N_6270);
nor U6486 (N_6486,N_6329,N_6338);
nand U6487 (N_6487,N_6346,N_6369);
nor U6488 (N_6488,N_6325,N_6362);
nor U6489 (N_6489,N_6327,N_6303);
or U6490 (N_6490,N_6328,N_6325);
nand U6491 (N_6491,N_6257,N_6371);
and U6492 (N_6492,N_6266,N_6359);
and U6493 (N_6493,N_6350,N_6374);
nor U6494 (N_6494,N_6265,N_6349);
nor U6495 (N_6495,N_6371,N_6260);
or U6496 (N_6496,N_6334,N_6324);
xor U6497 (N_6497,N_6348,N_6308);
xnor U6498 (N_6498,N_6253,N_6285);
and U6499 (N_6499,N_6281,N_6315);
or U6500 (N_6500,N_6421,N_6465);
nand U6501 (N_6501,N_6459,N_6482);
xor U6502 (N_6502,N_6411,N_6420);
and U6503 (N_6503,N_6432,N_6410);
nand U6504 (N_6504,N_6497,N_6478);
xor U6505 (N_6505,N_6377,N_6495);
and U6506 (N_6506,N_6426,N_6488);
and U6507 (N_6507,N_6448,N_6403);
and U6508 (N_6508,N_6485,N_6415);
nand U6509 (N_6509,N_6423,N_6436);
and U6510 (N_6510,N_6474,N_6491);
and U6511 (N_6511,N_6400,N_6463);
and U6512 (N_6512,N_6425,N_6406);
xnor U6513 (N_6513,N_6422,N_6378);
or U6514 (N_6514,N_6401,N_6455);
nand U6515 (N_6515,N_6392,N_6452);
or U6516 (N_6516,N_6384,N_6483);
nor U6517 (N_6517,N_6379,N_6453);
nand U6518 (N_6518,N_6461,N_6441);
and U6519 (N_6519,N_6434,N_6416);
or U6520 (N_6520,N_6383,N_6430);
nor U6521 (N_6521,N_6417,N_6462);
nor U6522 (N_6522,N_6396,N_6458);
and U6523 (N_6523,N_6380,N_6464);
and U6524 (N_6524,N_6414,N_6428);
nor U6525 (N_6525,N_6493,N_6399);
and U6526 (N_6526,N_6456,N_6443);
nand U6527 (N_6527,N_6389,N_6393);
nor U6528 (N_6528,N_6476,N_6437);
nor U6529 (N_6529,N_6447,N_6446);
and U6530 (N_6530,N_6398,N_6468);
nor U6531 (N_6531,N_6382,N_6466);
xor U6532 (N_6532,N_6407,N_6460);
and U6533 (N_6533,N_6376,N_6454);
or U6534 (N_6534,N_6405,N_6472);
xor U6535 (N_6535,N_6487,N_6467);
or U6536 (N_6536,N_6469,N_6387);
nor U6537 (N_6537,N_6494,N_6397);
nor U6538 (N_6538,N_6409,N_6438);
nand U6539 (N_6539,N_6386,N_6433);
and U6540 (N_6540,N_6489,N_6402);
or U6541 (N_6541,N_6427,N_6490);
nand U6542 (N_6542,N_6424,N_6470);
nand U6543 (N_6543,N_6475,N_6499);
nand U6544 (N_6544,N_6381,N_6419);
nand U6545 (N_6545,N_6484,N_6385);
xor U6546 (N_6546,N_6471,N_6457);
xor U6547 (N_6547,N_6435,N_6449);
nand U6548 (N_6548,N_6477,N_6480);
nand U6549 (N_6549,N_6440,N_6375);
xor U6550 (N_6550,N_6429,N_6451);
or U6551 (N_6551,N_6473,N_6486);
or U6552 (N_6552,N_6394,N_6388);
xor U6553 (N_6553,N_6390,N_6450);
nor U6554 (N_6554,N_6395,N_6496);
or U6555 (N_6555,N_6479,N_6412);
or U6556 (N_6556,N_6408,N_6492);
nor U6557 (N_6557,N_6444,N_6404);
or U6558 (N_6558,N_6391,N_6413);
nor U6559 (N_6559,N_6418,N_6431);
nand U6560 (N_6560,N_6439,N_6481);
xnor U6561 (N_6561,N_6498,N_6445);
nand U6562 (N_6562,N_6442,N_6459);
nand U6563 (N_6563,N_6407,N_6434);
xor U6564 (N_6564,N_6480,N_6439);
nand U6565 (N_6565,N_6401,N_6435);
nor U6566 (N_6566,N_6442,N_6478);
nor U6567 (N_6567,N_6499,N_6457);
nand U6568 (N_6568,N_6475,N_6394);
xor U6569 (N_6569,N_6391,N_6426);
xnor U6570 (N_6570,N_6475,N_6457);
and U6571 (N_6571,N_6376,N_6476);
nor U6572 (N_6572,N_6488,N_6473);
or U6573 (N_6573,N_6479,N_6415);
and U6574 (N_6574,N_6471,N_6380);
xor U6575 (N_6575,N_6488,N_6402);
or U6576 (N_6576,N_6398,N_6481);
nand U6577 (N_6577,N_6414,N_6490);
or U6578 (N_6578,N_6431,N_6450);
xor U6579 (N_6579,N_6433,N_6415);
and U6580 (N_6580,N_6410,N_6455);
and U6581 (N_6581,N_6408,N_6402);
xor U6582 (N_6582,N_6475,N_6417);
nand U6583 (N_6583,N_6435,N_6496);
nand U6584 (N_6584,N_6490,N_6429);
or U6585 (N_6585,N_6468,N_6466);
xor U6586 (N_6586,N_6414,N_6440);
or U6587 (N_6587,N_6409,N_6465);
nor U6588 (N_6588,N_6442,N_6382);
nand U6589 (N_6589,N_6381,N_6425);
xnor U6590 (N_6590,N_6388,N_6467);
or U6591 (N_6591,N_6495,N_6431);
and U6592 (N_6592,N_6440,N_6426);
nor U6593 (N_6593,N_6448,N_6423);
xnor U6594 (N_6594,N_6436,N_6464);
and U6595 (N_6595,N_6395,N_6441);
nor U6596 (N_6596,N_6406,N_6491);
nor U6597 (N_6597,N_6429,N_6489);
xnor U6598 (N_6598,N_6381,N_6472);
xor U6599 (N_6599,N_6413,N_6441);
or U6600 (N_6600,N_6494,N_6492);
or U6601 (N_6601,N_6494,N_6470);
nor U6602 (N_6602,N_6465,N_6459);
nand U6603 (N_6603,N_6462,N_6408);
nand U6604 (N_6604,N_6496,N_6467);
nor U6605 (N_6605,N_6384,N_6388);
xor U6606 (N_6606,N_6380,N_6406);
nor U6607 (N_6607,N_6409,N_6411);
nor U6608 (N_6608,N_6412,N_6399);
xor U6609 (N_6609,N_6445,N_6425);
and U6610 (N_6610,N_6407,N_6459);
or U6611 (N_6611,N_6468,N_6380);
nand U6612 (N_6612,N_6407,N_6386);
nor U6613 (N_6613,N_6461,N_6390);
or U6614 (N_6614,N_6472,N_6443);
nor U6615 (N_6615,N_6445,N_6383);
nand U6616 (N_6616,N_6437,N_6377);
nand U6617 (N_6617,N_6468,N_6381);
and U6618 (N_6618,N_6442,N_6427);
nand U6619 (N_6619,N_6447,N_6499);
nand U6620 (N_6620,N_6461,N_6478);
or U6621 (N_6621,N_6452,N_6465);
xor U6622 (N_6622,N_6436,N_6380);
xor U6623 (N_6623,N_6432,N_6473);
and U6624 (N_6624,N_6458,N_6431);
nand U6625 (N_6625,N_6517,N_6526);
or U6626 (N_6626,N_6581,N_6547);
nand U6627 (N_6627,N_6616,N_6593);
and U6628 (N_6628,N_6588,N_6500);
xor U6629 (N_6629,N_6503,N_6569);
nand U6630 (N_6630,N_6617,N_6521);
and U6631 (N_6631,N_6546,N_6505);
and U6632 (N_6632,N_6577,N_6591);
nand U6633 (N_6633,N_6557,N_6540);
and U6634 (N_6634,N_6544,N_6606);
or U6635 (N_6635,N_6536,N_6559);
nand U6636 (N_6636,N_6548,N_6598);
or U6637 (N_6637,N_6599,N_6549);
xnor U6638 (N_6638,N_6524,N_6613);
and U6639 (N_6639,N_6600,N_6501);
nor U6640 (N_6640,N_6513,N_6534);
nor U6641 (N_6641,N_6595,N_6525);
xor U6642 (N_6642,N_6572,N_6535);
nor U6643 (N_6643,N_6565,N_6570);
and U6644 (N_6644,N_6612,N_6596);
or U6645 (N_6645,N_6543,N_6550);
xor U6646 (N_6646,N_6597,N_6576);
nand U6647 (N_6647,N_6506,N_6589);
or U6648 (N_6648,N_6519,N_6518);
xor U6649 (N_6649,N_6527,N_6584);
nor U6650 (N_6650,N_6563,N_6532);
or U6651 (N_6651,N_6514,N_6578);
nand U6652 (N_6652,N_6562,N_6515);
or U6653 (N_6653,N_6571,N_6554);
and U6654 (N_6654,N_6539,N_6507);
xnor U6655 (N_6655,N_6528,N_6582);
or U6656 (N_6656,N_6583,N_6622);
and U6657 (N_6657,N_6620,N_6510);
nor U6658 (N_6658,N_6541,N_6556);
and U6659 (N_6659,N_6545,N_6566);
nand U6660 (N_6660,N_6608,N_6512);
nor U6661 (N_6661,N_6611,N_6522);
nand U6662 (N_6662,N_6533,N_6603);
nand U6663 (N_6663,N_6624,N_6586);
or U6664 (N_6664,N_6553,N_6551);
nor U6665 (N_6665,N_6511,N_6552);
or U6666 (N_6666,N_6567,N_6579);
or U6667 (N_6667,N_6575,N_6558);
or U6668 (N_6668,N_6604,N_6614);
or U6669 (N_6669,N_6504,N_6594);
or U6670 (N_6670,N_6580,N_6523);
or U6671 (N_6671,N_6538,N_6509);
xnor U6672 (N_6672,N_6516,N_6615);
nand U6673 (N_6673,N_6531,N_6508);
nand U6674 (N_6674,N_6621,N_6587);
nor U6675 (N_6675,N_6529,N_6590);
nand U6676 (N_6676,N_6605,N_6537);
xnor U6677 (N_6677,N_6574,N_6530);
nand U6678 (N_6678,N_6610,N_6609);
nand U6679 (N_6679,N_6619,N_6623);
or U6680 (N_6680,N_6601,N_6555);
or U6681 (N_6681,N_6568,N_6560);
nand U6682 (N_6682,N_6602,N_6607);
nand U6683 (N_6683,N_6561,N_6573);
nand U6684 (N_6684,N_6618,N_6502);
or U6685 (N_6685,N_6564,N_6542);
and U6686 (N_6686,N_6585,N_6520);
nand U6687 (N_6687,N_6592,N_6539);
xnor U6688 (N_6688,N_6555,N_6604);
nor U6689 (N_6689,N_6568,N_6587);
or U6690 (N_6690,N_6542,N_6621);
and U6691 (N_6691,N_6527,N_6574);
or U6692 (N_6692,N_6557,N_6539);
nor U6693 (N_6693,N_6535,N_6618);
xnor U6694 (N_6694,N_6553,N_6585);
or U6695 (N_6695,N_6562,N_6534);
or U6696 (N_6696,N_6593,N_6529);
and U6697 (N_6697,N_6570,N_6566);
nand U6698 (N_6698,N_6530,N_6572);
nand U6699 (N_6699,N_6515,N_6580);
or U6700 (N_6700,N_6578,N_6533);
or U6701 (N_6701,N_6507,N_6505);
nand U6702 (N_6702,N_6556,N_6615);
or U6703 (N_6703,N_6562,N_6542);
xnor U6704 (N_6704,N_6587,N_6524);
or U6705 (N_6705,N_6526,N_6524);
xnor U6706 (N_6706,N_6571,N_6510);
or U6707 (N_6707,N_6539,N_6590);
nand U6708 (N_6708,N_6598,N_6564);
nor U6709 (N_6709,N_6588,N_6503);
and U6710 (N_6710,N_6578,N_6583);
nand U6711 (N_6711,N_6601,N_6517);
and U6712 (N_6712,N_6569,N_6616);
nor U6713 (N_6713,N_6545,N_6576);
nor U6714 (N_6714,N_6563,N_6543);
xor U6715 (N_6715,N_6572,N_6533);
nor U6716 (N_6716,N_6570,N_6526);
nand U6717 (N_6717,N_6568,N_6600);
and U6718 (N_6718,N_6522,N_6542);
and U6719 (N_6719,N_6595,N_6501);
and U6720 (N_6720,N_6516,N_6534);
nand U6721 (N_6721,N_6617,N_6518);
nand U6722 (N_6722,N_6525,N_6588);
nor U6723 (N_6723,N_6607,N_6597);
or U6724 (N_6724,N_6501,N_6506);
or U6725 (N_6725,N_6619,N_6531);
xor U6726 (N_6726,N_6539,N_6618);
or U6727 (N_6727,N_6604,N_6567);
xor U6728 (N_6728,N_6560,N_6522);
nor U6729 (N_6729,N_6502,N_6520);
xor U6730 (N_6730,N_6570,N_6585);
xnor U6731 (N_6731,N_6518,N_6585);
and U6732 (N_6732,N_6607,N_6564);
xor U6733 (N_6733,N_6540,N_6536);
xor U6734 (N_6734,N_6585,N_6619);
nor U6735 (N_6735,N_6619,N_6561);
xnor U6736 (N_6736,N_6586,N_6601);
xor U6737 (N_6737,N_6554,N_6500);
and U6738 (N_6738,N_6569,N_6568);
nand U6739 (N_6739,N_6533,N_6587);
nor U6740 (N_6740,N_6539,N_6573);
nand U6741 (N_6741,N_6606,N_6579);
nor U6742 (N_6742,N_6557,N_6579);
and U6743 (N_6743,N_6618,N_6511);
xor U6744 (N_6744,N_6581,N_6579);
or U6745 (N_6745,N_6508,N_6500);
and U6746 (N_6746,N_6521,N_6620);
nor U6747 (N_6747,N_6561,N_6530);
nand U6748 (N_6748,N_6545,N_6556);
nor U6749 (N_6749,N_6517,N_6507);
and U6750 (N_6750,N_6733,N_6720);
xnor U6751 (N_6751,N_6678,N_6650);
and U6752 (N_6752,N_6696,N_6704);
or U6753 (N_6753,N_6698,N_6694);
nor U6754 (N_6754,N_6746,N_6711);
or U6755 (N_6755,N_6643,N_6743);
nor U6756 (N_6756,N_6684,N_6697);
and U6757 (N_6757,N_6744,N_6709);
and U6758 (N_6758,N_6625,N_6737);
xnor U6759 (N_6759,N_6652,N_6740);
or U6760 (N_6760,N_6707,N_6675);
or U6761 (N_6761,N_6725,N_6679);
or U6762 (N_6762,N_6681,N_6638);
or U6763 (N_6763,N_6708,N_6637);
xnor U6764 (N_6764,N_6686,N_6721);
and U6765 (N_6765,N_6644,N_6736);
xnor U6766 (N_6766,N_6648,N_6685);
xnor U6767 (N_6767,N_6723,N_6661);
nand U6768 (N_6768,N_6722,N_6664);
xnor U6769 (N_6769,N_6739,N_6668);
xor U6770 (N_6770,N_6651,N_6626);
or U6771 (N_6771,N_6689,N_6674);
nor U6772 (N_6772,N_6730,N_6646);
xnor U6773 (N_6773,N_6749,N_6640);
xnor U6774 (N_6774,N_6692,N_6635);
and U6775 (N_6775,N_6691,N_6690);
xnor U6776 (N_6776,N_6688,N_6731);
nand U6777 (N_6777,N_6683,N_6706);
xor U6778 (N_6778,N_6647,N_6734);
nor U6779 (N_6779,N_6702,N_6670);
xor U6780 (N_6780,N_6636,N_6666);
and U6781 (N_6781,N_6672,N_6732);
and U6782 (N_6782,N_6717,N_6710);
nor U6783 (N_6783,N_6662,N_6735);
nand U6784 (N_6784,N_6659,N_6695);
xnor U6785 (N_6785,N_6639,N_6649);
nand U6786 (N_6786,N_6715,N_6727);
nand U6787 (N_6787,N_6671,N_6656);
or U6788 (N_6788,N_6700,N_6642);
xnor U6789 (N_6789,N_6745,N_6645);
and U6790 (N_6790,N_6655,N_6687);
nand U6791 (N_6791,N_6673,N_6653);
and U6792 (N_6792,N_6631,N_6713);
nor U6793 (N_6793,N_6634,N_6705);
nor U6794 (N_6794,N_6701,N_6728);
and U6795 (N_6795,N_6724,N_6663);
or U6796 (N_6796,N_6627,N_6658);
or U6797 (N_6797,N_6693,N_6680);
or U6798 (N_6798,N_6667,N_6677);
nor U6799 (N_6799,N_6629,N_6729);
and U6800 (N_6800,N_6654,N_6719);
nor U6801 (N_6801,N_6676,N_6748);
nand U6802 (N_6802,N_6741,N_6738);
nand U6803 (N_6803,N_6726,N_6641);
xor U6804 (N_6804,N_6660,N_6718);
nand U6805 (N_6805,N_6669,N_6633);
or U6806 (N_6806,N_6714,N_6657);
or U6807 (N_6807,N_6628,N_6712);
nor U6808 (N_6808,N_6742,N_6716);
nor U6809 (N_6809,N_6747,N_6632);
nand U6810 (N_6810,N_6665,N_6682);
nand U6811 (N_6811,N_6703,N_6630);
xor U6812 (N_6812,N_6699,N_6665);
nand U6813 (N_6813,N_6737,N_6676);
nand U6814 (N_6814,N_6683,N_6643);
and U6815 (N_6815,N_6707,N_6646);
or U6816 (N_6816,N_6630,N_6683);
nand U6817 (N_6817,N_6748,N_6740);
and U6818 (N_6818,N_6743,N_6696);
and U6819 (N_6819,N_6670,N_6651);
or U6820 (N_6820,N_6634,N_6640);
nor U6821 (N_6821,N_6671,N_6681);
xnor U6822 (N_6822,N_6702,N_6672);
nand U6823 (N_6823,N_6636,N_6746);
xor U6824 (N_6824,N_6651,N_6636);
xor U6825 (N_6825,N_6702,N_6675);
and U6826 (N_6826,N_6714,N_6674);
nand U6827 (N_6827,N_6671,N_6699);
xnor U6828 (N_6828,N_6648,N_6635);
and U6829 (N_6829,N_6722,N_6749);
xor U6830 (N_6830,N_6739,N_6641);
nand U6831 (N_6831,N_6730,N_6710);
nor U6832 (N_6832,N_6642,N_6731);
xnor U6833 (N_6833,N_6680,N_6667);
nor U6834 (N_6834,N_6639,N_6710);
and U6835 (N_6835,N_6742,N_6652);
nor U6836 (N_6836,N_6657,N_6677);
or U6837 (N_6837,N_6644,N_6628);
or U6838 (N_6838,N_6681,N_6748);
nand U6839 (N_6839,N_6695,N_6671);
or U6840 (N_6840,N_6626,N_6737);
or U6841 (N_6841,N_6724,N_6719);
and U6842 (N_6842,N_6686,N_6667);
nor U6843 (N_6843,N_6713,N_6723);
xnor U6844 (N_6844,N_6687,N_6627);
nand U6845 (N_6845,N_6625,N_6746);
xor U6846 (N_6846,N_6690,N_6749);
nand U6847 (N_6847,N_6629,N_6653);
nor U6848 (N_6848,N_6738,N_6737);
or U6849 (N_6849,N_6626,N_6710);
nor U6850 (N_6850,N_6649,N_6682);
xnor U6851 (N_6851,N_6677,N_6703);
nand U6852 (N_6852,N_6663,N_6679);
xnor U6853 (N_6853,N_6656,N_6717);
nor U6854 (N_6854,N_6632,N_6662);
and U6855 (N_6855,N_6697,N_6729);
nand U6856 (N_6856,N_6699,N_6737);
xor U6857 (N_6857,N_6665,N_6659);
nor U6858 (N_6858,N_6656,N_6737);
or U6859 (N_6859,N_6652,N_6705);
nand U6860 (N_6860,N_6669,N_6645);
or U6861 (N_6861,N_6700,N_6701);
or U6862 (N_6862,N_6652,N_6665);
xnor U6863 (N_6863,N_6636,N_6708);
or U6864 (N_6864,N_6736,N_6671);
and U6865 (N_6865,N_6722,N_6694);
nor U6866 (N_6866,N_6698,N_6659);
or U6867 (N_6867,N_6641,N_6664);
nor U6868 (N_6868,N_6677,N_6628);
and U6869 (N_6869,N_6676,N_6668);
xor U6870 (N_6870,N_6746,N_6668);
nand U6871 (N_6871,N_6669,N_6734);
xnor U6872 (N_6872,N_6641,N_6670);
xor U6873 (N_6873,N_6710,N_6683);
or U6874 (N_6874,N_6742,N_6670);
nand U6875 (N_6875,N_6790,N_6794);
or U6876 (N_6876,N_6796,N_6761);
nor U6877 (N_6877,N_6789,N_6867);
or U6878 (N_6878,N_6871,N_6780);
nand U6879 (N_6879,N_6792,N_6852);
nor U6880 (N_6880,N_6754,N_6764);
nor U6881 (N_6881,N_6870,N_6837);
and U6882 (N_6882,N_6799,N_6822);
and U6883 (N_6883,N_6844,N_6843);
xnor U6884 (N_6884,N_6853,N_6866);
nand U6885 (N_6885,N_6856,N_6816);
nand U6886 (N_6886,N_6830,N_6858);
or U6887 (N_6887,N_6766,N_6833);
nor U6888 (N_6888,N_6762,N_6842);
nand U6889 (N_6889,N_6759,N_6810);
or U6890 (N_6890,N_6820,N_6801);
or U6891 (N_6891,N_6851,N_6765);
or U6892 (N_6892,N_6828,N_6786);
or U6893 (N_6893,N_6781,N_6873);
and U6894 (N_6894,N_6859,N_6845);
nand U6895 (N_6895,N_6753,N_6763);
xor U6896 (N_6896,N_6834,N_6756);
or U6897 (N_6897,N_6791,N_6836);
nand U6898 (N_6898,N_6768,N_6751);
and U6899 (N_6899,N_6798,N_6862);
nand U6900 (N_6900,N_6868,N_6802);
and U6901 (N_6901,N_6841,N_6803);
or U6902 (N_6902,N_6777,N_6850);
or U6903 (N_6903,N_6874,N_6819);
nor U6904 (N_6904,N_6847,N_6869);
xor U6905 (N_6905,N_6776,N_6865);
nand U6906 (N_6906,N_6872,N_6752);
nor U6907 (N_6907,N_6857,N_6808);
or U6908 (N_6908,N_6797,N_6784);
xor U6909 (N_6909,N_6832,N_6806);
nand U6910 (N_6910,N_6771,N_6825);
or U6911 (N_6911,N_6758,N_6757);
nor U6912 (N_6912,N_6779,N_6795);
nand U6913 (N_6913,N_6783,N_6849);
nand U6914 (N_6914,N_6827,N_6778);
nand U6915 (N_6915,N_6774,N_6826);
nand U6916 (N_6916,N_6773,N_6846);
xnor U6917 (N_6917,N_6814,N_6785);
or U6918 (N_6918,N_6812,N_6755);
nor U6919 (N_6919,N_6860,N_6823);
nand U6920 (N_6920,N_6760,N_6817);
or U6921 (N_6921,N_6804,N_6775);
nand U6922 (N_6922,N_6767,N_6809);
or U6923 (N_6923,N_6811,N_6831);
and U6924 (N_6924,N_6788,N_6824);
or U6925 (N_6925,N_6838,N_6815);
nor U6926 (N_6926,N_6848,N_6787);
and U6927 (N_6927,N_6782,N_6863);
xnor U6928 (N_6928,N_6770,N_6813);
xor U6929 (N_6929,N_6805,N_6821);
nor U6930 (N_6930,N_6861,N_6840);
xor U6931 (N_6931,N_6772,N_6835);
xor U6932 (N_6932,N_6750,N_6854);
and U6933 (N_6933,N_6769,N_6829);
nand U6934 (N_6934,N_6807,N_6839);
nand U6935 (N_6935,N_6855,N_6864);
xor U6936 (N_6936,N_6818,N_6793);
nand U6937 (N_6937,N_6800,N_6820);
and U6938 (N_6938,N_6794,N_6762);
or U6939 (N_6939,N_6757,N_6844);
or U6940 (N_6940,N_6846,N_6763);
or U6941 (N_6941,N_6804,N_6845);
and U6942 (N_6942,N_6841,N_6830);
nand U6943 (N_6943,N_6812,N_6858);
and U6944 (N_6944,N_6798,N_6796);
or U6945 (N_6945,N_6855,N_6800);
xor U6946 (N_6946,N_6754,N_6825);
and U6947 (N_6947,N_6809,N_6851);
nor U6948 (N_6948,N_6811,N_6752);
or U6949 (N_6949,N_6833,N_6828);
and U6950 (N_6950,N_6854,N_6820);
xnor U6951 (N_6951,N_6851,N_6873);
nand U6952 (N_6952,N_6800,N_6805);
or U6953 (N_6953,N_6761,N_6808);
or U6954 (N_6954,N_6757,N_6765);
nor U6955 (N_6955,N_6825,N_6818);
nand U6956 (N_6956,N_6763,N_6781);
xnor U6957 (N_6957,N_6766,N_6789);
xnor U6958 (N_6958,N_6758,N_6805);
nand U6959 (N_6959,N_6872,N_6817);
and U6960 (N_6960,N_6800,N_6846);
or U6961 (N_6961,N_6765,N_6872);
and U6962 (N_6962,N_6781,N_6770);
xnor U6963 (N_6963,N_6764,N_6795);
or U6964 (N_6964,N_6864,N_6826);
xor U6965 (N_6965,N_6759,N_6824);
xor U6966 (N_6966,N_6871,N_6788);
xnor U6967 (N_6967,N_6823,N_6869);
nand U6968 (N_6968,N_6854,N_6834);
nand U6969 (N_6969,N_6817,N_6795);
nor U6970 (N_6970,N_6854,N_6775);
nor U6971 (N_6971,N_6761,N_6836);
xor U6972 (N_6972,N_6770,N_6818);
nand U6973 (N_6973,N_6778,N_6813);
nand U6974 (N_6974,N_6810,N_6790);
nor U6975 (N_6975,N_6755,N_6866);
or U6976 (N_6976,N_6842,N_6853);
or U6977 (N_6977,N_6820,N_6847);
nand U6978 (N_6978,N_6860,N_6752);
and U6979 (N_6979,N_6803,N_6759);
nor U6980 (N_6980,N_6760,N_6816);
or U6981 (N_6981,N_6806,N_6777);
nor U6982 (N_6982,N_6810,N_6805);
nand U6983 (N_6983,N_6845,N_6787);
or U6984 (N_6984,N_6817,N_6860);
nand U6985 (N_6985,N_6788,N_6811);
xor U6986 (N_6986,N_6817,N_6750);
nor U6987 (N_6987,N_6827,N_6779);
and U6988 (N_6988,N_6780,N_6872);
or U6989 (N_6989,N_6864,N_6807);
xnor U6990 (N_6990,N_6829,N_6824);
xor U6991 (N_6991,N_6766,N_6771);
or U6992 (N_6992,N_6840,N_6775);
nand U6993 (N_6993,N_6864,N_6832);
and U6994 (N_6994,N_6802,N_6865);
or U6995 (N_6995,N_6868,N_6768);
or U6996 (N_6996,N_6870,N_6860);
and U6997 (N_6997,N_6798,N_6873);
and U6998 (N_6998,N_6835,N_6803);
or U6999 (N_6999,N_6863,N_6763);
nor U7000 (N_7000,N_6927,N_6906);
nand U7001 (N_7001,N_6982,N_6948);
xor U7002 (N_7002,N_6888,N_6967);
nand U7003 (N_7003,N_6878,N_6909);
nand U7004 (N_7004,N_6917,N_6955);
and U7005 (N_7005,N_6926,N_6968);
xor U7006 (N_7006,N_6987,N_6995);
xor U7007 (N_7007,N_6953,N_6876);
xnor U7008 (N_7008,N_6929,N_6935);
or U7009 (N_7009,N_6957,N_6974);
nand U7010 (N_7010,N_6951,N_6881);
or U7011 (N_7011,N_6898,N_6885);
nand U7012 (N_7012,N_6941,N_6994);
and U7013 (N_7013,N_6914,N_6972);
xnor U7014 (N_7014,N_6923,N_6999);
nor U7015 (N_7015,N_6933,N_6983);
nand U7016 (N_7016,N_6936,N_6961);
xor U7017 (N_7017,N_6997,N_6945);
xnor U7018 (N_7018,N_6976,N_6954);
nand U7019 (N_7019,N_6894,N_6977);
or U7020 (N_7020,N_6934,N_6942);
nand U7021 (N_7021,N_6964,N_6877);
and U7022 (N_7022,N_6993,N_6883);
or U7023 (N_7023,N_6899,N_6886);
xnor U7024 (N_7024,N_6890,N_6922);
nand U7025 (N_7025,N_6882,N_6973);
and U7026 (N_7026,N_6978,N_6902);
and U7027 (N_7027,N_6921,N_6998);
xnor U7028 (N_7028,N_6988,N_6875);
xnor U7029 (N_7029,N_6981,N_6912);
nor U7030 (N_7030,N_6958,N_6918);
and U7031 (N_7031,N_6956,N_6986);
xor U7032 (N_7032,N_6901,N_6897);
nand U7033 (N_7033,N_6992,N_6970);
xnor U7034 (N_7034,N_6907,N_6893);
or U7035 (N_7035,N_6880,N_6925);
and U7036 (N_7036,N_6965,N_6971);
nor U7037 (N_7037,N_6900,N_6931);
xnor U7038 (N_7038,N_6946,N_6947);
nor U7039 (N_7039,N_6944,N_6891);
and U7040 (N_7040,N_6963,N_6979);
nor U7041 (N_7041,N_6905,N_6989);
or U7042 (N_7042,N_6908,N_6915);
xor U7043 (N_7043,N_6928,N_6990);
or U7044 (N_7044,N_6916,N_6949);
or U7045 (N_7045,N_6924,N_6950);
nand U7046 (N_7046,N_6904,N_6903);
or U7047 (N_7047,N_6889,N_6938);
or U7048 (N_7048,N_6959,N_6932);
nor U7049 (N_7049,N_6975,N_6884);
and U7050 (N_7050,N_6887,N_6937);
xnor U7051 (N_7051,N_6991,N_6939);
xnor U7052 (N_7052,N_6960,N_6940);
xor U7053 (N_7053,N_6879,N_6952);
xnor U7054 (N_7054,N_6985,N_6910);
and U7055 (N_7055,N_6969,N_6996);
nand U7056 (N_7056,N_6984,N_6896);
nor U7057 (N_7057,N_6966,N_6920);
nand U7058 (N_7058,N_6895,N_6930);
xor U7059 (N_7059,N_6919,N_6943);
and U7060 (N_7060,N_6962,N_6911);
and U7061 (N_7061,N_6913,N_6892);
xor U7062 (N_7062,N_6980,N_6963);
nand U7063 (N_7063,N_6920,N_6970);
xor U7064 (N_7064,N_6907,N_6939);
and U7065 (N_7065,N_6996,N_6937);
nor U7066 (N_7066,N_6882,N_6981);
or U7067 (N_7067,N_6954,N_6886);
xnor U7068 (N_7068,N_6998,N_6964);
and U7069 (N_7069,N_6952,N_6975);
xnor U7070 (N_7070,N_6884,N_6930);
and U7071 (N_7071,N_6978,N_6895);
or U7072 (N_7072,N_6893,N_6955);
nand U7073 (N_7073,N_6929,N_6995);
xor U7074 (N_7074,N_6880,N_6881);
nor U7075 (N_7075,N_6912,N_6936);
or U7076 (N_7076,N_6936,N_6890);
and U7077 (N_7077,N_6927,N_6983);
nand U7078 (N_7078,N_6942,N_6888);
and U7079 (N_7079,N_6963,N_6928);
xor U7080 (N_7080,N_6960,N_6958);
nor U7081 (N_7081,N_6889,N_6895);
nor U7082 (N_7082,N_6876,N_6966);
xor U7083 (N_7083,N_6952,N_6951);
nor U7084 (N_7084,N_6947,N_6958);
xor U7085 (N_7085,N_6879,N_6953);
xnor U7086 (N_7086,N_6934,N_6977);
or U7087 (N_7087,N_6912,N_6993);
or U7088 (N_7088,N_6941,N_6973);
or U7089 (N_7089,N_6998,N_6989);
nor U7090 (N_7090,N_6999,N_6884);
and U7091 (N_7091,N_6986,N_6994);
nand U7092 (N_7092,N_6890,N_6973);
or U7093 (N_7093,N_6890,N_6969);
or U7094 (N_7094,N_6920,N_6983);
xnor U7095 (N_7095,N_6877,N_6932);
nand U7096 (N_7096,N_6918,N_6886);
and U7097 (N_7097,N_6987,N_6893);
or U7098 (N_7098,N_6885,N_6890);
and U7099 (N_7099,N_6947,N_6875);
xor U7100 (N_7100,N_6919,N_6958);
and U7101 (N_7101,N_6939,N_6943);
nand U7102 (N_7102,N_6887,N_6904);
or U7103 (N_7103,N_6985,N_6917);
nand U7104 (N_7104,N_6930,N_6910);
xor U7105 (N_7105,N_6934,N_6943);
nor U7106 (N_7106,N_6884,N_6905);
nor U7107 (N_7107,N_6884,N_6977);
or U7108 (N_7108,N_6879,N_6951);
xnor U7109 (N_7109,N_6939,N_6949);
xor U7110 (N_7110,N_6916,N_6929);
and U7111 (N_7111,N_6990,N_6946);
xnor U7112 (N_7112,N_6903,N_6882);
or U7113 (N_7113,N_6923,N_6990);
xnor U7114 (N_7114,N_6897,N_6938);
xor U7115 (N_7115,N_6884,N_6984);
xor U7116 (N_7116,N_6885,N_6990);
or U7117 (N_7117,N_6893,N_6986);
nor U7118 (N_7118,N_6958,N_6979);
or U7119 (N_7119,N_6936,N_6978);
and U7120 (N_7120,N_6898,N_6937);
nand U7121 (N_7121,N_6915,N_6988);
xor U7122 (N_7122,N_6926,N_6877);
nand U7123 (N_7123,N_6934,N_6881);
or U7124 (N_7124,N_6931,N_6880);
and U7125 (N_7125,N_7119,N_7073);
or U7126 (N_7126,N_7091,N_7087);
and U7127 (N_7127,N_7090,N_7021);
nor U7128 (N_7128,N_7032,N_7061);
or U7129 (N_7129,N_7059,N_7107);
and U7130 (N_7130,N_7044,N_7049);
and U7131 (N_7131,N_7072,N_7067);
nand U7132 (N_7132,N_7030,N_7106);
or U7133 (N_7133,N_7028,N_7024);
and U7134 (N_7134,N_7015,N_7054);
or U7135 (N_7135,N_7041,N_7010);
nor U7136 (N_7136,N_7113,N_7085);
or U7137 (N_7137,N_7017,N_7114);
xnor U7138 (N_7138,N_7084,N_7004);
xnor U7139 (N_7139,N_7120,N_7071);
or U7140 (N_7140,N_7093,N_7124);
and U7141 (N_7141,N_7042,N_7052);
xor U7142 (N_7142,N_7047,N_7063);
and U7143 (N_7143,N_7023,N_7108);
or U7144 (N_7144,N_7011,N_7116);
nand U7145 (N_7145,N_7051,N_7080);
or U7146 (N_7146,N_7038,N_7065);
or U7147 (N_7147,N_7097,N_7100);
nor U7148 (N_7148,N_7053,N_7086);
nand U7149 (N_7149,N_7070,N_7083);
xor U7150 (N_7150,N_7092,N_7013);
xor U7151 (N_7151,N_7068,N_7082);
nor U7152 (N_7152,N_7104,N_7101);
nor U7153 (N_7153,N_7098,N_7029);
and U7154 (N_7154,N_7007,N_7027);
xnor U7155 (N_7155,N_7094,N_7046);
xor U7156 (N_7156,N_7062,N_7048);
and U7157 (N_7157,N_7025,N_7075);
or U7158 (N_7158,N_7074,N_7018);
and U7159 (N_7159,N_7031,N_7112);
nor U7160 (N_7160,N_7055,N_7123);
nor U7161 (N_7161,N_7026,N_7008);
or U7162 (N_7162,N_7109,N_7060);
and U7163 (N_7163,N_7036,N_7020);
xor U7164 (N_7164,N_7105,N_7096);
xnor U7165 (N_7165,N_7079,N_7064);
xnor U7166 (N_7166,N_7043,N_7099);
nor U7167 (N_7167,N_7102,N_7005);
or U7168 (N_7168,N_7034,N_7006);
or U7169 (N_7169,N_7089,N_7122);
nand U7170 (N_7170,N_7022,N_7081);
nand U7171 (N_7171,N_7000,N_7040);
and U7172 (N_7172,N_7095,N_7066);
and U7173 (N_7173,N_7077,N_7057);
nand U7174 (N_7174,N_7117,N_7012);
xor U7175 (N_7175,N_7001,N_7118);
nand U7176 (N_7176,N_7039,N_7088);
nand U7177 (N_7177,N_7076,N_7103);
or U7178 (N_7178,N_7016,N_7069);
nor U7179 (N_7179,N_7121,N_7111);
nor U7180 (N_7180,N_7056,N_7014);
or U7181 (N_7181,N_7037,N_7019);
or U7182 (N_7182,N_7050,N_7115);
and U7183 (N_7183,N_7003,N_7009);
nand U7184 (N_7184,N_7045,N_7058);
and U7185 (N_7185,N_7035,N_7002);
nand U7186 (N_7186,N_7033,N_7110);
xor U7187 (N_7187,N_7078,N_7093);
or U7188 (N_7188,N_7084,N_7039);
and U7189 (N_7189,N_7121,N_7123);
nor U7190 (N_7190,N_7056,N_7098);
and U7191 (N_7191,N_7020,N_7053);
xnor U7192 (N_7192,N_7010,N_7034);
xnor U7193 (N_7193,N_7093,N_7090);
and U7194 (N_7194,N_7082,N_7102);
xnor U7195 (N_7195,N_7032,N_7062);
nand U7196 (N_7196,N_7103,N_7041);
and U7197 (N_7197,N_7111,N_7015);
and U7198 (N_7198,N_7041,N_7038);
and U7199 (N_7199,N_7044,N_7032);
xor U7200 (N_7200,N_7048,N_7094);
and U7201 (N_7201,N_7078,N_7011);
nor U7202 (N_7202,N_7026,N_7095);
or U7203 (N_7203,N_7001,N_7002);
xor U7204 (N_7204,N_7036,N_7047);
nand U7205 (N_7205,N_7015,N_7026);
nor U7206 (N_7206,N_7008,N_7030);
nand U7207 (N_7207,N_7107,N_7124);
nor U7208 (N_7208,N_7029,N_7012);
nand U7209 (N_7209,N_7003,N_7057);
nor U7210 (N_7210,N_7048,N_7053);
nor U7211 (N_7211,N_7118,N_7015);
nor U7212 (N_7212,N_7076,N_7016);
or U7213 (N_7213,N_7115,N_7106);
nor U7214 (N_7214,N_7093,N_7016);
and U7215 (N_7215,N_7023,N_7027);
nand U7216 (N_7216,N_7014,N_7039);
or U7217 (N_7217,N_7006,N_7114);
nor U7218 (N_7218,N_7098,N_7118);
xnor U7219 (N_7219,N_7123,N_7115);
and U7220 (N_7220,N_7094,N_7023);
and U7221 (N_7221,N_7009,N_7090);
nor U7222 (N_7222,N_7048,N_7105);
and U7223 (N_7223,N_7010,N_7095);
xor U7224 (N_7224,N_7077,N_7027);
xnor U7225 (N_7225,N_7026,N_7037);
or U7226 (N_7226,N_7001,N_7099);
nand U7227 (N_7227,N_7002,N_7034);
or U7228 (N_7228,N_7011,N_7067);
or U7229 (N_7229,N_7102,N_7110);
nand U7230 (N_7230,N_7106,N_7032);
or U7231 (N_7231,N_7046,N_7011);
nor U7232 (N_7232,N_7062,N_7122);
or U7233 (N_7233,N_7054,N_7032);
xor U7234 (N_7234,N_7119,N_7050);
and U7235 (N_7235,N_7068,N_7075);
and U7236 (N_7236,N_7091,N_7054);
nor U7237 (N_7237,N_7024,N_7074);
xor U7238 (N_7238,N_7025,N_7108);
nand U7239 (N_7239,N_7023,N_7035);
nand U7240 (N_7240,N_7121,N_7076);
or U7241 (N_7241,N_7115,N_7110);
xor U7242 (N_7242,N_7048,N_7088);
or U7243 (N_7243,N_7092,N_7006);
xnor U7244 (N_7244,N_7110,N_7101);
nand U7245 (N_7245,N_7084,N_7081);
xnor U7246 (N_7246,N_7091,N_7081);
nand U7247 (N_7247,N_7036,N_7121);
nor U7248 (N_7248,N_7117,N_7053);
or U7249 (N_7249,N_7060,N_7010);
nand U7250 (N_7250,N_7153,N_7196);
or U7251 (N_7251,N_7172,N_7178);
and U7252 (N_7252,N_7199,N_7132);
or U7253 (N_7253,N_7232,N_7246);
nand U7254 (N_7254,N_7181,N_7228);
or U7255 (N_7255,N_7194,N_7164);
and U7256 (N_7256,N_7218,N_7221);
nand U7257 (N_7257,N_7203,N_7226);
xnor U7258 (N_7258,N_7127,N_7209);
nand U7259 (N_7259,N_7236,N_7234);
and U7260 (N_7260,N_7242,N_7126);
and U7261 (N_7261,N_7185,N_7141);
xor U7262 (N_7262,N_7139,N_7193);
or U7263 (N_7263,N_7195,N_7150);
nor U7264 (N_7264,N_7171,N_7204);
nand U7265 (N_7265,N_7208,N_7245);
and U7266 (N_7266,N_7128,N_7187);
or U7267 (N_7267,N_7148,N_7248);
xor U7268 (N_7268,N_7176,N_7244);
and U7269 (N_7269,N_7147,N_7129);
xor U7270 (N_7270,N_7175,N_7184);
nand U7271 (N_7271,N_7180,N_7151);
and U7272 (N_7272,N_7169,N_7125);
nor U7273 (N_7273,N_7222,N_7217);
nor U7274 (N_7274,N_7238,N_7225);
nand U7275 (N_7275,N_7201,N_7186);
or U7276 (N_7276,N_7130,N_7131);
or U7277 (N_7277,N_7163,N_7231);
nand U7278 (N_7278,N_7198,N_7212);
or U7279 (N_7279,N_7134,N_7211);
nor U7280 (N_7280,N_7219,N_7136);
and U7281 (N_7281,N_7240,N_7189);
nor U7282 (N_7282,N_7177,N_7192);
or U7283 (N_7283,N_7162,N_7233);
or U7284 (N_7284,N_7156,N_7207);
or U7285 (N_7285,N_7224,N_7182);
nor U7286 (N_7286,N_7243,N_7216);
nand U7287 (N_7287,N_7214,N_7154);
xor U7288 (N_7288,N_7247,N_7229);
nor U7289 (N_7289,N_7145,N_7188);
and U7290 (N_7290,N_7168,N_7140);
and U7291 (N_7291,N_7142,N_7149);
and U7292 (N_7292,N_7210,N_7179);
nor U7293 (N_7293,N_7166,N_7206);
nor U7294 (N_7294,N_7190,N_7183);
and U7295 (N_7295,N_7197,N_7146);
nand U7296 (N_7296,N_7215,N_7133);
nor U7297 (N_7297,N_7161,N_7167);
or U7298 (N_7298,N_7160,N_7173);
xor U7299 (N_7299,N_7205,N_7152);
and U7300 (N_7300,N_7158,N_7165);
xnor U7301 (N_7301,N_7174,N_7227);
nand U7302 (N_7302,N_7230,N_7241);
and U7303 (N_7303,N_7239,N_7143);
xor U7304 (N_7304,N_7135,N_7137);
and U7305 (N_7305,N_7191,N_7157);
nor U7306 (N_7306,N_7200,N_7249);
and U7307 (N_7307,N_7155,N_7138);
xnor U7308 (N_7308,N_7170,N_7220);
xnor U7309 (N_7309,N_7235,N_7223);
xor U7310 (N_7310,N_7159,N_7237);
xnor U7311 (N_7311,N_7144,N_7213);
and U7312 (N_7312,N_7202,N_7232);
nand U7313 (N_7313,N_7131,N_7218);
nor U7314 (N_7314,N_7208,N_7178);
nor U7315 (N_7315,N_7217,N_7193);
nor U7316 (N_7316,N_7243,N_7233);
or U7317 (N_7317,N_7136,N_7153);
or U7318 (N_7318,N_7161,N_7247);
nand U7319 (N_7319,N_7210,N_7177);
nand U7320 (N_7320,N_7142,N_7198);
and U7321 (N_7321,N_7203,N_7156);
or U7322 (N_7322,N_7233,N_7178);
and U7323 (N_7323,N_7191,N_7170);
nand U7324 (N_7324,N_7191,N_7190);
and U7325 (N_7325,N_7237,N_7150);
and U7326 (N_7326,N_7227,N_7237);
and U7327 (N_7327,N_7211,N_7226);
nand U7328 (N_7328,N_7238,N_7196);
and U7329 (N_7329,N_7144,N_7170);
and U7330 (N_7330,N_7142,N_7201);
nor U7331 (N_7331,N_7187,N_7221);
xnor U7332 (N_7332,N_7196,N_7200);
xor U7333 (N_7333,N_7235,N_7184);
xnor U7334 (N_7334,N_7147,N_7189);
or U7335 (N_7335,N_7159,N_7126);
or U7336 (N_7336,N_7134,N_7166);
and U7337 (N_7337,N_7229,N_7243);
and U7338 (N_7338,N_7244,N_7146);
nor U7339 (N_7339,N_7209,N_7166);
xnor U7340 (N_7340,N_7187,N_7182);
or U7341 (N_7341,N_7142,N_7228);
nor U7342 (N_7342,N_7130,N_7187);
or U7343 (N_7343,N_7175,N_7219);
xor U7344 (N_7344,N_7184,N_7178);
nor U7345 (N_7345,N_7169,N_7179);
and U7346 (N_7346,N_7225,N_7199);
xor U7347 (N_7347,N_7138,N_7166);
nand U7348 (N_7348,N_7163,N_7218);
nand U7349 (N_7349,N_7216,N_7165);
and U7350 (N_7350,N_7229,N_7153);
xnor U7351 (N_7351,N_7163,N_7241);
xnor U7352 (N_7352,N_7206,N_7226);
and U7353 (N_7353,N_7242,N_7163);
xnor U7354 (N_7354,N_7209,N_7152);
nor U7355 (N_7355,N_7248,N_7178);
xor U7356 (N_7356,N_7159,N_7209);
and U7357 (N_7357,N_7161,N_7226);
nor U7358 (N_7358,N_7149,N_7206);
xnor U7359 (N_7359,N_7138,N_7205);
and U7360 (N_7360,N_7203,N_7141);
or U7361 (N_7361,N_7167,N_7187);
nand U7362 (N_7362,N_7233,N_7238);
nor U7363 (N_7363,N_7205,N_7170);
and U7364 (N_7364,N_7208,N_7184);
nor U7365 (N_7365,N_7179,N_7129);
and U7366 (N_7366,N_7232,N_7145);
and U7367 (N_7367,N_7168,N_7209);
or U7368 (N_7368,N_7130,N_7240);
xnor U7369 (N_7369,N_7142,N_7217);
or U7370 (N_7370,N_7135,N_7192);
and U7371 (N_7371,N_7231,N_7189);
or U7372 (N_7372,N_7203,N_7150);
and U7373 (N_7373,N_7136,N_7155);
and U7374 (N_7374,N_7141,N_7131);
and U7375 (N_7375,N_7363,N_7273);
xor U7376 (N_7376,N_7366,N_7311);
or U7377 (N_7377,N_7339,N_7261);
nor U7378 (N_7378,N_7283,N_7316);
or U7379 (N_7379,N_7351,N_7251);
nand U7380 (N_7380,N_7270,N_7319);
xor U7381 (N_7381,N_7272,N_7275);
xor U7382 (N_7382,N_7269,N_7356);
or U7383 (N_7383,N_7320,N_7347);
nor U7384 (N_7384,N_7262,N_7300);
and U7385 (N_7385,N_7292,N_7335);
nor U7386 (N_7386,N_7352,N_7312);
xor U7387 (N_7387,N_7253,N_7284);
nand U7388 (N_7388,N_7294,N_7289);
nand U7389 (N_7389,N_7370,N_7343);
or U7390 (N_7390,N_7345,N_7328);
or U7391 (N_7391,N_7288,N_7252);
and U7392 (N_7392,N_7260,N_7274);
xor U7393 (N_7393,N_7341,N_7333);
and U7394 (N_7394,N_7340,N_7315);
and U7395 (N_7395,N_7271,N_7280);
or U7396 (N_7396,N_7301,N_7346);
nor U7397 (N_7397,N_7338,N_7327);
xor U7398 (N_7398,N_7368,N_7317);
or U7399 (N_7399,N_7364,N_7255);
nor U7400 (N_7400,N_7296,N_7293);
nor U7401 (N_7401,N_7277,N_7325);
xor U7402 (N_7402,N_7314,N_7329);
or U7403 (N_7403,N_7265,N_7279);
xnor U7404 (N_7404,N_7302,N_7323);
and U7405 (N_7405,N_7344,N_7374);
and U7406 (N_7406,N_7290,N_7304);
or U7407 (N_7407,N_7254,N_7295);
nand U7408 (N_7408,N_7281,N_7258);
nand U7409 (N_7409,N_7362,N_7359);
nand U7410 (N_7410,N_7305,N_7267);
and U7411 (N_7411,N_7334,N_7318);
or U7412 (N_7412,N_7257,N_7259);
or U7413 (N_7413,N_7342,N_7256);
and U7414 (N_7414,N_7326,N_7310);
and U7415 (N_7415,N_7360,N_7336);
or U7416 (N_7416,N_7307,N_7285);
xnor U7417 (N_7417,N_7306,N_7299);
xnor U7418 (N_7418,N_7291,N_7324);
xnor U7419 (N_7419,N_7357,N_7353);
and U7420 (N_7420,N_7358,N_7263);
and U7421 (N_7421,N_7297,N_7266);
xor U7422 (N_7422,N_7264,N_7354);
nand U7423 (N_7423,N_7349,N_7321);
nor U7424 (N_7424,N_7331,N_7287);
nand U7425 (N_7425,N_7286,N_7348);
and U7426 (N_7426,N_7313,N_7282);
or U7427 (N_7427,N_7303,N_7372);
nor U7428 (N_7428,N_7332,N_7250);
or U7429 (N_7429,N_7276,N_7365);
and U7430 (N_7430,N_7373,N_7350);
and U7431 (N_7431,N_7322,N_7268);
nand U7432 (N_7432,N_7308,N_7371);
and U7433 (N_7433,N_7355,N_7369);
nand U7434 (N_7434,N_7330,N_7337);
and U7435 (N_7435,N_7298,N_7309);
and U7436 (N_7436,N_7278,N_7361);
xnor U7437 (N_7437,N_7367,N_7350);
nor U7438 (N_7438,N_7317,N_7269);
nand U7439 (N_7439,N_7305,N_7253);
nor U7440 (N_7440,N_7348,N_7274);
nor U7441 (N_7441,N_7356,N_7280);
xnor U7442 (N_7442,N_7374,N_7263);
or U7443 (N_7443,N_7368,N_7321);
and U7444 (N_7444,N_7314,N_7302);
or U7445 (N_7445,N_7328,N_7317);
nor U7446 (N_7446,N_7309,N_7307);
or U7447 (N_7447,N_7350,N_7362);
xnor U7448 (N_7448,N_7277,N_7304);
xnor U7449 (N_7449,N_7270,N_7300);
nand U7450 (N_7450,N_7287,N_7280);
xnor U7451 (N_7451,N_7336,N_7268);
nand U7452 (N_7452,N_7289,N_7359);
nand U7453 (N_7453,N_7356,N_7308);
nand U7454 (N_7454,N_7364,N_7254);
xnor U7455 (N_7455,N_7291,N_7277);
xor U7456 (N_7456,N_7362,N_7367);
xnor U7457 (N_7457,N_7330,N_7252);
and U7458 (N_7458,N_7296,N_7361);
xor U7459 (N_7459,N_7269,N_7288);
xnor U7460 (N_7460,N_7258,N_7270);
nor U7461 (N_7461,N_7277,N_7346);
xor U7462 (N_7462,N_7332,N_7313);
nor U7463 (N_7463,N_7340,N_7259);
and U7464 (N_7464,N_7273,N_7337);
xnor U7465 (N_7465,N_7335,N_7254);
and U7466 (N_7466,N_7331,N_7329);
nand U7467 (N_7467,N_7351,N_7335);
and U7468 (N_7468,N_7330,N_7268);
nand U7469 (N_7469,N_7272,N_7373);
nand U7470 (N_7470,N_7277,N_7349);
nor U7471 (N_7471,N_7355,N_7351);
xnor U7472 (N_7472,N_7372,N_7286);
nor U7473 (N_7473,N_7329,N_7319);
nand U7474 (N_7474,N_7313,N_7287);
xnor U7475 (N_7475,N_7266,N_7281);
or U7476 (N_7476,N_7307,N_7284);
nand U7477 (N_7477,N_7279,N_7314);
xnor U7478 (N_7478,N_7253,N_7276);
and U7479 (N_7479,N_7348,N_7345);
and U7480 (N_7480,N_7278,N_7337);
nand U7481 (N_7481,N_7358,N_7282);
or U7482 (N_7482,N_7256,N_7313);
nor U7483 (N_7483,N_7304,N_7317);
xor U7484 (N_7484,N_7254,N_7260);
nand U7485 (N_7485,N_7308,N_7324);
and U7486 (N_7486,N_7309,N_7279);
xor U7487 (N_7487,N_7274,N_7328);
or U7488 (N_7488,N_7344,N_7336);
xor U7489 (N_7489,N_7252,N_7274);
and U7490 (N_7490,N_7308,N_7251);
xnor U7491 (N_7491,N_7290,N_7294);
and U7492 (N_7492,N_7355,N_7346);
nor U7493 (N_7493,N_7320,N_7331);
xor U7494 (N_7494,N_7265,N_7259);
and U7495 (N_7495,N_7338,N_7314);
and U7496 (N_7496,N_7360,N_7309);
nor U7497 (N_7497,N_7295,N_7346);
or U7498 (N_7498,N_7280,N_7256);
xor U7499 (N_7499,N_7353,N_7342);
and U7500 (N_7500,N_7409,N_7425);
and U7501 (N_7501,N_7419,N_7451);
nand U7502 (N_7502,N_7388,N_7412);
xor U7503 (N_7503,N_7407,N_7395);
nand U7504 (N_7504,N_7455,N_7443);
nand U7505 (N_7505,N_7440,N_7488);
and U7506 (N_7506,N_7394,N_7447);
and U7507 (N_7507,N_7384,N_7452);
nor U7508 (N_7508,N_7450,N_7418);
nor U7509 (N_7509,N_7415,N_7390);
or U7510 (N_7510,N_7435,N_7422);
nor U7511 (N_7511,N_7434,N_7438);
nor U7512 (N_7512,N_7411,N_7480);
xnor U7513 (N_7513,N_7385,N_7483);
and U7514 (N_7514,N_7423,N_7458);
nor U7515 (N_7515,N_7485,N_7466);
or U7516 (N_7516,N_7470,N_7389);
or U7517 (N_7517,N_7437,N_7469);
nor U7518 (N_7518,N_7499,N_7392);
and U7519 (N_7519,N_7424,N_7404);
nor U7520 (N_7520,N_7401,N_7377);
xnor U7521 (N_7521,N_7433,N_7459);
or U7522 (N_7522,N_7448,N_7465);
and U7523 (N_7523,N_7479,N_7454);
nand U7524 (N_7524,N_7382,N_7387);
xor U7525 (N_7525,N_7474,N_7399);
nor U7526 (N_7526,N_7428,N_7376);
nand U7527 (N_7527,N_7468,N_7472);
nand U7528 (N_7528,N_7402,N_7431);
nor U7529 (N_7529,N_7498,N_7383);
or U7530 (N_7530,N_7453,N_7493);
nand U7531 (N_7531,N_7491,N_7490);
nor U7532 (N_7532,N_7496,N_7445);
nor U7533 (N_7533,N_7497,N_7439);
nor U7534 (N_7534,N_7430,N_7464);
xor U7535 (N_7535,N_7386,N_7410);
nand U7536 (N_7536,N_7403,N_7420);
and U7537 (N_7537,N_7473,N_7489);
nand U7538 (N_7538,N_7432,N_7408);
xnor U7539 (N_7539,N_7380,N_7475);
nand U7540 (N_7540,N_7476,N_7446);
nand U7541 (N_7541,N_7416,N_7456);
nand U7542 (N_7542,N_7495,N_7413);
xor U7543 (N_7543,N_7484,N_7494);
nand U7544 (N_7544,N_7405,N_7487);
nand U7545 (N_7545,N_7463,N_7481);
nor U7546 (N_7546,N_7426,N_7477);
nand U7547 (N_7547,N_7375,N_7471);
and U7548 (N_7548,N_7460,N_7478);
and U7549 (N_7549,N_7414,N_7442);
and U7550 (N_7550,N_7393,N_7444);
nand U7551 (N_7551,N_7449,N_7397);
nand U7552 (N_7552,N_7400,N_7406);
and U7553 (N_7553,N_7429,N_7486);
or U7554 (N_7554,N_7396,N_7391);
nand U7555 (N_7555,N_7492,N_7378);
xor U7556 (N_7556,N_7398,N_7441);
nand U7557 (N_7557,N_7436,N_7421);
and U7558 (N_7558,N_7381,N_7457);
nor U7559 (N_7559,N_7462,N_7461);
xor U7560 (N_7560,N_7427,N_7467);
nand U7561 (N_7561,N_7417,N_7482);
nor U7562 (N_7562,N_7379,N_7437);
nor U7563 (N_7563,N_7420,N_7481);
and U7564 (N_7564,N_7452,N_7434);
xnor U7565 (N_7565,N_7395,N_7472);
and U7566 (N_7566,N_7437,N_7492);
nand U7567 (N_7567,N_7421,N_7452);
and U7568 (N_7568,N_7454,N_7389);
nor U7569 (N_7569,N_7393,N_7480);
and U7570 (N_7570,N_7390,N_7434);
xor U7571 (N_7571,N_7425,N_7460);
nor U7572 (N_7572,N_7461,N_7496);
nand U7573 (N_7573,N_7457,N_7386);
nor U7574 (N_7574,N_7408,N_7463);
or U7575 (N_7575,N_7426,N_7424);
or U7576 (N_7576,N_7493,N_7402);
or U7577 (N_7577,N_7417,N_7435);
nand U7578 (N_7578,N_7486,N_7454);
nor U7579 (N_7579,N_7388,N_7485);
or U7580 (N_7580,N_7460,N_7421);
and U7581 (N_7581,N_7435,N_7446);
or U7582 (N_7582,N_7485,N_7473);
nand U7583 (N_7583,N_7382,N_7412);
or U7584 (N_7584,N_7417,N_7439);
nor U7585 (N_7585,N_7398,N_7382);
nand U7586 (N_7586,N_7396,N_7447);
nand U7587 (N_7587,N_7378,N_7395);
or U7588 (N_7588,N_7432,N_7470);
nor U7589 (N_7589,N_7446,N_7436);
xnor U7590 (N_7590,N_7412,N_7483);
xnor U7591 (N_7591,N_7396,N_7495);
xor U7592 (N_7592,N_7401,N_7473);
or U7593 (N_7593,N_7387,N_7404);
or U7594 (N_7594,N_7474,N_7460);
nor U7595 (N_7595,N_7479,N_7498);
and U7596 (N_7596,N_7422,N_7404);
xnor U7597 (N_7597,N_7428,N_7484);
and U7598 (N_7598,N_7460,N_7415);
xnor U7599 (N_7599,N_7422,N_7387);
nor U7600 (N_7600,N_7461,N_7394);
nor U7601 (N_7601,N_7453,N_7415);
nand U7602 (N_7602,N_7481,N_7449);
nand U7603 (N_7603,N_7440,N_7451);
nand U7604 (N_7604,N_7480,N_7383);
nor U7605 (N_7605,N_7429,N_7451);
or U7606 (N_7606,N_7493,N_7406);
xnor U7607 (N_7607,N_7490,N_7480);
and U7608 (N_7608,N_7475,N_7440);
and U7609 (N_7609,N_7498,N_7441);
or U7610 (N_7610,N_7454,N_7420);
nand U7611 (N_7611,N_7469,N_7379);
and U7612 (N_7612,N_7470,N_7486);
and U7613 (N_7613,N_7380,N_7387);
and U7614 (N_7614,N_7401,N_7472);
or U7615 (N_7615,N_7408,N_7425);
and U7616 (N_7616,N_7418,N_7496);
nor U7617 (N_7617,N_7375,N_7425);
and U7618 (N_7618,N_7448,N_7435);
or U7619 (N_7619,N_7465,N_7405);
nand U7620 (N_7620,N_7486,N_7481);
or U7621 (N_7621,N_7387,N_7406);
or U7622 (N_7622,N_7422,N_7476);
nand U7623 (N_7623,N_7465,N_7403);
and U7624 (N_7624,N_7399,N_7381);
nor U7625 (N_7625,N_7513,N_7609);
and U7626 (N_7626,N_7548,N_7611);
nor U7627 (N_7627,N_7524,N_7599);
or U7628 (N_7628,N_7571,N_7575);
nor U7629 (N_7629,N_7557,N_7560);
xor U7630 (N_7630,N_7546,N_7556);
or U7631 (N_7631,N_7563,N_7578);
nand U7632 (N_7632,N_7586,N_7504);
nand U7633 (N_7633,N_7606,N_7547);
and U7634 (N_7634,N_7584,N_7543);
xor U7635 (N_7635,N_7596,N_7558);
nand U7636 (N_7636,N_7534,N_7605);
or U7637 (N_7637,N_7589,N_7617);
or U7638 (N_7638,N_7554,N_7500);
xor U7639 (N_7639,N_7529,N_7542);
nand U7640 (N_7640,N_7537,N_7587);
nand U7641 (N_7641,N_7591,N_7572);
nor U7642 (N_7642,N_7614,N_7603);
nor U7643 (N_7643,N_7570,N_7601);
nand U7644 (N_7644,N_7518,N_7510);
nand U7645 (N_7645,N_7574,N_7559);
nor U7646 (N_7646,N_7536,N_7600);
nand U7647 (N_7647,N_7619,N_7527);
or U7648 (N_7648,N_7622,N_7541);
nand U7649 (N_7649,N_7568,N_7576);
and U7650 (N_7650,N_7561,N_7530);
xor U7651 (N_7651,N_7552,N_7506);
nor U7652 (N_7652,N_7612,N_7532);
xor U7653 (N_7653,N_7565,N_7615);
or U7654 (N_7654,N_7526,N_7519);
or U7655 (N_7655,N_7613,N_7585);
and U7656 (N_7656,N_7581,N_7621);
nor U7657 (N_7657,N_7577,N_7567);
xnor U7658 (N_7658,N_7608,N_7593);
xnor U7659 (N_7659,N_7618,N_7604);
xor U7660 (N_7660,N_7623,N_7590);
and U7661 (N_7661,N_7501,N_7594);
nand U7662 (N_7662,N_7509,N_7511);
or U7663 (N_7663,N_7508,N_7515);
xor U7664 (N_7664,N_7514,N_7592);
or U7665 (N_7665,N_7588,N_7569);
xnor U7666 (N_7666,N_7535,N_7573);
nand U7667 (N_7667,N_7522,N_7624);
nand U7668 (N_7668,N_7525,N_7566);
xnor U7669 (N_7669,N_7520,N_7550);
and U7670 (N_7670,N_7580,N_7583);
and U7671 (N_7671,N_7507,N_7533);
or U7672 (N_7672,N_7598,N_7597);
nand U7673 (N_7673,N_7595,N_7607);
nor U7674 (N_7674,N_7551,N_7602);
xor U7675 (N_7675,N_7545,N_7512);
or U7676 (N_7676,N_7531,N_7579);
or U7677 (N_7677,N_7553,N_7503);
or U7678 (N_7678,N_7549,N_7521);
nand U7679 (N_7679,N_7582,N_7540);
nand U7680 (N_7680,N_7620,N_7502);
nand U7681 (N_7681,N_7505,N_7538);
xor U7682 (N_7682,N_7564,N_7562);
xor U7683 (N_7683,N_7544,N_7539);
nand U7684 (N_7684,N_7517,N_7616);
or U7685 (N_7685,N_7528,N_7610);
and U7686 (N_7686,N_7516,N_7523);
xor U7687 (N_7687,N_7555,N_7551);
nor U7688 (N_7688,N_7522,N_7598);
nand U7689 (N_7689,N_7547,N_7601);
and U7690 (N_7690,N_7551,N_7559);
and U7691 (N_7691,N_7619,N_7542);
nor U7692 (N_7692,N_7504,N_7566);
xor U7693 (N_7693,N_7592,N_7598);
nor U7694 (N_7694,N_7582,N_7584);
nor U7695 (N_7695,N_7512,N_7531);
and U7696 (N_7696,N_7579,N_7570);
nand U7697 (N_7697,N_7606,N_7620);
nor U7698 (N_7698,N_7543,N_7570);
and U7699 (N_7699,N_7514,N_7511);
or U7700 (N_7700,N_7624,N_7543);
nor U7701 (N_7701,N_7505,N_7542);
xor U7702 (N_7702,N_7506,N_7618);
or U7703 (N_7703,N_7516,N_7601);
or U7704 (N_7704,N_7568,N_7615);
xnor U7705 (N_7705,N_7544,N_7569);
or U7706 (N_7706,N_7523,N_7597);
or U7707 (N_7707,N_7587,N_7605);
or U7708 (N_7708,N_7579,N_7545);
nand U7709 (N_7709,N_7542,N_7536);
nor U7710 (N_7710,N_7554,N_7511);
nor U7711 (N_7711,N_7619,N_7570);
xor U7712 (N_7712,N_7612,N_7531);
nand U7713 (N_7713,N_7593,N_7536);
and U7714 (N_7714,N_7572,N_7506);
nand U7715 (N_7715,N_7538,N_7516);
xnor U7716 (N_7716,N_7559,N_7572);
nand U7717 (N_7717,N_7552,N_7527);
or U7718 (N_7718,N_7592,N_7508);
or U7719 (N_7719,N_7568,N_7532);
xor U7720 (N_7720,N_7608,N_7616);
or U7721 (N_7721,N_7509,N_7593);
nand U7722 (N_7722,N_7564,N_7533);
or U7723 (N_7723,N_7506,N_7557);
or U7724 (N_7724,N_7548,N_7595);
nand U7725 (N_7725,N_7565,N_7508);
xor U7726 (N_7726,N_7529,N_7607);
xnor U7727 (N_7727,N_7521,N_7535);
or U7728 (N_7728,N_7563,N_7603);
or U7729 (N_7729,N_7554,N_7505);
or U7730 (N_7730,N_7500,N_7514);
nor U7731 (N_7731,N_7521,N_7570);
or U7732 (N_7732,N_7565,N_7571);
and U7733 (N_7733,N_7579,N_7532);
nor U7734 (N_7734,N_7501,N_7605);
xor U7735 (N_7735,N_7585,N_7583);
xor U7736 (N_7736,N_7543,N_7544);
and U7737 (N_7737,N_7617,N_7578);
and U7738 (N_7738,N_7523,N_7587);
and U7739 (N_7739,N_7621,N_7534);
and U7740 (N_7740,N_7607,N_7620);
and U7741 (N_7741,N_7513,N_7602);
or U7742 (N_7742,N_7537,N_7508);
nor U7743 (N_7743,N_7514,N_7605);
nor U7744 (N_7744,N_7551,N_7545);
xor U7745 (N_7745,N_7570,N_7572);
or U7746 (N_7746,N_7587,N_7601);
xor U7747 (N_7747,N_7541,N_7560);
or U7748 (N_7748,N_7529,N_7513);
or U7749 (N_7749,N_7525,N_7526);
nor U7750 (N_7750,N_7664,N_7724);
nand U7751 (N_7751,N_7746,N_7744);
or U7752 (N_7752,N_7709,N_7683);
nor U7753 (N_7753,N_7717,N_7633);
and U7754 (N_7754,N_7642,N_7681);
and U7755 (N_7755,N_7734,N_7736);
nand U7756 (N_7756,N_7728,N_7737);
or U7757 (N_7757,N_7667,N_7695);
or U7758 (N_7758,N_7647,N_7700);
nor U7759 (N_7759,N_7693,N_7722);
or U7760 (N_7760,N_7631,N_7650);
nand U7761 (N_7761,N_7676,N_7696);
nor U7762 (N_7762,N_7723,N_7743);
or U7763 (N_7763,N_7646,N_7662);
nor U7764 (N_7764,N_7718,N_7634);
nand U7765 (N_7765,N_7731,N_7730);
and U7766 (N_7766,N_7705,N_7688);
and U7767 (N_7767,N_7629,N_7686);
or U7768 (N_7768,N_7673,N_7658);
xor U7769 (N_7769,N_7725,N_7745);
nor U7770 (N_7770,N_7716,N_7689);
nor U7771 (N_7771,N_7741,N_7626);
or U7772 (N_7772,N_7733,N_7643);
and U7773 (N_7773,N_7685,N_7721);
xor U7774 (N_7774,N_7641,N_7719);
nor U7775 (N_7775,N_7742,N_7672);
nand U7776 (N_7776,N_7639,N_7694);
nand U7777 (N_7777,N_7714,N_7679);
and U7778 (N_7778,N_7635,N_7627);
nor U7779 (N_7779,N_7657,N_7652);
and U7780 (N_7780,N_7720,N_7653);
nand U7781 (N_7781,N_7748,N_7711);
xnor U7782 (N_7782,N_7677,N_7715);
and U7783 (N_7783,N_7659,N_7645);
and U7784 (N_7784,N_7628,N_7675);
and U7785 (N_7785,N_7727,N_7671);
or U7786 (N_7786,N_7691,N_7638);
or U7787 (N_7787,N_7668,N_7740);
or U7788 (N_7788,N_7713,N_7704);
nand U7789 (N_7789,N_7644,N_7701);
nor U7790 (N_7790,N_7735,N_7706);
or U7791 (N_7791,N_7674,N_7732);
nor U7792 (N_7792,N_7651,N_7697);
xnor U7793 (N_7793,N_7625,N_7699);
nand U7794 (N_7794,N_7710,N_7682);
nand U7795 (N_7795,N_7669,N_7670);
nand U7796 (N_7796,N_7684,N_7747);
xnor U7797 (N_7797,N_7648,N_7649);
xor U7798 (N_7798,N_7692,N_7637);
xor U7799 (N_7799,N_7698,N_7738);
xor U7800 (N_7800,N_7729,N_7749);
nor U7801 (N_7801,N_7708,N_7678);
nor U7802 (N_7802,N_7663,N_7665);
xnor U7803 (N_7803,N_7640,N_7702);
or U7804 (N_7804,N_7630,N_7739);
and U7805 (N_7805,N_7680,N_7703);
xor U7806 (N_7806,N_7666,N_7687);
xor U7807 (N_7807,N_7690,N_7726);
nor U7808 (N_7808,N_7712,N_7636);
nor U7809 (N_7809,N_7655,N_7654);
xnor U7810 (N_7810,N_7661,N_7707);
nand U7811 (N_7811,N_7632,N_7656);
or U7812 (N_7812,N_7660,N_7725);
and U7813 (N_7813,N_7704,N_7701);
xor U7814 (N_7814,N_7632,N_7641);
xnor U7815 (N_7815,N_7649,N_7653);
nor U7816 (N_7816,N_7741,N_7653);
or U7817 (N_7817,N_7692,N_7693);
nor U7818 (N_7818,N_7660,N_7705);
nand U7819 (N_7819,N_7705,N_7637);
xor U7820 (N_7820,N_7636,N_7692);
xnor U7821 (N_7821,N_7722,N_7641);
or U7822 (N_7822,N_7697,N_7741);
nor U7823 (N_7823,N_7658,N_7638);
nor U7824 (N_7824,N_7723,N_7661);
or U7825 (N_7825,N_7728,N_7727);
nor U7826 (N_7826,N_7709,N_7660);
and U7827 (N_7827,N_7633,N_7713);
or U7828 (N_7828,N_7646,N_7749);
xor U7829 (N_7829,N_7701,N_7734);
or U7830 (N_7830,N_7632,N_7629);
nor U7831 (N_7831,N_7742,N_7726);
nand U7832 (N_7832,N_7687,N_7681);
or U7833 (N_7833,N_7625,N_7658);
and U7834 (N_7834,N_7721,N_7718);
xnor U7835 (N_7835,N_7725,N_7641);
or U7836 (N_7836,N_7657,N_7688);
or U7837 (N_7837,N_7705,N_7676);
and U7838 (N_7838,N_7669,N_7731);
and U7839 (N_7839,N_7666,N_7631);
and U7840 (N_7840,N_7662,N_7723);
nand U7841 (N_7841,N_7736,N_7704);
nand U7842 (N_7842,N_7650,N_7712);
xor U7843 (N_7843,N_7721,N_7698);
xnor U7844 (N_7844,N_7634,N_7709);
and U7845 (N_7845,N_7744,N_7681);
and U7846 (N_7846,N_7640,N_7625);
nor U7847 (N_7847,N_7671,N_7668);
xor U7848 (N_7848,N_7639,N_7628);
and U7849 (N_7849,N_7651,N_7739);
and U7850 (N_7850,N_7713,N_7662);
and U7851 (N_7851,N_7633,N_7680);
and U7852 (N_7852,N_7653,N_7637);
or U7853 (N_7853,N_7749,N_7715);
or U7854 (N_7854,N_7694,N_7635);
and U7855 (N_7855,N_7638,N_7727);
or U7856 (N_7856,N_7655,N_7696);
xor U7857 (N_7857,N_7678,N_7641);
and U7858 (N_7858,N_7680,N_7744);
nor U7859 (N_7859,N_7716,N_7649);
xnor U7860 (N_7860,N_7735,N_7656);
or U7861 (N_7861,N_7729,N_7709);
or U7862 (N_7862,N_7633,N_7627);
and U7863 (N_7863,N_7674,N_7713);
nor U7864 (N_7864,N_7732,N_7681);
nor U7865 (N_7865,N_7735,N_7708);
nor U7866 (N_7866,N_7706,N_7627);
nor U7867 (N_7867,N_7660,N_7655);
nand U7868 (N_7868,N_7718,N_7697);
xor U7869 (N_7869,N_7673,N_7696);
nor U7870 (N_7870,N_7669,N_7748);
and U7871 (N_7871,N_7704,N_7632);
and U7872 (N_7872,N_7692,N_7662);
xor U7873 (N_7873,N_7732,N_7739);
or U7874 (N_7874,N_7727,N_7654);
or U7875 (N_7875,N_7843,N_7865);
nor U7876 (N_7876,N_7775,N_7854);
or U7877 (N_7877,N_7817,N_7849);
nor U7878 (N_7878,N_7783,N_7844);
xnor U7879 (N_7879,N_7795,N_7828);
nand U7880 (N_7880,N_7810,N_7769);
nand U7881 (N_7881,N_7848,N_7760);
nor U7882 (N_7882,N_7786,N_7797);
and U7883 (N_7883,N_7829,N_7812);
nor U7884 (N_7884,N_7868,N_7803);
nand U7885 (N_7885,N_7827,N_7867);
nor U7886 (N_7886,N_7825,N_7816);
nand U7887 (N_7887,N_7756,N_7784);
nor U7888 (N_7888,N_7873,N_7826);
and U7889 (N_7889,N_7837,N_7801);
or U7890 (N_7890,N_7766,N_7776);
or U7891 (N_7891,N_7855,N_7840);
xor U7892 (N_7892,N_7869,N_7822);
nand U7893 (N_7893,N_7832,N_7860);
nor U7894 (N_7894,N_7752,N_7830);
or U7895 (N_7895,N_7824,N_7793);
xor U7896 (N_7896,N_7819,N_7778);
nand U7897 (N_7897,N_7792,N_7774);
nand U7898 (N_7898,N_7850,N_7751);
xnor U7899 (N_7899,N_7808,N_7763);
nand U7900 (N_7900,N_7773,N_7862);
or U7901 (N_7901,N_7811,N_7753);
or U7902 (N_7902,N_7762,N_7789);
nand U7903 (N_7903,N_7804,N_7772);
or U7904 (N_7904,N_7799,N_7781);
and U7905 (N_7905,N_7856,N_7821);
and U7906 (N_7906,N_7833,N_7782);
or U7907 (N_7907,N_7761,N_7780);
nand U7908 (N_7908,N_7794,N_7791);
nor U7909 (N_7909,N_7777,N_7785);
nor U7910 (N_7910,N_7770,N_7755);
nand U7911 (N_7911,N_7765,N_7846);
and U7912 (N_7912,N_7767,N_7818);
nor U7913 (N_7913,N_7870,N_7861);
or U7914 (N_7914,N_7863,N_7857);
nor U7915 (N_7915,N_7754,N_7757);
nor U7916 (N_7916,N_7847,N_7788);
xor U7917 (N_7917,N_7866,N_7852);
and U7918 (N_7918,N_7805,N_7758);
and U7919 (N_7919,N_7838,N_7806);
nand U7920 (N_7920,N_7750,N_7851);
nor U7921 (N_7921,N_7815,N_7813);
nand U7922 (N_7922,N_7764,N_7853);
nor U7923 (N_7923,N_7872,N_7800);
nand U7924 (N_7924,N_7807,N_7809);
or U7925 (N_7925,N_7759,N_7836);
or U7926 (N_7926,N_7835,N_7858);
nor U7927 (N_7927,N_7768,N_7771);
nand U7928 (N_7928,N_7779,N_7802);
and U7929 (N_7929,N_7839,N_7859);
or U7930 (N_7930,N_7841,N_7834);
nand U7931 (N_7931,N_7814,N_7845);
and U7932 (N_7932,N_7871,N_7842);
or U7933 (N_7933,N_7874,N_7823);
and U7934 (N_7934,N_7787,N_7864);
nor U7935 (N_7935,N_7790,N_7798);
nand U7936 (N_7936,N_7831,N_7796);
nor U7937 (N_7937,N_7820,N_7836);
nor U7938 (N_7938,N_7855,N_7800);
nor U7939 (N_7939,N_7759,N_7779);
or U7940 (N_7940,N_7789,N_7830);
xnor U7941 (N_7941,N_7810,N_7823);
xor U7942 (N_7942,N_7821,N_7809);
xnor U7943 (N_7943,N_7753,N_7865);
nor U7944 (N_7944,N_7768,N_7798);
xnor U7945 (N_7945,N_7816,N_7839);
or U7946 (N_7946,N_7822,N_7792);
nand U7947 (N_7947,N_7764,N_7861);
and U7948 (N_7948,N_7834,N_7794);
xor U7949 (N_7949,N_7871,N_7788);
and U7950 (N_7950,N_7803,N_7787);
nor U7951 (N_7951,N_7801,N_7848);
or U7952 (N_7952,N_7846,N_7860);
or U7953 (N_7953,N_7791,N_7775);
nor U7954 (N_7954,N_7865,N_7785);
nand U7955 (N_7955,N_7871,N_7757);
nand U7956 (N_7956,N_7775,N_7837);
xor U7957 (N_7957,N_7804,N_7800);
xnor U7958 (N_7958,N_7756,N_7798);
nand U7959 (N_7959,N_7822,N_7821);
nand U7960 (N_7960,N_7755,N_7833);
nand U7961 (N_7961,N_7762,N_7815);
nand U7962 (N_7962,N_7755,N_7816);
and U7963 (N_7963,N_7790,N_7764);
or U7964 (N_7964,N_7838,N_7792);
nor U7965 (N_7965,N_7863,N_7781);
nand U7966 (N_7966,N_7789,N_7836);
and U7967 (N_7967,N_7824,N_7859);
or U7968 (N_7968,N_7752,N_7787);
nor U7969 (N_7969,N_7862,N_7755);
nor U7970 (N_7970,N_7786,N_7783);
nor U7971 (N_7971,N_7753,N_7844);
nand U7972 (N_7972,N_7832,N_7781);
nand U7973 (N_7973,N_7862,N_7764);
xnor U7974 (N_7974,N_7772,N_7852);
nand U7975 (N_7975,N_7836,N_7769);
nand U7976 (N_7976,N_7768,N_7854);
nand U7977 (N_7977,N_7758,N_7850);
xnor U7978 (N_7978,N_7783,N_7870);
xor U7979 (N_7979,N_7766,N_7812);
xnor U7980 (N_7980,N_7848,N_7759);
and U7981 (N_7981,N_7842,N_7810);
nand U7982 (N_7982,N_7824,N_7854);
or U7983 (N_7983,N_7809,N_7823);
or U7984 (N_7984,N_7830,N_7834);
and U7985 (N_7985,N_7861,N_7750);
or U7986 (N_7986,N_7792,N_7815);
nor U7987 (N_7987,N_7764,N_7810);
nor U7988 (N_7988,N_7851,N_7860);
nor U7989 (N_7989,N_7853,N_7772);
or U7990 (N_7990,N_7780,N_7750);
and U7991 (N_7991,N_7803,N_7851);
and U7992 (N_7992,N_7846,N_7872);
or U7993 (N_7993,N_7802,N_7871);
or U7994 (N_7994,N_7763,N_7849);
xnor U7995 (N_7995,N_7760,N_7826);
xnor U7996 (N_7996,N_7836,N_7764);
nor U7997 (N_7997,N_7785,N_7853);
and U7998 (N_7998,N_7792,N_7807);
xnor U7999 (N_7999,N_7851,N_7825);
or U8000 (N_8000,N_7971,N_7940);
or U8001 (N_8001,N_7957,N_7888);
or U8002 (N_8002,N_7889,N_7890);
xor U8003 (N_8003,N_7985,N_7961);
nand U8004 (N_8004,N_7952,N_7990);
or U8005 (N_8005,N_7905,N_7877);
xor U8006 (N_8006,N_7886,N_7975);
nand U8007 (N_8007,N_7893,N_7980);
nor U8008 (N_8008,N_7924,N_7934);
or U8009 (N_8009,N_7976,N_7931);
or U8010 (N_8010,N_7919,N_7891);
and U8011 (N_8011,N_7878,N_7963);
and U8012 (N_8012,N_7925,N_7883);
xor U8013 (N_8013,N_7974,N_7935);
nor U8014 (N_8014,N_7977,N_7922);
xor U8015 (N_8015,N_7987,N_7943);
and U8016 (N_8016,N_7950,N_7953);
or U8017 (N_8017,N_7946,N_7984);
or U8018 (N_8018,N_7970,N_7914);
or U8019 (N_8019,N_7875,N_7939);
and U8020 (N_8020,N_7880,N_7923);
or U8021 (N_8021,N_7920,N_7954);
and U8022 (N_8022,N_7962,N_7986);
nor U8023 (N_8023,N_7921,N_7973);
nor U8024 (N_8024,N_7978,N_7892);
nand U8025 (N_8025,N_7960,N_7927);
nor U8026 (N_8026,N_7898,N_7956);
nor U8027 (N_8027,N_7996,N_7979);
or U8028 (N_8028,N_7887,N_7951);
xnor U8029 (N_8029,N_7876,N_7910);
or U8030 (N_8030,N_7897,N_7901);
and U8031 (N_8031,N_7955,N_7879);
or U8032 (N_8032,N_7944,N_7884);
nand U8033 (N_8033,N_7983,N_7967);
or U8034 (N_8034,N_7917,N_7900);
nand U8035 (N_8035,N_7896,N_7928);
or U8036 (N_8036,N_7932,N_7993);
or U8037 (N_8037,N_7912,N_7948);
and U8038 (N_8038,N_7882,N_7949);
nand U8039 (N_8039,N_7969,N_7916);
and U8040 (N_8040,N_7959,N_7908);
nor U8041 (N_8041,N_7894,N_7964);
nor U8042 (N_8042,N_7972,N_7915);
nand U8043 (N_8043,N_7929,N_7913);
or U8044 (N_8044,N_7965,N_7997);
xor U8045 (N_8045,N_7904,N_7999);
or U8046 (N_8046,N_7991,N_7989);
and U8047 (N_8047,N_7994,N_7945);
and U8048 (N_8048,N_7988,N_7906);
or U8049 (N_8049,N_7992,N_7942);
nor U8050 (N_8050,N_7907,N_7938);
or U8051 (N_8051,N_7881,N_7995);
nand U8052 (N_8052,N_7998,N_7911);
and U8053 (N_8053,N_7930,N_7947);
or U8054 (N_8054,N_7903,N_7958);
or U8055 (N_8055,N_7885,N_7941);
or U8056 (N_8056,N_7902,N_7926);
and U8057 (N_8057,N_7968,N_7909);
or U8058 (N_8058,N_7936,N_7895);
or U8059 (N_8059,N_7982,N_7937);
xnor U8060 (N_8060,N_7918,N_7899);
and U8061 (N_8061,N_7933,N_7981);
xor U8062 (N_8062,N_7966,N_7932);
or U8063 (N_8063,N_7957,N_7913);
xnor U8064 (N_8064,N_7944,N_7918);
or U8065 (N_8065,N_7995,N_7965);
or U8066 (N_8066,N_7935,N_7920);
nor U8067 (N_8067,N_7878,N_7956);
nor U8068 (N_8068,N_7875,N_7914);
and U8069 (N_8069,N_7880,N_7981);
nor U8070 (N_8070,N_7918,N_7923);
or U8071 (N_8071,N_7948,N_7937);
xor U8072 (N_8072,N_7923,N_7932);
xnor U8073 (N_8073,N_7994,N_7942);
nand U8074 (N_8074,N_7909,N_7917);
or U8075 (N_8075,N_7901,N_7992);
xor U8076 (N_8076,N_7894,N_7966);
nor U8077 (N_8077,N_7937,N_7893);
or U8078 (N_8078,N_7917,N_7942);
nor U8079 (N_8079,N_7918,N_7963);
or U8080 (N_8080,N_7979,N_7947);
and U8081 (N_8081,N_7905,N_7984);
or U8082 (N_8082,N_7952,N_7981);
or U8083 (N_8083,N_7918,N_7975);
and U8084 (N_8084,N_7963,N_7901);
xnor U8085 (N_8085,N_7942,N_7920);
xnor U8086 (N_8086,N_7904,N_7908);
nand U8087 (N_8087,N_7948,N_7982);
nor U8088 (N_8088,N_7965,N_7945);
or U8089 (N_8089,N_7901,N_7935);
nor U8090 (N_8090,N_7887,N_7893);
xor U8091 (N_8091,N_7988,N_7963);
xnor U8092 (N_8092,N_7912,N_7924);
or U8093 (N_8093,N_7985,N_7905);
and U8094 (N_8094,N_7976,N_7932);
nand U8095 (N_8095,N_7927,N_7969);
nor U8096 (N_8096,N_7991,N_7965);
nor U8097 (N_8097,N_7899,N_7950);
nor U8098 (N_8098,N_7937,N_7876);
xor U8099 (N_8099,N_7884,N_7938);
xor U8100 (N_8100,N_7887,N_7947);
xnor U8101 (N_8101,N_7955,N_7893);
xor U8102 (N_8102,N_7967,N_7966);
nor U8103 (N_8103,N_7983,N_7928);
or U8104 (N_8104,N_7882,N_7902);
xnor U8105 (N_8105,N_7931,N_7985);
nor U8106 (N_8106,N_7927,N_7916);
or U8107 (N_8107,N_7920,N_7915);
nor U8108 (N_8108,N_7977,N_7984);
or U8109 (N_8109,N_7948,N_7876);
xnor U8110 (N_8110,N_7960,N_7980);
or U8111 (N_8111,N_7986,N_7958);
or U8112 (N_8112,N_7948,N_7943);
and U8113 (N_8113,N_7993,N_7905);
and U8114 (N_8114,N_7962,N_7950);
nor U8115 (N_8115,N_7936,N_7910);
xor U8116 (N_8116,N_7896,N_7982);
nand U8117 (N_8117,N_7893,N_7910);
and U8118 (N_8118,N_7995,N_7903);
and U8119 (N_8119,N_7883,N_7892);
or U8120 (N_8120,N_7930,N_7957);
and U8121 (N_8121,N_7886,N_7970);
xnor U8122 (N_8122,N_7946,N_7989);
and U8123 (N_8123,N_7982,N_7892);
xnor U8124 (N_8124,N_7939,N_7918);
nand U8125 (N_8125,N_8083,N_8023);
and U8126 (N_8126,N_8047,N_8091);
nor U8127 (N_8127,N_8019,N_8112);
nand U8128 (N_8128,N_8103,N_8082);
xnor U8129 (N_8129,N_8110,N_8105);
and U8130 (N_8130,N_8068,N_8115);
and U8131 (N_8131,N_8093,N_8101);
nor U8132 (N_8132,N_8048,N_8069);
nand U8133 (N_8133,N_8123,N_8099);
or U8134 (N_8134,N_8114,N_8071);
or U8135 (N_8135,N_8109,N_8086);
nor U8136 (N_8136,N_8122,N_8061);
xnor U8137 (N_8137,N_8058,N_8029);
or U8138 (N_8138,N_8098,N_8003);
and U8139 (N_8139,N_8117,N_8001);
nor U8140 (N_8140,N_8016,N_8056);
nand U8141 (N_8141,N_8054,N_8040);
or U8142 (N_8142,N_8038,N_8006);
nand U8143 (N_8143,N_8096,N_8090);
nand U8144 (N_8144,N_8067,N_8092);
or U8145 (N_8145,N_8076,N_8064);
and U8146 (N_8146,N_8031,N_8066);
and U8147 (N_8147,N_8059,N_8020);
xnor U8148 (N_8148,N_8012,N_8104);
and U8149 (N_8149,N_8044,N_8004);
nor U8150 (N_8150,N_8081,N_8107);
or U8151 (N_8151,N_8008,N_8011);
xnor U8152 (N_8152,N_8022,N_8030);
nor U8153 (N_8153,N_8032,N_8050);
nand U8154 (N_8154,N_8052,N_8106);
nand U8155 (N_8155,N_8095,N_8049);
and U8156 (N_8156,N_8010,N_8055);
or U8157 (N_8157,N_8014,N_8021);
nor U8158 (N_8158,N_8035,N_8041);
nand U8159 (N_8159,N_8039,N_8024);
nor U8160 (N_8160,N_8113,N_8088);
nand U8161 (N_8161,N_8034,N_8043);
nand U8162 (N_8162,N_8042,N_8025);
xor U8163 (N_8163,N_8057,N_8120);
nor U8164 (N_8164,N_8062,N_8051);
or U8165 (N_8165,N_8036,N_8075);
or U8166 (N_8166,N_8074,N_8037);
nor U8167 (N_8167,N_8085,N_8002);
nand U8168 (N_8168,N_8028,N_8063);
nand U8169 (N_8169,N_8026,N_8046);
xor U8170 (N_8170,N_8015,N_8000);
and U8171 (N_8171,N_8027,N_8013);
and U8172 (N_8172,N_8060,N_8072);
or U8173 (N_8173,N_8077,N_8073);
xnor U8174 (N_8174,N_8087,N_8009);
nand U8175 (N_8175,N_8111,N_8080);
nand U8176 (N_8176,N_8116,N_8053);
nor U8177 (N_8177,N_8033,N_8102);
and U8178 (N_8178,N_8018,N_8094);
or U8179 (N_8179,N_8108,N_8045);
or U8180 (N_8180,N_8079,N_8089);
xnor U8181 (N_8181,N_8005,N_8070);
or U8182 (N_8182,N_8065,N_8084);
xnor U8183 (N_8183,N_8007,N_8119);
xnor U8184 (N_8184,N_8100,N_8017);
nand U8185 (N_8185,N_8118,N_8097);
nor U8186 (N_8186,N_8078,N_8124);
and U8187 (N_8187,N_8121,N_8042);
and U8188 (N_8188,N_8120,N_8030);
and U8189 (N_8189,N_8025,N_8047);
and U8190 (N_8190,N_8090,N_8044);
xor U8191 (N_8191,N_8094,N_8036);
or U8192 (N_8192,N_8118,N_8020);
and U8193 (N_8193,N_8121,N_8045);
xnor U8194 (N_8194,N_8074,N_8086);
nand U8195 (N_8195,N_8094,N_8042);
and U8196 (N_8196,N_8051,N_8084);
or U8197 (N_8197,N_8035,N_8029);
xor U8198 (N_8198,N_8024,N_8081);
nor U8199 (N_8199,N_8039,N_8123);
xnor U8200 (N_8200,N_8086,N_8082);
nand U8201 (N_8201,N_8082,N_8070);
xnor U8202 (N_8202,N_8063,N_8038);
nor U8203 (N_8203,N_8119,N_8041);
or U8204 (N_8204,N_8105,N_8031);
and U8205 (N_8205,N_8094,N_8038);
xnor U8206 (N_8206,N_8066,N_8045);
nor U8207 (N_8207,N_8092,N_8099);
xnor U8208 (N_8208,N_8104,N_8029);
nand U8209 (N_8209,N_8058,N_8009);
and U8210 (N_8210,N_8107,N_8049);
nor U8211 (N_8211,N_8079,N_8036);
xor U8212 (N_8212,N_8091,N_8024);
nor U8213 (N_8213,N_8071,N_8027);
and U8214 (N_8214,N_8038,N_8060);
nor U8215 (N_8215,N_8000,N_8029);
and U8216 (N_8216,N_8005,N_8020);
and U8217 (N_8217,N_8014,N_8031);
or U8218 (N_8218,N_8084,N_8018);
xor U8219 (N_8219,N_8048,N_8014);
nor U8220 (N_8220,N_8056,N_8015);
xnor U8221 (N_8221,N_8000,N_8083);
nor U8222 (N_8222,N_8003,N_8036);
or U8223 (N_8223,N_8011,N_8023);
nor U8224 (N_8224,N_8009,N_8044);
nor U8225 (N_8225,N_8053,N_8039);
and U8226 (N_8226,N_8080,N_8061);
nor U8227 (N_8227,N_8006,N_8055);
or U8228 (N_8228,N_8080,N_8008);
nor U8229 (N_8229,N_8001,N_8057);
xnor U8230 (N_8230,N_8092,N_8051);
nand U8231 (N_8231,N_8081,N_8105);
or U8232 (N_8232,N_8109,N_8003);
or U8233 (N_8233,N_8022,N_8071);
nand U8234 (N_8234,N_8109,N_8093);
or U8235 (N_8235,N_8055,N_8002);
nor U8236 (N_8236,N_8038,N_8050);
or U8237 (N_8237,N_8098,N_8010);
nand U8238 (N_8238,N_8103,N_8018);
and U8239 (N_8239,N_8100,N_8055);
xor U8240 (N_8240,N_8060,N_8031);
nand U8241 (N_8241,N_8076,N_8062);
xnor U8242 (N_8242,N_8078,N_8002);
nor U8243 (N_8243,N_8094,N_8035);
nand U8244 (N_8244,N_8089,N_8016);
xor U8245 (N_8245,N_8053,N_8007);
or U8246 (N_8246,N_8024,N_8071);
xnor U8247 (N_8247,N_8003,N_8051);
xor U8248 (N_8248,N_8011,N_8120);
nand U8249 (N_8249,N_8088,N_8098);
or U8250 (N_8250,N_8140,N_8172);
and U8251 (N_8251,N_8233,N_8149);
xnor U8252 (N_8252,N_8143,N_8185);
or U8253 (N_8253,N_8153,N_8151);
nor U8254 (N_8254,N_8175,N_8199);
nor U8255 (N_8255,N_8194,N_8207);
nor U8256 (N_8256,N_8126,N_8201);
nor U8257 (N_8257,N_8220,N_8202);
and U8258 (N_8258,N_8137,N_8148);
xnor U8259 (N_8259,N_8181,N_8173);
nand U8260 (N_8260,N_8247,N_8241);
or U8261 (N_8261,N_8242,N_8188);
xnor U8262 (N_8262,N_8144,N_8171);
and U8263 (N_8263,N_8179,N_8127);
nor U8264 (N_8264,N_8128,N_8214);
nand U8265 (N_8265,N_8130,N_8204);
nor U8266 (N_8266,N_8203,N_8182);
nand U8267 (N_8267,N_8200,N_8211);
nor U8268 (N_8268,N_8229,N_8145);
xnor U8269 (N_8269,N_8174,N_8166);
xnor U8270 (N_8270,N_8139,N_8212);
nand U8271 (N_8271,N_8168,N_8219);
nor U8272 (N_8272,N_8152,N_8234);
xor U8273 (N_8273,N_8164,N_8158);
or U8274 (N_8274,N_8240,N_8192);
or U8275 (N_8275,N_8176,N_8142);
or U8276 (N_8276,N_8134,N_8210);
nand U8277 (N_8277,N_8184,N_8163);
nand U8278 (N_8278,N_8231,N_8141);
or U8279 (N_8279,N_8235,N_8155);
nand U8280 (N_8280,N_8189,N_8180);
xor U8281 (N_8281,N_8161,N_8165);
and U8282 (N_8282,N_8195,N_8232);
and U8283 (N_8283,N_8169,N_8131);
and U8284 (N_8284,N_8213,N_8226);
or U8285 (N_8285,N_8177,N_8125);
xnor U8286 (N_8286,N_8243,N_8248);
nor U8287 (N_8287,N_8205,N_8225);
xnor U8288 (N_8288,N_8230,N_8190);
or U8289 (N_8289,N_8160,N_8218);
or U8290 (N_8290,N_8147,N_8154);
or U8291 (N_8291,N_8237,N_8156);
nor U8292 (N_8292,N_8150,N_8245);
and U8293 (N_8293,N_8193,N_8206);
nand U8294 (N_8294,N_8157,N_8159);
or U8295 (N_8295,N_8249,N_8170);
nand U8296 (N_8296,N_8167,N_8222);
xnor U8297 (N_8297,N_8196,N_8228);
nor U8298 (N_8298,N_8136,N_8227);
or U8299 (N_8299,N_8244,N_8209);
nor U8300 (N_8300,N_8221,N_8238);
nand U8301 (N_8301,N_8191,N_8187);
nor U8302 (N_8302,N_8236,N_8215);
nand U8303 (N_8303,N_8224,N_8246);
nand U8304 (N_8304,N_8146,N_8135);
nand U8305 (N_8305,N_8129,N_8217);
xnor U8306 (N_8306,N_8183,N_8186);
nor U8307 (N_8307,N_8197,N_8132);
nor U8308 (N_8308,N_8239,N_8162);
xnor U8309 (N_8309,N_8198,N_8216);
xnor U8310 (N_8310,N_8178,N_8133);
or U8311 (N_8311,N_8138,N_8223);
and U8312 (N_8312,N_8208,N_8132);
nand U8313 (N_8313,N_8226,N_8192);
nand U8314 (N_8314,N_8127,N_8213);
or U8315 (N_8315,N_8247,N_8226);
or U8316 (N_8316,N_8203,N_8240);
nor U8317 (N_8317,N_8238,N_8210);
nor U8318 (N_8318,N_8205,N_8153);
or U8319 (N_8319,N_8160,N_8237);
or U8320 (N_8320,N_8243,N_8187);
and U8321 (N_8321,N_8221,N_8207);
nor U8322 (N_8322,N_8155,N_8152);
and U8323 (N_8323,N_8242,N_8234);
xor U8324 (N_8324,N_8190,N_8180);
xor U8325 (N_8325,N_8230,N_8188);
or U8326 (N_8326,N_8126,N_8244);
nor U8327 (N_8327,N_8175,N_8145);
nand U8328 (N_8328,N_8249,N_8141);
nor U8329 (N_8329,N_8142,N_8229);
and U8330 (N_8330,N_8132,N_8127);
nor U8331 (N_8331,N_8204,N_8158);
xnor U8332 (N_8332,N_8140,N_8179);
nand U8333 (N_8333,N_8158,N_8148);
nand U8334 (N_8334,N_8165,N_8227);
nor U8335 (N_8335,N_8126,N_8162);
or U8336 (N_8336,N_8168,N_8249);
or U8337 (N_8337,N_8159,N_8127);
xnor U8338 (N_8338,N_8233,N_8219);
nor U8339 (N_8339,N_8125,N_8139);
nor U8340 (N_8340,N_8150,N_8147);
xnor U8341 (N_8341,N_8168,N_8128);
and U8342 (N_8342,N_8197,N_8187);
nor U8343 (N_8343,N_8133,N_8241);
xor U8344 (N_8344,N_8193,N_8246);
xor U8345 (N_8345,N_8144,N_8235);
nor U8346 (N_8346,N_8192,N_8194);
xnor U8347 (N_8347,N_8157,N_8244);
nand U8348 (N_8348,N_8208,N_8169);
nor U8349 (N_8349,N_8177,N_8167);
nand U8350 (N_8350,N_8174,N_8144);
and U8351 (N_8351,N_8232,N_8137);
nor U8352 (N_8352,N_8140,N_8208);
or U8353 (N_8353,N_8199,N_8167);
or U8354 (N_8354,N_8141,N_8221);
nor U8355 (N_8355,N_8147,N_8226);
and U8356 (N_8356,N_8210,N_8241);
xor U8357 (N_8357,N_8214,N_8178);
or U8358 (N_8358,N_8197,N_8195);
nor U8359 (N_8359,N_8174,N_8164);
nor U8360 (N_8360,N_8239,N_8187);
or U8361 (N_8361,N_8228,N_8215);
or U8362 (N_8362,N_8143,N_8144);
nand U8363 (N_8363,N_8175,N_8179);
nand U8364 (N_8364,N_8190,N_8224);
and U8365 (N_8365,N_8235,N_8245);
and U8366 (N_8366,N_8141,N_8163);
and U8367 (N_8367,N_8132,N_8145);
or U8368 (N_8368,N_8204,N_8238);
nand U8369 (N_8369,N_8132,N_8217);
nand U8370 (N_8370,N_8220,N_8160);
and U8371 (N_8371,N_8182,N_8225);
xor U8372 (N_8372,N_8203,N_8207);
xnor U8373 (N_8373,N_8239,N_8126);
or U8374 (N_8374,N_8152,N_8229);
nor U8375 (N_8375,N_8341,N_8257);
xnor U8376 (N_8376,N_8258,N_8363);
and U8377 (N_8377,N_8350,N_8322);
and U8378 (N_8378,N_8367,N_8282);
xnor U8379 (N_8379,N_8329,N_8332);
nand U8380 (N_8380,N_8266,N_8336);
or U8381 (N_8381,N_8250,N_8356);
xnor U8382 (N_8382,N_8310,N_8278);
or U8383 (N_8383,N_8302,N_8326);
and U8384 (N_8384,N_8254,N_8365);
nor U8385 (N_8385,N_8308,N_8289);
and U8386 (N_8386,N_8304,N_8283);
nor U8387 (N_8387,N_8333,N_8372);
or U8388 (N_8388,N_8316,N_8296);
nand U8389 (N_8389,N_8265,N_8291);
or U8390 (N_8390,N_8277,N_8327);
or U8391 (N_8391,N_8342,N_8255);
or U8392 (N_8392,N_8284,N_8299);
nand U8393 (N_8393,N_8279,N_8267);
nor U8394 (N_8394,N_8294,N_8273);
nor U8395 (N_8395,N_8337,N_8335);
or U8396 (N_8396,N_8295,N_8264);
or U8397 (N_8397,N_8261,N_8251);
nor U8398 (N_8398,N_8370,N_8309);
and U8399 (N_8399,N_8339,N_8290);
or U8400 (N_8400,N_8351,N_8271);
nand U8401 (N_8401,N_8315,N_8312);
xnor U8402 (N_8402,N_8358,N_8260);
nor U8403 (N_8403,N_8253,N_8285);
nand U8404 (N_8404,N_8344,N_8357);
and U8405 (N_8405,N_8287,N_8288);
and U8406 (N_8406,N_8262,N_8325);
xor U8407 (N_8407,N_8355,N_8343);
nand U8408 (N_8408,N_8348,N_8252);
and U8409 (N_8409,N_8330,N_8286);
and U8410 (N_8410,N_8331,N_8259);
nand U8411 (N_8411,N_8318,N_8328);
nand U8412 (N_8412,N_8306,N_8256);
and U8413 (N_8413,N_8307,N_8361);
or U8414 (N_8414,N_8324,N_8298);
or U8415 (N_8415,N_8270,N_8320);
nor U8416 (N_8416,N_8305,N_8269);
nand U8417 (N_8417,N_8281,N_8345);
xnor U8418 (N_8418,N_8300,N_8268);
nor U8419 (N_8419,N_8352,N_8314);
or U8420 (N_8420,N_8275,N_8353);
xnor U8421 (N_8421,N_8369,N_8366);
nor U8422 (N_8422,N_8359,N_8263);
nand U8423 (N_8423,N_8334,N_8274);
nor U8424 (N_8424,N_8371,N_8347);
nor U8425 (N_8425,N_8292,N_8297);
and U8426 (N_8426,N_8349,N_8340);
xor U8427 (N_8427,N_8313,N_8373);
xor U8428 (N_8428,N_8272,N_8293);
or U8429 (N_8429,N_8311,N_8317);
and U8430 (N_8430,N_8276,N_8301);
or U8431 (N_8431,N_8303,N_8280);
nand U8432 (N_8432,N_8346,N_8374);
nor U8433 (N_8433,N_8362,N_8319);
and U8434 (N_8434,N_8338,N_8364);
nor U8435 (N_8435,N_8323,N_8368);
and U8436 (N_8436,N_8354,N_8360);
nand U8437 (N_8437,N_8321,N_8302);
nor U8438 (N_8438,N_8280,N_8349);
nand U8439 (N_8439,N_8327,N_8253);
and U8440 (N_8440,N_8292,N_8302);
or U8441 (N_8441,N_8316,N_8268);
nand U8442 (N_8442,N_8346,N_8258);
nand U8443 (N_8443,N_8259,N_8334);
nor U8444 (N_8444,N_8321,N_8291);
nor U8445 (N_8445,N_8321,N_8284);
xnor U8446 (N_8446,N_8263,N_8274);
and U8447 (N_8447,N_8324,N_8273);
or U8448 (N_8448,N_8253,N_8315);
nand U8449 (N_8449,N_8348,N_8370);
nor U8450 (N_8450,N_8277,N_8372);
nand U8451 (N_8451,N_8253,N_8273);
or U8452 (N_8452,N_8282,N_8252);
xor U8453 (N_8453,N_8350,N_8341);
xnor U8454 (N_8454,N_8262,N_8271);
nor U8455 (N_8455,N_8366,N_8285);
and U8456 (N_8456,N_8280,N_8333);
or U8457 (N_8457,N_8340,N_8365);
or U8458 (N_8458,N_8371,N_8317);
and U8459 (N_8459,N_8347,N_8273);
and U8460 (N_8460,N_8281,N_8295);
and U8461 (N_8461,N_8286,N_8373);
xnor U8462 (N_8462,N_8267,N_8330);
or U8463 (N_8463,N_8371,N_8308);
xnor U8464 (N_8464,N_8359,N_8369);
nor U8465 (N_8465,N_8347,N_8251);
nor U8466 (N_8466,N_8275,N_8304);
and U8467 (N_8467,N_8314,N_8355);
or U8468 (N_8468,N_8271,N_8272);
xor U8469 (N_8469,N_8360,N_8365);
or U8470 (N_8470,N_8294,N_8303);
nor U8471 (N_8471,N_8317,N_8312);
xor U8472 (N_8472,N_8368,N_8298);
and U8473 (N_8473,N_8322,N_8272);
or U8474 (N_8474,N_8303,N_8326);
and U8475 (N_8475,N_8297,N_8349);
and U8476 (N_8476,N_8291,N_8372);
nand U8477 (N_8477,N_8335,N_8332);
nand U8478 (N_8478,N_8365,N_8312);
xor U8479 (N_8479,N_8358,N_8290);
or U8480 (N_8480,N_8309,N_8321);
xor U8481 (N_8481,N_8301,N_8307);
or U8482 (N_8482,N_8309,N_8250);
and U8483 (N_8483,N_8368,N_8276);
nor U8484 (N_8484,N_8320,N_8260);
xnor U8485 (N_8485,N_8313,N_8325);
and U8486 (N_8486,N_8309,N_8264);
xor U8487 (N_8487,N_8364,N_8264);
or U8488 (N_8488,N_8361,N_8357);
and U8489 (N_8489,N_8308,N_8263);
xor U8490 (N_8490,N_8334,N_8284);
or U8491 (N_8491,N_8361,N_8302);
nor U8492 (N_8492,N_8323,N_8336);
nand U8493 (N_8493,N_8250,N_8301);
or U8494 (N_8494,N_8323,N_8310);
nand U8495 (N_8495,N_8252,N_8279);
and U8496 (N_8496,N_8272,N_8350);
nor U8497 (N_8497,N_8345,N_8351);
or U8498 (N_8498,N_8259,N_8369);
nand U8499 (N_8499,N_8294,N_8346);
and U8500 (N_8500,N_8483,N_8485);
xor U8501 (N_8501,N_8466,N_8487);
nor U8502 (N_8502,N_8404,N_8375);
xor U8503 (N_8503,N_8456,N_8478);
or U8504 (N_8504,N_8473,N_8412);
xnor U8505 (N_8505,N_8486,N_8495);
xnor U8506 (N_8506,N_8450,N_8471);
or U8507 (N_8507,N_8419,N_8428);
nand U8508 (N_8508,N_8446,N_8407);
xor U8509 (N_8509,N_8494,N_8457);
xor U8510 (N_8510,N_8401,N_8414);
or U8511 (N_8511,N_8384,N_8426);
xor U8512 (N_8512,N_8399,N_8382);
nand U8513 (N_8513,N_8415,N_8464);
nand U8514 (N_8514,N_8440,N_8441);
nand U8515 (N_8515,N_8387,N_8452);
and U8516 (N_8516,N_8492,N_8493);
nor U8517 (N_8517,N_8472,N_8458);
or U8518 (N_8518,N_8448,N_8439);
and U8519 (N_8519,N_8432,N_8391);
nor U8520 (N_8520,N_8388,N_8497);
or U8521 (N_8521,N_8468,N_8396);
or U8522 (N_8522,N_8376,N_8491);
nor U8523 (N_8523,N_8436,N_8397);
nor U8524 (N_8524,N_8479,N_8475);
xor U8525 (N_8525,N_8444,N_8403);
nand U8526 (N_8526,N_8449,N_8488);
and U8527 (N_8527,N_8380,N_8411);
and U8528 (N_8528,N_8377,N_8476);
xnor U8529 (N_8529,N_8421,N_8386);
or U8530 (N_8530,N_8385,N_8469);
nand U8531 (N_8531,N_8394,N_8484);
or U8532 (N_8532,N_8438,N_8470);
nand U8533 (N_8533,N_8383,N_8445);
or U8534 (N_8534,N_8465,N_8418);
or U8535 (N_8535,N_8395,N_8462);
and U8536 (N_8536,N_8453,N_8477);
nor U8537 (N_8537,N_8463,N_8454);
xor U8538 (N_8538,N_8442,N_8451);
xor U8539 (N_8539,N_8437,N_8480);
xor U8540 (N_8540,N_8474,N_8410);
xor U8541 (N_8541,N_8467,N_8400);
and U8542 (N_8542,N_8379,N_8489);
and U8543 (N_8543,N_8461,N_8378);
nor U8544 (N_8544,N_8424,N_8429);
xor U8545 (N_8545,N_8430,N_8433);
and U8546 (N_8546,N_8406,N_8425);
nand U8547 (N_8547,N_8498,N_8393);
nand U8548 (N_8548,N_8405,N_8402);
or U8549 (N_8549,N_8408,N_8417);
or U8550 (N_8550,N_8427,N_8496);
nor U8551 (N_8551,N_8460,N_8434);
and U8552 (N_8552,N_8435,N_8459);
xor U8553 (N_8553,N_8431,N_8389);
and U8554 (N_8554,N_8499,N_8413);
xnor U8555 (N_8555,N_8420,N_8481);
or U8556 (N_8556,N_8392,N_8443);
nor U8557 (N_8557,N_8381,N_8482);
or U8558 (N_8558,N_8455,N_8398);
nor U8559 (N_8559,N_8416,N_8423);
xnor U8560 (N_8560,N_8390,N_8422);
xor U8561 (N_8561,N_8409,N_8490);
nor U8562 (N_8562,N_8447,N_8434);
or U8563 (N_8563,N_8384,N_8438);
and U8564 (N_8564,N_8474,N_8421);
xnor U8565 (N_8565,N_8382,N_8494);
and U8566 (N_8566,N_8442,N_8495);
xor U8567 (N_8567,N_8382,N_8461);
nand U8568 (N_8568,N_8420,N_8462);
nor U8569 (N_8569,N_8402,N_8492);
nand U8570 (N_8570,N_8375,N_8402);
and U8571 (N_8571,N_8489,N_8407);
nand U8572 (N_8572,N_8416,N_8484);
or U8573 (N_8573,N_8381,N_8487);
or U8574 (N_8574,N_8391,N_8415);
nand U8575 (N_8575,N_8474,N_8494);
and U8576 (N_8576,N_8484,N_8435);
nor U8577 (N_8577,N_8383,N_8390);
or U8578 (N_8578,N_8403,N_8455);
nor U8579 (N_8579,N_8493,N_8479);
nor U8580 (N_8580,N_8480,N_8495);
nand U8581 (N_8581,N_8441,N_8480);
nand U8582 (N_8582,N_8412,N_8456);
xnor U8583 (N_8583,N_8418,N_8397);
nor U8584 (N_8584,N_8401,N_8400);
xnor U8585 (N_8585,N_8472,N_8399);
xor U8586 (N_8586,N_8444,N_8498);
nor U8587 (N_8587,N_8422,N_8378);
nand U8588 (N_8588,N_8436,N_8384);
or U8589 (N_8589,N_8388,N_8487);
and U8590 (N_8590,N_8392,N_8459);
xor U8591 (N_8591,N_8446,N_8492);
nor U8592 (N_8592,N_8468,N_8495);
or U8593 (N_8593,N_8489,N_8482);
or U8594 (N_8594,N_8396,N_8487);
nand U8595 (N_8595,N_8453,N_8420);
or U8596 (N_8596,N_8381,N_8470);
or U8597 (N_8597,N_8377,N_8435);
nor U8598 (N_8598,N_8439,N_8499);
and U8599 (N_8599,N_8460,N_8464);
and U8600 (N_8600,N_8496,N_8432);
xor U8601 (N_8601,N_8453,N_8464);
and U8602 (N_8602,N_8471,N_8452);
and U8603 (N_8603,N_8472,N_8465);
nand U8604 (N_8604,N_8481,N_8452);
xnor U8605 (N_8605,N_8452,N_8389);
nor U8606 (N_8606,N_8453,N_8411);
or U8607 (N_8607,N_8433,N_8438);
xnor U8608 (N_8608,N_8379,N_8380);
and U8609 (N_8609,N_8482,N_8396);
or U8610 (N_8610,N_8451,N_8433);
and U8611 (N_8611,N_8481,N_8436);
nor U8612 (N_8612,N_8413,N_8463);
nand U8613 (N_8613,N_8412,N_8431);
xnor U8614 (N_8614,N_8399,N_8418);
or U8615 (N_8615,N_8385,N_8436);
nor U8616 (N_8616,N_8404,N_8460);
and U8617 (N_8617,N_8464,N_8410);
and U8618 (N_8618,N_8434,N_8410);
xor U8619 (N_8619,N_8412,N_8435);
or U8620 (N_8620,N_8432,N_8456);
nand U8621 (N_8621,N_8473,N_8420);
and U8622 (N_8622,N_8488,N_8409);
or U8623 (N_8623,N_8473,N_8476);
or U8624 (N_8624,N_8488,N_8438);
xor U8625 (N_8625,N_8611,N_8620);
xor U8626 (N_8626,N_8578,N_8566);
and U8627 (N_8627,N_8622,N_8623);
nor U8628 (N_8628,N_8605,N_8568);
and U8629 (N_8629,N_8521,N_8522);
or U8630 (N_8630,N_8594,N_8505);
nor U8631 (N_8631,N_8576,N_8559);
or U8632 (N_8632,N_8532,N_8581);
or U8633 (N_8633,N_8603,N_8555);
nand U8634 (N_8634,N_8527,N_8590);
or U8635 (N_8635,N_8525,N_8604);
nor U8636 (N_8636,N_8552,N_8530);
or U8637 (N_8637,N_8565,N_8528);
xor U8638 (N_8638,N_8523,N_8613);
nor U8639 (N_8639,N_8567,N_8610);
and U8640 (N_8640,N_8538,N_8501);
nand U8641 (N_8641,N_8608,N_8540);
xnor U8642 (N_8642,N_8517,N_8511);
nor U8643 (N_8643,N_8516,N_8615);
and U8644 (N_8644,N_8507,N_8616);
and U8645 (N_8645,N_8564,N_8529);
nand U8646 (N_8646,N_8512,N_8543);
and U8647 (N_8647,N_8575,N_8600);
nand U8648 (N_8648,N_8602,N_8574);
nor U8649 (N_8649,N_8520,N_8544);
and U8650 (N_8650,N_8550,N_8504);
xor U8651 (N_8651,N_8515,N_8583);
and U8652 (N_8652,N_8500,N_8618);
xor U8653 (N_8653,N_8535,N_8601);
or U8654 (N_8654,N_8572,N_8526);
nand U8655 (N_8655,N_8617,N_8534);
nor U8656 (N_8656,N_8539,N_8570);
xor U8657 (N_8657,N_8563,N_8533);
xor U8658 (N_8658,N_8619,N_8551);
or U8659 (N_8659,N_8503,N_8524);
or U8660 (N_8660,N_8591,N_8599);
and U8661 (N_8661,N_8585,N_8569);
nor U8662 (N_8662,N_8549,N_8607);
xnor U8663 (N_8663,N_8509,N_8598);
nand U8664 (N_8664,N_8592,N_8545);
or U8665 (N_8665,N_8554,N_8621);
nand U8666 (N_8666,N_8560,N_8614);
xor U8667 (N_8667,N_8537,N_8584);
and U8668 (N_8668,N_8593,N_8573);
and U8669 (N_8669,N_8548,N_8596);
nand U8670 (N_8670,N_8577,N_8519);
and U8671 (N_8671,N_8597,N_8508);
nand U8672 (N_8672,N_8579,N_8609);
nand U8673 (N_8673,N_8606,N_8542);
nor U8674 (N_8674,N_8587,N_8595);
or U8675 (N_8675,N_8571,N_8589);
xnor U8676 (N_8676,N_8506,N_8547);
nor U8677 (N_8677,N_8612,N_8562);
xnor U8678 (N_8678,N_8586,N_8588);
xor U8679 (N_8679,N_8502,N_8510);
and U8680 (N_8680,N_8536,N_8541);
or U8681 (N_8681,N_8556,N_8513);
nand U8682 (N_8682,N_8558,N_8531);
nor U8683 (N_8683,N_8514,N_8624);
nand U8684 (N_8684,N_8582,N_8546);
or U8685 (N_8685,N_8580,N_8561);
or U8686 (N_8686,N_8557,N_8518);
nor U8687 (N_8687,N_8553,N_8615);
xor U8688 (N_8688,N_8579,N_8500);
or U8689 (N_8689,N_8523,N_8594);
nand U8690 (N_8690,N_8605,N_8509);
nor U8691 (N_8691,N_8509,N_8586);
nand U8692 (N_8692,N_8598,N_8550);
nand U8693 (N_8693,N_8611,N_8502);
and U8694 (N_8694,N_8624,N_8538);
nand U8695 (N_8695,N_8572,N_8599);
nand U8696 (N_8696,N_8595,N_8615);
and U8697 (N_8697,N_8518,N_8598);
nor U8698 (N_8698,N_8617,N_8565);
nor U8699 (N_8699,N_8548,N_8509);
or U8700 (N_8700,N_8571,N_8517);
nand U8701 (N_8701,N_8580,N_8551);
or U8702 (N_8702,N_8562,N_8502);
and U8703 (N_8703,N_8577,N_8518);
nand U8704 (N_8704,N_8546,N_8604);
and U8705 (N_8705,N_8564,N_8519);
and U8706 (N_8706,N_8542,N_8539);
nand U8707 (N_8707,N_8528,N_8507);
nand U8708 (N_8708,N_8596,N_8561);
xnor U8709 (N_8709,N_8585,N_8568);
xnor U8710 (N_8710,N_8551,N_8602);
and U8711 (N_8711,N_8510,N_8527);
or U8712 (N_8712,N_8520,N_8531);
or U8713 (N_8713,N_8620,N_8524);
nor U8714 (N_8714,N_8522,N_8569);
or U8715 (N_8715,N_8602,N_8518);
xnor U8716 (N_8716,N_8528,N_8589);
xnor U8717 (N_8717,N_8613,N_8548);
and U8718 (N_8718,N_8524,N_8593);
xor U8719 (N_8719,N_8610,N_8553);
and U8720 (N_8720,N_8528,N_8609);
or U8721 (N_8721,N_8555,N_8504);
or U8722 (N_8722,N_8598,N_8510);
xor U8723 (N_8723,N_8541,N_8617);
xor U8724 (N_8724,N_8622,N_8523);
xor U8725 (N_8725,N_8595,N_8602);
and U8726 (N_8726,N_8613,N_8511);
and U8727 (N_8727,N_8586,N_8571);
xnor U8728 (N_8728,N_8593,N_8622);
and U8729 (N_8729,N_8527,N_8575);
and U8730 (N_8730,N_8597,N_8541);
nand U8731 (N_8731,N_8532,N_8602);
nor U8732 (N_8732,N_8545,N_8538);
xor U8733 (N_8733,N_8516,N_8502);
and U8734 (N_8734,N_8593,N_8570);
xnor U8735 (N_8735,N_8598,N_8566);
xnor U8736 (N_8736,N_8583,N_8512);
xor U8737 (N_8737,N_8604,N_8587);
nand U8738 (N_8738,N_8588,N_8506);
nand U8739 (N_8739,N_8592,N_8624);
xor U8740 (N_8740,N_8507,N_8562);
xnor U8741 (N_8741,N_8614,N_8616);
nor U8742 (N_8742,N_8535,N_8574);
or U8743 (N_8743,N_8561,N_8589);
and U8744 (N_8744,N_8571,N_8557);
xor U8745 (N_8745,N_8606,N_8543);
xnor U8746 (N_8746,N_8513,N_8600);
or U8747 (N_8747,N_8540,N_8514);
xor U8748 (N_8748,N_8605,N_8592);
xor U8749 (N_8749,N_8562,N_8503);
nand U8750 (N_8750,N_8663,N_8657);
nand U8751 (N_8751,N_8668,N_8730);
xor U8752 (N_8752,N_8713,N_8705);
and U8753 (N_8753,N_8729,N_8728);
or U8754 (N_8754,N_8666,N_8688);
xor U8755 (N_8755,N_8731,N_8639);
and U8756 (N_8756,N_8679,N_8716);
nand U8757 (N_8757,N_8693,N_8649);
nor U8758 (N_8758,N_8734,N_8677);
nor U8759 (N_8759,N_8720,N_8640);
xnor U8760 (N_8760,N_8678,N_8667);
nand U8761 (N_8761,N_8721,N_8675);
nor U8762 (N_8762,N_8715,N_8690);
xor U8763 (N_8763,N_8691,N_8632);
xor U8764 (N_8764,N_8655,N_8631);
nor U8765 (N_8765,N_8653,N_8689);
and U8766 (N_8766,N_8749,N_8672);
nand U8767 (N_8767,N_8719,N_8647);
nand U8768 (N_8768,N_8747,N_8627);
nor U8769 (N_8769,N_8664,N_8698);
xnor U8770 (N_8770,N_8744,N_8743);
nor U8771 (N_8771,N_8638,N_8641);
xor U8772 (N_8772,N_8629,N_8685);
nand U8773 (N_8773,N_8634,N_8725);
and U8774 (N_8774,N_8711,N_8651);
or U8775 (N_8775,N_8736,N_8724);
and U8776 (N_8776,N_8656,N_8676);
xor U8777 (N_8777,N_8674,N_8704);
xor U8778 (N_8778,N_8741,N_8712);
nand U8779 (N_8779,N_8694,N_8733);
and U8780 (N_8780,N_8706,N_8660);
and U8781 (N_8781,N_8740,N_8659);
or U8782 (N_8782,N_8646,N_8645);
or U8783 (N_8783,N_8643,N_8686);
or U8784 (N_8784,N_8650,N_8708);
nor U8785 (N_8785,N_8746,N_8642);
and U8786 (N_8786,N_8681,N_8680);
nor U8787 (N_8787,N_8673,N_8709);
or U8788 (N_8788,N_8661,N_8723);
nor U8789 (N_8789,N_8671,N_8737);
xnor U8790 (N_8790,N_8700,N_8669);
or U8791 (N_8791,N_8717,N_8626);
or U8792 (N_8792,N_8637,N_8628);
nand U8793 (N_8793,N_8670,N_8697);
xnor U8794 (N_8794,N_8665,N_8718);
or U8795 (N_8795,N_8710,N_8630);
nand U8796 (N_8796,N_8648,N_8745);
nor U8797 (N_8797,N_8633,N_8625);
and U8798 (N_8798,N_8738,N_8699);
xor U8799 (N_8799,N_8714,N_8707);
and U8800 (N_8800,N_8662,N_8696);
nand U8801 (N_8801,N_8687,N_8636);
nand U8802 (N_8802,N_8695,N_8726);
nor U8803 (N_8803,N_8735,N_8683);
or U8804 (N_8804,N_8732,N_8644);
nor U8805 (N_8805,N_8682,N_8739);
and U8806 (N_8806,N_8635,N_8684);
nand U8807 (N_8807,N_8722,N_8703);
xnor U8808 (N_8808,N_8727,N_8654);
xnor U8809 (N_8809,N_8701,N_8702);
and U8810 (N_8810,N_8652,N_8692);
nand U8811 (N_8811,N_8748,N_8658);
and U8812 (N_8812,N_8742,N_8668);
and U8813 (N_8813,N_8662,N_8640);
xor U8814 (N_8814,N_8723,N_8726);
xnor U8815 (N_8815,N_8637,N_8716);
or U8816 (N_8816,N_8675,N_8723);
nor U8817 (N_8817,N_8652,N_8747);
nand U8818 (N_8818,N_8747,N_8671);
and U8819 (N_8819,N_8675,N_8673);
or U8820 (N_8820,N_8635,N_8650);
xor U8821 (N_8821,N_8683,N_8671);
and U8822 (N_8822,N_8625,N_8630);
nand U8823 (N_8823,N_8667,N_8703);
nand U8824 (N_8824,N_8628,N_8702);
nand U8825 (N_8825,N_8671,N_8630);
and U8826 (N_8826,N_8634,N_8734);
or U8827 (N_8827,N_8683,N_8725);
or U8828 (N_8828,N_8686,N_8664);
or U8829 (N_8829,N_8749,N_8681);
xnor U8830 (N_8830,N_8733,N_8739);
or U8831 (N_8831,N_8734,N_8635);
or U8832 (N_8832,N_8722,N_8705);
nor U8833 (N_8833,N_8701,N_8719);
xor U8834 (N_8834,N_8657,N_8700);
xnor U8835 (N_8835,N_8720,N_8715);
nand U8836 (N_8836,N_8692,N_8690);
or U8837 (N_8837,N_8625,N_8722);
xnor U8838 (N_8838,N_8710,N_8739);
xor U8839 (N_8839,N_8722,N_8666);
or U8840 (N_8840,N_8749,N_8707);
nor U8841 (N_8841,N_8653,N_8644);
xnor U8842 (N_8842,N_8738,N_8639);
xnor U8843 (N_8843,N_8691,N_8668);
and U8844 (N_8844,N_8736,N_8694);
nand U8845 (N_8845,N_8646,N_8676);
nand U8846 (N_8846,N_8746,N_8712);
or U8847 (N_8847,N_8697,N_8673);
and U8848 (N_8848,N_8724,N_8707);
nand U8849 (N_8849,N_8723,N_8646);
xnor U8850 (N_8850,N_8684,N_8641);
or U8851 (N_8851,N_8693,N_8703);
nand U8852 (N_8852,N_8736,N_8722);
or U8853 (N_8853,N_8631,N_8741);
nor U8854 (N_8854,N_8660,N_8736);
and U8855 (N_8855,N_8744,N_8692);
xnor U8856 (N_8856,N_8729,N_8638);
or U8857 (N_8857,N_8630,N_8656);
nor U8858 (N_8858,N_8671,N_8656);
or U8859 (N_8859,N_8700,N_8718);
nor U8860 (N_8860,N_8652,N_8701);
nor U8861 (N_8861,N_8714,N_8734);
xor U8862 (N_8862,N_8676,N_8681);
or U8863 (N_8863,N_8689,N_8748);
nor U8864 (N_8864,N_8666,N_8645);
xnor U8865 (N_8865,N_8732,N_8655);
nand U8866 (N_8866,N_8633,N_8736);
nor U8867 (N_8867,N_8729,N_8725);
xnor U8868 (N_8868,N_8686,N_8711);
nor U8869 (N_8869,N_8696,N_8651);
or U8870 (N_8870,N_8718,N_8725);
and U8871 (N_8871,N_8685,N_8643);
or U8872 (N_8872,N_8664,N_8703);
or U8873 (N_8873,N_8702,N_8667);
nor U8874 (N_8874,N_8664,N_8714);
or U8875 (N_8875,N_8821,N_8811);
and U8876 (N_8876,N_8792,N_8781);
or U8877 (N_8877,N_8776,N_8822);
or U8878 (N_8878,N_8857,N_8853);
or U8879 (N_8879,N_8805,N_8839);
nor U8880 (N_8880,N_8867,N_8830);
nor U8881 (N_8881,N_8856,N_8829);
and U8882 (N_8882,N_8774,N_8778);
or U8883 (N_8883,N_8801,N_8820);
nand U8884 (N_8884,N_8758,N_8837);
and U8885 (N_8885,N_8818,N_8849);
xnor U8886 (N_8886,N_8752,N_8844);
nor U8887 (N_8887,N_8841,N_8824);
and U8888 (N_8888,N_8794,N_8847);
xnor U8889 (N_8889,N_8799,N_8783);
or U8890 (N_8890,N_8751,N_8848);
xnor U8891 (N_8891,N_8814,N_8796);
nor U8892 (N_8892,N_8789,N_8858);
or U8893 (N_8893,N_8800,N_8851);
or U8894 (N_8894,N_8874,N_8835);
xnor U8895 (N_8895,N_8854,N_8803);
and U8896 (N_8896,N_8865,N_8775);
nor U8897 (N_8897,N_8842,N_8834);
nor U8898 (N_8898,N_8793,N_8873);
xnor U8899 (N_8899,N_8838,N_8760);
and U8900 (N_8900,N_8797,N_8755);
or U8901 (N_8901,N_8788,N_8808);
nand U8902 (N_8902,N_8872,N_8761);
xnor U8903 (N_8903,N_8816,N_8852);
or U8904 (N_8904,N_8772,N_8866);
and U8905 (N_8905,N_8862,N_8863);
nand U8906 (N_8906,N_8812,N_8769);
or U8907 (N_8907,N_8777,N_8764);
nor U8908 (N_8908,N_8828,N_8763);
and U8909 (N_8909,N_8871,N_8807);
nand U8910 (N_8910,N_8868,N_8790);
or U8911 (N_8911,N_8750,N_8827);
nand U8912 (N_8912,N_8840,N_8860);
or U8913 (N_8913,N_8766,N_8756);
nor U8914 (N_8914,N_8809,N_8798);
nor U8915 (N_8915,N_8831,N_8757);
nor U8916 (N_8916,N_8759,N_8819);
nor U8917 (N_8917,N_8869,N_8785);
nor U8918 (N_8918,N_8855,N_8791);
xor U8919 (N_8919,N_8833,N_8806);
and U8920 (N_8920,N_8753,N_8817);
xor U8921 (N_8921,N_8845,N_8787);
and U8922 (N_8922,N_8782,N_8795);
xor U8923 (N_8923,N_8836,N_8850);
nor U8924 (N_8924,N_8767,N_8765);
and U8925 (N_8925,N_8825,N_8802);
or U8926 (N_8926,N_8773,N_8846);
or U8927 (N_8927,N_8826,N_8815);
nand U8928 (N_8928,N_8754,N_8770);
xnor U8929 (N_8929,N_8786,N_8771);
xnor U8930 (N_8930,N_8859,N_8762);
nand U8931 (N_8931,N_8810,N_8861);
nand U8932 (N_8932,N_8780,N_8779);
and U8933 (N_8933,N_8870,N_8864);
or U8934 (N_8934,N_8823,N_8784);
or U8935 (N_8935,N_8843,N_8768);
xor U8936 (N_8936,N_8832,N_8804);
nor U8937 (N_8937,N_8813,N_8779);
xnor U8938 (N_8938,N_8820,N_8841);
nand U8939 (N_8939,N_8842,N_8862);
nand U8940 (N_8940,N_8862,N_8774);
nor U8941 (N_8941,N_8774,N_8831);
nor U8942 (N_8942,N_8795,N_8793);
or U8943 (N_8943,N_8814,N_8797);
nand U8944 (N_8944,N_8835,N_8822);
or U8945 (N_8945,N_8797,N_8786);
nor U8946 (N_8946,N_8814,N_8873);
xor U8947 (N_8947,N_8824,N_8872);
nor U8948 (N_8948,N_8846,N_8793);
xor U8949 (N_8949,N_8869,N_8792);
nor U8950 (N_8950,N_8856,N_8803);
nor U8951 (N_8951,N_8775,N_8864);
and U8952 (N_8952,N_8844,N_8861);
nor U8953 (N_8953,N_8854,N_8830);
xor U8954 (N_8954,N_8855,N_8849);
and U8955 (N_8955,N_8856,N_8771);
xnor U8956 (N_8956,N_8833,N_8771);
and U8957 (N_8957,N_8771,N_8826);
xor U8958 (N_8958,N_8794,N_8851);
or U8959 (N_8959,N_8863,N_8787);
nand U8960 (N_8960,N_8867,N_8874);
or U8961 (N_8961,N_8853,N_8874);
or U8962 (N_8962,N_8774,N_8788);
and U8963 (N_8963,N_8862,N_8850);
nand U8964 (N_8964,N_8824,N_8756);
or U8965 (N_8965,N_8847,N_8874);
or U8966 (N_8966,N_8799,N_8838);
nor U8967 (N_8967,N_8844,N_8820);
nand U8968 (N_8968,N_8855,N_8871);
nor U8969 (N_8969,N_8830,N_8801);
nand U8970 (N_8970,N_8810,N_8784);
and U8971 (N_8971,N_8834,N_8825);
and U8972 (N_8972,N_8871,N_8862);
and U8973 (N_8973,N_8754,N_8817);
xor U8974 (N_8974,N_8769,N_8791);
xnor U8975 (N_8975,N_8834,N_8788);
xor U8976 (N_8976,N_8874,N_8862);
nand U8977 (N_8977,N_8753,N_8784);
or U8978 (N_8978,N_8848,N_8802);
and U8979 (N_8979,N_8869,N_8775);
and U8980 (N_8980,N_8847,N_8791);
nand U8981 (N_8981,N_8835,N_8854);
or U8982 (N_8982,N_8834,N_8871);
nand U8983 (N_8983,N_8820,N_8866);
and U8984 (N_8984,N_8806,N_8794);
or U8985 (N_8985,N_8804,N_8769);
nor U8986 (N_8986,N_8847,N_8825);
nor U8987 (N_8987,N_8863,N_8794);
or U8988 (N_8988,N_8791,N_8869);
nand U8989 (N_8989,N_8762,N_8871);
xor U8990 (N_8990,N_8772,N_8789);
nand U8991 (N_8991,N_8859,N_8855);
xor U8992 (N_8992,N_8770,N_8836);
and U8993 (N_8993,N_8850,N_8824);
nand U8994 (N_8994,N_8861,N_8755);
xor U8995 (N_8995,N_8807,N_8842);
nor U8996 (N_8996,N_8815,N_8795);
or U8997 (N_8997,N_8818,N_8752);
nand U8998 (N_8998,N_8773,N_8844);
nor U8999 (N_8999,N_8853,N_8786);
nand U9000 (N_9000,N_8963,N_8959);
or U9001 (N_9001,N_8946,N_8895);
nor U9002 (N_9002,N_8961,N_8953);
nand U9003 (N_9003,N_8880,N_8938);
or U9004 (N_9004,N_8884,N_8913);
nand U9005 (N_9005,N_8893,N_8936);
nor U9006 (N_9006,N_8990,N_8902);
nand U9007 (N_9007,N_8889,N_8878);
nor U9008 (N_9008,N_8972,N_8877);
xnor U9009 (N_9009,N_8999,N_8932);
xor U9010 (N_9010,N_8887,N_8879);
xnor U9011 (N_9011,N_8916,N_8943);
and U9012 (N_9012,N_8928,N_8915);
and U9013 (N_9013,N_8917,N_8919);
or U9014 (N_9014,N_8897,N_8883);
nand U9015 (N_9015,N_8960,N_8992);
nand U9016 (N_9016,N_8996,N_8931);
nor U9017 (N_9017,N_8890,N_8912);
nor U9018 (N_9018,N_8981,N_8950);
and U9019 (N_9019,N_8979,N_8914);
xnor U9020 (N_9020,N_8966,N_8997);
xnor U9021 (N_9021,N_8969,N_8926);
nand U9022 (N_9022,N_8952,N_8982);
nand U9023 (N_9023,N_8930,N_8876);
nand U9024 (N_9024,N_8948,N_8989);
and U9025 (N_9025,N_8885,N_8900);
xor U9026 (N_9026,N_8882,N_8886);
nand U9027 (N_9027,N_8894,N_8904);
nand U9028 (N_9028,N_8905,N_8985);
or U9029 (N_9029,N_8964,N_8922);
nand U9030 (N_9030,N_8994,N_8941);
nand U9031 (N_9031,N_8881,N_8921);
and U9032 (N_9032,N_8958,N_8891);
nand U9033 (N_9033,N_8973,N_8975);
nand U9034 (N_9034,N_8906,N_8937);
xor U9035 (N_9035,N_8899,N_8910);
nor U9036 (N_9036,N_8933,N_8934);
and U9037 (N_9037,N_8984,N_8911);
nor U9038 (N_9038,N_8924,N_8896);
xor U9039 (N_9039,N_8986,N_8955);
nor U9040 (N_9040,N_8927,N_8968);
nor U9041 (N_9041,N_8908,N_8998);
and U9042 (N_9042,N_8976,N_8920);
and U9043 (N_9043,N_8962,N_8903);
nand U9044 (N_9044,N_8888,N_8940);
and U9045 (N_9045,N_8951,N_8957);
or U9046 (N_9046,N_8970,N_8991);
nand U9047 (N_9047,N_8978,N_8918);
xnor U9048 (N_9048,N_8944,N_8987);
or U9049 (N_9049,N_8935,N_8892);
nand U9050 (N_9050,N_8898,N_8980);
xnor U9051 (N_9051,N_8909,N_8988);
and U9052 (N_9052,N_8923,N_8949);
xor U9053 (N_9053,N_8947,N_8907);
and U9054 (N_9054,N_8956,N_8971);
nor U9055 (N_9055,N_8945,N_8965);
nor U9056 (N_9056,N_8995,N_8942);
nor U9057 (N_9057,N_8993,N_8901);
and U9058 (N_9058,N_8983,N_8967);
nand U9059 (N_9059,N_8875,N_8929);
or U9060 (N_9060,N_8974,N_8925);
nor U9061 (N_9061,N_8977,N_8939);
and U9062 (N_9062,N_8954,N_8937);
nand U9063 (N_9063,N_8882,N_8960);
or U9064 (N_9064,N_8900,N_8950);
xor U9065 (N_9065,N_8938,N_8883);
nand U9066 (N_9066,N_8975,N_8900);
or U9067 (N_9067,N_8921,N_8943);
or U9068 (N_9068,N_8923,N_8973);
nor U9069 (N_9069,N_8995,N_8965);
nor U9070 (N_9070,N_8958,N_8993);
or U9071 (N_9071,N_8955,N_8992);
or U9072 (N_9072,N_8935,N_8876);
nor U9073 (N_9073,N_8936,N_8999);
and U9074 (N_9074,N_8921,N_8937);
or U9075 (N_9075,N_8954,N_8931);
nand U9076 (N_9076,N_8887,N_8949);
xor U9077 (N_9077,N_8929,N_8905);
nand U9078 (N_9078,N_8921,N_8883);
nor U9079 (N_9079,N_8993,N_8977);
xor U9080 (N_9080,N_8907,N_8951);
and U9081 (N_9081,N_8879,N_8892);
and U9082 (N_9082,N_8957,N_8959);
or U9083 (N_9083,N_8907,N_8876);
xnor U9084 (N_9084,N_8941,N_8921);
and U9085 (N_9085,N_8944,N_8909);
or U9086 (N_9086,N_8990,N_8875);
or U9087 (N_9087,N_8920,N_8898);
nor U9088 (N_9088,N_8886,N_8897);
nor U9089 (N_9089,N_8947,N_8882);
xnor U9090 (N_9090,N_8997,N_8964);
or U9091 (N_9091,N_8892,N_8889);
nand U9092 (N_9092,N_8981,N_8897);
nor U9093 (N_9093,N_8905,N_8901);
nor U9094 (N_9094,N_8890,N_8935);
xor U9095 (N_9095,N_8997,N_8884);
or U9096 (N_9096,N_8910,N_8942);
xor U9097 (N_9097,N_8935,N_8878);
nor U9098 (N_9098,N_8922,N_8949);
or U9099 (N_9099,N_8956,N_8949);
nand U9100 (N_9100,N_8886,N_8934);
or U9101 (N_9101,N_8950,N_8956);
and U9102 (N_9102,N_8968,N_8889);
nor U9103 (N_9103,N_8970,N_8883);
nor U9104 (N_9104,N_8975,N_8977);
and U9105 (N_9105,N_8912,N_8940);
and U9106 (N_9106,N_8987,N_8887);
or U9107 (N_9107,N_8877,N_8905);
or U9108 (N_9108,N_8909,N_8991);
nor U9109 (N_9109,N_8974,N_8932);
nor U9110 (N_9110,N_8974,N_8875);
nor U9111 (N_9111,N_8970,N_8905);
and U9112 (N_9112,N_8993,N_8944);
nor U9113 (N_9113,N_8916,N_8929);
and U9114 (N_9114,N_8912,N_8969);
or U9115 (N_9115,N_8993,N_8999);
nor U9116 (N_9116,N_8914,N_8995);
xnor U9117 (N_9117,N_8935,N_8928);
nor U9118 (N_9118,N_8897,N_8960);
xnor U9119 (N_9119,N_8903,N_8981);
or U9120 (N_9120,N_8887,N_8977);
nand U9121 (N_9121,N_8893,N_8978);
or U9122 (N_9122,N_8942,N_8962);
or U9123 (N_9123,N_8969,N_8941);
xnor U9124 (N_9124,N_8919,N_8986);
and U9125 (N_9125,N_9059,N_9103);
nor U9126 (N_9126,N_9069,N_9044);
xnor U9127 (N_9127,N_9090,N_9082);
nor U9128 (N_9128,N_9064,N_9047);
or U9129 (N_9129,N_9094,N_9107);
or U9130 (N_9130,N_9115,N_9052);
nand U9131 (N_9131,N_9017,N_9116);
xnor U9132 (N_9132,N_9109,N_9053);
or U9133 (N_9133,N_9058,N_9014);
and U9134 (N_9134,N_9086,N_9001);
nor U9135 (N_9135,N_9009,N_9095);
nor U9136 (N_9136,N_9026,N_9111);
nor U9137 (N_9137,N_9114,N_9029);
nand U9138 (N_9138,N_9070,N_9106);
nor U9139 (N_9139,N_9006,N_9034);
nor U9140 (N_9140,N_9101,N_9057);
nor U9141 (N_9141,N_9062,N_9011);
xnor U9142 (N_9142,N_9007,N_9110);
nor U9143 (N_9143,N_9113,N_9022);
nor U9144 (N_9144,N_9043,N_9093);
and U9145 (N_9145,N_9077,N_9063);
nor U9146 (N_9146,N_9048,N_9019);
nor U9147 (N_9147,N_9087,N_9039);
xnor U9148 (N_9148,N_9102,N_9075);
xor U9149 (N_9149,N_9050,N_9012);
or U9150 (N_9150,N_9124,N_9054);
nor U9151 (N_9151,N_9003,N_9040);
and U9152 (N_9152,N_9088,N_9038);
and U9153 (N_9153,N_9083,N_9021);
nand U9154 (N_9154,N_9112,N_9060);
nor U9155 (N_9155,N_9018,N_9035);
and U9156 (N_9156,N_9032,N_9020);
and U9157 (N_9157,N_9123,N_9068);
nor U9158 (N_9158,N_9084,N_9016);
nor U9159 (N_9159,N_9000,N_9120);
nor U9160 (N_9160,N_9097,N_9091);
nand U9161 (N_9161,N_9061,N_9010);
xnor U9162 (N_9162,N_9072,N_9051);
xnor U9163 (N_9163,N_9108,N_9081);
nor U9164 (N_9164,N_9078,N_9027);
nand U9165 (N_9165,N_9079,N_9045);
xor U9166 (N_9166,N_9067,N_9030);
and U9167 (N_9167,N_9002,N_9037);
nor U9168 (N_9168,N_9031,N_9066);
xnor U9169 (N_9169,N_9105,N_9046);
and U9170 (N_9170,N_9004,N_9042);
nand U9171 (N_9171,N_9121,N_9033);
nand U9172 (N_9172,N_9118,N_9049);
and U9173 (N_9173,N_9104,N_9025);
nor U9174 (N_9174,N_9117,N_9008);
xnor U9175 (N_9175,N_9085,N_9074);
nand U9176 (N_9176,N_9089,N_9122);
nand U9177 (N_9177,N_9024,N_9073);
nor U9178 (N_9178,N_9092,N_9071);
nor U9179 (N_9179,N_9099,N_9080);
nand U9180 (N_9180,N_9023,N_9119);
nand U9181 (N_9181,N_9098,N_9015);
and U9182 (N_9182,N_9028,N_9065);
nor U9183 (N_9183,N_9005,N_9100);
nand U9184 (N_9184,N_9036,N_9013);
or U9185 (N_9185,N_9076,N_9041);
and U9186 (N_9186,N_9096,N_9056);
and U9187 (N_9187,N_9055,N_9078);
nor U9188 (N_9188,N_9014,N_9000);
or U9189 (N_9189,N_9061,N_9072);
and U9190 (N_9190,N_9087,N_9052);
nand U9191 (N_9191,N_9113,N_9063);
and U9192 (N_9192,N_9000,N_9082);
nand U9193 (N_9193,N_9032,N_9035);
nand U9194 (N_9194,N_9076,N_9090);
nand U9195 (N_9195,N_9023,N_9084);
nand U9196 (N_9196,N_9039,N_9001);
nor U9197 (N_9197,N_9109,N_9035);
xnor U9198 (N_9198,N_9099,N_9045);
xor U9199 (N_9199,N_9065,N_9021);
xor U9200 (N_9200,N_9056,N_9106);
nor U9201 (N_9201,N_9038,N_9121);
xnor U9202 (N_9202,N_9000,N_9107);
xor U9203 (N_9203,N_9054,N_9115);
or U9204 (N_9204,N_9049,N_9087);
and U9205 (N_9205,N_9035,N_9042);
nor U9206 (N_9206,N_9087,N_9095);
and U9207 (N_9207,N_9111,N_9000);
or U9208 (N_9208,N_9046,N_9056);
nand U9209 (N_9209,N_9076,N_9013);
xor U9210 (N_9210,N_9074,N_9022);
nand U9211 (N_9211,N_9047,N_9118);
nand U9212 (N_9212,N_9100,N_9103);
xnor U9213 (N_9213,N_9003,N_9013);
or U9214 (N_9214,N_9036,N_9046);
or U9215 (N_9215,N_9114,N_9000);
nor U9216 (N_9216,N_9124,N_9001);
nand U9217 (N_9217,N_9092,N_9016);
xnor U9218 (N_9218,N_9104,N_9083);
nand U9219 (N_9219,N_9054,N_9003);
nand U9220 (N_9220,N_9067,N_9116);
and U9221 (N_9221,N_9058,N_9051);
xnor U9222 (N_9222,N_9052,N_9041);
nand U9223 (N_9223,N_9004,N_9072);
and U9224 (N_9224,N_9114,N_9119);
and U9225 (N_9225,N_9121,N_9042);
nor U9226 (N_9226,N_9005,N_9068);
nand U9227 (N_9227,N_9071,N_9051);
or U9228 (N_9228,N_9075,N_9097);
and U9229 (N_9229,N_9061,N_9048);
nor U9230 (N_9230,N_9012,N_9011);
nand U9231 (N_9231,N_9105,N_9118);
and U9232 (N_9232,N_9031,N_9113);
nand U9233 (N_9233,N_9053,N_9006);
xnor U9234 (N_9234,N_9014,N_9072);
xnor U9235 (N_9235,N_9007,N_9061);
xor U9236 (N_9236,N_9058,N_9119);
nor U9237 (N_9237,N_9013,N_9115);
and U9238 (N_9238,N_9033,N_9027);
nand U9239 (N_9239,N_9053,N_9052);
nand U9240 (N_9240,N_9116,N_9091);
xor U9241 (N_9241,N_9063,N_9050);
nand U9242 (N_9242,N_9051,N_9108);
and U9243 (N_9243,N_9123,N_9030);
nand U9244 (N_9244,N_9102,N_9040);
and U9245 (N_9245,N_9011,N_9093);
nor U9246 (N_9246,N_9071,N_9005);
and U9247 (N_9247,N_9037,N_9031);
or U9248 (N_9248,N_9109,N_9111);
or U9249 (N_9249,N_9011,N_9104);
and U9250 (N_9250,N_9168,N_9219);
nor U9251 (N_9251,N_9195,N_9194);
and U9252 (N_9252,N_9203,N_9222);
nor U9253 (N_9253,N_9190,N_9186);
nor U9254 (N_9254,N_9246,N_9140);
and U9255 (N_9255,N_9125,N_9237);
xnor U9256 (N_9256,N_9242,N_9126);
and U9257 (N_9257,N_9175,N_9236);
nand U9258 (N_9258,N_9165,N_9234);
and U9259 (N_9259,N_9249,N_9241);
nand U9260 (N_9260,N_9180,N_9135);
nand U9261 (N_9261,N_9208,N_9161);
and U9262 (N_9262,N_9159,N_9215);
and U9263 (N_9263,N_9132,N_9164);
nand U9264 (N_9264,N_9224,N_9130);
and U9265 (N_9265,N_9151,N_9197);
nor U9266 (N_9266,N_9204,N_9171);
nor U9267 (N_9267,N_9213,N_9177);
and U9268 (N_9268,N_9225,N_9192);
or U9269 (N_9269,N_9143,N_9247);
and U9270 (N_9270,N_9205,N_9214);
nor U9271 (N_9271,N_9139,N_9157);
nand U9272 (N_9272,N_9131,N_9221);
and U9273 (N_9273,N_9141,N_9212);
and U9274 (N_9274,N_9240,N_9137);
nand U9275 (N_9275,N_9207,N_9245);
xnor U9276 (N_9276,N_9156,N_9149);
xor U9277 (N_9277,N_9223,N_9146);
and U9278 (N_9278,N_9170,N_9231);
and U9279 (N_9279,N_9174,N_9178);
nor U9280 (N_9280,N_9142,N_9188);
nand U9281 (N_9281,N_9152,N_9248);
or U9282 (N_9282,N_9172,N_9233);
nor U9283 (N_9283,N_9162,N_9179);
nor U9284 (N_9284,N_9182,N_9227);
xnor U9285 (N_9285,N_9138,N_9232);
nor U9286 (N_9286,N_9211,N_9201);
and U9287 (N_9287,N_9153,N_9155);
nand U9288 (N_9288,N_9191,N_9166);
and U9289 (N_9289,N_9216,N_9193);
or U9290 (N_9290,N_9200,N_9176);
nand U9291 (N_9291,N_9187,N_9169);
nand U9292 (N_9292,N_9198,N_9145);
nand U9293 (N_9293,N_9229,N_9217);
xnor U9294 (N_9294,N_9209,N_9150);
and U9295 (N_9295,N_9154,N_9185);
nor U9296 (N_9296,N_9230,N_9220);
nand U9297 (N_9297,N_9158,N_9238);
nor U9298 (N_9298,N_9181,N_9167);
xor U9299 (N_9299,N_9235,N_9163);
nor U9300 (N_9300,N_9189,N_9160);
nand U9301 (N_9301,N_9228,N_9218);
or U9302 (N_9302,N_9144,N_9210);
nor U9303 (N_9303,N_9239,N_9243);
or U9304 (N_9304,N_9202,N_9147);
xor U9305 (N_9305,N_9226,N_9199);
nand U9306 (N_9306,N_9196,N_9136);
xnor U9307 (N_9307,N_9129,N_9127);
and U9308 (N_9308,N_9148,N_9134);
nand U9309 (N_9309,N_9128,N_9173);
nor U9310 (N_9310,N_9183,N_9206);
or U9311 (N_9311,N_9184,N_9244);
nor U9312 (N_9312,N_9133,N_9168);
and U9313 (N_9313,N_9136,N_9228);
or U9314 (N_9314,N_9185,N_9125);
or U9315 (N_9315,N_9180,N_9208);
and U9316 (N_9316,N_9137,N_9158);
and U9317 (N_9317,N_9221,N_9152);
xor U9318 (N_9318,N_9226,N_9129);
nand U9319 (N_9319,N_9181,N_9212);
nand U9320 (N_9320,N_9159,N_9232);
nand U9321 (N_9321,N_9167,N_9136);
nand U9322 (N_9322,N_9207,N_9239);
nand U9323 (N_9323,N_9180,N_9217);
nand U9324 (N_9324,N_9146,N_9186);
xor U9325 (N_9325,N_9180,N_9235);
and U9326 (N_9326,N_9217,N_9134);
or U9327 (N_9327,N_9183,N_9145);
and U9328 (N_9328,N_9216,N_9202);
and U9329 (N_9329,N_9191,N_9141);
and U9330 (N_9330,N_9236,N_9171);
or U9331 (N_9331,N_9235,N_9134);
nor U9332 (N_9332,N_9151,N_9162);
nand U9333 (N_9333,N_9163,N_9148);
nand U9334 (N_9334,N_9215,N_9168);
nand U9335 (N_9335,N_9151,N_9205);
or U9336 (N_9336,N_9226,N_9245);
xor U9337 (N_9337,N_9190,N_9173);
nand U9338 (N_9338,N_9140,N_9202);
or U9339 (N_9339,N_9165,N_9224);
xnor U9340 (N_9340,N_9231,N_9161);
nor U9341 (N_9341,N_9125,N_9148);
nand U9342 (N_9342,N_9184,N_9182);
xor U9343 (N_9343,N_9127,N_9193);
and U9344 (N_9344,N_9146,N_9211);
xnor U9345 (N_9345,N_9195,N_9200);
or U9346 (N_9346,N_9201,N_9174);
or U9347 (N_9347,N_9178,N_9141);
nor U9348 (N_9348,N_9132,N_9134);
nor U9349 (N_9349,N_9211,N_9247);
and U9350 (N_9350,N_9125,N_9149);
xnor U9351 (N_9351,N_9175,N_9204);
or U9352 (N_9352,N_9151,N_9166);
xor U9353 (N_9353,N_9173,N_9242);
xnor U9354 (N_9354,N_9200,N_9127);
nor U9355 (N_9355,N_9225,N_9241);
nor U9356 (N_9356,N_9206,N_9130);
or U9357 (N_9357,N_9140,N_9158);
nor U9358 (N_9358,N_9227,N_9134);
and U9359 (N_9359,N_9244,N_9180);
and U9360 (N_9360,N_9155,N_9227);
xnor U9361 (N_9361,N_9198,N_9179);
and U9362 (N_9362,N_9130,N_9214);
and U9363 (N_9363,N_9180,N_9238);
nor U9364 (N_9364,N_9224,N_9245);
or U9365 (N_9365,N_9184,N_9157);
nor U9366 (N_9366,N_9197,N_9168);
xnor U9367 (N_9367,N_9245,N_9185);
nor U9368 (N_9368,N_9219,N_9146);
and U9369 (N_9369,N_9140,N_9223);
or U9370 (N_9370,N_9237,N_9198);
and U9371 (N_9371,N_9209,N_9149);
nor U9372 (N_9372,N_9194,N_9221);
or U9373 (N_9373,N_9140,N_9167);
or U9374 (N_9374,N_9243,N_9238);
xor U9375 (N_9375,N_9255,N_9278);
nor U9376 (N_9376,N_9304,N_9374);
nor U9377 (N_9377,N_9273,N_9351);
nand U9378 (N_9378,N_9325,N_9259);
and U9379 (N_9379,N_9342,N_9336);
or U9380 (N_9380,N_9302,N_9289);
nand U9381 (N_9381,N_9332,N_9275);
nand U9382 (N_9382,N_9290,N_9260);
nor U9383 (N_9383,N_9330,N_9321);
or U9384 (N_9384,N_9284,N_9264);
or U9385 (N_9385,N_9353,N_9363);
nor U9386 (N_9386,N_9272,N_9251);
or U9387 (N_9387,N_9349,N_9310);
or U9388 (N_9388,N_9303,N_9270);
nor U9389 (N_9389,N_9262,N_9311);
xor U9390 (N_9390,N_9291,N_9314);
and U9391 (N_9391,N_9366,N_9287);
nand U9392 (N_9392,N_9345,N_9315);
nand U9393 (N_9393,N_9250,N_9335);
nor U9394 (N_9394,N_9357,N_9316);
nand U9395 (N_9395,N_9322,N_9295);
nor U9396 (N_9396,N_9308,N_9373);
or U9397 (N_9397,N_9309,N_9326);
nor U9398 (N_9398,N_9276,N_9288);
or U9399 (N_9399,N_9263,N_9296);
xor U9400 (N_9400,N_9369,N_9372);
or U9401 (N_9401,N_9344,N_9318);
nor U9402 (N_9402,N_9313,N_9274);
nand U9403 (N_9403,N_9282,N_9347);
and U9404 (N_9404,N_9281,N_9319);
and U9405 (N_9405,N_9283,N_9271);
nor U9406 (N_9406,N_9305,N_9348);
nor U9407 (N_9407,N_9277,N_9368);
or U9408 (N_9408,N_9266,N_9298);
nor U9409 (N_9409,N_9359,N_9261);
nor U9410 (N_9410,N_9364,N_9370);
nor U9411 (N_9411,N_9286,N_9301);
xnor U9412 (N_9412,N_9360,N_9329);
and U9413 (N_9413,N_9267,N_9350);
and U9414 (N_9414,N_9361,N_9320);
and U9415 (N_9415,N_9293,N_9269);
nand U9416 (N_9416,N_9312,N_9337);
xnor U9417 (N_9417,N_9331,N_9323);
xnor U9418 (N_9418,N_9362,N_9352);
nand U9419 (N_9419,N_9268,N_9339);
and U9420 (N_9420,N_9285,N_9306);
xor U9421 (N_9421,N_9328,N_9367);
or U9422 (N_9422,N_9355,N_9341);
nand U9423 (N_9423,N_9343,N_9300);
xor U9424 (N_9424,N_9324,N_9257);
and U9425 (N_9425,N_9254,N_9299);
or U9426 (N_9426,N_9280,N_9253);
and U9427 (N_9427,N_9356,N_9317);
and U9428 (N_9428,N_9354,N_9258);
or U9429 (N_9429,N_9279,N_9294);
or U9430 (N_9430,N_9256,N_9371);
and U9431 (N_9431,N_9265,N_9338);
nor U9432 (N_9432,N_9252,N_9340);
nand U9433 (N_9433,N_9292,N_9327);
xnor U9434 (N_9434,N_9334,N_9307);
nand U9435 (N_9435,N_9365,N_9346);
or U9436 (N_9436,N_9297,N_9333);
and U9437 (N_9437,N_9358,N_9296);
xor U9438 (N_9438,N_9310,N_9287);
or U9439 (N_9439,N_9298,N_9320);
xnor U9440 (N_9440,N_9274,N_9271);
xnor U9441 (N_9441,N_9374,N_9344);
nand U9442 (N_9442,N_9259,N_9280);
and U9443 (N_9443,N_9338,N_9348);
nor U9444 (N_9444,N_9373,N_9270);
xor U9445 (N_9445,N_9337,N_9331);
nand U9446 (N_9446,N_9252,N_9348);
xnor U9447 (N_9447,N_9258,N_9360);
xor U9448 (N_9448,N_9374,N_9261);
nor U9449 (N_9449,N_9287,N_9296);
nor U9450 (N_9450,N_9332,N_9297);
and U9451 (N_9451,N_9348,N_9335);
nand U9452 (N_9452,N_9312,N_9300);
or U9453 (N_9453,N_9255,N_9343);
or U9454 (N_9454,N_9349,N_9255);
xor U9455 (N_9455,N_9272,N_9352);
or U9456 (N_9456,N_9317,N_9261);
nand U9457 (N_9457,N_9282,N_9365);
nor U9458 (N_9458,N_9352,N_9340);
xnor U9459 (N_9459,N_9295,N_9373);
nand U9460 (N_9460,N_9293,N_9311);
xor U9461 (N_9461,N_9374,N_9293);
nand U9462 (N_9462,N_9310,N_9283);
nor U9463 (N_9463,N_9358,N_9363);
nand U9464 (N_9464,N_9276,N_9339);
xor U9465 (N_9465,N_9299,N_9305);
nand U9466 (N_9466,N_9250,N_9327);
or U9467 (N_9467,N_9355,N_9353);
nor U9468 (N_9468,N_9329,N_9354);
nand U9469 (N_9469,N_9367,N_9262);
nor U9470 (N_9470,N_9309,N_9318);
and U9471 (N_9471,N_9250,N_9264);
nand U9472 (N_9472,N_9321,N_9282);
and U9473 (N_9473,N_9285,N_9345);
nor U9474 (N_9474,N_9347,N_9352);
xor U9475 (N_9475,N_9251,N_9291);
or U9476 (N_9476,N_9358,N_9369);
and U9477 (N_9477,N_9270,N_9371);
nand U9478 (N_9478,N_9299,N_9252);
or U9479 (N_9479,N_9359,N_9347);
xor U9480 (N_9480,N_9351,N_9315);
nand U9481 (N_9481,N_9276,N_9258);
nand U9482 (N_9482,N_9346,N_9315);
nor U9483 (N_9483,N_9374,N_9320);
nand U9484 (N_9484,N_9316,N_9368);
nor U9485 (N_9485,N_9320,N_9310);
xor U9486 (N_9486,N_9281,N_9354);
nand U9487 (N_9487,N_9259,N_9329);
nor U9488 (N_9488,N_9307,N_9326);
nand U9489 (N_9489,N_9365,N_9317);
or U9490 (N_9490,N_9351,N_9253);
nor U9491 (N_9491,N_9307,N_9360);
nand U9492 (N_9492,N_9315,N_9344);
xnor U9493 (N_9493,N_9306,N_9257);
and U9494 (N_9494,N_9319,N_9316);
or U9495 (N_9495,N_9346,N_9324);
nor U9496 (N_9496,N_9290,N_9275);
and U9497 (N_9497,N_9307,N_9295);
nand U9498 (N_9498,N_9285,N_9363);
and U9499 (N_9499,N_9258,N_9294);
nor U9500 (N_9500,N_9454,N_9376);
xnor U9501 (N_9501,N_9422,N_9496);
and U9502 (N_9502,N_9443,N_9438);
or U9503 (N_9503,N_9483,N_9453);
nand U9504 (N_9504,N_9381,N_9377);
and U9505 (N_9505,N_9406,N_9391);
or U9506 (N_9506,N_9449,N_9468);
and U9507 (N_9507,N_9413,N_9408);
nand U9508 (N_9508,N_9436,N_9489);
nor U9509 (N_9509,N_9421,N_9401);
xnor U9510 (N_9510,N_9462,N_9497);
and U9511 (N_9511,N_9380,N_9476);
nor U9512 (N_9512,N_9465,N_9472);
or U9513 (N_9513,N_9393,N_9437);
and U9514 (N_9514,N_9446,N_9473);
nand U9515 (N_9515,N_9490,N_9403);
or U9516 (N_9516,N_9418,N_9389);
or U9517 (N_9517,N_9407,N_9390);
xnor U9518 (N_9518,N_9460,N_9451);
nor U9519 (N_9519,N_9387,N_9416);
xnor U9520 (N_9520,N_9411,N_9447);
nand U9521 (N_9521,N_9481,N_9385);
or U9522 (N_9522,N_9457,N_9441);
nand U9523 (N_9523,N_9397,N_9498);
xor U9524 (N_9524,N_9433,N_9414);
and U9525 (N_9525,N_9431,N_9402);
nor U9526 (N_9526,N_9459,N_9435);
xnor U9527 (N_9527,N_9494,N_9450);
and U9528 (N_9528,N_9452,N_9426);
nand U9529 (N_9529,N_9458,N_9399);
xnor U9530 (N_9530,N_9429,N_9434);
nand U9531 (N_9531,N_9386,N_9392);
or U9532 (N_9532,N_9427,N_9463);
nand U9533 (N_9533,N_9445,N_9383);
or U9534 (N_9534,N_9382,N_9432);
and U9535 (N_9535,N_9479,N_9398);
nand U9536 (N_9536,N_9404,N_9424);
nor U9537 (N_9537,N_9420,N_9395);
and U9538 (N_9538,N_9495,N_9417);
nand U9539 (N_9539,N_9470,N_9448);
and U9540 (N_9540,N_9480,N_9430);
xnor U9541 (N_9541,N_9461,N_9477);
xnor U9542 (N_9542,N_9499,N_9474);
nor U9543 (N_9543,N_9425,N_9487);
nand U9544 (N_9544,N_9405,N_9415);
xnor U9545 (N_9545,N_9423,N_9478);
xnor U9546 (N_9546,N_9469,N_9466);
nand U9547 (N_9547,N_9444,N_9409);
and U9548 (N_9548,N_9456,N_9439);
or U9549 (N_9549,N_9442,N_9455);
nand U9550 (N_9550,N_9375,N_9486);
and U9551 (N_9551,N_9410,N_9396);
nand U9552 (N_9552,N_9419,N_9491);
and U9553 (N_9553,N_9471,N_9482);
nand U9554 (N_9554,N_9484,N_9440);
nor U9555 (N_9555,N_9485,N_9475);
and U9556 (N_9556,N_9428,N_9493);
or U9557 (N_9557,N_9412,N_9379);
nor U9558 (N_9558,N_9492,N_9388);
xnor U9559 (N_9559,N_9394,N_9400);
or U9560 (N_9560,N_9378,N_9467);
xor U9561 (N_9561,N_9464,N_9384);
or U9562 (N_9562,N_9488,N_9389);
or U9563 (N_9563,N_9453,N_9470);
nand U9564 (N_9564,N_9400,N_9488);
and U9565 (N_9565,N_9423,N_9498);
nand U9566 (N_9566,N_9399,N_9405);
nor U9567 (N_9567,N_9428,N_9424);
xor U9568 (N_9568,N_9403,N_9407);
xnor U9569 (N_9569,N_9477,N_9427);
xnor U9570 (N_9570,N_9451,N_9431);
xor U9571 (N_9571,N_9428,N_9427);
nor U9572 (N_9572,N_9486,N_9475);
nand U9573 (N_9573,N_9398,N_9385);
or U9574 (N_9574,N_9466,N_9474);
or U9575 (N_9575,N_9448,N_9463);
and U9576 (N_9576,N_9479,N_9428);
xnor U9577 (N_9577,N_9409,N_9467);
xnor U9578 (N_9578,N_9445,N_9382);
nor U9579 (N_9579,N_9434,N_9403);
or U9580 (N_9580,N_9376,N_9423);
nand U9581 (N_9581,N_9437,N_9466);
and U9582 (N_9582,N_9442,N_9414);
nor U9583 (N_9583,N_9499,N_9497);
or U9584 (N_9584,N_9435,N_9384);
xor U9585 (N_9585,N_9433,N_9496);
nor U9586 (N_9586,N_9491,N_9450);
or U9587 (N_9587,N_9496,N_9404);
nand U9588 (N_9588,N_9424,N_9490);
xnor U9589 (N_9589,N_9428,N_9395);
or U9590 (N_9590,N_9391,N_9409);
nand U9591 (N_9591,N_9406,N_9412);
or U9592 (N_9592,N_9479,N_9408);
xnor U9593 (N_9593,N_9391,N_9447);
nand U9594 (N_9594,N_9457,N_9482);
xnor U9595 (N_9595,N_9459,N_9452);
xnor U9596 (N_9596,N_9421,N_9444);
and U9597 (N_9597,N_9383,N_9477);
and U9598 (N_9598,N_9475,N_9457);
xnor U9599 (N_9599,N_9426,N_9424);
and U9600 (N_9600,N_9460,N_9385);
and U9601 (N_9601,N_9398,N_9381);
nand U9602 (N_9602,N_9432,N_9384);
nor U9603 (N_9603,N_9483,N_9499);
xor U9604 (N_9604,N_9411,N_9461);
and U9605 (N_9605,N_9436,N_9466);
nand U9606 (N_9606,N_9447,N_9471);
nand U9607 (N_9607,N_9472,N_9454);
xor U9608 (N_9608,N_9409,N_9434);
nand U9609 (N_9609,N_9448,N_9477);
nor U9610 (N_9610,N_9436,N_9420);
xnor U9611 (N_9611,N_9431,N_9498);
nor U9612 (N_9612,N_9375,N_9492);
nor U9613 (N_9613,N_9397,N_9420);
nor U9614 (N_9614,N_9493,N_9424);
nand U9615 (N_9615,N_9413,N_9453);
nand U9616 (N_9616,N_9474,N_9495);
nor U9617 (N_9617,N_9444,N_9436);
and U9618 (N_9618,N_9495,N_9394);
and U9619 (N_9619,N_9485,N_9377);
nand U9620 (N_9620,N_9478,N_9406);
or U9621 (N_9621,N_9486,N_9399);
and U9622 (N_9622,N_9466,N_9487);
and U9623 (N_9623,N_9493,N_9491);
nand U9624 (N_9624,N_9488,N_9408);
or U9625 (N_9625,N_9616,N_9528);
xor U9626 (N_9626,N_9600,N_9525);
or U9627 (N_9627,N_9579,N_9511);
nand U9628 (N_9628,N_9572,N_9597);
and U9629 (N_9629,N_9564,N_9553);
nor U9630 (N_9630,N_9523,N_9582);
or U9631 (N_9631,N_9574,N_9527);
xor U9632 (N_9632,N_9522,N_9573);
nor U9633 (N_9633,N_9541,N_9568);
nand U9634 (N_9634,N_9529,N_9514);
nand U9635 (N_9635,N_9614,N_9585);
or U9636 (N_9636,N_9502,N_9599);
or U9637 (N_9637,N_9567,N_9534);
nor U9638 (N_9638,N_9587,N_9557);
or U9639 (N_9639,N_9612,N_9510);
nand U9640 (N_9640,N_9537,N_9601);
nor U9641 (N_9641,N_9613,N_9507);
and U9642 (N_9642,N_9596,N_9565);
xor U9643 (N_9643,N_9593,N_9563);
or U9644 (N_9644,N_9536,N_9531);
xnor U9645 (N_9645,N_9543,N_9551);
nand U9646 (N_9646,N_9586,N_9583);
and U9647 (N_9647,N_9542,N_9546);
nand U9648 (N_9648,N_9519,N_9520);
or U9649 (N_9649,N_9544,N_9506);
nor U9650 (N_9650,N_9526,N_9516);
nor U9651 (N_9651,N_9577,N_9503);
xor U9652 (N_9652,N_9580,N_9539);
or U9653 (N_9653,N_9549,N_9504);
or U9654 (N_9654,N_9512,N_9594);
nand U9655 (N_9655,N_9615,N_9603);
nor U9656 (N_9656,N_9558,N_9576);
or U9657 (N_9657,N_9556,N_9588);
nand U9658 (N_9658,N_9578,N_9521);
and U9659 (N_9659,N_9535,N_9575);
nand U9660 (N_9660,N_9619,N_9561);
nand U9661 (N_9661,N_9562,N_9530);
and U9662 (N_9662,N_9584,N_9569);
nor U9663 (N_9663,N_9545,N_9622);
or U9664 (N_9664,N_9589,N_9501);
nand U9665 (N_9665,N_9513,N_9595);
xor U9666 (N_9666,N_9500,N_9610);
nor U9667 (N_9667,N_9602,N_9566);
nor U9668 (N_9668,N_9559,N_9509);
xor U9669 (N_9669,N_9532,N_9581);
and U9670 (N_9670,N_9552,N_9538);
or U9671 (N_9671,N_9508,N_9518);
nor U9672 (N_9672,N_9590,N_9555);
or U9673 (N_9673,N_9623,N_9624);
xor U9674 (N_9674,N_9620,N_9548);
xor U9675 (N_9675,N_9524,N_9604);
and U9676 (N_9676,N_9554,N_9550);
nor U9677 (N_9677,N_9605,N_9606);
or U9678 (N_9678,N_9598,N_9609);
nor U9679 (N_9679,N_9540,N_9621);
and U9680 (N_9680,N_9617,N_9547);
xnor U9681 (N_9681,N_9560,N_9608);
xnor U9682 (N_9682,N_9505,N_9611);
xnor U9683 (N_9683,N_9515,N_9607);
nor U9684 (N_9684,N_9571,N_9517);
and U9685 (N_9685,N_9591,N_9570);
and U9686 (N_9686,N_9618,N_9592);
or U9687 (N_9687,N_9533,N_9593);
and U9688 (N_9688,N_9575,N_9607);
nand U9689 (N_9689,N_9545,N_9621);
nor U9690 (N_9690,N_9591,N_9584);
and U9691 (N_9691,N_9516,N_9540);
nor U9692 (N_9692,N_9546,N_9552);
and U9693 (N_9693,N_9513,N_9616);
nand U9694 (N_9694,N_9624,N_9611);
and U9695 (N_9695,N_9578,N_9535);
nor U9696 (N_9696,N_9527,N_9589);
and U9697 (N_9697,N_9544,N_9584);
and U9698 (N_9698,N_9619,N_9599);
and U9699 (N_9699,N_9541,N_9561);
nand U9700 (N_9700,N_9528,N_9545);
and U9701 (N_9701,N_9574,N_9619);
xor U9702 (N_9702,N_9507,N_9618);
nand U9703 (N_9703,N_9624,N_9537);
and U9704 (N_9704,N_9569,N_9578);
nor U9705 (N_9705,N_9511,N_9559);
nand U9706 (N_9706,N_9619,N_9531);
and U9707 (N_9707,N_9545,N_9610);
nor U9708 (N_9708,N_9581,N_9535);
and U9709 (N_9709,N_9562,N_9577);
and U9710 (N_9710,N_9516,N_9618);
xor U9711 (N_9711,N_9556,N_9531);
nor U9712 (N_9712,N_9571,N_9618);
nor U9713 (N_9713,N_9532,N_9500);
xnor U9714 (N_9714,N_9564,N_9500);
nor U9715 (N_9715,N_9505,N_9556);
or U9716 (N_9716,N_9533,N_9550);
nand U9717 (N_9717,N_9532,N_9604);
or U9718 (N_9718,N_9581,N_9613);
xor U9719 (N_9719,N_9612,N_9549);
nor U9720 (N_9720,N_9595,N_9550);
and U9721 (N_9721,N_9518,N_9581);
nand U9722 (N_9722,N_9574,N_9570);
nor U9723 (N_9723,N_9600,N_9596);
or U9724 (N_9724,N_9594,N_9533);
nor U9725 (N_9725,N_9616,N_9615);
nor U9726 (N_9726,N_9530,N_9573);
and U9727 (N_9727,N_9528,N_9566);
and U9728 (N_9728,N_9623,N_9598);
and U9729 (N_9729,N_9560,N_9533);
or U9730 (N_9730,N_9580,N_9610);
xor U9731 (N_9731,N_9574,N_9552);
or U9732 (N_9732,N_9617,N_9574);
nand U9733 (N_9733,N_9575,N_9505);
or U9734 (N_9734,N_9608,N_9536);
nand U9735 (N_9735,N_9569,N_9532);
and U9736 (N_9736,N_9515,N_9566);
and U9737 (N_9737,N_9605,N_9585);
nand U9738 (N_9738,N_9611,N_9623);
or U9739 (N_9739,N_9539,N_9575);
and U9740 (N_9740,N_9583,N_9506);
nor U9741 (N_9741,N_9538,N_9574);
xor U9742 (N_9742,N_9584,N_9600);
and U9743 (N_9743,N_9579,N_9539);
xnor U9744 (N_9744,N_9589,N_9553);
and U9745 (N_9745,N_9620,N_9536);
or U9746 (N_9746,N_9570,N_9609);
xnor U9747 (N_9747,N_9600,N_9612);
xor U9748 (N_9748,N_9520,N_9624);
nor U9749 (N_9749,N_9517,N_9594);
and U9750 (N_9750,N_9657,N_9710);
nor U9751 (N_9751,N_9635,N_9689);
xnor U9752 (N_9752,N_9724,N_9744);
and U9753 (N_9753,N_9640,N_9666);
xor U9754 (N_9754,N_9648,N_9638);
nand U9755 (N_9755,N_9726,N_9727);
or U9756 (N_9756,N_9684,N_9745);
nor U9757 (N_9757,N_9705,N_9665);
and U9758 (N_9758,N_9682,N_9631);
and U9759 (N_9759,N_9693,N_9697);
nand U9760 (N_9760,N_9652,N_9700);
xor U9761 (N_9761,N_9644,N_9737);
or U9762 (N_9762,N_9720,N_9680);
and U9763 (N_9763,N_9625,N_9650);
nor U9764 (N_9764,N_9733,N_9659);
xnor U9765 (N_9765,N_9729,N_9695);
and U9766 (N_9766,N_9655,N_9694);
or U9767 (N_9767,N_9628,N_9641);
nor U9768 (N_9768,N_9662,N_9653);
nor U9769 (N_9769,N_9723,N_9637);
nor U9770 (N_9770,N_9677,N_9658);
nor U9771 (N_9771,N_9669,N_9742);
and U9772 (N_9772,N_9743,N_9746);
nand U9773 (N_9773,N_9676,N_9674);
xor U9774 (N_9774,N_9688,N_9725);
and U9775 (N_9775,N_9714,N_9654);
nor U9776 (N_9776,N_9696,N_9634);
and U9777 (N_9777,N_9656,N_9717);
xor U9778 (N_9778,N_9704,N_9702);
xnor U9779 (N_9779,N_9730,N_9639);
nand U9780 (N_9780,N_9691,N_9713);
nand U9781 (N_9781,N_9703,N_9651);
nand U9782 (N_9782,N_9670,N_9711);
nand U9783 (N_9783,N_9626,N_9671);
and U9784 (N_9784,N_9706,N_9740);
nand U9785 (N_9785,N_9686,N_9632);
or U9786 (N_9786,N_9649,N_9718);
nand U9787 (N_9787,N_9692,N_9630);
or U9788 (N_9788,N_9629,N_9647);
nor U9789 (N_9789,N_9715,N_9728);
nor U9790 (N_9790,N_9681,N_9690);
nand U9791 (N_9791,N_9683,N_9721);
and U9792 (N_9792,N_9716,N_9735);
nand U9793 (N_9793,N_9709,N_9642);
nand U9794 (N_9794,N_9738,N_9739);
xnor U9795 (N_9795,N_9661,N_9667);
nand U9796 (N_9796,N_9707,N_9673);
and U9797 (N_9797,N_9645,N_9660);
nand U9798 (N_9798,N_9643,N_9675);
nand U9799 (N_9799,N_9627,N_9736);
and U9800 (N_9800,N_9708,N_9636);
or U9801 (N_9801,N_9719,N_9679);
and U9802 (N_9802,N_9747,N_9687);
and U9803 (N_9803,N_9685,N_9633);
nand U9804 (N_9804,N_9698,N_9731);
and U9805 (N_9805,N_9646,N_9749);
nor U9806 (N_9806,N_9678,N_9701);
or U9807 (N_9807,N_9722,N_9672);
xnor U9808 (N_9808,N_9732,N_9663);
nor U9809 (N_9809,N_9699,N_9712);
or U9810 (N_9810,N_9748,N_9734);
or U9811 (N_9811,N_9741,N_9668);
nor U9812 (N_9812,N_9664,N_9723);
nor U9813 (N_9813,N_9630,N_9709);
or U9814 (N_9814,N_9660,N_9692);
nor U9815 (N_9815,N_9744,N_9729);
nand U9816 (N_9816,N_9659,N_9664);
nor U9817 (N_9817,N_9736,N_9651);
and U9818 (N_9818,N_9678,N_9693);
xor U9819 (N_9819,N_9675,N_9746);
and U9820 (N_9820,N_9703,N_9638);
or U9821 (N_9821,N_9666,N_9675);
nor U9822 (N_9822,N_9655,N_9692);
nand U9823 (N_9823,N_9740,N_9671);
and U9824 (N_9824,N_9723,N_9746);
and U9825 (N_9825,N_9664,N_9694);
nand U9826 (N_9826,N_9744,N_9675);
and U9827 (N_9827,N_9720,N_9742);
xnor U9828 (N_9828,N_9655,N_9630);
nor U9829 (N_9829,N_9707,N_9668);
or U9830 (N_9830,N_9749,N_9715);
or U9831 (N_9831,N_9654,N_9680);
xor U9832 (N_9832,N_9673,N_9684);
xor U9833 (N_9833,N_9720,N_9677);
xor U9834 (N_9834,N_9678,N_9728);
xor U9835 (N_9835,N_9734,N_9670);
nor U9836 (N_9836,N_9705,N_9743);
nor U9837 (N_9837,N_9637,N_9661);
xnor U9838 (N_9838,N_9662,N_9735);
and U9839 (N_9839,N_9673,N_9721);
nor U9840 (N_9840,N_9705,N_9644);
or U9841 (N_9841,N_9731,N_9643);
or U9842 (N_9842,N_9634,N_9695);
nand U9843 (N_9843,N_9668,N_9679);
nand U9844 (N_9844,N_9732,N_9669);
or U9845 (N_9845,N_9704,N_9712);
or U9846 (N_9846,N_9659,N_9712);
xor U9847 (N_9847,N_9663,N_9742);
and U9848 (N_9848,N_9643,N_9647);
and U9849 (N_9849,N_9728,N_9723);
xnor U9850 (N_9850,N_9690,N_9636);
xnor U9851 (N_9851,N_9734,N_9686);
nand U9852 (N_9852,N_9633,N_9639);
nand U9853 (N_9853,N_9680,N_9699);
xor U9854 (N_9854,N_9663,N_9720);
or U9855 (N_9855,N_9730,N_9725);
and U9856 (N_9856,N_9740,N_9628);
nand U9857 (N_9857,N_9721,N_9731);
xnor U9858 (N_9858,N_9735,N_9703);
nand U9859 (N_9859,N_9656,N_9743);
and U9860 (N_9860,N_9708,N_9669);
or U9861 (N_9861,N_9698,N_9694);
nand U9862 (N_9862,N_9665,N_9721);
and U9863 (N_9863,N_9644,N_9668);
nand U9864 (N_9864,N_9625,N_9638);
nand U9865 (N_9865,N_9678,N_9663);
or U9866 (N_9866,N_9634,N_9661);
nand U9867 (N_9867,N_9690,N_9654);
or U9868 (N_9868,N_9663,N_9731);
and U9869 (N_9869,N_9638,N_9680);
nor U9870 (N_9870,N_9683,N_9746);
nor U9871 (N_9871,N_9637,N_9669);
nor U9872 (N_9872,N_9700,N_9649);
and U9873 (N_9873,N_9647,N_9714);
and U9874 (N_9874,N_9697,N_9657);
nor U9875 (N_9875,N_9786,N_9761);
and U9876 (N_9876,N_9850,N_9817);
and U9877 (N_9877,N_9764,N_9752);
and U9878 (N_9878,N_9868,N_9814);
xor U9879 (N_9879,N_9765,N_9768);
or U9880 (N_9880,N_9856,N_9800);
nand U9881 (N_9881,N_9854,N_9840);
xnor U9882 (N_9882,N_9867,N_9796);
nor U9883 (N_9883,N_9847,N_9843);
xor U9884 (N_9884,N_9872,N_9763);
xnor U9885 (N_9885,N_9809,N_9837);
xnor U9886 (N_9886,N_9871,N_9826);
nand U9887 (N_9887,N_9873,N_9835);
or U9888 (N_9888,N_9853,N_9783);
xnor U9889 (N_9889,N_9827,N_9760);
nand U9890 (N_9890,N_9848,N_9804);
nor U9891 (N_9891,N_9788,N_9767);
and U9892 (N_9892,N_9836,N_9816);
nor U9893 (N_9893,N_9785,N_9820);
nand U9894 (N_9894,N_9863,N_9864);
nand U9895 (N_9895,N_9852,N_9813);
nor U9896 (N_9896,N_9772,N_9861);
xor U9897 (N_9897,N_9787,N_9869);
nor U9898 (N_9898,N_9754,N_9771);
nor U9899 (N_9899,N_9812,N_9781);
nor U9900 (N_9900,N_9857,N_9789);
nor U9901 (N_9901,N_9818,N_9756);
or U9902 (N_9902,N_9762,N_9792);
nand U9903 (N_9903,N_9831,N_9801);
or U9904 (N_9904,N_9791,N_9790);
or U9905 (N_9905,N_9777,N_9825);
nor U9906 (N_9906,N_9779,N_9815);
nor U9907 (N_9907,N_9776,N_9844);
nand U9908 (N_9908,N_9819,N_9822);
or U9909 (N_9909,N_9859,N_9811);
or U9910 (N_9910,N_9849,N_9828);
nor U9911 (N_9911,N_9865,N_9842);
xnor U9912 (N_9912,N_9832,N_9807);
or U9913 (N_9913,N_9851,N_9773);
and U9914 (N_9914,N_9793,N_9798);
and U9915 (N_9915,N_9751,N_9855);
nor U9916 (N_9916,N_9806,N_9803);
xnor U9917 (N_9917,N_9799,N_9846);
nand U9918 (N_9918,N_9759,N_9866);
xor U9919 (N_9919,N_9824,N_9770);
or U9920 (N_9920,N_9795,N_9810);
nand U9921 (N_9921,N_9874,N_9841);
nor U9922 (N_9922,N_9802,N_9784);
or U9923 (N_9923,N_9862,N_9780);
xor U9924 (N_9924,N_9829,N_9757);
xor U9925 (N_9925,N_9830,N_9823);
nor U9926 (N_9926,N_9833,N_9794);
nor U9927 (N_9927,N_9838,N_9778);
xor U9928 (N_9928,N_9808,N_9839);
nand U9929 (N_9929,N_9750,N_9775);
or U9930 (N_9930,N_9753,N_9766);
or U9931 (N_9931,N_9769,N_9845);
nor U9932 (N_9932,N_9805,N_9858);
or U9933 (N_9933,N_9821,N_9797);
nand U9934 (N_9934,N_9774,N_9755);
xnor U9935 (N_9935,N_9834,N_9782);
nor U9936 (N_9936,N_9870,N_9758);
or U9937 (N_9937,N_9860,N_9782);
nor U9938 (N_9938,N_9768,N_9856);
xor U9939 (N_9939,N_9770,N_9825);
nand U9940 (N_9940,N_9831,N_9754);
nand U9941 (N_9941,N_9834,N_9852);
nand U9942 (N_9942,N_9868,N_9800);
nand U9943 (N_9943,N_9837,N_9822);
xor U9944 (N_9944,N_9853,N_9795);
nand U9945 (N_9945,N_9833,N_9827);
nor U9946 (N_9946,N_9795,N_9809);
nor U9947 (N_9947,N_9826,N_9784);
or U9948 (N_9948,N_9872,N_9842);
nand U9949 (N_9949,N_9817,N_9764);
nand U9950 (N_9950,N_9775,N_9801);
nand U9951 (N_9951,N_9816,N_9809);
nor U9952 (N_9952,N_9800,N_9815);
nor U9953 (N_9953,N_9785,N_9792);
nor U9954 (N_9954,N_9846,N_9756);
xor U9955 (N_9955,N_9750,N_9863);
xor U9956 (N_9956,N_9759,N_9814);
xor U9957 (N_9957,N_9801,N_9807);
xor U9958 (N_9958,N_9774,N_9789);
and U9959 (N_9959,N_9786,N_9826);
xor U9960 (N_9960,N_9768,N_9828);
nand U9961 (N_9961,N_9840,N_9805);
and U9962 (N_9962,N_9824,N_9861);
nand U9963 (N_9963,N_9784,N_9843);
nand U9964 (N_9964,N_9752,N_9807);
and U9965 (N_9965,N_9841,N_9821);
and U9966 (N_9966,N_9755,N_9862);
xor U9967 (N_9967,N_9836,N_9819);
nor U9968 (N_9968,N_9780,N_9803);
and U9969 (N_9969,N_9757,N_9762);
nor U9970 (N_9970,N_9753,N_9867);
xnor U9971 (N_9971,N_9852,N_9750);
xnor U9972 (N_9972,N_9865,N_9836);
xnor U9973 (N_9973,N_9857,N_9818);
or U9974 (N_9974,N_9794,N_9823);
and U9975 (N_9975,N_9802,N_9821);
nor U9976 (N_9976,N_9835,N_9824);
xor U9977 (N_9977,N_9789,N_9817);
and U9978 (N_9978,N_9757,N_9807);
xnor U9979 (N_9979,N_9765,N_9845);
nor U9980 (N_9980,N_9753,N_9829);
xnor U9981 (N_9981,N_9813,N_9752);
nor U9982 (N_9982,N_9755,N_9810);
xnor U9983 (N_9983,N_9868,N_9770);
nor U9984 (N_9984,N_9812,N_9791);
or U9985 (N_9985,N_9855,N_9863);
or U9986 (N_9986,N_9782,N_9783);
xnor U9987 (N_9987,N_9862,N_9787);
nor U9988 (N_9988,N_9846,N_9778);
and U9989 (N_9989,N_9762,N_9861);
or U9990 (N_9990,N_9854,N_9769);
nor U9991 (N_9991,N_9837,N_9792);
and U9992 (N_9992,N_9852,N_9766);
nand U9993 (N_9993,N_9859,N_9775);
nor U9994 (N_9994,N_9767,N_9866);
and U9995 (N_9995,N_9798,N_9755);
nand U9996 (N_9996,N_9783,N_9771);
or U9997 (N_9997,N_9779,N_9756);
nand U9998 (N_9998,N_9867,N_9771);
nand U9999 (N_9999,N_9873,N_9803);
xnor U10000 (N_10000,N_9977,N_9934);
xor U10001 (N_10001,N_9926,N_9880);
xor U10002 (N_10002,N_9893,N_9996);
nor U10003 (N_10003,N_9952,N_9989);
or U10004 (N_10004,N_9892,N_9954);
and U10005 (N_10005,N_9899,N_9973);
and U10006 (N_10006,N_9990,N_9928);
and U10007 (N_10007,N_9909,N_9895);
xnor U10008 (N_10008,N_9936,N_9964);
or U10009 (N_10009,N_9901,N_9907);
or U10010 (N_10010,N_9962,N_9987);
xnor U10011 (N_10011,N_9882,N_9980);
xor U10012 (N_10012,N_9995,N_9883);
or U10013 (N_10013,N_9931,N_9966);
xnor U10014 (N_10014,N_9997,N_9921);
or U10015 (N_10015,N_9947,N_9920);
nand U10016 (N_10016,N_9992,N_9906);
nor U10017 (N_10017,N_9976,N_9933);
xor U10018 (N_10018,N_9956,N_9941);
or U10019 (N_10019,N_9913,N_9985);
xor U10020 (N_10020,N_9958,N_9878);
and U10021 (N_10021,N_9879,N_9972);
xor U10022 (N_10022,N_9946,N_9963);
xor U10023 (N_10023,N_9905,N_9960);
xnor U10024 (N_10024,N_9875,N_9981);
nand U10025 (N_10025,N_9876,N_9935);
or U10026 (N_10026,N_9927,N_9929);
nand U10027 (N_10027,N_9983,N_9967);
nor U10028 (N_10028,N_9922,N_9953);
and U10029 (N_10029,N_9937,N_9910);
nand U10030 (N_10030,N_9884,N_9993);
xor U10031 (N_10031,N_9896,N_9915);
or U10032 (N_10032,N_9877,N_9961);
or U10033 (N_10033,N_9994,N_9968);
xnor U10034 (N_10034,N_9897,N_9942);
nand U10035 (N_10035,N_9894,N_9945);
nor U10036 (N_10036,N_9885,N_9979);
and U10037 (N_10037,N_9944,N_9938);
nor U10038 (N_10038,N_9943,N_9919);
xnor U10039 (N_10039,N_9902,N_9940);
and U10040 (N_10040,N_9889,N_9881);
and U10041 (N_10041,N_9969,N_9887);
and U10042 (N_10042,N_9932,N_9903);
and U10043 (N_10043,N_9939,N_9971);
and U10044 (N_10044,N_9984,N_9908);
xor U10045 (N_10045,N_9918,N_9911);
nor U10046 (N_10046,N_9904,N_9988);
and U10047 (N_10047,N_9916,N_9890);
nor U10048 (N_10048,N_9912,N_9959);
or U10049 (N_10049,N_9917,N_9974);
nand U10050 (N_10050,N_9888,N_9965);
and U10051 (N_10051,N_9886,N_9900);
or U10052 (N_10052,N_9970,N_9978);
nor U10053 (N_10053,N_9975,N_9930);
and U10054 (N_10054,N_9925,N_9986);
nand U10055 (N_10055,N_9950,N_9949);
xnor U10056 (N_10056,N_9914,N_9948);
or U10057 (N_10057,N_9999,N_9957);
nor U10058 (N_10058,N_9998,N_9891);
and U10059 (N_10059,N_9991,N_9951);
xnor U10060 (N_10060,N_9955,N_9923);
xor U10061 (N_10061,N_9924,N_9898);
and U10062 (N_10062,N_9982,N_9980);
nor U10063 (N_10063,N_9908,N_9919);
and U10064 (N_10064,N_9931,N_9897);
nand U10065 (N_10065,N_9930,N_9916);
or U10066 (N_10066,N_9955,N_9993);
xnor U10067 (N_10067,N_9953,N_9899);
and U10068 (N_10068,N_9949,N_9908);
xnor U10069 (N_10069,N_9977,N_9880);
nor U10070 (N_10070,N_9960,N_9947);
nor U10071 (N_10071,N_9909,N_9993);
nand U10072 (N_10072,N_9994,N_9996);
nand U10073 (N_10073,N_9949,N_9991);
nor U10074 (N_10074,N_9886,N_9915);
xnor U10075 (N_10075,N_9912,N_9955);
nand U10076 (N_10076,N_9961,N_9898);
nor U10077 (N_10077,N_9940,N_9922);
or U10078 (N_10078,N_9906,N_9875);
or U10079 (N_10079,N_9965,N_9955);
nor U10080 (N_10080,N_9902,N_9995);
xor U10081 (N_10081,N_9969,N_9968);
xor U10082 (N_10082,N_9981,N_9944);
or U10083 (N_10083,N_9911,N_9965);
xnor U10084 (N_10084,N_9991,N_9916);
and U10085 (N_10085,N_9952,N_9940);
or U10086 (N_10086,N_9959,N_9883);
nand U10087 (N_10087,N_9990,N_9957);
nand U10088 (N_10088,N_9995,N_9975);
nor U10089 (N_10089,N_9906,N_9898);
nor U10090 (N_10090,N_9882,N_9938);
nor U10091 (N_10091,N_9990,N_9912);
nand U10092 (N_10092,N_9942,N_9890);
nor U10093 (N_10093,N_9941,N_9934);
and U10094 (N_10094,N_9984,N_9923);
or U10095 (N_10095,N_9999,N_9989);
xor U10096 (N_10096,N_9946,N_9878);
or U10097 (N_10097,N_9932,N_9920);
and U10098 (N_10098,N_9986,N_9916);
nor U10099 (N_10099,N_9889,N_9885);
and U10100 (N_10100,N_9984,N_9988);
nand U10101 (N_10101,N_9900,N_9957);
nand U10102 (N_10102,N_9965,N_9971);
nor U10103 (N_10103,N_9987,N_9881);
xnor U10104 (N_10104,N_9920,N_9953);
nor U10105 (N_10105,N_9962,N_9890);
nor U10106 (N_10106,N_9905,N_9899);
or U10107 (N_10107,N_9915,N_9930);
nor U10108 (N_10108,N_9946,N_9897);
nand U10109 (N_10109,N_9926,N_9882);
and U10110 (N_10110,N_9919,N_9968);
nor U10111 (N_10111,N_9955,N_9876);
nor U10112 (N_10112,N_9951,N_9881);
and U10113 (N_10113,N_9915,N_9995);
or U10114 (N_10114,N_9927,N_9940);
or U10115 (N_10115,N_9999,N_9917);
nand U10116 (N_10116,N_9911,N_9959);
and U10117 (N_10117,N_9929,N_9937);
xor U10118 (N_10118,N_9998,N_9900);
nand U10119 (N_10119,N_9960,N_9984);
or U10120 (N_10120,N_9994,N_9953);
and U10121 (N_10121,N_9987,N_9908);
nor U10122 (N_10122,N_9905,N_9910);
xor U10123 (N_10123,N_9941,N_9960);
and U10124 (N_10124,N_9961,N_9909);
nor U10125 (N_10125,N_10064,N_10025);
and U10126 (N_10126,N_10092,N_10103);
nand U10127 (N_10127,N_10122,N_10116);
or U10128 (N_10128,N_10088,N_10048);
nand U10129 (N_10129,N_10083,N_10005);
or U10130 (N_10130,N_10007,N_10120);
and U10131 (N_10131,N_10101,N_10084);
nor U10132 (N_10132,N_10080,N_10115);
and U10133 (N_10133,N_10072,N_10001);
nand U10134 (N_10134,N_10014,N_10010);
and U10135 (N_10135,N_10026,N_10065);
or U10136 (N_10136,N_10114,N_10036);
xnor U10137 (N_10137,N_10021,N_10118);
nand U10138 (N_10138,N_10110,N_10105);
and U10139 (N_10139,N_10035,N_10073);
and U10140 (N_10140,N_10032,N_10063);
and U10141 (N_10141,N_10070,N_10058);
or U10142 (N_10142,N_10075,N_10076);
nor U10143 (N_10143,N_10056,N_10046);
xor U10144 (N_10144,N_10112,N_10109);
xnor U10145 (N_10145,N_10038,N_10100);
nand U10146 (N_10146,N_10106,N_10027);
nand U10147 (N_10147,N_10111,N_10028);
xnor U10148 (N_10148,N_10003,N_10067);
nor U10149 (N_10149,N_10008,N_10091);
xor U10150 (N_10150,N_10013,N_10078);
nand U10151 (N_10151,N_10011,N_10051);
nand U10152 (N_10152,N_10069,N_10040);
and U10153 (N_10153,N_10085,N_10098);
nor U10154 (N_10154,N_10086,N_10081);
nand U10155 (N_10155,N_10079,N_10107);
xnor U10156 (N_10156,N_10044,N_10093);
xnor U10157 (N_10157,N_10059,N_10094);
and U10158 (N_10158,N_10006,N_10102);
and U10159 (N_10159,N_10113,N_10041);
and U10160 (N_10160,N_10000,N_10031);
or U10161 (N_10161,N_10023,N_10045);
xnor U10162 (N_10162,N_10121,N_10039);
nand U10163 (N_10163,N_10024,N_10119);
nand U10164 (N_10164,N_10124,N_10049);
and U10165 (N_10165,N_10087,N_10009);
xnor U10166 (N_10166,N_10037,N_10053);
or U10167 (N_10167,N_10004,N_10019);
nand U10168 (N_10168,N_10052,N_10090);
nand U10169 (N_10169,N_10016,N_10033);
nor U10170 (N_10170,N_10002,N_10066);
nor U10171 (N_10171,N_10017,N_10055);
and U10172 (N_10172,N_10104,N_10020);
nor U10173 (N_10173,N_10089,N_10117);
and U10174 (N_10174,N_10062,N_10022);
or U10175 (N_10175,N_10082,N_10047);
nor U10176 (N_10176,N_10042,N_10057);
xor U10177 (N_10177,N_10099,N_10077);
and U10178 (N_10178,N_10123,N_10018);
nand U10179 (N_10179,N_10097,N_10096);
nor U10180 (N_10180,N_10012,N_10061);
or U10181 (N_10181,N_10029,N_10060);
xnor U10182 (N_10182,N_10015,N_10095);
or U10183 (N_10183,N_10068,N_10034);
and U10184 (N_10184,N_10030,N_10071);
xnor U10185 (N_10185,N_10054,N_10050);
and U10186 (N_10186,N_10074,N_10043);
nand U10187 (N_10187,N_10108,N_10032);
or U10188 (N_10188,N_10089,N_10028);
nand U10189 (N_10189,N_10121,N_10089);
or U10190 (N_10190,N_10082,N_10049);
xnor U10191 (N_10191,N_10047,N_10102);
and U10192 (N_10192,N_10111,N_10116);
nor U10193 (N_10193,N_10102,N_10120);
nand U10194 (N_10194,N_10117,N_10011);
and U10195 (N_10195,N_10025,N_10075);
nor U10196 (N_10196,N_10042,N_10026);
nand U10197 (N_10197,N_10014,N_10008);
nand U10198 (N_10198,N_10082,N_10114);
or U10199 (N_10199,N_10009,N_10018);
nor U10200 (N_10200,N_10011,N_10025);
and U10201 (N_10201,N_10024,N_10096);
or U10202 (N_10202,N_10033,N_10028);
nor U10203 (N_10203,N_10037,N_10085);
nor U10204 (N_10204,N_10003,N_10092);
xor U10205 (N_10205,N_10091,N_10054);
nor U10206 (N_10206,N_10014,N_10044);
or U10207 (N_10207,N_10012,N_10023);
nand U10208 (N_10208,N_10102,N_10027);
nor U10209 (N_10209,N_10105,N_10047);
nand U10210 (N_10210,N_10001,N_10124);
nand U10211 (N_10211,N_10098,N_10032);
nor U10212 (N_10212,N_10117,N_10087);
and U10213 (N_10213,N_10046,N_10086);
nand U10214 (N_10214,N_10039,N_10016);
or U10215 (N_10215,N_10083,N_10078);
or U10216 (N_10216,N_10115,N_10124);
nand U10217 (N_10217,N_10105,N_10023);
or U10218 (N_10218,N_10068,N_10056);
nand U10219 (N_10219,N_10036,N_10028);
or U10220 (N_10220,N_10013,N_10070);
and U10221 (N_10221,N_10005,N_10093);
xnor U10222 (N_10222,N_10122,N_10035);
and U10223 (N_10223,N_10036,N_10045);
or U10224 (N_10224,N_10046,N_10120);
xor U10225 (N_10225,N_10092,N_10037);
or U10226 (N_10226,N_10014,N_10089);
xor U10227 (N_10227,N_10044,N_10054);
nor U10228 (N_10228,N_10047,N_10053);
nor U10229 (N_10229,N_10097,N_10043);
nand U10230 (N_10230,N_10072,N_10081);
and U10231 (N_10231,N_10022,N_10031);
nor U10232 (N_10232,N_10119,N_10004);
nand U10233 (N_10233,N_10021,N_10077);
and U10234 (N_10234,N_10105,N_10002);
nor U10235 (N_10235,N_10034,N_10092);
nor U10236 (N_10236,N_10122,N_10071);
nand U10237 (N_10237,N_10004,N_10091);
nand U10238 (N_10238,N_10027,N_10076);
and U10239 (N_10239,N_10011,N_10108);
or U10240 (N_10240,N_10012,N_10011);
xnor U10241 (N_10241,N_10045,N_10124);
or U10242 (N_10242,N_10010,N_10016);
and U10243 (N_10243,N_10105,N_10038);
or U10244 (N_10244,N_10048,N_10104);
nand U10245 (N_10245,N_10053,N_10001);
nor U10246 (N_10246,N_10080,N_10121);
nand U10247 (N_10247,N_10043,N_10072);
and U10248 (N_10248,N_10053,N_10081);
nand U10249 (N_10249,N_10035,N_10071);
xor U10250 (N_10250,N_10223,N_10184);
nand U10251 (N_10251,N_10133,N_10140);
or U10252 (N_10252,N_10201,N_10145);
and U10253 (N_10253,N_10134,N_10238);
xor U10254 (N_10254,N_10171,N_10217);
xor U10255 (N_10255,N_10172,N_10150);
nor U10256 (N_10256,N_10127,N_10245);
xnor U10257 (N_10257,N_10181,N_10174);
or U10258 (N_10258,N_10229,N_10227);
xnor U10259 (N_10259,N_10225,N_10210);
nand U10260 (N_10260,N_10149,N_10222);
and U10261 (N_10261,N_10239,N_10230);
and U10262 (N_10262,N_10207,N_10236);
nor U10263 (N_10263,N_10167,N_10205);
xnor U10264 (N_10264,N_10160,N_10211);
and U10265 (N_10265,N_10189,N_10125);
and U10266 (N_10266,N_10219,N_10138);
or U10267 (N_10267,N_10213,N_10154);
or U10268 (N_10268,N_10182,N_10148);
nand U10269 (N_10269,N_10224,N_10235);
nor U10270 (N_10270,N_10180,N_10214);
nor U10271 (N_10271,N_10247,N_10226);
xnor U10272 (N_10272,N_10212,N_10153);
nor U10273 (N_10273,N_10215,N_10168);
and U10274 (N_10274,N_10199,N_10204);
xnor U10275 (N_10275,N_10128,N_10129);
nand U10276 (N_10276,N_10203,N_10132);
nand U10277 (N_10277,N_10208,N_10157);
and U10278 (N_10278,N_10188,N_10232);
nand U10279 (N_10279,N_10241,N_10177);
xor U10280 (N_10280,N_10151,N_10244);
nor U10281 (N_10281,N_10146,N_10200);
nor U10282 (N_10282,N_10228,N_10193);
nand U10283 (N_10283,N_10152,N_10198);
nand U10284 (N_10284,N_10209,N_10173);
nor U10285 (N_10285,N_10143,N_10183);
nand U10286 (N_10286,N_10194,N_10165);
nand U10287 (N_10287,N_10195,N_10190);
nand U10288 (N_10288,N_10248,N_10186);
nor U10289 (N_10289,N_10162,N_10161);
nand U10290 (N_10290,N_10246,N_10220);
xor U10291 (N_10291,N_10136,N_10231);
and U10292 (N_10292,N_10192,N_10163);
and U10293 (N_10293,N_10155,N_10202);
and U10294 (N_10294,N_10130,N_10137);
nor U10295 (N_10295,N_10216,N_10131);
nand U10296 (N_10296,N_10142,N_10249);
xnor U10297 (N_10297,N_10126,N_10233);
nand U10298 (N_10298,N_10240,N_10139);
xnor U10299 (N_10299,N_10237,N_10141);
nand U10300 (N_10300,N_10164,N_10135);
nor U10301 (N_10301,N_10234,N_10243);
or U10302 (N_10302,N_10170,N_10187);
or U10303 (N_10303,N_10191,N_10158);
xor U10304 (N_10304,N_10179,N_10218);
or U10305 (N_10305,N_10185,N_10242);
and U10306 (N_10306,N_10178,N_10169);
and U10307 (N_10307,N_10144,N_10221);
xor U10308 (N_10308,N_10176,N_10197);
and U10309 (N_10309,N_10175,N_10147);
or U10310 (N_10310,N_10156,N_10206);
xor U10311 (N_10311,N_10159,N_10166);
or U10312 (N_10312,N_10196,N_10241);
and U10313 (N_10313,N_10227,N_10147);
and U10314 (N_10314,N_10220,N_10226);
and U10315 (N_10315,N_10196,N_10206);
xnor U10316 (N_10316,N_10217,N_10182);
or U10317 (N_10317,N_10225,N_10144);
xor U10318 (N_10318,N_10228,N_10238);
and U10319 (N_10319,N_10247,N_10228);
nor U10320 (N_10320,N_10242,N_10173);
and U10321 (N_10321,N_10242,N_10213);
nor U10322 (N_10322,N_10185,N_10172);
or U10323 (N_10323,N_10137,N_10231);
nor U10324 (N_10324,N_10159,N_10133);
or U10325 (N_10325,N_10145,N_10187);
or U10326 (N_10326,N_10141,N_10194);
or U10327 (N_10327,N_10168,N_10134);
nor U10328 (N_10328,N_10125,N_10137);
nor U10329 (N_10329,N_10126,N_10195);
or U10330 (N_10330,N_10205,N_10245);
xor U10331 (N_10331,N_10127,N_10220);
or U10332 (N_10332,N_10232,N_10141);
or U10333 (N_10333,N_10174,N_10240);
nor U10334 (N_10334,N_10131,N_10173);
and U10335 (N_10335,N_10135,N_10201);
and U10336 (N_10336,N_10137,N_10164);
nor U10337 (N_10337,N_10211,N_10224);
xor U10338 (N_10338,N_10152,N_10135);
and U10339 (N_10339,N_10200,N_10139);
and U10340 (N_10340,N_10211,N_10164);
xnor U10341 (N_10341,N_10183,N_10162);
or U10342 (N_10342,N_10169,N_10192);
nand U10343 (N_10343,N_10134,N_10202);
or U10344 (N_10344,N_10128,N_10184);
and U10345 (N_10345,N_10165,N_10137);
nor U10346 (N_10346,N_10187,N_10203);
nor U10347 (N_10347,N_10166,N_10200);
and U10348 (N_10348,N_10168,N_10204);
xor U10349 (N_10349,N_10230,N_10127);
nor U10350 (N_10350,N_10217,N_10193);
and U10351 (N_10351,N_10125,N_10231);
nor U10352 (N_10352,N_10173,N_10169);
xnor U10353 (N_10353,N_10186,N_10244);
nor U10354 (N_10354,N_10203,N_10159);
and U10355 (N_10355,N_10125,N_10180);
xor U10356 (N_10356,N_10241,N_10208);
xnor U10357 (N_10357,N_10131,N_10235);
nor U10358 (N_10358,N_10141,N_10138);
nor U10359 (N_10359,N_10198,N_10179);
and U10360 (N_10360,N_10225,N_10158);
or U10361 (N_10361,N_10211,N_10228);
and U10362 (N_10362,N_10221,N_10164);
nor U10363 (N_10363,N_10167,N_10175);
or U10364 (N_10364,N_10195,N_10162);
and U10365 (N_10365,N_10195,N_10225);
nor U10366 (N_10366,N_10233,N_10202);
and U10367 (N_10367,N_10134,N_10164);
xnor U10368 (N_10368,N_10158,N_10184);
and U10369 (N_10369,N_10211,N_10177);
nand U10370 (N_10370,N_10236,N_10227);
xnor U10371 (N_10371,N_10182,N_10155);
nand U10372 (N_10372,N_10166,N_10178);
or U10373 (N_10373,N_10163,N_10215);
xnor U10374 (N_10374,N_10160,N_10228);
xnor U10375 (N_10375,N_10337,N_10250);
nand U10376 (N_10376,N_10348,N_10283);
nor U10377 (N_10377,N_10274,N_10363);
nor U10378 (N_10378,N_10315,N_10260);
and U10379 (N_10379,N_10307,N_10281);
and U10380 (N_10380,N_10258,N_10264);
or U10381 (N_10381,N_10333,N_10361);
xor U10382 (N_10382,N_10343,N_10265);
and U10383 (N_10383,N_10278,N_10326);
nand U10384 (N_10384,N_10293,N_10341);
nand U10385 (N_10385,N_10295,N_10368);
xnor U10386 (N_10386,N_10325,N_10329);
or U10387 (N_10387,N_10310,N_10262);
xor U10388 (N_10388,N_10317,N_10279);
nor U10389 (N_10389,N_10339,N_10352);
or U10390 (N_10390,N_10273,N_10365);
and U10391 (N_10391,N_10320,N_10267);
nor U10392 (N_10392,N_10345,N_10327);
or U10393 (N_10393,N_10364,N_10312);
and U10394 (N_10394,N_10269,N_10266);
nor U10395 (N_10395,N_10271,N_10306);
and U10396 (N_10396,N_10372,N_10287);
xnor U10397 (N_10397,N_10336,N_10355);
xor U10398 (N_10398,N_10369,N_10297);
and U10399 (N_10399,N_10354,N_10370);
nand U10400 (N_10400,N_10276,N_10308);
nor U10401 (N_10401,N_10268,N_10334);
nor U10402 (N_10402,N_10322,N_10299);
or U10403 (N_10403,N_10255,N_10261);
or U10404 (N_10404,N_10351,N_10340);
or U10405 (N_10405,N_10374,N_10323);
nor U10406 (N_10406,N_10366,N_10263);
xnor U10407 (N_10407,N_10302,N_10290);
nand U10408 (N_10408,N_10304,N_10311);
or U10409 (N_10409,N_10277,N_10358);
xor U10410 (N_10410,N_10346,N_10252);
and U10411 (N_10411,N_10344,N_10331);
nor U10412 (N_10412,N_10257,N_10324);
nor U10413 (N_10413,N_10338,N_10305);
nor U10414 (N_10414,N_10301,N_10282);
nand U10415 (N_10415,N_10272,N_10330);
nor U10416 (N_10416,N_10280,N_10321);
nor U10417 (N_10417,N_10285,N_10319);
or U10418 (N_10418,N_10356,N_10291);
nand U10419 (N_10419,N_10303,N_10309);
nor U10420 (N_10420,N_10342,N_10298);
xnor U10421 (N_10421,N_10253,N_10300);
nor U10422 (N_10422,N_10349,N_10350);
and U10423 (N_10423,N_10288,N_10296);
nor U10424 (N_10424,N_10254,N_10332);
nand U10425 (N_10425,N_10373,N_10371);
and U10426 (N_10426,N_10316,N_10314);
nand U10427 (N_10427,N_10328,N_10259);
and U10428 (N_10428,N_10357,N_10251);
nand U10429 (N_10429,N_10335,N_10360);
and U10430 (N_10430,N_10275,N_10294);
xor U10431 (N_10431,N_10353,N_10359);
xnor U10432 (N_10432,N_10284,N_10362);
nand U10433 (N_10433,N_10270,N_10289);
or U10434 (N_10434,N_10318,N_10313);
nor U10435 (N_10435,N_10292,N_10347);
or U10436 (N_10436,N_10367,N_10256);
nand U10437 (N_10437,N_10286,N_10328);
nand U10438 (N_10438,N_10307,N_10254);
xor U10439 (N_10439,N_10335,N_10331);
xor U10440 (N_10440,N_10267,N_10265);
nand U10441 (N_10441,N_10285,N_10252);
and U10442 (N_10442,N_10370,N_10368);
nand U10443 (N_10443,N_10289,N_10340);
nand U10444 (N_10444,N_10283,N_10260);
xor U10445 (N_10445,N_10279,N_10353);
or U10446 (N_10446,N_10263,N_10293);
nand U10447 (N_10447,N_10299,N_10305);
nor U10448 (N_10448,N_10286,N_10278);
and U10449 (N_10449,N_10266,N_10319);
nand U10450 (N_10450,N_10359,N_10345);
or U10451 (N_10451,N_10291,N_10362);
and U10452 (N_10452,N_10373,N_10289);
and U10453 (N_10453,N_10301,N_10278);
nor U10454 (N_10454,N_10372,N_10303);
and U10455 (N_10455,N_10315,N_10300);
xor U10456 (N_10456,N_10303,N_10268);
or U10457 (N_10457,N_10279,N_10311);
and U10458 (N_10458,N_10329,N_10330);
nand U10459 (N_10459,N_10328,N_10332);
xnor U10460 (N_10460,N_10324,N_10267);
xnor U10461 (N_10461,N_10315,N_10270);
or U10462 (N_10462,N_10302,N_10330);
and U10463 (N_10463,N_10259,N_10290);
and U10464 (N_10464,N_10259,N_10373);
or U10465 (N_10465,N_10260,N_10250);
or U10466 (N_10466,N_10364,N_10297);
nor U10467 (N_10467,N_10295,N_10269);
nor U10468 (N_10468,N_10332,N_10325);
nor U10469 (N_10469,N_10341,N_10258);
xnor U10470 (N_10470,N_10301,N_10303);
nor U10471 (N_10471,N_10286,N_10254);
nor U10472 (N_10472,N_10354,N_10294);
and U10473 (N_10473,N_10323,N_10266);
and U10474 (N_10474,N_10274,N_10304);
nand U10475 (N_10475,N_10331,N_10352);
or U10476 (N_10476,N_10307,N_10348);
and U10477 (N_10477,N_10343,N_10349);
and U10478 (N_10478,N_10320,N_10317);
nand U10479 (N_10479,N_10321,N_10304);
nand U10480 (N_10480,N_10302,N_10356);
nand U10481 (N_10481,N_10365,N_10309);
or U10482 (N_10482,N_10265,N_10325);
xor U10483 (N_10483,N_10263,N_10272);
and U10484 (N_10484,N_10322,N_10359);
or U10485 (N_10485,N_10326,N_10271);
nand U10486 (N_10486,N_10311,N_10332);
nor U10487 (N_10487,N_10370,N_10281);
and U10488 (N_10488,N_10343,N_10323);
and U10489 (N_10489,N_10285,N_10342);
xor U10490 (N_10490,N_10292,N_10284);
or U10491 (N_10491,N_10255,N_10320);
nand U10492 (N_10492,N_10299,N_10263);
or U10493 (N_10493,N_10305,N_10344);
xor U10494 (N_10494,N_10296,N_10265);
and U10495 (N_10495,N_10333,N_10326);
xor U10496 (N_10496,N_10332,N_10266);
nand U10497 (N_10497,N_10360,N_10325);
nor U10498 (N_10498,N_10303,N_10359);
and U10499 (N_10499,N_10365,N_10280);
and U10500 (N_10500,N_10473,N_10408);
xor U10501 (N_10501,N_10461,N_10484);
and U10502 (N_10502,N_10451,N_10385);
xnor U10503 (N_10503,N_10420,N_10425);
and U10504 (N_10504,N_10431,N_10433);
nor U10505 (N_10505,N_10468,N_10384);
nor U10506 (N_10506,N_10470,N_10392);
and U10507 (N_10507,N_10496,N_10445);
nand U10508 (N_10508,N_10448,N_10409);
or U10509 (N_10509,N_10487,N_10395);
nand U10510 (N_10510,N_10377,N_10447);
or U10511 (N_10511,N_10383,N_10401);
nand U10512 (N_10512,N_10397,N_10486);
nor U10513 (N_10513,N_10480,N_10376);
or U10514 (N_10514,N_10426,N_10441);
nand U10515 (N_10515,N_10400,N_10458);
nor U10516 (N_10516,N_10378,N_10379);
or U10517 (N_10517,N_10396,N_10424);
nand U10518 (N_10518,N_10412,N_10485);
nand U10519 (N_10519,N_10499,N_10465);
nand U10520 (N_10520,N_10413,N_10483);
nor U10521 (N_10521,N_10399,N_10466);
and U10522 (N_10522,N_10454,N_10393);
and U10523 (N_10523,N_10435,N_10429);
nor U10524 (N_10524,N_10491,N_10398);
nand U10525 (N_10525,N_10423,N_10476);
nand U10526 (N_10526,N_10493,N_10416);
nor U10527 (N_10527,N_10471,N_10456);
and U10528 (N_10528,N_10481,N_10494);
nand U10529 (N_10529,N_10391,N_10449);
nor U10530 (N_10530,N_10453,N_10455);
or U10531 (N_10531,N_10452,N_10410);
and U10532 (N_10532,N_10404,N_10422);
or U10533 (N_10533,N_10469,N_10421);
and U10534 (N_10534,N_10442,N_10457);
or U10535 (N_10535,N_10459,N_10437);
nand U10536 (N_10536,N_10394,N_10406);
nor U10537 (N_10537,N_10430,N_10434);
xnor U10538 (N_10538,N_10482,N_10444);
xnor U10539 (N_10539,N_10477,N_10464);
or U10540 (N_10540,N_10415,N_10436);
nand U10541 (N_10541,N_10488,N_10386);
nand U10542 (N_10542,N_10495,N_10382);
and U10543 (N_10543,N_10478,N_10407);
xor U10544 (N_10544,N_10389,N_10450);
nor U10545 (N_10545,N_10402,N_10387);
or U10546 (N_10546,N_10432,N_10467);
nor U10547 (N_10547,N_10438,N_10446);
xor U10548 (N_10548,N_10475,N_10474);
and U10549 (N_10549,N_10489,N_10427);
nand U10550 (N_10550,N_10390,N_10381);
xor U10551 (N_10551,N_10497,N_10460);
nand U10552 (N_10552,N_10472,N_10380);
nand U10553 (N_10553,N_10479,N_10417);
nor U10554 (N_10554,N_10498,N_10462);
nand U10555 (N_10555,N_10492,N_10419);
nor U10556 (N_10556,N_10440,N_10463);
and U10557 (N_10557,N_10388,N_10418);
xnor U10558 (N_10558,N_10414,N_10490);
xor U10559 (N_10559,N_10411,N_10403);
nor U10560 (N_10560,N_10439,N_10375);
xor U10561 (N_10561,N_10443,N_10428);
or U10562 (N_10562,N_10405,N_10434);
or U10563 (N_10563,N_10499,N_10420);
and U10564 (N_10564,N_10403,N_10378);
and U10565 (N_10565,N_10484,N_10406);
nor U10566 (N_10566,N_10486,N_10442);
nor U10567 (N_10567,N_10439,N_10471);
nor U10568 (N_10568,N_10430,N_10483);
nand U10569 (N_10569,N_10489,N_10379);
xnor U10570 (N_10570,N_10406,N_10435);
nand U10571 (N_10571,N_10412,N_10421);
and U10572 (N_10572,N_10429,N_10424);
nand U10573 (N_10573,N_10436,N_10388);
nand U10574 (N_10574,N_10457,N_10392);
xor U10575 (N_10575,N_10475,N_10446);
and U10576 (N_10576,N_10492,N_10396);
or U10577 (N_10577,N_10458,N_10409);
and U10578 (N_10578,N_10445,N_10413);
nor U10579 (N_10579,N_10485,N_10469);
and U10580 (N_10580,N_10393,N_10475);
and U10581 (N_10581,N_10379,N_10392);
nor U10582 (N_10582,N_10407,N_10467);
or U10583 (N_10583,N_10492,N_10435);
and U10584 (N_10584,N_10416,N_10431);
nand U10585 (N_10585,N_10443,N_10385);
and U10586 (N_10586,N_10417,N_10387);
xnor U10587 (N_10587,N_10419,N_10456);
xor U10588 (N_10588,N_10393,N_10396);
xor U10589 (N_10589,N_10413,N_10422);
nor U10590 (N_10590,N_10490,N_10450);
nor U10591 (N_10591,N_10380,N_10424);
xnor U10592 (N_10592,N_10441,N_10438);
nor U10593 (N_10593,N_10418,N_10466);
xor U10594 (N_10594,N_10418,N_10497);
nor U10595 (N_10595,N_10470,N_10378);
nor U10596 (N_10596,N_10462,N_10427);
nor U10597 (N_10597,N_10420,N_10462);
and U10598 (N_10598,N_10386,N_10427);
and U10599 (N_10599,N_10419,N_10485);
nor U10600 (N_10600,N_10477,N_10408);
nand U10601 (N_10601,N_10463,N_10399);
xnor U10602 (N_10602,N_10457,N_10391);
and U10603 (N_10603,N_10405,N_10416);
xor U10604 (N_10604,N_10444,N_10384);
xnor U10605 (N_10605,N_10400,N_10492);
and U10606 (N_10606,N_10420,N_10406);
xnor U10607 (N_10607,N_10435,N_10439);
nor U10608 (N_10608,N_10450,N_10382);
or U10609 (N_10609,N_10379,N_10394);
or U10610 (N_10610,N_10398,N_10418);
or U10611 (N_10611,N_10487,N_10405);
nor U10612 (N_10612,N_10472,N_10496);
nand U10613 (N_10613,N_10396,N_10445);
or U10614 (N_10614,N_10475,N_10489);
nor U10615 (N_10615,N_10415,N_10403);
xor U10616 (N_10616,N_10444,N_10439);
or U10617 (N_10617,N_10413,N_10484);
nor U10618 (N_10618,N_10411,N_10435);
nor U10619 (N_10619,N_10439,N_10388);
and U10620 (N_10620,N_10453,N_10469);
nand U10621 (N_10621,N_10453,N_10489);
nand U10622 (N_10622,N_10395,N_10429);
nor U10623 (N_10623,N_10483,N_10403);
xor U10624 (N_10624,N_10390,N_10389);
nor U10625 (N_10625,N_10522,N_10600);
or U10626 (N_10626,N_10501,N_10549);
or U10627 (N_10627,N_10507,N_10580);
and U10628 (N_10628,N_10534,N_10526);
nor U10629 (N_10629,N_10506,N_10578);
nand U10630 (N_10630,N_10556,N_10574);
or U10631 (N_10631,N_10546,N_10570);
nor U10632 (N_10632,N_10528,N_10518);
and U10633 (N_10633,N_10609,N_10510);
xnor U10634 (N_10634,N_10604,N_10531);
and U10635 (N_10635,N_10512,N_10591);
nor U10636 (N_10636,N_10513,N_10595);
nand U10637 (N_10637,N_10532,N_10523);
or U10638 (N_10638,N_10589,N_10542);
or U10639 (N_10639,N_10582,N_10541);
or U10640 (N_10640,N_10588,N_10547);
and U10641 (N_10641,N_10535,N_10552);
or U10642 (N_10642,N_10607,N_10605);
nor U10643 (N_10643,N_10515,N_10621);
nor U10644 (N_10644,N_10606,N_10553);
xnor U10645 (N_10645,N_10503,N_10576);
nor U10646 (N_10646,N_10573,N_10587);
or U10647 (N_10647,N_10601,N_10554);
or U10648 (N_10648,N_10530,N_10505);
and U10649 (N_10649,N_10559,N_10598);
or U10650 (N_10650,N_10525,N_10536);
and U10651 (N_10651,N_10514,N_10551);
nor U10652 (N_10652,N_10623,N_10516);
and U10653 (N_10653,N_10548,N_10584);
or U10654 (N_10654,N_10543,N_10555);
nor U10655 (N_10655,N_10557,N_10617);
and U10656 (N_10656,N_10565,N_10561);
and U10657 (N_10657,N_10544,N_10524);
nor U10658 (N_10658,N_10567,N_10614);
or U10659 (N_10659,N_10602,N_10519);
or U10660 (N_10660,N_10599,N_10593);
and U10661 (N_10661,N_10564,N_10579);
nand U10662 (N_10662,N_10571,N_10608);
xor U10663 (N_10663,N_10615,N_10618);
xnor U10664 (N_10664,N_10517,N_10619);
nand U10665 (N_10665,N_10533,N_10572);
nand U10666 (N_10666,N_10622,N_10502);
nor U10667 (N_10667,N_10500,N_10583);
and U10668 (N_10668,N_10624,N_10611);
nand U10669 (N_10669,N_10529,N_10566);
nor U10670 (N_10670,N_10597,N_10537);
and U10671 (N_10671,N_10545,N_10575);
nand U10672 (N_10672,N_10508,N_10568);
and U10673 (N_10673,N_10563,N_10550);
nor U10674 (N_10674,N_10616,N_10596);
nor U10675 (N_10675,N_10592,N_10585);
nor U10676 (N_10676,N_10540,N_10577);
nor U10677 (N_10677,N_10586,N_10539);
xor U10678 (N_10678,N_10511,N_10569);
and U10679 (N_10679,N_10603,N_10590);
nand U10680 (N_10680,N_10594,N_10504);
or U10681 (N_10681,N_10521,N_10527);
or U10682 (N_10682,N_10538,N_10520);
or U10683 (N_10683,N_10558,N_10620);
nand U10684 (N_10684,N_10610,N_10509);
nor U10685 (N_10685,N_10613,N_10612);
nor U10686 (N_10686,N_10562,N_10581);
or U10687 (N_10687,N_10560,N_10524);
nand U10688 (N_10688,N_10564,N_10573);
nor U10689 (N_10689,N_10567,N_10557);
and U10690 (N_10690,N_10619,N_10532);
nand U10691 (N_10691,N_10589,N_10571);
xnor U10692 (N_10692,N_10620,N_10500);
nand U10693 (N_10693,N_10594,N_10503);
and U10694 (N_10694,N_10514,N_10553);
or U10695 (N_10695,N_10621,N_10558);
or U10696 (N_10696,N_10596,N_10594);
and U10697 (N_10697,N_10529,N_10624);
nor U10698 (N_10698,N_10613,N_10611);
nor U10699 (N_10699,N_10507,N_10556);
nor U10700 (N_10700,N_10618,N_10532);
nand U10701 (N_10701,N_10512,N_10562);
nand U10702 (N_10702,N_10617,N_10531);
or U10703 (N_10703,N_10513,N_10591);
nor U10704 (N_10704,N_10512,N_10540);
or U10705 (N_10705,N_10515,N_10547);
nand U10706 (N_10706,N_10581,N_10595);
nand U10707 (N_10707,N_10569,N_10595);
xor U10708 (N_10708,N_10598,N_10523);
or U10709 (N_10709,N_10508,N_10511);
and U10710 (N_10710,N_10611,N_10569);
or U10711 (N_10711,N_10527,N_10556);
or U10712 (N_10712,N_10619,N_10513);
xnor U10713 (N_10713,N_10594,N_10606);
nand U10714 (N_10714,N_10519,N_10542);
and U10715 (N_10715,N_10603,N_10607);
nand U10716 (N_10716,N_10574,N_10553);
or U10717 (N_10717,N_10573,N_10524);
and U10718 (N_10718,N_10568,N_10585);
or U10719 (N_10719,N_10618,N_10597);
nand U10720 (N_10720,N_10622,N_10587);
nand U10721 (N_10721,N_10515,N_10583);
xnor U10722 (N_10722,N_10609,N_10535);
nor U10723 (N_10723,N_10617,N_10587);
or U10724 (N_10724,N_10620,N_10539);
xor U10725 (N_10725,N_10562,N_10619);
or U10726 (N_10726,N_10503,N_10582);
xor U10727 (N_10727,N_10578,N_10591);
xnor U10728 (N_10728,N_10553,N_10565);
xor U10729 (N_10729,N_10577,N_10616);
nand U10730 (N_10730,N_10585,N_10603);
nand U10731 (N_10731,N_10523,N_10581);
or U10732 (N_10732,N_10585,N_10605);
nand U10733 (N_10733,N_10608,N_10525);
and U10734 (N_10734,N_10561,N_10553);
nor U10735 (N_10735,N_10504,N_10559);
nand U10736 (N_10736,N_10555,N_10619);
nand U10737 (N_10737,N_10562,N_10526);
nand U10738 (N_10738,N_10525,N_10505);
and U10739 (N_10739,N_10596,N_10605);
and U10740 (N_10740,N_10512,N_10585);
xor U10741 (N_10741,N_10580,N_10581);
and U10742 (N_10742,N_10562,N_10555);
xor U10743 (N_10743,N_10624,N_10511);
xor U10744 (N_10744,N_10615,N_10596);
or U10745 (N_10745,N_10602,N_10597);
xnor U10746 (N_10746,N_10517,N_10602);
nor U10747 (N_10747,N_10579,N_10622);
or U10748 (N_10748,N_10581,N_10507);
nor U10749 (N_10749,N_10511,N_10502);
and U10750 (N_10750,N_10727,N_10693);
or U10751 (N_10751,N_10655,N_10731);
xnor U10752 (N_10752,N_10742,N_10637);
xor U10753 (N_10753,N_10721,N_10636);
nand U10754 (N_10754,N_10642,N_10625);
or U10755 (N_10755,N_10639,N_10699);
nor U10756 (N_10756,N_10681,N_10658);
and U10757 (N_10757,N_10669,N_10653);
or U10758 (N_10758,N_10654,N_10712);
and U10759 (N_10759,N_10703,N_10735);
or U10760 (N_10760,N_10663,N_10733);
xor U10761 (N_10761,N_10747,N_10729);
nand U10762 (N_10762,N_10738,N_10662);
or U10763 (N_10763,N_10652,N_10661);
and U10764 (N_10764,N_10726,N_10660);
and U10765 (N_10765,N_10723,N_10626);
and U10766 (N_10766,N_10667,N_10666);
or U10767 (N_10767,N_10691,N_10739);
xor U10768 (N_10768,N_10675,N_10629);
nand U10769 (N_10769,N_10685,N_10734);
nor U10770 (N_10770,N_10670,N_10646);
or U10771 (N_10771,N_10705,N_10640);
xor U10772 (N_10772,N_10746,N_10635);
or U10773 (N_10773,N_10745,N_10722);
xor U10774 (N_10774,N_10680,N_10668);
nand U10775 (N_10775,N_10704,N_10673);
and U10776 (N_10776,N_10650,N_10744);
nand U10777 (N_10777,N_10695,N_10730);
and U10778 (N_10778,N_10719,N_10737);
nor U10779 (N_10779,N_10716,N_10686);
and U10780 (N_10780,N_10725,N_10720);
nor U10781 (N_10781,N_10656,N_10678);
nor U10782 (N_10782,N_10664,N_10740);
nor U10783 (N_10783,N_10702,N_10648);
and U10784 (N_10784,N_10694,N_10707);
nor U10785 (N_10785,N_10687,N_10713);
and U10786 (N_10786,N_10676,N_10748);
and U10787 (N_10787,N_10647,N_10645);
xnor U10788 (N_10788,N_10711,N_10672);
nor U10789 (N_10789,N_10659,N_10628);
or U10790 (N_10790,N_10697,N_10732);
or U10791 (N_10791,N_10706,N_10715);
nand U10792 (N_10792,N_10728,N_10714);
xnor U10793 (N_10793,N_10651,N_10741);
or U10794 (N_10794,N_10633,N_10709);
or U10795 (N_10795,N_10708,N_10690);
or U10796 (N_10796,N_10698,N_10688);
or U10797 (N_10797,N_10684,N_10677);
xnor U10798 (N_10798,N_10718,N_10671);
nor U10799 (N_10799,N_10692,N_10717);
or U10800 (N_10800,N_10641,N_10736);
nor U10801 (N_10801,N_10749,N_10657);
nor U10802 (N_10802,N_10683,N_10631);
nor U10803 (N_10803,N_10665,N_10643);
and U10804 (N_10804,N_10724,N_10743);
nand U10805 (N_10805,N_10630,N_10638);
or U10806 (N_10806,N_10679,N_10674);
nor U10807 (N_10807,N_10644,N_10710);
xor U10808 (N_10808,N_10689,N_10696);
and U10809 (N_10809,N_10701,N_10634);
and U10810 (N_10810,N_10649,N_10632);
nor U10811 (N_10811,N_10627,N_10700);
nor U10812 (N_10812,N_10682,N_10739);
nor U10813 (N_10813,N_10736,N_10658);
xor U10814 (N_10814,N_10647,N_10660);
nor U10815 (N_10815,N_10679,N_10632);
xnor U10816 (N_10816,N_10715,N_10720);
nor U10817 (N_10817,N_10713,N_10700);
nand U10818 (N_10818,N_10691,N_10698);
nor U10819 (N_10819,N_10699,N_10682);
nand U10820 (N_10820,N_10666,N_10649);
nand U10821 (N_10821,N_10698,N_10749);
nand U10822 (N_10822,N_10716,N_10673);
nor U10823 (N_10823,N_10648,N_10643);
nand U10824 (N_10824,N_10693,N_10749);
or U10825 (N_10825,N_10734,N_10729);
xnor U10826 (N_10826,N_10691,N_10740);
nor U10827 (N_10827,N_10732,N_10645);
xor U10828 (N_10828,N_10727,N_10747);
nor U10829 (N_10829,N_10663,N_10684);
and U10830 (N_10830,N_10738,N_10663);
nand U10831 (N_10831,N_10738,N_10641);
nand U10832 (N_10832,N_10652,N_10724);
or U10833 (N_10833,N_10718,N_10731);
or U10834 (N_10834,N_10679,N_10640);
and U10835 (N_10835,N_10727,N_10733);
or U10836 (N_10836,N_10700,N_10639);
nand U10837 (N_10837,N_10698,N_10635);
xnor U10838 (N_10838,N_10699,N_10638);
and U10839 (N_10839,N_10628,N_10633);
and U10840 (N_10840,N_10661,N_10708);
nand U10841 (N_10841,N_10737,N_10715);
or U10842 (N_10842,N_10652,N_10743);
and U10843 (N_10843,N_10706,N_10722);
and U10844 (N_10844,N_10718,N_10685);
and U10845 (N_10845,N_10679,N_10697);
or U10846 (N_10846,N_10718,N_10724);
xor U10847 (N_10847,N_10731,N_10688);
nor U10848 (N_10848,N_10736,N_10744);
and U10849 (N_10849,N_10708,N_10743);
xor U10850 (N_10850,N_10629,N_10734);
or U10851 (N_10851,N_10643,N_10636);
nor U10852 (N_10852,N_10631,N_10744);
and U10853 (N_10853,N_10681,N_10647);
xnor U10854 (N_10854,N_10651,N_10705);
and U10855 (N_10855,N_10723,N_10740);
nor U10856 (N_10856,N_10653,N_10637);
and U10857 (N_10857,N_10647,N_10686);
nand U10858 (N_10858,N_10698,N_10628);
xor U10859 (N_10859,N_10742,N_10651);
nand U10860 (N_10860,N_10728,N_10639);
or U10861 (N_10861,N_10684,N_10727);
xor U10862 (N_10862,N_10680,N_10684);
nand U10863 (N_10863,N_10692,N_10641);
or U10864 (N_10864,N_10677,N_10634);
nand U10865 (N_10865,N_10686,N_10684);
nor U10866 (N_10866,N_10727,N_10709);
or U10867 (N_10867,N_10635,N_10745);
nor U10868 (N_10868,N_10715,N_10697);
nor U10869 (N_10869,N_10742,N_10699);
nor U10870 (N_10870,N_10643,N_10712);
nor U10871 (N_10871,N_10702,N_10644);
or U10872 (N_10872,N_10710,N_10669);
nand U10873 (N_10873,N_10715,N_10674);
nor U10874 (N_10874,N_10723,N_10665);
xor U10875 (N_10875,N_10868,N_10843);
or U10876 (N_10876,N_10783,N_10803);
xnor U10877 (N_10877,N_10802,N_10825);
xnor U10878 (N_10878,N_10821,N_10835);
xor U10879 (N_10879,N_10829,N_10798);
or U10880 (N_10880,N_10832,N_10862);
and U10881 (N_10881,N_10750,N_10861);
xor U10882 (N_10882,N_10845,N_10785);
nor U10883 (N_10883,N_10838,N_10761);
nor U10884 (N_10884,N_10807,N_10859);
nand U10885 (N_10885,N_10782,N_10819);
or U10886 (N_10886,N_10853,N_10813);
xnor U10887 (N_10887,N_10772,N_10799);
or U10888 (N_10888,N_10758,N_10797);
nand U10889 (N_10889,N_10780,N_10834);
xor U10890 (N_10890,N_10786,N_10846);
nand U10891 (N_10891,N_10787,N_10827);
and U10892 (N_10892,N_10765,N_10842);
nand U10893 (N_10893,N_10863,N_10837);
or U10894 (N_10894,N_10823,N_10852);
and U10895 (N_10895,N_10831,N_10800);
nor U10896 (N_10896,N_10828,N_10796);
and U10897 (N_10897,N_10850,N_10849);
xor U10898 (N_10898,N_10820,N_10840);
nor U10899 (N_10899,N_10830,N_10801);
or U10900 (N_10900,N_10779,N_10757);
xnor U10901 (N_10901,N_10767,N_10822);
xor U10902 (N_10902,N_10841,N_10762);
nor U10903 (N_10903,N_10809,N_10826);
and U10904 (N_10904,N_10766,N_10759);
nor U10905 (N_10905,N_10771,N_10760);
xor U10906 (N_10906,N_10773,N_10769);
nand U10907 (N_10907,N_10806,N_10812);
and U10908 (N_10908,N_10789,N_10790);
and U10909 (N_10909,N_10870,N_10858);
or U10910 (N_10910,N_10778,N_10872);
and U10911 (N_10911,N_10781,N_10794);
and U10912 (N_10912,N_10754,N_10763);
or U10913 (N_10913,N_10836,N_10756);
or U10914 (N_10914,N_10815,N_10851);
nand U10915 (N_10915,N_10810,N_10865);
nand U10916 (N_10916,N_10805,N_10874);
nor U10917 (N_10917,N_10777,N_10791);
nand U10918 (N_10918,N_10866,N_10795);
or U10919 (N_10919,N_10864,N_10775);
and U10920 (N_10920,N_10804,N_10788);
and U10921 (N_10921,N_10808,N_10792);
xnor U10922 (N_10922,N_10776,N_10824);
or U10923 (N_10923,N_10774,N_10764);
xor U10924 (N_10924,N_10816,N_10854);
nor U10925 (N_10925,N_10855,N_10784);
or U10926 (N_10926,N_10839,N_10755);
xor U10927 (N_10927,N_10847,N_10856);
and U10928 (N_10928,N_10860,N_10811);
or U10929 (N_10929,N_10814,N_10833);
or U10930 (N_10930,N_10770,N_10817);
nor U10931 (N_10931,N_10848,N_10753);
and U10932 (N_10932,N_10818,N_10844);
nor U10933 (N_10933,N_10857,N_10752);
and U10934 (N_10934,N_10793,N_10869);
xnor U10935 (N_10935,N_10871,N_10873);
nor U10936 (N_10936,N_10751,N_10867);
or U10937 (N_10937,N_10768,N_10847);
nand U10938 (N_10938,N_10832,N_10791);
and U10939 (N_10939,N_10858,N_10785);
nand U10940 (N_10940,N_10836,N_10873);
nand U10941 (N_10941,N_10840,N_10818);
nor U10942 (N_10942,N_10785,N_10754);
nor U10943 (N_10943,N_10862,N_10792);
and U10944 (N_10944,N_10855,N_10791);
xor U10945 (N_10945,N_10840,N_10815);
nor U10946 (N_10946,N_10828,N_10873);
xor U10947 (N_10947,N_10798,N_10776);
and U10948 (N_10948,N_10754,N_10835);
or U10949 (N_10949,N_10822,N_10850);
or U10950 (N_10950,N_10774,N_10841);
nand U10951 (N_10951,N_10807,N_10813);
xor U10952 (N_10952,N_10769,N_10817);
nor U10953 (N_10953,N_10752,N_10761);
nand U10954 (N_10954,N_10771,N_10759);
nand U10955 (N_10955,N_10874,N_10851);
nand U10956 (N_10956,N_10868,N_10762);
nor U10957 (N_10957,N_10839,N_10786);
nor U10958 (N_10958,N_10872,N_10835);
nor U10959 (N_10959,N_10820,N_10836);
or U10960 (N_10960,N_10776,N_10827);
or U10961 (N_10961,N_10867,N_10758);
xnor U10962 (N_10962,N_10832,N_10868);
or U10963 (N_10963,N_10859,N_10842);
and U10964 (N_10964,N_10791,N_10830);
and U10965 (N_10965,N_10835,N_10757);
and U10966 (N_10966,N_10866,N_10817);
xor U10967 (N_10967,N_10751,N_10769);
nand U10968 (N_10968,N_10765,N_10808);
xor U10969 (N_10969,N_10793,N_10809);
nor U10970 (N_10970,N_10783,N_10829);
xor U10971 (N_10971,N_10758,N_10834);
xnor U10972 (N_10972,N_10759,N_10850);
xnor U10973 (N_10973,N_10772,N_10874);
or U10974 (N_10974,N_10813,N_10824);
or U10975 (N_10975,N_10787,N_10806);
nor U10976 (N_10976,N_10803,N_10784);
and U10977 (N_10977,N_10832,N_10783);
xor U10978 (N_10978,N_10821,N_10763);
and U10979 (N_10979,N_10861,N_10829);
or U10980 (N_10980,N_10778,N_10867);
and U10981 (N_10981,N_10863,N_10841);
nor U10982 (N_10982,N_10774,N_10840);
and U10983 (N_10983,N_10780,N_10752);
xnor U10984 (N_10984,N_10810,N_10796);
nor U10985 (N_10985,N_10873,N_10865);
and U10986 (N_10986,N_10770,N_10860);
nand U10987 (N_10987,N_10803,N_10766);
xor U10988 (N_10988,N_10775,N_10788);
or U10989 (N_10989,N_10767,N_10783);
and U10990 (N_10990,N_10871,N_10791);
and U10991 (N_10991,N_10802,N_10797);
nor U10992 (N_10992,N_10847,N_10831);
and U10993 (N_10993,N_10868,N_10789);
nand U10994 (N_10994,N_10854,N_10840);
nor U10995 (N_10995,N_10843,N_10864);
xor U10996 (N_10996,N_10830,N_10822);
or U10997 (N_10997,N_10781,N_10765);
nand U10998 (N_10998,N_10835,N_10826);
xor U10999 (N_10999,N_10867,N_10764);
xor U11000 (N_11000,N_10926,N_10965);
nor U11001 (N_11001,N_10887,N_10913);
and U11002 (N_11002,N_10898,N_10936);
xor U11003 (N_11003,N_10950,N_10877);
xor U11004 (N_11004,N_10984,N_10939);
xor U11005 (N_11005,N_10893,N_10964);
xnor U11006 (N_11006,N_10895,N_10875);
and U11007 (N_11007,N_10907,N_10882);
or U11008 (N_11008,N_10920,N_10906);
xor U11009 (N_11009,N_10916,N_10962);
and U11010 (N_11010,N_10903,N_10971);
and U11011 (N_11011,N_10989,N_10952);
nand U11012 (N_11012,N_10957,N_10929);
xor U11013 (N_11013,N_10998,N_10885);
xnor U11014 (N_11014,N_10992,N_10925);
and U11015 (N_11015,N_10908,N_10986);
nand U11016 (N_11016,N_10892,N_10933);
nor U11017 (N_11017,N_10966,N_10997);
xnor U11018 (N_11018,N_10890,N_10889);
nand U11019 (N_11019,N_10899,N_10960);
nor U11020 (N_11020,N_10937,N_10995);
nand U11021 (N_11021,N_10944,N_10955);
xnor U11022 (N_11022,N_10968,N_10958);
or U11023 (N_11023,N_10987,N_10918);
nand U11024 (N_11024,N_10961,N_10881);
nand U11025 (N_11025,N_10972,N_10981);
and U11026 (N_11026,N_10980,N_10945);
nand U11027 (N_11027,N_10973,N_10967);
nor U11028 (N_11028,N_10910,N_10946);
and U11029 (N_11029,N_10876,N_10923);
nor U11030 (N_11030,N_10879,N_10935);
nand U11031 (N_11031,N_10909,N_10993);
xnor U11032 (N_11032,N_10991,N_10891);
nand U11033 (N_11033,N_10990,N_10896);
nor U11034 (N_11034,N_10915,N_10927);
nor U11035 (N_11035,N_10931,N_10941);
or U11036 (N_11036,N_10996,N_10943);
nand U11037 (N_11037,N_10948,N_10938);
or U11038 (N_11038,N_10983,N_10954);
or U11039 (N_11039,N_10894,N_10884);
xor U11040 (N_11040,N_10963,N_10951);
and U11041 (N_11041,N_10940,N_10977);
nand U11042 (N_11042,N_10928,N_10959);
or U11043 (N_11043,N_10878,N_10999);
xnor U11044 (N_11044,N_10985,N_10947);
nor U11045 (N_11045,N_10974,N_10888);
xor U11046 (N_11046,N_10994,N_10982);
xnor U11047 (N_11047,N_10900,N_10934);
xnor U11048 (N_11048,N_10902,N_10988);
nand U11049 (N_11049,N_10922,N_10904);
nand U11050 (N_11050,N_10975,N_10953);
xnor U11051 (N_11051,N_10921,N_10919);
and U11052 (N_11052,N_10912,N_10978);
or U11053 (N_11053,N_10949,N_10883);
nand U11054 (N_11054,N_10930,N_10924);
or U11055 (N_11055,N_10886,N_10969);
xor U11056 (N_11056,N_10914,N_10905);
and U11057 (N_11057,N_10979,N_10897);
xor U11058 (N_11058,N_10911,N_10932);
and U11059 (N_11059,N_10956,N_10942);
nor U11060 (N_11060,N_10917,N_10976);
nand U11061 (N_11061,N_10880,N_10970);
and U11062 (N_11062,N_10901,N_10984);
and U11063 (N_11063,N_10906,N_10958);
xor U11064 (N_11064,N_10928,N_10884);
or U11065 (N_11065,N_10890,N_10929);
nor U11066 (N_11066,N_10971,N_10907);
xor U11067 (N_11067,N_10939,N_10906);
nand U11068 (N_11068,N_10959,N_10979);
and U11069 (N_11069,N_10883,N_10994);
nand U11070 (N_11070,N_10880,N_10902);
xor U11071 (N_11071,N_10893,N_10948);
xnor U11072 (N_11072,N_10911,N_10987);
xor U11073 (N_11073,N_10982,N_10969);
xor U11074 (N_11074,N_10894,N_10898);
nand U11075 (N_11075,N_10925,N_10981);
xnor U11076 (N_11076,N_10960,N_10953);
xor U11077 (N_11077,N_10957,N_10877);
or U11078 (N_11078,N_10993,N_10881);
nor U11079 (N_11079,N_10903,N_10931);
and U11080 (N_11080,N_10899,N_10957);
or U11081 (N_11081,N_10991,N_10952);
nand U11082 (N_11082,N_10938,N_10937);
nand U11083 (N_11083,N_10900,N_10958);
nor U11084 (N_11084,N_10990,N_10927);
nor U11085 (N_11085,N_10918,N_10919);
nand U11086 (N_11086,N_10906,N_10914);
xor U11087 (N_11087,N_10977,N_10951);
or U11088 (N_11088,N_10984,N_10953);
nand U11089 (N_11089,N_10895,N_10908);
or U11090 (N_11090,N_10885,N_10976);
nor U11091 (N_11091,N_10991,N_10886);
and U11092 (N_11092,N_10985,N_10964);
xnor U11093 (N_11093,N_10980,N_10932);
nor U11094 (N_11094,N_10950,N_10953);
or U11095 (N_11095,N_10945,N_10994);
nand U11096 (N_11096,N_10954,N_10985);
nor U11097 (N_11097,N_10887,N_10996);
nor U11098 (N_11098,N_10902,N_10921);
nand U11099 (N_11099,N_10974,N_10904);
and U11100 (N_11100,N_10977,N_10921);
or U11101 (N_11101,N_10960,N_10951);
or U11102 (N_11102,N_10931,N_10886);
and U11103 (N_11103,N_10890,N_10885);
xnor U11104 (N_11104,N_10927,N_10953);
nor U11105 (N_11105,N_10950,N_10876);
xor U11106 (N_11106,N_10924,N_10991);
xor U11107 (N_11107,N_10939,N_10885);
nand U11108 (N_11108,N_10921,N_10968);
and U11109 (N_11109,N_10901,N_10937);
and U11110 (N_11110,N_10968,N_10989);
nand U11111 (N_11111,N_10887,N_10941);
or U11112 (N_11112,N_10926,N_10906);
xnor U11113 (N_11113,N_10970,N_10919);
or U11114 (N_11114,N_10943,N_10886);
nand U11115 (N_11115,N_10994,N_10893);
nand U11116 (N_11116,N_10950,N_10961);
xnor U11117 (N_11117,N_10983,N_10885);
and U11118 (N_11118,N_10939,N_10883);
nor U11119 (N_11119,N_10908,N_10999);
and U11120 (N_11120,N_10879,N_10976);
or U11121 (N_11121,N_10909,N_10879);
xnor U11122 (N_11122,N_10911,N_10956);
or U11123 (N_11123,N_10968,N_10993);
nand U11124 (N_11124,N_10905,N_10952);
nor U11125 (N_11125,N_11113,N_11086);
nor U11126 (N_11126,N_11093,N_11087);
nand U11127 (N_11127,N_11099,N_11081);
nor U11128 (N_11128,N_11071,N_11123);
or U11129 (N_11129,N_11085,N_11070);
xnor U11130 (N_11130,N_11026,N_11058);
xor U11131 (N_11131,N_11124,N_11032);
and U11132 (N_11132,N_11065,N_11028);
xor U11133 (N_11133,N_11042,N_11013);
xor U11134 (N_11134,N_11056,N_11005);
and U11135 (N_11135,N_11089,N_11035);
xnor U11136 (N_11136,N_11053,N_11030);
nand U11137 (N_11137,N_11074,N_11025);
nor U11138 (N_11138,N_11051,N_11002);
and U11139 (N_11139,N_11061,N_11116);
or U11140 (N_11140,N_11018,N_11069);
nor U11141 (N_11141,N_11041,N_11102);
or U11142 (N_11142,N_11078,N_11082);
and U11143 (N_11143,N_11054,N_11080);
or U11144 (N_11144,N_11077,N_11066);
nand U11145 (N_11145,N_11022,N_11015);
and U11146 (N_11146,N_11055,N_11038);
or U11147 (N_11147,N_11079,N_11118);
or U11148 (N_11148,N_11114,N_11084);
nor U11149 (N_11149,N_11090,N_11039);
nor U11150 (N_11150,N_11046,N_11104);
nand U11151 (N_11151,N_11047,N_11117);
and U11152 (N_11152,N_11036,N_11003);
and U11153 (N_11153,N_11027,N_11006);
nor U11154 (N_11154,N_11064,N_11043);
and U11155 (N_11155,N_11020,N_11050);
or U11156 (N_11156,N_11098,N_11034);
xnor U11157 (N_11157,N_11045,N_11110);
nand U11158 (N_11158,N_11048,N_11115);
or U11159 (N_11159,N_11008,N_11031);
xnor U11160 (N_11160,N_11009,N_11092);
nand U11161 (N_11161,N_11122,N_11109);
nor U11162 (N_11162,N_11068,N_11108);
xor U11163 (N_11163,N_11059,N_11121);
or U11164 (N_11164,N_11057,N_11021);
xnor U11165 (N_11165,N_11040,N_11052);
nor U11166 (N_11166,N_11111,N_11010);
and U11167 (N_11167,N_11103,N_11073);
or U11168 (N_11168,N_11100,N_11094);
nor U11169 (N_11169,N_11017,N_11000);
nor U11170 (N_11170,N_11105,N_11095);
or U11171 (N_11171,N_11019,N_11007);
xnor U11172 (N_11172,N_11011,N_11049);
and U11173 (N_11173,N_11067,N_11088);
and U11174 (N_11174,N_11107,N_11091);
xor U11175 (N_11175,N_11033,N_11037);
nor U11176 (N_11176,N_11072,N_11023);
xor U11177 (N_11177,N_11004,N_11106);
or U11178 (N_11178,N_11112,N_11083);
nand U11179 (N_11179,N_11014,N_11101);
or U11180 (N_11180,N_11075,N_11120);
nor U11181 (N_11181,N_11096,N_11016);
xnor U11182 (N_11182,N_11060,N_11063);
or U11183 (N_11183,N_11119,N_11076);
nor U11184 (N_11184,N_11044,N_11001);
nor U11185 (N_11185,N_11062,N_11024);
nor U11186 (N_11186,N_11029,N_11012);
or U11187 (N_11187,N_11097,N_11102);
and U11188 (N_11188,N_11030,N_11079);
xor U11189 (N_11189,N_11021,N_11118);
nor U11190 (N_11190,N_11112,N_11079);
and U11191 (N_11191,N_11081,N_11048);
nor U11192 (N_11192,N_11047,N_11019);
nand U11193 (N_11193,N_11045,N_11118);
nor U11194 (N_11194,N_11011,N_11089);
and U11195 (N_11195,N_11008,N_11046);
nand U11196 (N_11196,N_11118,N_11049);
or U11197 (N_11197,N_11075,N_11005);
nor U11198 (N_11198,N_11065,N_11039);
or U11199 (N_11199,N_11049,N_11065);
nand U11200 (N_11200,N_11074,N_11110);
nand U11201 (N_11201,N_11088,N_11022);
nor U11202 (N_11202,N_11035,N_11107);
nor U11203 (N_11203,N_11029,N_11118);
or U11204 (N_11204,N_11061,N_11047);
xnor U11205 (N_11205,N_11000,N_11063);
or U11206 (N_11206,N_11063,N_11094);
and U11207 (N_11207,N_11025,N_11088);
or U11208 (N_11208,N_11001,N_11057);
nor U11209 (N_11209,N_11095,N_11119);
nor U11210 (N_11210,N_11060,N_11029);
xor U11211 (N_11211,N_11083,N_11056);
nand U11212 (N_11212,N_11006,N_11083);
or U11213 (N_11213,N_11032,N_11112);
nand U11214 (N_11214,N_11022,N_11117);
xnor U11215 (N_11215,N_11006,N_11063);
xnor U11216 (N_11216,N_11078,N_11071);
or U11217 (N_11217,N_11051,N_11081);
nor U11218 (N_11218,N_11096,N_11077);
nand U11219 (N_11219,N_11031,N_11087);
nor U11220 (N_11220,N_11099,N_11051);
xor U11221 (N_11221,N_11030,N_11021);
xor U11222 (N_11222,N_11098,N_11069);
nand U11223 (N_11223,N_11020,N_11093);
xnor U11224 (N_11224,N_11021,N_11076);
and U11225 (N_11225,N_11044,N_11115);
nor U11226 (N_11226,N_11114,N_11093);
nor U11227 (N_11227,N_11078,N_11000);
nand U11228 (N_11228,N_11037,N_11051);
nand U11229 (N_11229,N_11077,N_11116);
or U11230 (N_11230,N_11035,N_11097);
nand U11231 (N_11231,N_11049,N_11054);
xnor U11232 (N_11232,N_11062,N_11090);
xnor U11233 (N_11233,N_11023,N_11015);
or U11234 (N_11234,N_11111,N_11107);
nor U11235 (N_11235,N_11121,N_11019);
xnor U11236 (N_11236,N_11105,N_11025);
or U11237 (N_11237,N_11116,N_11071);
xor U11238 (N_11238,N_11037,N_11042);
xor U11239 (N_11239,N_11022,N_11073);
nand U11240 (N_11240,N_11027,N_11079);
nand U11241 (N_11241,N_11046,N_11025);
and U11242 (N_11242,N_11071,N_11090);
nor U11243 (N_11243,N_11118,N_11120);
xor U11244 (N_11244,N_11058,N_11069);
xor U11245 (N_11245,N_11052,N_11043);
nand U11246 (N_11246,N_11086,N_11100);
or U11247 (N_11247,N_11059,N_11002);
and U11248 (N_11248,N_11086,N_11112);
and U11249 (N_11249,N_11056,N_11089);
nor U11250 (N_11250,N_11129,N_11153);
xnor U11251 (N_11251,N_11248,N_11159);
nor U11252 (N_11252,N_11240,N_11191);
or U11253 (N_11253,N_11221,N_11199);
xnor U11254 (N_11254,N_11242,N_11176);
xor U11255 (N_11255,N_11128,N_11198);
nor U11256 (N_11256,N_11212,N_11226);
nor U11257 (N_11257,N_11234,N_11203);
nand U11258 (N_11258,N_11136,N_11138);
or U11259 (N_11259,N_11205,N_11151);
and U11260 (N_11260,N_11246,N_11243);
nor U11261 (N_11261,N_11141,N_11161);
and U11262 (N_11262,N_11180,N_11170);
nor U11263 (N_11263,N_11204,N_11225);
nand U11264 (N_11264,N_11183,N_11163);
nor U11265 (N_11265,N_11168,N_11201);
and U11266 (N_11266,N_11171,N_11166);
and U11267 (N_11267,N_11185,N_11134);
xor U11268 (N_11268,N_11233,N_11137);
or U11269 (N_11269,N_11175,N_11218);
and U11270 (N_11270,N_11144,N_11178);
nor U11271 (N_11271,N_11164,N_11239);
or U11272 (N_11272,N_11238,N_11214);
nand U11273 (N_11273,N_11209,N_11192);
and U11274 (N_11274,N_11177,N_11152);
xnor U11275 (N_11275,N_11142,N_11208);
nand U11276 (N_11276,N_11145,N_11135);
and U11277 (N_11277,N_11206,N_11179);
nor U11278 (N_11278,N_11229,N_11162);
nor U11279 (N_11279,N_11130,N_11143);
nand U11280 (N_11280,N_11196,N_11236);
xnor U11281 (N_11281,N_11244,N_11186);
nand U11282 (N_11282,N_11247,N_11169);
nor U11283 (N_11283,N_11182,N_11193);
or U11284 (N_11284,N_11202,N_11184);
and U11285 (N_11285,N_11217,N_11207);
xor U11286 (N_11286,N_11227,N_11222);
nor U11287 (N_11287,N_11140,N_11150);
or U11288 (N_11288,N_11132,N_11173);
or U11289 (N_11289,N_11165,N_11228);
nand U11290 (N_11290,N_11197,N_11219);
nand U11291 (N_11291,N_11149,N_11213);
and U11292 (N_11292,N_11126,N_11223);
nand U11293 (N_11293,N_11232,N_11160);
and U11294 (N_11294,N_11154,N_11133);
or U11295 (N_11295,N_11181,N_11200);
xor U11296 (N_11296,N_11230,N_11156);
nand U11297 (N_11297,N_11245,N_11210);
nand U11298 (N_11298,N_11216,N_11188);
xnor U11299 (N_11299,N_11215,N_11155);
and U11300 (N_11300,N_11220,N_11158);
nor U11301 (N_11301,N_11194,N_11189);
nor U11302 (N_11302,N_11125,N_11174);
xor U11303 (N_11303,N_11147,N_11235);
nor U11304 (N_11304,N_11241,N_11131);
nand U11305 (N_11305,N_11190,N_11195);
nand U11306 (N_11306,N_11167,N_11237);
or U11307 (N_11307,N_11127,N_11139);
or U11308 (N_11308,N_11148,N_11157);
or U11309 (N_11309,N_11211,N_11146);
and U11310 (N_11310,N_11172,N_11231);
nor U11311 (N_11311,N_11224,N_11249);
xor U11312 (N_11312,N_11187,N_11151);
or U11313 (N_11313,N_11223,N_11213);
xnor U11314 (N_11314,N_11216,N_11211);
nor U11315 (N_11315,N_11138,N_11165);
nor U11316 (N_11316,N_11142,N_11135);
and U11317 (N_11317,N_11132,N_11138);
and U11318 (N_11318,N_11227,N_11190);
nand U11319 (N_11319,N_11196,N_11158);
xnor U11320 (N_11320,N_11177,N_11185);
xnor U11321 (N_11321,N_11170,N_11247);
or U11322 (N_11322,N_11134,N_11247);
or U11323 (N_11323,N_11227,N_11196);
xor U11324 (N_11324,N_11208,N_11235);
xnor U11325 (N_11325,N_11157,N_11132);
or U11326 (N_11326,N_11181,N_11136);
or U11327 (N_11327,N_11146,N_11173);
xnor U11328 (N_11328,N_11220,N_11147);
xnor U11329 (N_11329,N_11176,N_11164);
xnor U11330 (N_11330,N_11229,N_11246);
and U11331 (N_11331,N_11169,N_11126);
or U11332 (N_11332,N_11162,N_11218);
and U11333 (N_11333,N_11244,N_11245);
or U11334 (N_11334,N_11182,N_11149);
and U11335 (N_11335,N_11184,N_11191);
and U11336 (N_11336,N_11160,N_11208);
nand U11337 (N_11337,N_11198,N_11160);
nor U11338 (N_11338,N_11183,N_11153);
nand U11339 (N_11339,N_11193,N_11153);
xnor U11340 (N_11340,N_11146,N_11153);
xor U11341 (N_11341,N_11154,N_11168);
xor U11342 (N_11342,N_11149,N_11134);
nor U11343 (N_11343,N_11198,N_11199);
nor U11344 (N_11344,N_11234,N_11147);
nor U11345 (N_11345,N_11203,N_11226);
and U11346 (N_11346,N_11133,N_11159);
nor U11347 (N_11347,N_11236,N_11160);
nor U11348 (N_11348,N_11212,N_11204);
xnor U11349 (N_11349,N_11227,N_11225);
nor U11350 (N_11350,N_11163,N_11164);
and U11351 (N_11351,N_11226,N_11132);
xor U11352 (N_11352,N_11156,N_11205);
or U11353 (N_11353,N_11194,N_11211);
and U11354 (N_11354,N_11240,N_11170);
nand U11355 (N_11355,N_11151,N_11242);
nor U11356 (N_11356,N_11177,N_11170);
and U11357 (N_11357,N_11243,N_11207);
xor U11358 (N_11358,N_11132,N_11206);
or U11359 (N_11359,N_11160,N_11219);
xnor U11360 (N_11360,N_11231,N_11141);
nand U11361 (N_11361,N_11154,N_11163);
nand U11362 (N_11362,N_11194,N_11135);
nor U11363 (N_11363,N_11230,N_11245);
or U11364 (N_11364,N_11165,N_11196);
xnor U11365 (N_11365,N_11188,N_11192);
or U11366 (N_11366,N_11164,N_11137);
nand U11367 (N_11367,N_11189,N_11244);
nor U11368 (N_11368,N_11142,N_11236);
nor U11369 (N_11369,N_11209,N_11198);
nor U11370 (N_11370,N_11170,N_11215);
nand U11371 (N_11371,N_11138,N_11245);
nand U11372 (N_11372,N_11212,N_11203);
xor U11373 (N_11373,N_11171,N_11192);
and U11374 (N_11374,N_11195,N_11196);
and U11375 (N_11375,N_11280,N_11254);
or U11376 (N_11376,N_11264,N_11327);
or U11377 (N_11377,N_11357,N_11286);
nand U11378 (N_11378,N_11257,N_11367);
or U11379 (N_11379,N_11340,N_11322);
nor U11380 (N_11380,N_11373,N_11360);
nor U11381 (N_11381,N_11290,N_11291);
xor U11382 (N_11382,N_11362,N_11354);
nor U11383 (N_11383,N_11301,N_11266);
or U11384 (N_11384,N_11253,N_11273);
and U11385 (N_11385,N_11331,N_11293);
nor U11386 (N_11386,N_11368,N_11258);
xor U11387 (N_11387,N_11259,N_11268);
or U11388 (N_11388,N_11316,N_11256);
xor U11389 (N_11389,N_11308,N_11363);
nand U11390 (N_11390,N_11370,N_11343);
and U11391 (N_11391,N_11319,N_11346);
nor U11392 (N_11392,N_11282,N_11279);
xor U11393 (N_11393,N_11277,N_11332);
and U11394 (N_11394,N_11295,N_11355);
or U11395 (N_11395,N_11260,N_11315);
nand U11396 (N_11396,N_11339,N_11285);
nor U11397 (N_11397,N_11314,N_11321);
nand U11398 (N_11398,N_11338,N_11281);
nand U11399 (N_11399,N_11313,N_11278);
xor U11400 (N_11400,N_11250,N_11329);
nand U11401 (N_11401,N_11265,N_11305);
and U11402 (N_11402,N_11296,N_11270);
and U11403 (N_11403,N_11302,N_11311);
or U11404 (N_11404,N_11334,N_11267);
nor U11405 (N_11405,N_11274,N_11261);
nor U11406 (N_11406,N_11304,N_11317);
and U11407 (N_11407,N_11349,N_11287);
and U11408 (N_11408,N_11288,N_11312);
and U11409 (N_11409,N_11365,N_11283);
nand U11410 (N_11410,N_11325,N_11252);
nor U11411 (N_11411,N_11352,N_11297);
or U11412 (N_11412,N_11372,N_11310);
or U11413 (N_11413,N_11272,N_11276);
and U11414 (N_11414,N_11348,N_11347);
nor U11415 (N_11415,N_11309,N_11262);
nand U11416 (N_11416,N_11275,N_11371);
nand U11417 (N_11417,N_11366,N_11337);
nor U11418 (N_11418,N_11361,N_11263);
and U11419 (N_11419,N_11328,N_11289);
nand U11420 (N_11420,N_11251,N_11345);
and U11421 (N_11421,N_11298,N_11323);
and U11422 (N_11422,N_11374,N_11351);
xor U11423 (N_11423,N_11306,N_11303);
xor U11424 (N_11424,N_11294,N_11356);
nor U11425 (N_11425,N_11284,N_11255);
nor U11426 (N_11426,N_11341,N_11364);
and U11427 (N_11427,N_11359,N_11300);
nor U11428 (N_11428,N_11292,N_11320);
nor U11429 (N_11429,N_11350,N_11358);
nand U11430 (N_11430,N_11335,N_11369);
xor U11431 (N_11431,N_11330,N_11326);
or U11432 (N_11432,N_11307,N_11269);
or U11433 (N_11433,N_11299,N_11344);
and U11434 (N_11434,N_11318,N_11271);
xnor U11435 (N_11435,N_11324,N_11353);
or U11436 (N_11436,N_11333,N_11342);
nand U11437 (N_11437,N_11336,N_11353);
nand U11438 (N_11438,N_11292,N_11293);
nor U11439 (N_11439,N_11334,N_11264);
nand U11440 (N_11440,N_11281,N_11310);
or U11441 (N_11441,N_11315,N_11356);
and U11442 (N_11442,N_11363,N_11361);
nor U11443 (N_11443,N_11361,N_11279);
nand U11444 (N_11444,N_11268,N_11333);
nand U11445 (N_11445,N_11347,N_11268);
nor U11446 (N_11446,N_11318,N_11332);
or U11447 (N_11447,N_11325,N_11265);
nor U11448 (N_11448,N_11276,N_11306);
and U11449 (N_11449,N_11289,N_11357);
nor U11450 (N_11450,N_11307,N_11253);
or U11451 (N_11451,N_11358,N_11297);
nand U11452 (N_11452,N_11339,N_11367);
xor U11453 (N_11453,N_11336,N_11371);
nor U11454 (N_11454,N_11364,N_11367);
or U11455 (N_11455,N_11319,N_11328);
and U11456 (N_11456,N_11373,N_11266);
nand U11457 (N_11457,N_11334,N_11268);
nor U11458 (N_11458,N_11302,N_11288);
and U11459 (N_11459,N_11368,N_11293);
nand U11460 (N_11460,N_11297,N_11262);
nand U11461 (N_11461,N_11253,N_11328);
or U11462 (N_11462,N_11260,N_11348);
xnor U11463 (N_11463,N_11355,N_11256);
and U11464 (N_11464,N_11373,N_11262);
and U11465 (N_11465,N_11252,N_11267);
nand U11466 (N_11466,N_11317,N_11322);
nand U11467 (N_11467,N_11271,N_11329);
and U11468 (N_11468,N_11257,N_11360);
nor U11469 (N_11469,N_11368,N_11283);
nor U11470 (N_11470,N_11373,N_11253);
nand U11471 (N_11471,N_11327,N_11325);
nor U11472 (N_11472,N_11351,N_11260);
nand U11473 (N_11473,N_11309,N_11266);
xnor U11474 (N_11474,N_11300,N_11256);
or U11475 (N_11475,N_11255,N_11350);
and U11476 (N_11476,N_11337,N_11356);
or U11477 (N_11477,N_11313,N_11272);
nand U11478 (N_11478,N_11358,N_11271);
or U11479 (N_11479,N_11266,N_11348);
xnor U11480 (N_11480,N_11351,N_11252);
and U11481 (N_11481,N_11296,N_11339);
xnor U11482 (N_11482,N_11272,N_11296);
or U11483 (N_11483,N_11257,N_11336);
nand U11484 (N_11484,N_11263,N_11286);
xnor U11485 (N_11485,N_11353,N_11335);
and U11486 (N_11486,N_11288,N_11309);
xor U11487 (N_11487,N_11272,N_11261);
nand U11488 (N_11488,N_11292,N_11281);
nor U11489 (N_11489,N_11350,N_11353);
or U11490 (N_11490,N_11335,N_11312);
nor U11491 (N_11491,N_11343,N_11314);
or U11492 (N_11492,N_11374,N_11372);
xnor U11493 (N_11493,N_11300,N_11326);
and U11494 (N_11494,N_11261,N_11313);
nand U11495 (N_11495,N_11339,N_11320);
xor U11496 (N_11496,N_11291,N_11254);
and U11497 (N_11497,N_11325,N_11273);
nor U11498 (N_11498,N_11295,N_11323);
nand U11499 (N_11499,N_11250,N_11314);
nand U11500 (N_11500,N_11442,N_11427);
or U11501 (N_11501,N_11447,N_11418);
nand U11502 (N_11502,N_11429,N_11379);
nand U11503 (N_11503,N_11496,N_11397);
or U11504 (N_11504,N_11382,N_11398);
xor U11505 (N_11505,N_11487,N_11431);
or U11506 (N_11506,N_11482,N_11473);
nand U11507 (N_11507,N_11445,N_11448);
nand U11508 (N_11508,N_11444,N_11396);
nand U11509 (N_11509,N_11404,N_11395);
xor U11510 (N_11510,N_11381,N_11462);
nand U11511 (N_11511,N_11416,N_11423);
xnor U11512 (N_11512,N_11394,N_11459);
and U11513 (N_11513,N_11375,N_11483);
nor U11514 (N_11514,N_11426,N_11497);
nor U11515 (N_11515,N_11475,N_11468);
xor U11516 (N_11516,N_11490,N_11452);
nand U11517 (N_11517,N_11408,N_11386);
xnor U11518 (N_11518,N_11390,N_11485);
nor U11519 (N_11519,N_11453,N_11493);
nor U11520 (N_11520,N_11410,N_11432);
and U11521 (N_11521,N_11474,N_11441);
xor U11522 (N_11522,N_11480,N_11455);
nand U11523 (N_11523,N_11392,N_11383);
or U11524 (N_11524,N_11457,N_11466);
nor U11525 (N_11525,N_11405,N_11385);
nand U11526 (N_11526,N_11436,N_11389);
or U11527 (N_11527,N_11451,N_11401);
and U11528 (N_11528,N_11478,N_11495);
nand U11529 (N_11529,N_11489,N_11486);
or U11530 (N_11530,N_11471,N_11402);
and U11531 (N_11531,N_11417,N_11461);
xor U11532 (N_11532,N_11440,N_11422);
or U11533 (N_11533,N_11454,N_11492);
or U11534 (N_11534,N_11477,N_11449);
and U11535 (N_11535,N_11443,N_11469);
nor U11536 (N_11536,N_11433,N_11494);
nand U11537 (N_11537,N_11463,N_11428);
or U11538 (N_11538,N_11446,N_11470);
or U11539 (N_11539,N_11450,N_11488);
and U11540 (N_11540,N_11491,N_11465);
nand U11541 (N_11541,N_11484,N_11403);
nand U11542 (N_11542,N_11499,N_11380);
nand U11543 (N_11543,N_11407,N_11435);
nand U11544 (N_11544,N_11476,N_11388);
xor U11545 (N_11545,N_11414,N_11387);
or U11546 (N_11546,N_11393,N_11399);
xnor U11547 (N_11547,N_11439,N_11498);
and U11548 (N_11548,N_11434,N_11481);
nor U11549 (N_11549,N_11424,N_11409);
nor U11550 (N_11550,N_11458,N_11467);
nor U11551 (N_11551,N_11391,N_11400);
nand U11552 (N_11552,N_11415,N_11384);
and U11553 (N_11553,N_11413,N_11378);
and U11554 (N_11554,N_11460,N_11377);
nor U11555 (N_11555,N_11411,N_11421);
xnor U11556 (N_11556,N_11464,N_11406);
xnor U11557 (N_11557,N_11479,N_11425);
or U11558 (N_11558,N_11419,N_11437);
xor U11559 (N_11559,N_11412,N_11438);
xnor U11560 (N_11560,N_11420,N_11430);
xnor U11561 (N_11561,N_11456,N_11472);
or U11562 (N_11562,N_11376,N_11472);
nand U11563 (N_11563,N_11488,N_11415);
or U11564 (N_11564,N_11403,N_11467);
nor U11565 (N_11565,N_11423,N_11392);
and U11566 (N_11566,N_11426,N_11455);
xnor U11567 (N_11567,N_11415,N_11452);
xor U11568 (N_11568,N_11411,N_11388);
nand U11569 (N_11569,N_11408,N_11441);
xor U11570 (N_11570,N_11442,N_11458);
or U11571 (N_11571,N_11401,N_11436);
nand U11572 (N_11572,N_11471,N_11481);
and U11573 (N_11573,N_11488,N_11408);
and U11574 (N_11574,N_11384,N_11455);
and U11575 (N_11575,N_11409,N_11390);
and U11576 (N_11576,N_11411,N_11401);
xnor U11577 (N_11577,N_11385,N_11377);
or U11578 (N_11578,N_11380,N_11400);
and U11579 (N_11579,N_11379,N_11470);
and U11580 (N_11580,N_11443,N_11426);
or U11581 (N_11581,N_11455,N_11399);
and U11582 (N_11582,N_11431,N_11399);
nor U11583 (N_11583,N_11440,N_11418);
nand U11584 (N_11584,N_11427,N_11464);
or U11585 (N_11585,N_11427,N_11389);
nor U11586 (N_11586,N_11468,N_11431);
or U11587 (N_11587,N_11490,N_11461);
and U11588 (N_11588,N_11392,N_11499);
xnor U11589 (N_11589,N_11428,N_11424);
nand U11590 (N_11590,N_11468,N_11411);
or U11591 (N_11591,N_11413,N_11407);
nand U11592 (N_11592,N_11488,N_11478);
nor U11593 (N_11593,N_11416,N_11448);
or U11594 (N_11594,N_11418,N_11469);
and U11595 (N_11595,N_11381,N_11457);
nor U11596 (N_11596,N_11480,N_11419);
nor U11597 (N_11597,N_11422,N_11498);
and U11598 (N_11598,N_11433,N_11390);
nand U11599 (N_11599,N_11487,N_11465);
nand U11600 (N_11600,N_11375,N_11455);
nor U11601 (N_11601,N_11387,N_11389);
nand U11602 (N_11602,N_11465,N_11375);
nor U11603 (N_11603,N_11386,N_11498);
nor U11604 (N_11604,N_11483,N_11383);
xor U11605 (N_11605,N_11443,N_11452);
nor U11606 (N_11606,N_11495,N_11491);
and U11607 (N_11607,N_11421,N_11425);
or U11608 (N_11608,N_11460,N_11470);
nor U11609 (N_11609,N_11403,N_11456);
and U11610 (N_11610,N_11379,N_11475);
nor U11611 (N_11611,N_11400,N_11402);
nor U11612 (N_11612,N_11461,N_11484);
nand U11613 (N_11613,N_11388,N_11460);
nand U11614 (N_11614,N_11416,N_11489);
or U11615 (N_11615,N_11454,N_11447);
nand U11616 (N_11616,N_11415,N_11419);
and U11617 (N_11617,N_11488,N_11496);
xor U11618 (N_11618,N_11427,N_11497);
nand U11619 (N_11619,N_11410,N_11417);
nand U11620 (N_11620,N_11474,N_11478);
and U11621 (N_11621,N_11435,N_11466);
nor U11622 (N_11622,N_11489,N_11456);
xor U11623 (N_11623,N_11417,N_11406);
or U11624 (N_11624,N_11487,N_11401);
or U11625 (N_11625,N_11505,N_11513);
and U11626 (N_11626,N_11564,N_11538);
or U11627 (N_11627,N_11587,N_11574);
nand U11628 (N_11628,N_11595,N_11544);
and U11629 (N_11629,N_11549,N_11583);
nand U11630 (N_11630,N_11581,N_11525);
xor U11631 (N_11631,N_11591,N_11559);
or U11632 (N_11632,N_11576,N_11558);
nand U11633 (N_11633,N_11511,N_11611);
xor U11634 (N_11634,N_11590,N_11605);
nand U11635 (N_11635,N_11579,N_11596);
nand U11636 (N_11636,N_11504,N_11537);
or U11637 (N_11637,N_11589,N_11506);
or U11638 (N_11638,N_11528,N_11569);
xor U11639 (N_11639,N_11602,N_11593);
xor U11640 (N_11640,N_11586,N_11550);
xor U11641 (N_11641,N_11619,N_11568);
and U11642 (N_11642,N_11536,N_11571);
nand U11643 (N_11643,N_11609,N_11530);
xor U11644 (N_11644,N_11557,N_11577);
xor U11645 (N_11645,N_11523,N_11603);
nor U11646 (N_11646,N_11510,N_11514);
nand U11647 (N_11647,N_11612,N_11507);
xor U11648 (N_11648,N_11500,N_11545);
nand U11649 (N_11649,N_11565,N_11524);
nand U11650 (N_11650,N_11582,N_11508);
or U11651 (N_11651,N_11526,N_11618);
or U11652 (N_11652,N_11624,N_11599);
nand U11653 (N_11653,N_11515,N_11570);
or U11654 (N_11654,N_11563,N_11533);
xnor U11655 (N_11655,N_11501,N_11518);
and U11656 (N_11656,N_11512,N_11584);
and U11657 (N_11657,N_11592,N_11607);
nand U11658 (N_11658,N_11585,N_11621);
nor U11659 (N_11659,N_11555,N_11623);
or U11660 (N_11660,N_11617,N_11532);
and U11661 (N_11661,N_11604,N_11541);
or U11662 (N_11662,N_11552,N_11553);
xor U11663 (N_11663,N_11519,N_11503);
nand U11664 (N_11664,N_11598,N_11542);
xor U11665 (N_11665,N_11572,N_11551);
and U11666 (N_11666,N_11560,N_11548);
nor U11667 (N_11667,N_11535,N_11562);
nor U11668 (N_11668,N_11588,N_11554);
nand U11669 (N_11669,N_11622,N_11522);
and U11670 (N_11670,N_11580,N_11516);
or U11671 (N_11671,N_11567,N_11600);
and U11672 (N_11672,N_11546,N_11502);
or U11673 (N_11673,N_11527,N_11597);
and U11674 (N_11674,N_11575,N_11531);
or U11675 (N_11675,N_11616,N_11517);
nand U11676 (N_11676,N_11534,N_11613);
nor U11677 (N_11677,N_11556,N_11615);
nand U11678 (N_11678,N_11594,N_11529);
nor U11679 (N_11679,N_11614,N_11606);
nand U11680 (N_11680,N_11608,N_11573);
nor U11681 (N_11681,N_11578,N_11610);
and U11682 (N_11682,N_11520,N_11561);
nand U11683 (N_11683,N_11543,N_11620);
and U11684 (N_11684,N_11601,N_11540);
nor U11685 (N_11685,N_11509,N_11521);
or U11686 (N_11686,N_11547,N_11566);
nand U11687 (N_11687,N_11539,N_11588);
and U11688 (N_11688,N_11512,N_11608);
nor U11689 (N_11689,N_11537,N_11553);
and U11690 (N_11690,N_11597,N_11501);
and U11691 (N_11691,N_11593,N_11599);
nand U11692 (N_11692,N_11521,N_11549);
nor U11693 (N_11693,N_11512,N_11528);
nor U11694 (N_11694,N_11501,N_11623);
and U11695 (N_11695,N_11581,N_11503);
nand U11696 (N_11696,N_11509,N_11604);
xnor U11697 (N_11697,N_11562,N_11615);
and U11698 (N_11698,N_11567,N_11560);
nand U11699 (N_11699,N_11541,N_11596);
nand U11700 (N_11700,N_11555,N_11503);
nor U11701 (N_11701,N_11619,N_11581);
nand U11702 (N_11702,N_11540,N_11594);
xor U11703 (N_11703,N_11519,N_11588);
and U11704 (N_11704,N_11514,N_11529);
nand U11705 (N_11705,N_11530,N_11596);
nor U11706 (N_11706,N_11525,N_11504);
and U11707 (N_11707,N_11587,N_11597);
xnor U11708 (N_11708,N_11523,N_11568);
and U11709 (N_11709,N_11510,N_11542);
or U11710 (N_11710,N_11507,N_11585);
and U11711 (N_11711,N_11583,N_11541);
xnor U11712 (N_11712,N_11589,N_11564);
nor U11713 (N_11713,N_11512,N_11504);
or U11714 (N_11714,N_11515,N_11532);
or U11715 (N_11715,N_11571,N_11517);
nand U11716 (N_11716,N_11533,N_11550);
and U11717 (N_11717,N_11622,N_11566);
and U11718 (N_11718,N_11584,N_11558);
xor U11719 (N_11719,N_11610,N_11548);
xnor U11720 (N_11720,N_11537,N_11623);
nor U11721 (N_11721,N_11531,N_11578);
nand U11722 (N_11722,N_11599,N_11539);
and U11723 (N_11723,N_11544,N_11538);
and U11724 (N_11724,N_11510,N_11540);
and U11725 (N_11725,N_11614,N_11543);
xnor U11726 (N_11726,N_11589,N_11578);
nor U11727 (N_11727,N_11608,N_11590);
or U11728 (N_11728,N_11564,N_11537);
or U11729 (N_11729,N_11503,N_11541);
and U11730 (N_11730,N_11559,N_11503);
and U11731 (N_11731,N_11583,N_11580);
nor U11732 (N_11732,N_11619,N_11592);
nor U11733 (N_11733,N_11573,N_11613);
xor U11734 (N_11734,N_11528,N_11614);
xnor U11735 (N_11735,N_11608,N_11596);
xor U11736 (N_11736,N_11595,N_11537);
xnor U11737 (N_11737,N_11611,N_11594);
nor U11738 (N_11738,N_11573,N_11529);
or U11739 (N_11739,N_11559,N_11506);
xor U11740 (N_11740,N_11608,N_11519);
or U11741 (N_11741,N_11532,N_11565);
xor U11742 (N_11742,N_11613,N_11550);
nand U11743 (N_11743,N_11566,N_11556);
xnor U11744 (N_11744,N_11587,N_11592);
xor U11745 (N_11745,N_11512,N_11535);
xnor U11746 (N_11746,N_11511,N_11520);
nand U11747 (N_11747,N_11528,N_11535);
or U11748 (N_11748,N_11513,N_11616);
xor U11749 (N_11749,N_11530,N_11592);
nand U11750 (N_11750,N_11638,N_11719);
nand U11751 (N_11751,N_11636,N_11666);
nor U11752 (N_11752,N_11692,N_11688);
and U11753 (N_11753,N_11704,N_11731);
and U11754 (N_11754,N_11732,N_11662);
nand U11755 (N_11755,N_11693,N_11641);
nor U11756 (N_11756,N_11680,N_11657);
and U11757 (N_11757,N_11716,N_11709);
nand U11758 (N_11758,N_11739,N_11679);
nor U11759 (N_11759,N_11733,N_11724);
or U11760 (N_11760,N_11713,N_11726);
nand U11761 (N_11761,N_11743,N_11670);
or U11762 (N_11762,N_11632,N_11729);
or U11763 (N_11763,N_11736,N_11695);
or U11764 (N_11764,N_11708,N_11627);
nor U11765 (N_11765,N_11691,N_11698);
and U11766 (N_11766,N_11746,N_11712);
and U11767 (N_11767,N_11673,N_11660);
and U11768 (N_11768,N_11625,N_11669);
xor U11769 (N_11769,N_11705,N_11690);
and U11770 (N_11770,N_11628,N_11676);
nor U11771 (N_11771,N_11634,N_11686);
xor U11772 (N_11772,N_11639,N_11715);
nand U11773 (N_11773,N_11656,N_11701);
and U11774 (N_11774,N_11717,N_11742);
and U11775 (N_11775,N_11720,N_11689);
and U11776 (N_11776,N_11740,N_11672);
xnor U11777 (N_11777,N_11749,N_11647);
or U11778 (N_11778,N_11718,N_11741);
nand U11779 (N_11779,N_11677,N_11682);
or U11780 (N_11780,N_11629,N_11661);
nor U11781 (N_11781,N_11725,N_11697);
nand U11782 (N_11782,N_11687,N_11667);
xor U11783 (N_11783,N_11702,N_11707);
or U11784 (N_11784,N_11745,N_11674);
nand U11785 (N_11785,N_11747,N_11722);
or U11786 (N_11786,N_11654,N_11649);
or U11787 (N_11787,N_11700,N_11748);
nand U11788 (N_11788,N_11664,N_11706);
or U11789 (N_11789,N_11694,N_11714);
xor U11790 (N_11790,N_11630,N_11721);
nand U11791 (N_11791,N_11658,N_11631);
or U11792 (N_11792,N_11650,N_11646);
nand U11793 (N_11793,N_11643,N_11699);
and U11794 (N_11794,N_11684,N_11648);
and U11795 (N_11795,N_11678,N_11728);
nor U11796 (N_11796,N_11642,N_11633);
nand U11797 (N_11797,N_11734,N_11681);
and U11798 (N_11798,N_11644,N_11685);
nand U11799 (N_11799,N_11663,N_11696);
nor U11800 (N_11800,N_11655,N_11730);
xnor U11801 (N_11801,N_11703,N_11737);
or U11802 (N_11802,N_11735,N_11635);
or U11803 (N_11803,N_11645,N_11727);
nor U11804 (N_11804,N_11675,N_11683);
and U11805 (N_11805,N_11671,N_11744);
nor U11806 (N_11806,N_11626,N_11723);
xnor U11807 (N_11807,N_11659,N_11711);
and U11808 (N_11808,N_11640,N_11651);
nand U11809 (N_11809,N_11668,N_11637);
nand U11810 (N_11810,N_11652,N_11653);
or U11811 (N_11811,N_11665,N_11710);
or U11812 (N_11812,N_11738,N_11647);
nand U11813 (N_11813,N_11747,N_11716);
nand U11814 (N_11814,N_11692,N_11697);
and U11815 (N_11815,N_11734,N_11706);
xnor U11816 (N_11816,N_11707,N_11681);
nand U11817 (N_11817,N_11695,N_11687);
nor U11818 (N_11818,N_11689,N_11648);
xnor U11819 (N_11819,N_11685,N_11743);
nor U11820 (N_11820,N_11705,N_11639);
nor U11821 (N_11821,N_11645,N_11705);
nor U11822 (N_11822,N_11691,N_11723);
or U11823 (N_11823,N_11706,N_11632);
and U11824 (N_11824,N_11698,N_11701);
xnor U11825 (N_11825,N_11709,N_11675);
xor U11826 (N_11826,N_11748,N_11636);
nand U11827 (N_11827,N_11654,N_11674);
and U11828 (N_11828,N_11719,N_11668);
or U11829 (N_11829,N_11734,N_11650);
nand U11830 (N_11830,N_11698,N_11629);
and U11831 (N_11831,N_11676,N_11718);
nand U11832 (N_11832,N_11747,N_11663);
and U11833 (N_11833,N_11716,N_11745);
or U11834 (N_11834,N_11632,N_11662);
nand U11835 (N_11835,N_11699,N_11666);
or U11836 (N_11836,N_11689,N_11721);
nand U11837 (N_11837,N_11633,N_11656);
or U11838 (N_11838,N_11630,N_11742);
nand U11839 (N_11839,N_11693,N_11710);
or U11840 (N_11840,N_11717,N_11718);
or U11841 (N_11841,N_11712,N_11671);
nand U11842 (N_11842,N_11721,N_11715);
and U11843 (N_11843,N_11726,N_11715);
xor U11844 (N_11844,N_11695,N_11709);
nand U11845 (N_11845,N_11719,N_11671);
or U11846 (N_11846,N_11749,N_11707);
nand U11847 (N_11847,N_11631,N_11676);
or U11848 (N_11848,N_11658,N_11660);
nand U11849 (N_11849,N_11720,N_11706);
nor U11850 (N_11850,N_11743,N_11715);
and U11851 (N_11851,N_11707,N_11672);
nor U11852 (N_11852,N_11647,N_11635);
nor U11853 (N_11853,N_11662,N_11708);
nand U11854 (N_11854,N_11650,N_11654);
nor U11855 (N_11855,N_11661,N_11660);
nand U11856 (N_11856,N_11711,N_11716);
xor U11857 (N_11857,N_11685,N_11635);
or U11858 (N_11858,N_11669,N_11671);
nor U11859 (N_11859,N_11673,N_11697);
or U11860 (N_11860,N_11748,N_11736);
or U11861 (N_11861,N_11645,N_11634);
xor U11862 (N_11862,N_11686,N_11721);
or U11863 (N_11863,N_11717,N_11692);
nor U11864 (N_11864,N_11743,N_11686);
nand U11865 (N_11865,N_11681,N_11652);
or U11866 (N_11866,N_11742,N_11633);
and U11867 (N_11867,N_11691,N_11663);
or U11868 (N_11868,N_11642,N_11690);
xor U11869 (N_11869,N_11717,N_11721);
nor U11870 (N_11870,N_11676,N_11656);
nand U11871 (N_11871,N_11643,N_11625);
xnor U11872 (N_11872,N_11707,N_11670);
xor U11873 (N_11873,N_11710,N_11688);
xor U11874 (N_11874,N_11672,N_11637);
xnor U11875 (N_11875,N_11818,N_11836);
nand U11876 (N_11876,N_11873,N_11791);
and U11877 (N_11877,N_11823,N_11852);
nand U11878 (N_11878,N_11763,N_11814);
xor U11879 (N_11879,N_11773,N_11808);
and U11880 (N_11880,N_11753,N_11831);
and U11881 (N_11881,N_11806,N_11841);
nand U11882 (N_11882,N_11760,N_11775);
and U11883 (N_11883,N_11768,N_11864);
xnor U11884 (N_11884,N_11787,N_11803);
xor U11885 (N_11885,N_11860,N_11856);
xnor U11886 (N_11886,N_11862,N_11783);
or U11887 (N_11887,N_11772,N_11751);
or U11888 (N_11888,N_11788,N_11833);
xor U11889 (N_11889,N_11770,N_11798);
and U11890 (N_11890,N_11779,N_11758);
xnor U11891 (N_11891,N_11867,N_11871);
nor U11892 (N_11892,N_11825,N_11854);
and U11893 (N_11893,N_11790,N_11802);
nor U11894 (N_11894,N_11769,N_11811);
nor U11895 (N_11895,N_11781,N_11778);
nand U11896 (N_11896,N_11858,N_11816);
nand U11897 (N_11897,N_11771,N_11776);
nand U11898 (N_11898,N_11872,N_11774);
xnor U11899 (N_11899,N_11866,N_11839);
and U11900 (N_11900,N_11801,N_11809);
nor U11901 (N_11901,N_11846,N_11777);
or U11902 (N_11902,N_11804,N_11797);
nand U11903 (N_11903,N_11847,N_11869);
nor U11904 (N_11904,N_11759,N_11799);
xor U11905 (N_11905,N_11765,N_11780);
nor U11906 (N_11906,N_11840,N_11812);
nor U11907 (N_11907,N_11756,N_11817);
nor U11908 (N_11908,N_11834,N_11850);
and U11909 (N_11909,N_11785,N_11784);
or U11910 (N_11910,N_11870,N_11832);
nor U11911 (N_11911,N_11766,N_11849);
or U11912 (N_11912,N_11827,N_11754);
and U11913 (N_11913,N_11755,N_11767);
or U11914 (N_11914,N_11868,N_11835);
nor U11915 (N_11915,N_11810,N_11837);
xor U11916 (N_11916,N_11819,N_11828);
and U11917 (N_11917,N_11786,N_11824);
or U11918 (N_11918,N_11843,N_11821);
xnor U11919 (N_11919,N_11842,N_11851);
xor U11920 (N_11920,N_11807,N_11750);
nor U11921 (N_11921,N_11859,N_11752);
and U11922 (N_11922,N_11826,N_11815);
nor U11923 (N_11923,N_11830,N_11829);
nor U11924 (N_11924,N_11796,N_11793);
and U11925 (N_11925,N_11845,N_11874);
xnor U11926 (N_11926,N_11855,N_11757);
xnor U11927 (N_11927,N_11813,N_11805);
nand U11928 (N_11928,N_11800,N_11792);
or U11929 (N_11929,N_11838,N_11782);
nor U11930 (N_11930,N_11861,N_11863);
and U11931 (N_11931,N_11865,N_11822);
or U11932 (N_11932,N_11853,N_11764);
or U11933 (N_11933,N_11844,N_11848);
and U11934 (N_11934,N_11820,N_11762);
xnor U11935 (N_11935,N_11794,N_11795);
or U11936 (N_11936,N_11789,N_11857);
xor U11937 (N_11937,N_11761,N_11777);
xnor U11938 (N_11938,N_11872,N_11844);
and U11939 (N_11939,N_11810,N_11786);
or U11940 (N_11940,N_11825,N_11764);
xor U11941 (N_11941,N_11842,N_11831);
or U11942 (N_11942,N_11753,N_11815);
xnor U11943 (N_11943,N_11783,N_11850);
xnor U11944 (N_11944,N_11798,N_11755);
and U11945 (N_11945,N_11758,N_11818);
and U11946 (N_11946,N_11843,N_11848);
nor U11947 (N_11947,N_11790,N_11804);
nor U11948 (N_11948,N_11822,N_11853);
nor U11949 (N_11949,N_11793,N_11860);
nor U11950 (N_11950,N_11811,N_11807);
xor U11951 (N_11951,N_11842,N_11857);
and U11952 (N_11952,N_11794,N_11867);
nor U11953 (N_11953,N_11784,N_11799);
nand U11954 (N_11954,N_11799,N_11850);
nand U11955 (N_11955,N_11804,N_11821);
or U11956 (N_11956,N_11753,N_11770);
or U11957 (N_11957,N_11784,N_11856);
nor U11958 (N_11958,N_11833,N_11812);
xor U11959 (N_11959,N_11874,N_11862);
or U11960 (N_11960,N_11786,N_11774);
xor U11961 (N_11961,N_11868,N_11857);
and U11962 (N_11962,N_11751,N_11797);
or U11963 (N_11963,N_11835,N_11847);
nor U11964 (N_11964,N_11753,N_11821);
and U11965 (N_11965,N_11857,N_11803);
nor U11966 (N_11966,N_11817,N_11758);
or U11967 (N_11967,N_11857,N_11833);
nor U11968 (N_11968,N_11828,N_11838);
and U11969 (N_11969,N_11861,N_11751);
nand U11970 (N_11970,N_11807,N_11824);
nor U11971 (N_11971,N_11829,N_11817);
and U11972 (N_11972,N_11844,N_11805);
xor U11973 (N_11973,N_11775,N_11870);
nor U11974 (N_11974,N_11854,N_11755);
xnor U11975 (N_11975,N_11816,N_11760);
nand U11976 (N_11976,N_11753,N_11789);
nand U11977 (N_11977,N_11842,N_11778);
xor U11978 (N_11978,N_11791,N_11872);
nand U11979 (N_11979,N_11773,N_11842);
nor U11980 (N_11980,N_11796,N_11862);
nor U11981 (N_11981,N_11835,N_11770);
or U11982 (N_11982,N_11839,N_11796);
nor U11983 (N_11983,N_11790,N_11800);
and U11984 (N_11984,N_11856,N_11761);
and U11985 (N_11985,N_11790,N_11784);
xnor U11986 (N_11986,N_11765,N_11851);
or U11987 (N_11987,N_11853,N_11815);
nor U11988 (N_11988,N_11803,N_11853);
nor U11989 (N_11989,N_11764,N_11847);
and U11990 (N_11990,N_11772,N_11841);
nand U11991 (N_11991,N_11782,N_11833);
and U11992 (N_11992,N_11811,N_11788);
nor U11993 (N_11993,N_11866,N_11828);
xnor U11994 (N_11994,N_11847,N_11765);
and U11995 (N_11995,N_11820,N_11759);
and U11996 (N_11996,N_11843,N_11804);
or U11997 (N_11997,N_11851,N_11837);
xnor U11998 (N_11998,N_11859,N_11798);
nand U11999 (N_11999,N_11833,N_11842);
and U12000 (N_12000,N_11897,N_11930);
nand U12001 (N_12001,N_11880,N_11964);
xor U12002 (N_12002,N_11912,N_11972);
nand U12003 (N_12003,N_11876,N_11933);
nor U12004 (N_12004,N_11960,N_11909);
nand U12005 (N_12005,N_11996,N_11913);
and U12006 (N_12006,N_11941,N_11886);
xnor U12007 (N_12007,N_11956,N_11998);
nand U12008 (N_12008,N_11899,N_11881);
nand U12009 (N_12009,N_11918,N_11890);
nor U12010 (N_12010,N_11985,N_11993);
xnor U12011 (N_12011,N_11932,N_11939);
and U12012 (N_12012,N_11907,N_11896);
xnor U12013 (N_12013,N_11953,N_11948);
or U12014 (N_12014,N_11962,N_11955);
xnor U12015 (N_12015,N_11914,N_11936);
and U12016 (N_12016,N_11879,N_11944);
and U12017 (N_12017,N_11893,N_11999);
nor U12018 (N_12018,N_11892,N_11987);
nor U12019 (N_12019,N_11977,N_11984);
and U12020 (N_12020,N_11888,N_11940);
or U12021 (N_12021,N_11973,N_11928);
or U12022 (N_12022,N_11905,N_11951);
nor U12023 (N_12023,N_11954,N_11875);
nand U12024 (N_12024,N_11937,N_11885);
nor U12025 (N_12025,N_11898,N_11986);
and U12026 (N_12026,N_11910,N_11916);
nand U12027 (N_12027,N_11903,N_11882);
nand U12028 (N_12028,N_11908,N_11974);
nor U12029 (N_12029,N_11924,N_11929);
or U12030 (N_12030,N_11963,N_11971);
or U12031 (N_12031,N_11980,N_11877);
nand U12032 (N_12032,N_11883,N_11878);
and U12033 (N_12033,N_11966,N_11995);
and U12034 (N_12034,N_11949,N_11887);
or U12035 (N_12035,N_11981,N_11957);
nor U12036 (N_12036,N_11884,N_11978);
or U12037 (N_12037,N_11889,N_11931);
or U12038 (N_12038,N_11979,N_11935);
xnor U12039 (N_12039,N_11994,N_11959);
and U12040 (N_12040,N_11946,N_11983);
nor U12041 (N_12041,N_11967,N_11900);
nor U12042 (N_12042,N_11922,N_11919);
nor U12043 (N_12043,N_11961,N_11923);
and U12044 (N_12044,N_11945,N_11917);
or U12045 (N_12045,N_11988,N_11952);
nand U12046 (N_12046,N_11906,N_11989);
nor U12047 (N_12047,N_11991,N_11942);
nand U12048 (N_12048,N_11925,N_11982);
and U12049 (N_12049,N_11976,N_11926);
xnor U12050 (N_12050,N_11990,N_11965);
nand U12051 (N_12051,N_11938,N_11950);
or U12052 (N_12052,N_11958,N_11943);
and U12053 (N_12053,N_11992,N_11901);
nand U12054 (N_12054,N_11934,N_11891);
xor U12055 (N_12055,N_11915,N_11969);
xor U12056 (N_12056,N_11902,N_11895);
and U12057 (N_12057,N_11920,N_11927);
or U12058 (N_12058,N_11947,N_11968);
or U12059 (N_12059,N_11997,N_11970);
nand U12060 (N_12060,N_11975,N_11921);
and U12061 (N_12061,N_11911,N_11894);
nor U12062 (N_12062,N_11904,N_11909);
nor U12063 (N_12063,N_11994,N_11910);
and U12064 (N_12064,N_11998,N_11885);
nand U12065 (N_12065,N_11974,N_11960);
and U12066 (N_12066,N_11981,N_11922);
nor U12067 (N_12067,N_11956,N_11967);
xor U12068 (N_12068,N_11936,N_11983);
nand U12069 (N_12069,N_11999,N_11956);
and U12070 (N_12070,N_11946,N_11955);
or U12071 (N_12071,N_11894,N_11875);
nor U12072 (N_12072,N_11944,N_11973);
xor U12073 (N_12073,N_11913,N_11985);
nor U12074 (N_12074,N_11887,N_11911);
nand U12075 (N_12075,N_11976,N_11994);
nor U12076 (N_12076,N_11998,N_11941);
and U12077 (N_12077,N_11960,N_11913);
and U12078 (N_12078,N_11939,N_11962);
and U12079 (N_12079,N_11876,N_11949);
or U12080 (N_12080,N_11983,N_11999);
xor U12081 (N_12081,N_11893,N_11911);
xor U12082 (N_12082,N_11966,N_11924);
nor U12083 (N_12083,N_11949,N_11890);
xnor U12084 (N_12084,N_11965,N_11880);
xnor U12085 (N_12085,N_11939,N_11902);
nor U12086 (N_12086,N_11932,N_11936);
nor U12087 (N_12087,N_11962,N_11938);
nand U12088 (N_12088,N_11883,N_11999);
and U12089 (N_12089,N_11940,N_11911);
xnor U12090 (N_12090,N_11913,N_11878);
nor U12091 (N_12091,N_11979,N_11926);
and U12092 (N_12092,N_11942,N_11878);
and U12093 (N_12093,N_11946,N_11989);
xnor U12094 (N_12094,N_11992,N_11882);
nand U12095 (N_12095,N_11938,N_11960);
and U12096 (N_12096,N_11926,N_11970);
nor U12097 (N_12097,N_11890,N_11925);
nand U12098 (N_12098,N_11992,N_11951);
nor U12099 (N_12099,N_11966,N_11889);
nor U12100 (N_12100,N_11964,N_11910);
nor U12101 (N_12101,N_11948,N_11924);
xnor U12102 (N_12102,N_11944,N_11910);
xor U12103 (N_12103,N_11907,N_11973);
xnor U12104 (N_12104,N_11889,N_11920);
nor U12105 (N_12105,N_11948,N_11985);
nand U12106 (N_12106,N_11925,N_11971);
xnor U12107 (N_12107,N_11906,N_11956);
and U12108 (N_12108,N_11993,N_11920);
or U12109 (N_12109,N_11999,N_11954);
and U12110 (N_12110,N_11942,N_11902);
and U12111 (N_12111,N_11899,N_11919);
nand U12112 (N_12112,N_11908,N_11922);
nand U12113 (N_12113,N_11875,N_11898);
xnor U12114 (N_12114,N_11887,N_11937);
or U12115 (N_12115,N_11916,N_11997);
nor U12116 (N_12116,N_11894,N_11883);
xnor U12117 (N_12117,N_11961,N_11997);
nor U12118 (N_12118,N_11998,N_11929);
or U12119 (N_12119,N_11924,N_11906);
or U12120 (N_12120,N_11893,N_11935);
and U12121 (N_12121,N_11914,N_11993);
or U12122 (N_12122,N_11990,N_11887);
nand U12123 (N_12123,N_11937,N_11898);
or U12124 (N_12124,N_11988,N_11885);
nand U12125 (N_12125,N_12016,N_12042);
or U12126 (N_12126,N_12011,N_12046);
and U12127 (N_12127,N_12080,N_12112);
nor U12128 (N_12128,N_12121,N_12054);
nand U12129 (N_12129,N_12087,N_12118);
and U12130 (N_12130,N_12015,N_12033);
or U12131 (N_12131,N_12041,N_12063);
nor U12132 (N_12132,N_12071,N_12006);
nor U12133 (N_12133,N_12057,N_12044);
xnor U12134 (N_12134,N_12020,N_12089);
nand U12135 (N_12135,N_12052,N_12120);
nor U12136 (N_12136,N_12085,N_12068);
or U12137 (N_12137,N_12022,N_12083);
xnor U12138 (N_12138,N_12109,N_12058);
xor U12139 (N_12139,N_12017,N_12123);
xnor U12140 (N_12140,N_12019,N_12053);
xor U12141 (N_12141,N_12060,N_12021);
xnor U12142 (N_12142,N_12105,N_12094);
or U12143 (N_12143,N_12029,N_12078);
or U12144 (N_12144,N_12073,N_12075);
and U12145 (N_12145,N_12050,N_12014);
nand U12146 (N_12146,N_12047,N_12103);
nand U12147 (N_12147,N_12090,N_12099);
xor U12148 (N_12148,N_12107,N_12001);
or U12149 (N_12149,N_12061,N_12114);
nor U12150 (N_12150,N_12030,N_12082);
and U12151 (N_12151,N_12034,N_12024);
nand U12152 (N_12152,N_12023,N_12088);
xor U12153 (N_12153,N_12067,N_12056);
nor U12154 (N_12154,N_12074,N_12101);
nor U12155 (N_12155,N_12081,N_12095);
nand U12156 (N_12156,N_12038,N_12048);
and U12157 (N_12157,N_12027,N_12059);
nand U12158 (N_12158,N_12069,N_12003);
nor U12159 (N_12159,N_12000,N_12025);
or U12160 (N_12160,N_12004,N_12039);
xor U12161 (N_12161,N_12010,N_12117);
or U12162 (N_12162,N_12093,N_12012);
and U12163 (N_12163,N_12049,N_12035);
and U12164 (N_12164,N_12124,N_12102);
and U12165 (N_12165,N_12066,N_12045);
nand U12166 (N_12166,N_12122,N_12108);
xnor U12167 (N_12167,N_12013,N_12115);
nor U12168 (N_12168,N_12065,N_12104);
or U12169 (N_12169,N_12100,N_12043);
nor U12170 (N_12170,N_12111,N_12005);
and U12171 (N_12171,N_12076,N_12062);
nand U12172 (N_12172,N_12032,N_12113);
nor U12173 (N_12173,N_12079,N_12070);
xor U12174 (N_12174,N_12072,N_12036);
nand U12175 (N_12175,N_12002,N_12096);
or U12176 (N_12176,N_12055,N_12092);
nor U12177 (N_12177,N_12110,N_12119);
nor U12178 (N_12178,N_12018,N_12051);
xor U12179 (N_12179,N_12026,N_12116);
nand U12180 (N_12180,N_12031,N_12098);
nand U12181 (N_12181,N_12007,N_12077);
or U12182 (N_12182,N_12084,N_12106);
xor U12183 (N_12183,N_12064,N_12086);
and U12184 (N_12184,N_12097,N_12091);
nor U12185 (N_12185,N_12037,N_12009);
nand U12186 (N_12186,N_12008,N_12040);
xnor U12187 (N_12187,N_12028,N_12095);
and U12188 (N_12188,N_12090,N_12113);
or U12189 (N_12189,N_12025,N_12107);
and U12190 (N_12190,N_12011,N_12064);
nor U12191 (N_12191,N_12119,N_12048);
and U12192 (N_12192,N_12103,N_12082);
or U12193 (N_12193,N_12084,N_12015);
or U12194 (N_12194,N_12002,N_12010);
xor U12195 (N_12195,N_12053,N_12001);
nand U12196 (N_12196,N_12014,N_12069);
and U12197 (N_12197,N_12020,N_12114);
nor U12198 (N_12198,N_12065,N_12050);
nor U12199 (N_12199,N_12036,N_12026);
or U12200 (N_12200,N_12078,N_12039);
and U12201 (N_12201,N_12002,N_12039);
or U12202 (N_12202,N_12011,N_12109);
xor U12203 (N_12203,N_12102,N_12068);
and U12204 (N_12204,N_12072,N_12005);
nand U12205 (N_12205,N_12063,N_12011);
nor U12206 (N_12206,N_12008,N_12080);
nand U12207 (N_12207,N_12091,N_12062);
or U12208 (N_12208,N_12087,N_12060);
nor U12209 (N_12209,N_12067,N_12003);
or U12210 (N_12210,N_12102,N_12044);
xor U12211 (N_12211,N_12050,N_12082);
xnor U12212 (N_12212,N_12003,N_12016);
nor U12213 (N_12213,N_12025,N_12060);
xor U12214 (N_12214,N_12104,N_12019);
or U12215 (N_12215,N_12074,N_12005);
nor U12216 (N_12216,N_12049,N_12010);
nor U12217 (N_12217,N_12014,N_12092);
nand U12218 (N_12218,N_12077,N_12013);
xor U12219 (N_12219,N_12016,N_12111);
and U12220 (N_12220,N_12119,N_12096);
xor U12221 (N_12221,N_12090,N_12060);
and U12222 (N_12222,N_12093,N_12036);
and U12223 (N_12223,N_12064,N_12016);
nand U12224 (N_12224,N_12086,N_12060);
or U12225 (N_12225,N_12003,N_12101);
nand U12226 (N_12226,N_12100,N_12047);
nor U12227 (N_12227,N_12001,N_12009);
and U12228 (N_12228,N_12029,N_12034);
xor U12229 (N_12229,N_12070,N_12043);
nor U12230 (N_12230,N_12103,N_12066);
xor U12231 (N_12231,N_12058,N_12112);
nor U12232 (N_12232,N_12099,N_12027);
and U12233 (N_12233,N_12060,N_12077);
nand U12234 (N_12234,N_12039,N_12022);
xor U12235 (N_12235,N_12008,N_12086);
nor U12236 (N_12236,N_12093,N_12044);
and U12237 (N_12237,N_12071,N_12048);
or U12238 (N_12238,N_12020,N_12102);
and U12239 (N_12239,N_12061,N_12010);
or U12240 (N_12240,N_12086,N_12110);
nand U12241 (N_12241,N_12041,N_12044);
and U12242 (N_12242,N_12022,N_12110);
xnor U12243 (N_12243,N_12027,N_12046);
or U12244 (N_12244,N_12114,N_12022);
and U12245 (N_12245,N_12078,N_12072);
nor U12246 (N_12246,N_12004,N_12029);
nand U12247 (N_12247,N_12056,N_12090);
xor U12248 (N_12248,N_12045,N_12092);
nand U12249 (N_12249,N_12037,N_12008);
nor U12250 (N_12250,N_12129,N_12198);
xnor U12251 (N_12251,N_12164,N_12156);
xor U12252 (N_12252,N_12233,N_12180);
nand U12253 (N_12253,N_12151,N_12135);
or U12254 (N_12254,N_12216,N_12138);
xor U12255 (N_12255,N_12172,N_12195);
nand U12256 (N_12256,N_12249,N_12136);
nand U12257 (N_12257,N_12197,N_12147);
nand U12258 (N_12258,N_12179,N_12132);
and U12259 (N_12259,N_12226,N_12165);
and U12260 (N_12260,N_12144,N_12240);
and U12261 (N_12261,N_12182,N_12178);
nor U12262 (N_12262,N_12148,N_12228);
nor U12263 (N_12263,N_12183,N_12139);
nor U12264 (N_12264,N_12208,N_12238);
nor U12265 (N_12265,N_12199,N_12169);
nand U12266 (N_12266,N_12171,N_12205);
nor U12267 (N_12267,N_12157,N_12215);
nand U12268 (N_12268,N_12154,N_12152);
or U12269 (N_12269,N_12186,N_12159);
nor U12270 (N_12270,N_12125,N_12213);
and U12271 (N_12271,N_12146,N_12174);
nor U12272 (N_12272,N_12194,N_12243);
nor U12273 (N_12273,N_12241,N_12234);
or U12274 (N_12274,N_12224,N_12206);
nor U12275 (N_12275,N_12184,N_12229);
and U12276 (N_12276,N_12202,N_12221);
or U12277 (N_12277,N_12133,N_12158);
nor U12278 (N_12278,N_12155,N_12160);
nand U12279 (N_12279,N_12141,N_12212);
nand U12280 (N_12280,N_12219,N_12126);
and U12281 (N_12281,N_12227,N_12204);
xnor U12282 (N_12282,N_12127,N_12170);
nand U12283 (N_12283,N_12223,N_12232);
nand U12284 (N_12284,N_12220,N_12150);
nor U12285 (N_12285,N_12218,N_12231);
nor U12286 (N_12286,N_12207,N_12214);
or U12287 (N_12287,N_12193,N_12190);
and U12288 (N_12288,N_12203,N_12167);
xnor U12289 (N_12289,N_12187,N_12225);
nand U12290 (N_12290,N_12185,N_12153);
and U12291 (N_12291,N_12149,N_12191);
nor U12292 (N_12292,N_12210,N_12188);
nand U12293 (N_12293,N_12217,N_12245);
and U12294 (N_12294,N_12173,N_12128);
xnor U12295 (N_12295,N_12239,N_12181);
nor U12296 (N_12296,N_12230,N_12196);
nand U12297 (N_12297,N_12211,N_12237);
and U12298 (N_12298,N_12246,N_12222);
or U12299 (N_12299,N_12235,N_12131);
or U12300 (N_12300,N_12242,N_12248);
and U12301 (N_12301,N_12201,N_12200);
nand U12302 (N_12302,N_12236,N_12140);
xor U12303 (N_12303,N_12175,N_12168);
nand U12304 (N_12304,N_12143,N_12134);
and U12305 (N_12305,N_12166,N_12142);
nand U12306 (N_12306,N_12145,N_12161);
nor U12307 (N_12307,N_12244,N_12162);
nor U12308 (N_12308,N_12209,N_12137);
or U12309 (N_12309,N_12177,N_12192);
nor U12310 (N_12310,N_12247,N_12163);
nand U12311 (N_12311,N_12176,N_12189);
nor U12312 (N_12312,N_12130,N_12245);
nand U12313 (N_12313,N_12243,N_12249);
nand U12314 (N_12314,N_12200,N_12129);
and U12315 (N_12315,N_12184,N_12216);
and U12316 (N_12316,N_12171,N_12154);
xnor U12317 (N_12317,N_12166,N_12220);
or U12318 (N_12318,N_12230,N_12176);
nor U12319 (N_12319,N_12127,N_12148);
nor U12320 (N_12320,N_12232,N_12241);
and U12321 (N_12321,N_12157,N_12163);
xor U12322 (N_12322,N_12141,N_12161);
nand U12323 (N_12323,N_12178,N_12227);
and U12324 (N_12324,N_12161,N_12183);
nand U12325 (N_12325,N_12185,N_12234);
and U12326 (N_12326,N_12151,N_12137);
or U12327 (N_12327,N_12171,N_12209);
or U12328 (N_12328,N_12175,N_12229);
and U12329 (N_12329,N_12157,N_12130);
or U12330 (N_12330,N_12232,N_12136);
and U12331 (N_12331,N_12208,N_12166);
nor U12332 (N_12332,N_12139,N_12163);
nor U12333 (N_12333,N_12137,N_12217);
nand U12334 (N_12334,N_12161,N_12158);
nor U12335 (N_12335,N_12140,N_12128);
nor U12336 (N_12336,N_12233,N_12230);
or U12337 (N_12337,N_12192,N_12140);
and U12338 (N_12338,N_12149,N_12151);
and U12339 (N_12339,N_12226,N_12146);
nand U12340 (N_12340,N_12175,N_12194);
and U12341 (N_12341,N_12140,N_12145);
or U12342 (N_12342,N_12196,N_12167);
or U12343 (N_12343,N_12152,N_12146);
nand U12344 (N_12344,N_12180,N_12157);
nor U12345 (N_12345,N_12184,N_12141);
nand U12346 (N_12346,N_12190,N_12158);
nand U12347 (N_12347,N_12133,N_12219);
or U12348 (N_12348,N_12193,N_12189);
nor U12349 (N_12349,N_12135,N_12175);
xor U12350 (N_12350,N_12185,N_12201);
xnor U12351 (N_12351,N_12158,N_12152);
nand U12352 (N_12352,N_12130,N_12152);
and U12353 (N_12353,N_12204,N_12195);
and U12354 (N_12354,N_12200,N_12231);
nand U12355 (N_12355,N_12212,N_12166);
and U12356 (N_12356,N_12176,N_12190);
and U12357 (N_12357,N_12224,N_12227);
and U12358 (N_12358,N_12212,N_12227);
nand U12359 (N_12359,N_12233,N_12173);
or U12360 (N_12360,N_12249,N_12192);
nand U12361 (N_12361,N_12221,N_12171);
xnor U12362 (N_12362,N_12141,N_12196);
nor U12363 (N_12363,N_12126,N_12183);
xor U12364 (N_12364,N_12173,N_12133);
nor U12365 (N_12365,N_12197,N_12136);
xnor U12366 (N_12366,N_12199,N_12239);
xnor U12367 (N_12367,N_12225,N_12126);
and U12368 (N_12368,N_12131,N_12188);
or U12369 (N_12369,N_12139,N_12153);
and U12370 (N_12370,N_12219,N_12147);
and U12371 (N_12371,N_12148,N_12144);
or U12372 (N_12372,N_12186,N_12160);
nor U12373 (N_12373,N_12145,N_12139);
and U12374 (N_12374,N_12231,N_12179);
xor U12375 (N_12375,N_12278,N_12373);
or U12376 (N_12376,N_12309,N_12302);
nor U12377 (N_12377,N_12319,N_12300);
nand U12378 (N_12378,N_12253,N_12329);
or U12379 (N_12379,N_12252,N_12335);
and U12380 (N_12380,N_12352,N_12327);
xnor U12381 (N_12381,N_12356,N_12343);
and U12382 (N_12382,N_12261,N_12273);
nand U12383 (N_12383,N_12360,N_12315);
or U12384 (N_12384,N_12367,N_12330);
xnor U12385 (N_12385,N_12279,N_12320);
nor U12386 (N_12386,N_12358,N_12306);
xnor U12387 (N_12387,N_12298,N_12256);
and U12388 (N_12388,N_12342,N_12281);
nor U12389 (N_12389,N_12304,N_12296);
nor U12390 (N_12390,N_12332,N_12303);
xnor U12391 (N_12391,N_12372,N_12322);
nand U12392 (N_12392,N_12338,N_12266);
and U12393 (N_12393,N_12346,N_12365);
and U12394 (N_12394,N_12254,N_12314);
and U12395 (N_12395,N_12313,N_12262);
or U12396 (N_12396,N_12287,N_12270);
or U12397 (N_12397,N_12350,N_12265);
nor U12398 (N_12398,N_12277,N_12308);
and U12399 (N_12399,N_12361,N_12347);
xnor U12400 (N_12400,N_12299,N_12301);
and U12401 (N_12401,N_12328,N_12364);
and U12402 (N_12402,N_12251,N_12286);
and U12403 (N_12403,N_12258,N_12267);
and U12404 (N_12404,N_12316,N_12374);
and U12405 (N_12405,N_12250,N_12255);
nand U12406 (N_12406,N_12268,N_12354);
and U12407 (N_12407,N_12333,N_12331);
or U12408 (N_12408,N_12311,N_12282);
or U12409 (N_12409,N_12368,N_12289);
nand U12410 (N_12410,N_12344,N_12284);
or U12411 (N_12411,N_12359,N_12326);
xor U12412 (N_12412,N_12293,N_12325);
xnor U12413 (N_12413,N_12260,N_12341);
and U12414 (N_12414,N_12280,N_12272);
or U12415 (N_12415,N_12305,N_12259);
and U12416 (N_12416,N_12351,N_12292);
nor U12417 (N_12417,N_12257,N_12357);
nand U12418 (N_12418,N_12339,N_12263);
nand U12419 (N_12419,N_12353,N_12283);
nand U12420 (N_12420,N_12294,N_12317);
xor U12421 (N_12421,N_12291,N_12271);
or U12422 (N_12422,N_12337,N_12371);
or U12423 (N_12423,N_12290,N_12323);
nand U12424 (N_12424,N_12307,N_12340);
xnor U12425 (N_12425,N_12297,N_12348);
xnor U12426 (N_12426,N_12324,N_12321);
nor U12427 (N_12427,N_12295,N_12349);
nand U12428 (N_12428,N_12312,N_12362);
nor U12429 (N_12429,N_12366,N_12355);
nor U12430 (N_12430,N_12264,N_12274);
and U12431 (N_12431,N_12370,N_12310);
or U12432 (N_12432,N_12345,N_12276);
xor U12433 (N_12433,N_12336,N_12285);
nor U12434 (N_12434,N_12318,N_12288);
nor U12435 (N_12435,N_12369,N_12275);
or U12436 (N_12436,N_12363,N_12269);
xnor U12437 (N_12437,N_12334,N_12330);
nand U12438 (N_12438,N_12351,N_12250);
and U12439 (N_12439,N_12301,N_12369);
and U12440 (N_12440,N_12315,N_12272);
nand U12441 (N_12441,N_12254,N_12287);
or U12442 (N_12442,N_12293,N_12354);
xor U12443 (N_12443,N_12312,N_12274);
nor U12444 (N_12444,N_12339,N_12301);
or U12445 (N_12445,N_12274,N_12296);
or U12446 (N_12446,N_12266,N_12311);
or U12447 (N_12447,N_12294,N_12285);
nand U12448 (N_12448,N_12303,N_12319);
nand U12449 (N_12449,N_12327,N_12332);
and U12450 (N_12450,N_12307,N_12299);
nand U12451 (N_12451,N_12335,N_12352);
or U12452 (N_12452,N_12301,N_12281);
and U12453 (N_12453,N_12269,N_12291);
or U12454 (N_12454,N_12318,N_12253);
and U12455 (N_12455,N_12251,N_12282);
nor U12456 (N_12456,N_12341,N_12306);
xor U12457 (N_12457,N_12332,N_12253);
or U12458 (N_12458,N_12351,N_12298);
or U12459 (N_12459,N_12341,N_12258);
and U12460 (N_12460,N_12326,N_12318);
nand U12461 (N_12461,N_12374,N_12289);
xnor U12462 (N_12462,N_12253,N_12285);
nand U12463 (N_12463,N_12298,N_12287);
and U12464 (N_12464,N_12261,N_12300);
nand U12465 (N_12465,N_12369,N_12300);
nand U12466 (N_12466,N_12349,N_12294);
xnor U12467 (N_12467,N_12343,N_12335);
and U12468 (N_12468,N_12328,N_12283);
nand U12469 (N_12469,N_12347,N_12362);
or U12470 (N_12470,N_12330,N_12263);
nor U12471 (N_12471,N_12309,N_12301);
nand U12472 (N_12472,N_12272,N_12332);
and U12473 (N_12473,N_12290,N_12281);
nor U12474 (N_12474,N_12263,N_12285);
and U12475 (N_12475,N_12279,N_12259);
nand U12476 (N_12476,N_12326,N_12271);
nand U12477 (N_12477,N_12258,N_12353);
or U12478 (N_12478,N_12335,N_12348);
xor U12479 (N_12479,N_12351,N_12328);
and U12480 (N_12480,N_12354,N_12338);
or U12481 (N_12481,N_12251,N_12365);
nand U12482 (N_12482,N_12323,N_12287);
nand U12483 (N_12483,N_12288,N_12322);
or U12484 (N_12484,N_12338,N_12267);
or U12485 (N_12485,N_12366,N_12258);
xnor U12486 (N_12486,N_12368,N_12326);
nor U12487 (N_12487,N_12259,N_12299);
or U12488 (N_12488,N_12278,N_12263);
or U12489 (N_12489,N_12346,N_12288);
or U12490 (N_12490,N_12253,N_12362);
nor U12491 (N_12491,N_12372,N_12315);
nor U12492 (N_12492,N_12343,N_12332);
nand U12493 (N_12493,N_12268,N_12277);
and U12494 (N_12494,N_12259,N_12373);
xor U12495 (N_12495,N_12325,N_12373);
and U12496 (N_12496,N_12325,N_12354);
nand U12497 (N_12497,N_12334,N_12307);
nand U12498 (N_12498,N_12343,N_12350);
nor U12499 (N_12499,N_12307,N_12372);
nor U12500 (N_12500,N_12489,N_12410);
or U12501 (N_12501,N_12461,N_12480);
or U12502 (N_12502,N_12465,N_12469);
or U12503 (N_12503,N_12488,N_12479);
and U12504 (N_12504,N_12445,N_12422);
and U12505 (N_12505,N_12402,N_12484);
nand U12506 (N_12506,N_12476,N_12440);
nand U12507 (N_12507,N_12456,N_12482);
nand U12508 (N_12508,N_12483,N_12494);
nor U12509 (N_12509,N_12408,N_12398);
nor U12510 (N_12510,N_12405,N_12437);
xor U12511 (N_12511,N_12397,N_12430);
xnor U12512 (N_12512,N_12384,N_12428);
nand U12513 (N_12513,N_12477,N_12485);
xnor U12514 (N_12514,N_12418,N_12468);
and U12515 (N_12515,N_12406,N_12481);
or U12516 (N_12516,N_12470,N_12420);
nor U12517 (N_12517,N_12453,N_12424);
or U12518 (N_12518,N_12492,N_12446);
nand U12519 (N_12519,N_12383,N_12382);
nor U12520 (N_12520,N_12423,N_12433);
xnor U12521 (N_12521,N_12381,N_12444);
or U12522 (N_12522,N_12415,N_12394);
and U12523 (N_12523,N_12390,N_12464);
nor U12524 (N_12524,N_12458,N_12407);
nand U12525 (N_12525,N_12435,N_12409);
or U12526 (N_12526,N_12391,N_12447);
or U12527 (N_12527,N_12425,N_12442);
or U12528 (N_12528,N_12459,N_12376);
nand U12529 (N_12529,N_12416,N_12493);
or U12530 (N_12530,N_12414,N_12475);
nand U12531 (N_12531,N_12491,N_12497);
nor U12532 (N_12532,N_12432,N_12378);
and U12533 (N_12533,N_12380,N_12448);
nand U12534 (N_12534,N_12439,N_12411);
and U12535 (N_12535,N_12457,N_12388);
or U12536 (N_12536,N_12441,N_12421);
or U12537 (N_12537,N_12431,N_12496);
or U12538 (N_12538,N_12389,N_12434);
and U12539 (N_12539,N_12379,N_12499);
xnor U12540 (N_12540,N_12443,N_12377);
and U12541 (N_12541,N_12399,N_12385);
nand U12542 (N_12542,N_12392,N_12473);
nand U12543 (N_12543,N_12474,N_12472);
or U12544 (N_12544,N_12467,N_12436);
xor U12545 (N_12545,N_12463,N_12478);
or U12546 (N_12546,N_12490,N_12452);
and U12547 (N_12547,N_12417,N_12396);
nor U12548 (N_12548,N_12419,N_12454);
nand U12549 (N_12549,N_12451,N_12449);
and U12550 (N_12550,N_12400,N_12487);
or U12551 (N_12551,N_12462,N_12387);
xor U12552 (N_12552,N_12426,N_12429);
nor U12553 (N_12553,N_12486,N_12427);
xor U12554 (N_12554,N_12395,N_12495);
nand U12555 (N_12555,N_12404,N_12403);
nor U12556 (N_12556,N_12438,N_12401);
nand U12557 (N_12557,N_12413,N_12375);
nor U12558 (N_12558,N_12466,N_12412);
xnor U12559 (N_12559,N_12460,N_12450);
xor U12560 (N_12560,N_12393,N_12471);
xnor U12561 (N_12561,N_12386,N_12498);
nor U12562 (N_12562,N_12455,N_12475);
nand U12563 (N_12563,N_12495,N_12412);
and U12564 (N_12564,N_12486,N_12464);
and U12565 (N_12565,N_12386,N_12435);
nor U12566 (N_12566,N_12454,N_12387);
or U12567 (N_12567,N_12415,N_12401);
nor U12568 (N_12568,N_12429,N_12427);
xnor U12569 (N_12569,N_12485,N_12415);
nor U12570 (N_12570,N_12452,N_12485);
xnor U12571 (N_12571,N_12434,N_12410);
xor U12572 (N_12572,N_12446,N_12426);
or U12573 (N_12573,N_12493,N_12483);
nand U12574 (N_12574,N_12434,N_12494);
nand U12575 (N_12575,N_12389,N_12423);
and U12576 (N_12576,N_12466,N_12454);
nand U12577 (N_12577,N_12449,N_12476);
xnor U12578 (N_12578,N_12440,N_12444);
and U12579 (N_12579,N_12422,N_12415);
xnor U12580 (N_12580,N_12430,N_12407);
or U12581 (N_12581,N_12392,N_12468);
nand U12582 (N_12582,N_12487,N_12423);
xnor U12583 (N_12583,N_12380,N_12402);
or U12584 (N_12584,N_12446,N_12449);
nand U12585 (N_12585,N_12493,N_12413);
xor U12586 (N_12586,N_12381,N_12431);
or U12587 (N_12587,N_12475,N_12398);
and U12588 (N_12588,N_12435,N_12399);
and U12589 (N_12589,N_12388,N_12497);
nand U12590 (N_12590,N_12469,N_12460);
or U12591 (N_12591,N_12414,N_12379);
nor U12592 (N_12592,N_12430,N_12436);
nor U12593 (N_12593,N_12430,N_12387);
and U12594 (N_12594,N_12420,N_12392);
or U12595 (N_12595,N_12467,N_12409);
or U12596 (N_12596,N_12406,N_12403);
xnor U12597 (N_12597,N_12466,N_12497);
nor U12598 (N_12598,N_12486,N_12416);
and U12599 (N_12599,N_12450,N_12475);
nand U12600 (N_12600,N_12454,N_12377);
xnor U12601 (N_12601,N_12402,N_12436);
xnor U12602 (N_12602,N_12408,N_12466);
nor U12603 (N_12603,N_12488,N_12450);
xor U12604 (N_12604,N_12455,N_12391);
xor U12605 (N_12605,N_12467,N_12422);
or U12606 (N_12606,N_12470,N_12387);
or U12607 (N_12607,N_12401,N_12411);
nand U12608 (N_12608,N_12412,N_12434);
nand U12609 (N_12609,N_12388,N_12444);
or U12610 (N_12610,N_12478,N_12409);
nor U12611 (N_12611,N_12470,N_12479);
or U12612 (N_12612,N_12426,N_12403);
or U12613 (N_12613,N_12380,N_12427);
nor U12614 (N_12614,N_12383,N_12453);
xnor U12615 (N_12615,N_12403,N_12382);
xor U12616 (N_12616,N_12488,N_12442);
and U12617 (N_12617,N_12496,N_12471);
and U12618 (N_12618,N_12442,N_12416);
or U12619 (N_12619,N_12421,N_12472);
nand U12620 (N_12620,N_12445,N_12497);
nor U12621 (N_12621,N_12378,N_12472);
nor U12622 (N_12622,N_12492,N_12412);
and U12623 (N_12623,N_12469,N_12479);
xnor U12624 (N_12624,N_12432,N_12447);
or U12625 (N_12625,N_12565,N_12577);
or U12626 (N_12626,N_12620,N_12535);
and U12627 (N_12627,N_12573,N_12513);
or U12628 (N_12628,N_12509,N_12517);
or U12629 (N_12629,N_12603,N_12562);
nand U12630 (N_12630,N_12530,N_12623);
or U12631 (N_12631,N_12518,N_12540);
and U12632 (N_12632,N_12617,N_12606);
nor U12633 (N_12633,N_12571,N_12561);
nor U12634 (N_12634,N_12549,N_12615);
and U12635 (N_12635,N_12546,N_12578);
or U12636 (N_12636,N_12526,N_12541);
and U12637 (N_12637,N_12551,N_12527);
and U12638 (N_12638,N_12503,N_12575);
or U12639 (N_12639,N_12579,N_12607);
nor U12640 (N_12640,N_12563,N_12505);
xor U12641 (N_12641,N_12616,N_12609);
xor U12642 (N_12642,N_12508,N_12512);
nor U12643 (N_12643,N_12608,N_12558);
and U12644 (N_12644,N_12548,N_12582);
nor U12645 (N_12645,N_12572,N_12554);
xnor U12646 (N_12646,N_12566,N_12567);
nand U12647 (N_12647,N_12515,N_12506);
nor U12648 (N_12648,N_12531,N_12619);
xnor U12649 (N_12649,N_12590,N_12564);
or U12650 (N_12650,N_12595,N_12502);
xnor U12651 (N_12651,N_12592,N_12585);
xor U12652 (N_12652,N_12611,N_12574);
xor U12653 (N_12653,N_12604,N_12613);
nor U12654 (N_12654,N_12587,N_12538);
or U12655 (N_12655,N_12624,N_12622);
xnor U12656 (N_12656,N_12570,N_12599);
or U12657 (N_12657,N_12522,N_12507);
and U12658 (N_12658,N_12610,N_12542);
nand U12659 (N_12659,N_12576,N_12614);
and U12660 (N_12660,N_12524,N_12591);
nor U12661 (N_12661,N_12580,N_12500);
or U12662 (N_12662,N_12553,N_12583);
xor U12663 (N_12663,N_12501,N_12534);
and U12664 (N_12664,N_12525,N_12504);
nor U12665 (N_12665,N_12516,N_12514);
nor U12666 (N_12666,N_12533,N_12543);
and U12667 (N_12667,N_12556,N_12597);
nand U12668 (N_12668,N_12569,N_12547);
or U12669 (N_12669,N_12539,N_12511);
nand U12670 (N_12670,N_12621,N_12605);
nand U12671 (N_12671,N_12588,N_12602);
and U12672 (N_12672,N_12557,N_12555);
or U12673 (N_12673,N_12600,N_12532);
xor U12674 (N_12674,N_12618,N_12559);
nand U12675 (N_12675,N_12581,N_12529);
and U12676 (N_12676,N_12545,N_12589);
nor U12677 (N_12677,N_12523,N_12596);
xor U12678 (N_12678,N_12568,N_12528);
xor U12679 (N_12679,N_12536,N_12510);
nor U12680 (N_12680,N_12560,N_12519);
xnor U12681 (N_12681,N_12544,N_12537);
nor U12682 (N_12682,N_12521,N_12520);
or U12683 (N_12683,N_12552,N_12586);
nand U12684 (N_12684,N_12550,N_12594);
nand U12685 (N_12685,N_12612,N_12598);
or U12686 (N_12686,N_12601,N_12593);
and U12687 (N_12687,N_12584,N_12562);
nand U12688 (N_12688,N_12537,N_12623);
nor U12689 (N_12689,N_12617,N_12539);
nor U12690 (N_12690,N_12543,N_12597);
nand U12691 (N_12691,N_12573,N_12596);
nor U12692 (N_12692,N_12527,N_12624);
xnor U12693 (N_12693,N_12515,N_12569);
nor U12694 (N_12694,N_12556,N_12534);
xor U12695 (N_12695,N_12532,N_12569);
nand U12696 (N_12696,N_12611,N_12530);
nand U12697 (N_12697,N_12546,N_12543);
and U12698 (N_12698,N_12577,N_12510);
nor U12699 (N_12699,N_12544,N_12548);
xor U12700 (N_12700,N_12583,N_12563);
nor U12701 (N_12701,N_12579,N_12566);
or U12702 (N_12702,N_12504,N_12517);
nand U12703 (N_12703,N_12545,N_12558);
xor U12704 (N_12704,N_12527,N_12580);
and U12705 (N_12705,N_12500,N_12614);
xnor U12706 (N_12706,N_12595,N_12539);
or U12707 (N_12707,N_12504,N_12599);
nor U12708 (N_12708,N_12507,N_12511);
and U12709 (N_12709,N_12523,N_12607);
xor U12710 (N_12710,N_12560,N_12529);
and U12711 (N_12711,N_12515,N_12573);
xor U12712 (N_12712,N_12551,N_12549);
or U12713 (N_12713,N_12616,N_12540);
and U12714 (N_12714,N_12507,N_12525);
or U12715 (N_12715,N_12509,N_12555);
and U12716 (N_12716,N_12571,N_12621);
or U12717 (N_12717,N_12533,N_12617);
nor U12718 (N_12718,N_12548,N_12574);
and U12719 (N_12719,N_12608,N_12609);
nand U12720 (N_12720,N_12578,N_12616);
nor U12721 (N_12721,N_12565,N_12544);
nor U12722 (N_12722,N_12517,N_12555);
and U12723 (N_12723,N_12559,N_12588);
and U12724 (N_12724,N_12533,N_12623);
and U12725 (N_12725,N_12594,N_12586);
nand U12726 (N_12726,N_12619,N_12566);
nor U12727 (N_12727,N_12590,N_12556);
or U12728 (N_12728,N_12537,N_12548);
nand U12729 (N_12729,N_12594,N_12576);
xor U12730 (N_12730,N_12566,N_12591);
nor U12731 (N_12731,N_12505,N_12576);
nand U12732 (N_12732,N_12525,N_12587);
nand U12733 (N_12733,N_12605,N_12588);
nor U12734 (N_12734,N_12541,N_12523);
xnor U12735 (N_12735,N_12538,N_12511);
and U12736 (N_12736,N_12515,N_12526);
xnor U12737 (N_12737,N_12524,N_12584);
nor U12738 (N_12738,N_12521,N_12602);
and U12739 (N_12739,N_12558,N_12522);
nor U12740 (N_12740,N_12579,N_12622);
nand U12741 (N_12741,N_12580,N_12622);
and U12742 (N_12742,N_12594,N_12503);
xnor U12743 (N_12743,N_12523,N_12554);
xor U12744 (N_12744,N_12531,N_12527);
xor U12745 (N_12745,N_12521,N_12553);
nor U12746 (N_12746,N_12529,N_12590);
or U12747 (N_12747,N_12517,N_12578);
nor U12748 (N_12748,N_12605,N_12575);
or U12749 (N_12749,N_12611,N_12553);
nor U12750 (N_12750,N_12717,N_12654);
xor U12751 (N_12751,N_12740,N_12700);
and U12752 (N_12752,N_12636,N_12715);
xor U12753 (N_12753,N_12704,N_12660);
or U12754 (N_12754,N_12659,N_12625);
xor U12755 (N_12755,N_12698,N_12670);
nand U12756 (N_12756,N_12734,N_12653);
xnor U12757 (N_12757,N_12741,N_12747);
nand U12758 (N_12758,N_12690,N_12629);
and U12759 (N_12759,N_12724,N_12693);
or U12760 (N_12760,N_12664,N_12637);
nor U12761 (N_12761,N_12682,N_12691);
nand U12762 (N_12762,N_12671,N_12735);
or U12763 (N_12763,N_12685,N_12721);
and U12764 (N_12764,N_12661,N_12650);
or U12765 (N_12765,N_12713,N_12710);
or U12766 (N_12766,N_12663,N_12729);
xor U12767 (N_12767,N_12667,N_12728);
nor U12768 (N_12768,N_12695,N_12744);
and U12769 (N_12769,N_12697,N_12716);
nor U12770 (N_12770,N_12677,N_12687);
and U12771 (N_12771,N_12706,N_12648);
or U12772 (N_12772,N_12632,N_12641);
nor U12773 (N_12773,N_12646,N_12733);
nor U12774 (N_12774,N_12643,N_12631);
nand U12775 (N_12775,N_12658,N_12694);
and U12776 (N_12776,N_12652,N_12678);
nor U12777 (N_12777,N_12692,N_12718);
or U12778 (N_12778,N_12679,N_12703);
nor U12779 (N_12779,N_12651,N_12688);
nor U12780 (N_12780,N_12676,N_12745);
xor U12781 (N_12781,N_12668,N_12645);
nand U12782 (N_12782,N_12674,N_12673);
nand U12783 (N_12783,N_12689,N_12705);
nor U12784 (N_12784,N_12746,N_12630);
or U12785 (N_12785,N_12627,N_12626);
nand U12786 (N_12786,N_12657,N_12701);
or U12787 (N_12787,N_12649,N_12708);
xor U12788 (N_12788,N_12711,N_12638);
nor U12789 (N_12789,N_12712,N_12748);
or U12790 (N_12790,N_12749,N_12655);
nor U12791 (N_12791,N_12635,N_12666);
xnor U12792 (N_12792,N_12699,N_12739);
xor U12793 (N_12793,N_12714,N_12656);
xnor U12794 (N_12794,N_12742,N_12640);
or U12795 (N_12795,N_12633,N_12743);
xor U12796 (N_12796,N_12730,N_12634);
nor U12797 (N_12797,N_12628,N_12672);
nor U12798 (N_12798,N_12686,N_12639);
nand U12799 (N_12799,N_12702,N_12669);
xnor U12800 (N_12800,N_12684,N_12683);
xor U12801 (N_12801,N_12732,N_12727);
nand U12802 (N_12802,N_12731,N_12725);
nor U12803 (N_12803,N_12738,N_12722);
xnor U12804 (N_12804,N_12696,N_12719);
nor U12805 (N_12805,N_12709,N_12681);
and U12806 (N_12806,N_12647,N_12642);
and U12807 (N_12807,N_12720,N_12707);
xnor U12808 (N_12808,N_12726,N_12680);
xnor U12809 (N_12809,N_12675,N_12662);
and U12810 (N_12810,N_12737,N_12723);
and U12811 (N_12811,N_12665,N_12644);
or U12812 (N_12812,N_12736,N_12667);
nand U12813 (N_12813,N_12741,N_12719);
and U12814 (N_12814,N_12738,N_12678);
and U12815 (N_12815,N_12666,N_12731);
xnor U12816 (N_12816,N_12680,N_12728);
and U12817 (N_12817,N_12689,N_12709);
and U12818 (N_12818,N_12748,N_12693);
and U12819 (N_12819,N_12719,N_12633);
xnor U12820 (N_12820,N_12712,N_12646);
nand U12821 (N_12821,N_12717,N_12644);
xor U12822 (N_12822,N_12632,N_12655);
or U12823 (N_12823,N_12686,N_12668);
and U12824 (N_12824,N_12654,N_12689);
xnor U12825 (N_12825,N_12712,N_12686);
nor U12826 (N_12826,N_12740,N_12653);
xor U12827 (N_12827,N_12667,N_12666);
and U12828 (N_12828,N_12628,N_12636);
nor U12829 (N_12829,N_12731,N_12696);
nand U12830 (N_12830,N_12681,N_12663);
xor U12831 (N_12831,N_12625,N_12749);
or U12832 (N_12832,N_12697,N_12679);
xnor U12833 (N_12833,N_12715,N_12711);
nor U12834 (N_12834,N_12738,N_12693);
nor U12835 (N_12835,N_12730,N_12743);
and U12836 (N_12836,N_12706,N_12685);
and U12837 (N_12837,N_12683,N_12634);
and U12838 (N_12838,N_12690,N_12665);
or U12839 (N_12839,N_12634,N_12741);
xor U12840 (N_12840,N_12642,N_12645);
and U12841 (N_12841,N_12698,N_12681);
and U12842 (N_12842,N_12628,N_12645);
and U12843 (N_12843,N_12744,N_12626);
or U12844 (N_12844,N_12688,N_12643);
nor U12845 (N_12845,N_12682,N_12678);
and U12846 (N_12846,N_12748,N_12699);
or U12847 (N_12847,N_12658,N_12746);
and U12848 (N_12848,N_12632,N_12668);
nand U12849 (N_12849,N_12717,N_12670);
nor U12850 (N_12850,N_12728,N_12675);
and U12851 (N_12851,N_12727,N_12642);
or U12852 (N_12852,N_12640,N_12653);
xor U12853 (N_12853,N_12748,N_12704);
and U12854 (N_12854,N_12715,N_12695);
nor U12855 (N_12855,N_12731,N_12707);
and U12856 (N_12856,N_12635,N_12651);
nor U12857 (N_12857,N_12744,N_12683);
or U12858 (N_12858,N_12696,N_12701);
or U12859 (N_12859,N_12652,N_12631);
or U12860 (N_12860,N_12716,N_12746);
or U12861 (N_12861,N_12685,N_12651);
or U12862 (N_12862,N_12658,N_12729);
xor U12863 (N_12863,N_12679,N_12647);
nand U12864 (N_12864,N_12662,N_12742);
nor U12865 (N_12865,N_12718,N_12707);
nor U12866 (N_12866,N_12732,N_12637);
nor U12867 (N_12867,N_12714,N_12718);
xor U12868 (N_12868,N_12630,N_12709);
nand U12869 (N_12869,N_12689,N_12642);
xor U12870 (N_12870,N_12677,N_12669);
nand U12871 (N_12871,N_12675,N_12697);
nor U12872 (N_12872,N_12643,N_12743);
nor U12873 (N_12873,N_12701,N_12748);
xor U12874 (N_12874,N_12643,N_12719);
nor U12875 (N_12875,N_12788,N_12817);
xnor U12876 (N_12876,N_12868,N_12766);
or U12877 (N_12877,N_12785,N_12815);
or U12878 (N_12878,N_12825,N_12800);
or U12879 (N_12879,N_12750,N_12813);
nand U12880 (N_12880,N_12839,N_12762);
nor U12881 (N_12881,N_12824,N_12768);
or U12882 (N_12882,N_12793,N_12756);
xnor U12883 (N_12883,N_12866,N_12770);
nand U12884 (N_12884,N_12847,N_12852);
nor U12885 (N_12885,N_12761,N_12832);
nor U12886 (N_12886,N_12873,N_12810);
or U12887 (N_12887,N_12821,N_12843);
or U12888 (N_12888,N_12780,N_12872);
nand U12889 (N_12889,N_12794,N_12833);
or U12890 (N_12890,N_12850,N_12798);
and U12891 (N_12891,N_12835,N_12755);
nor U12892 (N_12892,N_12757,N_12784);
or U12893 (N_12893,N_12830,N_12857);
xor U12894 (N_12894,N_12865,N_12860);
nand U12895 (N_12895,N_12783,N_12797);
nor U12896 (N_12896,N_12804,N_12816);
nand U12897 (N_12897,N_12769,N_12841);
or U12898 (N_12898,N_12751,N_12811);
xor U12899 (N_12899,N_12838,N_12764);
and U12900 (N_12900,N_12808,N_12782);
or U12901 (N_12901,N_12807,N_12760);
xor U12902 (N_12902,N_12829,N_12767);
and U12903 (N_12903,N_12846,N_12796);
and U12904 (N_12904,N_12859,N_12856);
xnor U12905 (N_12905,N_12790,N_12781);
xor U12906 (N_12906,N_12871,N_12848);
and U12907 (N_12907,N_12840,N_12864);
nor U12908 (N_12908,N_12836,N_12822);
nand U12909 (N_12909,N_12845,N_12758);
or U12910 (N_12910,N_12814,N_12826);
and U12911 (N_12911,N_12851,N_12773);
nor U12912 (N_12912,N_12753,N_12862);
nand U12913 (N_12913,N_12805,N_12752);
xnor U12914 (N_12914,N_12775,N_12763);
xor U12915 (N_12915,N_12870,N_12795);
nor U12916 (N_12916,N_12831,N_12820);
and U12917 (N_12917,N_12771,N_12819);
nand U12918 (N_12918,N_12792,N_12834);
nand U12919 (N_12919,N_12799,N_12854);
nand U12920 (N_12920,N_12806,N_12809);
nor U12921 (N_12921,N_12772,N_12827);
xor U12922 (N_12922,N_12874,N_12791);
and U12923 (N_12923,N_12802,N_12869);
nand U12924 (N_12924,N_12858,N_12828);
nor U12925 (N_12925,N_12776,N_12863);
nor U12926 (N_12926,N_12765,N_12774);
and U12927 (N_12927,N_12801,N_12844);
xnor U12928 (N_12928,N_12853,N_12812);
and U12929 (N_12929,N_12861,N_12842);
nand U12930 (N_12930,N_12823,N_12777);
xnor U12931 (N_12931,N_12867,N_12789);
xnor U12932 (N_12932,N_12849,N_12754);
nand U12933 (N_12933,N_12818,N_12837);
nor U12934 (N_12934,N_12855,N_12803);
or U12935 (N_12935,N_12779,N_12778);
and U12936 (N_12936,N_12759,N_12786);
nand U12937 (N_12937,N_12787,N_12849);
nand U12938 (N_12938,N_12858,N_12760);
xnor U12939 (N_12939,N_12802,N_12826);
nand U12940 (N_12940,N_12756,N_12831);
nand U12941 (N_12941,N_12863,N_12802);
nand U12942 (N_12942,N_12840,N_12852);
xnor U12943 (N_12943,N_12780,N_12825);
xor U12944 (N_12944,N_12808,N_12795);
or U12945 (N_12945,N_12799,N_12796);
nor U12946 (N_12946,N_12835,N_12857);
or U12947 (N_12947,N_12800,N_12755);
nor U12948 (N_12948,N_12786,N_12831);
or U12949 (N_12949,N_12765,N_12784);
or U12950 (N_12950,N_12803,N_12836);
or U12951 (N_12951,N_12851,N_12762);
nor U12952 (N_12952,N_12760,N_12831);
nand U12953 (N_12953,N_12867,N_12768);
nand U12954 (N_12954,N_12773,N_12820);
and U12955 (N_12955,N_12813,N_12756);
or U12956 (N_12956,N_12841,N_12873);
nor U12957 (N_12957,N_12826,N_12858);
and U12958 (N_12958,N_12762,N_12823);
xor U12959 (N_12959,N_12789,N_12777);
nand U12960 (N_12960,N_12807,N_12857);
xor U12961 (N_12961,N_12801,N_12770);
or U12962 (N_12962,N_12766,N_12762);
or U12963 (N_12963,N_12819,N_12762);
or U12964 (N_12964,N_12759,N_12795);
or U12965 (N_12965,N_12802,N_12756);
xor U12966 (N_12966,N_12760,N_12839);
xor U12967 (N_12967,N_12817,N_12865);
nor U12968 (N_12968,N_12873,N_12859);
nor U12969 (N_12969,N_12794,N_12829);
or U12970 (N_12970,N_12761,N_12784);
xor U12971 (N_12971,N_12831,N_12865);
nand U12972 (N_12972,N_12793,N_12828);
or U12973 (N_12973,N_12753,N_12848);
xor U12974 (N_12974,N_12782,N_12843);
nand U12975 (N_12975,N_12798,N_12815);
nand U12976 (N_12976,N_12767,N_12820);
nand U12977 (N_12977,N_12821,N_12808);
nor U12978 (N_12978,N_12854,N_12780);
xor U12979 (N_12979,N_12810,N_12862);
nor U12980 (N_12980,N_12772,N_12869);
or U12981 (N_12981,N_12857,N_12811);
nand U12982 (N_12982,N_12770,N_12771);
or U12983 (N_12983,N_12845,N_12772);
nor U12984 (N_12984,N_12816,N_12774);
or U12985 (N_12985,N_12774,N_12779);
xor U12986 (N_12986,N_12798,N_12755);
xnor U12987 (N_12987,N_12827,N_12858);
and U12988 (N_12988,N_12855,N_12840);
xnor U12989 (N_12989,N_12790,N_12833);
nor U12990 (N_12990,N_12808,N_12815);
nor U12991 (N_12991,N_12779,N_12872);
xnor U12992 (N_12992,N_12771,N_12834);
or U12993 (N_12993,N_12787,N_12831);
or U12994 (N_12994,N_12769,N_12864);
nor U12995 (N_12995,N_12847,N_12826);
nor U12996 (N_12996,N_12863,N_12807);
xor U12997 (N_12997,N_12834,N_12863);
and U12998 (N_12998,N_12784,N_12832);
nor U12999 (N_12999,N_12774,N_12826);
nor U13000 (N_13000,N_12984,N_12992);
xnor U13001 (N_13001,N_12939,N_12876);
and U13002 (N_13002,N_12978,N_12981);
or U13003 (N_13003,N_12943,N_12965);
or U13004 (N_13004,N_12923,N_12997);
or U13005 (N_13005,N_12950,N_12947);
xnor U13006 (N_13006,N_12916,N_12956);
xor U13007 (N_13007,N_12961,N_12878);
xnor U13008 (N_13008,N_12946,N_12974);
nor U13009 (N_13009,N_12910,N_12907);
xor U13010 (N_13010,N_12970,N_12881);
or U13011 (N_13011,N_12914,N_12976);
and U13012 (N_13012,N_12903,N_12975);
or U13013 (N_13013,N_12888,N_12902);
and U13014 (N_13014,N_12882,N_12936);
nor U13015 (N_13015,N_12924,N_12959);
and U13016 (N_13016,N_12889,N_12900);
and U13017 (N_13017,N_12886,N_12894);
nor U13018 (N_13018,N_12987,N_12990);
and U13019 (N_13019,N_12906,N_12962);
nand U13020 (N_13020,N_12989,N_12945);
nand U13021 (N_13021,N_12938,N_12931);
xor U13022 (N_13022,N_12905,N_12994);
or U13023 (N_13023,N_12898,N_12968);
or U13024 (N_13024,N_12957,N_12911);
xor U13025 (N_13025,N_12944,N_12885);
nand U13026 (N_13026,N_12896,N_12913);
or U13027 (N_13027,N_12912,N_12948);
nor U13028 (N_13028,N_12988,N_12937);
nand U13029 (N_13029,N_12929,N_12891);
xor U13030 (N_13030,N_12879,N_12935);
or U13031 (N_13031,N_12960,N_12986);
or U13032 (N_13032,N_12892,N_12991);
and U13033 (N_13033,N_12915,N_12880);
and U13034 (N_13034,N_12996,N_12999);
nand U13035 (N_13035,N_12998,N_12893);
xnor U13036 (N_13036,N_12955,N_12979);
nor U13037 (N_13037,N_12890,N_12899);
xor U13038 (N_13038,N_12908,N_12941);
or U13039 (N_13039,N_12993,N_12977);
nand U13040 (N_13040,N_12928,N_12930);
nor U13041 (N_13041,N_12958,N_12932);
nand U13042 (N_13042,N_12884,N_12887);
or U13043 (N_13043,N_12954,N_12966);
nor U13044 (N_13044,N_12904,N_12940);
nand U13045 (N_13045,N_12877,N_12895);
nand U13046 (N_13046,N_12933,N_12963);
nand U13047 (N_13047,N_12926,N_12973);
nand U13048 (N_13048,N_12925,N_12953);
xnor U13049 (N_13049,N_12969,N_12934);
nand U13050 (N_13050,N_12901,N_12918);
nand U13051 (N_13051,N_12897,N_12917);
xnor U13052 (N_13052,N_12995,N_12971);
or U13053 (N_13053,N_12980,N_12967);
nand U13054 (N_13054,N_12949,N_12942);
xor U13055 (N_13055,N_12983,N_12875);
nor U13056 (N_13056,N_12927,N_12921);
nand U13057 (N_13057,N_12920,N_12952);
and U13058 (N_13058,N_12985,N_12922);
xnor U13059 (N_13059,N_12964,N_12972);
nand U13060 (N_13060,N_12982,N_12951);
nand U13061 (N_13061,N_12919,N_12883);
and U13062 (N_13062,N_12909,N_12993);
nand U13063 (N_13063,N_12967,N_12988);
nand U13064 (N_13064,N_12949,N_12998);
and U13065 (N_13065,N_12967,N_12993);
nor U13066 (N_13066,N_12987,N_12998);
xnor U13067 (N_13067,N_12974,N_12877);
xor U13068 (N_13068,N_12956,N_12951);
or U13069 (N_13069,N_12972,N_12998);
nor U13070 (N_13070,N_12946,N_12943);
nand U13071 (N_13071,N_12897,N_12977);
nand U13072 (N_13072,N_12953,N_12946);
xnor U13073 (N_13073,N_12894,N_12879);
nor U13074 (N_13074,N_12927,N_12943);
or U13075 (N_13075,N_12904,N_12945);
and U13076 (N_13076,N_12885,N_12948);
nand U13077 (N_13077,N_12986,N_12934);
and U13078 (N_13078,N_12930,N_12963);
xor U13079 (N_13079,N_12927,N_12983);
nand U13080 (N_13080,N_12954,N_12946);
and U13081 (N_13081,N_12991,N_12990);
nor U13082 (N_13082,N_12876,N_12962);
and U13083 (N_13083,N_12900,N_12983);
nand U13084 (N_13084,N_12881,N_12952);
or U13085 (N_13085,N_12988,N_12902);
nor U13086 (N_13086,N_12895,N_12943);
and U13087 (N_13087,N_12877,N_12875);
and U13088 (N_13088,N_12959,N_12880);
and U13089 (N_13089,N_12937,N_12991);
and U13090 (N_13090,N_12918,N_12903);
xor U13091 (N_13091,N_12988,N_12955);
nand U13092 (N_13092,N_12978,N_12878);
and U13093 (N_13093,N_12887,N_12956);
nor U13094 (N_13094,N_12961,N_12900);
xor U13095 (N_13095,N_12991,N_12984);
nand U13096 (N_13096,N_12933,N_12951);
or U13097 (N_13097,N_12984,N_12963);
xor U13098 (N_13098,N_12953,N_12880);
xor U13099 (N_13099,N_12987,N_12911);
or U13100 (N_13100,N_12890,N_12999);
nand U13101 (N_13101,N_12967,N_12983);
nand U13102 (N_13102,N_12904,N_12880);
xnor U13103 (N_13103,N_12877,N_12948);
or U13104 (N_13104,N_12951,N_12953);
xor U13105 (N_13105,N_12941,N_12931);
xnor U13106 (N_13106,N_12952,N_12934);
or U13107 (N_13107,N_12894,N_12963);
nand U13108 (N_13108,N_12944,N_12995);
nand U13109 (N_13109,N_12965,N_12979);
nor U13110 (N_13110,N_12947,N_12909);
and U13111 (N_13111,N_12958,N_12967);
or U13112 (N_13112,N_12980,N_12961);
and U13113 (N_13113,N_12931,N_12910);
xor U13114 (N_13114,N_12960,N_12939);
or U13115 (N_13115,N_12980,N_12915);
nand U13116 (N_13116,N_12875,N_12970);
xor U13117 (N_13117,N_12954,N_12945);
and U13118 (N_13118,N_12880,N_12914);
or U13119 (N_13119,N_12950,N_12955);
nand U13120 (N_13120,N_12993,N_12974);
nand U13121 (N_13121,N_12924,N_12962);
nor U13122 (N_13122,N_12936,N_12963);
xor U13123 (N_13123,N_12973,N_12965);
and U13124 (N_13124,N_12974,N_12932);
and U13125 (N_13125,N_13116,N_13101);
and U13126 (N_13126,N_13067,N_13071);
or U13127 (N_13127,N_13049,N_13023);
xnor U13128 (N_13128,N_13094,N_13001);
xor U13129 (N_13129,N_13099,N_13084);
or U13130 (N_13130,N_13098,N_13031);
and U13131 (N_13131,N_13075,N_13006);
nor U13132 (N_13132,N_13106,N_13062);
nand U13133 (N_13133,N_13038,N_13081);
or U13134 (N_13134,N_13059,N_13109);
xnor U13135 (N_13135,N_13057,N_13121);
nand U13136 (N_13136,N_13072,N_13043);
or U13137 (N_13137,N_13092,N_13015);
nor U13138 (N_13138,N_13060,N_13091);
nand U13139 (N_13139,N_13083,N_13028);
nor U13140 (N_13140,N_13063,N_13024);
xor U13141 (N_13141,N_13104,N_13102);
xor U13142 (N_13142,N_13004,N_13120);
or U13143 (N_13143,N_13090,N_13052);
and U13144 (N_13144,N_13086,N_13111);
or U13145 (N_13145,N_13118,N_13051);
or U13146 (N_13146,N_13113,N_13093);
xor U13147 (N_13147,N_13122,N_13068);
nand U13148 (N_13148,N_13074,N_13019);
and U13149 (N_13149,N_13009,N_13014);
xnor U13150 (N_13150,N_13034,N_13008);
xor U13151 (N_13151,N_13030,N_13105);
nand U13152 (N_13152,N_13100,N_13089);
nand U13153 (N_13153,N_13087,N_13026);
or U13154 (N_13154,N_13058,N_13069);
and U13155 (N_13155,N_13123,N_13005);
xnor U13156 (N_13156,N_13112,N_13103);
nand U13157 (N_13157,N_13065,N_13044);
xor U13158 (N_13158,N_13036,N_13070);
nand U13159 (N_13159,N_13061,N_13037);
nor U13160 (N_13160,N_13117,N_13055);
or U13161 (N_13161,N_13003,N_13045);
and U13162 (N_13162,N_13097,N_13064);
or U13163 (N_13163,N_13047,N_13076);
nand U13164 (N_13164,N_13040,N_13078);
or U13165 (N_13165,N_13011,N_13050);
and U13166 (N_13166,N_13119,N_13018);
and U13167 (N_13167,N_13096,N_13027);
xor U13168 (N_13168,N_13088,N_13002);
xnor U13169 (N_13169,N_13022,N_13032);
xor U13170 (N_13170,N_13016,N_13042);
xor U13171 (N_13171,N_13108,N_13114);
nand U13172 (N_13172,N_13066,N_13073);
nor U13173 (N_13173,N_13124,N_13013);
nor U13174 (N_13174,N_13085,N_13095);
nor U13175 (N_13175,N_13082,N_13007);
xor U13176 (N_13176,N_13020,N_13012);
nor U13177 (N_13177,N_13035,N_13080);
or U13178 (N_13178,N_13046,N_13056);
and U13179 (N_13179,N_13048,N_13079);
nand U13180 (N_13180,N_13110,N_13054);
nor U13181 (N_13181,N_13010,N_13029);
and U13182 (N_13182,N_13025,N_13115);
nand U13183 (N_13183,N_13077,N_13041);
or U13184 (N_13184,N_13033,N_13000);
and U13185 (N_13185,N_13039,N_13053);
nand U13186 (N_13186,N_13017,N_13021);
nand U13187 (N_13187,N_13107,N_13075);
and U13188 (N_13188,N_13093,N_13111);
and U13189 (N_13189,N_13045,N_13093);
nor U13190 (N_13190,N_13041,N_13050);
nor U13191 (N_13191,N_13106,N_13089);
xor U13192 (N_13192,N_13067,N_13025);
xor U13193 (N_13193,N_13060,N_13097);
nand U13194 (N_13194,N_13092,N_13088);
nand U13195 (N_13195,N_13079,N_13065);
xnor U13196 (N_13196,N_13010,N_13049);
xnor U13197 (N_13197,N_13124,N_13037);
and U13198 (N_13198,N_13062,N_13098);
nand U13199 (N_13199,N_13095,N_13017);
xnor U13200 (N_13200,N_13065,N_13095);
nand U13201 (N_13201,N_13090,N_13008);
xnor U13202 (N_13202,N_13081,N_13095);
and U13203 (N_13203,N_13089,N_13063);
nand U13204 (N_13204,N_13044,N_13000);
or U13205 (N_13205,N_13123,N_13081);
or U13206 (N_13206,N_13004,N_13089);
and U13207 (N_13207,N_13122,N_13058);
or U13208 (N_13208,N_13028,N_13026);
or U13209 (N_13209,N_13086,N_13067);
xnor U13210 (N_13210,N_13030,N_13019);
nor U13211 (N_13211,N_13016,N_13080);
and U13212 (N_13212,N_13046,N_13120);
and U13213 (N_13213,N_13072,N_13112);
nand U13214 (N_13214,N_13099,N_13091);
or U13215 (N_13215,N_13051,N_13048);
nand U13216 (N_13216,N_13052,N_13019);
xnor U13217 (N_13217,N_13022,N_13083);
or U13218 (N_13218,N_13051,N_13084);
nor U13219 (N_13219,N_13090,N_13041);
or U13220 (N_13220,N_13095,N_13092);
xor U13221 (N_13221,N_13074,N_13048);
and U13222 (N_13222,N_13063,N_13074);
xor U13223 (N_13223,N_13079,N_13107);
nor U13224 (N_13224,N_13038,N_13059);
xnor U13225 (N_13225,N_13072,N_13045);
or U13226 (N_13226,N_13117,N_13072);
and U13227 (N_13227,N_13086,N_13049);
nor U13228 (N_13228,N_13025,N_13076);
nand U13229 (N_13229,N_13100,N_13106);
nor U13230 (N_13230,N_13027,N_13083);
or U13231 (N_13231,N_13105,N_13084);
nand U13232 (N_13232,N_13059,N_13076);
and U13233 (N_13233,N_13091,N_13078);
and U13234 (N_13234,N_13068,N_13017);
nand U13235 (N_13235,N_13114,N_13023);
xnor U13236 (N_13236,N_13077,N_13109);
or U13237 (N_13237,N_13101,N_13008);
nand U13238 (N_13238,N_13067,N_13007);
xor U13239 (N_13239,N_13115,N_13057);
nand U13240 (N_13240,N_13104,N_13043);
xnor U13241 (N_13241,N_13038,N_13088);
and U13242 (N_13242,N_13118,N_13110);
or U13243 (N_13243,N_13065,N_13062);
or U13244 (N_13244,N_13081,N_13031);
nor U13245 (N_13245,N_13101,N_13038);
nand U13246 (N_13246,N_13090,N_13032);
or U13247 (N_13247,N_13079,N_13057);
xor U13248 (N_13248,N_13012,N_13088);
or U13249 (N_13249,N_13034,N_13012);
nand U13250 (N_13250,N_13232,N_13166);
nor U13251 (N_13251,N_13172,N_13208);
nand U13252 (N_13252,N_13164,N_13244);
nand U13253 (N_13253,N_13138,N_13204);
or U13254 (N_13254,N_13202,N_13245);
nand U13255 (N_13255,N_13219,N_13185);
xor U13256 (N_13256,N_13129,N_13225);
nand U13257 (N_13257,N_13151,N_13141);
nor U13258 (N_13258,N_13159,N_13228);
or U13259 (N_13259,N_13125,N_13193);
nor U13260 (N_13260,N_13189,N_13134);
and U13261 (N_13261,N_13221,N_13184);
or U13262 (N_13262,N_13145,N_13139);
nand U13263 (N_13263,N_13161,N_13143);
or U13264 (N_13264,N_13224,N_13194);
or U13265 (N_13265,N_13237,N_13212);
nand U13266 (N_13266,N_13190,N_13222);
nand U13267 (N_13267,N_13183,N_13211);
nand U13268 (N_13268,N_13127,N_13176);
or U13269 (N_13269,N_13210,N_13249);
and U13270 (N_13270,N_13246,N_13216);
nand U13271 (N_13271,N_13170,N_13180);
xor U13272 (N_13272,N_13186,N_13135);
nand U13273 (N_13273,N_13206,N_13217);
nor U13274 (N_13274,N_13243,N_13230);
xor U13275 (N_13275,N_13160,N_13226);
nor U13276 (N_13276,N_13240,N_13150);
or U13277 (N_13277,N_13142,N_13199);
nand U13278 (N_13278,N_13136,N_13148);
nand U13279 (N_13279,N_13152,N_13131);
or U13280 (N_13280,N_13165,N_13144);
nand U13281 (N_13281,N_13173,N_13153);
nand U13282 (N_13282,N_13220,N_13223);
nand U13283 (N_13283,N_13209,N_13179);
or U13284 (N_13284,N_13235,N_13181);
and U13285 (N_13285,N_13157,N_13214);
or U13286 (N_13286,N_13233,N_13147);
nor U13287 (N_13287,N_13207,N_13197);
or U13288 (N_13288,N_13191,N_13187);
xnor U13289 (N_13289,N_13158,N_13198);
or U13290 (N_13290,N_13215,N_13218);
nand U13291 (N_13291,N_13154,N_13203);
and U13292 (N_13292,N_13140,N_13236);
or U13293 (N_13293,N_13155,N_13168);
and U13294 (N_13294,N_13196,N_13231);
and U13295 (N_13295,N_13242,N_13128);
xnor U13296 (N_13296,N_13234,N_13182);
or U13297 (N_13297,N_13146,N_13239);
nand U13298 (N_13298,N_13213,N_13133);
nand U13299 (N_13299,N_13126,N_13171);
or U13300 (N_13300,N_13195,N_13174);
nor U13301 (N_13301,N_13132,N_13178);
nand U13302 (N_13302,N_13137,N_13241);
xnor U13303 (N_13303,N_13149,N_13200);
nand U13304 (N_13304,N_13169,N_13227);
nor U13305 (N_13305,N_13130,N_13201);
xnor U13306 (N_13306,N_13162,N_13163);
or U13307 (N_13307,N_13177,N_13192);
and U13308 (N_13308,N_13248,N_13167);
xor U13309 (N_13309,N_13229,N_13156);
or U13310 (N_13310,N_13247,N_13205);
or U13311 (N_13311,N_13175,N_13188);
nor U13312 (N_13312,N_13238,N_13176);
nand U13313 (N_13313,N_13174,N_13228);
and U13314 (N_13314,N_13167,N_13184);
nand U13315 (N_13315,N_13149,N_13228);
nand U13316 (N_13316,N_13187,N_13244);
and U13317 (N_13317,N_13186,N_13239);
or U13318 (N_13318,N_13209,N_13142);
and U13319 (N_13319,N_13198,N_13187);
nand U13320 (N_13320,N_13235,N_13201);
xnor U13321 (N_13321,N_13217,N_13216);
nor U13322 (N_13322,N_13239,N_13196);
nand U13323 (N_13323,N_13127,N_13219);
and U13324 (N_13324,N_13193,N_13162);
or U13325 (N_13325,N_13192,N_13241);
nand U13326 (N_13326,N_13225,N_13218);
xnor U13327 (N_13327,N_13154,N_13241);
xnor U13328 (N_13328,N_13148,N_13213);
or U13329 (N_13329,N_13173,N_13207);
nand U13330 (N_13330,N_13192,N_13217);
nor U13331 (N_13331,N_13151,N_13190);
or U13332 (N_13332,N_13217,N_13243);
nor U13333 (N_13333,N_13133,N_13245);
and U13334 (N_13334,N_13133,N_13183);
nor U13335 (N_13335,N_13247,N_13246);
xor U13336 (N_13336,N_13137,N_13158);
and U13337 (N_13337,N_13244,N_13210);
or U13338 (N_13338,N_13132,N_13244);
and U13339 (N_13339,N_13168,N_13198);
and U13340 (N_13340,N_13161,N_13175);
nor U13341 (N_13341,N_13163,N_13173);
xnor U13342 (N_13342,N_13159,N_13160);
nand U13343 (N_13343,N_13149,N_13236);
nand U13344 (N_13344,N_13239,N_13162);
nand U13345 (N_13345,N_13248,N_13236);
nor U13346 (N_13346,N_13217,N_13179);
nor U13347 (N_13347,N_13186,N_13204);
xnor U13348 (N_13348,N_13174,N_13222);
and U13349 (N_13349,N_13237,N_13247);
or U13350 (N_13350,N_13234,N_13129);
or U13351 (N_13351,N_13150,N_13169);
xnor U13352 (N_13352,N_13139,N_13190);
nand U13353 (N_13353,N_13247,N_13131);
and U13354 (N_13354,N_13229,N_13226);
and U13355 (N_13355,N_13227,N_13187);
xnor U13356 (N_13356,N_13144,N_13140);
nand U13357 (N_13357,N_13220,N_13157);
xnor U13358 (N_13358,N_13235,N_13151);
and U13359 (N_13359,N_13173,N_13223);
xor U13360 (N_13360,N_13248,N_13207);
nor U13361 (N_13361,N_13231,N_13156);
nor U13362 (N_13362,N_13197,N_13181);
xnor U13363 (N_13363,N_13206,N_13177);
xor U13364 (N_13364,N_13241,N_13199);
xnor U13365 (N_13365,N_13207,N_13151);
and U13366 (N_13366,N_13198,N_13178);
and U13367 (N_13367,N_13181,N_13193);
nor U13368 (N_13368,N_13230,N_13130);
and U13369 (N_13369,N_13234,N_13157);
or U13370 (N_13370,N_13205,N_13234);
nor U13371 (N_13371,N_13248,N_13177);
and U13372 (N_13372,N_13150,N_13248);
and U13373 (N_13373,N_13148,N_13229);
or U13374 (N_13374,N_13130,N_13223);
nor U13375 (N_13375,N_13352,N_13259);
and U13376 (N_13376,N_13299,N_13324);
xor U13377 (N_13377,N_13345,N_13374);
and U13378 (N_13378,N_13360,N_13281);
or U13379 (N_13379,N_13250,N_13322);
nand U13380 (N_13380,N_13350,N_13265);
nor U13381 (N_13381,N_13315,N_13316);
or U13382 (N_13382,N_13373,N_13288);
or U13383 (N_13383,N_13252,N_13364);
xor U13384 (N_13384,N_13307,N_13260);
nand U13385 (N_13385,N_13329,N_13349);
nor U13386 (N_13386,N_13358,N_13334);
and U13387 (N_13387,N_13273,N_13268);
nor U13388 (N_13388,N_13256,N_13339);
or U13389 (N_13389,N_13300,N_13279);
xnor U13390 (N_13390,N_13280,N_13310);
and U13391 (N_13391,N_13314,N_13355);
nor U13392 (N_13392,N_13317,N_13289);
xor U13393 (N_13393,N_13342,N_13351);
nand U13394 (N_13394,N_13291,N_13276);
or U13395 (N_13395,N_13326,N_13347);
or U13396 (N_13396,N_13287,N_13292);
nand U13397 (N_13397,N_13284,N_13304);
or U13398 (N_13398,N_13356,N_13264);
or U13399 (N_13399,N_13325,N_13261);
xnor U13400 (N_13400,N_13330,N_13363);
or U13401 (N_13401,N_13362,N_13286);
nand U13402 (N_13402,N_13369,N_13309);
nand U13403 (N_13403,N_13251,N_13366);
and U13404 (N_13404,N_13321,N_13283);
nor U13405 (N_13405,N_13277,N_13295);
nand U13406 (N_13406,N_13253,N_13372);
xor U13407 (N_13407,N_13274,N_13327);
or U13408 (N_13408,N_13343,N_13336);
or U13409 (N_13409,N_13370,N_13319);
and U13410 (N_13410,N_13278,N_13328);
or U13411 (N_13411,N_13272,N_13365);
nand U13412 (N_13412,N_13320,N_13332);
or U13413 (N_13413,N_13294,N_13303);
and U13414 (N_13414,N_13335,N_13312);
xnor U13415 (N_13415,N_13338,N_13257);
or U13416 (N_13416,N_13353,N_13371);
and U13417 (N_13417,N_13301,N_13290);
or U13418 (N_13418,N_13341,N_13331);
nor U13419 (N_13419,N_13275,N_13302);
or U13420 (N_13420,N_13266,N_13346);
nor U13421 (N_13421,N_13270,N_13263);
or U13422 (N_13422,N_13282,N_13311);
and U13423 (N_13423,N_13297,N_13285);
xnor U13424 (N_13424,N_13361,N_13357);
nor U13425 (N_13425,N_13337,N_13255);
and U13426 (N_13426,N_13306,N_13340);
and U13427 (N_13427,N_13258,N_13305);
nor U13428 (N_13428,N_13318,N_13269);
or U13429 (N_13429,N_13296,N_13359);
xnor U13430 (N_13430,N_13354,N_13333);
or U13431 (N_13431,N_13348,N_13298);
nor U13432 (N_13432,N_13262,N_13271);
or U13433 (N_13433,N_13323,N_13254);
xnor U13434 (N_13434,N_13267,N_13313);
and U13435 (N_13435,N_13293,N_13368);
xor U13436 (N_13436,N_13308,N_13367);
nand U13437 (N_13437,N_13344,N_13368);
or U13438 (N_13438,N_13320,N_13371);
xnor U13439 (N_13439,N_13371,N_13314);
nor U13440 (N_13440,N_13293,N_13370);
and U13441 (N_13441,N_13365,N_13355);
and U13442 (N_13442,N_13344,N_13305);
nor U13443 (N_13443,N_13369,N_13284);
nand U13444 (N_13444,N_13327,N_13339);
or U13445 (N_13445,N_13262,N_13311);
and U13446 (N_13446,N_13278,N_13361);
or U13447 (N_13447,N_13261,N_13303);
and U13448 (N_13448,N_13321,N_13295);
xnor U13449 (N_13449,N_13339,N_13324);
nor U13450 (N_13450,N_13330,N_13293);
xor U13451 (N_13451,N_13360,N_13312);
and U13452 (N_13452,N_13364,N_13352);
nand U13453 (N_13453,N_13283,N_13280);
xor U13454 (N_13454,N_13346,N_13357);
xnor U13455 (N_13455,N_13307,N_13315);
or U13456 (N_13456,N_13342,N_13353);
xor U13457 (N_13457,N_13360,N_13269);
xnor U13458 (N_13458,N_13309,N_13363);
and U13459 (N_13459,N_13295,N_13256);
and U13460 (N_13460,N_13346,N_13324);
or U13461 (N_13461,N_13329,N_13332);
xor U13462 (N_13462,N_13315,N_13297);
and U13463 (N_13463,N_13322,N_13341);
xnor U13464 (N_13464,N_13315,N_13303);
nand U13465 (N_13465,N_13302,N_13289);
nand U13466 (N_13466,N_13287,N_13321);
nand U13467 (N_13467,N_13321,N_13345);
nor U13468 (N_13468,N_13270,N_13373);
and U13469 (N_13469,N_13363,N_13340);
nor U13470 (N_13470,N_13336,N_13348);
or U13471 (N_13471,N_13338,N_13285);
xnor U13472 (N_13472,N_13353,N_13364);
and U13473 (N_13473,N_13294,N_13340);
xor U13474 (N_13474,N_13300,N_13250);
or U13475 (N_13475,N_13364,N_13368);
xnor U13476 (N_13476,N_13316,N_13326);
xor U13477 (N_13477,N_13259,N_13310);
nand U13478 (N_13478,N_13271,N_13318);
nor U13479 (N_13479,N_13298,N_13350);
and U13480 (N_13480,N_13314,N_13361);
and U13481 (N_13481,N_13303,N_13283);
xor U13482 (N_13482,N_13279,N_13356);
nor U13483 (N_13483,N_13327,N_13304);
nand U13484 (N_13484,N_13348,N_13339);
nor U13485 (N_13485,N_13320,N_13257);
and U13486 (N_13486,N_13354,N_13318);
and U13487 (N_13487,N_13271,N_13320);
nand U13488 (N_13488,N_13269,N_13349);
nor U13489 (N_13489,N_13332,N_13313);
and U13490 (N_13490,N_13285,N_13256);
or U13491 (N_13491,N_13335,N_13363);
xor U13492 (N_13492,N_13268,N_13331);
nor U13493 (N_13493,N_13370,N_13263);
or U13494 (N_13494,N_13310,N_13297);
xnor U13495 (N_13495,N_13304,N_13252);
nand U13496 (N_13496,N_13341,N_13355);
and U13497 (N_13497,N_13365,N_13268);
or U13498 (N_13498,N_13315,N_13254);
xor U13499 (N_13499,N_13373,N_13255);
xnor U13500 (N_13500,N_13414,N_13483);
and U13501 (N_13501,N_13457,N_13425);
nand U13502 (N_13502,N_13382,N_13491);
nand U13503 (N_13503,N_13380,N_13401);
or U13504 (N_13504,N_13431,N_13490);
nand U13505 (N_13505,N_13443,N_13389);
and U13506 (N_13506,N_13489,N_13424);
or U13507 (N_13507,N_13482,N_13444);
xor U13508 (N_13508,N_13477,N_13473);
nand U13509 (N_13509,N_13390,N_13422);
and U13510 (N_13510,N_13450,N_13497);
nor U13511 (N_13511,N_13452,N_13494);
nor U13512 (N_13512,N_13476,N_13421);
or U13513 (N_13513,N_13384,N_13415);
or U13514 (N_13514,N_13420,N_13432);
nor U13515 (N_13515,N_13498,N_13437);
nand U13516 (N_13516,N_13413,N_13385);
nor U13517 (N_13517,N_13493,N_13469);
nor U13518 (N_13518,N_13449,N_13462);
xnor U13519 (N_13519,N_13471,N_13461);
xor U13520 (N_13520,N_13398,N_13379);
nor U13521 (N_13521,N_13453,N_13427);
xnor U13522 (N_13522,N_13378,N_13439);
nor U13523 (N_13523,N_13438,N_13441);
or U13524 (N_13524,N_13451,N_13492);
nand U13525 (N_13525,N_13377,N_13395);
xor U13526 (N_13526,N_13403,N_13375);
nor U13527 (N_13527,N_13436,N_13468);
nand U13528 (N_13528,N_13404,N_13459);
nor U13529 (N_13529,N_13376,N_13470);
or U13530 (N_13530,N_13411,N_13460);
nor U13531 (N_13531,N_13487,N_13463);
xnor U13532 (N_13532,N_13381,N_13399);
nand U13533 (N_13533,N_13387,N_13406);
or U13534 (N_13534,N_13392,N_13388);
and U13535 (N_13535,N_13408,N_13410);
and U13536 (N_13536,N_13495,N_13496);
nand U13537 (N_13537,N_13446,N_13472);
nand U13538 (N_13538,N_13455,N_13466);
nand U13539 (N_13539,N_13478,N_13423);
xor U13540 (N_13540,N_13391,N_13485);
xnor U13541 (N_13541,N_13430,N_13488);
nand U13542 (N_13542,N_13428,N_13393);
nand U13543 (N_13543,N_13445,N_13475);
or U13544 (N_13544,N_13435,N_13433);
xor U13545 (N_13545,N_13397,N_13442);
nor U13546 (N_13546,N_13440,N_13426);
nor U13547 (N_13547,N_13407,N_13409);
or U13548 (N_13548,N_13480,N_13434);
and U13549 (N_13549,N_13481,N_13429);
and U13550 (N_13550,N_13402,N_13412);
xnor U13551 (N_13551,N_13465,N_13474);
or U13552 (N_13552,N_13419,N_13386);
nor U13553 (N_13553,N_13396,N_13400);
xor U13554 (N_13554,N_13454,N_13484);
and U13555 (N_13555,N_13486,N_13394);
xor U13556 (N_13556,N_13448,N_13418);
and U13557 (N_13557,N_13417,N_13499);
xor U13558 (N_13558,N_13458,N_13405);
and U13559 (N_13559,N_13464,N_13447);
xnor U13560 (N_13560,N_13416,N_13467);
xor U13561 (N_13561,N_13479,N_13383);
or U13562 (N_13562,N_13456,N_13472);
nand U13563 (N_13563,N_13376,N_13386);
and U13564 (N_13564,N_13433,N_13388);
and U13565 (N_13565,N_13451,N_13453);
nor U13566 (N_13566,N_13464,N_13439);
nand U13567 (N_13567,N_13436,N_13443);
xor U13568 (N_13568,N_13470,N_13416);
or U13569 (N_13569,N_13478,N_13432);
nand U13570 (N_13570,N_13497,N_13402);
xor U13571 (N_13571,N_13386,N_13469);
and U13572 (N_13572,N_13394,N_13417);
or U13573 (N_13573,N_13397,N_13416);
and U13574 (N_13574,N_13423,N_13477);
xnor U13575 (N_13575,N_13458,N_13488);
nor U13576 (N_13576,N_13452,N_13474);
and U13577 (N_13577,N_13411,N_13402);
and U13578 (N_13578,N_13448,N_13471);
and U13579 (N_13579,N_13407,N_13446);
nor U13580 (N_13580,N_13400,N_13381);
or U13581 (N_13581,N_13382,N_13462);
nand U13582 (N_13582,N_13472,N_13409);
or U13583 (N_13583,N_13432,N_13449);
nor U13584 (N_13584,N_13476,N_13377);
xnor U13585 (N_13585,N_13410,N_13376);
and U13586 (N_13586,N_13460,N_13445);
or U13587 (N_13587,N_13493,N_13484);
xor U13588 (N_13588,N_13496,N_13439);
nand U13589 (N_13589,N_13411,N_13465);
and U13590 (N_13590,N_13490,N_13473);
nor U13591 (N_13591,N_13480,N_13462);
nor U13592 (N_13592,N_13394,N_13436);
or U13593 (N_13593,N_13478,N_13391);
xnor U13594 (N_13594,N_13391,N_13474);
nand U13595 (N_13595,N_13386,N_13415);
nand U13596 (N_13596,N_13442,N_13490);
xor U13597 (N_13597,N_13498,N_13394);
nor U13598 (N_13598,N_13410,N_13483);
nand U13599 (N_13599,N_13433,N_13497);
xnor U13600 (N_13600,N_13419,N_13467);
or U13601 (N_13601,N_13394,N_13396);
xor U13602 (N_13602,N_13385,N_13433);
nand U13603 (N_13603,N_13408,N_13401);
nand U13604 (N_13604,N_13406,N_13401);
nor U13605 (N_13605,N_13399,N_13475);
xnor U13606 (N_13606,N_13397,N_13377);
nor U13607 (N_13607,N_13401,N_13394);
nand U13608 (N_13608,N_13398,N_13441);
and U13609 (N_13609,N_13470,N_13496);
xor U13610 (N_13610,N_13432,N_13476);
xor U13611 (N_13611,N_13462,N_13498);
nand U13612 (N_13612,N_13484,N_13421);
nand U13613 (N_13613,N_13459,N_13406);
or U13614 (N_13614,N_13481,N_13378);
xor U13615 (N_13615,N_13378,N_13449);
xor U13616 (N_13616,N_13454,N_13445);
nand U13617 (N_13617,N_13407,N_13478);
nor U13618 (N_13618,N_13378,N_13493);
nor U13619 (N_13619,N_13459,N_13464);
or U13620 (N_13620,N_13484,N_13425);
or U13621 (N_13621,N_13381,N_13397);
and U13622 (N_13622,N_13456,N_13462);
nor U13623 (N_13623,N_13409,N_13428);
nor U13624 (N_13624,N_13486,N_13438);
nand U13625 (N_13625,N_13552,N_13570);
nand U13626 (N_13626,N_13535,N_13521);
xnor U13627 (N_13627,N_13567,N_13520);
xnor U13628 (N_13628,N_13507,N_13550);
nand U13629 (N_13629,N_13577,N_13545);
xnor U13630 (N_13630,N_13572,N_13519);
nand U13631 (N_13631,N_13529,N_13538);
nand U13632 (N_13632,N_13605,N_13503);
or U13633 (N_13633,N_13506,N_13618);
and U13634 (N_13634,N_13585,N_13561);
and U13635 (N_13635,N_13500,N_13597);
nor U13636 (N_13636,N_13525,N_13591);
xnor U13637 (N_13637,N_13514,N_13607);
or U13638 (N_13638,N_13536,N_13556);
or U13639 (N_13639,N_13562,N_13539);
or U13640 (N_13640,N_13617,N_13576);
xnor U13641 (N_13641,N_13606,N_13516);
nand U13642 (N_13642,N_13615,N_13543);
nand U13643 (N_13643,N_13616,N_13553);
nor U13644 (N_13644,N_13600,N_13610);
nand U13645 (N_13645,N_13557,N_13505);
and U13646 (N_13646,N_13544,N_13622);
nor U13647 (N_13647,N_13586,N_13568);
or U13648 (N_13648,N_13579,N_13564);
nor U13649 (N_13649,N_13604,N_13512);
nand U13650 (N_13650,N_13554,N_13620);
nor U13651 (N_13651,N_13595,N_13571);
nor U13652 (N_13652,N_13548,N_13517);
nand U13653 (N_13653,N_13527,N_13608);
nor U13654 (N_13654,N_13588,N_13612);
or U13655 (N_13655,N_13541,N_13504);
xnor U13656 (N_13656,N_13526,N_13611);
nand U13657 (N_13657,N_13533,N_13589);
nor U13658 (N_13658,N_13566,N_13621);
and U13659 (N_13659,N_13614,N_13601);
nand U13660 (N_13660,N_13540,N_13534);
and U13661 (N_13661,N_13569,N_13609);
nor U13662 (N_13662,N_13558,N_13596);
or U13663 (N_13663,N_13623,N_13590);
nor U13664 (N_13664,N_13593,N_13624);
nand U13665 (N_13665,N_13559,N_13581);
nand U13666 (N_13666,N_13549,N_13546);
nand U13667 (N_13667,N_13532,N_13575);
xnor U13668 (N_13668,N_13582,N_13508);
and U13669 (N_13669,N_13518,N_13599);
nand U13670 (N_13670,N_13528,N_13594);
or U13671 (N_13671,N_13513,N_13547);
or U13672 (N_13672,N_13537,N_13511);
nor U13673 (N_13673,N_13578,N_13515);
or U13674 (N_13674,N_13565,N_13530);
and U13675 (N_13675,N_13501,N_13510);
nor U13676 (N_13676,N_13584,N_13613);
nand U13677 (N_13677,N_13560,N_13573);
and U13678 (N_13678,N_13542,N_13522);
or U13679 (N_13679,N_13583,N_13523);
nor U13680 (N_13680,N_13502,N_13574);
or U13681 (N_13681,N_13551,N_13555);
and U13682 (N_13682,N_13602,N_13509);
nor U13683 (N_13683,N_13580,N_13592);
nor U13684 (N_13684,N_13531,N_13563);
or U13685 (N_13685,N_13524,N_13587);
xnor U13686 (N_13686,N_13598,N_13603);
nor U13687 (N_13687,N_13619,N_13559);
nand U13688 (N_13688,N_13520,N_13571);
and U13689 (N_13689,N_13581,N_13584);
or U13690 (N_13690,N_13521,N_13530);
or U13691 (N_13691,N_13613,N_13551);
and U13692 (N_13692,N_13612,N_13571);
and U13693 (N_13693,N_13621,N_13517);
nand U13694 (N_13694,N_13614,N_13510);
xnor U13695 (N_13695,N_13611,N_13523);
and U13696 (N_13696,N_13587,N_13577);
xor U13697 (N_13697,N_13580,N_13583);
nand U13698 (N_13698,N_13523,N_13554);
nor U13699 (N_13699,N_13523,N_13559);
xor U13700 (N_13700,N_13539,N_13607);
xnor U13701 (N_13701,N_13582,N_13545);
nor U13702 (N_13702,N_13524,N_13609);
xnor U13703 (N_13703,N_13614,N_13607);
and U13704 (N_13704,N_13579,N_13508);
and U13705 (N_13705,N_13539,N_13538);
nand U13706 (N_13706,N_13580,N_13567);
xor U13707 (N_13707,N_13523,N_13517);
xnor U13708 (N_13708,N_13587,N_13541);
and U13709 (N_13709,N_13609,N_13545);
or U13710 (N_13710,N_13604,N_13596);
xnor U13711 (N_13711,N_13554,N_13540);
nand U13712 (N_13712,N_13559,N_13538);
nor U13713 (N_13713,N_13548,N_13612);
xnor U13714 (N_13714,N_13569,N_13542);
or U13715 (N_13715,N_13608,N_13528);
and U13716 (N_13716,N_13526,N_13589);
or U13717 (N_13717,N_13527,N_13530);
nor U13718 (N_13718,N_13616,N_13615);
nor U13719 (N_13719,N_13536,N_13573);
and U13720 (N_13720,N_13530,N_13526);
nand U13721 (N_13721,N_13547,N_13620);
or U13722 (N_13722,N_13558,N_13527);
nor U13723 (N_13723,N_13623,N_13531);
and U13724 (N_13724,N_13530,N_13598);
nor U13725 (N_13725,N_13505,N_13621);
nor U13726 (N_13726,N_13602,N_13532);
xor U13727 (N_13727,N_13617,N_13541);
and U13728 (N_13728,N_13594,N_13607);
and U13729 (N_13729,N_13551,N_13535);
nand U13730 (N_13730,N_13616,N_13582);
xor U13731 (N_13731,N_13586,N_13519);
xnor U13732 (N_13732,N_13619,N_13543);
and U13733 (N_13733,N_13603,N_13513);
and U13734 (N_13734,N_13622,N_13551);
xor U13735 (N_13735,N_13520,N_13531);
and U13736 (N_13736,N_13526,N_13538);
nand U13737 (N_13737,N_13555,N_13531);
and U13738 (N_13738,N_13522,N_13527);
and U13739 (N_13739,N_13617,N_13517);
nand U13740 (N_13740,N_13559,N_13605);
and U13741 (N_13741,N_13578,N_13554);
nand U13742 (N_13742,N_13557,N_13614);
and U13743 (N_13743,N_13601,N_13517);
nor U13744 (N_13744,N_13596,N_13560);
and U13745 (N_13745,N_13597,N_13620);
and U13746 (N_13746,N_13539,N_13524);
and U13747 (N_13747,N_13623,N_13540);
nand U13748 (N_13748,N_13517,N_13541);
nand U13749 (N_13749,N_13580,N_13570);
or U13750 (N_13750,N_13730,N_13693);
or U13751 (N_13751,N_13652,N_13627);
and U13752 (N_13752,N_13679,N_13633);
xor U13753 (N_13753,N_13715,N_13626);
and U13754 (N_13754,N_13635,N_13639);
or U13755 (N_13755,N_13732,N_13727);
nor U13756 (N_13756,N_13670,N_13697);
xor U13757 (N_13757,N_13643,N_13700);
or U13758 (N_13758,N_13745,N_13704);
and U13759 (N_13759,N_13660,N_13649);
nand U13760 (N_13760,N_13655,N_13699);
xnor U13761 (N_13761,N_13721,N_13664);
xnor U13762 (N_13762,N_13651,N_13739);
or U13763 (N_13763,N_13666,N_13650);
nand U13764 (N_13764,N_13701,N_13676);
nand U13765 (N_13765,N_13681,N_13736);
nand U13766 (N_13766,N_13682,N_13625);
and U13767 (N_13767,N_13710,N_13647);
xor U13768 (N_13768,N_13658,N_13740);
xor U13769 (N_13769,N_13719,N_13632);
nand U13770 (N_13770,N_13687,N_13672);
and U13771 (N_13771,N_13690,N_13694);
and U13772 (N_13772,N_13638,N_13634);
or U13773 (N_13773,N_13703,N_13656);
nand U13774 (N_13774,N_13686,N_13702);
or U13775 (N_13775,N_13706,N_13734);
nand U13776 (N_13776,N_13661,N_13744);
nor U13777 (N_13777,N_13657,N_13677);
xor U13778 (N_13778,N_13628,N_13668);
xor U13779 (N_13779,N_13637,N_13631);
nor U13780 (N_13780,N_13748,N_13728);
or U13781 (N_13781,N_13691,N_13733);
or U13782 (N_13782,N_13688,N_13713);
nor U13783 (N_13783,N_13674,N_13685);
nor U13784 (N_13784,N_13737,N_13707);
nand U13785 (N_13785,N_13636,N_13720);
nor U13786 (N_13786,N_13729,N_13683);
xnor U13787 (N_13787,N_13642,N_13724);
and U13788 (N_13788,N_13726,N_13709);
nand U13789 (N_13789,N_13718,N_13696);
and U13790 (N_13790,N_13705,N_13711);
nor U13791 (N_13791,N_13747,N_13738);
xor U13792 (N_13792,N_13716,N_13742);
or U13793 (N_13793,N_13684,N_13722);
nor U13794 (N_13794,N_13654,N_13648);
and U13795 (N_13795,N_13714,N_13712);
nand U13796 (N_13796,N_13671,N_13725);
or U13797 (N_13797,N_13659,N_13630);
nor U13798 (N_13798,N_13741,N_13662);
nor U13799 (N_13799,N_13673,N_13669);
nand U13800 (N_13800,N_13667,N_13743);
nand U13801 (N_13801,N_13675,N_13695);
or U13802 (N_13802,N_13678,N_13641);
nor U13803 (N_13803,N_13723,N_13640);
or U13804 (N_13804,N_13717,N_13653);
nor U13805 (N_13805,N_13746,N_13735);
xnor U13806 (N_13806,N_13645,N_13629);
or U13807 (N_13807,N_13689,N_13708);
nor U13808 (N_13808,N_13680,N_13749);
nand U13809 (N_13809,N_13692,N_13698);
and U13810 (N_13810,N_13665,N_13644);
nand U13811 (N_13811,N_13731,N_13663);
and U13812 (N_13812,N_13646,N_13704);
nand U13813 (N_13813,N_13670,N_13647);
nand U13814 (N_13814,N_13719,N_13700);
or U13815 (N_13815,N_13671,N_13723);
or U13816 (N_13816,N_13720,N_13661);
or U13817 (N_13817,N_13747,N_13748);
and U13818 (N_13818,N_13726,N_13637);
xnor U13819 (N_13819,N_13736,N_13713);
and U13820 (N_13820,N_13708,N_13736);
or U13821 (N_13821,N_13736,N_13702);
nand U13822 (N_13822,N_13707,N_13722);
and U13823 (N_13823,N_13672,N_13628);
or U13824 (N_13824,N_13640,N_13681);
nand U13825 (N_13825,N_13722,N_13709);
and U13826 (N_13826,N_13726,N_13725);
xnor U13827 (N_13827,N_13697,N_13669);
xor U13828 (N_13828,N_13729,N_13742);
xnor U13829 (N_13829,N_13728,N_13641);
and U13830 (N_13830,N_13690,N_13674);
nand U13831 (N_13831,N_13683,N_13703);
nand U13832 (N_13832,N_13712,N_13696);
or U13833 (N_13833,N_13674,N_13732);
and U13834 (N_13834,N_13655,N_13716);
or U13835 (N_13835,N_13738,N_13652);
or U13836 (N_13836,N_13656,N_13653);
xnor U13837 (N_13837,N_13708,N_13726);
xor U13838 (N_13838,N_13668,N_13656);
xor U13839 (N_13839,N_13695,N_13676);
nor U13840 (N_13840,N_13625,N_13657);
and U13841 (N_13841,N_13712,N_13632);
and U13842 (N_13842,N_13734,N_13657);
or U13843 (N_13843,N_13664,N_13633);
nand U13844 (N_13844,N_13685,N_13666);
and U13845 (N_13845,N_13738,N_13672);
or U13846 (N_13846,N_13688,N_13732);
or U13847 (N_13847,N_13714,N_13680);
xor U13848 (N_13848,N_13749,N_13682);
or U13849 (N_13849,N_13724,N_13625);
nand U13850 (N_13850,N_13737,N_13744);
nand U13851 (N_13851,N_13686,N_13649);
and U13852 (N_13852,N_13644,N_13697);
nor U13853 (N_13853,N_13706,N_13694);
or U13854 (N_13854,N_13644,N_13729);
and U13855 (N_13855,N_13663,N_13691);
nor U13856 (N_13856,N_13730,N_13745);
and U13857 (N_13857,N_13702,N_13630);
xor U13858 (N_13858,N_13723,N_13735);
xnor U13859 (N_13859,N_13666,N_13668);
nor U13860 (N_13860,N_13726,N_13719);
nor U13861 (N_13861,N_13675,N_13717);
nand U13862 (N_13862,N_13706,N_13714);
or U13863 (N_13863,N_13711,N_13684);
and U13864 (N_13864,N_13676,N_13725);
and U13865 (N_13865,N_13724,N_13635);
and U13866 (N_13866,N_13745,N_13715);
xnor U13867 (N_13867,N_13659,N_13664);
nor U13868 (N_13868,N_13713,N_13636);
and U13869 (N_13869,N_13745,N_13708);
and U13870 (N_13870,N_13658,N_13633);
xor U13871 (N_13871,N_13668,N_13646);
or U13872 (N_13872,N_13661,N_13672);
xor U13873 (N_13873,N_13682,N_13681);
xnor U13874 (N_13874,N_13692,N_13697);
xnor U13875 (N_13875,N_13849,N_13824);
and U13876 (N_13876,N_13766,N_13773);
and U13877 (N_13877,N_13769,N_13752);
xnor U13878 (N_13878,N_13858,N_13813);
and U13879 (N_13879,N_13810,N_13863);
nor U13880 (N_13880,N_13831,N_13833);
nor U13881 (N_13881,N_13862,N_13848);
nand U13882 (N_13882,N_13847,N_13856);
nand U13883 (N_13883,N_13854,N_13771);
or U13884 (N_13884,N_13796,N_13795);
nand U13885 (N_13885,N_13861,N_13853);
and U13886 (N_13886,N_13756,N_13793);
and U13887 (N_13887,N_13778,N_13834);
nor U13888 (N_13888,N_13774,N_13832);
nor U13889 (N_13889,N_13826,N_13782);
and U13890 (N_13890,N_13822,N_13841);
nor U13891 (N_13891,N_13823,N_13792);
nand U13892 (N_13892,N_13855,N_13837);
nand U13893 (N_13893,N_13815,N_13874);
xnor U13894 (N_13894,N_13768,N_13784);
nand U13895 (N_13895,N_13844,N_13839);
nand U13896 (N_13896,N_13787,N_13867);
or U13897 (N_13897,N_13765,N_13788);
or U13898 (N_13898,N_13779,N_13757);
nor U13899 (N_13899,N_13750,N_13772);
nor U13900 (N_13900,N_13835,N_13754);
or U13901 (N_13901,N_13764,N_13770);
nand U13902 (N_13902,N_13842,N_13827);
xor U13903 (N_13903,N_13808,N_13818);
xor U13904 (N_13904,N_13860,N_13789);
xor U13905 (N_13905,N_13819,N_13851);
or U13906 (N_13906,N_13828,N_13864);
or U13907 (N_13907,N_13843,N_13783);
nor U13908 (N_13908,N_13814,N_13868);
nor U13909 (N_13909,N_13776,N_13803);
and U13910 (N_13910,N_13845,N_13805);
nand U13911 (N_13911,N_13816,N_13873);
nand U13912 (N_13912,N_13790,N_13820);
and U13913 (N_13913,N_13817,N_13786);
xor U13914 (N_13914,N_13807,N_13785);
nor U13915 (N_13915,N_13809,N_13852);
nor U13916 (N_13916,N_13800,N_13799);
nor U13917 (N_13917,N_13872,N_13798);
and U13918 (N_13918,N_13821,N_13838);
or U13919 (N_13919,N_13806,N_13836);
nor U13920 (N_13920,N_13850,N_13781);
nand U13921 (N_13921,N_13794,N_13767);
or U13922 (N_13922,N_13780,N_13811);
nor U13923 (N_13923,N_13829,N_13804);
and U13924 (N_13924,N_13762,N_13865);
xor U13925 (N_13925,N_13751,N_13871);
and U13926 (N_13926,N_13758,N_13846);
or U13927 (N_13927,N_13801,N_13759);
or U13928 (N_13928,N_13763,N_13775);
nor U13929 (N_13929,N_13791,N_13812);
nor U13930 (N_13930,N_13870,N_13830);
xor U13931 (N_13931,N_13859,N_13869);
nand U13932 (N_13932,N_13797,N_13755);
or U13933 (N_13933,N_13825,N_13761);
and U13934 (N_13934,N_13753,N_13760);
nor U13935 (N_13935,N_13866,N_13840);
nor U13936 (N_13936,N_13777,N_13857);
and U13937 (N_13937,N_13802,N_13772);
nor U13938 (N_13938,N_13771,N_13768);
nor U13939 (N_13939,N_13796,N_13820);
or U13940 (N_13940,N_13869,N_13753);
and U13941 (N_13941,N_13838,N_13825);
xor U13942 (N_13942,N_13777,N_13855);
xnor U13943 (N_13943,N_13834,N_13770);
and U13944 (N_13944,N_13835,N_13751);
or U13945 (N_13945,N_13826,N_13830);
nor U13946 (N_13946,N_13822,N_13759);
and U13947 (N_13947,N_13816,N_13784);
nor U13948 (N_13948,N_13825,N_13750);
xor U13949 (N_13949,N_13826,N_13838);
nor U13950 (N_13950,N_13759,N_13784);
nor U13951 (N_13951,N_13797,N_13766);
nor U13952 (N_13952,N_13751,N_13787);
nand U13953 (N_13953,N_13873,N_13874);
and U13954 (N_13954,N_13868,N_13792);
xnor U13955 (N_13955,N_13784,N_13793);
or U13956 (N_13956,N_13757,N_13805);
nor U13957 (N_13957,N_13819,N_13830);
nand U13958 (N_13958,N_13780,N_13752);
nor U13959 (N_13959,N_13836,N_13788);
and U13960 (N_13960,N_13856,N_13828);
or U13961 (N_13961,N_13759,N_13854);
and U13962 (N_13962,N_13805,N_13855);
or U13963 (N_13963,N_13801,N_13812);
nor U13964 (N_13964,N_13870,N_13834);
and U13965 (N_13965,N_13808,N_13824);
xnor U13966 (N_13966,N_13808,N_13848);
and U13967 (N_13967,N_13845,N_13829);
and U13968 (N_13968,N_13796,N_13834);
or U13969 (N_13969,N_13774,N_13797);
nand U13970 (N_13970,N_13856,N_13782);
xor U13971 (N_13971,N_13793,N_13805);
and U13972 (N_13972,N_13844,N_13825);
and U13973 (N_13973,N_13854,N_13845);
nor U13974 (N_13974,N_13800,N_13757);
nand U13975 (N_13975,N_13804,N_13756);
and U13976 (N_13976,N_13769,N_13773);
and U13977 (N_13977,N_13837,N_13753);
or U13978 (N_13978,N_13802,N_13807);
and U13979 (N_13979,N_13767,N_13857);
nand U13980 (N_13980,N_13818,N_13851);
xor U13981 (N_13981,N_13810,N_13847);
or U13982 (N_13982,N_13836,N_13866);
nand U13983 (N_13983,N_13780,N_13845);
nor U13984 (N_13984,N_13863,N_13753);
nand U13985 (N_13985,N_13873,N_13836);
or U13986 (N_13986,N_13761,N_13754);
nor U13987 (N_13987,N_13811,N_13854);
xor U13988 (N_13988,N_13813,N_13854);
or U13989 (N_13989,N_13760,N_13870);
nor U13990 (N_13990,N_13789,N_13843);
nor U13991 (N_13991,N_13790,N_13792);
or U13992 (N_13992,N_13755,N_13764);
xor U13993 (N_13993,N_13868,N_13870);
xnor U13994 (N_13994,N_13765,N_13779);
nor U13995 (N_13995,N_13764,N_13825);
and U13996 (N_13996,N_13852,N_13756);
nand U13997 (N_13997,N_13835,N_13810);
nand U13998 (N_13998,N_13869,N_13870);
and U13999 (N_13999,N_13790,N_13768);
and U14000 (N_14000,N_13900,N_13907);
nand U14001 (N_14001,N_13993,N_13881);
xor U14002 (N_14002,N_13968,N_13920);
and U14003 (N_14003,N_13953,N_13942);
and U14004 (N_14004,N_13912,N_13891);
xnor U14005 (N_14005,N_13987,N_13928);
xnor U14006 (N_14006,N_13897,N_13981);
or U14007 (N_14007,N_13940,N_13916);
or U14008 (N_14008,N_13882,N_13931);
or U14009 (N_14009,N_13941,N_13967);
xnor U14010 (N_14010,N_13996,N_13909);
nand U14011 (N_14011,N_13974,N_13925);
or U14012 (N_14012,N_13998,N_13951);
and U14013 (N_14013,N_13956,N_13877);
or U14014 (N_14014,N_13893,N_13876);
or U14015 (N_14015,N_13963,N_13976);
and U14016 (N_14016,N_13904,N_13908);
xnor U14017 (N_14017,N_13914,N_13934);
xor U14018 (N_14018,N_13984,N_13949);
nor U14019 (N_14019,N_13911,N_13936);
xor U14020 (N_14020,N_13926,N_13921);
nor U14021 (N_14021,N_13983,N_13997);
xor U14022 (N_14022,N_13950,N_13885);
xnor U14023 (N_14023,N_13994,N_13886);
xnor U14024 (N_14024,N_13895,N_13905);
xor U14025 (N_14025,N_13927,N_13948);
xnor U14026 (N_14026,N_13959,N_13875);
or U14027 (N_14027,N_13910,N_13992);
and U14028 (N_14028,N_13999,N_13892);
and U14029 (N_14029,N_13924,N_13903);
xnor U14030 (N_14030,N_13947,N_13991);
and U14031 (N_14031,N_13988,N_13957);
xnor U14032 (N_14032,N_13961,N_13937);
nor U14033 (N_14033,N_13955,N_13896);
nand U14034 (N_14034,N_13888,N_13995);
nand U14035 (N_14035,N_13917,N_13899);
nand U14036 (N_14036,N_13954,N_13977);
xor U14037 (N_14037,N_13939,N_13966);
nand U14038 (N_14038,N_13915,N_13943);
nor U14039 (N_14039,N_13980,N_13880);
nor U14040 (N_14040,N_13944,N_13978);
or U14041 (N_14041,N_13973,N_13965);
xnor U14042 (N_14042,N_13913,N_13883);
or U14043 (N_14043,N_13986,N_13889);
nand U14044 (N_14044,N_13918,N_13929);
nor U14045 (N_14045,N_13922,N_13898);
or U14046 (N_14046,N_13960,N_13945);
xnor U14047 (N_14047,N_13878,N_13989);
xnor U14048 (N_14048,N_13982,N_13969);
nor U14049 (N_14049,N_13902,N_13938);
xnor U14050 (N_14050,N_13985,N_13958);
or U14051 (N_14051,N_13906,N_13964);
nor U14052 (N_14052,N_13971,N_13990);
nor U14053 (N_14053,N_13933,N_13884);
xnor U14054 (N_14054,N_13970,N_13975);
nor U14055 (N_14055,N_13932,N_13919);
and U14056 (N_14056,N_13901,N_13894);
nand U14057 (N_14057,N_13979,N_13930);
xor U14058 (N_14058,N_13952,N_13946);
and U14059 (N_14059,N_13972,N_13890);
nor U14060 (N_14060,N_13923,N_13879);
xor U14061 (N_14061,N_13887,N_13935);
or U14062 (N_14062,N_13962,N_13905);
and U14063 (N_14063,N_13989,N_13992);
nor U14064 (N_14064,N_13970,N_13938);
nor U14065 (N_14065,N_13997,N_13981);
xor U14066 (N_14066,N_13904,N_13877);
nor U14067 (N_14067,N_13988,N_13880);
xnor U14068 (N_14068,N_13926,N_13924);
or U14069 (N_14069,N_13905,N_13922);
xor U14070 (N_14070,N_13991,N_13930);
nand U14071 (N_14071,N_13976,N_13962);
nor U14072 (N_14072,N_13983,N_13945);
and U14073 (N_14073,N_13993,N_13901);
nand U14074 (N_14074,N_13966,N_13880);
xor U14075 (N_14075,N_13962,N_13920);
or U14076 (N_14076,N_13981,N_13951);
nor U14077 (N_14077,N_13896,N_13952);
nor U14078 (N_14078,N_13879,N_13999);
or U14079 (N_14079,N_13925,N_13932);
nor U14080 (N_14080,N_13986,N_13905);
xnor U14081 (N_14081,N_13966,N_13927);
or U14082 (N_14082,N_13906,N_13982);
xnor U14083 (N_14083,N_13936,N_13976);
xor U14084 (N_14084,N_13927,N_13925);
xnor U14085 (N_14085,N_13885,N_13982);
or U14086 (N_14086,N_13983,N_13887);
nor U14087 (N_14087,N_13897,N_13949);
nand U14088 (N_14088,N_13971,N_13895);
nor U14089 (N_14089,N_13968,N_13902);
nand U14090 (N_14090,N_13967,N_13899);
or U14091 (N_14091,N_13943,N_13995);
nor U14092 (N_14092,N_13901,N_13966);
and U14093 (N_14093,N_13890,N_13981);
xnor U14094 (N_14094,N_13882,N_13934);
nand U14095 (N_14095,N_13936,N_13983);
nand U14096 (N_14096,N_13994,N_13916);
nand U14097 (N_14097,N_13969,N_13962);
and U14098 (N_14098,N_13986,N_13891);
xor U14099 (N_14099,N_13985,N_13916);
xnor U14100 (N_14100,N_13933,N_13953);
nor U14101 (N_14101,N_13975,N_13914);
or U14102 (N_14102,N_13986,N_13919);
nand U14103 (N_14103,N_13908,N_13921);
and U14104 (N_14104,N_13886,N_13987);
or U14105 (N_14105,N_13895,N_13899);
nand U14106 (N_14106,N_13908,N_13945);
and U14107 (N_14107,N_13999,N_13958);
nor U14108 (N_14108,N_13938,N_13944);
nor U14109 (N_14109,N_13941,N_13920);
and U14110 (N_14110,N_13885,N_13918);
nor U14111 (N_14111,N_13889,N_13979);
nor U14112 (N_14112,N_13878,N_13978);
or U14113 (N_14113,N_13908,N_13910);
or U14114 (N_14114,N_13877,N_13924);
xnor U14115 (N_14115,N_13995,N_13987);
nand U14116 (N_14116,N_13938,N_13977);
or U14117 (N_14117,N_13915,N_13892);
nand U14118 (N_14118,N_13961,N_13948);
xor U14119 (N_14119,N_13981,N_13977);
xor U14120 (N_14120,N_13943,N_13990);
or U14121 (N_14121,N_13899,N_13945);
and U14122 (N_14122,N_13915,N_13991);
or U14123 (N_14123,N_13897,N_13890);
nor U14124 (N_14124,N_13891,N_13975);
and U14125 (N_14125,N_14062,N_14067);
and U14126 (N_14126,N_14104,N_14059);
or U14127 (N_14127,N_14048,N_14095);
nor U14128 (N_14128,N_14113,N_14093);
nor U14129 (N_14129,N_14014,N_14052);
nor U14130 (N_14130,N_14084,N_14118);
nor U14131 (N_14131,N_14009,N_14072);
or U14132 (N_14132,N_14082,N_14066);
or U14133 (N_14133,N_14026,N_14080);
nor U14134 (N_14134,N_14016,N_14089);
xor U14135 (N_14135,N_14045,N_14123);
nand U14136 (N_14136,N_14030,N_14090);
and U14137 (N_14137,N_14117,N_14038);
nand U14138 (N_14138,N_14021,N_14019);
xnor U14139 (N_14139,N_14079,N_14006);
nand U14140 (N_14140,N_14124,N_14029);
nor U14141 (N_14141,N_14047,N_14083);
nand U14142 (N_14142,N_14071,N_14017);
xnor U14143 (N_14143,N_14037,N_14022);
or U14144 (N_14144,N_14041,N_14060);
xnor U14145 (N_14145,N_14069,N_14043);
nor U14146 (N_14146,N_14114,N_14042);
and U14147 (N_14147,N_14112,N_14070);
xnor U14148 (N_14148,N_14056,N_14098);
xor U14149 (N_14149,N_14119,N_14106);
nand U14150 (N_14150,N_14064,N_14122);
and U14151 (N_14151,N_14103,N_14002);
and U14152 (N_14152,N_14065,N_14110);
nand U14153 (N_14153,N_14087,N_14091);
xor U14154 (N_14154,N_14057,N_14108);
or U14155 (N_14155,N_14003,N_14024);
xnor U14156 (N_14156,N_14076,N_14063);
or U14157 (N_14157,N_14078,N_14010);
nor U14158 (N_14158,N_14001,N_14092);
and U14159 (N_14159,N_14025,N_14011);
nand U14160 (N_14160,N_14007,N_14055);
or U14161 (N_14161,N_14008,N_14058);
nor U14162 (N_14162,N_14032,N_14121);
xor U14163 (N_14163,N_14049,N_14040);
and U14164 (N_14164,N_14068,N_14023);
or U14165 (N_14165,N_14053,N_14099);
nor U14166 (N_14166,N_14086,N_14111);
or U14167 (N_14167,N_14102,N_14012);
nor U14168 (N_14168,N_14105,N_14088);
nor U14169 (N_14169,N_14039,N_14081);
nand U14170 (N_14170,N_14034,N_14073);
and U14171 (N_14171,N_14074,N_14018);
nand U14172 (N_14172,N_14120,N_14035);
or U14173 (N_14173,N_14054,N_14020);
nor U14174 (N_14174,N_14031,N_14050);
nor U14175 (N_14175,N_14101,N_14000);
nor U14176 (N_14176,N_14094,N_14015);
or U14177 (N_14177,N_14107,N_14046);
nor U14178 (N_14178,N_14004,N_14077);
xor U14179 (N_14179,N_14100,N_14051);
nor U14180 (N_14180,N_14027,N_14085);
nor U14181 (N_14181,N_14096,N_14097);
nor U14182 (N_14182,N_14036,N_14061);
nand U14183 (N_14183,N_14115,N_14028);
or U14184 (N_14184,N_14044,N_14109);
or U14185 (N_14185,N_14075,N_14033);
xnor U14186 (N_14186,N_14116,N_14013);
xor U14187 (N_14187,N_14005,N_14011);
or U14188 (N_14188,N_14062,N_14009);
nand U14189 (N_14189,N_14043,N_14121);
nor U14190 (N_14190,N_14058,N_14118);
and U14191 (N_14191,N_14059,N_14007);
and U14192 (N_14192,N_14037,N_14049);
and U14193 (N_14193,N_14108,N_14060);
nor U14194 (N_14194,N_14016,N_14096);
or U14195 (N_14195,N_14072,N_14086);
or U14196 (N_14196,N_14005,N_14007);
or U14197 (N_14197,N_14030,N_14010);
or U14198 (N_14198,N_14088,N_14072);
or U14199 (N_14199,N_14019,N_14032);
nor U14200 (N_14200,N_14071,N_14023);
nand U14201 (N_14201,N_14051,N_14086);
xor U14202 (N_14202,N_14115,N_14058);
and U14203 (N_14203,N_14012,N_14057);
nor U14204 (N_14204,N_14029,N_14002);
or U14205 (N_14205,N_14015,N_14018);
or U14206 (N_14206,N_14083,N_14068);
nand U14207 (N_14207,N_14078,N_14120);
nor U14208 (N_14208,N_14124,N_14122);
nor U14209 (N_14209,N_14014,N_14035);
nand U14210 (N_14210,N_14051,N_14091);
nor U14211 (N_14211,N_14110,N_14039);
and U14212 (N_14212,N_14102,N_14056);
xor U14213 (N_14213,N_14106,N_14113);
and U14214 (N_14214,N_14066,N_14059);
and U14215 (N_14215,N_14091,N_14011);
xnor U14216 (N_14216,N_14038,N_14082);
nand U14217 (N_14217,N_14116,N_14006);
xor U14218 (N_14218,N_14070,N_14015);
or U14219 (N_14219,N_14083,N_14098);
and U14220 (N_14220,N_14034,N_14032);
xnor U14221 (N_14221,N_14086,N_14018);
and U14222 (N_14222,N_14070,N_14087);
nor U14223 (N_14223,N_14006,N_14044);
nand U14224 (N_14224,N_14119,N_14101);
or U14225 (N_14225,N_14033,N_14022);
nor U14226 (N_14226,N_14020,N_14042);
nor U14227 (N_14227,N_14113,N_14011);
or U14228 (N_14228,N_14081,N_14018);
and U14229 (N_14229,N_14006,N_14029);
or U14230 (N_14230,N_14075,N_14069);
and U14231 (N_14231,N_14049,N_14030);
xor U14232 (N_14232,N_14071,N_14033);
and U14233 (N_14233,N_14078,N_14086);
xnor U14234 (N_14234,N_14115,N_14060);
nand U14235 (N_14235,N_14019,N_14006);
xnor U14236 (N_14236,N_14020,N_14077);
and U14237 (N_14237,N_14048,N_14015);
and U14238 (N_14238,N_14078,N_14053);
and U14239 (N_14239,N_14003,N_14053);
nor U14240 (N_14240,N_14027,N_14010);
or U14241 (N_14241,N_14109,N_14026);
xor U14242 (N_14242,N_14005,N_14117);
and U14243 (N_14243,N_14039,N_14070);
nor U14244 (N_14244,N_14063,N_14016);
and U14245 (N_14245,N_14108,N_14015);
nand U14246 (N_14246,N_14116,N_14103);
or U14247 (N_14247,N_14036,N_14105);
and U14248 (N_14248,N_14069,N_14121);
nor U14249 (N_14249,N_14018,N_14052);
nor U14250 (N_14250,N_14224,N_14192);
xor U14251 (N_14251,N_14196,N_14207);
nor U14252 (N_14252,N_14145,N_14156);
and U14253 (N_14253,N_14144,N_14165);
or U14254 (N_14254,N_14172,N_14139);
xnor U14255 (N_14255,N_14230,N_14129);
nor U14256 (N_14256,N_14199,N_14211);
and U14257 (N_14257,N_14136,N_14248);
nand U14258 (N_14258,N_14197,N_14232);
and U14259 (N_14259,N_14215,N_14154);
nor U14260 (N_14260,N_14236,N_14168);
and U14261 (N_14261,N_14245,N_14220);
xnor U14262 (N_14262,N_14243,N_14208);
and U14263 (N_14263,N_14130,N_14181);
nand U14264 (N_14264,N_14221,N_14174);
nor U14265 (N_14265,N_14231,N_14244);
or U14266 (N_14266,N_14193,N_14188);
nand U14267 (N_14267,N_14135,N_14131);
xor U14268 (N_14268,N_14182,N_14153);
nor U14269 (N_14269,N_14246,N_14143);
nand U14270 (N_14270,N_14198,N_14206);
or U14271 (N_14271,N_14158,N_14157);
xor U14272 (N_14272,N_14177,N_14223);
nand U14273 (N_14273,N_14152,N_14146);
and U14274 (N_14274,N_14235,N_14164);
xnor U14275 (N_14275,N_14141,N_14125);
nor U14276 (N_14276,N_14155,N_14227);
nand U14277 (N_14277,N_14201,N_14163);
and U14278 (N_14278,N_14187,N_14234);
xnor U14279 (N_14279,N_14205,N_14180);
nand U14280 (N_14280,N_14218,N_14217);
nor U14281 (N_14281,N_14184,N_14173);
xnor U14282 (N_14282,N_14179,N_14228);
and U14283 (N_14283,N_14203,N_14190);
or U14284 (N_14284,N_14132,N_14225);
or U14285 (N_14285,N_14191,N_14166);
nor U14286 (N_14286,N_14189,N_14222);
and U14287 (N_14287,N_14212,N_14133);
nor U14288 (N_14288,N_14140,N_14186);
or U14289 (N_14289,N_14229,N_14167);
or U14290 (N_14290,N_14160,N_14176);
nand U14291 (N_14291,N_14151,N_14127);
and U14292 (N_14292,N_14238,N_14242);
nand U14293 (N_14293,N_14202,N_14204);
and U14294 (N_14294,N_14161,N_14134);
or U14295 (N_14295,N_14126,N_14169);
nand U14296 (N_14296,N_14148,N_14149);
nor U14297 (N_14297,N_14183,N_14178);
or U14298 (N_14298,N_14137,N_14209);
or U14299 (N_14299,N_14159,N_14233);
nor U14300 (N_14300,N_14237,N_14249);
xnor U14301 (N_14301,N_14194,N_14200);
xnor U14302 (N_14302,N_14239,N_14195);
xnor U14303 (N_14303,N_14142,N_14226);
nand U14304 (N_14304,N_14171,N_14175);
and U14305 (N_14305,N_14214,N_14170);
xnor U14306 (N_14306,N_14147,N_14247);
nand U14307 (N_14307,N_14241,N_14150);
and U14308 (N_14308,N_14162,N_14128);
nor U14309 (N_14309,N_14216,N_14210);
xor U14310 (N_14310,N_14213,N_14219);
or U14311 (N_14311,N_14185,N_14240);
xnor U14312 (N_14312,N_14138,N_14220);
xor U14313 (N_14313,N_14164,N_14129);
xor U14314 (N_14314,N_14217,N_14140);
nand U14315 (N_14315,N_14145,N_14163);
nor U14316 (N_14316,N_14155,N_14189);
nand U14317 (N_14317,N_14184,N_14240);
nor U14318 (N_14318,N_14203,N_14135);
and U14319 (N_14319,N_14152,N_14187);
or U14320 (N_14320,N_14158,N_14221);
and U14321 (N_14321,N_14201,N_14166);
or U14322 (N_14322,N_14228,N_14181);
xnor U14323 (N_14323,N_14199,N_14172);
nor U14324 (N_14324,N_14224,N_14126);
nand U14325 (N_14325,N_14147,N_14138);
nor U14326 (N_14326,N_14229,N_14239);
nor U14327 (N_14327,N_14191,N_14138);
xnor U14328 (N_14328,N_14176,N_14132);
nor U14329 (N_14329,N_14209,N_14184);
nor U14330 (N_14330,N_14229,N_14180);
and U14331 (N_14331,N_14205,N_14140);
nor U14332 (N_14332,N_14190,N_14145);
or U14333 (N_14333,N_14187,N_14146);
xor U14334 (N_14334,N_14229,N_14179);
nand U14335 (N_14335,N_14227,N_14191);
nor U14336 (N_14336,N_14130,N_14172);
and U14337 (N_14337,N_14236,N_14181);
xnor U14338 (N_14338,N_14233,N_14132);
and U14339 (N_14339,N_14234,N_14134);
or U14340 (N_14340,N_14199,N_14194);
xnor U14341 (N_14341,N_14219,N_14244);
or U14342 (N_14342,N_14149,N_14163);
and U14343 (N_14343,N_14236,N_14206);
nand U14344 (N_14344,N_14137,N_14215);
nor U14345 (N_14345,N_14240,N_14201);
or U14346 (N_14346,N_14139,N_14189);
or U14347 (N_14347,N_14176,N_14192);
and U14348 (N_14348,N_14198,N_14211);
xnor U14349 (N_14349,N_14146,N_14198);
xnor U14350 (N_14350,N_14193,N_14161);
xor U14351 (N_14351,N_14218,N_14170);
xnor U14352 (N_14352,N_14220,N_14190);
xnor U14353 (N_14353,N_14158,N_14217);
nor U14354 (N_14354,N_14164,N_14169);
nor U14355 (N_14355,N_14243,N_14157);
nor U14356 (N_14356,N_14141,N_14191);
nand U14357 (N_14357,N_14165,N_14192);
nand U14358 (N_14358,N_14232,N_14171);
nand U14359 (N_14359,N_14234,N_14173);
xnor U14360 (N_14360,N_14180,N_14164);
or U14361 (N_14361,N_14236,N_14200);
or U14362 (N_14362,N_14195,N_14126);
and U14363 (N_14363,N_14192,N_14126);
nand U14364 (N_14364,N_14173,N_14157);
or U14365 (N_14365,N_14175,N_14246);
nand U14366 (N_14366,N_14217,N_14227);
nor U14367 (N_14367,N_14137,N_14193);
nor U14368 (N_14368,N_14200,N_14247);
or U14369 (N_14369,N_14181,N_14240);
xnor U14370 (N_14370,N_14230,N_14126);
nor U14371 (N_14371,N_14214,N_14206);
nand U14372 (N_14372,N_14135,N_14234);
and U14373 (N_14373,N_14143,N_14226);
or U14374 (N_14374,N_14229,N_14145);
nand U14375 (N_14375,N_14259,N_14317);
nor U14376 (N_14376,N_14371,N_14274);
and U14377 (N_14377,N_14284,N_14257);
and U14378 (N_14378,N_14270,N_14354);
or U14379 (N_14379,N_14286,N_14344);
or U14380 (N_14380,N_14287,N_14306);
and U14381 (N_14381,N_14256,N_14345);
nand U14382 (N_14382,N_14280,N_14313);
or U14383 (N_14383,N_14361,N_14319);
xor U14384 (N_14384,N_14326,N_14364);
xor U14385 (N_14385,N_14324,N_14298);
or U14386 (N_14386,N_14258,N_14297);
xor U14387 (N_14387,N_14304,N_14312);
or U14388 (N_14388,N_14362,N_14295);
nor U14389 (N_14389,N_14340,N_14268);
or U14390 (N_14390,N_14305,N_14363);
nor U14391 (N_14391,N_14315,N_14282);
xor U14392 (N_14392,N_14329,N_14325);
and U14393 (N_14393,N_14254,N_14262);
xnor U14394 (N_14394,N_14308,N_14311);
and U14395 (N_14395,N_14369,N_14367);
nor U14396 (N_14396,N_14307,N_14302);
xnor U14397 (N_14397,N_14271,N_14346);
and U14398 (N_14398,N_14294,N_14252);
nor U14399 (N_14399,N_14261,N_14360);
xnor U14400 (N_14400,N_14330,N_14342);
nand U14401 (N_14401,N_14293,N_14368);
xnor U14402 (N_14402,N_14323,N_14290);
or U14403 (N_14403,N_14366,N_14275);
xor U14404 (N_14404,N_14296,N_14322);
or U14405 (N_14405,N_14372,N_14343);
nor U14406 (N_14406,N_14338,N_14299);
xnor U14407 (N_14407,N_14337,N_14273);
nor U14408 (N_14408,N_14318,N_14320);
and U14409 (N_14409,N_14339,N_14267);
nor U14410 (N_14410,N_14351,N_14336);
xnor U14411 (N_14411,N_14250,N_14263);
nand U14412 (N_14412,N_14279,N_14285);
xor U14413 (N_14413,N_14352,N_14277);
and U14414 (N_14414,N_14292,N_14253);
xnor U14415 (N_14415,N_14355,N_14373);
and U14416 (N_14416,N_14269,N_14301);
or U14417 (N_14417,N_14365,N_14289);
xor U14418 (N_14418,N_14291,N_14347);
nand U14419 (N_14419,N_14356,N_14341);
nor U14420 (N_14420,N_14255,N_14260);
and U14421 (N_14421,N_14334,N_14374);
and U14422 (N_14422,N_14328,N_14309);
xnor U14423 (N_14423,N_14350,N_14370);
and U14424 (N_14424,N_14300,N_14358);
or U14425 (N_14425,N_14276,N_14265);
xor U14426 (N_14426,N_14335,N_14348);
or U14427 (N_14427,N_14332,N_14281);
nor U14428 (N_14428,N_14314,N_14321);
xnor U14429 (N_14429,N_14278,N_14272);
and U14430 (N_14430,N_14283,N_14251);
nand U14431 (N_14431,N_14349,N_14353);
or U14432 (N_14432,N_14288,N_14266);
xnor U14433 (N_14433,N_14331,N_14359);
or U14434 (N_14434,N_14327,N_14333);
or U14435 (N_14435,N_14303,N_14310);
nor U14436 (N_14436,N_14264,N_14357);
nor U14437 (N_14437,N_14316,N_14368);
nor U14438 (N_14438,N_14363,N_14258);
xnor U14439 (N_14439,N_14291,N_14312);
or U14440 (N_14440,N_14332,N_14259);
nor U14441 (N_14441,N_14274,N_14272);
or U14442 (N_14442,N_14352,N_14320);
nor U14443 (N_14443,N_14318,N_14372);
xor U14444 (N_14444,N_14343,N_14253);
and U14445 (N_14445,N_14302,N_14334);
nand U14446 (N_14446,N_14358,N_14311);
nand U14447 (N_14447,N_14325,N_14332);
nand U14448 (N_14448,N_14326,N_14371);
nor U14449 (N_14449,N_14309,N_14254);
nand U14450 (N_14450,N_14281,N_14315);
or U14451 (N_14451,N_14287,N_14263);
and U14452 (N_14452,N_14297,N_14269);
nor U14453 (N_14453,N_14296,N_14286);
nor U14454 (N_14454,N_14280,N_14291);
or U14455 (N_14455,N_14373,N_14287);
nor U14456 (N_14456,N_14356,N_14294);
xnor U14457 (N_14457,N_14296,N_14341);
xnor U14458 (N_14458,N_14349,N_14295);
nand U14459 (N_14459,N_14275,N_14258);
xor U14460 (N_14460,N_14262,N_14346);
and U14461 (N_14461,N_14362,N_14290);
nor U14462 (N_14462,N_14365,N_14264);
nand U14463 (N_14463,N_14256,N_14357);
and U14464 (N_14464,N_14290,N_14302);
or U14465 (N_14465,N_14359,N_14266);
or U14466 (N_14466,N_14316,N_14335);
nor U14467 (N_14467,N_14265,N_14262);
nor U14468 (N_14468,N_14365,N_14361);
or U14469 (N_14469,N_14316,N_14309);
nand U14470 (N_14470,N_14340,N_14262);
or U14471 (N_14471,N_14268,N_14362);
nor U14472 (N_14472,N_14365,N_14371);
or U14473 (N_14473,N_14259,N_14284);
nand U14474 (N_14474,N_14298,N_14314);
nand U14475 (N_14475,N_14283,N_14328);
or U14476 (N_14476,N_14368,N_14313);
nand U14477 (N_14477,N_14310,N_14302);
nor U14478 (N_14478,N_14304,N_14285);
nand U14479 (N_14479,N_14301,N_14263);
xnor U14480 (N_14480,N_14354,N_14294);
nand U14481 (N_14481,N_14331,N_14276);
or U14482 (N_14482,N_14255,N_14360);
nor U14483 (N_14483,N_14254,N_14327);
nand U14484 (N_14484,N_14323,N_14325);
nand U14485 (N_14485,N_14250,N_14319);
or U14486 (N_14486,N_14296,N_14302);
xor U14487 (N_14487,N_14280,N_14279);
nand U14488 (N_14488,N_14305,N_14357);
and U14489 (N_14489,N_14288,N_14323);
and U14490 (N_14490,N_14299,N_14281);
or U14491 (N_14491,N_14331,N_14291);
and U14492 (N_14492,N_14359,N_14334);
nor U14493 (N_14493,N_14369,N_14359);
xnor U14494 (N_14494,N_14336,N_14341);
xnor U14495 (N_14495,N_14266,N_14342);
or U14496 (N_14496,N_14296,N_14271);
and U14497 (N_14497,N_14323,N_14365);
nor U14498 (N_14498,N_14347,N_14299);
nand U14499 (N_14499,N_14342,N_14315);
or U14500 (N_14500,N_14471,N_14385);
nor U14501 (N_14501,N_14483,N_14408);
nand U14502 (N_14502,N_14447,N_14437);
or U14503 (N_14503,N_14469,N_14497);
xnor U14504 (N_14504,N_14394,N_14495);
nand U14505 (N_14505,N_14392,N_14444);
and U14506 (N_14506,N_14451,N_14388);
nand U14507 (N_14507,N_14404,N_14440);
nand U14508 (N_14508,N_14474,N_14414);
nand U14509 (N_14509,N_14435,N_14393);
or U14510 (N_14510,N_14411,N_14465);
or U14511 (N_14511,N_14425,N_14432);
and U14512 (N_14512,N_14413,N_14454);
nand U14513 (N_14513,N_14446,N_14496);
nand U14514 (N_14514,N_14375,N_14416);
nor U14515 (N_14515,N_14433,N_14493);
xnor U14516 (N_14516,N_14485,N_14412);
nor U14517 (N_14517,N_14439,N_14463);
xor U14518 (N_14518,N_14452,N_14475);
or U14519 (N_14519,N_14383,N_14409);
and U14520 (N_14520,N_14426,N_14498);
or U14521 (N_14521,N_14405,N_14396);
or U14522 (N_14522,N_14479,N_14420);
xor U14523 (N_14523,N_14407,N_14478);
nand U14524 (N_14524,N_14494,N_14389);
nor U14525 (N_14525,N_14418,N_14459);
nand U14526 (N_14526,N_14427,N_14380);
xor U14527 (N_14527,N_14424,N_14441);
nor U14528 (N_14528,N_14430,N_14415);
nand U14529 (N_14529,N_14448,N_14434);
nor U14530 (N_14530,N_14403,N_14467);
or U14531 (N_14531,N_14488,N_14491);
or U14532 (N_14532,N_14436,N_14395);
nand U14533 (N_14533,N_14431,N_14450);
nand U14534 (N_14534,N_14386,N_14398);
xor U14535 (N_14535,N_14401,N_14445);
nor U14536 (N_14536,N_14382,N_14406);
nand U14537 (N_14537,N_14473,N_14455);
nand U14538 (N_14538,N_14423,N_14468);
and U14539 (N_14539,N_14453,N_14422);
nand U14540 (N_14540,N_14486,N_14438);
xor U14541 (N_14541,N_14460,N_14482);
and U14542 (N_14542,N_14429,N_14417);
xnor U14543 (N_14543,N_14410,N_14489);
or U14544 (N_14544,N_14421,N_14378);
and U14545 (N_14545,N_14443,N_14499);
xnor U14546 (N_14546,N_14457,N_14477);
nand U14547 (N_14547,N_14428,N_14400);
and U14548 (N_14548,N_14481,N_14458);
xor U14549 (N_14549,N_14456,N_14464);
xnor U14550 (N_14550,N_14480,N_14419);
nor U14551 (N_14551,N_14442,N_14487);
xnor U14552 (N_14552,N_14390,N_14384);
nor U14553 (N_14553,N_14461,N_14376);
nand U14554 (N_14554,N_14391,N_14449);
nor U14555 (N_14555,N_14476,N_14472);
and U14556 (N_14556,N_14387,N_14470);
nor U14557 (N_14557,N_14399,N_14377);
or U14558 (N_14558,N_14379,N_14484);
or U14559 (N_14559,N_14492,N_14381);
or U14560 (N_14560,N_14397,N_14462);
nand U14561 (N_14561,N_14402,N_14490);
nor U14562 (N_14562,N_14466,N_14454);
xnor U14563 (N_14563,N_14478,N_14390);
nor U14564 (N_14564,N_14480,N_14477);
and U14565 (N_14565,N_14421,N_14430);
and U14566 (N_14566,N_14429,N_14385);
or U14567 (N_14567,N_14405,N_14472);
xor U14568 (N_14568,N_14423,N_14481);
or U14569 (N_14569,N_14487,N_14405);
nor U14570 (N_14570,N_14458,N_14455);
xor U14571 (N_14571,N_14487,N_14412);
and U14572 (N_14572,N_14495,N_14435);
xor U14573 (N_14573,N_14409,N_14451);
xnor U14574 (N_14574,N_14395,N_14450);
or U14575 (N_14575,N_14389,N_14393);
and U14576 (N_14576,N_14461,N_14405);
and U14577 (N_14577,N_14380,N_14493);
nor U14578 (N_14578,N_14410,N_14466);
nand U14579 (N_14579,N_14477,N_14441);
and U14580 (N_14580,N_14384,N_14490);
nand U14581 (N_14581,N_14418,N_14487);
xnor U14582 (N_14582,N_14402,N_14428);
and U14583 (N_14583,N_14464,N_14420);
nand U14584 (N_14584,N_14394,N_14387);
xnor U14585 (N_14585,N_14420,N_14487);
or U14586 (N_14586,N_14471,N_14493);
and U14587 (N_14587,N_14470,N_14393);
and U14588 (N_14588,N_14472,N_14430);
xor U14589 (N_14589,N_14466,N_14432);
xnor U14590 (N_14590,N_14454,N_14487);
or U14591 (N_14591,N_14433,N_14442);
nand U14592 (N_14592,N_14396,N_14448);
nand U14593 (N_14593,N_14389,N_14380);
xor U14594 (N_14594,N_14467,N_14461);
nor U14595 (N_14595,N_14458,N_14482);
nand U14596 (N_14596,N_14401,N_14413);
or U14597 (N_14597,N_14386,N_14459);
nor U14598 (N_14598,N_14483,N_14464);
or U14599 (N_14599,N_14481,N_14447);
nor U14600 (N_14600,N_14475,N_14444);
xnor U14601 (N_14601,N_14410,N_14440);
nand U14602 (N_14602,N_14460,N_14407);
and U14603 (N_14603,N_14487,N_14479);
nand U14604 (N_14604,N_14428,N_14491);
or U14605 (N_14605,N_14499,N_14472);
and U14606 (N_14606,N_14464,N_14463);
or U14607 (N_14607,N_14455,N_14424);
or U14608 (N_14608,N_14389,N_14410);
or U14609 (N_14609,N_14494,N_14447);
or U14610 (N_14610,N_14379,N_14495);
or U14611 (N_14611,N_14466,N_14405);
or U14612 (N_14612,N_14491,N_14492);
nand U14613 (N_14613,N_14482,N_14389);
nor U14614 (N_14614,N_14399,N_14419);
nor U14615 (N_14615,N_14473,N_14488);
xor U14616 (N_14616,N_14489,N_14418);
xor U14617 (N_14617,N_14429,N_14399);
or U14618 (N_14618,N_14445,N_14435);
nand U14619 (N_14619,N_14483,N_14395);
or U14620 (N_14620,N_14378,N_14486);
nor U14621 (N_14621,N_14403,N_14472);
and U14622 (N_14622,N_14377,N_14376);
nor U14623 (N_14623,N_14414,N_14461);
nor U14624 (N_14624,N_14472,N_14412);
or U14625 (N_14625,N_14615,N_14507);
or U14626 (N_14626,N_14504,N_14591);
nand U14627 (N_14627,N_14607,N_14575);
and U14628 (N_14628,N_14579,N_14604);
xor U14629 (N_14629,N_14537,N_14602);
nor U14630 (N_14630,N_14552,N_14563);
nand U14631 (N_14631,N_14609,N_14570);
xor U14632 (N_14632,N_14542,N_14582);
xnor U14633 (N_14633,N_14555,N_14515);
nand U14634 (N_14634,N_14562,N_14532);
xnor U14635 (N_14635,N_14508,N_14600);
xnor U14636 (N_14636,N_14501,N_14623);
and U14637 (N_14637,N_14611,N_14536);
and U14638 (N_14638,N_14605,N_14583);
or U14639 (N_14639,N_14543,N_14523);
xnor U14640 (N_14640,N_14593,N_14619);
and U14641 (N_14641,N_14585,N_14574);
nand U14642 (N_14642,N_14594,N_14546);
xor U14643 (N_14643,N_14502,N_14618);
nand U14644 (N_14644,N_14587,N_14512);
nand U14645 (N_14645,N_14530,N_14576);
and U14646 (N_14646,N_14520,N_14557);
xnor U14647 (N_14647,N_14534,N_14572);
nor U14648 (N_14648,N_14566,N_14533);
nor U14649 (N_14649,N_14526,N_14578);
xor U14650 (N_14650,N_14521,N_14539);
nor U14651 (N_14651,N_14588,N_14516);
and U14652 (N_14652,N_14549,N_14599);
and U14653 (N_14653,N_14511,N_14624);
xnor U14654 (N_14654,N_14571,N_14554);
or U14655 (N_14655,N_14596,N_14548);
nor U14656 (N_14656,N_14553,N_14517);
or U14657 (N_14657,N_14513,N_14561);
nand U14658 (N_14658,N_14538,N_14527);
nor U14659 (N_14659,N_14586,N_14590);
xnor U14660 (N_14660,N_14514,N_14608);
nor U14661 (N_14661,N_14518,N_14616);
xnor U14662 (N_14662,N_14510,N_14509);
xnor U14663 (N_14663,N_14597,N_14540);
or U14664 (N_14664,N_14617,N_14592);
nand U14665 (N_14665,N_14564,N_14584);
xor U14666 (N_14666,N_14541,N_14545);
nand U14667 (N_14667,N_14622,N_14528);
nor U14668 (N_14668,N_14620,N_14567);
nand U14669 (N_14669,N_14522,N_14558);
or U14670 (N_14670,N_14500,N_14519);
and U14671 (N_14671,N_14544,N_14503);
and U14672 (N_14672,N_14529,N_14589);
nand U14673 (N_14673,N_14505,N_14613);
nor U14674 (N_14674,N_14547,N_14550);
and U14675 (N_14675,N_14559,N_14565);
or U14676 (N_14676,N_14595,N_14612);
and U14677 (N_14677,N_14621,N_14525);
nand U14678 (N_14678,N_14551,N_14610);
and U14679 (N_14679,N_14531,N_14524);
xor U14680 (N_14680,N_14577,N_14601);
and U14681 (N_14681,N_14581,N_14580);
nand U14682 (N_14682,N_14606,N_14603);
or U14683 (N_14683,N_14598,N_14506);
and U14684 (N_14684,N_14556,N_14560);
and U14685 (N_14685,N_14573,N_14535);
nor U14686 (N_14686,N_14614,N_14569);
xor U14687 (N_14687,N_14568,N_14598);
nor U14688 (N_14688,N_14555,N_14580);
xnor U14689 (N_14689,N_14513,N_14515);
or U14690 (N_14690,N_14618,N_14610);
or U14691 (N_14691,N_14618,N_14536);
nor U14692 (N_14692,N_14620,N_14590);
or U14693 (N_14693,N_14550,N_14592);
or U14694 (N_14694,N_14518,N_14541);
nand U14695 (N_14695,N_14532,N_14558);
or U14696 (N_14696,N_14599,N_14577);
nand U14697 (N_14697,N_14612,N_14589);
nor U14698 (N_14698,N_14613,N_14610);
nor U14699 (N_14699,N_14599,N_14517);
xor U14700 (N_14700,N_14507,N_14572);
nor U14701 (N_14701,N_14540,N_14583);
nor U14702 (N_14702,N_14558,N_14572);
or U14703 (N_14703,N_14591,N_14530);
and U14704 (N_14704,N_14588,N_14579);
xnor U14705 (N_14705,N_14593,N_14613);
nand U14706 (N_14706,N_14525,N_14578);
or U14707 (N_14707,N_14532,N_14621);
and U14708 (N_14708,N_14546,N_14561);
xor U14709 (N_14709,N_14524,N_14544);
xnor U14710 (N_14710,N_14534,N_14620);
nor U14711 (N_14711,N_14510,N_14593);
xnor U14712 (N_14712,N_14563,N_14573);
nand U14713 (N_14713,N_14534,N_14542);
nand U14714 (N_14714,N_14581,N_14529);
xnor U14715 (N_14715,N_14619,N_14504);
nand U14716 (N_14716,N_14622,N_14547);
or U14717 (N_14717,N_14586,N_14518);
nor U14718 (N_14718,N_14598,N_14559);
nor U14719 (N_14719,N_14622,N_14503);
or U14720 (N_14720,N_14556,N_14574);
or U14721 (N_14721,N_14515,N_14600);
and U14722 (N_14722,N_14513,N_14581);
or U14723 (N_14723,N_14605,N_14586);
or U14724 (N_14724,N_14598,N_14610);
xnor U14725 (N_14725,N_14520,N_14539);
nand U14726 (N_14726,N_14502,N_14521);
xor U14727 (N_14727,N_14571,N_14592);
nand U14728 (N_14728,N_14591,N_14607);
xnor U14729 (N_14729,N_14591,N_14562);
xnor U14730 (N_14730,N_14573,N_14559);
nor U14731 (N_14731,N_14572,N_14599);
or U14732 (N_14732,N_14603,N_14586);
nand U14733 (N_14733,N_14608,N_14569);
nand U14734 (N_14734,N_14548,N_14623);
and U14735 (N_14735,N_14575,N_14525);
xnor U14736 (N_14736,N_14622,N_14510);
nor U14737 (N_14737,N_14576,N_14597);
and U14738 (N_14738,N_14612,N_14510);
nand U14739 (N_14739,N_14543,N_14569);
and U14740 (N_14740,N_14549,N_14575);
or U14741 (N_14741,N_14618,N_14608);
and U14742 (N_14742,N_14555,N_14501);
xor U14743 (N_14743,N_14606,N_14554);
nor U14744 (N_14744,N_14502,N_14605);
and U14745 (N_14745,N_14541,N_14613);
nand U14746 (N_14746,N_14531,N_14567);
nand U14747 (N_14747,N_14577,N_14511);
and U14748 (N_14748,N_14617,N_14571);
or U14749 (N_14749,N_14616,N_14531);
and U14750 (N_14750,N_14719,N_14743);
xor U14751 (N_14751,N_14715,N_14628);
or U14752 (N_14752,N_14643,N_14634);
and U14753 (N_14753,N_14669,N_14657);
nor U14754 (N_14754,N_14749,N_14641);
and U14755 (N_14755,N_14637,N_14650);
nor U14756 (N_14756,N_14716,N_14666);
nor U14757 (N_14757,N_14709,N_14706);
nand U14758 (N_14758,N_14701,N_14662);
nand U14759 (N_14759,N_14627,N_14654);
nand U14760 (N_14760,N_14705,N_14732);
nand U14761 (N_14761,N_14632,N_14676);
nor U14762 (N_14762,N_14635,N_14723);
nand U14763 (N_14763,N_14718,N_14711);
nand U14764 (N_14764,N_14714,N_14693);
nand U14765 (N_14765,N_14661,N_14724);
or U14766 (N_14766,N_14675,N_14713);
nand U14767 (N_14767,N_14748,N_14678);
and U14768 (N_14768,N_14665,N_14636);
and U14769 (N_14769,N_14647,N_14737);
and U14770 (N_14770,N_14689,N_14648);
nand U14771 (N_14771,N_14655,N_14646);
nand U14772 (N_14772,N_14679,N_14645);
nand U14773 (N_14773,N_14673,N_14736);
xnor U14774 (N_14774,N_14690,N_14687);
and U14775 (N_14775,N_14729,N_14702);
nor U14776 (N_14776,N_14660,N_14683);
nor U14777 (N_14777,N_14688,N_14722);
nor U14778 (N_14778,N_14725,N_14742);
and U14779 (N_14779,N_14664,N_14659);
nor U14780 (N_14780,N_14695,N_14727);
nor U14781 (N_14781,N_14745,N_14730);
nor U14782 (N_14782,N_14710,N_14656);
nand U14783 (N_14783,N_14703,N_14653);
xnor U14784 (N_14784,N_14717,N_14728);
nand U14785 (N_14785,N_14698,N_14696);
nor U14786 (N_14786,N_14704,N_14644);
nand U14787 (N_14787,N_14741,N_14658);
or U14788 (N_14788,N_14649,N_14746);
nand U14789 (N_14789,N_14733,N_14692);
nor U14790 (N_14790,N_14699,N_14630);
and U14791 (N_14791,N_14668,N_14720);
and U14792 (N_14792,N_14734,N_14744);
nor U14793 (N_14793,N_14726,N_14629);
xnor U14794 (N_14794,N_14651,N_14691);
nand U14795 (N_14795,N_14663,N_14721);
xnor U14796 (N_14796,N_14639,N_14672);
nor U14797 (N_14797,N_14707,N_14694);
nand U14798 (N_14798,N_14735,N_14747);
or U14799 (N_14799,N_14740,N_14671);
or U14800 (N_14800,N_14633,N_14674);
and U14801 (N_14801,N_14631,N_14652);
xor U14802 (N_14802,N_14712,N_14667);
nand U14803 (N_14803,N_14739,N_14685);
xnor U14804 (N_14804,N_14738,N_14682);
nand U14805 (N_14805,N_14642,N_14686);
and U14806 (N_14806,N_14684,N_14626);
and U14807 (N_14807,N_14670,N_14625);
nand U14808 (N_14808,N_14677,N_14700);
and U14809 (N_14809,N_14640,N_14638);
or U14810 (N_14810,N_14708,N_14681);
or U14811 (N_14811,N_14731,N_14697);
xnor U14812 (N_14812,N_14680,N_14677);
xnor U14813 (N_14813,N_14633,N_14644);
nor U14814 (N_14814,N_14712,N_14746);
xnor U14815 (N_14815,N_14692,N_14744);
and U14816 (N_14816,N_14677,N_14641);
nand U14817 (N_14817,N_14652,N_14729);
nor U14818 (N_14818,N_14659,N_14662);
xnor U14819 (N_14819,N_14642,N_14659);
or U14820 (N_14820,N_14655,N_14666);
nor U14821 (N_14821,N_14680,N_14726);
nand U14822 (N_14822,N_14736,N_14682);
nand U14823 (N_14823,N_14708,N_14633);
xnor U14824 (N_14824,N_14726,N_14651);
xnor U14825 (N_14825,N_14742,N_14726);
nor U14826 (N_14826,N_14662,N_14707);
xnor U14827 (N_14827,N_14744,N_14663);
xor U14828 (N_14828,N_14656,N_14686);
or U14829 (N_14829,N_14740,N_14694);
xnor U14830 (N_14830,N_14745,N_14742);
nand U14831 (N_14831,N_14669,N_14648);
or U14832 (N_14832,N_14680,N_14682);
or U14833 (N_14833,N_14690,N_14741);
and U14834 (N_14834,N_14705,N_14680);
nand U14835 (N_14835,N_14681,N_14645);
or U14836 (N_14836,N_14712,N_14628);
nor U14837 (N_14837,N_14654,N_14745);
nand U14838 (N_14838,N_14746,N_14636);
nand U14839 (N_14839,N_14631,N_14637);
xor U14840 (N_14840,N_14661,N_14719);
nand U14841 (N_14841,N_14712,N_14745);
xor U14842 (N_14842,N_14679,N_14739);
xor U14843 (N_14843,N_14718,N_14703);
or U14844 (N_14844,N_14716,N_14654);
nor U14845 (N_14845,N_14727,N_14640);
or U14846 (N_14846,N_14664,N_14746);
nand U14847 (N_14847,N_14691,N_14657);
xor U14848 (N_14848,N_14649,N_14680);
nand U14849 (N_14849,N_14698,N_14688);
xnor U14850 (N_14850,N_14641,N_14705);
nor U14851 (N_14851,N_14708,N_14700);
nand U14852 (N_14852,N_14692,N_14695);
xnor U14853 (N_14853,N_14712,N_14655);
and U14854 (N_14854,N_14652,N_14651);
nor U14855 (N_14855,N_14703,N_14663);
nand U14856 (N_14856,N_14634,N_14698);
nand U14857 (N_14857,N_14708,N_14671);
nand U14858 (N_14858,N_14695,N_14735);
nor U14859 (N_14859,N_14713,N_14728);
xnor U14860 (N_14860,N_14716,N_14747);
and U14861 (N_14861,N_14733,N_14636);
nand U14862 (N_14862,N_14634,N_14701);
nor U14863 (N_14863,N_14712,N_14724);
nor U14864 (N_14864,N_14730,N_14682);
nand U14865 (N_14865,N_14644,N_14741);
and U14866 (N_14866,N_14693,N_14697);
and U14867 (N_14867,N_14701,N_14749);
nand U14868 (N_14868,N_14748,N_14711);
nand U14869 (N_14869,N_14725,N_14642);
and U14870 (N_14870,N_14671,N_14654);
nand U14871 (N_14871,N_14673,N_14701);
or U14872 (N_14872,N_14712,N_14674);
nor U14873 (N_14873,N_14649,N_14657);
or U14874 (N_14874,N_14628,N_14695);
or U14875 (N_14875,N_14754,N_14792);
xnor U14876 (N_14876,N_14827,N_14787);
xnor U14877 (N_14877,N_14802,N_14850);
xnor U14878 (N_14878,N_14811,N_14835);
xor U14879 (N_14879,N_14791,N_14818);
xnor U14880 (N_14880,N_14801,N_14821);
nor U14881 (N_14881,N_14793,N_14800);
or U14882 (N_14882,N_14865,N_14790);
nor U14883 (N_14883,N_14779,N_14848);
nand U14884 (N_14884,N_14775,N_14776);
nor U14885 (N_14885,N_14796,N_14770);
and U14886 (N_14886,N_14816,N_14763);
or U14887 (N_14887,N_14863,N_14788);
nor U14888 (N_14888,N_14812,N_14862);
nand U14889 (N_14889,N_14871,N_14766);
nor U14890 (N_14890,N_14784,N_14852);
or U14891 (N_14891,N_14778,N_14771);
xor U14892 (N_14892,N_14782,N_14872);
nand U14893 (N_14893,N_14867,N_14866);
or U14894 (N_14894,N_14750,N_14768);
nor U14895 (N_14895,N_14855,N_14781);
xor U14896 (N_14896,N_14806,N_14815);
nor U14897 (N_14897,N_14842,N_14832);
and U14898 (N_14898,N_14869,N_14772);
xnor U14899 (N_14899,N_14823,N_14861);
nand U14900 (N_14900,N_14847,N_14830);
or U14901 (N_14901,N_14758,N_14769);
nand U14902 (N_14902,N_14783,N_14834);
nand U14903 (N_14903,N_14759,N_14810);
nor U14904 (N_14904,N_14798,N_14809);
nand U14905 (N_14905,N_14761,N_14805);
nand U14906 (N_14906,N_14825,N_14860);
nand U14907 (N_14907,N_14803,N_14837);
nor U14908 (N_14908,N_14757,N_14773);
nor U14909 (N_14909,N_14794,N_14795);
xnor U14910 (N_14910,N_14765,N_14829);
nand U14911 (N_14911,N_14857,N_14822);
or U14912 (N_14912,N_14845,N_14841);
or U14913 (N_14913,N_14836,N_14762);
nand U14914 (N_14914,N_14752,N_14785);
and U14915 (N_14915,N_14824,N_14786);
xor U14916 (N_14916,N_14828,N_14839);
nor U14917 (N_14917,N_14760,N_14856);
xor U14918 (N_14918,N_14764,N_14819);
and U14919 (N_14919,N_14833,N_14804);
nor U14920 (N_14920,N_14826,N_14751);
or U14921 (N_14921,N_14780,N_14756);
xor U14922 (N_14922,N_14874,N_14844);
nand U14923 (N_14923,N_14868,N_14755);
or U14924 (N_14924,N_14859,N_14774);
or U14925 (N_14925,N_14799,N_14864);
nor U14926 (N_14926,N_14840,N_14767);
nand U14927 (N_14927,N_14808,N_14807);
nor U14928 (N_14928,N_14854,N_14813);
nand U14929 (N_14929,N_14817,N_14838);
nand U14930 (N_14930,N_14846,N_14820);
nor U14931 (N_14931,N_14858,N_14849);
nand U14932 (N_14932,N_14797,N_14851);
and U14933 (N_14933,N_14789,N_14873);
xnor U14934 (N_14934,N_14753,N_14777);
nor U14935 (N_14935,N_14870,N_14853);
and U14936 (N_14936,N_14831,N_14814);
nor U14937 (N_14937,N_14843,N_14757);
nor U14938 (N_14938,N_14771,N_14769);
xor U14939 (N_14939,N_14755,N_14854);
nand U14940 (N_14940,N_14833,N_14874);
and U14941 (N_14941,N_14821,N_14755);
nor U14942 (N_14942,N_14764,N_14755);
and U14943 (N_14943,N_14750,N_14870);
xnor U14944 (N_14944,N_14871,N_14869);
nand U14945 (N_14945,N_14854,N_14855);
and U14946 (N_14946,N_14824,N_14760);
nand U14947 (N_14947,N_14867,N_14821);
nand U14948 (N_14948,N_14798,N_14845);
nand U14949 (N_14949,N_14754,N_14845);
xor U14950 (N_14950,N_14774,N_14826);
nor U14951 (N_14951,N_14798,N_14857);
or U14952 (N_14952,N_14813,N_14779);
xor U14953 (N_14953,N_14765,N_14793);
xor U14954 (N_14954,N_14865,N_14847);
nor U14955 (N_14955,N_14816,N_14755);
xor U14956 (N_14956,N_14841,N_14761);
nand U14957 (N_14957,N_14835,N_14843);
nor U14958 (N_14958,N_14751,N_14829);
xnor U14959 (N_14959,N_14855,N_14761);
and U14960 (N_14960,N_14834,N_14814);
or U14961 (N_14961,N_14770,N_14753);
or U14962 (N_14962,N_14750,N_14821);
and U14963 (N_14963,N_14854,N_14848);
or U14964 (N_14964,N_14835,N_14806);
nor U14965 (N_14965,N_14810,N_14854);
and U14966 (N_14966,N_14852,N_14828);
nand U14967 (N_14967,N_14765,N_14772);
xnor U14968 (N_14968,N_14812,N_14761);
nor U14969 (N_14969,N_14842,N_14864);
or U14970 (N_14970,N_14774,N_14802);
and U14971 (N_14971,N_14832,N_14795);
xnor U14972 (N_14972,N_14819,N_14776);
nand U14973 (N_14973,N_14770,N_14872);
or U14974 (N_14974,N_14788,N_14800);
or U14975 (N_14975,N_14855,N_14786);
nor U14976 (N_14976,N_14830,N_14814);
nand U14977 (N_14977,N_14867,N_14865);
xnor U14978 (N_14978,N_14845,N_14800);
nor U14979 (N_14979,N_14797,N_14871);
nor U14980 (N_14980,N_14828,N_14874);
or U14981 (N_14981,N_14782,N_14771);
nand U14982 (N_14982,N_14870,N_14751);
nor U14983 (N_14983,N_14770,N_14838);
or U14984 (N_14984,N_14769,N_14856);
or U14985 (N_14985,N_14771,N_14774);
nor U14986 (N_14986,N_14816,N_14805);
and U14987 (N_14987,N_14791,N_14816);
nor U14988 (N_14988,N_14825,N_14830);
xnor U14989 (N_14989,N_14861,N_14772);
nor U14990 (N_14990,N_14830,N_14868);
nor U14991 (N_14991,N_14759,N_14868);
or U14992 (N_14992,N_14797,N_14791);
or U14993 (N_14993,N_14854,N_14872);
or U14994 (N_14994,N_14753,N_14865);
nand U14995 (N_14995,N_14801,N_14850);
and U14996 (N_14996,N_14753,N_14791);
xor U14997 (N_14997,N_14870,N_14763);
nand U14998 (N_14998,N_14819,N_14829);
xor U14999 (N_14999,N_14834,N_14837);
nor UO_0 (O_0,N_14986,N_14966);
and UO_1 (O_1,N_14977,N_14932);
nor UO_2 (O_2,N_14885,N_14921);
xnor UO_3 (O_3,N_14887,N_14916);
and UO_4 (O_4,N_14883,N_14991);
or UO_5 (O_5,N_14948,N_14965);
or UO_6 (O_6,N_14931,N_14918);
nand UO_7 (O_7,N_14999,N_14930);
nor UO_8 (O_8,N_14996,N_14886);
and UO_9 (O_9,N_14953,N_14968);
xor UO_10 (O_10,N_14954,N_14935);
nand UO_11 (O_11,N_14945,N_14879);
nor UO_12 (O_12,N_14904,N_14944);
or UO_13 (O_13,N_14995,N_14969);
nand UO_14 (O_14,N_14978,N_14951);
xnor UO_15 (O_15,N_14946,N_14892);
nand UO_16 (O_16,N_14898,N_14922);
and UO_17 (O_17,N_14952,N_14983);
and UO_18 (O_18,N_14962,N_14924);
nor UO_19 (O_19,N_14875,N_14956);
nor UO_20 (O_20,N_14972,N_14909);
nand UO_21 (O_21,N_14890,N_14998);
or UO_22 (O_22,N_14888,N_14941);
and UO_23 (O_23,N_14975,N_14915);
xor UO_24 (O_24,N_14876,N_14893);
nand UO_25 (O_25,N_14906,N_14895);
or UO_26 (O_26,N_14907,N_14979);
nand UO_27 (O_27,N_14889,N_14940);
or UO_28 (O_28,N_14896,N_14912);
or UO_29 (O_29,N_14911,N_14936);
nor UO_30 (O_30,N_14994,N_14997);
xor UO_31 (O_31,N_14943,N_14988);
nor UO_32 (O_32,N_14908,N_14963);
xor UO_33 (O_33,N_14891,N_14985);
xnor UO_34 (O_34,N_14938,N_14913);
nor UO_35 (O_35,N_14880,N_14984);
or UO_36 (O_36,N_14981,N_14877);
and UO_37 (O_37,N_14937,N_14964);
and UO_38 (O_38,N_14971,N_14958);
or UO_39 (O_39,N_14974,N_14970);
or UO_40 (O_40,N_14955,N_14894);
or UO_41 (O_41,N_14920,N_14982);
nor UO_42 (O_42,N_14927,N_14933);
or UO_43 (O_43,N_14910,N_14987);
xnor UO_44 (O_44,N_14897,N_14976);
and UO_45 (O_45,N_14950,N_14923);
xor UO_46 (O_46,N_14881,N_14993);
or UO_47 (O_47,N_14960,N_14939);
and UO_48 (O_48,N_14919,N_14989);
xor UO_49 (O_49,N_14905,N_14934);
xnor UO_50 (O_50,N_14917,N_14900);
or UO_51 (O_51,N_14899,N_14878);
or UO_52 (O_52,N_14884,N_14928);
nor UO_53 (O_53,N_14929,N_14925);
nand UO_54 (O_54,N_14926,N_14957);
xnor UO_55 (O_55,N_14961,N_14992);
nor UO_56 (O_56,N_14949,N_14914);
or UO_57 (O_57,N_14882,N_14942);
and UO_58 (O_58,N_14902,N_14967);
xor UO_59 (O_59,N_14959,N_14973);
and UO_60 (O_60,N_14901,N_14980);
xor UO_61 (O_61,N_14947,N_14990);
xnor UO_62 (O_62,N_14903,N_14986);
and UO_63 (O_63,N_14897,N_14938);
nand UO_64 (O_64,N_14938,N_14933);
and UO_65 (O_65,N_14916,N_14906);
and UO_66 (O_66,N_14938,N_14907);
nand UO_67 (O_67,N_14945,N_14952);
nor UO_68 (O_68,N_14921,N_14977);
xor UO_69 (O_69,N_14914,N_14967);
nor UO_70 (O_70,N_14880,N_14994);
xnor UO_71 (O_71,N_14962,N_14911);
nor UO_72 (O_72,N_14967,N_14981);
and UO_73 (O_73,N_14950,N_14953);
or UO_74 (O_74,N_14876,N_14980);
nand UO_75 (O_75,N_14942,N_14970);
nor UO_76 (O_76,N_14901,N_14940);
nand UO_77 (O_77,N_14916,N_14902);
and UO_78 (O_78,N_14931,N_14941);
and UO_79 (O_79,N_14889,N_14909);
nor UO_80 (O_80,N_14981,N_14996);
nand UO_81 (O_81,N_14930,N_14993);
and UO_82 (O_82,N_14919,N_14929);
nor UO_83 (O_83,N_14950,N_14960);
nand UO_84 (O_84,N_14906,N_14945);
and UO_85 (O_85,N_14901,N_14875);
and UO_86 (O_86,N_14897,N_14921);
nor UO_87 (O_87,N_14933,N_14895);
xnor UO_88 (O_88,N_14948,N_14898);
nand UO_89 (O_89,N_14958,N_14930);
nor UO_90 (O_90,N_14882,N_14884);
nor UO_91 (O_91,N_14940,N_14956);
nor UO_92 (O_92,N_14927,N_14957);
and UO_93 (O_93,N_14926,N_14905);
nand UO_94 (O_94,N_14931,N_14888);
and UO_95 (O_95,N_14971,N_14940);
nor UO_96 (O_96,N_14991,N_14956);
or UO_97 (O_97,N_14907,N_14968);
xor UO_98 (O_98,N_14995,N_14910);
xnor UO_99 (O_99,N_14978,N_14896);
or UO_100 (O_100,N_14962,N_14887);
nor UO_101 (O_101,N_14959,N_14895);
nor UO_102 (O_102,N_14916,N_14968);
xnor UO_103 (O_103,N_14898,N_14921);
nor UO_104 (O_104,N_14925,N_14962);
and UO_105 (O_105,N_14985,N_14965);
xnor UO_106 (O_106,N_14976,N_14948);
nor UO_107 (O_107,N_14970,N_14961);
nand UO_108 (O_108,N_14959,N_14964);
xor UO_109 (O_109,N_14984,N_14920);
or UO_110 (O_110,N_14901,N_14883);
and UO_111 (O_111,N_14885,N_14882);
nand UO_112 (O_112,N_14902,N_14962);
nor UO_113 (O_113,N_14909,N_14899);
or UO_114 (O_114,N_14964,N_14928);
and UO_115 (O_115,N_14928,N_14908);
xnor UO_116 (O_116,N_14954,N_14884);
xor UO_117 (O_117,N_14931,N_14920);
and UO_118 (O_118,N_14942,N_14892);
xor UO_119 (O_119,N_14970,N_14972);
and UO_120 (O_120,N_14910,N_14929);
or UO_121 (O_121,N_14913,N_14987);
nor UO_122 (O_122,N_14968,N_14946);
or UO_123 (O_123,N_14903,N_14959);
xor UO_124 (O_124,N_14978,N_14994);
nand UO_125 (O_125,N_14936,N_14964);
or UO_126 (O_126,N_14967,N_14892);
nand UO_127 (O_127,N_14970,N_14962);
nand UO_128 (O_128,N_14880,N_14877);
nand UO_129 (O_129,N_14932,N_14999);
nand UO_130 (O_130,N_14907,N_14951);
and UO_131 (O_131,N_14908,N_14904);
nor UO_132 (O_132,N_14878,N_14994);
and UO_133 (O_133,N_14973,N_14944);
or UO_134 (O_134,N_14905,N_14939);
nand UO_135 (O_135,N_14956,N_14896);
nor UO_136 (O_136,N_14996,N_14922);
xnor UO_137 (O_137,N_14918,N_14906);
nand UO_138 (O_138,N_14942,N_14961);
or UO_139 (O_139,N_14890,N_14977);
xnor UO_140 (O_140,N_14908,N_14891);
nand UO_141 (O_141,N_14984,N_14985);
and UO_142 (O_142,N_14896,N_14932);
or UO_143 (O_143,N_14890,N_14930);
or UO_144 (O_144,N_14962,N_14918);
nand UO_145 (O_145,N_14996,N_14906);
nand UO_146 (O_146,N_14974,N_14923);
and UO_147 (O_147,N_14928,N_14930);
or UO_148 (O_148,N_14949,N_14920);
or UO_149 (O_149,N_14958,N_14998);
or UO_150 (O_150,N_14925,N_14944);
nor UO_151 (O_151,N_14992,N_14957);
nor UO_152 (O_152,N_14965,N_14954);
nor UO_153 (O_153,N_14922,N_14892);
or UO_154 (O_154,N_14977,N_14908);
xnor UO_155 (O_155,N_14981,N_14940);
and UO_156 (O_156,N_14980,N_14993);
xnor UO_157 (O_157,N_14880,N_14937);
nand UO_158 (O_158,N_14973,N_14967);
xor UO_159 (O_159,N_14926,N_14970);
xnor UO_160 (O_160,N_14941,N_14997);
nor UO_161 (O_161,N_14899,N_14978);
or UO_162 (O_162,N_14962,N_14907);
xnor UO_163 (O_163,N_14997,N_14883);
xnor UO_164 (O_164,N_14995,N_14973);
nand UO_165 (O_165,N_14940,N_14929);
or UO_166 (O_166,N_14993,N_14887);
nor UO_167 (O_167,N_14986,N_14994);
nand UO_168 (O_168,N_14894,N_14889);
or UO_169 (O_169,N_14906,N_14939);
and UO_170 (O_170,N_14882,N_14893);
nor UO_171 (O_171,N_14897,N_14915);
nand UO_172 (O_172,N_14897,N_14995);
nor UO_173 (O_173,N_14919,N_14925);
xnor UO_174 (O_174,N_14969,N_14976);
nor UO_175 (O_175,N_14909,N_14976);
nand UO_176 (O_176,N_14924,N_14906);
and UO_177 (O_177,N_14876,N_14959);
nor UO_178 (O_178,N_14956,N_14942);
nand UO_179 (O_179,N_14927,N_14917);
and UO_180 (O_180,N_14964,N_14982);
nand UO_181 (O_181,N_14894,N_14926);
xnor UO_182 (O_182,N_14991,N_14907);
nand UO_183 (O_183,N_14926,N_14923);
and UO_184 (O_184,N_14934,N_14947);
xnor UO_185 (O_185,N_14982,N_14896);
xnor UO_186 (O_186,N_14918,N_14898);
and UO_187 (O_187,N_14942,N_14900);
nand UO_188 (O_188,N_14881,N_14996);
and UO_189 (O_189,N_14962,N_14895);
nand UO_190 (O_190,N_14914,N_14972);
nand UO_191 (O_191,N_14918,N_14919);
and UO_192 (O_192,N_14996,N_14915);
and UO_193 (O_193,N_14903,N_14973);
nor UO_194 (O_194,N_14992,N_14885);
xnor UO_195 (O_195,N_14914,N_14927);
nor UO_196 (O_196,N_14924,N_14907);
nor UO_197 (O_197,N_14994,N_14949);
nand UO_198 (O_198,N_14958,N_14990);
nor UO_199 (O_199,N_14917,N_14904);
nand UO_200 (O_200,N_14990,N_14892);
or UO_201 (O_201,N_14915,N_14980);
xor UO_202 (O_202,N_14979,N_14887);
xnor UO_203 (O_203,N_14959,N_14946);
nand UO_204 (O_204,N_14895,N_14999);
and UO_205 (O_205,N_14940,N_14946);
and UO_206 (O_206,N_14903,N_14902);
nor UO_207 (O_207,N_14940,N_14886);
xor UO_208 (O_208,N_14927,N_14975);
nand UO_209 (O_209,N_14931,N_14890);
xnor UO_210 (O_210,N_14916,N_14878);
and UO_211 (O_211,N_14985,N_14928);
or UO_212 (O_212,N_14996,N_14999);
or UO_213 (O_213,N_14927,N_14995);
nand UO_214 (O_214,N_14906,N_14988);
xor UO_215 (O_215,N_14953,N_14976);
and UO_216 (O_216,N_14984,N_14969);
or UO_217 (O_217,N_14890,N_14979);
or UO_218 (O_218,N_14892,N_14972);
nor UO_219 (O_219,N_14894,N_14957);
or UO_220 (O_220,N_14933,N_14901);
nand UO_221 (O_221,N_14934,N_14998);
xnor UO_222 (O_222,N_14964,N_14960);
nor UO_223 (O_223,N_14980,N_14879);
nor UO_224 (O_224,N_14925,N_14915);
and UO_225 (O_225,N_14890,N_14918);
nor UO_226 (O_226,N_14906,N_14975);
or UO_227 (O_227,N_14991,N_14895);
nor UO_228 (O_228,N_14882,N_14977);
xnor UO_229 (O_229,N_14930,N_14949);
or UO_230 (O_230,N_14986,N_14891);
nor UO_231 (O_231,N_14925,N_14899);
or UO_232 (O_232,N_14990,N_14916);
nand UO_233 (O_233,N_14901,N_14939);
or UO_234 (O_234,N_14878,N_14910);
and UO_235 (O_235,N_14922,N_14994);
and UO_236 (O_236,N_14992,N_14930);
and UO_237 (O_237,N_14945,N_14979);
xor UO_238 (O_238,N_14995,N_14908);
or UO_239 (O_239,N_14880,N_14934);
and UO_240 (O_240,N_14923,N_14889);
nor UO_241 (O_241,N_14981,N_14887);
or UO_242 (O_242,N_14970,N_14955);
and UO_243 (O_243,N_14977,N_14939);
xnor UO_244 (O_244,N_14938,N_14878);
xnor UO_245 (O_245,N_14971,N_14990);
nor UO_246 (O_246,N_14896,N_14924);
nand UO_247 (O_247,N_14998,N_14940);
nand UO_248 (O_248,N_14998,N_14975);
xnor UO_249 (O_249,N_14973,N_14910);
or UO_250 (O_250,N_14915,N_14883);
or UO_251 (O_251,N_14944,N_14912);
nor UO_252 (O_252,N_14959,N_14995);
xor UO_253 (O_253,N_14906,N_14929);
xnor UO_254 (O_254,N_14949,N_14974);
nor UO_255 (O_255,N_14904,N_14930);
and UO_256 (O_256,N_14953,N_14910);
or UO_257 (O_257,N_14994,N_14933);
or UO_258 (O_258,N_14963,N_14999);
nor UO_259 (O_259,N_14915,N_14971);
nand UO_260 (O_260,N_14918,N_14888);
nor UO_261 (O_261,N_14947,N_14909);
nor UO_262 (O_262,N_14979,N_14917);
nand UO_263 (O_263,N_14999,N_14919);
or UO_264 (O_264,N_14940,N_14995);
nand UO_265 (O_265,N_14984,N_14974);
or UO_266 (O_266,N_14935,N_14900);
xor UO_267 (O_267,N_14919,N_14980);
nand UO_268 (O_268,N_14962,N_14933);
nand UO_269 (O_269,N_14943,N_14944);
xnor UO_270 (O_270,N_14931,N_14883);
xnor UO_271 (O_271,N_14937,N_14989);
nor UO_272 (O_272,N_14985,N_14907);
and UO_273 (O_273,N_14892,N_14999);
or UO_274 (O_274,N_14916,N_14991);
or UO_275 (O_275,N_14974,N_14890);
nand UO_276 (O_276,N_14911,N_14930);
or UO_277 (O_277,N_14951,N_14939);
nor UO_278 (O_278,N_14929,N_14952);
xor UO_279 (O_279,N_14996,N_14893);
nor UO_280 (O_280,N_14940,N_14892);
or UO_281 (O_281,N_14991,N_14965);
and UO_282 (O_282,N_14945,N_14968);
xnor UO_283 (O_283,N_14952,N_14890);
nand UO_284 (O_284,N_14967,N_14880);
or UO_285 (O_285,N_14902,N_14929);
nor UO_286 (O_286,N_14943,N_14889);
xnor UO_287 (O_287,N_14930,N_14984);
nand UO_288 (O_288,N_14891,N_14886);
nor UO_289 (O_289,N_14906,N_14925);
and UO_290 (O_290,N_14966,N_14942);
nor UO_291 (O_291,N_14919,N_14985);
xor UO_292 (O_292,N_14879,N_14968);
and UO_293 (O_293,N_14966,N_14943);
and UO_294 (O_294,N_14880,N_14887);
and UO_295 (O_295,N_14887,N_14965);
nand UO_296 (O_296,N_14967,N_14930);
nor UO_297 (O_297,N_14894,N_14935);
nand UO_298 (O_298,N_14882,N_14989);
or UO_299 (O_299,N_14926,N_14908);
xor UO_300 (O_300,N_14926,N_14875);
or UO_301 (O_301,N_14892,N_14970);
nand UO_302 (O_302,N_14923,N_14955);
nor UO_303 (O_303,N_14894,N_14989);
nand UO_304 (O_304,N_14899,N_14923);
and UO_305 (O_305,N_14978,N_14937);
nor UO_306 (O_306,N_14902,N_14885);
or UO_307 (O_307,N_14905,N_14992);
and UO_308 (O_308,N_14911,N_14958);
or UO_309 (O_309,N_14923,N_14902);
or UO_310 (O_310,N_14898,N_14939);
and UO_311 (O_311,N_14944,N_14999);
nand UO_312 (O_312,N_14894,N_14893);
or UO_313 (O_313,N_14978,N_14959);
xnor UO_314 (O_314,N_14935,N_14960);
xor UO_315 (O_315,N_14931,N_14975);
xor UO_316 (O_316,N_14985,N_14925);
nand UO_317 (O_317,N_14929,N_14971);
nand UO_318 (O_318,N_14949,N_14966);
xor UO_319 (O_319,N_14891,N_14975);
or UO_320 (O_320,N_14875,N_14885);
and UO_321 (O_321,N_14937,N_14980);
xnor UO_322 (O_322,N_14906,N_14961);
or UO_323 (O_323,N_14997,N_14978);
xnor UO_324 (O_324,N_14913,N_14993);
nand UO_325 (O_325,N_14884,N_14976);
nand UO_326 (O_326,N_14945,N_14933);
or UO_327 (O_327,N_14979,N_14989);
nand UO_328 (O_328,N_14900,N_14968);
nand UO_329 (O_329,N_14908,N_14956);
nand UO_330 (O_330,N_14995,N_14879);
nor UO_331 (O_331,N_14955,N_14979);
or UO_332 (O_332,N_14933,N_14952);
xor UO_333 (O_333,N_14980,N_14903);
xnor UO_334 (O_334,N_14938,N_14948);
nand UO_335 (O_335,N_14955,N_14912);
and UO_336 (O_336,N_14886,N_14918);
and UO_337 (O_337,N_14945,N_14882);
nand UO_338 (O_338,N_14922,N_14987);
nand UO_339 (O_339,N_14902,N_14936);
nor UO_340 (O_340,N_14990,N_14997);
nand UO_341 (O_341,N_14995,N_14950);
and UO_342 (O_342,N_14932,N_14886);
or UO_343 (O_343,N_14957,N_14879);
nor UO_344 (O_344,N_14963,N_14957);
or UO_345 (O_345,N_14951,N_14950);
xnor UO_346 (O_346,N_14934,N_14970);
xnor UO_347 (O_347,N_14895,N_14916);
and UO_348 (O_348,N_14946,N_14890);
or UO_349 (O_349,N_14976,N_14954);
nor UO_350 (O_350,N_14966,N_14878);
nor UO_351 (O_351,N_14979,N_14891);
nor UO_352 (O_352,N_14876,N_14995);
or UO_353 (O_353,N_14915,N_14935);
and UO_354 (O_354,N_14961,N_14952);
and UO_355 (O_355,N_14993,N_14997);
or UO_356 (O_356,N_14977,N_14919);
and UO_357 (O_357,N_14994,N_14912);
nand UO_358 (O_358,N_14969,N_14955);
or UO_359 (O_359,N_14943,N_14971);
and UO_360 (O_360,N_14893,N_14895);
xor UO_361 (O_361,N_14932,N_14971);
xor UO_362 (O_362,N_14974,N_14911);
nand UO_363 (O_363,N_14948,N_14995);
or UO_364 (O_364,N_14956,N_14886);
nand UO_365 (O_365,N_14890,N_14901);
xor UO_366 (O_366,N_14972,N_14912);
nor UO_367 (O_367,N_14881,N_14883);
and UO_368 (O_368,N_14935,N_14963);
xor UO_369 (O_369,N_14989,N_14891);
and UO_370 (O_370,N_14967,N_14942);
or UO_371 (O_371,N_14943,N_14911);
nor UO_372 (O_372,N_14963,N_14937);
xnor UO_373 (O_373,N_14919,N_14938);
nor UO_374 (O_374,N_14977,N_14980);
xor UO_375 (O_375,N_14919,N_14891);
or UO_376 (O_376,N_14974,N_14886);
or UO_377 (O_377,N_14994,N_14906);
nand UO_378 (O_378,N_14890,N_14951);
xnor UO_379 (O_379,N_14886,N_14939);
nor UO_380 (O_380,N_14935,N_14977);
and UO_381 (O_381,N_14882,N_14904);
xor UO_382 (O_382,N_14908,N_14947);
or UO_383 (O_383,N_14891,N_14931);
and UO_384 (O_384,N_14900,N_14962);
and UO_385 (O_385,N_14890,N_14926);
or UO_386 (O_386,N_14933,N_14970);
nand UO_387 (O_387,N_14947,N_14937);
nor UO_388 (O_388,N_14963,N_14994);
nand UO_389 (O_389,N_14969,N_14989);
and UO_390 (O_390,N_14898,N_14978);
nor UO_391 (O_391,N_14916,N_14894);
nor UO_392 (O_392,N_14962,N_14930);
nor UO_393 (O_393,N_14887,N_14935);
nor UO_394 (O_394,N_14942,N_14950);
nor UO_395 (O_395,N_14992,N_14897);
nand UO_396 (O_396,N_14938,N_14917);
nor UO_397 (O_397,N_14975,N_14970);
and UO_398 (O_398,N_14948,N_14979);
nor UO_399 (O_399,N_14885,N_14998);
and UO_400 (O_400,N_14989,N_14988);
nand UO_401 (O_401,N_14997,N_14939);
nor UO_402 (O_402,N_14893,N_14960);
xnor UO_403 (O_403,N_14991,N_14959);
nand UO_404 (O_404,N_14879,N_14963);
or UO_405 (O_405,N_14974,N_14995);
and UO_406 (O_406,N_14897,N_14896);
nand UO_407 (O_407,N_14932,N_14942);
nor UO_408 (O_408,N_14919,N_14941);
xor UO_409 (O_409,N_14889,N_14995);
xor UO_410 (O_410,N_14928,N_14971);
nor UO_411 (O_411,N_14969,N_14931);
and UO_412 (O_412,N_14988,N_14905);
nand UO_413 (O_413,N_14922,N_14901);
nand UO_414 (O_414,N_14882,N_14892);
xor UO_415 (O_415,N_14997,N_14936);
or UO_416 (O_416,N_14890,N_14932);
nor UO_417 (O_417,N_14895,N_14897);
xnor UO_418 (O_418,N_14989,N_14908);
or UO_419 (O_419,N_14971,N_14970);
nand UO_420 (O_420,N_14943,N_14900);
and UO_421 (O_421,N_14964,N_14974);
nor UO_422 (O_422,N_14987,N_14907);
or UO_423 (O_423,N_14934,N_14969);
xnor UO_424 (O_424,N_14942,N_14989);
and UO_425 (O_425,N_14883,N_14957);
nand UO_426 (O_426,N_14912,N_14982);
nor UO_427 (O_427,N_14966,N_14934);
or UO_428 (O_428,N_14946,N_14939);
xnor UO_429 (O_429,N_14998,N_14876);
nor UO_430 (O_430,N_14895,N_14929);
and UO_431 (O_431,N_14953,N_14993);
nor UO_432 (O_432,N_14877,N_14931);
nand UO_433 (O_433,N_14902,N_14909);
xnor UO_434 (O_434,N_14922,N_14881);
nand UO_435 (O_435,N_14987,N_14916);
xnor UO_436 (O_436,N_14988,N_14923);
and UO_437 (O_437,N_14940,N_14958);
or UO_438 (O_438,N_14989,N_14971);
nand UO_439 (O_439,N_14946,N_14879);
or UO_440 (O_440,N_14970,N_14950);
nand UO_441 (O_441,N_14960,N_14981);
and UO_442 (O_442,N_14940,N_14910);
and UO_443 (O_443,N_14908,N_14992);
or UO_444 (O_444,N_14930,N_14991);
or UO_445 (O_445,N_14965,N_14997);
nor UO_446 (O_446,N_14984,N_14925);
nand UO_447 (O_447,N_14965,N_14930);
or UO_448 (O_448,N_14960,N_14895);
xor UO_449 (O_449,N_14887,N_14952);
or UO_450 (O_450,N_14937,N_14899);
or UO_451 (O_451,N_14970,N_14925);
and UO_452 (O_452,N_14910,N_14908);
nand UO_453 (O_453,N_14942,N_14899);
xnor UO_454 (O_454,N_14942,N_14949);
or UO_455 (O_455,N_14975,N_14876);
and UO_456 (O_456,N_14931,N_14972);
and UO_457 (O_457,N_14875,N_14941);
and UO_458 (O_458,N_14986,N_14952);
nand UO_459 (O_459,N_14967,N_14936);
and UO_460 (O_460,N_14935,N_14931);
nor UO_461 (O_461,N_14951,N_14987);
nor UO_462 (O_462,N_14917,N_14930);
xnor UO_463 (O_463,N_14911,N_14885);
xnor UO_464 (O_464,N_14877,N_14912);
and UO_465 (O_465,N_14875,N_14973);
or UO_466 (O_466,N_14985,N_14901);
nor UO_467 (O_467,N_14998,N_14980);
and UO_468 (O_468,N_14982,N_14886);
and UO_469 (O_469,N_14947,N_14955);
or UO_470 (O_470,N_14899,N_14912);
or UO_471 (O_471,N_14903,N_14897);
or UO_472 (O_472,N_14959,N_14948);
or UO_473 (O_473,N_14924,N_14888);
and UO_474 (O_474,N_14930,N_14923);
nand UO_475 (O_475,N_14881,N_14895);
nand UO_476 (O_476,N_14902,N_14947);
and UO_477 (O_477,N_14987,N_14970);
nand UO_478 (O_478,N_14995,N_14929);
nor UO_479 (O_479,N_14885,N_14912);
nor UO_480 (O_480,N_14921,N_14925);
nor UO_481 (O_481,N_14986,N_14976);
xor UO_482 (O_482,N_14878,N_14958);
nor UO_483 (O_483,N_14979,N_14970);
xnor UO_484 (O_484,N_14881,N_14887);
nor UO_485 (O_485,N_14997,N_14974);
or UO_486 (O_486,N_14952,N_14889);
nand UO_487 (O_487,N_14897,N_14880);
or UO_488 (O_488,N_14998,N_14899);
xor UO_489 (O_489,N_14917,N_14892);
nor UO_490 (O_490,N_14956,N_14944);
and UO_491 (O_491,N_14973,N_14980);
nand UO_492 (O_492,N_14913,N_14970);
nor UO_493 (O_493,N_14945,N_14972);
xnor UO_494 (O_494,N_14959,N_14937);
nor UO_495 (O_495,N_14944,N_14993);
nor UO_496 (O_496,N_14931,N_14932);
and UO_497 (O_497,N_14946,N_14984);
xnor UO_498 (O_498,N_14876,N_14892);
xnor UO_499 (O_499,N_14982,N_14975);
nand UO_500 (O_500,N_14941,N_14905);
and UO_501 (O_501,N_14962,N_14961);
nor UO_502 (O_502,N_14897,N_14980);
xor UO_503 (O_503,N_14919,N_14902);
and UO_504 (O_504,N_14900,N_14947);
xor UO_505 (O_505,N_14994,N_14890);
nand UO_506 (O_506,N_14995,N_14962);
or UO_507 (O_507,N_14969,N_14904);
and UO_508 (O_508,N_14990,N_14951);
and UO_509 (O_509,N_14956,N_14917);
or UO_510 (O_510,N_14931,N_14934);
nand UO_511 (O_511,N_14901,N_14957);
nand UO_512 (O_512,N_14979,N_14909);
or UO_513 (O_513,N_14909,N_14929);
nor UO_514 (O_514,N_14989,N_14946);
and UO_515 (O_515,N_14904,N_14979);
nor UO_516 (O_516,N_14945,N_14885);
nor UO_517 (O_517,N_14985,N_14889);
nor UO_518 (O_518,N_14949,N_14950);
or UO_519 (O_519,N_14978,N_14957);
or UO_520 (O_520,N_14990,N_14904);
nand UO_521 (O_521,N_14895,N_14968);
and UO_522 (O_522,N_14920,N_14966);
and UO_523 (O_523,N_14941,N_14904);
nor UO_524 (O_524,N_14919,N_14991);
or UO_525 (O_525,N_14957,N_14896);
nor UO_526 (O_526,N_14903,N_14963);
nor UO_527 (O_527,N_14907,N_14897);
nand UO_528 (O_528,N_14939,N_14902);
and UO_529 (O_529,N_14979,N_14943);
nand UO_530 (O_530,N_14937,N_14884);
and UO_531 (O_531,N_14981,N_14933);
or UO_532 (O_532,N_14914,N_14973);
xor UO_533 (O_533,N_14901,N_14938);
nand UO_534 (O_534,N_14972,N_14881);
or UO_535 (O_535,N_14985,N_14900);
and UO_536 (O_536,N_14964,N_14953);
nand UO_537 (O_537,N_14976,N_14913);
or UO_538 (O_538,N_14898,N_14970);
xnor UO_539 (O_539,N_14962,N_14886);
nand UO_540 (O_540,N_14912,N_14959);
or UO_541 (O_541,N_14940,N_14953);
nor UO_542 (O_542,N_14925,N_14889);
and UO_543 (O_543,N_14990,N_14983);
xor UO_544 (O_544,N_14946,N_14953);
nor UO_545 (O_545,N_14953,N_14959);
nand UO_546 (O_546,N_14985,N_14896);
xnor UO_547 (O_547,N_14911,N_14881);
nor UO_548 (O_548,N_14960,N_14894);
and UO_549 (O_549,N_14910,N_14899);
xnor UO_550 (O_550,N_14967,N_14888);
nand UO_551 (O_551,N_14947,N_14962);
and UO_552 (O_552,N_14961,N_14889);
nor UO_553 (O_553,N_14979,N_14897);
or UO_554 (O_554,N_14943,N_14894);
and UO_555 (O_555,N_14984,N_14965);
nand UO_556 (O_556,N_14901,N_14889);
nor UO_557 (O_557,N_14909,N_14910);
nand UO_558 (O_558,N_14881,N_14893);
xor UO_559 (O_559,N_14895,N_14942);
nand UO_560 (O_560,N_14990,N_14931);
nand UO_561 (O_561,N_14963,N_14909);
nand UO_562 (O_562,N_14933,N_14942);
and UO_563 (O_563,N_14933,N_14953);
or UO_564 (O_564,N_14978,N_14886);
or UO_565 (O_565,N_14938,N_14937);
nor UO_566 (O_566,N_14933,N_14916);
or UO_567 (O_567,N_14990,N_14946);
or UO_568 (O_568,N_14898,N_14963);
xor UO_569 (O_569,N_14938,N_14984);
nor UO_570 (O_570,N_14912,N_14943);
or UO_571 (O_571,N_14899,N_14911);
or UO_572 (O_572,N_14906,N_14893);
or UO_573 (O_573,N_14985,N_14927);
nand UO_574 (O_574,N_14977,N_14941);
and UO_575 (O_575,N_14953,N_14955);
and UO_576 (O_576,N_14920,N_14980);
and UO_577 (O_577,N_14949,N_14883);
and UO_578 (O_578,N_14976,N_14983);
nand UO_579 (O_579,N_14920,N_14935);
xor UO_580 (O_580,N_14951,N_14914);
and UO_581 (O_581,N_14976,N_14925);
xor UO_582 (O_582,N_14941,N_14947);
nor UO_583 (O_583,N_14887,N_14950);
xnor UO_584 (O_584,N_14925,N_14930);
and UO_585 (O_585,N_14959,N_14880);
nand UO_586 (O_586,N_14920,N_14904);
and UO_587 (O_587,N_14932,N_14953);
nor UO_588 (O_588,N_14962,N_14994);
xor UO_589 (O_589,N_14910,N_14934);
nor UO_590 (O_590,N_14999,N_14971);
nor UO_591 (O_591,N_14975,N_14942);
xor UO_592 (O_592,N_14969,N_14972);
nor UO_593 (O_593,N_14941,N_14934);
and UO_594 (O_594,N_14890,N_14922);
nor UO_595 (O_595,N_14926,N_14973);
and UO_596 (O_596,N_14947,N_14989);
or UO_597 (O_597,N_14930,N_14956);
nor UO_598 (O_598,N_14887,N_14940);
xnor UO_599 (O_599,N_14899,N_14996);
and UO_600 (O_600,N_14927,N_14891);
nand UO_601 (O_601,N_14943,N_14932);
and UO_602 (O_602,N_14886,N_14899);
nor UO_603 (O_603,N_14915,N_14924);
nor UO_604 (O_604,N_14979,N_14985);
nor UO_605 (O_605,N_14988,N_14926);
nand UO_606 (O_606,N_14970,N_14888);
nor UO_607 (O_607,N_14947,N_14967);
nor UO_608 (O_608,N_14880,N_14996);
nand UO_609 (O_609,N_14883,N_14897);
or UO_610 (O_610,N_14887,N_14894);
and UO_611 (O_611,N_14951,N_14927);
and UO_612 (O_612,N_14893,N_14966);
and UO_613 (O_613,N_14882,N_14896);
xor UO_614 (O_614,N_14957,N_14946);
and UO_615 (O_615,N_14921,N_14916);
or UO_616 (O_616,N_14878,N_14987);
nand UO_617 (O_617,N_14925,N_14956);
nor UO_618 (O_618,N_14953,N_14952);
xnor UO_619 (O_619,N_14937,N_14936);
or UO_620 (O_620,N_14982,N_14994);
and UO_621 (O_621,N_14931,N_14927);
or UO_622 (O_622,N_14878,N_14882);
nand UO_623 (O_623,N_14978,N_14908);
nor UO_624 (O_624,N_14968,N_14963);
or UO_625 (O_625,N_14956,N_14983);
or UO_626 (O_626,N_14926,N_14910);
or UO_627 (O_627,N_14954,N_14947);
nor UO_628 (O_628,N_14875,N_14968);
nor UO_629 (O_629,N_14875,N_14896);
xnor UO_630 (O_630,N_14923,N_14986);
or UO_631 (O_631,N_14941,N_14895);
nor UO_632 (O_632,N_14881,N_14984);
xor UO_633 (O_633,N_14952,N_14905);
or UO_634 (O_634,N_14982,N_14938);
or UO_635 (O_635,N_14999,N_14975);
and UO_636 (O_636,N_14936,N_14935);
or UO_637 (O_637,N_14909,N_14944);
and UO_638 (O_638,N_14997,N_14905);
or UO_639 (O_639,N_14902,N_14948);
or UO_640 (O_640,N_14982,N_14883);
nor UO_641 (O_641,N_14924,N_14902);
or UO_642 (O_642,N_14945,N_14920);
xor UO_643 (O_643,N_14941,N_14883);
nor UO_644 (O_644,N_14921,N_14900);
xor UO_645 (O_645,N_14989,N_14880);
and UO_646 (O_646,N_14913,N_14928);
and UO_647 (O_647,N_14930,N_14953);
and UO_648 (O_648,N_14916,N_14918);
or UO_649 (O_649,N_14914,N_14948);
nand UO_650 (O_650,N_14932,N_14973);
xor UO_651 (O_651,N_14953,N_14956);
and UO_652 (O_652,N_14977,N_14956);
and UO_653 (O_653,N_14891,N_14955);
nor UO_654 (O_654,N_14980,N_14918);
xnor UO_655 (O_655,N_14923,N_14917);
nand UO_656 (O_656,N_14965,N_14922);
xor UO_657 (O_657,N_14934,N_14904);
nor UO_658 (O_658,N_14889,N_14893);
nand UO_659 (O_659,N_14999,N_14879);
nor UO_660 (O_660,N_14963,N_14917);
and UO_661 (O_661,N_14914,N_14922);
or UO_662 (O_662,N_14875,N_14994);
xnor UO_663 (O_663,N_14917,N_14896);
and UO_664 (O_664,N_14955,N_14996);
nor UO_665 (O_665,N_14945,N_14953);
nor UO_666 (O_666,N_14921,N_14906);
nor UO_667 (O_667,N_14875,N_14951);
or UO_668 (O_668,N_14967,N_14926);
and UO_669 (O_669,N_14884,N_14952);
nor UO_670 (O_670,N_14927,N_14979);
xnor UO_671 (O_671,N_14898,N_14953);
or UO_672 (O_672,N_14986,N_14930);
nand UO_673 (O_673,N_14875,N_14971);
nand UO_674 (O_674,N_14951,N_14996);
or UO_675 (O_675,N_14952,N_14928);
nor UO_676 (O_676,N_14917,N_14922);
and UO_677 (O_677,N_14971,N_14904);
or UO_678 (O_678,N_14958,N_14989);
nand UO_679 (O_679,N_14985,N_14981);
xor UO_680 (O_680,N_14981,N_14902);
nand UO_681 (O_681,N_14963,N_14962);
nand UO_682 (O_682,N_14899,N_14885);
xor UO_683 (O_683,N_14978,N_14930);
xor UO_684 (O_684,N_14985,N_14921);
and UO_685 (O_685,N_14984,N_14976);
and UO_686 (O_686,N_14896,N_14887);
or UO_687 (O_687,N_14915,N_14999);
or UO_688 (O_688,N_14945,N_14886);
xor UO_689 (O_689,N_14925,N_14926);
nand UO_690 (O_690,N_14999,N_14877);
nor UO_691 (O_691,N_14876,N_14966);
nand UO_692 (O_692,N_14888,N_14977);
or UO_693 (O_693,N_14975,N_14986);
xnor UO_694 (O_694,N_14912,N_14910);
xnor UO_695 (O_695,N_14917,N_14913);
and UO_696 (O_696,N_14909,N_14975);
xnor UO_697 (O_697,N_14988,N_14933);
or UO_698 (O_698,N_14946,N_14875);
nor UO_699 (O_699,N_14945,N_14905);
nand UO_700 (O_700,N_14912,N_14942);
xor UO_701 (O_701,N_14906,N_14958);
xnor UO_702 (O_702,N_14893,N_14884);
and UO_703 (O_703,N_14955,N_14911);
xnor UO_704 (O_704,N_14900,N_14887);
nand UO_705 (O_705,N_14987,N_14883);
and UO_706 (O_706,N_14889,N_14963);
xnor UO_707 (O_707,N_14889,N_14960);
or UO_708 (O_708,N_14981,N_14931);
nor UO_709 (O_709,N_14932,N_14888);
nor UO_710 (O_710,N_14938,N_14884);
nand UO_711 (O_711,N_14983,N_14926);
and UO_712 (O_712,N_14990,N_14982);
nor UO_713 (O_713,N_14973,N_14925);
nand UO_714 (O_714,N_14912,N_14891);
and UO_715 (O_715,N_14885,N_14970);
and UO_716 (O_716,N_14935,N_14918);
nor UO_717 (O_717,N_14893,N_14929);
or UO_718 (O_718,N_14901,N_14929);
and UO_719 (O_719,N_14993,N_14935);
xor UO_720 (O_720,N_14912,N_14932);
and UO_721 (O_721,N_14986,N_14924);
and UO_722 (O_722,N_14899,N_14936);
or UO_723 (O_723,N_14990,N_14979);
xor UO_724 (O_724,N_14896,N_14939);
nor UO_725 (O_725,N_14982,N_14948);
nand UO_726 (O_726,N_14946,N_14975);
and UO_727 (O_727,N_14886,N_14979);
nand UO_728 (O_728,N_14952,N_14988);
nand UO_729 (O_729,N_14891,N_14945);
and UO_730 (O_730,N_14909,N_14933);
nand UO_731 (O_731,N_14909,N_14966);
xor UO_732 (O_732,N_14923,N_14893);
nor UO_733 (O_733,N_14908,N_14964);
or UO_734 (O_734,N_14966,N_14955);
or UO_735 (O_735,N_14986,N_14967);
nand UO_736 (O_736,N_14884,N_14916);
nor UO_737 (O_737,N_14949,N_14899);
and UO_738 (O_738,N_14886,N_14977);
xnor UO_739 (O_739,N_14877,N_14917);
nor UO_740 (O_740,N_14921,N_14939);
xor UO_741 (O_741,N_14929,N_14928);
or UO_742 (O_742,N_14963,N_14991);
nor UO_743 (O_743,N_14903,N_14989);
nand UO_744 (O_744,N_14985,N_14975);
or UO_745 (O_745,N_14943,N_14934);
nor UO_746 (O_746,N_14973,N_14989);
and UO_747 (O_747,N_14928,N_14881);
and UO_748 (O_748,N_14889,N_14984);
xnor UO_749 (O_749,N_14923,N_14929);
or UO_750 (O_750,N_14939,N_14919);
and UO_751 (O_751,N_14893,N_14967);
nand UO_752 (O_752,N_14904,N_14940);
nand UO_753 (O_753,N_14919,N_14995);
xor UO_754 (O_754,N_14922,N_14926);
nor UO_755 (O_755,N_14993,N_14878);
nand UO_756 (O_756,N_14952,N_14925);
or UO_757 (O_757,N_14975,N_14958);
nand UO_758 (O_758,N_14906,N_14959);
xor UO_759 (O_759,N_14970,N_14982);
and UO_760 (O_760,N_14946,N_14997);
xor UO_761 (O_761,N_14892,N_14954);
xor UO_762 (O_762,N_14895,N_14969);
nor UO_763 (O_763,N_14992,N_14911);
nand UO_764 (O_764,N_14984,N_14885);
and UO_765 (O_765,N_14998,N_14990);
and UO_766 (O_766,N_14985,N_14935);
and UO_767 (O_767,N_14974,N_14979);
or UO_768 (O_768,N_14950,N_14922);
or UO_769 (O_769,N_14990,N_14876);
nand UO_770 (O_770,N_14977,N_14972);
and UO_771 (O_771,N_14926,N_14892);
or UO_772 (O_772,N_14921,N_14945);
and UO_773 (O_773,N_14945,N_14938);
or UO_774 (O_774,N_14973,N_14909);
and UO_775 (O_775,N_14917,N_14918);
and UO_776 (O_776,N_14883,N_14972);
or UO_777 (O_777,N_14904,N_14928);
nor UO_778 (O_778,N_14900,N_14885);
xor UO_779 (O_779,N_14954,N_14950);
and UO_780 (O_780,N_14970,N_14918);
and UO_781 (O_781,N_14907,N_14978);
xnor UO_782 (O_782,N_14882,N_14921);
nand UO_783 (O_783,N_14957,N_14902);
nand UO_784 (O_784,N_14958,N_14985);
nand UO_785 (O_785,N_14996,N_14911);
nand UO_786 (O_786,N_14911,N_14917);
nand UO_787 (O_787,N_14946,N_14972);
or UO_788 (O_788,N_14887,N_14878);
nor UO_789 (O_789,N_14925,N_14898);
or UO_790 (O_790,N_14885,N_14894);
xor UO_791 (O_791,N_14891,N_14887);
and UO_792 (O_792,N_14961,N_14880);
nand UO_793 (O_793,N_14893,N_14892);
or UO_794 (O_794,N_14963,N_14942);
xor UO_795 (O_795,N_14989,N_14962);
or UO_796 (O_796,N_14939,N_14932);
nand UO_797 (O_797,N_14905,N_14936);
nand UO_798 (O_798,N_14999,N_14947);
nor UO_799 (O_799,N_14965,N_14891);
nand UO_800 (O_800,N_14994,N_14901);
xor UO_801 (O_801,N_14893,N_14943);
nand UO_802 (O_802,N_14983,N_14966);
or UO_803 (O_803,N_14936,N_14897);
nor UO_804 (O_804,N_14957,N_14918);
nor UO_805 (O_805,N_14934,N_14965);
xnor UO_806 (O_806,N_14899,N_14898);
and UO_807 (O_807,N_14883,N_14914);
nand UO_808 (O_808,N_14963,N_14880);
nor UO_809 (O_809,N_14965,N_14905);
nor UO_810 (O_810,N_14980,N_14934);
xor UO_811 (O_811,N_14909,N_14903);
nor UO_812 (O_812,N_14969,N_14954);
xnor UO_813 (O_813,N_14987,N_14905);
nand UO_814 (O_814,N_14907,N_14953);
or UO_815 (O_815,N_14898,N_14947);
nand UO_816 (O_816,N_14913,N_14916);
or UO_817 (O_817,N_14959,N_14886);
nand UO_818 (O_818,N_14998,N_14910);
xnor UO_819 (O_819,N_14929,N_14967);
nand UO_820 (O_820,N_14922,N_14876);
or UO_821 (O_821,N_14929,N_14904);
or UO_822 (O_822,N_14898,N_14927);
nor UO_823 (O_823,N_14979,N_14876);
xor UO_824 (O_824,N_14906,N_14991);
and UO_825 (O_825,N_14922,N_14998);
or UO_826 (O_826,N_14881,N_14882);
nand UO_827 (O_827,N_14954,N_14953);
and UO_828 (O_828,N_14908,N_14999);
and UO_829 (O_829,N_14889,N_14970);
xor UO_830 (O_830,N_14923,N_14892);
xor UO_831 (O_831,N_14992,N_14902);
xnor UO_832 (O_832,N_14939,N_14878);
xnor UO_833 (O_833,N_14950,N_14875);
xor UO_834 (O_834,N_14925,N_14978);
or UO_835 (O_835,N_14896,N_14890);
and UO_836 (O_836,N_14879,N_14992);
nor UO_837 (O_837,N_14967,N_14878);
and UO_838 (O_838,N_14991,N_14964);
and UO_839 (O_839,N_14985,N_14970);
nand UO_840 (O_840,N_14936,N_14901);
nor UO_841 (O_841,N_14949,N_14965);
nor UO_842 (O_842,N_14886,N_14881);
nand UO_843 (O_843,N_14939,N_14957);
or UO_844 (O_844,N_14932,N_14948);
and UO_845 (O_845,N_14916,N_14898);
and UO_846 (O_846,N_14971,N_14965);
xor UO_847 (O_847,N_14990,N_14977);
nor UO_848 (O_848,N_14978,N_14962);
or UO_849 (O_849,N_14976,N_14977);
xnor UO_850 (O_850,N_14977,N_14957);
and UO_851 (O_851,N_14979,N_14884);
and UO_852 (O_852,N_14881,N_14888);
nand UO_853 (O_853,N_14911,N_14938);
xor UO_854 (O_854,N_14908,N_14954);
nor UO_855 (O_855,N_14906,N_14923);
and UO_856 (O_856,N_14940,N_14936);
and UO_857 (O_857,N_14948,N_14984);
and UO_858 (O_858,N_14998,N_14887);
or UO_859 (O_859,N_14875,N_14929);
and UO_860 (O_860,N_14887,N_14892);
nor UO_861 (O_861,N_14875,N_14895);
nand UO_862 (O_862,N_14998,N_14987);
or UO_863 (O_863,N_14923,N_14936);
xnor UO_864 (O_864,N_14960,N_14931);
xnor UO_865 (O_865,N_14971,N_14912);
or UO_866 (O_866,N_14991,N_14896);
and UO_867 (O_867,N_14973,N_14893);
nand UO_868 (O_868,N_14897,N_14971);
xor UO_869 (O_869,N_14919,N_14914);
xnor UO_870 (O_870,N_14999,N_14894);
xnor UO_871 (O_871,N_14885,N_14915);
or UO_872 (O_872,N_14936,N_14966);
nand UO_873 (O_873,N_14957,N_14971);
and UO_874 (O_874,N_14908,N_14971);
or UO_875 (O_875,N_14910,N_14900);
or UO_876 (O_876,N_14897,N_14989);
nor UO_877 (O_877,N_14899,N_14970);
xor UO_878 (O_878,N_14910,N_14985);
nor UO_879 (O_879,N_14938,N_14887);
nor UO_880 (O_880,N_14906,N_14915);
or UO_881 (O_881,N_14890,N_14888);
or UO_882 (O_882,N_14981,N_14995);
and UO_883 (O_883,N_14932,N_14983);
or UO_884 (O_884,N_14944,N_14988);
nand UO_885 (O_885,N_14977,N_14907);
xor UO_886 (O_886,N_14890,N_14942);
or UO_887 (O_887,N_14919,N_14996);
nand UO_888 (O_888,N_14959,N_14938);
xnor UO_889 (O_889,N_14994,N_14917);
and UO_890 (O_890,N_14989,N_14875);
and UO_891 (O_891,N_14997,N_14906);
or UO_892 (O_892,N_14921,N_14905);
nor UO_893 (O_893,N_14995,N_14909);
nand UO_894 (O_894,N_14973,N_14912);
or UO_895 (O_895,N_14886,N_14925);
and UO_896 (O_896,N_14916,N_14914);
or UO_897 (O_897,N_14954,N_14936);
or UO_898 (O_898,N_14950,N_14972);
xnor UO_899 (O_899,N_14991,N_14994);
nand UO_900 (O_900,N_14991,N_14979);
xor UO_901 (O_901,N_14986,N_14961);
xnor UO_902 (O_902,N_14950,N_14984);
xor UO_903 (O_903,N_14975,N_14935);
nand UO_904 (O_904,N_14942,N_14940);
nand UO_905 (O_905,N_14923,N_14940);
and UO_906 (O_906,N_14894,N_14928);
xnor UO_907 (O_907,N_14890,N_14937);
or UO_908 (O_908,N_14875,N_14886);
or UO_909 (O_909,N_14875,N_14949);
nand UO_910 (O_910,N_14990,N_14999);
or UO_911 (O_911,N_14993,N_14899);
xnor UO_912 (O_912,N_14881,N_14877);
and UO_913 (O_913,N_14972,N_14935);
and UO_914 (O_914,N_14959,N_14944);
xnor UO_915 (O_915,N_14901,N_14903);
and UO_916 (O_916,N_14924,N_14875);
xnor UO_917 (O_917,N_14884,N_14913);
nor UO_918 (O_918,N_14983,N_14920);
nor UO_919 (O_919,N_14983,N_14889);
nand UO_920 (O_920,N_14891,N_14928);
nand UO_921 (O_921,N_14932,N_14905);
xor UO_922 (O_922,N_14973,N_14966);
nand UO_923 (O_923,N_14964,N_14969);
nand UO_924 (O_924,N_14933,N_14915);
or UO_925 (O_925,N_14944,N_14949);
nand UO_926 (O_926,N_14954,N_14975);
or UO_927 (O_927,N_14941,N_14991);
and UO_928 (O_928,N_14930,N_14987);
nor UO_929 (O_929,N_14904,N_14924);
nand UO_930 (O_930,N_14939,N_14933);
xor UO_931 (O_931,N_14920,N_14886);
nor UO_932 (O_932,N_14877,N_14975);
nor UO_933 (O_933,N_14993,N_14877);
nor UO_934 (O_934,N_14902,N_14908);
nand UO_935 (O_935,N_14985,N_14942);
nand UO_936 (O_936,N_14954,N_14897);
xor UO_937 (O_937,N_14891,N_14959);
nand UO_938 (O_938,N_14905,N_14914);
or UO_939 (O_939,N_14967,N_14877);
nand UO_940 (O_940,N_14936,N_14875);
nand UO_941 (O_941,N_14991,N_14887);
or UO_942 (O_942,N_14949,N_14902);
or UO_943 (O_943,N_14985,N_14941);
nand UO_944 (O_944,N_14986,N_14907);
nor UO_945 (O_945,N_14940,N_14943);
and UO_946 (O_946,N_14895,N_14904);
nand UO_947 (O_947,N_14966,N_14947);
or UO_948 (O_948,N_14885,N_14918);
xor UO_949 (O_949,N_14938,N_14900);
and UO_950 (O_950,N_14938,N_14943);
or UO_951 (O_951,N_14988,N_14984);
nor UO_952 (O_952,N_14999,N_14876);
and UO_953 (O_953,N_14938,N_14889);
nand UO_954 (O_954,N_14890,N_14880);
or UO_955 (O_955,N_14940,N_14963);
xor UO_956 (O_956,N_14900,N_14953);
and UO_957 (O_957,N_14935,N_14919);
and UO_958 (O_958,N_14946,N_14896);
nor UO_959 (O_959,N_14932,N_14899);
and UO_960 (O_960,N_14914,N_14996);
nand UO_961 (O_961,N_14951,N_14925);
nor UO_962 (O_962,N_14895,N_14931);
nor UO_963 (O_963,N_14965,N_14990);
or UO_964 (O_964,N_14975,N_14971);
and UO_965 (O_965,N_14892,N_14971);
xnor UO_966 (O_966,N_14917,N_14966);
xor UO_967 (O_967,N_14995,N_14964);
xnor UO_968 (O_968,N_14951,N_14942);
and UO_969 (O_969,N_14950,N_14947);
nor UO_970 (O_970,N_14889,N_14987);
nor UO_971 (O_971,N_14943,N_14952);
and UO_972 (O_972,N_14932,N_14981);
and UO_973 (O_973,N_14887,N_14877);
nor UO_974 (O_974,N_14930,N_14973);
nor UO_975 (O_975,N_14941,N_14965);
or UO_976 (O_976,N_14999,N_14934);
xnor UO_977 (O_977,N_14987,N_14959);
nand UO_978 (O_978,N_14886,N_14894);
or UO_979 (O_979,N_14938,N_14880);
nand UO_980 (O_980,N_14909,N_14881);
or UO_981 (O_981,N_14946,N_14950);
or UO_982 (O_982,N_14937,N_14952);
xor UO_983 (O_983,N_14897,N_14912);
nand UO_984 (O_984,N_14896,N_14891);
and UO_985 (O_985,N_14919,N_14982);
or UO_986 (O_986,N_14925,N_14959);
nor UO_987 (O_987,N_14885,N_14919);
and UO_988 (O_988,N_14979,N_14895);
xor UO_989 (O_989,N_14988,N_14892);
nand UO_990 (O_990,N_14915,N_14976);
nor UO_991 (O_991,N_14927,N_14955);
xor UO_992 (O_992,N_14992,N_14892);
nand UO_993 (O_993,N_14976,N_14938);
xnor UO_994 (O_994,N_14964,N_14897);
nand UO_995 (O_995,N_14983,N_14909);
xnor UO_996 (O_996,N_14908,N_14875);
and UO_997 (O_997,N_14966,N_14881);
xor UO_998 (O_998,N_14937,N_14961);
nor UO_999 (O_999,N_14944,N_14992);
and UO_1000 (O_1000,N_14947,N_14935);
nor UO_1001 (O_1001,N_14944,N_14976);
or UO_1002 (O_1002,N_14945,N_14880);
and UO_1003 (O_1003,N_14996,N_14937);
xnor UO_1004 (O_1004,N_14932,N_14908);
nor UO_1005 (O_1005,N_14877,N_14926);
xnor UO_1006 (O_1006,N_14956,N_14966);
and UO_1007 (O_1007,N_14888,N_14939);
nand UO_1008 (O_1008,N_14877,N_14919);
or UO_1009 (O_1009,N_14928,N_14944);
and UO_1010 (O_1010,N_14971,N_14966);
xnor UO_1011 (O_1011,N_14982,N_14908);
nand UO_1012 (O_1012,N_14940,N_14884);
xnor UO_1013 (O_1013,N_14923,N_14916);
nor UO_1014 (O_1014,N_14893,N_14997);
nand UO_1015 (O_1015,N_14973,N_14986);
and UO_1016 (O_1016,N_14879,N_14917);
nor UO_1017 (O_1017,N_14967,N_14882);
or UO_1018 (O_1018,N_14962,N_14944);
nor UO_1019 (O_1019,N_14979,N_14967);
and UO_1020 (O_1020,N_14978,N_14942);
xnor UO_1021 (O_1021,N_14932,N_14882);
and UO_1022 (O_1022,N_14959,N_14940);
and UO_1023 (O_1023,N_14884,N_14898);
nor UO_1024 (O_1024,N_14937,N_14904);
xor UO_1025 (O_1025,N_14882,N_14924);
and UO_1026 (O_1026,N_14951,N_14944);
nor UO_1027 (O_1027,N_14956,N_14955);
nor UO_1028 (O_1028,N_14878,N_14935);
nand UO_1029 (O_1029,N_14876,N_14996);
and UO_1030 (O_1030,N_14928,N_14986);
xor UO_1031 (O_1031,N_14963,N_14993);
nand UO_1032 (O_1032,N_14906,N_14907);
and UO_1033 (O_1033,N_14934,N_14936);
or UO_1034 (O_1034,N_14972,N_14886);
nand UO_1035 (O_1035,N_14923,N_14924);
xor UO_1036 (O_1036,N_14992,N_14998);
nand UO_1037 (O_1037,N_14878,N_14908);
or UO_1038 (O_1038,N_14933,N_14892);
nand UO_1039 (O_1039,N_14996,N_14978);
or UO_1040 (O_1040,N_14972,N_14934);
xor UO_1041 (O_1041,N_14919,N_14913);
or UO_1042 (O_1042,N_14948,N_14968);
xor UO_1043 (O_1043,N_14922,N_14894);
nor UO_1044 (O_1044,N_14900,N_14967);
xor UO_1045 (O_1045,N_14888,N_14917);
or UO_1046 (O_1046,N_14909,N_14924);
xnor UO_1047 (O_1047,N_14902,N_14888);
and UO_1048 (O_1048,N_14963,N_14980);
and UO_1049 (O_1049,N_14913,N_14933);
nand UO_1050 (O_1050,N_14946,N_14969);
and UO_1051 (O_1051,N_14878,N_14925);
nor UO_1052 (O_1052,N_14981,N_14890);
nand UO_1053 (O_1053,N_14890,N_14899);
nand UO_1054 (O_1054,N_14948,N_14977);
and UO_1055 (O_1055,N_14913,N_14951);
nand UO_1056 (O_1056,N_14891,N_14951);
xnor UO_1057 (O_1057,N_14907,N_14939);
xor UO_1058 (O_1058,N_14953,N_14985);
and UO_1059 (O_1059,N_14992,N_14936);
and UO_1060 (O_1060,N_14998,N_14965);
nor UO_1061 (O_1061,N_14978,N_14972);
nor UO_1062 (O_1062,N_14894,N_14899);
xnor UO_1063 (O_1063,N_14946,N_14962);
xor UO_1064 (O_1064,N_14921,N_14908);
xor UO_1065 (O_1065,N_14967,N_14920);
nand UO_1066 (O_1066,N_14983,N_14941);
xnor UO_1067 (O_1067,N_14980,N_14982);
and UO_1068 (O_1068,N_14962,N_14979);
and UO_1069 (O_1069,N_14934,N_14967);
nor UO_1070 (O_1070,N_14984,N_14960);
nor UO_1071 (O_1071,N_14994,N_14914);
nor UO_1072 (O_1072,N_14952,N_14965);
xnor UO_1073 (O_1073,N_14984,N_14923);
or UO_1074 (O_1074,N_14955,N_14878);
and UO_1075 (O_1075,N_14916,N_14955);
nand UO_1076 (O_1076,N_14976,N_14932);
and UO_1077 (O_1077,N_14996,N_14879);
or UO_1078 (O_1078,N_14989,N_14999);
or UO_1079 (O_1079,N_14988,N_14947);
or UO_1080 (O_1080,N_14878,N_14969);
nor UO_1081 (O_1081,N_14933,N_14883);
or UO_1082 (O_1082,N_14923,N_14945);
or UO_1083 (O_1083,N_14965,N_14919);
and UO_1084 (O_1084,N_14987,N_14890);
nor UO_1085 (O_1085,N_14972,N_14966);
or UO_1086 (O_1086,N_14992,N_14982);
and UO_1087 (O_1087,N_14932,N_14992);
nor UO_1088 (O_1088,N_14877,N_14902);
nor UO_1089 (O_1089,N_14934,N_14930);
and UO_1090 (O_1090,N_14880,N_14949);
and UO_1091 (O_1091,N_14986,N_14935);
and UO_1092 (O_1092,N_14935,N_14907);
xnor UO_1093 (O_1093,N_14922,N_14918);
xnor UO_1094 (O_1094,N_14896,N_14926);
nand UO_1095 (O_1095,N_14985,N_14887);
or UO_1096 (O_1096,N_14884,N_14925);
xnor UO_1097 (O_1097,N_14922,N_14972);
nand UO_1098 (O_1098,N_14963,N_14971);
nand UO_1099 (O_1099,N_14979,N_14882);
nand UO_1100 (O_1100,N_14953,N_14962);
nor UO_1101 (O_1101,N_14875,N_14915);
nor UO_1102 (O_1102,N_14898,N_14950);
xnor UO_1103 (O_1103,N_14888,N_14915);
or UO_1104 (O_1104,N_14950,N_14891);
nand UO_1105 (O_1105,N_14942,N_14897);
nand UO_1106 (O_1106,N_14917,N_14910);
nand UO_1107 (O_1107,N_14969,N_14994);
xor UO_1108 (O_1108,N_14877,N_14994);
or UO_1109 (O_1109,N_14902,N_14907);
nand UO_1110 (O_1110,N_14916,N_14959);
xnor UO_1111 (O_1111,N_14950,N_14965);
and UO_1112 (O_1112,N_14998,N_14924);
nand UO_1113 (O_1113,N_14916,N_14994);
nor UO_1114 (O_1114,N_14947,N_14892);
nand UO_1115 (O_1115,N_14969,N_14893);
xor UO_1116 (O_1116,N_14953,N_14958);
nor UO_1117 (O_1117,N_14907,N_14880);
xor UO_1118 (O_1118,N_14928,N_14949);
nor UO_1119 (O_1119,N_14930,N_14884);
and UO_1120 (O_1120,N_14948,N_14944);
nand UO_1121 (O_1121,N_14885,N_14935);
and UO_1122 (O_1122,N_14875,N_14967);
and UO_1123 (O_1123,N_14884,N_14876);
nand UO_1124 (O_1124,N_14879,N_14979);
xnor UO_1125 (O_1125,N_14928,N_14936);
xor UO_1126 (O_1126,N_14964,N_14888);
and UO_1127 (O_1127,N_14983,N_14895);
nand UO_1128 (O_1128,N_14904,N_14912);
xor UO_1129 (O_1129,N_14915,N_14878);
or UO_1130 (O_1130,N_14992,N_14931);
xnor UO_1131 (O_1131,N_14962,N_14897);
or UO_1132 (O_1132,N_14998,N_14900);
nand UO_1133 (O_1133,N_14908,N_14882);
and UO_1134 (O_1134,N_14934,N_14895);
and UO_1135 (O_1135,N_14900,N_14980);
xor UO_1136 (O_1136,N_14882,N_14990);
nand UO_1137 (O_1137,N_14881,N_14907);
xnor UO_1138 (O_1138,N_14879,N_14967);
nor UO_1139 (O_1139,N_14928,N_14886);
or UO_1140 (O_1140,N_14908,N_14901);
nand UO_1141 (O_1141,N_14914,N_14898);
nand UO_1142 (O_1142,N_14973,N_14928);
nand UO_1143 (O_1143,N_14892,N_14996);
xnor UO_1144 (O_1144,N_14895,N_14919);
nand UO_1145 (O_1145,N_14996,N_14877);
and UO_1146 (O_1146,N_14979,N_14888);
or UO_1147 (O_1147,N_14884,N_14888);
nand UO_1148 (O_1148,N_14993,N_14901);
nor UO_1149 (O_1149,N_14877,N_14989);
xor UO_1150 (O_1150,N_14888,N_14929);
nand UO_1151 (O_1151,N_14995,N_14924);
or UO_1152 (O_1152,N_14889,N_14908);
and UO_1153 (O_1153,N_14968,N_14999);
nor UO_1154 (O_1154,N_14950,N_14892);
or UO_1155 (O_1155,N_14931,N_14938);
and UO_1156 (O_1156,N_14968,N_14939);
or UO_1157 (O_1157,N_14982,N_14954);
nor UO_1158 (O_1158,N_14953,N_14991);
xnor UO_1159 (O_1159,N_14917,N_14958);
nor UO_1160 (O_1160,N_14923,N_14939);
nor UO_1161 (O_1161,N_14894,N_14953);
and UO_1162 (O_1162,N_14980,N_14971);
or UO_1163 (O_1163,N_14878,N_14930);
and UO_1164 (O_1164,N_14933,N_14989);
nand UO_1165 (O_1165,N_14965,N_14963);
xnor UO_1166 (O_1166,N_14999,N_14881);
xnor UO_1167 (O_1167,N_14892,N_14976);
nand UO_1168 (O_1168,N_14920,N_14919);
nand UO_1169 (O_1169,N_14904,N_14997);
or UO_1170 (O_1170,N_14976,N_14910);
or UO_1171 (O_1171,N_14953,N_14924);
or UO_1172 (O_1172,N_14876,N_14887);
or UO_1173 (O_1173,N_14944,N_14963);
or UO_1174 (O_1174,N_14976,N_14964);
and UO_1175 (O_1175,N_14889,N_14930);
nor UO_1176 (O_1176,N_14965,N_14908);
or UO_1177 (O_1177,N_14879,N_14965);
nand UO_1178 (O_1178,N_14914,N_14938);
and UO_1179 (O_1179,N_14886,N_14993);
or UO_1180 (O_1180,N_14959,N_14945);
or UO_1181 (O_1181,N_14960,N_14875);
nor UO_1182 (O_1182,N_14982,N_14909);
or UO_1183 (O_1183,N_14905,N_14960);
nor UO_1184 (O_1184,N_14914,N_14992);
nand UO_1185 (O_1185,N_14915,N_14934);
or UO_1186 (O_1186,N_14962,N_14952);
nor UO_1187 (O_1187,N_14934,N_14901);
nor UO_1188 (O_1188,N_14951,N_14926);
nand UO_1189 (O_1189,N_14893,N_14921);
and UO_1190 (O_1190,N_14928,N_14998);
or UO_1191 (O_1191,N_14961,N_14998);
xnor UO_1192 (O_1192,N_14974,N_14925);
nand UO_1193 (O_1193,N_14981,N_14924);
nor UO_1194 (O_1194,N_14885,N_14975);
and UO_1195 (O_1195,N_14943,N_14950);
nor UO_1196 (O_1196,N_14904,N_14935);
or UO_1197 (O_1197,N_14948,N_14924);
or UO_1198 (O_1198,N_14892,N_14945);
nor UO_1199 (O_1199,N_14992,N_14937);
nor UO_1200 (O_1200,N_14956,N_14941);
nand UO_1201 (O_1201,N_14922,N_14902);
xor UO_1202 (O_1202,N_14909,N_14974);
xor UO_1203 (O_1203,N_14944,N_14888);
or UO_1204 (O_1204,N_14916,N_14910);
and UO_1205 (O_1205,N_14980,N_14916);
nand UO_1206 (O_1206,N_14960,N_14936);
xnor UO_1207 (O_1207,N_14978,N_14961);
xnor UO_1208 (O_1208,N_14918,N_14901);
or UO_1209 (O_1209,N_14896,N_14934);
or UO_1210 (O_1210,N_14946,N_14889);
and UO_1211 (O_1211,N_14988,N_14916);
or UO_1212 (O_1212,N_14971,N_14906);
xnor UO_1213 (O_1213,N_14983,N_14888);
xnor UO_1214 (O_1214,N_14877,N_14908);
and UO_1215 (O_1215,N_14948,N_14974);
xnor UO_1216 (O_1216,N_14970,N_14959);
or UO_1217 (O_1217,N_14886,N_14935);
nand UO_1218 (O_1218,N_14996,N_14967);
nor UO_1219 (O_1219,N_14974,N_14969);
nor UO_1220 (O_1220,N_14911,N_14978);
xnor UO_1221 (O_1221,N_14891,N_14889);
nor UO_1222 (O_1222,N_14945,N_14961);
xnor UO_1223 (O_1223,N_14930,N_14996);
nand UO_1224 (O_1224,N_14998,N_14982);
xor UO_1225 (O_1225,N_14940,N_14912);
or UO_1226 (O_1226,N_14969,N_14988);
nor UO_1227 (O_1227,N_14960,N_14982);
and UO_1228 (O_1228,N_14893,N_14927);
nand UO_1229 (O_1229,N_14934,N_14944);
xor UO_1230 (O_1230,N_14926,N_14930);
nand UO_1231 (O_1231,N_14926,N_14985);
nor UO_1232 (O_1232,N_14936,N_14989);
and UO_1233 (O_1233,N_14961,N_14916);
nor UO_1234 (O_1234,N_14916,N_14896);
and UO_1235 (O_1235,N_14914,N_14888);
and UO_1236 (O_1236,N_14888,N_14959);
xnor UO_1237 (O_1237,N_14945,N_14974);
xor UO_1238 (O_1238,N_14998,N_14950);
nand UO_1239 (O_1239,N_14941,N_14877);
nand UO_1240 (O_1240,N_14986,N_14939);
and UO_1241 (O_1241,N_14997,N_14927);
nor UO_1242 (O_1242,N_14978,N_14892);
nor UO_1243 (O_1243,N_14902,N_14910);
nor UO_1244 (O_1244,N_14918,N_14982);
xor UO_1245 (O_1245,N_14875,N_14945);
nor UO_1246 (O_1246,N_14939,N_14982);
or UO_1247 (O_1247,N_14969,N_14920);
and UO_1248 (O_1248,N_14899,N_14934);
xor UO_1249 (O_1249,N_14993,N_14967);
nand UO_1250 (O_1250,N_14921,N_14987);
or UO_1251 (O_1251,N_14898,N_14980);
and UO_1252 (O_1252,N_14911,N_14975);
xor UO_1253 (O_1253,N_14881,N_14939);
nand UO_1254 (O_1254,N_14951,N_14916);
nand UO_1255 (O_1255,N_14979,N_14912);
xnor UO_1256 (O_1256,N_14957,N_14893);
xor UO_1257 (O_1257,N_14919,N_14896);
and UO_1258 (O_1258,N_14991,N_14951);
nand UO_1259 (O_1259,N_14972,N_14898);
nor UO_1260 (O_1260,N_14879,N_14955);
nand UO_1261 (O_1261,N_14970,N_14953);
nand UO_1262 (O_1262,N_14976,N_14931);
nor UO_1263 (O_1263,N_14907,N_14916);
and UO_1264 (O_1264,N_14998,N_14973);
nor UO_1265 (O_1265,N_14978,N_14987);
and UO_1266 (O_1266,N_14878,N_14920);
and UO_1267 (O_1267,N_14892,N_14935);
nor UO_1268 (O_1268,N_14927,N_14911);
and UO_1269 (O_1269,N_14914,N_14997);
nand UO_1270 (O_1270,N_14965,N_14890);
nand UO_1271 (O_1271,N_14908,N_14888);
xor UO_1272 (O_1272,N_14976,N_14961);
or UO_1273 (O_1273,N_14971,N_14934);
nor UO_1274 (O_1274,N_14998,N_14875);
nand UO_1275 (O_1275,N_14984,N_14971);
and UO_1276 (O_1276,N_14936,N_14912);
and UO_1277 (O_1277,N_14983,N_14942);
and UO_1278 (O_1278,N_14918,N_14876);
nor UO_1279 (O_1279,N_14875,N_14988);
xnor UO_1280 (O_1280,N_14911,N_14994);
nor UO_1281 (O_1281,N_14888,N_14992);
nor UO_1282 (O_1282,N_14987,N_14968);
and UO_1283 (O_1283,N_14947,N_14928);
and UO_1284 (O_1284,N_14939,N_14913);
or UO_1285 (O_1285,N_14890,N_14945);
nor UO_1286 (O_1286,N_14968,N_14929);
and UO_1287 (O_1287,N_14893,N_14911);
nor UO_1288 (O_1288,N_14964,N_14904);
nor UO_1289 (O_1289,N_14966,N_14999);
and UO_1290 (O_1290,N_14963,N_14923);
nand UO_1291 (O_1291,N_14895,N_14975);
and UO_1292 (O_1292,N_14957,N_14941);
nor UO_1293 (O_1293,N_14886,N_14888);
or UO_1294 (O_1294,N_14906,N_14976);
nand UO_1295 (O_1295,N_14930,N_14908);
nand UO_1296 (O_1296,N_14878,N_14959);
or UO_1297 (O_1297,N_14925,N_14920);
and UO_1298 (O_1298,N_14958,N_14896);
xnor UO_1299 (O_1299,N_14889,N_14949);
nand UO_1300 (O_1300,N_14979,N_14976);
and UO_1301 (O_1301,N_14995,N_14977);
xnor UO_1302 (O_1302,N_14921,N_14967);
nand UO_1303 (O_1303,N_14971,N_14954);
xor UO_1304 (O_1304,N_14971,N_14899);
or UO_1305 (O_1305,N_14949,N_14987);
nor UO_1306 (O_1306,N_14939,N_14930);
and UO_1307 (O_1307,N_14911,N_14894);
and UO_1308 (O_1308,N_14886,N_14906);
nand UO_1309 (O_1309,N_14966,N_14895);
nand UO_1310 (O_1310,N_14877,N_14951);
or UO_1311 (O_1311,N_14881,N_14879);
or UO_1312 (O_1312,N_14961,N_14999);
nand UO_1313 (O_1313,N_14903,N_14960);
and UO_1314 (O_1314,N_14964,N_14894);
nor UO_1315 (O_1315,N_14951,N_14882);
xor UO_1316 (O_1316,N_14946,N_14960);
nor UO_1317 (O_1317,N_14901,N_14953);
nand UO_1318 (O_1318,N_14922,N_14923);
nor UO_1319 (O_1319,N_14916,N_14880);
and UO_1320 (O_1320,N_14985,N_14882);
xnor UO_1321 (O_1321,N_14960,N_14948);
and UO_1322 (O_1322,N_14994,N_14905);
nand UO_1323 (O_1323,N_14905,N_14975);
and UO_1324 (O_1324,N_14905,N_14884);
and UO_1325 (O_1325,N_14879,N_14901);
nor UO_1326 (O_1326,N_14956,N_14920);
and UO_1327 (O_1327,N_14888,N_14887);
nor UO_1328 (O_1328,N_14926,N_14931);
and UO_1329 (O_1329,N_14920,N_14944);
and UO_1330 (O_1330,N_14896,N_14901);
xnor UO_1331 (O_1331,N_14981,N_14953);
nor UO_1332 (O_1332,N_14930,N_14948);
nor UO_1333 (O_1333,N_14973,N_14890);
xnor UO_1334 (O_1334,N_14899,N_14975);
nand UO_1335 (O_1335,N_14991,N_14891);
nor UO_1336 (O_1336,N_14980,N_14990);
and UO_1337 (O_1337,N_14904,N_14962);
nand UO_1338 (O_1338,N_14893,N_14918);
nor UO_1339 (O_1339,N_14965,N_14942);
and UO_1340 (O_1340,N_14908,N_14924);
nor UO_1341 (O_1341,N_14902,N_14977);
nor UO_1342 (O_1342,N_14953,N_14921);
and UO_1343 (O_1343,N_14889,N_14953);
and UO_1344 (O_1344,N_14938,N_14895);
and UO_1345 (O_1345,N_14995,N_14943);
xor UO_1346 (O_1346,N_14999,N_14901);
nand UO_1347 (O_1347,N_14904,N_14901);
or UO_1348 (O_1348,N_14950,N_14916);
and UO_1349 (O_1349,N_14958,N_14904);
xnor UO_1350 (O_1350,N_14934,N_14928);
or UO_1351 (O_1351,N_14916,N_14893);
xor UO_1352 (O_1352,N_14971,N_14968);
nor UO_1353 (O_1353,N_14957,N_14981);
or UO_1354 (O_1354,N_14911,N_14910);
or UO_1355 (O_1355,N_14936,N_14971);
xor UO_1356 (O_1356,N_14897,N_14958);
nor UO_1357 (O_1357,N_14940,N_14915);
xor UO_1358 (O_1358,N_14926,N_14995);
and UO_1359 (O_1359,N_14883,N_14928);
or UO_1360 (O_1360,N_14972,N_14916);
nand UO_1361 (O_1361,N_14939,N_14885);
or UO_1362 (O_1362,N_14925,N_14875);
nand UO_1363 (O_1363,N_14934,N_14997);
nor UO_1364 (O_1364,N_14974,N_14977);
and UO_1365 (O_1365,N_14975,N_14938);
nand UO_1366 (O_1366,N_14994,N_14972);
nor UO_1367 (O_1367,N_14939,N_14927);
or UO_1368 (O_1368,N_14983,N_14962);
xor UO_1369 (O_1369,N_14953,N_14914);
and UO_1370 (O_1370,N_14933,N_14917);
xor UO_1371 (O_1371,N_14978,N_14910);
and UO_1372 (O_1372,N_14952,N_14976);
nand UO_1373 (O_1373,N_14932,N_14930);
or UO_1374 (O_1374,N_14954,N_14922);
nand UO_1375 (O_1375,N_14880,N_14901);
or UO_1376 (O_1376,N_14911,N_14935);
nor UO_1377 (O_1377,N_14906,N_14894);
nor UO_1378 (O_1378,N_14993,N_14975);
xor UO_1379 (O_1379,N_14938,N_14988);
and UO_1380 (O_1380,N_14876,N_14913);
or UO_1381 (O_1381,N_14988,N_14912);
xnor UO_1382 (O_1382,N_14973,N_14971);
xnor UO_1383 (O_1383,N_14894,N_14907);
nand UO_1384 (O_1384,N_14888,N_14968);
nor UO_1385 (O_1385,N_14957,N_14912);
and UO_1386 (O_1386,N_14909,N_14875);
nor UO_1387 (O_1387,N_14973,N_14960);
nand UO_1388 (O_1388,N_14935,N_14875);
nor UO_1389 (O_1389,N_14927,N_14974);
or UO_1390 (O_1390,N_14910,N_14896);
xor UO_1391 (O_1391,N_14901,N_14984);
nand UO_1392 (O_1392,N_14913,N_14980);
nor UO_1393 (O_1393,N_14996,N_14988);
xor UO_1394 (O_1394,N_14907,N_14901);
nor UO_1395 (O_1395,N_14960,N_14987);
nor UO_1396 (O_1396,N_14945,N_14876);
and UO_1397 (O_1397,N_14905,N_14885);
nor UO_1398 (O_1398,N_14982,N_14890);
or UO_1399 (O_1399,N_14940,N_14988);
xnor UO_1400 (O_1400,N_14882,N_14937);
nand UO_1401 (O_1401,N_14947,N_14983);
nand UO_1402 (O_1402,N_14900,N_14892);
nand UO_1403 (O_1403,N_14944,N_14986);
nor UO_1404 (O_1404,N_14994,N_14951);
or UO_1405 (O_1405,N_14910,N_14888);
or UO_1406 (O_1406,N_14937,N_14916);
xor UO_1407 (O_1407,N_14930,N_14901);
nand UO_1408 (O_1408,N_14978,N_14973);
and UO_1409 (O_1409,N_14958,N_14996);
xnor UO_1410 (O_1410,N_14965,N_14876);
xor UO_1411 (O_1411,N_14880,N_14903);
and UO_1412 (O_1412,N_14978,N_14968);
and UO_1413 (O_1413,N_14960,N_14958);
and UO_1414 (O_1414,N_14877,N_14933);
nand UO_1415 (O_1415,N_14985,N_14916);
xnor UO_1416 (O_1416,N_14909,N_14925);
and UO_1417 (O_1417,N_14991,N_14954);
xnor UO_1418 (O_1418,N_14889,N_14887);
nor UO_1419 (O_1419,N_14976,N_14900);
nor UO_1420 (O_1420,N_14996,N_14949);
and UO_1421 (O_1421,N_14944,N_14989);
or UO_1422 (O_1422,N_14911,N_14986);
or UO_1423 (O_1423,N_14999,N_14949);
xnor UO_1424 (O_1424,N_14993,N_14920);
and UO_1425 (O_1425,N_14994,N_14945);
nand UO_1426 (O_1426,N_14938,N_14899);
and UO_1427 (O_1427,N_14967,N_14948);
nor UO_1428 (O_1428,N_14982,N_14949);
and UO_1429 (O_1429,N_14965,N_14992);
or UO_1430 (O_1430,N_14985,N_14982);
nor UO_1431 (O_1431,N_14937,N_14924);
or UO_1432 (O_1432,N_14952,N_14882);
and UO_1433 (O_1433,N_14921,N_14991);
nand UO_1434 (O_1434,N_14949,N_14989);
nand UO_1435 (O_1435,N_14878,N_14909);
nor UO_1436 (O_1436,N_14885,N_14978);
nand UO_1437 (O_1437,N_14912,N_14964);
xor UO_1438 (O_1438,N_14963,N_14947);
nor UO_1439 (O_1439,N_14895,N_14930);
or UO_1440 (O_1440,N_14896,N_14880);
and UO_1441 (O_1441,N_14958,N_14965);
xnor UO_1442 (O_1442,N_14931,N_14991);
or UO_1443 (O_1443,N_14988,N_14954);
nor UO_1444 (O_1444,N_14893,N_14914);
or UO_1445 (O_1445,N_14950,N_14933);
nand UO_1446 (O_1446,N_14986,N_14880);
nand UO_1447 (O_1447,N_14888,N_14960);
xnor UO_1448 (O_1448,N_14948,N_14954);
xnor UO_1449 (O_1449,N_14938,N_14903);
nand UO_1450 (O_1450,N_14984,N_14926);
and UO_1451 (O_1451,N_14926,N_14935);
and UO_1452 (O_1452,N_14913,N_14991);
and UO_1453 (O_1453,N_14932,N_14887);
and UO_1454 (O_1454,N_14876,N_14941);
xor UO_1455 (O_1455,N_14969,N_14889);
xnor UO_1456 (O_1456,N_14963,N_14996);
xor UO_1457 (O_1457,N_14925,N_14999);
and UO_1458 (O_1458,N_14973,N_14933);
nor UO_1459 (O_1459,N_14922,N_14934);
or UO_1460 (O_1460,N_14891,N_14921);
and UO_1461 (O_1461,N_14935,N_14987);
or UO_1462 (O_1462,N_14971,N_14890);
nor UO_1463 (O_1463,N_14909,N_14911);
nor UO_1464 (O_1464,N_14895,N_14888);
nand UO_1465 (O_1465,N_14876,N_14907);
xor UO_1466 (O_1466,N_14917,N_14987);
nand UO_1467 (O_1467,N_14893,N_14999);
nand UO_1468 (O_1468,N_14893,N_14922);
nand UO_1469 (O_1469,N_14956,N_14899);
nand UO_1470 (O_1470,N_14988,N_14974);
nand UO_1471 (O_1471,N_14938,N_14956);
nand UO_1472 (O_1472,N_14970,N_14920);
nand UO_1473 (O_1473,N_14939,N_14974);
nor UO_1474 (O_1474,N_14933,N_14929);
xnor UO_1475 (O_1475,N_14878,N_14883);
xor UO_1476 (O_1476,N_14995,N_14987);
and UO_1477 (O_1477,N_14918,N_14891);
and UO_1478 (O_1478,N_14994,N_14919);
and UO_1479 (O_1479,N_14931,N_14916);
and UO_1480 (O_1480,N_14905,N_14880);
nor UO_1481 (O_1481,N_14885,N_14991);
and UO_1482 (O_1482,N_14990,N_14895);
and UO_1483 (O_1483,N_14992,N_14916);
and UO_1484 (O_1484,N_14905,N_14954);
nand UO_1485 (O_1485,N_14991,N_14944);
nor UO_1486 (O_1486,N_14882,N_14922);
and UO_1487 (O_1487,N_14879,N_14924);
nor UO_1488 (O_1488,N_14965,N_14915);
and UO_1489 (O_1489,N_14952,N_14881);
or UO_1490 (O_1490,N_14964,N_14915);
xnor UO_1491 (O_1491,N_14962,N_14980);
or UO_1492 (O_1492,N_14884,N_14943);
xor UO_1493 (O_1493,N_14881,N_14933);
xor UO_1494 (O_1494,N_14887,N_14915);
nor UO_1495 (O_1495,N_14976,N_14886);
nor UO_1496 (O_1496,N_14947,N_14905);
and UO_1497 (O_1497,N_14912,N_14965);
or UO_1498 (O_1498,N_14922,N_14978);
or UO_1499 (O_1499,N_14996,N_14895);
xnor UO_1500 (O_1500,N_14975,N_14988);
and UO_1501 (O_1501,N_14898,N_14905);
nand UO_1502 (O_1502,N_14971,N_14964);
nand UO_1503 (O_1503,N_14978,N_14963);
xnor UO_1504 (O_1504,N_14919,N_14915);
xnor UO_1505 (O_1505,N_14889,N_14905);
nand UO_1506 (O_1506,N_14998,N_14898);
nor UO_1507 (O_1507,N_14959,N_14932);
nand UO_1508 (O_1508,N_14951,N_14885);
nor UO_1509 (O_1509,N_14953,N_14937);
and UO_1510 (O_1510,N_14877,N_14980);
nand UO_1511 (O_1511,N_14966,N_14912);
xor UO_1512 (O_1512,N_14955,N_14888);
nand UO_1513 (O_1513,N_14953,N_14891);
or UO_1514 (O_1514,N_14959,N_14877);
and UO_1515 (O_1515,N_14969,N_14876);
and UO_1516 (O_1516,N_14901,N_14988);
or UO_1517 (O_1517,N_14906,N_14964);
nor UO_1518 (O_1518,N_14979,N_14911);
or UO_1519 (O_1519,N_14912,N_14952);
nor UO_1520 (O_1520,N_14908,N_14969);
and UO_1521 (O_1521,N_14912,N_14894);
or UO_1522 (O_1522,N_14927,N_14950);
nor UO_1523 (O_1523,N_14936,N_14882);
xnor UO_1524 (O_1524,N_14955,N_14944);
nor UO_1525 (O_1525,N_14996,N_14987);
nor UO_1526 (O_1526,N_14952,N_14972);
and UO_1527 (O_1527,N_14970,N_14995);
or UO_1528 (O_1528,N_14944,N_14979);
nand UO_1529 (O_1529,N_14951,N_14905);
nand UO_1530 (O_1530,N_14957,N_14984);
nand UO_1531 (O_1531,N_14979,N_14993);
or UO_1532 (O_1532,N_14958,N_14931);
xor UO_1533 (O_1533,N_14878,N_14884);
or UO_1534 (O_1534,N_14944,N_14990);
and UO_1535 (O_1535,N_14915,N_14917);
and UO_1536 (O_1536,N_14950,N_14894);
xnor UO_1537 (O_1537,N_14908,N_14998);
nor UO_1538 (O_1538,N_14967,N_14957);
and UO_1539 (O_1539,N_14948,N_14883);
nand UO_1540 (O_1540,N_14920,N_14934);
nor UO_1541 (O_1541,N_14907,N_14895);
xor UO_1542 (O_1542,N_14995,N_14985);
or UO_1543 (O_1543,N_14914,N_14960);
and UO_1544 (O_1544,N_14936,N_14968);
and UO_1545 (O_1545,N_14979,N_14946);
xnor UO_1546 (O_1546,N_14908,N_14916);
xnor UO_1547 (O_1547,N_14920,N_14901);
xnor UO_1548 (O_1548,N_14967,N_14887);
and UO_1549 (O_1549,N_14962,N_14883);
and UO_1550 (O_1550,N_14896,N_14879);
or UO_1551 (O_1551,N_14939,N_14893);
or UO_1552 (O_1552,N_14929,N_14999);
or UO_1553 (O_1553,N_14879,N_14885);
xnor UO_1554 (O_1554,N_14972,N_14997);
xnor UO_1555 (O_1555,N_14965,N_14883);
nor UO_1556 (O_1556,N_14882,N_14995);
and UO_1557 (O_1557,N_14945,N_14895);
nor UO_1558 (O_1558,N_14924,N_14980);
xnor UO_1559 (O_1559,N_14975,N_14881);
and UO_1560 (O_1560,N_14971,N_14998);
or UO_1561 (O_1561,N_14996,N_14954);
and UO_1562 (O_1562,N_14931,N_14945);
and UO_1563 (O_1563,N_14938,N_14898);
nor UO_1564 (O_1564,N_14966,N_14962);
nor UO_1565 (O_1565,N_14886,N_14889);
and UO_1566 (O_1566,N_14992,N_14906);
nand UO_1567 (O_1567,N_14900,N_14889);
nand UO_1568 (O_1568,N_14924,N_14895);
or UO_1569 (O_1569,N_14957,N_14924);
nor UO_1570 (O_1570,N_14962,N_14955);
xor UO_1571 (O_1571,N_14915,N_14957);
nand UO_1572 (O_1572,N_14999,N_14900);
or UO_1573 (O_1573,N_14907,N_14887);
xor UO_1574 (O_1574,N_14940,N_14949);
and UO_1575 (O_1575,N_14991,N_14952);
xor UO_1576 (O_1576,N_14877,N_14997);
nor UO_1577 (O_1577,N_14990,N_14914);
nor UO_1578 (O_1578,N_14920,N_14973);
or UO_1579 (O_1579,N_14918,N_14968);
or UO_1580 (O_1580,N_14979,N_14951);
or UO_1581 (O_1581,N_14962,N_14975);
or UO_1582 (O_1582,N_14942,N_14894);
nor UO_1583 (O_1583,N_14897,N_14949);
nor UO_1584 (O_1584,N_14973,N_14905);
nor UO_1585 (O_1585,N_14927,N_14960);
or UO_1586 (O_1586,N_14976,N_14920);
or UO_1587 (O_1587,N_14959,N_14928);
and UO_1588 (O_1588,N_14884,N_14939);
nor UO_1589 (O_1589,N_14913,N_14921);
and UO_1590 (O_1590,N_14914,N_14917);
or UO_1591 (O_1591,N_14931,N_14998);
nor UO_1592 (O_1592,N_14969,N_14948);
nand UO_1593 (O_1593,N_14915,N_14977);
xnor UO_1594 (O_1594,N_14910,N_14898);
or UO_1595 (O_1595,N_14880,N_14977);
nor UO_1596 (O_1596,N_14896,N_14998);
xor UO_1597 (O_1597,N_14973,N_14898);
nor UO_1598 (O_1598,N_14958,N_14875);
nor UO_1599 (O_1599,N_14934,N_14889);
and UO_1600 (O_1600,N_14986,N_14875);
xor UO_1601 (O_1601,N_14954,N_14961);
nand UO_1602 (O_1602,N_14896,N_14878);
and UO_1603 (O_1603,N_14900,N_14920);
or UO_1604 (O_1604,N_14949,N_14893);
and UO_1605 (O_1605,N_14915,N_14947);
and UO_1606 (O_1606,N_14983,N_14915);
and UO_1607 (O_1607,N_14997,N_14926);
nand UO_1608 (O_1608,N_14935,N_14880);
xnor UO_1609 (O_1609,N_14935,N_14940);
or UO_1610 (O_1610,N_14988,N_14949);
nor UO_1611 (O_1611,N_14943,N_14899);
and UO_1612 (O_1612,N_14981,N_14976);
nor UO_1613 (O_1613,N_14972,N_14988);
and UO_1614 (O_1614,N_14908,N_14966);
xor UO_1615 (O_1615,N_14999,N_14939);
and UO_1616 (O_1616,N_14920,N_14927);
nand UO_1617 (O_1617,N_14901,N_14969);
nor UO_1618 (O_1618,N_14885,N_14908);
xnor UO_1619 (O_1619,N_14899,N_14915);
and UO_1620 (O_1620,N_14949,N_14894);
or UO_1621 (O_1621,N_14958,N_14934);
nand UO_1622 (O_1622,N_14898,N_14957);
xor UO_1623 (O_1623,N_14899,N_14888);
or UO_1624 (O_1624,N_14880,N_14919);
xnor UO_1625 (O_1625,N_14917,N_14901);
xor UO_1626 (O_1626,N_14991,N_14912);
nor UO_1627 (O_1627,N_14936,N_14894);
or UO_1628 (O_1628,N_14922,N_14959);
xnor UO_1629 (O_1629,N_14903,N_14898);
or UO_1630 (O_1630,N_14919,N_14899);
xnor UO_1631 (O_1631,N_14905,N_14878);
or UO_1632 (O_1632,N_14938,N_14961);
nand UO_1633 (O_1633,N_14997,N_14899);
nor UO_1634 (O_1634,N_14920,N_14916);
or UO_1635 (O_1635,N_14888,N_14963);
or UO_1636 (O_1636,N_14904,N_14952);
nor UO_1637 (O_1637,N_14987,N_14948);
or UO_1638 (O_1638,N_14906,N_14876);
nand UO_1639 (O_1639,N_14885,N_14959);
and UO_1640 (O_1640,N_14950,N_14902);
nor UO_1641 (O_1641,N_14948,N_14956);
or UO_1642 (O_1642,N_14894,N_14959);
xnor UO_1643 (O_1643,N_14920,N_14939);
or UO_1644 (O_1644,N_14898,N_14882);
xor UO_1645 (O_1645,N_14951,N_14938);
nor UO_1646 (O_1646,N_14915,N_14910);
nor UO_1647 (O_1647,N_14938,N_14924);
or UO_1648 (O_1648,N_14911,N_14880);
or UO_1649 (O_1649,N_14956,N_14978);
nand UO_1650 (O_1650,N_14899,N_14939);
nand UO_1651 (O_1651,N_14945,N_14937);
nand UO_1652 (O_1652,N_14945,N_14977);
nor UO_1653 (O_1653,N_14916,N_14974);
xor UO_1654 (O_1654,N_14902,N_14927);
nor UO_1655 (O_1655,N_14997,N_14955);
nor UO_1656 (O_1656,N_14939,N_14891);
nor UO_1657 (O_1657,N_14971,N_14893);
nor UO_1658 (O_1658,N_14955,N_14957);
nor UO_1659 (O_1659,N_14979,N_14987);
nand UO_1660 (O_1660,N_14918,N_14892);
nor UO_1661 (O_1661,N_14996,N_14990);
nor UO_1662 (O_1662,N_14915,N_14953);
and UO_1663 (O_1663,N_14953,N_14895);
nand UO_1664 (O_1664,N_14917,N_14993);
nand UO_1665 (O_1665,N_14927,N_14943);
or UO_1666 (O_1666,N_14981,N_14917);
xnor UO_1667 (O_1667,N_14978,N_14953);
nand UO_1668 (O_1668,N_14905,N_14922);
xor UO_1669 (O_1669,N_14902,N_14897);
nand UO_1670 (O_1670,N_14982,N_14930);
nand UO_1671 (O_1671,N_14988,N_14977);
nor UO_1672 (O_1672,N_14993,N_14998);
or UO_1673 (O_1673,N_14894,N_14975);
xor UO_1674 (O_1674,N_14880,N_14985);
and UO_1675 (O_1675,N_14937,N_14895);
nand UO_1676 (O_1676,N_14966,N_14913);
nor UO_1677 (O_1677,N_14979,N_14901);
xor UO_1678 (O_1678,N_14906,N_14878);
nor UO_1679 (O_1679,N_14986,N_14963);
xnor UO_1680 (O_1680,N_14894,N_14969);
or UO_1681 (O_1681,N_14975,N_14886);
and UO_1682 (O_1682,N_14987,N_14881);
or UO_1683 (O_1683,N_14958,N_14899);
or UO_1684 (O_1684,N_14901,N_14964);
nand UO_1685 (O_1685,N_14878,N_14963);
or UO_1686 (O_1686,N_14954,N_14987);
xnor UO_1687 (O_1687,N_14996,N_14890);
xor UO_1688 (O_1688,N_14950,N_14967);
xnor UO_1689 (O_1689,N_14913,N_14958);
nand UO_1690 (O_1690,N_14979,N_14915);
and UO_1691 (O_1691,N_14909,N_14965);
nand UO_1692 (O_1692,N_14875,N_14878);
and UO_1693 (O_1693,N_14877,N_14984);
xor UO_1694 (O_1694,N_14919,N_14978);
nor UO_1695 (O_1695,N_14921,N_14902);
or UO_1696 (O_1696,N_14939,N_14965);
nand UO_1697 (O_1697,N_14928,N_14954);
nor UO_1698 (O_1698,N_14967,N_14901);
or UO_1699 (O_1699,N_14941,N_14935);
and UO_1700 (O_1700,N_14916,N_14886);
or UO_1701 (O_1701,N_14994,N_14942);
nand UO_1702 (O_1702,N_14972,N_14882);
and UO_1703 (O_1703,N_14896,N_14987);
or UO_1704 (O_1704,N_14910,N_14907);
nor UO_1705 (O_1705,N_14888,N_14980);
nand UO_1706 (O_1706,N_14968,N_14880);
nor UO_1707 (O_1707,N_14896,N_14942);
xnor UO_1708 (O_1708,N_14979,N_14996);
nor UO_1709 (O_1709,N_14876,N_14956);
nor UO_1710 (O_1710,N_14923,N_14987);
nand UO_1711 (O_1711,N_14958,N_14962);
or UO_1712 (O_1712,N_14953,N_14979);
nor UO_1713 (O_1713,N_14900,N_14896);
xnor UO_1714 (O_1714,N_14996,N_14894);
and UO_1715 (O_1715,N_14932,N_14958);
nand UO_1716 (O_1716,N_14953,N_14909);
xor UO_1717 (O_1717,N_14900,N_14992);
or UO_1718 (O_1718,N_14978,N_14918);
nand UO_1719 (O_1719,N_14983,N_14980);
xnor UO_1720 (O_1720,N_14889,N_14990);
or UO_1721 (O_1721,N_14945,N_14954);
nand UO_1722 (O_1722,N_14997,N_14930);
xor UO_1723 (O_1723,N_14949,N_14926);
nor UO_1724 (O_1724,N_14964,N_14932);
nor UO_1725 (O_1725,N_14918,N_14908);
nand UO_1726 (O_1726,N_14945,N_14962);
nand UO_1727 (O_1727,N_14986,N_14980);
xor UO_1728 (O_1728,N_14989,N_14991);
and UO_1729 (O_1729,N_14919,N_14934);
nand UO_1730 (O_1730,N_14970,N_14935);
nor UO_1731 (O_1731,N_14907,N_14885);
nand UO_1732 (O_1732,N_14962,N_14948);
and UO_1733 (O_1733,N_14879,N_14969);
or UO_1734 (O_1734,N_14951,N_14928);
or UO_1735 (O_1735,N_14912,N_14908);
nor UO_1736 (O_1736,N_14923,N_14985);
nand UO_1737 (O_1737,N_14984,N_14944);
and UO_1738 (O_1738,N_14947,N_14951);
or UO_1739 (O_1739,N_14983,N_14897);
nand UO_1740 (O_1740,N_14973,N_14921);
or UO_1741 (O_1741,N_14938,N_14926);
nor UO_1742 (O_1742,N_14991,N_14892);
xor UO_1743 (O_1743,N_14878,N_14893);
and UO_1744 (O_1744,N_14914,N_14964);
or UO_1745 (O_1745,N_14968,N_14995);
or UO_1746 (O_1746,N_14930,N_14966);
or UO_1747 (O_1747,N_14934,N_14925);
xor UO_1748 (O_1748,N_14978,N_14924);
nor UO_1749 (O_1749,N_14908,N_14959);
or UO_1750 (O_1750,N_14917,N_14936);
or UO_1751 (O_1751,N_14933,N_14923);
nor UO_1752 (O_1752,N_14997,N_14975);
or UO_1753 (O_1753,N_14953,N_14995);
or UO_1754 (O_1754,N_14916,N_14979);
and UO_1755 (O_1755,N_14900,N_14907);
xnor UO_1756 (O_1756,N_14919,N_14993);
xnor UO_1757 (O_1757,N_14888,N_14972);
nor UO_1758 (O_1758,N_14898,N_14988);
or UO_1759 (O_1759,N_14907,N_14994);
and UO_1760 (O_1760,N_14939,N_14988);
nor UO_1761 (O_1761,N_14932,N_14960);
nand UO_1762 (O_1762,N_14946,N_14956);
or UO_1763 (O_1763,N_14899,N_14974);
and UO_1764 (O_1764,N_14953,N_14977);
or UO_1765 (O_1765,N_14910,N_14875);
xnor UO_1766 (O_1766,N_14927,N_14876);
nor UO_1767 (O_1767,N_14907,N_14965);
nor UO_1768 (O_1768,N_14907,N_14934);
xor UO_1769 (O_1769,N_14984,N_14935);
nor UO_1770 (O_1770,N_14975,N_14932);
nand UO_1771 (O_1771,N_14995,N_14954);
xor UO_1772 (O_1772,N_14971,N_14967);
or UO_1773 (O_1773,N_14914,N_14878);
xnor UO_1774 (O_1774,N_14957,N_14914);
nand UO_1775 (O_1775,N_14990,N_14928);
and UO_1776 (O_1776,N_14957,N_14920);
nor UO_1777 (O_1777,N_14943,N_14982);
and UO_1778 (O_1778,N_14920,N_14958);
or UO_1779 (O_1779,N_14997,N_14876);
and UO_1780 (O_1780,N_14986,N_14936);
or UO_1781 (O_1781,N_14890,N_14938);
and UO_1782 (O_1782,N_14996,N_14985);
nand UO_1783 (O_1783,N_14984,N_14886);
xor UO_1784 (O_1784,N_14990,N_14921);
and UO_1785 (O_1785,N_14936,N_14963);
and UO_1786 (O_1786,N_14943,N_14996);
xor UO_1787 (O_1787,N_14953,N_14960);
nor UO_1788 (O_1788,N_14943,N_14989);
and UO_1789 (O_1789,N_14898,N_14975);
nand UO_1790 (O_1790,N_14881,N_14903);
nor UO_1791 (O_1791,N_14995,N_14960);
xor UO_1792 (O_1792,N_14961,N_14985);
and UO_1793 (O_1793,N_14963,N_14913);
nor UO_1794 (O_1794,N_14936,N_14908);
nor UO_1795 (O_1795,N_14970,N_14897);
or UO_1796 (O_1796,N_14933,N_14937);
xnor UO_1797 (O_1797,N_14897,N_14898);
nor UO_1798 (O_1798,N_14923,N_14897);
nand UO_1799 (O_1799,N_14980,N_14948);
or UO_1800 (O_1800,N_14990,N_14967);
or UO_1801 (O_1801,N_14896,N_14913);
or UO_1802 (O_1802,N_14898,N_14889);
and UO_1803 (O_1803,N_14994,N_14902);
and UO_1804 (O_1804,N_14995,N_14982);
or UO_1805 (O_1805,N_14920,N_14938);
or UO_1806 (O_1806,N_14878,N_14929);
nor UO_1807 (O_1807,N_14984,N_14888);
nand UO_1808 (O_1808,N_14964,N_14992);
nor UO_1809 (O_1809,N_14936,N_14876);
or UO_1810 (O_1810,N_14931,N_14995);
or UO_1811 (O_1811,N_14888,N_14998);
nand UO_1812 (O_1812,N_14972,N_14879);
nor UO_1813 (O_1813,N_14885,N_14982);
and UO_1814 (O_1814,N_14987,N_14994);
or UO_1815 (O_1815,N_14942,N_14968);
xor UO_1816 (O_1816,N_14931,N_14961);
or UO_1817 (O_1817,N_14940,N_14913);
nand UO_1818 (O_1818,N_14970,N_14939);
xor UO_1819 (O_1819,N_14927,N_14890);
nor UO_1820 (O_1820,N_14879,N_14911);
or UO_1821 (O_1821,N_14988,N_14896);
xor UO_1822 (O_1822,N_14916,N_14876);
and UO_1823 (O_1823,N_14881,N_14905);
xor UO_1824 (O_1824,N_14947,N_14958);
nand UO_1825 (O_1825,N_14875,N_14997);
or UO_1826 (O_1826,N_14946,N_14881);
nand UO_1827 (O_1827,N_14983,N_14938);
xnor UO_1828 (O_1828,N_14896,N_14980);
or UO_1829 (O_1829,N_14957,N_14905);
nand UO_1830 (O_1830,N_14999,N_14994);
nor UO_1831 (O_1831,N_14969,N_14875);
and UO_1832 (O_1832,N_14992,N_14939);
xnor UO_1833 (O_1833,N_14960,N_14941);
or UO_1834 (O_1834,N_14927,N_14907);
or UO_1835 (O_1835,N_14971,N_14918);
nand UO_1836 (O_1836,N_14911,N_14991);
or UO_1837 (O_1837,N_14902,N_14999);
or UO_1838 (O_1838,N_14912,N_14990);
nor UO_1839 (O_1839,N_14898,N_14900);
and UO_1840 (O_1840,N_14898,N_14890);
nand UO_1841 (O_1841,N_14919,N_14886);
or UO_1842 (O_1842,N_14879,N_14890);
and UO_1843 (O_1843,N_14941,N_14916);
nand UO_1844 (O_1844,N_14899,N_14883);
and UO_1845 (O_1845,N_14998,N_14979);
xor UO_1846 (O_1846,N_14937,N_14887);
or UO_1847 (O_1847,N_14894,N_14892);
nand UO_1848 (O_1848,N_14882,N_14913);
nor UO_1849 (O_1849,N_14957,N_14932);
nor UO_1850 (O_1850,N_14909,N_14946);
xor UO_1851 (O_1851,N_14973,N_14907);
nor UO_1852 (O_1852,N_14939,N_14882);
nor UO_1853 (O_1853,N_14973,N_14984);
and UO_1854 (O_1854,N_14936,N_14949);
and UO_1855 (O_1855,N_14962,N_14991);
or UO_1856 (O_1856,N_14948,N_14917);
nand UO_1857 (O_1857,N_14889,N_14922);
nor UO_1858 (O_1858,N_14932,N_14966);
nand UO_1859 (O_1859,N_14978,N_14995);
and UO_1860 (O_1860,N_14971,N_14878);
nand UO_1861 (O_1861,N_14891,N_14977);
xor UO_1862 (O_1862,N_14931,N_14925);
nand UO_1863 (O_1863,N_14904,N_14921);
and UO_1864 (O_1864,N_14923,N_14942);
xnor UO_1865 (O_1865,N_14947,N_14881);
xor UO_1866 (O_1866,N_14924,N_14933);
and UO_1867 (O_1867,N_14927,N_14921);
xor UO_1868 (O_1868,N_14963,N_14975);
nand UO_1869 (O_1869,N_14895,N_14920);
xor UO_1870 (O_1870,N_14890,N_14990);
or UO_1871 (O_1871,N_14954,N_14906);
xor UO_1872 (O_1872,N_14966,N_14996);
nand UO_1873 (O_1873,N_14904,N_14959);
nor UO_1874 (O_1874,N_14925,N_14980);
and UO_1875 (O_1875,N_14983,N_14890);
nor UO_1876 (O_1876,N_14932,N_14875);
and UO_1877 (O_1877,N_14991,N_14948);
and UO_1878 (O_1878,N_14893,N_14946);
xor UO_1879 (O_1879,N_14952,N_14902);
nand UO_1880 (O_1880,N_14991,N_14980);
nand UO_1881 (O_1881,N_14898,N_14949);
xnor UO_1882 (O_1882,N_14951,N_14963);
or UO_1883 (O_1883,N_14914,N_14944);
and UO_1884 (O_1884,N_14888,N_14903);
and UO_1885 (O_1885,N_14919,N_14947);
nand UO_1886 (O_1886,N_14955,N_14906);
or UO_1887 (O_1887,N_14921,N_14950);
or UO_1888 (O_1888,N_14881,N_14942);
nor UO_1889 (O_1889,N_14998,N_14960);
nand UO_1890 (O_1890,N_14928,N_14965);
nand UO_1891 (O_1891,N_14890,N_14948);
nand UO_1892 (O_1892,N_14886,N_14914);
and UO_1893 (O_1893,N_14969,N_14992);
xor UO_1894 (O_1894,N_14938,N_14949);
and UO_1895 (O_1895,N_14993,N_14988);
and UO_1896 (O_1896,N_14959,N_14887);
and UO_1897 (O_1897,N_14952,N_14913);
and UO_1898 (O_1898,N_14999,N_14995);
xnor UO_1899 (O_1899,N_14917,N_14920);
xnor UO_1900 (O_1900,N_14885,N_14881);
and UO_1901 (O_1901,N_14893,N_14959);
and UO_1902 (O_1902,N_14893,N_14978);
xor UO_1903 (O_1903,N_14877,N_14882);
and UO_1904 (O_1904,N_14938,N_14986);
and UO_1905 (O_1905,N_14878,N_14940);
and UO_1906 (O_1906,N_14929,N_14944);
xor UO_1907 (O_1907,N_14897,N_14894);
or UO_1908 (O_1908,N_14890,N_14980);
and UO_1909 (O_1909,N_14927,N_14915);
and UO_1910 (O_1910,N_14947,N_14920);
or UO_1911 (O_1911,N_14987,N_14986);
nand UO_1912 (O_1912,N_14876,N_14944);
and UO_1913 (O_1913,N_14965,N_14996);
and UO_1914 (O_1914,N_14992,N_14883);
nand UO_1915 (O_1915,N_14996,N_14997);
nor UO_1916 (O_1916,N_14999,N_14924);
nand UO_1917 (O_1917,N_14906,N_14920);
nand UO_1918 (O_1918,N_14981,N_14977);
or UO_1919 (O_1919,N_14997,N_14959);
nand UO_1920 (O_1920,N_14976,N_14937);
xnor UO_1921 (O_1921,N_14944,N_14879);
xnor UO_1922 (O_1922,N_14995,N_14967);
nor UO_1923 (O_1923,N_14932,N_14921);
nand UO_1924 (O_1924,N_14944,N_14926);
xor UO_1925 (O_1925,N_14928,N_14903);
or UO_1926 (O_1926,N_14994,N_14936);
nand UO_1927 (O_1927,N_14998,N_14999);
and UO_1928 (O_1928,N_14984,N_14884);
xnor UO_1929 (O_1929,N_14934,N_14954);
nand UO_1930 (O_1930,N_14960,N_14912);
or UO_1931 (O_1931,N_14910,N_14974);
and UO_1932 (O_1932,N_14994,N_14961);
xnor UO_1933 (O_1933,N_14951,N_14962);
and UO_1934 (O_1934,N_14986,N_14933);
or UO_1935 (O_1935,N_14909,N_14952);
nor UO_1936 (O_1936,N_14923,N_14956);
nand UO_1937 (O_1937,N_14952,N_14900);
nand UO_1938 (O_1938,N_14950,N_14883);
xor UO_1939 (O_1939,N_14885,N_14906);
nor UO_1940 (O_1940,N_14979,N_14896);
nor UO_1941 (O_1941,N_14964,N_14999);
xor UO_1942 (O_1942,N_14950,N_14979);
xnor UO_1943 (O_1943,N_14951,N_14892);
nor UO_1944 (O_1944,N_14939,N_14931);
and UO_1945 (O_1945,N_14945,N_14988);
or UO_1946 (O_1946,N_14995,N_14875);
nor UO_1947 (O_1947,N_14909,N_14943);
xnor UO_1948 (O_1948,N_14939,N_14944);
and UO_1949 (O_1949,N_14951,N_14899);
nor UO_1950 (O_1950,N_14956,N_14932);
and UO_1951 (O_1951,N_14964,N_14951);
nor UO_1952 (O_1952,N_14981,N_14966);
xnor UO_1953 (O_1953,N_14902,N_14954);
and UO_1954 (O_1954,N_14943,N_14957);
or UO_1955 (O_1955,N_14928,N_14922);
xnor UO_1956 (O_1956,N_14951,N_14999);
xor UO_1957 (O_1957,N_14876,N_14948);
or UO_1958 (O_1958,N_14971,N_14985);
nor UO_1959 (O_1959,N_14909,N_14919);
nand UO_1960 (O_1960,N_14941,N_14898);
xor UO_1961 (O_1961,N_14909,N_14883);
nand UO_1962 (O_1962,N_14947,N_14890);
or UO_1963 (O_1963,N_14893,N_14924);
xnor UO_1964 (O_1964,N_14960,N_14886);
or UO_1965 (O_1965,N_14890,N_14905);
nand UO_1966 (O_1966,N_14979,N_14918);
xor UO_1967 (O_1967,N_14927,N_14984);
and UO_1968 (O_1968,N_14906,N_14944);
nand UO_1969 (O_1969,N_14907,N_14913);
xor UO_1970 (O_1970,N_14900,N_14986);
or UO_1971 (O_1971,N_14975,N_14879);
xnor UO_1972 (O_1972,N_14951,N_14941);
nor UO_1973 (O_1973,N_14876,N_14992);
nor UO_1974 (O_1974,N_14971,N_14944);
and UO_1975 (O_1975,N_14948,N_14993);
xnor UO_1976 (O_1976,N_14981,N_14919);
or UO_1977 (O_1977,N_14894,N_14985);
xnor UO_1978 (O_1978,N_14901,N_14966);
nor UO_1979 (O_1979,N_14963,N_14877);
nor UO_1980 (O_1980,N_14877,N_14929);
or UO_1981 (O_1981,N_14965,N_14975);
nand UO_1982 (O_1982,N_14940,N_14945);
nor UO_1983 (O_1983,N_14900,N_14989);
xnor UO_1984 (O_1984,N_14884,N_14912);
xor UO_1985 (O_1985,N_14973,N_14931);
nor UO_1986 (O_1986,N_14954,N_14889);
or UO_1987 (O_1987,N_14945,N_14901);
and UO_1988 (O_1988,N_14966,N_14918);
or UO_1989 (O_1989,N_14942,N_14996);
nand UO_1990 (O_1990,N_14909,N_14961);
and UO_1991 (O_1991,N_14980,N_14912);
or UO_1992 (O_1992,N_14906,N_14933);
xor UO_1993 (O_1993,N_14946,N_14951);
nor UO_1994 (O_1994,N_14966,N_14900);
nand UO_1995 (O_1995,N_14919,N_14966);
nor UO_1996 (O_1996,N_14941,N_14903);
nor UO_1997 (O_1997,N_14917,N_14959);
nor UO_1998 (O_1998,N_14943,N_14947);
and UO_1999 (O_1999,N_14959,N_14947);
endmodule